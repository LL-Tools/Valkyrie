

module b17_C_gen_AntiSAT_k_128_6 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput_f0, keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, 
        keyinput_f5, keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, 
        keyinput_f10, keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, 
        keyinput_f15, keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, 
        keyinput_f20, keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, 
        keyinput_f25, keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, 
        keyinput_f30, keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, 
        keyinput_f35, keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, 
        keyinput_f40, keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, 
        keyinput_f45, keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, 
        keyinput_f50, keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, 
        keyinput_f55, keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, 
        keyinput_f60, keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, 
        keyinput_g1, keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, 
        keyinput_g6, keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, 
        keyinput_g11, keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, 
        keyinput_g16, keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, 
        keyinput_g21, keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, 
        keyinput_g26, keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, 
        keyinput_g31, keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, 
        keyinput_g36, keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, 
        keyinput_g41, keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, 
        keyinput_g46, keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, 
        keyinput_g51, keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, 
        keyinput_g56, keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, 
        keyinput_g61, keyinput_g62, keyinput_g63, U355, U356, U357, U358, U359, 
        U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, 
        U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, 
        U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, 
        U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, 
        U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, 
        U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, 
        U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, 
        U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9653, n9654, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13686, n13687, n13688, n13689, n13690, n13691, n13692,
         n13693, n13694, n13695, n13696, n13697, n13698, n13699, n13700,
         n13701, n13702, n13703, n13704, n13705, n13706, n13707, n13708,
         n13709, n13710, n13711, n13712, n13713, n13714, n13715, n13716,
         n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
         n13725, n13726, n13727, n13728, n13729, n13730, n13731, n13732,
         n13733, n13734, n13735, n13736, n13737, n13738, n13739, n13740,
         n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
         n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756,
         n13757, n13758, n13759, n13760, n13761, n13762, n13763, n13764,
         n13765, n13766, n13767, n13768, n13769, n13770, n13771, n13772,
         n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780,
         n13781, n13782, n13783, n13784, n13785, n13786, n13787, n13788,
         n13789, n13790, n13791, n13792, n13793, n13794, n13795, n13796,
         n13797, n13798, n13799, n13800, n13801, n13802, n13803, n13804,
         n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812,
         n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
         n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
         n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836,
         n13837, n13838, n13839, n13840, n13841, n13842, n13843, n13844,
         n13845, n13846, n13847, n13848, n13849, n13850, n13851, n13852,
         n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
         n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868,
         n13869, n13870, n13871, n13872, n13873, n13874, n13875, n13876,
         n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884,
         n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
         n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900,
         n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908,
         n13909, n13910, n13911, n13912, n13913, n13914, n13915, n13916,
         n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
         n13925, n13926, n13927, n13928, n13929, n13930, n13931, n13932,
         n13933, n13934, n13935, n13936, n13937, n13938, n13939, n13940,
         n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948,
         n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956,
         n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126,
         n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
         n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
         n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
         n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
         n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174,
         n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
         n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
         n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198,
         n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
         n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214,
         n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222,
         n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
         n21231, n21232, n21233;

  NAND2_X1 U11097 ( .A1(n18024), .A2(n17929), .ZN(n18170) );
  AND2_X1 U11098 ( .A1(n14166), .A2(n14737), .ZN(n20338) );
  AND2_X1 U11099 ( .A1(n13230), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13229) );
  NOR2_X1 U11100 ( .A1(n15750), .A2(n15884), .ZN(n15751) );
  NOR2_X1 U11101 ( .A1(n16035), .A2(n16042), .ZN(n16002) );
  NOR2_X1 U11102 ( .A1(n15535), .A2(n10781), .ZN(n15714) );
  NOR2_X1 U11103 ( .A1(n17782), .A2(n17604), .ZN(n17603) );
  INV_X2 U11104 ( .A(n18240), .ZN(n18966) );
  AOI21_X1 U11105 ( .B1(n15233), .B2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10075), .ZN(n10074) );
  AND2_X1 U11107 ( .A1(n15529), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15531) );
  INV_X2 U11108 ( .A(n18080), .ZN(n18066) );
  NAND2_X1 U11109 ( .A1(n12815), .A2(n12814), .ZN(n13741) );
  BUF_X1 U11110 ( .A(n16274), .Z(n9725) );
  NOR2_X1 U11111 ( .A1(n12055), .A2(n13954), .ZN(n12091) );
  OR2_X1 U11112 ( .A1(n13915), .A2(n13914), .ZN(n9895) );
  OR2_X1 U11113 ( .A1(n10334), .A2(n10352), .ZN(n10483) );
  AND2_X1 U11114 ( .A1(n9734), .A2(n10340), .ZN(n10114) );
  OR2_X1 U11115 ( .A1(n14391), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11971) );
  NAND2_X1 U11116 ( .A1(n11945), .A2(n13296), .ZN(n11972) );
  INV_X4 U11117 ( .A(n17511), .ZN(n16175) );
  XNOR2_X1 U11118 ( .A(n13612), .B(n11406), .ZN(n13627) );
  AND2_X1 U11119 ( .A1(n13609), .A2(n13610), .ZN(n13612) );
  BUF_X2 U11120 ( .A(n10961), .Z(n17476) );
  CLKBUF_X1 U11121 ( .A(n10981), .Z(n17339) );
  CLKBUF_X2 U11122 ( .A(n11823), .Z(n12508) );
  NAND2_X1 U11123 ( .A1(n11389), .A2(n9908), .ZN(n11632) );
  AND3_X1 U11124 ( .A1(n9684), .A2(n10248), .A3(n20195), .ZN(n11602) );
  INV_X2 U11125 ( .A(n17455), .ZN(n11129) );
  INV_X1 U11126 ( .A(n12896), .ZN(n12960) );
  INV_X2 U11127 ( .A(n10109), .ZN(n17420) );
  AND2_X1 U11128 ( .A1(n14039), .A2(n10371), .ZN(n10385) );
  AND2_X1 U11129 ( .A1(n12976), .A2(n10370), .ZN(n10396) );
  AND2_X1 U11130 ( .A1(n14039), .A2(n12976), .ZN(n10384) );
  CLKBUF_X2 U11131 ( .A(n11774), .Z(n12396) );
  INV_X1 U11132 ( .A(n10948), .ZN(n17403) );
  INV_X1 U11133 ( .A(n9752), .ZN(n9671) );
  INV_X1 U11134 ( .A(n16118), .ZN(n17457) );
  AND2_X1 U11135 ( .A1(n9686), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12907) );
  AND2_X1 U11136 ( .A1(n13150), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12906) );
  INV_X2 U11137 ( .A(n10949), .ZN(n17495) );
  AND2_X1 U11138 ( .A1(n10194), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12904) );
  CLKBUF_X2 U11139 ( .A(n11804), .Z(n12384) );
  AND2_X1 U11140 ( .A1(n10188), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12965) );
  AND2_X1 U11141 ( .A1(n10372), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12964) );
  INV_X1 U11142 ( .A(n13128), .ZN(n13162) );
  NOR2_X1 U11143 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12976) );
  INV_X1 U11144 ( .A(n13134), .ZN(n13128) );
  NOR2_X1 U11145 ( .A1(n9997), .A2(n10935), .ZN(n18984) );
  OR2_X2 U11146 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10933), .ZN(
        n17472) );
  NAND2_X2 U11148 ( .A1(n10221), .A2(n10454), .ZN(n11336) );
  INV_X1 U11149 ( .A(n11336), .ZN(n10646) );
  NAND4_X2 U11150 ( .A1(n11786), .A2(n11785), .A3(n11784), .A4(n11783), .ZN(
        n12589) );
  INV_X2 U11151 ( .A(n13115), .ZN(n14000) );
  AND2_X2 U11152 ( .A1(n10370), .A2(n14006), .ZN(n10194) );
  INV_X1 U11154 ( .A(n20014), .ZN(n9653) );
  NOR2_X1 U11155 ( .A1(n9654), .A2(n16035), .ZN(n13230) );
  NAND2_X1 U11156 ( .A1(n9806), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9654) );
  NAND2_X1 U11157 ( .A1(n10113), .A2(n10346), .ZN(n20018) );
  AOI22_X2 U11158 ( .A1(n11077), .A2(n11076), .B1(n11075), .B2(n11074), .ZN(
        n11700) );
  OR2_X2 U11159 ( .A1(n18102), .A2(n18423), .ZN(n11058) );
  NAND2_X2 U11160 ( .A1(n14157), .A2(n14159), .ZN(n14158) );
  NOR2_X4 U11161 ( .A1(n13925), .A2(n16021), .ZN(n14157) );
  NAND2_X2 U11162 ( .A1(n13667), .A2(n13666), .ZN(n13722) );
  NOR2_X2 U11163 ( .A1(n15632), .A2(n15633), .ZN(n15536) );
  NOR2_X2 U11164 ( .A1(n14158), .A2(n9896), .ZN(n14433) );
  NOR2_X2 U11165 ( .A1(n10378), .A2(n10377), .ZN(n11395) );
  NAND2_X2 U11166 ( .A1(n14708), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9849) );
  OAI22_X2 U11167 ( .A1(n16757), .A2(n14147), .B1(n21177), .B2(n14146), .ZN(
        n20901) );
  NAND2_X2 U11168 ( .A1(n16364), .A2(n14104), .ZN(n14146) );
  NAND2_X2 U11169 ( .A1(n16364), .A2(n14699), .ZN(n14147) );
  INV_X1 U11171 ( .A(n21233), .ZN(n9656) );
  NOR2_X2 U11173 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11744) );
  OR2_X1 U11174 ( .A1(n11972), .A2(n11974), .ZN(n11975) );
  AND2_X2 U11175 ( .A1(n11744), .A2(n13857), .ZN(n12542) );
  AND4_X1 U11176 ( .A1(n11756), .A2(n11755), .A3(n11754), .A4(n11753), .ZN(
        n10088) );
  AND2_X1 U11177 ( .A1(n11971), .A2(n11970), .ZN(n13237) );
  INV_X1 U11178 ( .A(n12904), .ZN(n12955) );
  NAND2_X1 U11179 ( .A1(n9737), .A2(n10359), .ZN(n12963) );
  OAI21_X1 U11180 ( .B1(n10661), .B2(n10290), .A(n10289), .ZN(n10291) );
  INV_X1 U11181 ( .A(n10352), .ZN(n10346) );
  NAND2_X1 U11182 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n10935), .ZN(
        n10927) );
  NOR2_X1 U11183 ( .A1(n17567), .A2(n18542), .ZN(n11234) );
  INV_X1 U11184 ( .A(n12091), .ZN(n12079) );
  OR2_X1 U11185 ( .A1(n15559), .A2(n10017), .ZN(n10020) );
  OAI21_X1 U11187 ( .B1(n10808), .B2(n14818), .A(n19414), .ZN(n10809) );
  AND2_X1 U11188 ( .A1(n10368), .A2(n10371), .ZN(n10383) );
  AND2_X2 U11189 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10637) );
  INV_X2 U11190 ( .A(n10978), .ZN(n17514) );
  INV_X1 U11191 ( .A(n10948), .ZN(n9667) );
  NAND2_X1 U11192 ( .A1(n9997), .A2(n9998), .ZN(n10931) );
  NAND2_X1 U11193 ( .A1(n14133), .A2(n11889), .ZN(n13658) );
  INV_X1 U11194 ( .A(n9738), .ZN(n9674) );
  AOI21_X1 U11195 ( .B1(n10074), .B2(n10072), .A(n10071), .ZN(n10070) );
  NAND2_X1 U11196 ( .A1(n11986), .A2(n11985), .ZN(n12036) );
  INV_X1 U11197 ( .A(n11889), .ZN(n11941) );
  INV_X1 U11198 ( .A(n19551), .ZN(n14815) );
  AOI21_X1 U11199 ( .B1(n12817), .B2(n13745), .A(n12816), .ZN(n12818) );
  INV_X1 U11200 ( .A(n10454), .ZN(n9684) );
  XNOR2_X1 U11201 ( .A(n10311), .B(n10310), .ZN(n10312) );
  NAND2_X1 U11202 ( .A1(n17765), .A2(n11237), .ZN(n16855) );
  INV_X1 U11203 ( .A(n9752), .ZN(n9670) );
  NAND2_X1 U11204 ( .A1(n10115), .A2(n11795), .ZN(n11877) );
  INV_X1 U11205 ( .A(n15968), .ZN(n14598) );
  OR2_X1 U11206 ( .A1(n9709), .A2(n9710), .ZN(n17588) );
  INV_X2 U11207 ( .A(n10946), .ZN(n17421) );
  AOI221_X1 U11208 ( .B1(n17901), .B2(n18238), .C1(n17901), .C2(n9675), .A(
        n17935), .ZN(n17902) );
  INV_X1 U11209 ( .A(n20338), .ZN(n20306) );
  INV_X1 U11210 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11741) );
  AOI211_X1 U11211 ( .C1(n17421), .C2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n10958), .B(n10957), .ZN(n17704) );
  INV_X1 U11212 ( .A(n18170), .ZN(n18160) );
  INV_X1 U11213 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9832) );
  INV_X1 U11214 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14006) );
  NAND2_X2 U11215 ( .A1(n11757), .A2(n10088), .ZN(n13678) );
  INV_X1 U11216 ( .A(n13678), .ZN(n12770) );
  NAND3_X2 U11217 ( .A1(n9832), .A2(n10118), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13007) );
  NOR2_X2 U11218 ( .A1(n17789), .A2(n17588), .ZN(n17582) );
  NOR2_X2 U11219 ( .A1(n18112), .A2(n18113), .ZN(n18082) );
  AND2_X4 U11220 ( .A1(n11740), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11750) );
  AND2_X2 U11221 ( .A1(n15708), .A2(n15711), .ZN(n10096) );
  OR2_X2 U11222 ( .A1(n13997), .A2(n20218), .ZN(n9657) );
  INV_X1 U11223 ( .A(n10747), .ZN(n9658) );
  INV_X1 U11224 ( .A(n9657), .ZN(n9659) );
  NOR2_X2 U11226 ( .A1(n17965), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17964) );
  BUF_X1 U11227 ( .A(n14856), .Z(n9660) );
  NOR2_X2 U11228 ( .A1(n10862), .A2(n10861), .ZN(n10863) );
  NOR2_X2 U11229 ( .A1(n12057), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11743) );
  AND2_X4 U11230 ( .A1(n11752), .A2(n13875), .ZN(n11860) );
  AND2_X2 U11231 ( .A1(n10066), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11752) );
  AND2_X1 U11233 ( .A1(n13875), .A2(n13858), .ZN(n9661) );
  AND2_X1 U11234 ( .A1(n13875), .A2(n13858), .ZN(n11823) );
  NAND2_X2 U11235 ( .A1(n13557), .A2(n11887), .ZN(n13692) );
  AND2_X2 U11236 ( .A1(n11744), .A2(n13857), .ZN(n9662) );
  AND2_X4 U11239 ( .A1(n13559), .A2(n13858), .ZN(n11824) );
  INV_X2 U11240 ( .A(n13106), .ZN(n9665) );
  INV_X1 U11241 ( .A(n13106), .ZN(n9666) );
  NAND2_X4 U11242 ( .A1(n10637), .A2(n10016), .ZN(n13106) );
  INV_X2 U11243 ( .A(n11350), .ZN(n19543) );
  INV_X2 U11244 ( .A(n10219), .ZN(n11350) );
  AND2_X4 U11246 ( .A1(n11750), .A2(n13875), .ZN(n11804) );
  NAND2_X2 U11247 ( .A1(n15709), .A2(n10096), .ZN(n15731) );
  AND2_X1 U11248 ( .A1(n10370), .A2(n14006), .ZN(n9668) );
  NOR2_X2 U11249 ( .A1(n15600), .A2(n15601), .ZN(n13004) );
  NAND2_X2 U11250 ( .A1(n10599), .A2(n9760), .ZN(n10601) );
  INV_X4 U11251 ( .A(n16111), .ZN(n17512) );
  AND2_X4 U11252 ( .A1(n10117), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10368) );
  AND2_X4 U11253 ( .A1(n11752), .A2(n11751), .ZN(n11774) );
  AND2_X2 U11254 ( .A1(n11742), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11751) );
  XNOR2_X1 U11255 ( .A(n11701), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n17205) );
  NAND2_X1 U11256 ( .A1(n11875), .A2(n9852), .ZN(n9669) );
  INV_X1 U11257 ( .A(n9671), .ZN(n9672) );
  OR3_X1 U11258 ( .A1(n18989), .A2(n10936), .A3(n10935), .ZN(n9752) );
  NOR2_X2 U11259 ( .A1(n14893), .A2(n14895), .ZN(n14881) );
  XNOR2_X2 U11260 ( .A(n9909), .B(n10660), .ZN(n12808) );
  NAND2_X2 U11261 ( .A1(n9831), .A2(n10297), .ZN(n9909) );
  INV_X1 U11262 ( .A(n9738), .ZN(n9673) );
  INV_X2 U11263 ( .A(n9738), .ZN(n15449) );
  CLKBUF_X3 U11264 ( .A(n17973), .Z(n9675) );
  NAND2_X1 U11265 ( .A1(n15230), .A2(n10072), .ZN(n9845) );
  AND2_X1 U11266 ( .A1(n15576), .A2(n13053), .ZN(n13077) );
  AOI21_X1 U11267 ( .B1(n15232), .B2(n15244), .A(n13312), .ZN(n15233) );
  OR2_X1 U11268 ( .A1(n17864), .A2(n11067), .ZN(n11069) );
  AOI221_X1 U11269 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17946), 
        .C1(n17936), .C2(n17957), .A(n17935), .ZN(n17937) );
  AOI22_X1 U11270 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14838), .B1(n15698), 
        .B2(n20218), .ZN(n14305) );
  OAI21_X1 U11271 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19179), .A(n16856), 
        .ZN(n18176) );
  NAND2_X1 U11273 ( .A1(n10114), .A2(n10346), .ZN(n10479) );
  NAND2_X1 U11274 ( .A1(n10114), .A2(n10352), .ZN(n10480) );
  NOR2_X1 U11275 ( .A1(n14500), .A2(n15088), .ZN(n20917) );
  NOR2_X1 U11276 ( .A1(n14500), .A2(n15103), .ZN(n20899) );
  NOR2_X1 U11277 ( .A1(n14500), .A2(n15093), .ZN(n20911) );
  NOR2_X1 U11278 ( .A1(n14500), .A2(n15098), .ZN(n20905) );
  NOR2_X1 U11279 ( .A1(n15076), .A2(n14500), .ZN(n20932) );
  NOR2_X1 U11280 ( .A1(n14500), .A2(n15117), .ZN(n20882) );
  NOR2_X1 U11281 ( .A1(n14500), .A2(n15108), .ZN(n20893) );
  AND2_X1 U11282 ( .A1(n15527), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15529) );
  OAI21_X1 U11283 ( .B1(n16277), .B2(n16276), .A(n19180), .ZN(n17720) );
  NOR2_X1 U11285 ( .A1(n19186), .A2(n17820), .ZN(n17821) );
  NOR2_X1 U11286 ( .A1(n10824), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n19366) );
  NOR2_X1 U11287 ( .A1(n10790), .A2(n10783), .ZN(n10782) );
  INV_X1 U11288 ( .A(n18548), .ZN(n17691) );
  CLKBUF_X1 U11289 ( .A(n10256), .Z(n13406) );
  NAND2_X1 U11290 ( .A1(n14185), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15513) );
  INV_X2 U11291 ( .A(n11354), .ZN(n10221) );
  NOR2_X1 U11292 ( .A1(n10248), .A2(n10454), .ZN(n11389) );
  BUF_X1 U11293 ( .A(n10236), .Z(n13746) );
  NOR2_X2 U11294 ( .A1(n14183), .A2(n19381), .ZN(n14185) );
  NAND2_X1 U11295 ( .A1(n10129), .A2(n10130), .ZN(n10454) );
  INV_X2 U11296 ( .A(n12897), .ZN(n12961) );
  INV_X1 U11297 ( .A(n11891), .ZN(n12636) );
  NAND2_X1 U11298 ( .A1(n14184), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14183) );
  INV_X4 U11299 ( .A(n17256), .ZN(n17508) );
  BUF_X2 U11301 ( .A(n12378), .Z(n12543) );
  BUF_X2 U11302 ( .A(n11859), .Z(n12526) );
  CLKBUF_X2 U11303 ( .A(n12527), .Z(n12224) );
  AND2_X1 U11304 ( .A1(n14000), .A2(n10359), .ZN(n12905) );
  CLKBUF_X2 U11305 ( .A(n12549), .Z(n12507) );
  BUF_X2 U11306 ( .A(n11796), .Z(n9866) );
  AND2_X1 U11307 ( .A1(n13859), .A2(n13559), .ZN(n11796) );
  INV_X1 U11308 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10936) );
  NAND2_X1 U11309 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18989) );
  INV_X1 U11310 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16678) );
  NAND2_X1 U11311 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14178) );
  INV_X2 U11312 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11740) );
  NAND2_X1 U11314 ( .A1(n9927), .A2(n9926), .ZN(n11279) );
  AND2_X1 U11315 ( .A1(n9835), .A2(n9834), .ZN(n9833) );
  NAND2_X1 U11316 ( .A1(n10064), .A2(n9782), .ZN(n15810) );
  AND2_X1 U11317 ( .A1(n15845), .A2(n9934), .ZN(n9933) );
  NAND2_X1 U11318 ( .A1(n10910), .A2(n10909), .ZN(n15712) );
  AOI21_X1 U11319 ( .B1(n15704), .B2(n16700), .A(n14843), .ZN(n14844) );
  CLKBUF_X1 U11320 ( .A(n15734), .Z(n15735) );
  NOR2_X1 U11321 ( .A1(n15965), .A2(n9838), .ZN(n15986) );
  NAND2_X1 U11322 ( .A1(n13204), .A2(n16016), .ZN(n15989) );
  NAND2_X1 U11323 ( .A1(n15146), .A2(n10068), .ZN(n10069) );
  NOR2_X1 U11324 ( .A1(n15717), .A2(n14830), .ZN(n14822) );
  INV_X1 U11325 ( .A(n15717), .ZN(n15738) );
  NAND2_X1 U11326 ( .A1(n16599), .A2(n16601), .ZN(n16600) );
  NOR2_X1 U11327 ( .A1(n15996), .A2(n15985), .ZN(n15963) );
  AOI21_X1 U11328 ( .B1(n12767), .B2(n12765), .A(n12766), .ZN(n15129) );
  XNOR2_X1 U11329 ( .A(n12766), .B(n12568), .ZN(n15054) );
  NAND2_X1 U11330 ( .A1(n15997), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15996) );
  CLKBUF_X1 U11331 ( .A(n15915), .Z(n9687) );
  NOR2_X1 U11332 ( .A1(n15559), .A2(n15558), .ZN(n15557) );
  NAND2_X1 U11333 ( .A1(n16484), .A2(n16485), .ZN(n16483) );
  XNOR2_X1 U11334 ( .A(n13101), .B(n13099), .ZN(n15559) );
  NAND2_X1 U11335 ( .A1(n15567), .A2(n10095), .ZN(n13101) );
  AND2_X1 U11336 ( .A1(n9704), .A2(n9705), .ZN(n13318) );
  NAND2_X1 U11337 ( .A1(n10829), .A2(n16042), .ZN(n13198) );
  NAND2_X1 U11338 ( .A1(n16496), .A2(n16497), .ZN(n16495) );
  NAND2_X1 U11339 ( .A1(n10070), .A2(n9845), .ZN(n15194) );
  OR2_X1 U11340 ( .A1(n13077), .A2(n13078), .ZN(n10095) );
  OAI21_X1 U11341 ( .B1(n11270), .B2(n16255), .A(n18080), .ZN(n11076) );
  AOI21_X1 U11342 ( .B1(n16710), .B2(n11648), .A(n14676), .ZN(n11649) );
  AOI21_X1 U11343 ( .B1(n16493), .B2(n16710), .A(n9937), .ZN(n9936) );
  NAND2_X1 U11344 ( .A1(n10081), .A2(n10080), .ZN(n15277) );
  AND2_X1 U11345 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16052), .ZN(
        n10615) );
  NOR2_X1 U11346 ( .A1(n11686), .A2(n16200), .ZN(n11072) );
  NAND2_X1 U11347 ( .A1(n17835), .A2(n10102), .ZN(n11686) );
  NOR2_X1 U11348 ( .A1(n11663), .A2(n11728), .ZN(n11717) );
  AOI21_X1 U11349 ( .B1(n10749), .B2(n15508), .A(n10748), .ZN(n16494) );
  NAND2_X1 U11350 ( .A1(n16512), .A2(n16513), .ZN(n16511) );
  OR2_X1 U11351 ( .A1(n10606), .A2(n16638), .ZN(n10609) );
  XNOR2_X1 U11352 ( .A(n14827), .B(n14826), .ZN(n19448) );
  AND2_X1 U11353 ( .A1(n16051), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16052) );
  INV_X1 U11354 ( .A(n10058), .ZN(n10057) );
  NOR2_X1 U11355 ( .A1(n11725), .A2(n18196), .ZN(n17835) );
  XNOR2_X1 U11356 ( .A(n14835), .B(n14834), .ZN(n16481) );
  XNOR2_X1 U11357 ( .A(n10578), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16638) );
  OAI21_X1 U11358 ( .B1(n11725), .B2(n9994), .A(n9993), .ZN(n11663) );
  OR2_X1 U11359 ( .A1(n10614), .A2(n16642), .ZN(n16051) );
  AND2_X1 U11360 ( .A1(n13315), .A2(n10073), .ZN(n10072) );
  OAI21_X1 U11361 ( .B1(n11681), .B2(n11735), .A(n11680), .ZN(n11682) );
  XNOR2_X1 U11362 ( .A(n10613), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16642) );
  NAND3_X1 U11363 ( .A1(n10598), .A2(n14444), .A3(n10597), .ZN(n14449) );
  NAND2_X1 U11364 ( .A1(n10796), .A2(n14453), .ZN(n14369) );
  NOR2_X1 U11365 ( .A1(n15245), .A2(n15249), .ZN(n13315) );
  OR2_X1 U11366 ( .A1(n10576), .A2(n10577), .ZN(n10612) );
  OR2_X1 U11367 ( .A1(n10576), .A2(n10781), .ZN(n10613) );
  AND2_X1 U11368 ( .A1(n13303), .A2(n13305), .ZN(n9697) );
  NAND2_X1 U11369 ( .A1(n17275), .A2(n17551), .ZN(n17279) );
  NAND2_X1 U11370 ( .A1(n16539), .A2(n16540), .ZN(n16538) );
  NAND2_X1 U11371 ( .A1(n14378), .A2(n10589), .ZN(n16086) );
  NAND2_X1 U11372 ( .A1(n17286), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n17275) );
  NAND2_X1 U11373 ( .A1(n10075), .A2(n9805), .ZN(n10073) );
  INV_X1 U11374 ( .A(n17281), .ZN(n17286) );
  NOR3_X1 U11375 ( .A1(n18230), .A2(n11666), .A3(n17989), .ZN(n17841) );
  AND2_X1 U11376 ( .A1(n15449), .A2(n15481), .ZN(n15262) );
  INV_X1 U11377 ( .A(n17578), .ZN(n17573) );
  AOI211_X1 U11378 ( .C1(n18966), .C2(n11723), .A(n18489), .B(n16193), .ZN(
        n11724) );
  AOI211_X1 U11379 ( .C1(n18966), .C2(n18357), .A(n18377), .B(n18356), .ZN(
        n18364) );
  AOI211_X1 U11380 ( .C1(n19002), .C2(n18378), .A(n18377), .B(n18388), .ZN(
        n18379) );
  AOI211_X1 U11381 ( .C1(n18966), .C2(n18220), .A(n18489), .B(n18219), .ZN(
        n18221) );
  NAND2_X1 U11382 ( .A1(n16565), .A2(n16566), .ZN(n16564) );
  AOI22_X1 U11383 ( .A1(n18090), .A2(n18004), .B1(n18150), .B2(n18011), .ZN(
        n18078) );
  NOR2_X1 U11384 ( .A1(n17786), .A2(n17598), .ZN(n17592) );
  NAND2_X1 U11385 ( .A1(n10904), .A2(n16531), .ZN(n10907) );
  NAND2_X1 U11386 ( .A1(n9856), .A2(n9855), .ZN(n13298) );
  OR2_X1 U11387 ( .A1(n14331), .A2(n14422), .ZN(n14472) );
  NOR2_X2 U11388 ( .A1(n10898), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10904) );
  OR2_X1 U11389 ( .A1(n17784), .A2(n17597), .ZN(n17598) );
  OR2_X1 U11390 ( .A1(n17597), .A2(n17784), .ZN(n9709) );
  NOR2_X2 U11391 ( .A1(n17692), .A2(n18179), .ZN(n18090) );
  CLKBUF_X2 U11392 ( .A(n14305), .Z(n19384) );
  NOR2_X1 U11393 ( .A1(n19941), .A2(n19811), .ZN(n19867) );
  NOR2_X1 U11394 ( .A1(n10483), .A2(n12845), .ZN(n10336) );
  CLKBUF_X1 U11395 ( .A(n13246), .Z(n13949) );
  AOI22_X1 U11396 ( .A1(n18967), .A2(n18966), .B1(n18971), .B2(n11732), .ZN(
        n11664) );
  AND2_X1 U11397 ( .A1(n11055), .A2(n9995), .ZN(n18014) );
  NAND2_X1 U11398 ( .A1(n10333), .A2(n10343), .ZN(n10486) );
  AOI211_X1 U11399 ( .C1(n19002), .C2(n18186), .A(n18204), .B(n18185), .ZN(
        n18187) );
  INV_X1 U11400 ( .A(n11255), .ZN(n11055) );
  INV_X1 U11401 ( .A(n20905), .ZN(n9676) );
  NAND2_X1 U11402 ( .A1(n19186), .A2(n18451), .ZN(n18240) );
  INV_X1 U11403 ( .A(n20911), .ZN(n9677) );
  INV_X1 U11404 ( .A(n20893), .ZN(n9678) );
  INV_X1 U11405 ( .A(n20899), .ZN(n9679) );
  INV_X1 U11406 ( .A(n20882), .ZN(n9680) );
  AND2_X1 U11407 ( .A1(n13638), .A2(n12802), .ZN(n13641) );
  NOR2_X1 U11408 ( .A1(n16278), .A2(n17720), .ZN(n17718) );
  INV_X1 U11409 ( .A(n20932), .ZN(n9681) );
  INV_X1 U11410 ( .A(n20917), .ZN(n9682) );
  AND2_X1 U11411 ( .A1(n12054), .A2(n12053), .ZN(n13954) );
  AND2_X1 U11412 ( .A1(n9823), .A2(n9724), .ZN(n13398) );
  NOR2_X2 U11413 ( .A1(n18447), .A2(n19000), .ZN(n18451) );
  OR2_X1 U11414 ( .A1(n11053), .A2(n11052), .ZN(n11059) );
  NAND2_X1 U11415 ( .A1(n12794), .A2(n12793), .ZN(n12805) );
  NOR4_X1 U11416 ( .A1(n17467), .A2(n17395), .A3(n17396), .A4(n16186), .ZN(
        n17415) );
  INV_X4 U11417 ( .A(n19002), .ZN(n18992) );
  NAND2_X1 U11418 ( .A1(n12800), .A2(n12799), .ZN(n14792) );
  OR2_X2 U11419 ( .A1(n15037), .A2(n15052), .ZN(n15040) );
  AND2_X1 U11420 ( .A1(n14346), .A2(n10319), .ZN(n10340) );
  NOR2_X2 U11421 ( .A1(n19533), .A2(n19947), .ZN(n19534) );
  NOR2_X2 U11422 ( .A1(n19523), .A2(n19947), .ZN(n19524) );
  INV_X1 U11423 ( .A(n14346), .ZN(n13467) );
  INV_X1 U11424 ( .A(n18977), .ZN(n19004) );
  NAND2_X1 U11425 ( .A1(n16995), .A2(n10085), .ZN(n13362) );
  NAND2_X1 U11426 ( .A1(n15526), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15528) );
  NAND2_X2 U11427 ( .A1(n13337), .A2(n13336), .ZN(n13835) );
  NOR2_X2 U11428 ( .A1(n15525), .A2(n9812), .ZN(n15526) );
  OR2_X1 U11429 ( .A1(n14099), .A2(n11968), .ZN(n11990) );
  AND2_X2 U11430 ( .A1(n10322), .A2(n10317), .ZN(n14346) );
  XNOR2_X1 U11431 ( .A(n11965), .B(n11978), .ZN(n14099) );
  NAND2_X1 U11432 ( .A1(n15524), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15525) );
  CLKBUF_X1 U11433 ( .A(n10314), .Z(n10322) );
  NAND2_X1 U11434 ( .A1(n10766), .A2(n14815), .ZN(n10906) );
  AND2_X1 U11435 ( .A1(n9749), .A2(n13968), .ZN(n9894) );
  INV_X2 U11436 ( .A(n17205), .ZN(n17175) );
  NAND2_X1 U11437 ( .A1(n10294), .A2(n10293), .ZN(n10310) );
  XNOR2_X1 U11438 ( .A(n11046), .B(n11045), .ZN(n18131) );
  CLKBUF_X1 U11439 ( .A(n17557), .Z(n9732) );
  NAND2_X2 U11440 ( .A1(n19186), .A2(n17766), .ZN(n17831) );
  NOR2_X1 U11441 ( .A1(n16275), .A2(n9967), .ZN(n17557) );
  NOR2_X1 U11442 ( .A1(n10006), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10005) );
  NOR2_X1 U11443 ( .A1(n10000), .A2(n10002), .ZN(n9999) );
  AND2_X1 U11444 ( .A1(n18533), .A2(n11235), .ZN(n11241) );
  NOR2_X1 U11445 ( .A1(n18123), .A2(n18439), .ZN(n9991) );
  NAND2_X1 U11446 ( .A1(n13379), .A2(n11673), .ZN(n11693) );
  CLKBUF_X1 U11447 ( .A(n10274), .Z(n11345) );
  NOR3_X1 U11448 ( .A1(n11254), .A2(n11253), .A3(n18982), .ZN(n16093) );
  NOR2_X1 U11449 ( .A1(n10009), .A2(n10008), .ZN(n10007) );
  NOR2_X1 U11450 ( .A1(n11668), .A2(n17857), .ZN(n17845) );
  AND2_X1 U11451 ( .A1(n9983), .A2(n9751), .ZN(n18156) );
  INV_X2 U11452 ( .A(n16274), .ZN(n19186) );
  AOI21_X1 U11453 ( .B1(n10642), .B2(n10245), .A(n10244), .ZN(n11384) );
  NAND2_X1 U11454 ( .A1(n11142), .A2(n11141), .ZN(n17567) );
  NAND2_X2 U11455 ( .A1(n10224), .A2(n11354), .ZN(n11314) );
  XNOR2_X1 U11456 ( .A(n11210), .B(n17712), .ZN(n11039) );
  OR2_X1 U11457 ( .A1(n18167), .A2(n18174), .ZN(n9983) );
  OR2_X1 U11458 ( .A1(n13552), .A2(n13686), .ZN(n10116) );
  INV_X1 U11459 ( .A(n11143), .ZN(n18542) );
  AND3_X1 U11460 ( .A1(n11834), .A2(n14093), .A3(n11833), .ZN(n13551) );
  INV_X1 U11461 ( .A(n18524), .ZN(n11186) );
  OAI211_X1 U11462 ( .C1(n19495), .C2(n9718), .A(n11401), .B(n11400), .ZN(
        n11406) );
  NOR2_X1 U11463 ( .A1(n11879), .A2(n12006), .ZN(n12247) );
  CLKBUF_X1 U11464 ( .A(n11896), .Z(n11897) );
  INV_X1 U11465 ( .A(n17717), .ZN(n11210) );
  OAI211_X1 U11466 ( .C1(n9672), .C2(n17544), .A(n11003), .B(n11002), .ZN(
        n11205) );
  NOR2_X1 U11467 ( .A1(n11889), .A2(n9669), .ZN(n14856) );
  NAND2_X1 U11468 ( .A1(n19565), .A2(n20195), .ZN(n11421) );
  AOI211_X1 U11469 ( .C1(n17512), .C2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A(
        n11012), .B(n11011), .ZN(n11013) );
  INV_X1 U11470 ( .A(n9735), .ZN(n9683) );
  AND2_X2 U11471 ( .A1(n11889), .A2(n13675), .ZN(n14857) );
  NAND3_X1 U11472 ( .A1(n10976), .A2(n10975), .A3(n10974), .ZN(n17717) );
  CLKBUF_X3 U11473 ( .A(n9685), .Z(n19551) );
  INV_X1 U11474 ( .A(n11315), .ZN(n11321) );
  BUF_X2 U11475 ( .A(n10454), .Z(n15586) );
  AND2_X2 U11476 ( .A1(n11910), .A2(n12589), .ZN(n9717) );
  INV_X1 U11477 ( .A(n10236), .ZN(n10203) );
  AND2_X2 U11478 ( .A1(n10155), .A2(n10154), .ZN(n11315) );
  NAND2_X1 U11479 ( .A1(n11941), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12042) );
  NAND2_X1 U11480 ( .A1(n12770), .A2(n11891), .ZN(n13321) );
  NAND2_X2 U11482 ( .A1(n11875), .A2(n9852), .ZN(n13675) );
  NAND3_X1 U11483 ( .A1(n11037), .A2(n11038), .A3(n9771), .ZN(n18175) );
  NOR2_X1 U11484 ( .A1(n9854), .A2(n9853), .ZN(n9852) );
  AND2_X1 U11485 ( .A1(n10201), .A2(n10200), .ZN(n10219) );
  AND2_X2 U11486 ( .A1(n10218), .A2(n10217), .ZN(n19538) );
  NAND2_X1 U11487 ( .A1(n9974), .A2(n9972), .ZN(n10236) );
  OR2_X2 U11488 ( .A1(n16805), .A2(n16747), .ZN(n16807) );
  INV_X2 U11489 ( .A(U212), .ZN(n16791) );
  OR2_X1 U11490 ( .A1(n10991), .A2(n10990), .ZN(n10992) );
  OR2_X1 U11491 ( .A1(n10964), .A2(n10963), .ZN(n10965) );
  BUF_X1 U11492 ( .A(n11890), .Z(n14106) );
  AND2_X1 U11493 ( .A1(n9698), .A2(n11877), .ZN(n11876) );
  INV_X1 U11494 ( .A(n12589), .ZN(n14148) );
  AND2_X1 U11495 ( .A1(n9713), .A2(n9714), .ZN(n11147) );
  NOR2_X1 U11496 ( .A1(n17975), .A2(n17982), .ZN(n17963) );
  INV_X1 U11497 ( .A(n10248), .ZN(n9685) );
  NAND2_X2 U11498 ( .A1(n9739), .A2(n10087), .ZN(n11891) );
  NAND4_X2 U11499 ( .A1(n11854), .A2(n11853), .A3(n11852), .A4(n11851), .ZN(
        n11889) );
  AND4_X1 U11500 ( .A1(n11832), .A2(n11831), .A3(n11830), .A4(n11829), .ZN(
        n11890) );
  NAND2_X2 U11501 ( .A1(n13162), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12897) );
  AND4_X1 U11502 ( .A1(n11765), .A2(n11764), .A3(n11763), .A4(n11762), .ZN(
        n10087) );
  AND4_X1 U11503 ( .A1(n11794), .A2(n11793), .A3(n11792), .A4(n11791), .ZN(
        n11795) );
  AND4_X1 U11504 ( .A1(n11778), .A2(n11777), .A3(n11776), .A4(n11775), .ZN(
        n11784) );
  AND4_X1 U11505 ( .A1(n11748), .A2(n11747), .A3(n11746), .A4(n11745), .ZN(
        n11757) );
  AND4_X1 U11506 ( .A1(n11782), .A2(n11781), .A3(n11780), .A4(n11779), .ZN(
        n11783) );
  AND4_X1 U11507 ( .A1(n11842), .A2(n11841), .A3(n11840), .A4(n11839), .ZN(
        n11853) );
  AND4_X1 U11508 ( .A1(n11838), .A2(n11837), .A3(n11836), .A4(n11835), .ZN(
        n11854) );
  AND4_X1 U11509 ( .A1(n11769), .A2(n11768), .A3(n11767), .A4(n11766), .ZN(
        n11786) );
  AND3_X1 U11510 ( .A1(n11855), .A2(n11858), .A3(n11869), .ZN(n9851) );
  AND4_X1 U11511 ( .A1(n11874), .A2(n11873), .A3(n11872), .A4(n11871), .ZN(
        n11875) );
  AND4_X1 U11512 ( .A1(n11850), .A2(n11849), .A3(n11848), .A4(n11847), .ZN(
        n11851) );
  AND4_X1 U11513 ( .A1(n11846), .A2(n11845), .A3(n11844), .A4(n11843), .ZN(
        n11852) );
  AND4_X1 U11514 ( .A1(n11773), .A2(n11772), .A3(n11771), .A4(n11770), .ZN(
        n11785) );
  AND4_X1 U11515 ( .A1(n11828), .A2(n11827), .A3(n11826), .A4(n11825), .ZN(
        n11829) );
  AND4_X1 U11516 ( .A1(n11822), .A2(n11821), .A3(n11820), .A4(n11819), .ZN(
        n11830) );
  AND4_X1 U11518 ( .A1(n11818), .A2(n11817), .A3(n11816), .A4(n11815), .ZN(
        n11831) );
  AND4_X1 U11519 ( .A1(n11800), .A2(n11799), .A3(n11798), .A4(n11797), .ZN(
        n11810) );
  AOI22_X1 U11520 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11823), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11794) );
  NAND2_X2 U11521 ( .A1(n19126), .A2(n19065), .ZN(n19124) );
  NAND2_X2 U11522 ( .A1(n20233), .A2(n20101), .ZN(n20151) );
  CLKBUF_X2 U11523 ( .A(n11860), .Z(n12235) );
  NAND2_X1 U11524 ( .A1(n13090), .A2(n10359), .ZN(n12896) );
  CLKBUF_X1 U11525 ( .A(n10194), .Z(n13146) );
  CLKBUF_X1 U11526 ( .A(n13498), .Z(n19519) );
  INV_X2 U11527 ( .A(n16846), .ZN(n16848) );
  INV_X2 U11528 ( .A(n13007), .ZN(n12982) );
  OR2_X2 U11529 ( .A1(n10932), .A2(n18989), .ZN(n10946) );
  AND2_X2 U11530 ( .A1(n11743), .A2(n13857), .ZN(n9722) );
  AND2_X2 U11531 ( .A1(n11743), .A2(n13857), .ZN(n9723) );
  OAI21_X1 U11532 ( .B1(n13186), .B2(n13185), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13498) );
  OR2_X1 U11533 ( .A1(n10936), .A2(n10933), .ZN(n10948) );
  INV_X2 U11534 ( .A(n20234), .ZN(n20233) );
  NOR3_X2 U11535 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n10931), .ZN(n11156) );
  OR3_X1 U11536 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n10934), .ZN(n16118) );
  AND2_X1 U11537 ( .A1(n11741), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11749) );
  INV_X1 U11538 ( .A(n13115), .ZN(n13150) );
  NAND2_X1 U11539 ( .A1(n10369), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10142) );
  INV_X2 U11540 ( .A(n13007), .ZN(n9686) );
  NAND2_X1 U11541 ( .A1(n17155), .A2(n10091), .ZN(n18112) );
  OR3_X2 U11542 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n18989), .ZN(n11006) );
  NAND2_X1 U11543 ( .A1(n10936), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10932) );
  NAND4_X1 U11544 ( .A1(n10936), .A2(n9997), .A3(n10935), .A4(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n17455) );
  INV_X1 U11545 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10117) );
  AND2_X1 U11546 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10370) );
  INV_X2 U11547 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n20195) );
  INV_X1 U11548 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9715) );
  INV_X1 U11549 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9716) );
  INV_X1 U11550 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9998) );
  NOR2_X2 U11551 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13859) );
  AND2_X4 U11552 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13857) );
  AND2_X1 U11553 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13858) );
  AND2_X4 U11554 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13559) );
  NAND2_X1 U11555 ( .A1(n14476), .A2(n9697), .ZN(n9694) );
  AOI211_X1 U11556 ( .C1(n17508), .C2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n17318), .B(n17317), .ZN(n17319) );
  NAND2_X2 U11557 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18138), .ZN(n18024) );
  NAND2_X1 U11558 ( .A1(n13201), .A2(n9691), .ZN(n9688) );
  AND2_X1 U11559 ( .A1(n9688), .A2(n9689), .ZN(n13204) );
  OR2_X1 U11560 ( .A1(n9690), .A2(n16601), .ZN(n9689) );
  INV_X1 U11561 ( .A(n10065), .ZN(n9690) );
  AND2_X1 U11562 ( .A1(n16023), .A2(n10065), .ZN(n9691) );
  NAND2_X1 U11563 ( .A1(n10264), .A2(n10255), .ZN(n9692) );
  NAND2_X1 U11564 ( .A1(n10264), .A2(n10255), .ZN(n10292) );
  OAI21_X1 U11566 ( .B1(n15557), .B2(n15552), .A(n13142), .ZN(n15546) );
  XNOR2_X1 U11567 ( .A(n13740), .B(n13744), .ZN(n20167) );
  AND2_X1 U11568 ( .A1(n10221), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n20224) );
  NAND2_X1 U11569 ( .A1(n10244), .A2(n10221), .ZN(n10256) );
  XNOR2_X1 U11570 ( .A(n9693), .B(n11279), .ZN(n15846) );
  AND2_X1 U11571 ( .A1(n11278), .A2(n14809), .ZN(n9693) );
  AND2_X4 U11572 ( .A1(n9694), .A2(n9695), .ZN(n15230) );
  OR2_X1 U11573 ( .A1(n9696), .A2(n10080), .ZN(n9695) );
  INV_X1 U11574 ( .A(n13305), .ZN(n9696) );
  NAND4_X1 U11575 ( .A1(n11832), .A2(n11831), .A3(n11830), .A4(n11829), .ZN(
        n9698) );
  OR2_X1 U11576 ( .A1(n15225), .A2(n13317), .ZN(n9764) );
  NAND2_X1 U11577 ( .A1(n9764), .A2(n10075), .ZN(n15186) );
  XNOR2_X1 U11578 ( .A(n11053), .B(n11052), .ZN(n18102) );
  CLKBUF_X1 U11579 ( .A(n15186), .Z(n9699) );
  OAI21_X1 U11580 ( .B1(n15230), .B2(n10074), .A(n10072), .ZN(n9700) );
  OAI21_X1 U11581 ( .B1(n15230), .B2(n10074), .A(n10072), .ZN(n15225) );
  NAND2_X1 U11582 ( .A1(n17691), .A2(n11245), .ZN(n11254) );
  OAI21_X2 U11583 ( .B1(n15827), .B2(n10059), .A(n10057), .ZN(n9701) );
  OAI21_X1 U11584 ( .B1(n15827), .B2(n10059), .A(n10057), .ZN(n9702) );
  OAI21_X1 U11585 ( .B1(n15827), .B2(n10059), .A(n10057), .ZN(n16037) );
  OR2_X1 U11586 ( .A1(n10425), .A2(n10424), .ZN(n10427) );
  OAI211_X1 U11587 ( .C1(n10605), .C2(n10808), .A(n10603), .B(n9979), .ZN(
        n15830) );
  AND2_X1 U11588 ( .A1(n9807), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9703) );
  NAND2_X1 U11589 ( .A1(n9845), .A2(n9707), .ZN(n9704) );
  OR2_X1 U11590 ( .A1(n9706), .A2(n9674), .ZN(n9705) );
  INV_X1 U11591 ( .A(n9762), .ZN(n9706) );
  AND2_X1 U11592 ( .A1(n10070), .A2(n9762), .ZN(n9707) );
  NAND2_X1 U11593 ( .A1(n14476), .A2(n13303), .ZN(n9708) );
  NAND2_X1 U11594 ( .A1(n14476), .A2(n13303), .ZN(n10081) );
  AND4_X1 U11595 ( .A1(n11814), .A2(n11813), .A3(n11812), .A4(n11811), .ZN(
        n11832) );
  NOR2_X2 U11596 ( .A1(n13722), .A2(n9904), .ZN(n13889) );
  NOR3_X4 U11597 ( .A1(n15673), .A2(n9889), .A3(n9891), .ZN(n15641) );
  AND2_X1 U11598 ( .A1(n11390), .A2(n20195), .ZN(n9908) );
  AND4_X1 U11599 ( .A1(n19565), .A2(n9685), .A3(n13746), .A4(n11315), .ZN(
        n13172) );
  INV_X1 U11600 ( .A(n9717), .ZN(n11906) );
  OR2_X1 U11601 ( .A1(n9711), .A2(n17786), .ZN(n9710) );
  INV_X1 U11602 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n9711) );
  NAND2_X1 U11603 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17573), .ZN(n9712) );
  NAND2_X1 U11604 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n9713) );
  NAND2_X1 U11605 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17508), .ZN(
        n9714) );
  NOR2_X2 U11606 ( .A1(n11893), .A2(n13550), .ZN(n11915) );
  OR2_X1 U11607 ( .A1(n15837), .A2(n16668), .ZN(n9978) );
  NAND2_X2 U11608 ( .A1(n14592), .A2(n14593), .ZN(n15827) );
  NAND2_X2 U11609 ( .A1(n10806), .A2(n10805), .ZN(n14592) );
  NOR2_X4 U11610 ( .A1(n13836), .A2(n12820), .ZN(n13838) );
  OAI21_X2 U11611 ( .B1(n13740), .B2(n12819), .A(n12818), .ZN(n13836) );
  NAND2_X1 U11612 ( .A1(n19565), .A2(n20195), .ZN(n9718) );
  NAND2_X2 U11613 ( .A1(n11884), .A2(n11883), .ZN(n11900) );
  AOI21_X2 U11614 ( .B1(n11896), .B2(n11878), .A(n15052), .ZN(n11884) );
  OAI22_X1 U11615 ( .A1(n12843), .A2(n10492), .B1(n10487), .B2(n10323), .ZN(
        n10324) );
  AND2_X1 U11616 ( .A1(n13859), .A2(n13559), .ZN(n9719) );
  NOR2_X1 U11617 ( .A1(n10932), .A2(n10931), .ZN(n10977) );
  NAND2_X1 U11618 ( .A1(n19538), .A2(n10219), .ZN(n10271) );
  INV_X2 U11619 ( .A(n13007), .ZN(n9721) );
  NAND2_X1 U11620 ( .A1(n9850), .A2(n10069), .ZN(n15124) );
  INV_X1 U11621 ( .A(n10601), .ZN(n9843) );
  AND2_X2 U11622 ( .A1(n11743), .A2(n13857), .ZN(n12509) );
  NOR2_X2 U11623 ( .A1(n15776), .A2(n15775), .ZN(n15781) );
  XNOR2_X1 U11624 ( .A(n11701), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9724) );
  OAI211_X1 U11625 ( .C1(n10109), .C2(n17492), .A(n11087), .B(n11086), .ZN(
        n16274) );
  XNOR2_X2 U11626 ( .A(n10804), .B(n14462), .ZN(n14442) );
  NAND2_X2 U11627 ( .A1(n10780), .A2(n19435), .ZN(n10804) );
  AND2_X4 U11628 ( .A1(n11751), .A2(n11750), .ZN(n11866) );
  AND2_X1 U11629 ( .A1(n11751), .A2(n13858), .ZN(n9726) );
  AND2_X2 U11630 ( .A1(n11751), .A2(n13858), .ZN(n12527) );
  NAND2_X2 U11631 ( .A1(n13295), .A2(n16369), .ZN(n14476) );
  AOI22_X1 U11632 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14838), .B1(n15698), 
        .B2(n20218), .ZN(n9727) );
  AOI22_X1 U11633 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n14838), .B1(n15698), 
        .B2(n20218), .ZN(n9728) );
  NAND2_X2 U11634 ( .A1(n20420), .A2(n13266), .ZN(n16381) );
  NAND2_X2 U11635 ( .A1(n20418), .A2(n20417), .ZN(n20420) );
  NAND2_X2 U11636 ( .A1(n13671), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13672) );
  AND2_X4 U11637 ( .A1(n11750), .A2(n13559), .ZN(n11861) );
  NAND2_X2 U11638 ( .A1(n13897), .A2(n13896), .ZN(n13898) );
  XNOR2_X2 U11639 ( .A(n13252), .B(n20464), .ZN(n13897) );
  OAI222_X1 U11640 ( .A1(n17554), .A2(n17559), .B1(n17553), .B2(n9732), .C1(
        n17552), .C2(n17551), .ZN(P3_U2702) );
  AOI221_X1 U11641 ( .B1(n17547), .B2(n9732), .C1(n17691), .C2(n9732), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17549) );
  NAND2_X2 U11642 ( .A1(n13672), .A2(n13245), .ZN(n13252) );
  XNOR2_X2 U11643 ( .A(n13243), .B(n13710), .ZN(n13671) );
  NOR2_X4 U11644 ( .A1(n11900), .A2(n11886), .ZN(n12572) );
  NAND2_X2 U11645 ( .A1(n12572), .A2(n14133), .ZN(n13557) );
  NAND2_X2 U11646 ( .A1(n13711), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13710) );
  OAI21_X2 U11647 ( .B1(n13236), .B2(n13235), .A(n13234), .ZN(n13711) );
  BUF_X1 U11648 ( .A(n12808), .Z(n9733) );
  BUF_X4 U11649 ( .A(n12808), .Z(n9734) );
  OAI21_X2 U11650 ( .B1(n11888), .B2(n13692), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11964) );
  NAND2_X2 U11651 ( .A1(n11964), .A2(n11903), .ZN(n11979) );
  XNOR2_X2 U11652 ( .A(n13258), .B(n20447), .ZN(n13962) );
  NAND2_X2 U11653 ( .A1(n13898), .A2(n13253), .ZN(n13258) );
  AND2_X4 U11654 ( .A1(n10368), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13091) );
  NAND2_X2 U11655 ( .A1(n11905), .A2(n11904), .ZN(n11967) );
  NOR2_X1 U11656 ( .A1(n9684), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n9735) );
  NOR2_X1 U11657 ( .A1(n9684), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11397) );
  AND4_X1 U11658 ( .A1(n10561), .A2(n10560), .A3(n10559), .A4(n10558), .ZN(
        n10574) );
  AND2_X1 U11659 ( .A1(n15561), .A2(n15562), .ZN(n15564) );
  AND2_X1 U11660 ( .A1(n11335), .A2(n13336), .ZN(n11388) );
  INV_X1 U11661 ( .A(n12111), .ZN(n9856) );
  OAI21_X1 U11662 ( .B1(n12630), .B2(n12746), .A(n10116), .ZN(n11888) );
  NOR2_X1 U11663 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n12578), .ZN(
        n12580) );
  NOR2_X1 U11664 ( .A1(n15759), .A2(n9917), .ZN(n9916) );
  INV_X1 U11665 ( .A(n9918), .ZN(n9917) );
  OAI211_X1 U11666 ( .C1(n10239), .C2(n10238), .A(n11354), .B(n10237), .ZN(
        n11360) );
  AND3_X1 U11667 ( .A1(n9685), .A2(n10203), .A3(n11390), .ZN(n10220) );
  INV_X1 U11668 ( .A(n12537), .ZN(n12631) );
  INV_X1 U11669 ( .A(n12631), .ZN(n12560) );
  NOR2_X1 U11670 ( .A1(n14705), .A2(n15303), .ZN(n10068) );
  OR2_X1 U11671 ( .A1(n9886), .A2(n9796), .ZN(n14931) );
  NOR2_X1 U11672 ( .A1(n12663), .A2(n9865), .ZN(n9864) );
  INV_X1 U11673 ( .A(n14382), .ZN(n9865) );
  NAND2_X1 U11674 ( .A1(n12739), .A2(n14857), .ZN(n12738) );
  OR2_X1 U11675 ( .A1(n9698), .A2(n21023), .ZN(n12041) );
  NAND2_X1 U11676 ( .A1(n12042), .A2(n12041), .ZN(n12596) );
  AND3_X1 U11677 ( .A1(n9698), .A2(n11889), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12619) );
  NOR2_X1 U11678 ( .A1(n15819), .A2(n10063), .ZN(n10062) );
  INV_X1 U11679 ( .A(n15988), .ZN(n10063) );
  OR2_X1 U11680 ( .A1(n16009), .A2(n9898), .ZN(n9897) );
  INV_X1 U11681 ( .A(n14354), .ZN(n9898) );
  NOR2_X1 U11682 ( .A1(n13723), .A2(n9907), .ZN(n9906) );
  INV_X1 U11683 ( .A(n13760), .ZN(n9907) );
  NAND2_X1 U11684 ( .A1(n9715), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10934) );
  NOR2_X1 U11685 ( .A1(n17697), .A2(n11049), .ZN(n11715) );
  NAND2_X1 U11686 ( .A1(n9982), .A2(n9981), .ZN(n11042) );
  INV_X1 U11687 ( .A(n13682), .ZN(n14851) );
  NAND2_X1 U11688 ( .A1(n13682), .A2(n14860), .ZN(n14086) );
  INV_X1 U11689 ( .A(n13811), .ZN(n12769) );
  AND2_X1 U11690 ( .A1(n14871), .A2(n14687), .ZN(n14689) );
  NOR2_X1 U11691 ( .A1(n14891), .A2(n9888), .ZN(n14871) );
  OR2_X1 U11692 ( .A1(n14884), .A2(n14872), .ZN(n9888) );
  INV_X1 U11693 ( .A(n13983), .ZN(n12658) );
  INV_X1 U11694 ( .A(n14065), .ZN(n12659) );
  INV_X1 U11695 ( .A(n14857), .ZN(n14084) );
  AND3_X1 U11696 ( .A1(n11627), .A2(n11626), .A3(n11625), .ZN(n15659) );
  NOR2_X1 U11697 ( .A1(n10013), .A2(n10849), .ZN(n10012) );
  INV_X1 U11698 ( .A(n10014), .ZN(n10013) );
  NAND2_X1 U11699 ( .A1(n10229), .A2(n13172), .ZN(n13997) );
  NOR2_X1 U11700 ( .A1(n11336), .A2(n10271), .ZN(n10229) );
  NAND2_X1 U11701 ( .A1(n11644), .A2(n11643), .ZN(n14827) );
  OR2_X1 U11702 ( .A1(n9892), .A2(n15659), .ZN(n9891) );
  NAND2_X1 U11704 ( .A1(n15564), .A2(n9955), .ZN(n14835) );
  NOR2_X1 U11705 ( .A1(n10749), .A2(n9956), .ZN(n9955) );
  INV_X1 U11706 ( .A(n15509), .ZN(n9956) );
  AND4_X1 U11707 ( .A1(n10565), .A2(n10564), .A3(n10563), .A4(n10562), .ZN(
        n10573) );
  NOR2_X1 U11708 ( .A1(n11637), .A2(n15730), .ZN(n9928) );
  NAND2_X1 U11709 ( .A1(n9766), .A2(n9930), .ZN(n9929) );
  INV_X1 U11710 ( .A(n15712), .ZN(n10913) );
  AND2_X1 U11711 ( .A1(n9924), .A2(n15714), .ZN(n9921) );
  OAI21_X1 U11712 ( .B1(n9941), .B2(n16716), .A(n9936), .ZN(n9935) );
  INV_X1 U11713 ( .A(n16494), .ZN(n9941) );
  OR2_X1 U11714 ( .A1(n15844), .A2(n9938), .ZN(n9937) );
  AOI21_X1 U11715 ( .B1(n15848), .B2(n16710), .A(n15847), .ZN(n15849) );
  AOI22_X1 U11716 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14148), .B1(n12596), 
        .B2(n9669), .ZN(n12603) );
  NOR2_X1 U11717 ( .A1(n15584), .A2(n13027), .ZN(n10025) );
  NAND2_X1 U11718 ( .A1(n12576), .A2(n12575), .ZN(n12583) );
  AND2_X1 U11719 ( .A1(n12186), .A2(n14487), .ZN(n10044) );
  INV_X1 U11720 ( .A(n11897), .ZN(n13673) );
  OR2_X1 U11721 ( .A1(n12001), .A2(n12000), .ZN(n12002) );
  INV_X1 U11722 ( .A(n12002), .ZN(n13255) );
  NAND2_X1 U11723 ( .A1(n12589), .A2(n11890), .ZN(n13323) );
  XNOR2_X1 U11724 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10631) );
  NAND2_X1 U11725 ( .A1(n10621), .A2(n10627), .ZN(n10632) );
  AND2_X1 U11726 ( .A1(n10554), .A2(n10553), .ZN(n11429) );
  AND2_X1 U11727 ( .A1(n19538), .A2(n15586), .ZN(n10245) );
  NAND2_X1 U11728 ( .A1(n10449), .A2(n10448), .ZN(n10450) );
  INV_X1 U11729 ( .A(n10436), .ZN(n10437) );
  NOR2_X1 U11730 ( .A1(n17704), .A2(n11216), .ZN(n11204) );
  NAND2_X1 U11731 ( .A1(n18175), .A2(n17717), .ZN(n11207) );
  AOI21_X1 U11732 ( .B1(n19010), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11167), .ZN(n11173) );
  NOR2_X1 U11733 ( .A1(n11186), .A2(n11234), .ZN(n11235) );
  INV_X1 U11734 ( .A(n14918), .ZN(n10052) );
  AND2_X1 U11735 ( .A1(n10054), .A2(n14930), .ZN(n10053) );
  NAND2_X1 U11736 ( .A1(n12285), .A2(n10040), .ZN(n10039) );
  INV_X1 U11737 ( .A(n15005), .ZN(n10040) );
  NAND2_X1 U11738 ( .A1(n13673), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12563) );
  AND2_X1 U11739 ( .A1(n10042), .A2(n14571), .ZN(n10041) );
  XNOR2_X1 U11740 ( .A(n13298), .B(n12133), .ZN(n13292) );
  NAND2_X1 U11741 ( .A1(n14587), .A2(n9883), .ZN(n9886) );
  NOR2_X1 U11742 ( .A1(n9885), .A2(n12706), .ZN(n9883) );
  NOR2_X1 U11743 ( .A1(n14589), .A2(n14588), .ZN(n14587) );
  INV_X1 U11744 ( .A(n12738), .ZN(n12730) );
  AND2_X1 U11745 ( .A1(n13285), .A2(n16380), .ZN(n10077) );
  INV_X1 U11746 ( .A(n13277), .ZN(n10079) );
  NAND2_X1 U11747 ( .A1(n10067), .A2(n13242), .ZN(n13243) );
  AND3_X1 U11748 ( .A1(n11960), .A2(n11959), .A3(n11958), .ZN(n11973) );
  OR2_X1 U11749 ( .A1(n12052), .A2(n12051), .ZN(n13270) );
  AOI21_X1 U11750 ( .B1(n11902), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11901), 
        .ZN(n11903) );
  AND2_X1 U11751 ( .A1(n11900), .A2(n12003), .ZN(n11901) );
  NOR2_X2 U11752 ( .A1(n10907), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10915) );
  NAND2_X1 U11753 ( .A1(n10890), .A2(n10906), .ZN(n10838) );
  NOR2_X1 U11754 ( .A1(n10854), .A2(n10015), .ZN(n10014) );
  INV_X1 U11755 ( .A(n10831), .ZN(n10015) );
  INV_X1 U11756 ( .A(n10810), .ZN(n10008) );
  INV_X1 U11757 ( .A(n10812), .ZN(n10009) );
  OAI211_X1 U11758 ( .C1(n9657), .C2(n10287), .A(n10286), .B(n10285), .ZN(
        n10288) );
  INV_X1 U11759 ( .A(n12906), .ZN(n12951) );
  INV_X1 U11760 ( .A(n12905), .ZN(n12956) );
  NOR2_X2 U11761 ( .A1(n15619), .A2(n15620), .ZN(n11644) );
  NOR2_X1 U11762 ( .A1(n14624), .A2(n14642), .ZN(n10024) );
  AND2_X1 U11763 ( .A1(n12795), .A2(n10203), .ZN(n13750) );
  AND2_X1 U11764 ( .A1(n15586), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12795) );
  NOR2_X1 U11765 ( .A1(n10454), .A2(n10221), .ZN(n10225) );
  NAND2_X1 U11766 ( .A1(n10737), .A2(n9951), .ZN(n9950) );
  INV_X1 U11767 ( .A(n15581), .ZN(n9951) );
  NAND2_X1 U11768 ( .A1(n9947), .A2(n13851), .ZN(n9946) );
  INV_X1 U11769 ( .A(n13831), .ZN(n9947) );
  OR2_X1 U11770 ( .A1(n9932), .A2(n11637), .ZN(n9931) );
  INV_X1 U11771 ( .A(n15714), .ZN(n9932) );
  NAND2_X1 U11772 ( .A1(n16520), .A2(n14818), .ZN(n10920) );
  AND2_X1 U11773 ( .A1(n9914), .A2(n15760), .ZN(n9913) );
  NOR2_X1 U11774 ( .A1(n14628), .A2(n14627), .ZN(n14626) );
  NAND2_X1 U11775 ( .A1(n9701), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10868) );
  NAND2_X1 U11776 ( .A1(n13889), .A2(n13926), .ZN(n13925) );
  OR2_X1 U11777 ( .A1(n10821), .A2(n10060), .ZN(n10059) );
  INV_X1 U11778 ( .A(n16624), .ZN(n10060) );
  NAND2_X1 U11779 ( .A1(n9945), .A2(n13907), .ZN(n9944) );
  INV_X1 U11780 ( .A(n9946), .ZN(n9945) );
  OAI211_X1 U11781 ( .C1(n9843), .C2(n10781), .A(n9842), .B(n9841), .ZN(n10575) );
  NAND2_X1 U11782 ( .A1(n10602), .A2(n14818), .ZN(n9842) );
  NAND2_X1 U11783 ( .A1(n9843), .A2(n9759), .ZN(n9841) );
  AOI21_X1 U11784 ( .B1(n10654), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10302), .ZN(n10306) );
  NAND2_X1 U11785 ( .A1(n10306), .A2(n10307), .ZN(n10658) );
  NAND2_X1 U11786 ( .A1(n10202), .A2(n19543), .ZN(n10204) );
  OR2_X1 U11787 ( .A1(n11365), .A2(n11364), .ZN(n13999) );
  INV_X1 U11788 ( .A(n10345), .ZN(n10350) );
  AOI211_X1 U11789 ( .C1(n17403), .C2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n11134), .B(n11133), .ZN(n11135) );
  INV_X1 U11790 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17419) );
  NOR2_X1 U11791 ( .A1(n17935), .A2(n17920), .ZN(n17921) );
  NAND2_X1 U11792 ( .A1(n17765), .A2(n14655), .ZN(n13364) );
  NAND2_X1 U11793 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18094), .ZN(
        n11229) );
  NOR2_X1 U11794 ( .A1(n18109), .A2(n11051), .ZN(n11053) );
  AND2_X1 U11795 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11050), .ZN(
        n11051) );
  NOR2_X1 U11796 ( .A1(n17704), .A2(n11044), .ZN(n11048) );
  NOR2_X1 U11797 ( .A1(n11043), .A2(n18142), .ZN(n11046) );
  XNOR2_X1 U11798 ( .A(n11207), .B(n9813), .ZN(n11208) );
  INV_X1 U11799 ( .A(n17712), .ZN(n9813) );
  INV_X1 U11800 ( .A(n11165), .ZN(n9965) );
  NAND2_X1 U11801 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n9964) );
  INV_X1 U11802 ( .A(n11164), .ZN(n9966) );
  NAND2_X1 U11803 ( .A1(n20334), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n14163) );
  NAND2_X1 U11804 ( .A1(n14551), .A2(n9875), .ZN(n14589) );
  NOR2_X1 U11805 ( .A1(n9876), .A2(n9882), .ZN(n9875) );
  INV_X1 U11806 ( .A(n14576), .ZN(n9882) );
  INV_X1 U11807 ( .A(n9877), .ZN(n9876) );
  OR2_X1 U11808 ( .A1(n13699), .A2(n12776), .ZN(n14850) );
  AOI21_X1 U11809 ( .B1(n12010), .B2(n12264), .A(n10035), .ZN(n10034) );
  INV_X1 U11810 ( .A(n12032), .ZN(n10035) );
  OR2_X1 U11811 ( .A1(n13572), .A2(n14160), .ZN(n14088) );
  OR2_X1 U11812 ( .A1(n12353), .A2(n14978), .ZN(n12374) );
  OAI211_X1 U11813 ( .C1(n12127), .C2(n20363), .A(n12126), .B(n12125), .ZN(
        n14281) );
  NAND2_X1 U11814 ( .A1(n12084), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12105) );
  NAND2_X1 U11815 ( .A1(n14911), .A2(n14892), .ZN(n14891) );
  NOR2_X1 U11816 ( .A1(n14933), .A2(n14920), .ZN(n14919) );
  INV_X1 U11817 ( .A(n15224), .ZN(n10071) );
  OR2_X1 U11818 ( .A1(n14431), .A2(n14430), .ZN(n14558) );
  AND2_X1 U11819 ( .A1(n12667), .A2(n12666), .ZN(n14382) );
  NAND2_X1 U11820 ( .A1(n9863), .A2(n9864), .ZN(n14407) );
  INV_X1 U11821 ( .A(n13903), .ZN(n9871) );
  NOR2_X1 U11822 ( .A1(n9874), .A2(n9873), .ZN(n9872) );
  INV_X1 U11823 ( .A(n13827), .ZN(n9874) );
  NAND2_X1 U11824 ( .A1(n13691), .A2(n13690), .ZN(n13703) );
  INV_X1 U11825 ( .A(n11938), .ZN(n11939) );
  NOR2_X2 U11826 ( .A1(n11891), .A2(n13678), .ZN(n13865) );
  NAND2_X1 U11827 ( .A1(n14388), .A2(n13254), .ZN(n20580) );
  INV_X1 U11828 ( .A(n13949), .ZN(n14388) );
  NAND2_X1 U11829 ( .A1(n13949), .A2(n13954), .ZN(n20649) );
  NOR2_X1 U11830 ( .A1(n14500), .A2(n20674), .ZN(n20773) );
  OR2_X1 U11831 ( .A1(n13254), .A2(n13949), .ZN(n20812) );
  NOR2_X1 U11832 ( .A1(n20771), .A2(n14500), .ZN(n20847) );
  OR2_X1 U11833 ( .A1(n15489), .A2(n13236), .ZN(n20739) );
  NAND2_X1 U11834 ( .A1(n15489), .A2(n13236), .ZN(n20839) );
  NOR2_X1 U11835 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14105), .ZN(n14117) );
  INV_X1 U11836 ( .A(n14117), .ZN(n14500) );
  NAND2_X1 U11837 ( .A1(n15489), .A2(n14232), .ZN(n20579) );
  NAND2_X1 U11838 ( .A1(n13949), .A2(n13950), .ZN(n20885) );
  NAND2_X1 U11839 ( .A1(n12629), .A2(n12628), .ZN(n13682) );
  OR2_X1 U11840 ( .A1(n12615), .A2(n12590), .ZN(n12629) );
  INV_X1 U11841 ( .A(n10003), .ZN(n16534) );
  INV_X1 U11842 ( .A(n10779), .ZN(n10002) );
  NAND2_X1 U11843 ( .A1(n10782), .A2(n10798), .ZN(n10801) );
  NAND2_X1 U11844 ( .A1(n10283), .A2(n10282), .ZN(n10309) );
  INV_X1 U11845 ( .A(n14021), .ZN(n13408) );
  INV_X1 U11846 ( .A(n12907), .ZN(n12953) );
  NAND2_X1 U11847 ( .A1(n9745), .A2(n10018), .ZN(n10017) );
  INV_X1 U11848 ( .A(n15558), .ZN(n10018) );
  OR2_X1 U11849 ( .A1(n15674), .A2(n9890), .ZN(n9889) );
  INV_X1 U11850 ( .A(n15651), .ZN(n9890) );
  OR2_X1 U11851 ( .A1(n15593), .A2(n15594), .ZN(n10029) );
  AND4_X1 U11852 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n16009) );
  OR2_X1 U11853 ( .A1(n11566), .A2(n11565), .ZN(n14159) );
  AND4_X1 U11854 ( .A1(n11456), .A2(n11455), .A3(n11454), .A4(n11453), .ZN(
        n13723) );
  INV_X1 U11855 ( .A(n19210), .ZN(n13336) );
  AND2_X1 U11856 ( .A1(n9958), .A2(n14300), .ZN(n9957) );
  NAND2_X1 U11857 ( .A1(n15707), .A2(n15714), .ZN(n9926) );
  NAND2_X1 U11858 ( .A1(n14433), .A2(n15971), .ZN(n14628) );
  AND2_X1 U11859 ( .A1(n13210), .A2(n13209), .ZN(n15811) );
  INV_X1 U11860 ( .A(n15992), .ZN(n9840) );
  OR3_X1 U11861 ( .A1(n10881), .A2(n10781), .A3(n15966), .ZN(n15987) );
  NAND2_X1 U11862 ( .A1(n10611), .A2(n10610), .ZN(n16053) );
  NAND2_X1 U11863 ( .A1(n15831), .A2(n10607), .ZN(n10608) );
  INV_X1 U11864 ( .A(n14219), .ZN(n9893) );
  INV_X1 U11865 ( .A(n14792), .ZN(n13622) );
  XNOR2_X1 U11866 ( .A(n14792), .B(n12801), .ZN(n13636) );
  AOI21_X1 U11867 ( .B1(n14327), .B2(n12809), .A(n12797), .ZN(n13635) );
  NAND2_X1 U11868 ( .A1(n13635), .A2(n13636), .ZN(n13638) );
  AND2_X1 U11869 ( .A1(n20218), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12809) );
  NAND2_X1 U11870 ( .A1(n20167), .A2(n20197), .ZN(n19719) );
  AND2_X1 U11871 ( .A1(n20167), .A2(n19779), .ZN(n19758) );
  OR2_X1 U11872 ( .A1(n20178), .A2(n20190), .ZN(n19940) );
  NAND2_X1 U11873 ( .A1(n10153), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10154) );
  OR2_X1 U11874 ( .A1(n20167), .A2(n20197), .ZN(n19941) );
  OAI21_X2 U11875 ( .B1(n20161), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16271), 
        .ZN(n20022) );
  INV_X1 U11876 ( .A(n20022), .ZN(n19947) );
  NAND2_X1 U11877 ( .A1(n19942), .A2(n20195), .ZN(n20016) );
  NOR2_X1 U11878 ( .A1(n11311), .A2(n11310), .ZN(n14310) );
  AND2_X1 U11879 ( .A1(n11309), .A2(n20224), .ZN(n11310) );
  INV_X1 U11880 ( .A(n11181), .ZN(n18970) );
  NOR2_X1 U11881 ( .A1(n17175), .A2(n17005), .ZN(n17030) );
  NOR2_X1 U11882 ( .A1(n10985), .A2(n10984), .ZN(n10988) );
  NOR2_X1 U11883 ( .A1(n10949), .A2(n17353), .ZN(n10984) );
  OR2_X1 U11884 ( .A1(n10983), .A2(n10982), .ZN(n10985) );
  AOI21_X1 U11885 ( .B1(n16093), .B2(n18967), .A(n9969), .ZN(n16275) );
  NOR2_X1 U11886 ( .A1(n16092), .A2(n9970), .ZN(n9969) );
  NAND2_X1 U11887 ( .A1(n18548), .A2(n18533), .ZN(n9970) );
  AND2_X1 U11888 ( .A1(n17512), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n10963) );
  NOR2_X1 U11889 ( .A1(n10946), .A2(n17493), .ZN(n10968) );
  AND2_X1 U11890 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10972) );
  NOR2_X1 U11891 ( .A1(n11693), .A2(n16901), .ZN(n16733) );
  NOR2_X1 U11892 ( .A1(n17907), .A2(n17908), .ZN(n17887) );
  NAND2_X1 U11893 ( .A1(n13359), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n17907) );
  AND2_X1 U11894 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U11895 ( .A1(n17403), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11087) );
  AOI211_X1 U11896 ( .C1(n17512), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(
        n11085), .B(n11084), .ZN(n11086) );
  XNOR2_X1 U11897 ( .A(n11208), .B(n11027), .ZN(n18158) );
  OR2_X1 U11898 ( .A1(n9675), .A2(n17878), .ZN(n11065) );
  NAND2_X1 U11899 ( .A1(n18011), .A2(n18280), .ZN(n18312) );
  NAND2_X1 U11900 ( .A1(n18524), .A2(n18529), .ZN(n18981) );
  AND2_X1 U11901 ( .A1(n10103), .A2(n18378), .ZN(n9996) );
  INV_X1 U11902 ( .A(n9818), .ZN(n11217) );
  OR2_X1 U11903 ( .A1(n18121), .A2(n18120), .ZN(n9819) );
  INV_X1 U11904 ( .A(n19036), .ZN(n19180) );
  NOR2_X2 U11905 ( .A1(n14737), .A2(n14165), .ZN(n20287) );
  XNOR2_X1 U11906 ( .A(n12744), .B(n12743), .ZN(n15016) );
  NAND2_X1 U11907 ( .A1(n12742), .A2(n12741), .ZN(n12744) );
  OR2_X1 U11908 ( .A1(n14689), .A2(n12739), .ZN(n12742) );
  OAI21_X1 U11909 ( .B1(n9846), .B2(n15124), .A(n9847), .ZN(n14710) );
  OR2_X1 U11910 ( .A1(n13324), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20432) );
  CLKBUF_X1 U11911 ( .A(n14391), .Z(n14392) );
  NAND2_X1 U11912 ( .A1(n14097), .A2(n20766), .ZN(n20810) );
  INV_X1 U11913 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n20226) );
  NAND2_X1 U11914 ( .A1(n11331), .A2(n10653), .ZN(n19212) );
  OR2_X1 U11915 ( .A1(n19462), .A2(n13188), .ZN(n15692) );
  OR2_X1 U11916 ( .A1(n19462), .A2(n13193), .ZN(n15690) );
  INV_X2 U11917 ( .A(n19462), .ZN(n15689) );
  INV_X1 U11918 ( .A(n20197), .ZN(n19779) );
  AND2_X1 U11919 ( .A1(n16677), .A2(n13460), .ZN(n16667) );
  AND2_X1 U11920 ( .A1(n16677), .A2(n20184), .ZN(n19504) );
  NOR2_X1 U11921 ( .A1(n14835), .A2(n14834), .ZN(n14840) );
  AND2_X1 U11922 ( .A1(n14833), .A2(n14832), .ZN(n14842) );
  AOI21_X1 U11923 ( .B1(n19448), .B2(n16710), .A(n15700), .ZN(n14833) );
  XNOR2_X1 U11924 ( .A(n14822), .B(n14838), .ZN(n15704) );
  OAI211_X1 U11925 ( .C1(n9927), .C2(n9923), .A(n14811), .B(n9922), .ZN(n14821) );
  NOR2_X1 U11926 ( .A1(n15857), .A2(n15852), .ZN(n9901) );
  NAND2_X1 U11927 ( .A1(n15853), .A2(n16700), .ZN(n9899) );
  NOR2_X1 U11928 ( .A1(n15729), .A2(n15713), .ZN(n15716) );
  NAND2_X1 U11929 ( .A1(n9836), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9835) );
  NAND2_X1 U11930 ( .A1(n15986), .A2(n9837), .ZN(n9836) );
  NAND2_X1 U11931 ( .A1(n14598), .A2(n15985), .ZN(n9837) );
  AND2_X1 U11932 ( .A1(n11388), .A2(n20206), .ZN(n16700) );
  NAND2_X1 U11933 ( .A1(n11388), .A2(n11347), .ZN(n16716) );
  AND2_X1 U11934 ( .A1(n11388), .A2(n20207), .ZN(n16721) );
  INV_X1 U11935 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20202) );
  INV_X1 U11936 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20193) );
  INV_X1 U11937 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20175) );
  NAND2_X1 U11938 ( .A1(n16893), .A2(n17233), .ZN(n9827) );
  NAND2_X1 U11939 ( .A1(n17270), .A2(n17269), .ZN(n9961) );
  NAND2_X1 U11940 ( .A1(n17279), .A2(n9795), .ZN(n17267) );
  NOR2_X1 U11941 ( .A1(n17323), .A2(n16974), .ZN(n17290) );
  NAND2_X1 U11942 ( .A1(n17336), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n17323) );
  INV_X1 U11943 ( .A(n18090), .ZN(n18027) );
  NAND2_X1 U11944 ( .A1(n17692), .A2(n9729), .ZN(n18093) );
  AND2_X1 U11945 ( .A1(n11727), .A2(n11726), .ZN(n11730) );
  NAND2_X1 U11946 ( .A1(n18258), .A2(n9814), .ZN(n18250) );
  INV_X1 U11947 ( .A(n9815), .ZN(n9814) );
  OAI21_X1 U11948 ( .B1(n18386), .B2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n9816), .ZN(n9815) );
  AOI21_X1 U11949 ( .B1(n19002), .B2(n18249), .A(n9817), .ZN(n9816) );
  AND2_X1 U11950 ( .A1(n9868), .A2(n9867), .ZN(n12484) );
  NAND2_X1 U11951 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n9867) );
  NAND2_X1 U11952 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n9868) );
  AOI21_X1 U11953 ( .B1(n12507), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A(n9794), .ZN(n12398) );
  AND2_X1 U11954 ( .A1(n9870), .A2(n9869), .ZN(n12098) );
  NAND2_X1 U11955 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n9869) );
  NAND2_X1 U11956 ( .A1(n12508), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n9870) );
  OAI22_X1 U11957 ( .A1(n10429), .A2(n19576), .B1(n19664), .B2(n13054), .ZN(
        n10430) );
  OAI22_X1 U11958 ( .A1(n10487), .A2(n13060), .B1(n11513), .B2(n10486), .ZN(
        n10420) );
  OAI21_X1 U11959 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n10935), .A(
        n11168), .ZN(n11169) );
  OR2_X1 U11960 ( .A1(n11172), .A2(n11173), .ZN(n11168) );
  AOI21_X1 U11961 ( .B1(n9866), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A(n9804), 
        .ZN(n12451) );
  AOI21_X1 U11962 ( .B1(n12508), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n9801), .ZN(n12379) );
  AOI21_X1 U11963 ( .B1(n12548), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A(
        n9802), .ZN(n12362) );
  AOI21_X1 U11964 ( .B1(n9866), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A(n9803), 
        .ZN(n12326) );
  AOI21_X1 U11965 ( .B1(n12396), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A(n9791), .ZN(n12286) );
  AOI21_X1 U11966 ( .B1(n12526), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A(n9792), .ZN(n12272) );
  AOI21_X1 U11967 ( .B1(n12235), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A(n9793), .ZN(n12256) );
  BUF_X1 U11968 ( .A(n11861), .Z(n12467) );
  INV_X1 U11969 ( .A(n11964), .ZN(n11978) );
  OR3_X1 U11970 ( .A1(n12610), .A2(n12609), .A3(n12608), .ZN(n12611) );
  AND2_X1 U11971 ( .A1(n10620), .A2(n10619), .ZN(n10629) );
  OR2_X1 U11972 ( .A1(n11294), .A2(n10634), .ZN(n10620) );
  OAI211_X1 U11973 ( .C1(n15593), .C2(n10027), .A(n10026), .B(n13028), .ZN(
        n13052) );
  OR2_X1 U11974 ( .A1(n15584), .A2(n15594), .ZN(n10027) );
  NAND2_X1 U11975 ( .A1(n9843), .A2(n10557), .ZN(n10576) );
  INV_X1 U11976 ( .A(n10580), .ZN(n10458) );
  NAND2_X1 U11977 ( .A1(n10267), .A2(n19522), .ZN(n10240) );
  NAND2_X1 U11978 ( .A1(n11350), .A2(n10249), .ZN(n10235) );
  NAND2_X1 U11979 ( .A1(n11048), .A2(n11203), .ZN(n11049) );
  INV_X1 U11980 ( .A(n14853), .ZN(n13576) );
  AND2_X1 U11981 ( .A1(n12581), .A2(n12580), .ZN(n12617) );
  NAND2_X1 U11982 ( .A1(n9719), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11849) );
  NOR2_X1 U11983 ( .A1(n10051), .A2(n10048), .ZN(n10047) );
  INV_X1 U11984 ( .A(n10049), .ZN(n10048) );
  INV_X1 U11985 ( .A(n13331), .ZN(n10051) );
  NOR2_X1 U11986 ( .A1(n14870), .A2(n10050), .ZN(n10049) );
  INV_X1 U11987 ( .A(n14882), .ZN(n10050) );
  NAND2_X1 U11988 ( .A1(n14904), .A2(n14906), .ZN(n14893) );
  AND2_X1 U11989 ( .A1(n12395), .A2(n12373), .ZN(n10054) );
  AND2_X1 U11990 ( .A1(n10043), .A2(n9797), .ZN(n10042) );
  OR2_X1 U11991 ( .A1(n9783), .A2(n10044), .ZN(n10043) );
  NAND2_X1 U11992 ( .A1(n15449), .A2(n14728), .ZN(n9844) );
  OR2_X1 U11993 ( .A1(n15449), .A2(n16393), .ZN(n15248) );
  NOR2_X1 U11994 ( .A1(n14534), .A2(n9878), .ZN(n9877) );
  INV_X1 U11995 ( .A(n9879), .ZN(n9878) );
  NOR2_X1 U11996 ( .A1(n9881), .A2(n9880), .ZN(n9879) );
  INV_X1 U11997 ( .A(n14493), .ZN(n9880) );
  NOR2_X1 U11998 ( .A1(n14558), .A2(n14557), .ZN(n14551) );
  NAND2_X1 U11999 ( .A1(n9856), .A2(n12112), .ZN(n12128) );
  AND2_X1 U12000 ( .A1(n12130), .A2(n12112), .ZN(n9855) );
  INV_X1 U12001 ( .A(n14062), .ZN(n9873) );
  NAND2_X1 U12002 ( .A1(n12637), .A2(n14857), .ZN(n12727) );
  AND2_X1 U12003 ( .A1(n12775), .A2(n12774), .ZN(n13546) );
  OR2_X1 U12004 ( .A1(n11937), .A2(n11936), .ZN(n13238) );
  OR2_X1 U12005 ( .A1(n11926), .A2(n11925), .ZN(n13300) );
  OR2_X1 U12006 ( .A1(n11956), .A2(n11955), .ZN(n13239) );
  XNOR2_X1 U12007 ( .A(n12005), .B(n12004), .ZN(n12034) );
  NAND2_X1 U12008 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11874) );
  NAND2_X1 U12009 ( .A1(n11885), .A2(n13678), .ZN(n11882) );
  AOI21_X1 U12010 ( .B1(n11979), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11980), .ZN(n11989) );
  AOI21_X1 U12011 ( .B1(n21022), .B2(n16467), .A(n13882), .ZN(n14105) );
  INV_X1 U12012 ( .A(n13236), .ZN(n14232) );
  INV_X1 U12013 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20532) );
  AOI21_X1 U12014 ( .B1(n12581), .B2(n12579), .A(n12580), .ZN(n12591) );
  NAND2_X1 U12015 ( .A1(n12619), .A2(n13291), .ZN(n12615) );
  NOR2_X1 U12016 ( .A1(n10632), .A2(n10622), .ZN(n10623) );
  INV_X1 U12017 ( .A(n10631), .ZN(n10622) );
  NAND2_X1 U12018 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20202), .ZN(
        n10634) );
  NAND2_X1 U12019 ( .A1(n10773), .A2(n10914), .ZN(n10919) );
  NAND2_X1 U12020 ( .A1(n10764), .A2(n10763), .ZN(n10783) );
  NAND2_X1 U12021 ( .A1(n19551), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10763) );
  OR2_X1 U12022 ( .A1(n10762), .A2(n19551), .ZN(n10764) );
  NOR2_X1 U12023 ( .A1(n10233), .A2(n10232), .ZN(n10280) );
  NOR2_X1 U12024 ( .A1(n10284), .A2(n14308), .ZN(n10233) );
  INV_X1 U12025 ( .A(n15668), .ZN(n9892) );
  NAND2_X1 U12026 ( .A1(n15520), .A2(n9808), .ZN(n9811) );
  NOR2_X1 U12027 ( .A1(n15813), .A2(n9809), .ZN(n9808) );
  AND2_X1 U12028 ( .A1(n10413), .A2(n10412), .ZN(n10643) );
  NAND2_X1 U12029 ( .A1(n15714), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9930) );
  INV_X1 U12030 ( .A(n11278), .ZN(n9925) );
  NAND2_X1 U12031 ( .A1(n15751), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15717) );
  AOI21_X1 U12032 ( .B1(n10905), .B2(n19551), .A(n10004), .ZN(n10003) );
  NAND2_X1 U12033 ( .A1(n10907), .A2(n10906), .ZN(n10004) );
  AND2_X1 U12034 ( .A1(n14070), .A2(n13989), .ZN(n9958) );
  INV_X1 U12035 ( .A(n10606), .ZN(n10607) );
  NAND2_X1 U12036 ( .A1(n14450), .A2(n11431), .ZN(n13670) );
  XNOR2_X1 U12037 ( .A(n10599), .B(n9760), .ZN(n10600) );
  NAND2_X1 U12038 ( .A1(n10251), .A2(n19543), .ZN(n10252) );
  INV_X1 U12039 ( .A(n13172), .ZN(n10251) );
  NOR2_X1 U12040 ( .A1(n13627), .A2(n11405), .ZN(n11408) );
  NAND2_X1 U12041 ( .A1(n10453), .A2(n10452), .ZN(n11416) );
  NOR2_X1 U12042 ( .A1(n10329), .A2(n10350), .ZN(n19749) );
  NAND2_X1 U12043 ( .A1(n10113), .A2(n10352), .ZN(n19876) );
  NAND2_X1 U12044 ( .A1(n20183), .A2(n20022), .ZN(n19520) );
  NAND2_X2 U12045 ( .A1(n10140), .A2(n10139), .ZN(n11354) );
  INV_X1 U12046 ( .A(n18981), .ZN(n11233) );
  INV_X1 U12047 ( .A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17492) );
  AND2_X1 U12048 ( .A1(n9819), .A2(n9786), .ZN(n11221) );
  INV_X1 U12049 ( .A(n9991), .ZN(n9990) );
  OR2_X1 U12050 ( .A1(n18144), .A2(n11215), .ZN(n9818) );
  INV_X1 U12051 ( .A(n16278), .ZN(n19003) );
  OAI211_X1 U12052 ( .C1(n10949), .C2(n17419), .A(n11107), .B(n11106), .ZN(
        n11143) );
  AOI211_X1 U12053 ( .C1(n17512), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n11105), .B(n11104), .ZN(n11106) );
  INV_X1 U12054 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n16334) );
  INV_X1 U12055 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20260) );
  AND2_X1 U12056 ( .A1(n14148), .A2(n11877), .ZN(n14093) );
  NAND2_X1 U12057 ( .A1(n15116), .A2(n14094), .ZN(n14700) );
  AND2_X1 U12058 ( .A1(n13584), .A2(n13688), .ZN(n20352) );
  AND2_X1 U12059 ( .A1(n12006), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12566) );
  AND2_X1 U12060 ( .A1(n14881), .A2(n10045), .ZN(n12766) );
  AND2_X1 U12061 ( .A1(n10047), .A2(n10046), .ZN(n10045) );
  INV_X1 U12062 ( .A(n12767), .ZN(n10046) );
  OR2_X1 U12063 ( .A1(n12498), .A2(n15143), .ZN(n12499) );
  OR2_X1 U12064 ( .A1(n12499), .A2(n14873), .ZN(n12540) );
  NOR2_X1 U12065 ( .A1(n12461), .A2(n15165), .ZN(n12462) );
  NAND2_X1 U12066 ( .A1(n12462), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12498) );
  INV_X1 U12067 ( .A(n12422), .ZN(n12423) );
  OR2_X1 U12068 ( .A1(n12424), .A2(n14921), .ZN(n12461) );
  CLKBUF_X1 U12069 ( .A(n14904), .Z(n14905) );
  INV_X1 U12070 ( .A(n12374), .ZN(n12375) );
  NAND2_X1 U12071 ( .A1(n12352), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12353) );
  INV_X1 U12072 ( .A(n12351), .ZN(n12352) );
  INV_X1 U12073 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n14978) );
  OR2_X1 U12074 ( .A1(n15209), .A2(n12631), .ZN(n12355) );
  AND2_X1 U12075 ( .A1(n12336), .A2(n12335), .ZN(n14987) );
  AND2_X1 U12076 ( .A1(n12314), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12315) );
  INV_X1 U12077 ( .A(n12313), .ZN(n12314) );
  NAND2_X1 U12078 ( .A1(n10037), .A2(n12320), .ZN(n10036) );
  INV_X1 U12079 ( .A(n10039), .ZN(n10037) );
  NOR2_X1 U12080 ( .A1(n12281), .A2(n16301), .ZN(n12282) );
  INV_X1 U12081 ( .A(n14583), .ZN(n10038) );
  NAND2_X1 U12082 ( .A1(n12250), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12281) );
  NOR2_X1 U12083 ( .A1(n12234), .A2(n16321), .ZN(n12250) );
  OR2_X1 U12084 ( .A1(n12218), .A2(n16334), .ZN(n12234) );
  AND2_X1 U12085 ( .A1(n12189), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12190) );
  NOR2_X1 U12086 ( .A1(n12154), .A2(n20260), .ZN(n12189) );
  OR2_X1 U12087 ( .A1(n14404), .A2(n14405), .ZN(n14427) );
  NAND2_X1 U12088 ( .A1(n12134), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12170) );
  INV_X1 U12089 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12107) );
  NOR2_X1 U12090 ( .A1(n12105), .A2(n12107), .ZN(n12123) );
  AND2_X1 U12091 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n12058), .ZN(
        n12084) );
  NAND2_X1 U12092 ( .A1(n14689), .A2(n12783), .ZN(n12741) );
  INV_X1 U12093 ( .A(n10069), .ZN(n14708) );
  NAND2_X1 U12094 ( .A1(n10075), .A2(n15288), .ZN(n9848) );
  AND2_X1 U12095 ( .A1(n14919), .A2(n14913), .ZN(n14911) );
  AND2_X1 U12096 ( .A1(n12721), .A2(n12720), .ZN(n14920) );
  OR2_X1 U12097 ( .A1(n14931), .A2(n12716), .ZN(n14933) );
  NAND2_X1 U12098 ( .A1(n14587), .A2(n9884), .ZN(n15035) );
  NAND2_X1 U12099 ( .A1(n14587), .A2(n12696), .ZN(n15046) );
  INV_X1 U12100 ( .A(n15248), .ZN(n15249) );
  NOR2_X1 U12101 ( .A1(n15262), .A2(n15264), .ZN(n15445) );
  NAND2_X1 U12102 ( .A1(n9738), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15447) );
  NAND2_X1 U12103 ( .A1(n14551), .A2(n9879), .ZN(n14535) );
  AND2_X1 U12104 ( .A1(n9773), .A2(n13304), .ZN(n10080) );
  NAND2_X1 U12105 ( .A1(n9863), .A2(n9861), .ZN(n14431) );
  NOR2_X1 U12106 ( .A1(n12671), .A2(n9862), .ZN(n9861) );
  INV_X1 U12107 ( .A(n9864), .ZN(n9862) );
  AOI21_X1 U12108 ( .B1(n13285), .B2(n10079), .A(n9765), .ZN(n10078) );
  OR2_X1 U12109 ( .A1(n20464), .A2(n20465), .ZN(n16424) );
  NOR2_X1 U12110 ( .A1(n13903), .A2(n13904), .ZN(n14063) );
  NOR2_X1 U12111 ( .A1(n16404), .A2(n14725), .ZN(n15479) );
  AND2_X1 U12112 ( .A1(n12644), .A2(n12643), .ZN(n13828) );
  NAND2_X1 U12113 ( .A1(n13828), .A2(n13827), .ZN(n13904) );
  AND2_X1 U12114 ( .A1(n20455), .A2(n20475), .ZN(n14725) );
  NAND2_X1 U12115 ( .A1(n13703), .A2(n13698), .ZN(n20428) );
  AND2_X1 U12116 ( .A1(n12642), .A2(n12641), .ZN(n13810) );
  AND2_X1 U12117 ( .A1(n12637), .A2(n12650), .ZN(n13811) );
  CLKBUF_X1 U12118 ( .A(n11824), .Z(n12432) );
  NAND2_X1 U12119 ( .A1(n13580), .A2(n13579), .ZN(n13877) );
  NOR2_X1 U12120 ( .A1(n11808), .A2(n11807), .ZN(n11809) );
  NOR2_X1 U12121 ( .A1(n13693), .A2(n14851), .ZN(n16235) );
  NAND2_X1 U12122 ( .A1(n10141), .A2(n11336), .ZN(n11352) );
  OR2_X1 U12123 ( .A1(n15533), .A2(n10756), .ZN(n14678) );
  NAND2_X1 U12124 ( .A1(n15531), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15533) );
  NOR2_X2 U12125 ( .A1(n15528), .A2(n16533), .ZN(n15527) );
  NAND2_X1 U12126 ( .A1(n9727), .A2(n9780), .ZN(n16210) );
  NAND2_X1 U12127 ( .A1(n16210), .A2(n16585), .ZN(n16209) );
  NAND2_X1 U12128 ( .A1(n10863), .A2(n9775), .ZN(n10836) );
  OR2_X1 U12129 ( .A1(n10839), .A2(n10769), .ZN(n10842) );
  NAND2_X1 U12130 ( .A1(n10771), .A2(n10770), .ZN(n10862) );
  INV_X1 U12131 ( .A(n10841), .ZN(n10770) );
  INV_X1 U12132 ( .A(n10842), .ZN(n10771) );
  NAND2_X1 U12133 ( .A1(n15520), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15519) );
  NAND2_X1 U12134 ( .A1(n19367), .A2(n10014), .ZN(n10850) );
  INV_X1 U12135 ( .A(n10007), .ZN(n10006) );
  NAND2_X1 U12136 ( .A1(n10813), .A2(n10007), .ZN(n10820) );
  AND2_X1 U12137 ( .A1(n12823), .A2(n9744), .ZN(n10032) );
  AND2_X1 U12138 ( .A1(n12822), .A2(n13849), .ZN(n13985) );
  INV_X1 U12139 ( .A(n11421), .ZN(n14823) );
  INV_X1 U12140 ( .A(n11644), .ZN(n11646) );
  NAND2_X1 U12141 ( .A1(n15536), .A2(n15537), .ZN(n15619) );
  XNOR2_X1 U12142 ( .A(n13077), .B(n13075), .ZN(n15569) );
  NAND2_X1 U12143 ( .A1(n15569), .A2(n15568), .ZN(n15567) );
  NOR2_X1 U12144 ( .A1(n10023), .A2(n10022), .ZN(n10021) );
  INV_X1 U12145 ( .A(n15612), .ZN(n10022) );
  INV_X1 U12146 ( .A(n10024), .ZN(n10023) );
  OR2_X1 U12147 ( .A1(n11525), .A2(n11524), .ZN(n13926) );
  INV_X1 U12148 ( .A(n10249), .ZN(n13176) );
  AND2_X1 U12149 ( .A1(n13408), .A2(n13407), .ZN(n14191) );
  INV_X1 U12150 ( .A(n13498), .ZN(n19521) );
  NAND2_X1 U12151 ( .A1(n9949), .A2(n15571), .ZN(n9948) );
  INV_X1 U12152 ( .A(n15597), .ZN(n9949) );
  NOR2_X1 U12153 ( .A1(n15522), .A2(n14670), .ZN(n15524) );
  NAND2_X1 U12154 ( .A1(n15523), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15522) );
  NOR2_X2 U12155 ( .A1(n15511), .A2(n15794), .ZN(n15523) );
  NAND2_X1 U12156 ( .A1(n14645), .A2(n9953), .ZN(n9952) );
  NOR2_X1 U12157 ( .A1(n14473), .A2(n14651), .ZN(n9953) );
  NOR2_X1 U12158 ( .A1(n15517), .A2(n16591), .ZN(n15520) );
  INV_X1 U12159 ( .A(n16005), .ZN(n15997) );
  NAND2_X1 U12160 ( .A1(n15518), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15517) );
  INV_X1 U12161 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15512) );
  NOR2_X1 U12162 ( .A1(n15515), .A2(n15512), .ZN(n15518) );
  NAND2_X1 U12163 ( .A1(n15516), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15515) );
  AND2_X1 U12164 ( .A1(n10693), .A2(n10692), .ZN(n13942) );
  AND2_X1 U12165 ( .A1(n10669), .A2(n10668), .ZN(n14456) );
  INV_X1 U12166 ( .A(n9924), .ZN(n9923) );
  AND2_X1 U12167 ( .A1(n14810), .A2(n14809), .ZN(n14811) );
  NOR2_X2 U12168 ( .A1(n15717), .A2(n15842), .ZN(n15718) );
  INV_X1 U12169 ( .A(n9939), .ZN(n9938) );
  AOI21_X1 U12170 ( .B1(n15860), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n9940), .ZN(n9939) );
  INV_X1 U12171 ( .A(n15840), .ZN(n9940) );
  NOR2_X1 U12172 ( .A1(n15737), .A2(n15746), .ZN(n10909) );
  AND2_X1 U12173 ( .A1(n15747), .A2(n10922), .ZN(n15711) );
  OR2_X1 U12174 ( .A1(n16505), .A2(n10781), .ZN(n15710) );
  XNOR2_X1 U12175 ( .A(n10920), .B(n15872), .ZN(n15737) );
  AND2_X1 U12176 ( .A1(n10908), .A2(n15884), .ZN(n15746) );
  NAND2_X1 U12177 ( .A1(n10003), .A2(n14818), .ZN(n10908) );
  OR3_X1 U12178 ( .A1(n16534), .A2(n10781), .A3(n15884), .ZN(n15747) );
  AOI21_X1 U12179 ( .B1(n15771), .B2(n9919), .A(n9763), .ZN(n9918) );
  INV_X1 U12180 ( .A(n15917), .ZN(n9919) );
  INV_X1 U12181 ( .A(n15771), .ZN(n9920) );
  NAND2_X1 U12182 ( .A1(n10894), .A2(n15917), .ZN(n15772) );
  NAND2_X1 U12183 ( .A1(n13229), .A2(n9746), .ZN(n15767) );
  OAI21_X1 U12184 ( .B1(n10870), .B2(n10781), .A(n13224), .ZN(n13215) );
  NOR2_X1 U12185 ( .A1(n13212), .A2(n13211), .ZN(n10056) );
  AND3_X1 U12186 ( .A1(n11615), .A2(n11614), .A3(n11613), .ZN(n14634) );
  OR2_X1 U12187 ( .A1(n9897), .A2(n14434), .ZN(n9896) );
  AND2_X1 U12188 ( .A1(n16015), .A2(n13203), .ZN(n10065) );
  NAND2_X1 U12189 ( .A1(n16002), .A2(n11655), .ZN(n16005) );
  NAND2_X1 U12190 ( .A1(n10877), .A2(n16007), .ZN(n16015) );
  NOR2_X1 U12191 ( .A1(n16040), .A2(n16695), .ZN(n16680) );
  AND2_X1 U12192 ( .A1(n13943), .A2(n9958), .ZN(n14301) );
  AND2_X1 U12193 ( .A1(n10835), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16024) );
  AND2_X1 U12194 ( .A1(n11372), .A2(n16693), .ZN(n16028) );
  AND4_X1 U12195 ( .A1(n11545), .A2(n11544), .A3(n11543), .A4(n11542), .ZN(
        n16021) );
  CLKBUF_X1 U12196 ( .A(n16002), .Z(n16003) );
  NAND2_X1 U12197 ( .A1(n9906), .A2(n9905), .ZN(n9904) );
  INV_X1 U12198 ( .A(n13888), .ZN(n9905) );
  NAND2_X1 U12199 ( .A1(n9943), .A2(n13931), .ZN(n9942) );
  INV_X1 U12200 ( .A(n9944), .ZN(n9943) );
  INV_X1 U12201 ( .A(n13722), .ZN(n9903) );
  AND2_X1 U12202 ( .A1(n10677), .A2(n10676), .ZN(n13831) );
  INV_X1 U12203 ( .A(n10575), .ZN(n10578) );
  INV_X1 U12204 ( .A(n14449), .ZN(n9980) );
  AND4_X1 U12205 ( .A1(n11425), .A2(n11424), .A3(n11423), .A4(n11422), .ZN(
        n14219) );
  AOI21_X1 U12206 ( .B1(n14288), .B2(n14818), .A(n14453), .ZN(n9911) );
  INV_X1 U12207 ( .A(n10795), .ZN(n10796) );
  AND2_X1 U12208 ( .A1(n10308), .A2(n10658), .ZN(n10660) );
  AND2_X1 U12209 ( .A1(n13528), .A2(n13527), .ZN(n14046) );
  INV_X1 U12210 ( .A(n19636), .ZN(n19630) );
  AND2_X1 U12211 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19979), .ZN(
        n12810) );
  OR2_X1 U12212 ( .A1(n20167), .A2(n19779), .ZN(n19978) );
  NOR2_X2 U12213 ( .A1(n19519), .A2(n19520), .ZN(n19563) );
  OR2_X1 U12214 ( .A1(n20178), .A2(n19513), .ZN(n20020) );
  NAND2_X1 U12215 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n20022), .ZN(n19564) );
  INV_X1 U12216 ( .A(n20221), .ZN(n20215) );
  NOR2_X1 U12217 ( .A1(n18991), .A2(n13364), .ZN(n18969) );
  AND2_X1 U12218 ( .A1(n9828), .A2(n9724), .ZN(n13391) );
  OR2_X1 U12219 ( .A1(n16944), .A2(n16938), .ZN(n9828) );
  NAND2_X1 U12220 ( .A1(n9822), .A2(n9821), .ZN(n9823) );
  AOI21_X1 U12221 ( .B1(n9724), .B2(n17933), .A(n16970), .ZN(n9821) );
  NAND2_X1 U12222 ( .A1(n13362), .A2(n9724), .ZN(n9822) );
  OR2_X1 U12223 ( .A1(n13362), .A2(n17933), .ZN(n9824) );
  NAND2_X1 U12224 ( .A1(n17338), .A2(P3_EBX_REG_19__SCAN_IN), .ZN(n17225) );
  NAND2_X1 U12225 ( .A1(n17415), .A2(P3_EBX_REG_15__SCAN_IN), .ZN(n17384) );
  NOR2_X1 U12226 ( .A1(n11140), .A2(n11139), .ZN(n11141) );
  INV_X1 U12227 ( .A(n11137), .ZN(n11142) );
  AND2_X1 U12228 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11139) );
  INV_X1 U12229 ( .A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17412) );
  CLKBUF_X1 U12230 ( .A(n16111), .Z(n17460) );
  INV_X1 U12231 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17452) );
  CLKBUF_X1 U12232 ( .A(n10948), .Z(n17474) );
  NAND2_X1 U12233 ( .A1(n17567), .A2(n18542), .ZN(n16278) );
  AOI211_X1 U12234 ( .C1(n17512), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n11115), .B(n11114), .ZN(n11116) );
  NOR2_X1 U12235 ( .A1(n17764), .A2(n17726), .ZN(n17745) );
  INV_X1 U12236 ( .A(n13379), .ZN(n16876) );
  NOR2_X1 U12237 ( .A1(n17942), .A2(n9830), .ZN(n9829) );
  INV_X1 U12238 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9830) );
  NOR2_X1 U12239 ( .A1(n16199), .A2(n16258), .ZN(n16739) );
  NOR2_X1 U12240 ( .A1(n16258), .A2(n18190), .ZN(n16738) );
  NAND2_X1 U12241 ( .A1(n17836), .A2(n10086), .ZN(n11687) );
  NAND2_X1 U12242 ( .A1(n11734), .A2(n18241), .ZN(n18190) );
  INV_X1 U12243 ( .A(n17876), .ZN(n11068) );
  NAND2_X1 U12244 ( .A1(n17877), .A2(n17881), .ZN(n17876) );
  NOR2_X1 U12245 ( .A1(n17921), .A2(n11258), .ZN(n17882) );
  OAI21_X1 U12246 ( .B1(n18469), .B2(n18259), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n9817) );
  NOR2_X1 U12247 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17922), .ZN(
        n17900) );
  INV_X1 U12248 ( .A(n18313), .ZN(n18242) );
  INV_X1 U12249 ( .A(n18312), .ZN(n18241) );
  NOR2_X1 U12250 ( .A1(n11060), .A2(n11061), .ZN(n17973) );
  INV_X1 U12251 ( .A(n11665), .ZN(n18280) );
  OR2_X1 U12252 ( .A1(n18088), .A2(n11231), .ZN(n18011) );
  AND2_X1 U12253 ( .A1(n9754), .A2(n18333), .ZN(n9995) );
  AOI21_X1 U12254 ( .B1(n11250), .B2(n11254), .A(n11249), .ZN(n18980) );
  INV_X1 U12255 ( .A(n11247), .ZN(n18993) );
  NAND2_X1 U12256 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18079), .ZN(
        n18370) );
  INV_X1 U12257 ( .A(n18011), .ZN(n18372) );
  INV_X1 U12258 ( .A(n18029), .ZN(n17990) );
  INV_X1 U12259 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18278) );
  NOR2_X1 U12260 ( .A1(n9820), .A2(n11228), .ZN(n18089) );
  AND2_X1 U12261 ( .A1(n11229), .A2(n11230), .ZN(n9820) );
  NOR2_X1 U12262 ( .A1(n18089), .A2(n18278), .ZN(n18088) );
  NAND2_X1 U12263 ( .A1(n18414), .A2(n18080), .ZN(n18079) );
  XNOR2_X1 U12264 ( .A(n11221), .B(n11222), .ZN(n18107) );
  NOR2_X1 U12265 ( .A1(n18107), .A2(n18433), .ZN(n18106) );
  XNOR2_X1 U12266 ( .A(n9818), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18135) );
  NOR2_X1 U12267 ( .A1(n11212), .A2(n11213), .ZN(n18146) );
  NOR2_X1 U12268 ( .A1(n18146), .A2(n18145), .ZN(n18144) );
  NOR2_X1 U12269 ( .A1(n11200), .A2(n11190), .ZN(n11732) );
  OAI21_X1 U12270 ( .B1(n11177), .B2(n11193), .A(n11194), .ZN(n11181) );
  AOI21_X1 U12271 ( .B1(n11197), .B2(n11196), .A(n11195), .ZN(n18967) );
  NOR2_X1 U12272 ( .A1(n13363), .A2(n18993), .ZN(n18991) );
  INV_X1 U12273 ( .A(n18991), .ZN(n14657) );
  AND2_X1 U12274 ( .A1(n11162), .A2(n9962), .ZN(n18529) );
  NOR2_X1 U12275 ( .A1(n9966), .A2(n9963), .ZN(n9962) );
  INV_X1 U12276 ( .A(n17567), .ZN(n18538) );
  INV_X1 U12277 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n19039) );
  OR2_X1 U12278 ( .A1(n13468), .A2(n14081), .ZN(n13457) );
  NAND2_X1 U12279 ( .A1(n13457), .A2(n13660), .ZN(n21025) );
  INV_X1 U12280 ( .A(n20323), .ZN(n20335) );
  AND2_X1 U12281 ( .A1(n20334), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20323) );
  INV_X1 U12282 ( .A(n20340), .ZN(n20321) );
  AND2_X1 U12283 ( .A1(n12757), .A2(n12745), .ZN(n20320) );
  XNOR2_X1 U12284 ( .A(n12643), .B(n13810), .ZN(n20350) );
  INV_X1 U12285 ( .A(n20320), .ZN(n20351) );
  NAND2_X1 U12286 ( .A1(n12779), .A2(n14860), .ZN(n15037) );
  INV_X1 U12287 ( .A(n15037), .ZN(n15047) );
  OR2_X1 U12288 ( .A1(n15037), .A2(n11877), .ZN(n15048) );
  AOI21_X1 U12289 ( .B1(n14083), .B2(n14082), .A(n14081), .ZN(n14090) );
  AOI21_X1 U12290 ( .B1(n14088), .B2(n14087), .A(n14086), .ZN(n14089) );
  INV_X2 U12291 ( .A(n15115), .ZN(n15113) );
  CLKBUF_X1 U12292 ( .A(n20373), .Z(n21028) );
  XNOR2_X1 U12293 ( .A(n12571), .B(n12758), .ZN(n14737) );
  NAND2_X1 U12294 ( .A1(n12765), .A2(n13332), .ZN(n14686) );
  OR2_X1 U12295 ( .A1(n13330), .A2(n13331), .ZN(n13332) );
  INV_X1 U12296 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16301) );
  AND2_X1 U12297 ( .A1(n14404), .A2(n14358), .ZN(n20278) );
  INV_X1 U12298 ( .A(n15254), .ZN(n20416) );
  AND2_X1 U12299 ( .A1(n16235), .A2(n14860), .ZN(n20422) );
  XNOR2_X1 U12300 ( .A(n9860), .B(n12783), .ZN(n15285) );
  INV_X1 U12301 ( .A(n12782), .ZN(n9860) );
  INV_X1 U12302 ( .A(n14871), .ZN(n12781) );
  OR2_X1 U12303 ( .A1(n15424), .A2(n14730), .ZN(n15357) );
  OAI21_X1 U12304 ( .B1(n15194), .B2(n14728), .A(n15449), .ZN(n15187) );
  INV_X1 U12305 ( .A(n16446), .ZN(n15474) );
  NOR2_X1 U12306 ( .A1(n14284), .A2(n12663), .ZN(n14383) );
  INV_X1 U12307 ( .A(n20470), .ZN(n20452) );
  AND2_X1 U12308 ( .A1(n13703), .A2(n13701), .ZN(n20466) );
  INV_X1 U12309 ( .A(n20428), .ZN(n20467) );
  INV_X1 U12310 ( .A(n20432), .ZN(n20473) );
  NAND2_X1 U12311 ( .A1(n12013), .A2(n12012), .ZN(n12014) );
  INV_X1 U12312 ( .A(n13237), .ZN(n12013) );
  NAND2_X1 U12313 ( .A1(n12036), .A2(n11991), .ZN(n13542) );
  INV_X1 U12314 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20768) );
  INV_X1 U12315 ( .A(n16251), .ZN(n13882) );
  NOR2_X1 U12316 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n15498) );
  NOR2_X1 U12317 ( .A1(n12036), .A2(n14233), .ZN(n13876) );
  INV_X1 U12318 ( .A(n20511), .ZN(n20526) );
  OAI21_X1 U12319 ( .B1(n20639), .B2(n20623), .A(n20847), .ZN(n20641) );
  OAI21_X1 U12320 ( .B1(n20682), .B2(n20681), .A(n20680), .ZN(n20700) );
  OAI211_X1 U12321 ( .C1(n20774), .C2(n20728), .A(n20712), .B(n20773), .ZN(
        n20730) );
  INV_X1 U12322 ( .A(n20778), .ZN(n20801) );
  NOR2_X2 U12323 ( .A1(n20812), .A2(n20739), .ZN(n20800) );
  OAI21_X1 U12324 ( .B1(n20817), .B2(n20816), .A(n20815), .ZN(n20835) );
  INV_X1 U12325 ( .A(n20838), .ZN(n14545) );
  AOI22_X1 U12326 ( .A1(n14504), .A2(n14501), .B1(n20706), .B2(n20674), .ZN(
        n14547) );
  OAI211_X1 U12327 ( .C1(n20848), .C2(n20870), .A(n20847), .B(n20846), .ZN(
        n20872) );
  NOR2_X2 U12328 ( .A1(n20885), .A2(n20739), .ZN(n20871) );
  AND2_X1 U12329 ( .A1(n15081), .A2(n14117), .ZN(n20923) );
  INV_X1 U12330 ( .A(n20929), .ZN(n20936) );
  OR2_X1 U12331 ( .A1(n20885), .A2(n20579), .ZN(n20940) );
  NAND2_X1 U12332 ( .A1(n13682), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16251) );
  AND2_X1 U12333 ( .A1(n20942), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16248) );
  INV_X1 U12334 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20774) );
  CLKBUF_X1 U12335 ( .A(n11352), .Z(n11353) );
  AND2_X1 U12336 ( .A1(n10641), .A2(n10640), .ZN(n20208) );
  NAND2_X1 U12337 ( .A1(n16495), .A2(n19384), .ZN(n16484) );
  NAND2_X1 U12338 ( .A1(n15534), .A2(n15721), .ZN(n16469) );
  NAND2_X1 U12339 ( .A1(n16524), .A2(n19384), .ZN(n16512) );
  NAND2_X1 U12340 ( .A1(n16525), .A2(n16526), .ZN(n16524) );
  NAND2_X1 U12341 ( .A1(n16538), .A2(n19384), .ZN(n16525) );
  AND2_X1 U12342 ( .A1(n14816), .A2(n10903), .ZN(n16520) );
  NAND2_X1 U12343 ( .A1(n16209), .A2(n9728), .ZN(n16565) );
  AND2_X1 U12344 ( .A1(n14195), .A2(n14192), .ZN(n19361) );
  NAND2_X1 U12345 ( .A1(n19417), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19397) );
  INV_X1 U12346 ( .A(n19397), .ZN(n19431) );
  NAND2_X1 U12347 ( .A1(n10778), .A2(n10001), .ZN(n19435) );
  INV_X1 U12348 ( .A(n19411), .ZN(n19443) );
  INV_X1 U12349 ( .A(n19361), .ZN(n19447) );
  INV_X1 U12350 ( .A(n19422), .ZN(n19441) );
  AND2_X1 U12351 ( .A1(n11474), .A2(n11473), .ZN(n13909) );
  INV_X1 U12352 ( .A(n14786), .ZN(n15618) );
  AND2_X1 U12353 ( .A1(n15616), .A2(n13338), .ZN(n14786) );
  XNOR2_X1 U12354 ( .A(n13171), .B(n13170), .ZN(n13339) );
  NAND2_X1 U12355 ( .A1(n10020), .A2(n10019), .ZN(n13171) );
  NOR3_X1 U12356 ( .A1(n15673), .A2(n9891), .A3(n15674), .ZN(n15650) );
  NAND2_X1 U12357 ( .A1(n13004), .A2(n13002), .ZN(n10028) );
  INV_X1 U12358 ( .A(n15692), .ZN(n19450) );
  AND2_X1 U12359 ( .A1(n15675), .A2(n19465), .ZN(n19471) );
  INV_X1 U12360 ( .A(n15675), .ZN(n19449) );
  OR2_X1 U12361 ( .A1(n13524), .A2(n13174), .ZN(n13175) );
  INV_X1 U12362 ( .A(n14356), .ZN(n19464) );
  NOR2_X1 U12363 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16270), .ZN(n13737) );
  BUF_X1 U12364 ( .A(n19484), .Z(n19496) );
  INV_X1 U12365 ( .A(n20214), .ZN(n19497) );
  AND2_X1 U12366 ( .A1(n14191), .A2(n9730), .ZN(n14195) );
  AOI21_X1 U12367 ( .B1(n14191), .B2(n20221), .A(n14195), .ZN(n13483) );
  CLKBUF_X1 U12368 ( .A(n13483), .Z(n13517) );
  INV_X1 U12369 ( .A(n14835), .ZN(n10748) );
  INV_X1 U12370 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19381) );
  INV_X1 U12371 ( .A(n16667), .ZN(n19510) );
  NAND2_X1 U12372 ( .A1(n19212), .A2(n10750), .ZN(n16677) );
  OR2_X1 U12373 ( .A1(n19212), .A2(n15586), .ZN(n16668) );
  XNOR2_X1 U12374 ( .A(n11287), .B(n10082), .ZN(n14685) );
  NAND2_X1 U12375 ( .A1(n11279), .A2(n11278), .ZN(n14813) );
  NAND2_X1 U12376 ( .A1(n15772), .A2(n15771), .ZN(n15909) );
  NAND2_X1 U12377 ( .A1(n9840), .A2(n9839), .ZN(n9838) );
  NAND2_X1 U12378 ( .A1(n15967), .A2(n15966), .ZN(n9839) );
  NAND2_X1 U12379 ( .A1(n13206), .A2(n15988), .ZN(n15820) );
  AND2_X1 U12380 ( .A1(n10598), .A2(n10597), .ZN(n14447) );
  AND2_X1 U12381 ( .A1(n11388), .A2(n11387), .ZN(n16710) );
  INV_X1 U12382 ( .A(n16716), .ZN(n16699) );
  NAND2_X1 U12383 ( .A1(n13622), .A2(n13621), .ZN(n20197) );
  NAND2_X1 U12384 ( .A1(n13638), .A2(n13637), .ZN(n20190) );
  INV_X1 U12385 ( .A(n20190), .ZN(n19513) );
  XNOR2_X1 U12386 ( .A(n13640), .B(n13641), .ZN(n20178) );
  INV_X1 U12387 ( .A(n14314), .ZN(n20162) );
  AND2_X1 U12388 ( .A1(n19518), .A2(n19517), .ZN(n19539) );
  INV_X1 U12389 ( .A(n19539), .ZN(n19569) );
  INV_X1 U12390 ( .A(n19661), .ZN(n19652) );
  OR2_X1 U12391 ( .A1(n19719), .A2(n19871), .ZN(n19661) );
  OAI21_X1 U12392 ( .B1(n19639), .B2(n19638), .A(n19637), .ZN(n19657) );
  INV_X1 U12393 ( .A(n19670), .ZN(n19688) );
  AND2_X1 U12394 ( .A1(n19758), .A2(n20164), .ZN(n19687) );
  OR3_X1 U12395 ( .A1(n19727), .A2(n19947), .A3(n19726), .ZN(n19746) );
  NOR2_X1 U12396 ( .A1(n20020), .A2(n19719), .ZN(n19767) );
  NAND2_X1 U12397 ( .A1(n19788), .A2(n19787), .ZN(n19806) );
  INV_X1 U12398 ( .A(n19838), .ZN(n19829) );
  OAI21_X1 U12399 ( .B1(n19818), .B2(n19817), .A(n19816), .ZN(n19834) );
  NOR2_X1 U12400 ( .A1(n19941), .A2(n19871), .ZN(n19909) );
  INV_X1 U12401 ( .A(n20028), .ZN(n19914) );
  INV_X1 U12402 ( .A(n19909), .ZN(n19939) );
  NOR2_X2 U12403 ( .A1(n19978), .A2(n19940), .ZN(n19973) );
  NOR2_X1 U12404 ( .A1(n19946), .A2(n19945), .ZN(n19971) );
  INV_X1 U12405 ( .A(n19923), .ZN(n20036) );
  INV_X1 U12406 ( .A(n20002), .ZN(n20048) );
  OAI22_X1 U12407 ( .A1(n19550), .A2(n19555), .B1(n15681), .B2(n19557), .ZN(
        n20054) );
  INV_X1 U12408 ( .A(n20075), .ZN(n20061) );
  OAI22_X1 U12409 ( .A1(n19558), .A2(n19557), .B1(n19556), .B2(n19555), .ZN(
        n20060) );
  AND2_X1 U12410 ( .A1(n12810), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20067) );
  INV_X1 U12411 ( .A(n20064), .ZN(n20071) );
  OR2_X1 U12412 ( .A1(n19978), .A2(n20020), .ZN(n20075) );
  NAND2_X1 U12413 ( .A1(n14196), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19210) );
  INV_X1 U12414 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n20218) );
  OR2_X1 U12415 ( .A1(n14310), .A2(n20195), .ZN(n20161) );
  NAND2_X1 U12416 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20086), .ZN(n20234) );
  INV_X1 U12417 ( .A(n19202), .ZN(n19198) );
  NAND2_X1 U12418 ( .A1(n19180), .A2(n18970), .ZN(n17764) );
  NOR2_X1 U12419 ( .A1(n18969), .A2(n17764), .ZN(n19202) );
  AND2_X1 U12420 ( .A1(n16944), .A2(n9724), .ZN(n16937) );
  AND2_X1 U12421 ( .A1(n9824), .A2(n17205), .ZN(n16969) );
  NOR2_X1 U12422 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17011), .ZN(n16996) );
  NOR2_X1 U12423 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17034), .ZN(n17019) );
  INV_X1 U12424 ( .A(n17030), .ZN(n17022) );
  NOR3_X1 U12425 ( .A1(n17210), .A2(n19093), .A3(n17040), .ZN(n17033) );
  NOR2_X1 U12426 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17080), .ZN(n17061) );
  NOR2_X2 U12427 ( .A1(n19138), .A2(n17204), .ZN(n17192) );
  NOR2_X1 U12428 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17151), .ZN(n17134) );
  INV_X1 U12429 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17532) );
  INV_X1 U12430 ( .A(n17165), .ZN(n17210) );
  INV_X1 U12431 ( .A(n17219), .ZN(n17216) );
  OAI211_X1 U12432 ( .C1(n19041), .C2(n18795), .A(n17172), .B(n19198), .ZN(
        n17221) );
  NAND2_X1 U12433 ( .A1(n17289), .A2(P3_EBX_REG_25__SCAN_IN), .ZN(n17281) );
  AND2_X1 U12434 ( .A1(n17295), .A2(P3_EBX_REG_24__SCAN_IN), .ZN(n17289) );
  AND2_X1 U12435 ( .A1(n17290), .A2(n9971), .ZN(n17295) );
  NOR2_X1 U12436 ( .A1(n16096), .A2(n16963), .ZN(n9971) );
  NOR2_X1 U12437 ( .A1(n17225), .A2(n17691), .ZN(n17336) );
  NOR2_X1 U12438 ( .A1(n17369), .A2(n17365), .ZN(n17338) );
  NOR2_X1 U12439 ( .A1(n17400), .A2(n17384), .ZN(n17370) );
  NOR2_X1 U12440 ( .A1(n17486), .A2(n17489), .ZN(n17468) );
  NAND2_X1 U12441 ( .A1(n17468), .A2(P3_EBX_REG_11__SCAN_IN), .ZN(n17467) );
  NOR2_X1 U12442 ( .A1(n17121), .A2(n17507), .ZN(n17526) );
  INV_X1 U12443 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17537) );
  INV_X1 U12444 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17544) );
  NAND2_X1 U12445 ( .A1(n17727), .A2(n9968), .ZN(n9967) );
  INV_X1 U12446 ( .A(n16094), .ZN(n9968) );
  NOR2_X1 U12447 ( .A1(n17770), .A2(n17634), .ZN(n17635) );
  NOR2_X1 U12448 ( .A1(n17813), .A2(n17693), .ZN(n17688) );
  INV_X1 U12449 ( .A(n10945), .ZN(n17697) );
  NOR2_X1 U12450 ( .A1(n17803), .A2(n17707), .ZN(n17710) );
  AND2_X1 U12451 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10990) );
  NAND2_X1 U12452 ( .A1(n16278), .A2(n17684), .ZN(n17716) );
  NOR2_X1 U12453 ( .A1(n10973), .A2(n10972), .ZN(n10974) );
  NOR2_X1 U12454 ( .A1(n10969), .A2(n10968), .ZN(n10975) );
  NOR2_X1 U12455 ( .A1(n10966), .A2(n10965), .ZN(n10976) );
  INV_X1 U12456 ( .A(n17720), .ZN(n17690) );
  INV_X1 U12457 ( .A(n17716), .ZN(n17719) );
  CLKBUF_X1 U12458 ( .A(n17828), .Z(n17820) );
  OAI21_X1 U12459 ( .B1(n19186), .B2(n19187), .A(n17766), .ZN(n17828) );
  NAND2_X1 U12461 ( .A1(n18080), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9993) );
  NOR2_X1 U12462 ( .A1(n18080), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9994) );
  NAND2_X1 U12463 ( .A1(n18004), .A2(n18280), .ZN(n18313) );
  INV_X1 U12464 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18045) );
  INV_X1 U12465 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n18058) );
  NOR2_X1 U12466 ( .A1(n18118), .A2(n17976), .ZN(n18138) );
  AND2_X1 U12467 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10091) );
  INV_X1 U12468 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n18113) );
  INV_X1 U12469 ( .A(n17155), .ZN(n18132) );
  INV_X1 U12470 ( .A(n18150), .ZN(n18180) );
  XNOR2_X1 U12471 ( .A(n11688), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16204) );
  NAND2_X1 U12472 ( .A1(n11687), .A2(n11686), .ZN(n11688) );
  NOR2_X1 U12473 ( .A1(n18265), .A2(n18248), .ZN(n18258) );
  NOR2_X1 U12474 ( .A1(n18278), .A2(n18409), .ZN(n18347) );
  INV_X1 U12475 ( .A(n18482), .ZN(n18349) );
  OAI21_X2 U12476 ( .B1(n18981), .B2(n18993), .A(n18980), .ZN(n19002) );
  AND2_X1 U12477 ( .A1(n11055), .A2(n9996), .ZN(n18050) );
  INV_X1 U12478 ( .A(n18303), .ZN(n18386) );
  NAND2_X1 U12479 ( .A1(n11055), .A2(n10103), .ZN(n18055) );
  AND2_X1 U12480 ( .A1(n17990), .A2(n11255), .ZN(n18414) );
  NAND2_X1 U12481 ( .A1(n17692), .A2(n18487), .ZN(n18418) );
  INV_X1 U12482 ( .A(n18494), .ZN(n18429) );
  NAND2_X1 U12483 ( .A1(n9790), .A2(n18123), .ZN(n18122) );
  INV_X1 U12484 ( .A(n9819), .ZN(n18119) );
  NOR2_X1 U12485 ( .A1(n18156), .A2(n18155), .ZN(n18154) );
  INV_X1 U12486 ( .A(n18503), .ZN(n18487) );
  INV_X1 U12487 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19015) );
  INV_X1 U12488 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n19019) );
  AOI211_X1 U12489 ( .C1(n19180), .C2(n19001), .A(n18516), .B(n14661), .ZN(
        n19166) );
  NOR2_X1 U12490 ( .A1(n19039), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n19033) );
  INV_X1 U12491 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n19138) );
  AND2_X2 U12492 ( .A1(n13355), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14699)
         );
  CLKBUF_X1 U12493 ( .A(n16836), .Z(n16842) );
  NOR4_X1 U12494 ( .A1(n14733), .A2(n14732), .A3(n14735), .A4(n14731), .ZN(
        n14734) );
  OAI21_X1 U12495 ( .B1(n15291), .B2(n20470), .A(n9857), .ZN(P1_U3001) );
  INV_X1 U12496 ( .A(n9858), .ZN(n9857) );
  OAI21_X1 U12497 ( .B1(n15285), .B2(n20469), .A(n9859), .ZN(n9858) );
  NOR2_X1 U12498 ( .A1(n15289), .A2(n15290), .ZN(n9859) );
  NAND2_X1 U12499 ( .A1(n14842), .A2(n14841), .ZN(n14843) );
  OR2_X1 U12500 ( .A1(n15702), .A2(n16716), .ZN(n14841) );
  OAI21_X1 U12501 ( .B1(n15846), .B2(n16704), .A(n9933), .ZN(P2_U3017) );
  INV_X1 U12502 ( .A(n9935), .ZN(n9934) );
  OAI21_X1 U12503 ( .B1(n15854), .B2(n16704), .A(n9761), .ZN(P2_U3018) );
  AOI21_X1 U12504 ( .B1(n15860), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n9901), .ZN(n9900) );
  INV_X1 U12505 ( .A(n15851), .ZN(n9902) );
  OAI21_X1 U12506 ( .B1(n15976), .B2(n16704), .A(n9833), .ZN(P2_U3029) );
  NOR2_X1 U12507 ( .A1(n15975), .A2(n15974), .ZN(n9834) );
  OAI21_X1 U12508 ( .B1(n16887), .B2(n9800), .A(n9825), .ZN(P3_U2640) );
  NOR2_X1 U12509 ( .A1(n16883), .A2(n9826), .ZN(n9825) );
  NAND2_X1 U12510 ( .A1(n9960), .A2(n9959), .ZN(n17271) );
  NAND2_X1 U12511 ( .A1(n9961), .A2(n17268), .ZN(n9960) );
  OR2_X1 U12512 ( .A1(n17267), .A2(n17268), .ZN(n9959) );
  INV_X1 U12513 ( .A(n17290), .ZN(n17308) );
  AND2_X1 U12514 ( .A1(n11712), .A2(n11711), .ZN(n11713) );
  NOR2_X1 U12515 ( .A1(n10089), .A2(n11710), .ZN(n11711) );
  NAND2_X1 U12516 ( .A1(n11738), .A2(n11739), .ZN(n9984) );
  NOR2_X2 U12517 ( .A1(n18989), .A2(n10927), .ZN(n10961) );
  OR2_X1 U12518 ( .A1(n9991), .A2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n9736) );
  INV_X1 U12519 ( .A(n11632), .ZN(n14824) );
  AND2_X1 U12520 ( .A1(n10368), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9737) );
  INV_X1 U12521 ( .A(n15449), .ZN(n10075) );
  NOR2_X1 U12522 ( .A1(n14583), .A2(n10039), .ZN(n15004) );
  AND3_X1 U12523 ( .A1(n12187), .A2(n12188), .A3(n10042), .ZN(n14525) );
  AND3_X1 U12524 ( .A1(n12187), .A2(n12188), .A3(n12186), .ZN(n14486) );
  AND2_X1 U12525 ( .A1(n14953), .A2(n10054), .ZN(n14929) );
  AND4_X1 U12526 ( .A1(n11761), .A2(n11760), .A3(n11759), .A4(n11758), .ZN(
        n9739) );
  OR3_X1 U12527 ( .A1(n15596), .A2(n15597), .A3(n15588), .ZN(n9740) );
  AND2_X1 U12528 ( .A1(n10061), .A2(n13208), .ZN(n15809) );
  OR3_X1 U12529 ( .A1(n15673), .A2(n15674), .A3(n9892), .ZN(n9741) );
  NAND2_X1 U12530 ( .A1(n15641), .A2(n15642), .ZN(n15632) );
  NAND2_X1 U12531 ( .A1(n10556), .A2(n10555), .ZN(n10602) );
  AND2_X1 U12532 ( .A1(n9776), .A2(n14421), .ZN(n9742) );
  OR2_X1 U12533 ( .A1(n9992), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9743) );
  INV_X2 U12534 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10359) );
  INV_X2 U12535 ( .A(n10661), .ZN(n10654) );
  NAND2_X1 U12536 ( .A1(n9903), .A2(n9906), .ZN(n13759) );
  AND2_X1 U12537 ( .A1(n12875), .A2(n10024), .ZN(n14641) );
  NOR2_X1 U12538 ( .A1(n14158), .A2(n16009), .ZN(n14353) );
  INV_X1 U12539 ( .A(n10030), .ZN(n14335) );
  OR2_X1 U12540 ( .A1(n11583), .A2(n11582), .ZN(n9744) );
  INV_X1 U12541 ( .A(n10031), .ZN(n14298) );
  NOR2_X1 U12542 ( .A1(n15547), .A2(n15553), .ZN(n9745) );
  AND2_X1 U12543 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n9746) );
  AND2_X1 U12544 ( .A1(n10617), .A2(n11655), .ZN(n9747) );
  AND2_X2 U12545 ( .A1(n12976), .A2(n10369), .ZN(n10395) );
  OR2_X1 U12546 ( .A1(n14472), .A2(n9952), .ZN(n9748) );
  OR2_X1 U12547 ( .A1(n11415), .A2(n11414), .ZN(n9749) );
  OR2_X2 U12548 ( .A1(n10334), .A2(n10346), .ZN(n9750) );
  NAND2_X1 U12549 ( .A1(n16002), .A2(n9747), .ZN(n15782) );
  XNOR2_X1 U12550 ( .A(n12805), .B(n12803), .ZN(n13640) );
  XNOR2_X1 U12551 ( .A(n12033), .B(n12034), .ZN(n13246) );
  NAND2_X1 U12552 ( .A1(n14953), .A2(n10053), .ZN(n14917) );
  OR2_X1 U12553 ( .A1(n17717), .A2(n19145), .ZN(n9751) );
  INV_X1 U12554 ( .A(n12788), .ZN(n10352) );
  OR2_X1 U12555 ( .A1(n11070), .A2(n18080), .ZN(n9753) );
  INV_X1 U12556 ( .A(n17727), .ZN(n18517) );
  AND2_X1 U12557 ( .A1(n9996), .A2(n18052), .ZN(n9754) );
  OAI21_X1 U12558 ( .B1(n10894), .B2(n9920), .A(n9918), .ZN(n15758) );
  NAND2_X1 U12559 ( .A1(n16600), .A2(n13203), .ZN(n16014) );
  NAND2_X1 U12560 ( .A1(n12807), .A2(n12806), .ZN(n13740) );
  AND2_X1 U12561 ( .A1(n10813), .A2(n10812), .ZN(n10766) );
  INV_X1 U12562 ( .A(n13323), .ZN(n11885) );
  AND4_X1 U12563 ( .A1(n13210), .A2(n15988), .A3(n16015), .A4(n13203), .ZN(
        n9755) );
  OR2_X1 U12564 ( .A1(n14686), .A2(n15258), .ZN(n9756) );
  AOI21_X1 U12565 ( .B1(n15827), .B2(n10822), .A(n10821), .ZN(n16620) );
  NOR3_X1 U12566 ( .A1(n15596), .A2(n9950), .A3(n9948), .ZN(n15561) );
  NAND2_X1 U12567 ( .A1(n9733), .A2(n13467), .ZN(n10341) );
  NAND2_X1 U12568 ( .A1(n14953), .A2(n12373), .ZN(n9757) );
  NAND2_X1 U12569 ( .A1(n14827), .A2(n11647), .ZN(n13189) );
  NAND2_X1 U12570 ( .A1(n13219), .A2(n15603), .ZN(n15596) );
  OAI21_X1 U12571 ( .B1(n12738), .B2(P1_EBX_REG_1__SCAN_IN), .A(n12640), .ZN(
        n12643) );
  OR2_X1 U12572 ( .A1(n11027), .A2(n11039), .ZN(n9758) );
  AND2_X1 U12573 ( .A1(n10557), .A2(n10781), .ZN(n9759) );
  AND2_X1 U12574 ( .A1(n10517), .A2(n10516), .ZN(n9760) );
  AND3_X1 U12575 ( .A1(n9902), .A2(n9900), .A3(n9899), .ZN(n9761) );
  AND2_X1 U12576 ( .A1(n9844), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9762) );
  NOR2_X1 U12577 ( .A1(n10897), .A2(n15906), .ZN(n9763) );
  AND2_X1 U12578 ( .A1(n16375), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9765) );
  NAND2_X1 U12579 ( .A1(n19367), .A2(n10831), .ZN(n10833) );
  AND2_X1 U12580 ( .A1(n9931), .A2(n15711), .ZN(n9766) );
  INV_X1 U12581 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10016) );
  NOR3_X1 U12582 ( .A1(n11730), .A2(n11729), .A3(n9984), .ZN(n9767) );
  AND2_X1 U12583 ( .A1(n15146), .A2(n15293), .ZN(n9768) );
  AND2_X1 U12584 ( .A1(n15124), .A2(n15288), .ZN(n9769) );
  AND3_X1 U12585 ( .A1(n11863), .A2(n11864), .A3(n11865), .ZN(n9770) );
  OR2_X1 U12586 ( .A1(n10109), .A2(n16131), .ZN(n9771) );
  OR2_X1 U12587 ( .A1(n13255), .A2(n12041), .ZN(n9772) );
  OR2_X1 U12588 ( .A1(n15449), .A2(n16420), .ZN(n9773) );
  INV_X1 U12589 ( .A(n10298), .ZN(n10670) );
  NOR3_X1 U12590 ( .A1(n15596), .A2(n9950), .A3(n15597), .ZN(n15570) );
  OR2_X1 U12591 ( .A1(n9811), .A2(n9810), .ZN(n15511) );
  NAND2_X1 U12592 ( .A1(n11055), .A2(n9754), .ZN(n18028) );
  AND2_X1 U12593 ( .A1(n17963), .A2(n9829), .ZN(n13359) );
  NAND2_X1 U12594 ( .A1(n12875), .A2(n12874), .ZN(n14623) );
  OR3_X1 U12595 ( .A1(n14472), .A2(n9954), .A3(n14473), .ZN(n9774) );
  NOR2_X1 U12596 ( .A1(n15673), .A2(n15674), .ZN(n15667) );
  AND2_X1 U12597 ( .A1(n10858), .A2(n19248), .ZN(n9775) );
  AND2_X1 U12598 ( .A1(n10032), .A2(n14336), .ZN(n9776) );
  AND2_X1 U12599 ( .A1(n14626), .A2(n11616), .ZN(n14636) );
  NOR2_X1 U12600 ( .A1(n14583), .A2(n10036), .ZN(n14986) );
  OR2_X1 U12601 ( .A1(n14158), .A2(n9897), .ZN(n9777) );
  NAND2_X1 U12602 ( .A1(n17963), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13361) );
  NOR2_X1 U12603 ( .A1(n15688), .A2(n15687), .ZN(n9778) );
  AND2_X1 U12604 ( .A1(n10029), .A2(n10028), .ZN(n9779) );
  NAND2_X1 U12605 ( .A1(n13826), .A2(n12032), .ZN(n13901) );
  NOR2_X1 U12606 ( .A1(n13980), .A2(n13981), .ZN(n13979) );
  NAND2_X1 U12607 ( .A1(n10076), .A2(n10078), .ZN(n16368) );
  NAND2_X1 U12608 ( .A1(n9708), .A2(n13304), .ZN(n14617) );
  NAND2_X1 U12609 ( .A1(n16379), .A2(n13277), .ZN(n16374) );
  INV_X1 U12610 ( .A(n10798), .ZN(n10000) );
  OR2_X1 U12611 ( .A1(n19237), .A2(n19245), .ZN(n9780) );
  INV_X1 U12612 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10066) );
  INV_X1 U12613 ( .A(n15759), .ZN(n9915) );
  OR2_X1 U12614 ( .A1(n17206), .A2(n16885), .ZN(n9781) );
  AND2_X1 U12615 ( .A1(n15811), .A2(n13208), .ZN(n9782) );
  NAND2_X1 U12616 ( .A1(n10038), .A2(n12285), .ZN(n15003) );
  NOR2_X1 U12617 ( .A1(n9748), .A2(n15613), .ZN(n13220) );
  INV_X1 U12618 ( .A(n9887), .ZN(n14883) );
  NOR2_X1 U12619 ( .A1(n14891), .A2(n14884), .ZN(n9887) );
  INV_X1 U12620 ( .A(n9885), .ZN(n9884) );
  OR2_X1 U12621 ( .A1(n15007), .A2(n15043), .ZN(n9885) );
  INV_X1 U12622 ( .A(n14953), .ZN(n14969) );
  AND2_X1 U12623 ( .A1(n12186), .A2(n12204), .ZN(n9783) );
  AND2_X1 U12624 ( .A1(n13220), .A2(n13221), .ZN(n13219) );
  NOR2_X1 U12625 ( .A1(n16937), .A2(n16938), .ZN(n9784) );
  AND2_X1 U12626 ( .A1(n10053), .A2(n10052), .ZN(n9785) );
  AOI21_X1 U12627 ( .B1(n16494), .B2(n19504), .A(n10757), .ZN(n10758) );
  INV_X1 U12628 ( .A(n15043), .ZN(n12696) );
  NAND2_X1 U12629 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11219), .ZN(
        n9786) );
  AND2_X1 U12630 ( .A1(n9775), .A2(n10011), .ZN(n9787) );
  OR2_X1 U12631 ( .A1(n15596), .A2(n15597), .ZN(n9788) );
  INV_X1 U12632 ( .A(n13795), .ZN(n20383) );
  AND2_X1 U12633 ( .A1(n13943), .A2(n13989), .ZN(n13988) );
  NOR2_X1 U12634 ( .A1(n13932), .A2(n13942), .ZN(n13943) );
  NAND2_X1 U12635 ( .A1(n9894), .A2(n9895), .ZN(n13969) );
  NOR2_X1 U12636 ( .A1(n13830), .A2(n13831), .ZN(n13832) );
  INV_X1 U12637 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11742) );
  NOR2_X1 U12638 ( .A1(n13722), .A2(n13723), .ZN(n13721) );
  NAND2_X2 U12639 ( .A1(n11715), .A2(n17692), .ZN(n18080) );
  NOR2_X1 U12640 ( .A1(n13830), .A2(n9946), .ZN(n13850) );
  NOR2_X1 U12641 ( .A1(n14455), .A2(n14456), .ZN(n14457) );
  OR2_X1 U12642 ( .A1(n13830), .A2(n9942), .ZN(n13932) );
  AND2_X1 U12643 ( .A1(n14551), .A2(n9877), .ZN(n9789) );
  NOR2_X1 U12644 ( .A1(n13830), .A2(n9944), .ZN(n13906) );
  NOR2_X1 U12645 ( .A1(n18130), .A2(n11047), .ZN(n9790) );
  AND2_X1 U12646 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n9791)
         );
  AND2_X1 U12647 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n9792)
         );
  AND2_X1 U12648 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n9793)
         );
  AND2_X1 U12649 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n9794)
         );
  AND2_X1 U12650 ( .A1(n14551), .A2(n14550), .ZN(n14492) );
  OR2_X1 U12651 ( .A1(n17559), .A2(n17269), .ZN(n9795) );
  NAND2_X1 U12652 ( .A1(n12659), .A2(n12658), .ZN(n14284) );
  INV_X1 U12653 ( .A(n14284), .ZN(n9863) );
  OR2_X1 U12654 ( .A1(n14977), .A2(n14959), .ZN(n9796) );
  NAND2_X1 U12655 ( .A1(n13838), .A2(n9776), .ZN(n10030) );
  NAND2_X1 U12656 ( .A1(n13838), .A2(n10032), .ZN(n10031) );
  AND2_X1 U12657 ( .A1(n14524), .A2(n14489), .ZN(n9797) );
  NOR2_X1 U12658 ( .A1(n13145), .A2(n13144), .ZN(n9798) );
  AND2_X1 U12659 ( .A1(n9895), .A2(n9749), .ZN(n9799) );
  INV_X1 U12660 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n21023) );
  OR3_X1 U12661 ( .A1(n17175), .A2(n16888), .A3(n17176), .ZN(n9800) );
  AND2_X1 U12662 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n9801)
         );
  AND2_X1 U12663 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n9802)
         );
  AND2_X1 U12664 ( .A1(n17845), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11672) );
  AND2_X1 U12665 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n9803) );
  AND2_X1 U12666 ( .A1(n12681), .A2(n12680), .ZN(n14550) );
  INV_X1 U12667 ( .A(n14550), .ZN(n9881) );
  AND2_X1 U12668 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n9804) );
  INV_X1 U12669 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10010) );
  OR2_X1 U12670 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n9805) );
  NOR2_X1 U12671 ( .A1(n18006), .A2(n18045), .ZN(n17979) );
  INV_X1 U12672 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n9812) );
  AND2_X1 U12673 ( .A1(n9747), .A2(n15928), .ZN(n9806) );
  AND2_X1 U12674 ( .A1(n9746), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9807) );
  INV_X1 U12675 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10011) );
  INV_X1 U12676 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9810) );
  INV_X1 U12677 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n9809) );
  AOI22_X2 U12678 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19563), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19562), .ZN(n20051) );
  NOR2_X2 U12679 ( .A1(n19521), .A2(n19520), .ZN(n19562) );
  OAI22_X2 U12680 ( .A1(n16748), .A2(n14147), .B1(n21140), .B2(n14146), .ZN(
        n20935) );
  INV_X1 U12681 ( .A(n9811), .ZN(n15521) );
  NOR2_X2 U12682 ( .A1(n14181), .A2(n19396), .ZN(n14184) );
  NAND2_X1 U12683 ( .A1(n14182), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14181) );
  NAND2_X1 U12684 ( .A1(n16469), .A2(n19384), .ZN(n16496) );
  NAND2_X1 U12685 ( .A1(n16552), .A2(n14305), .ZN(n16539) );
  NOR2_X2 U12686 ( .A1(n14178), .A2(n16678), .ZN(n14180) );
  NOR2_X2 U12687 ( .A1(n15513), .A2(n16619), .ZN(n15516) );
  INV_X1 U12688 ( .A(n9824), .ZN(n13386) );
  INV_X1 U12689 ( .A(n9823), .ZN(n16968) );
  AND2_X2 U12690 ( .A1(n11672), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13379) );
  NAND3_X1 U12691 ( .A1(n16884), .A2(n9827), .A3(n9781), .ZN(n9826) );
  AND2_X1 U12692 ( .A1(n16897), .A2(n17205), .ZN(n16887) );
  NOR2_X1 U12693 ( .A1(n13391), .A2(n17846), .ZN(n16877) );
  AOI21_X2 U12694 ( .B1(n17005), .B2(n16983), .A(n17175), .ZN(n16984) );
  INV_X1 U12695 ( .A(n16984), .ZN(n16995) );
  NAND2_X1 U12696 ( .A1(n10309), .A2(n10295), .ZN(n9831) );
  AND3_X4 U12697 ( .A1(n14807), .A2(n9832), .A3(n10118), .ZN(n10188) );
  NAND2_X2 U12698 ( .A1(n13318), .A2(n15186), .ZN(n15131) );
  INV_X1 U12699 ( .A(n9849), .ZN(n9846) );
  NAND2_X1 U12700 ( .A1(n9849), .A2(n9848), .ZN(n9847) );
  NAND2_X1 U12701 ( .A1(n14707), .A2(n14706), .ZN(n9850) );
  NAND4_X1 U12702 ( .A1(n9770), .A2(n11867), .A3(n11862), .A4(n11870), .ZN(
        n9853) );
  NAND4_X1 U12703 ( .A1(n9851), .A2(n11868), .A3(n11856), .A4(n11857), .ZN(
        n9854) );
  AND2_X2 U12704 ( .A1(n11891), .A2(n13675), .ZN(n12739) );
  NAND2_X1 U12705 ( .A1(n13306), .A2(n15447), .ZN(n15264) );
  XNOR2_X2 U12706 ( .A(n12036), .B(n14098), .ZN(n13856) );
  NAND3_X1 U12707 ( .A1(n9871), .A2(n13828), .A3(n9872), .ZN(n14065) );
  INV_X1 U12708 ( .A(n9886), .ZN(n14993) );
  AND3_X2 U12709 ( .A1(n9894), .A2(n9895), .A3(n9893), .ZN(n14452) );
  AND2_X1 U12710 ( .A1(n15538), .A2(n15619), .ZN(n15848) );
  NAND2_X2 U12711 ( .A1(n10166), .A2(n10167), .ZN(n11390) );
  NAND2_X2 U12712 ( .A1(n10179), .A2(n10178), .ZN(n10248) );
  NAND2_X1 U12713 ( .A1(n10203), .A2(n10248), .ZN(n10249) );
  AOI21_X1 U12714 ( .B1(n9909), .B2(n10660), .A(n10659), .ZN(n13755) );
  OAI21_X1 U12715 ( .B1(n9977), .B2(n14818), .A(n14288), .ZN(n10795) );
  NAND2_X1 U12716 ( .A1(n9910), .A2(n9911), .ZN(n14368) );
  NAND2_X1 U12717 ( .A1(n9977), .A2(n14288), .ZN(n9910) );
  NAND2_X1 U12718 ( .A1(n10894), .A2(n9916), .ZN(n9912) );
  NAND2_X1 U12719 ( .A1(n9912), .A2(n9913), .ZN(n15734) );
  NAND3_X1 U12720 ( .A1(n9915), .A2(n9918), .A3(n9920), .ZN(n9914) );
  NAND2_X1 U12721 ( .A1(n15707), .A2(n9921), .ZN(n9922) );
  NOR2_X2 U12722 ( .A1(n14812), .A2(n9925), .ZN(n9924) );
  AOI21_X2 U12723 ( .B1(n10913), .B2(n9928), .A(n9929), .ZN(n9927) );
  NOR2_X1 U12724 ( .A1(n14472), .A2(n14473), .ZN(n14646) );
  INV_X1 U12725 ( .A(n14645), .ZN(n9954) );
  NAND2_X1 U12726 ( .A1(n15564), .A2(n15509), .ZN(n15508) );
  NAND2_X1 U12727 ( .A1(n13943), .A2(n9957), .ZN(n14333) );
  INV_X1 U12728 ( .A(n14333), .ZN(n10708) );
  INV_X2 U12729 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10935) );
  NAND3_X1 U12730 ( .A1(n11163), .A2(n9965), .A3(n9964), .ZN(n9963) );
  NAND2_X1 U12731 ( .A1(n10457), .A2(n10456), .ZN(n10580) );
  NAND2_X1 U12732 ( .A1(n9973), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9972) );
  NAND4_X1 U12733 ( .A1(n10183), .A2(n10182), .A3(n10181), .A4(n10180), .ZN(
        n9973) );
  NAND2_X1 U12734 ( .A1(n9975), .A2(n10359), .ZN(n9974) );
  NAND4_X1 U12735 ( .A1(n10187), .A2(n10186), .A3(n10184), .A4(n10185), .ZN(
        n9975) );
  NAND2_X1 U12736 ( .A1(n9703), .A2(n13230), .ZN(n15750) );
  AND2_X1 U12737 ( .A1(n13229), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15766) );
  NAND2_X1 U12738 ( .A1(n10581), .A2(n10591), .ZN(n9977) );
  NAND3_X1 U12739 ( .A1(n10581), .A2(n10591), .A3(n14377), .ZN(n14378) );
  AND2_X1 U12740 ( .A1(n9977), .A2(n9976), .ZN(n16670) );
  INV_X1 U12741 ( .A(n14377), .ZN(n9976) );
  NAND3_X1 U12742 ( .A1(n10925), .A2(n9978), .A3(n10758), .ZN(P2_U2985) );
  XNOR2_X1 U12743 ( .A(n15718), .B(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15837) );
  NAND2_X1 U12744 ( .A1(n9980), .A2(n10808), .ZN(n9979) );
  NAND2_X1 U12745 ( .A1(n14449), .A2(n14445), .ZN(n10605) );
  NAND2_X1 U12746 ( .A1(n9758), .A2(n18155), .ZN(n9981) );
  XNOR2_X1 U12747 ( .A(n11039), .B(n11027), .ZN(n18155) );
  NAND2_X1 U12748 ( .A1(n9758), .A2(n18156), .ZN(n9982) );
  INV_X1 U12749 ( .A(n9983), .ZN(n18166) );
  NAND2_X1 U12750 ( .A1(n9985), .A2(n9767), .ZN(P3_U2834) );
  NAND2_X1 U12751 ( .A1(n9986), .A2(n11731), .ZN(n9985) );
  NAND2_X1 U12752 ( .A1(n9987), .A2(n11724), .ZN(n9986) );
  NAND2_X1 U12753 ( .A1(n11721), .A2(n11720), .ZN(n9987) );
  NAND3_X1 U12754 ( .A1(n9988), .A2(n18131), .A3(n9990), .ZN(n9989) );
  INV_X1 U12755 ( .A(n11047), .ZN(n9988) );
  OAI211_X1 U12756 ( .C1(n9736), .C2(n11047), .A(n9989), .B(n9743), .ZN(n18111) );
  NOR2_X1 U12757 ( .A1(n18131), .A2(n18450), .ZN(n18130) );
  INV_X1 U12758 ( .A(n18123), .ZN(n9992) );
  AND2_X2 U12759 ( .A1(n11725), .A2(n18196), .ZN(n17836) );
  NAND4_X2 U12760 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(n9998), .A4(n9997), .ZN(
        n10949) );
  INV_X2 U12761 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9997) );
  NAND2_X1 U12762 ( .A1(n10782), .A2(n9999), .ZN(n10778) );
  NAND2_X1 U12763 ( .A1(n10801), .A2(n10002), .ZN(n10001) );
  NAND2_X1 U12764 ( .A1(n10813), .A2(n10005), .ZN(n10824) );
  AND2_X1 U12765 ( .A1(n10863), .A2(n10858), .ZN(n10866) );
  NAND2_X1 U12766 ( .A1(n10863), .A2(n9787), .ZN(n10890) );
  AND2_X2 U12767 ( .A1(n19367), .A2(n10012), .ZN(n10852) );
  NAND2_X2 U12768 ( .A1(n10830), .A2(n10906), .ZN(n19367) );
  INV_X2 U12769 ( .A(n13106), .ZN(n13090) );
  AOI21_X1 U12770 ( .B1(n15552), .B2(n9745), .A(n9798), .ZN(n10019) );
  INV_X1 U12771 ( .A(n15607), .ZN(n12928) );
  NAND2_X1 U12772 ( .A1(n12875), .A2(n10021), .ZN(n15607) );
  NAND2_X1 U12773 ( .A1(n13004), .A2(n10025), .ZN(n10026) );
  INV_X1 U12774 ( .A(n10029), .ZN(n15592) );
  XNOR2_X1 U12775 ( .A(n13052), .B(n13050), .ZN(n15575) );
  NAND2_X1 U12776 ( .A1(n13838), .A2(n9742), .ZN(n14420) );
  NAND2_X1 U12777 ( .A1(n13838), .A2(n12823), .ZN(n14074) );
  NAND2_X1 U12778 ( .A1(n10033), .A2(n9772), .ZN(n12005) );
  NAND3_X1 U12779 ( .A1(n12036), .A2(n21023), .A3(n11991), .ZN(n10033) );
  OAI21_X1 U12780 ( .B1(n13246), .B2(n12009), .A(n10034), .ZN(n13824) );
  AND3_X2 U12781 ( .A1(n12187), .A2(n12188), .A3(n10041), .ZN(n14572) );
  NAND3_X1 U12782 ( .A1(n12187), .A2(n12188), .A3(n10044), .ZN(n14488) );
  AND2_X1 U12783 ( .A1(n14881), .A2(n10049), .ZN(n13330) );
  NAND2_X1 U12784 ( .A1(n14881), .A2(n10047), .ZN(n12765) );
  NAND2_X1 U12785 ( .A1(n14881), .A2(n14882), .ZN(n14869) );
  XNOR2_X1 U12787 ( .A(n10055), .B(n10083), .ZN(n14675) );
  OAI21_X2 U12788 ( .B1(n15776), .B2(n13213), .A(n15777), .ZN(n10055) );
  AND2_X2 U12789 ( .A1(n15799), .A2(n10056), .ZN(n15776) );
  NAND2_X1 U12790 ( .A1(n15799), .A2(n15801), .ZN(n15789) );
  OAI21_X1 U12791 ( .B1(n10822), .B2(n10059), .A(n10828), .ZN(n10058) );
  NAND2_X1 U12792 ( .A1(n13206), .A2(n10062), .ZN(n10064) );
  CLKBUF_X1 U12793 ( .A(n10064), .Z(n10061) );
  INV_X1 U12794 ( .A(n10061), .ZN(n15818) );
  NAND2_X1 U12795 ( .A1(n10459), .A2(n10458), .ZN(n10591) );
  INV_X1 U12796 ( .A(n10600), .ZN(n10777) );
  AND3_X2 U12797 ( .A1(n10458), .A2(n10459), .A3(n11420), .ZN(n10599) );
  AND2_X2 U12798 ( .A1(n11752), .A2(n13559), .ZN(n11803) );
  NAND2_X1 U12799 ( .A1(n13237), .A2(n9669), .ZN(n10067) );
  NAND2_X1 U12800 ( .A1(n16381), .A2(n16380), .ZN(n16379) );
  NAND2_X1 U12801 ( .A1(n16381), .A2(n10077), .ZN(n10076) );
  NOR2_X2 U12803 ( .A1(n17964), .A2(n18066), .ZN(n17935) );
  NOR2_X1 U12804 ( .A1(n10438), .A2(n10437), .ZN(n10453) );
  AND2_X1 U12805 ( .A1(n12788), .A2(n10342), .ZN(n10343) );
  OAI211_X1 U12806 ( .C1(n9750), .C2(n12882), .A(n10418), .B(n10417), .ZN(
        n10419) );
  NOR2_X1 U12807 ( .A1(n9750), .A2(n12846), .ZN(n10335) );
  NAND2_X1 U12808 ( .A1(n10204), .A2(n10235), .ZN(n10205) );
  AOI22_X1 U12809 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11117) );
  NOR2_X1 U12810 ( .A1(n10451), .A2(n10450), .ZN(n10452) );
  AND2_X1 U12811 ( .A1(n10226), .A2(n10225), .ZN(n13173) );
  INV_X2 U12812 ( .A(n11910), .ZN(n11879) );
  AND2_X2 U12813 ( .A1(n11810), .A2(n11809), .ZN(n11910) );
  NAND2_X1 U12814 ( .A1(n11880), .A2(n12770), .ZN(n11881) );
  AOI22_X1 U12815 ( .A1(n9721), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10194), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10174) );
  AOI22_X1 U12816 ( .A1(n9721), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9668), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10136) );
  OR2_X2 U12817 ( .A1(n10329), .A2(n10328), .ZN(n19721) );
  NOR2_X1 U12818 ( .A1(n15146), .A2(n10108), .ZN(n14707) );
  NAND2_X1 U12819 ( .A1(n15147), .A2(n15153), .ZN(n15146) );
  INV_X1 U12820 ( .A(n10967), .ZN(n10969) );
  NAND2_X1 U12821 ( .A1(n15054), .A2(n15053), .ZN(n15056) );
  AND2_X1 U12822 ( .A1(n15160), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15171) );
  CLKBUF_X1 U12823 ( .A(n10599), .Z(n10590) );
  NAND2_X1 U12824 ( .A1(n10259), .A2(n10258), .ZN(n10279) );
  AOI22_X1 U12825 ( .A1(n10358), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14000), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10119) );
  NAND2_X1 U12826 ( .A1(n10092), .A2(n10357), .ZN(n10415) );
  AOI211_X1 U12827 ( .C1(n17421), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n11025), .B(n11024), .ZN(n11716) );
  INV_X1 U12828 ( .A(n11716), .ZN(n17692) );
  INV_X1 U12829 ( .A(n15116), .ZN(n15080) );
  OR2_X2 U12830 ( .A1(n14090), .A2(n14089), .ZN(n15116) );
  NAND2_X1 U12831 ( .A1(n10646), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10272) );
  AND2_X1 U12833 ( .A1(n14808), .A2(n14810), .ZN(n10082) );
  AND2_X1 U12834 ( .A1(n13215), .A2(n13214), .ZN(n10083) );
  NAND2_X1 U12835 ( .A1(n10852), .A2(n10846), .ZN(n10839) );
  NOR3_X1 U12836 ( .A1(n13229), .A2(n14671), .A3(n16717), .ZN(n10084) );
  OR2_X1 U12837 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17175), .ZN(
        n10085) );
  AND2_X1 U12838 ( .A1(n18080), .A2(n11726), .ZN(n10086) );
  INV_X1 U12839 ( .A(n18545), .ZN(n18741) );
  AND2_X1 U12840 ( .A1(n11708), .A2(n18150), .ZN(n10089) );
  NOR2_X1 U12841 ( .A1(n13988), .A2(n13990), .ZN(n10090) );
  AND2_X1 U12842 ( .A1(n10349), .A2(n10348), .ZN(n10092) );
  OR2_X1 U12843 ( .A1(n10760), .A2(n19551), .ZN(n10093) );
  AND2_X1 U12844 ( .A1(n11321), .A2(n13338), .ZN(n10094) );
  AND2_X1 U12845 ( .A1(n10131), .A2(n10359), .ZN(n10097) );
  AND2_X1 U12846 ( .A1(n11276), .A2(n11275), .ZN(n10098) );
  NAND2_X1 U12847 ( .A1(n10372), .A2(n10359), .ZN(n10099) );
  OR2_X1 U12848 ( .A1(n18066), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10100) );
  AND3_X1 U12849 ( .A1(n18362), .A2(n18328), .A3(n11056), .ZN(n10101) );
  INV_X1 U12850 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14709) );
  AND2_X1 U12851 ( .A1(n18066), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10102) );
  NAND2_X1 U12852 ( .A1(n10249), .A2(n9684), .ZN(n10267) );
  INV_X1 U12853 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11027) );
  NOR2_X1 U12854 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18066), .ZN(
        n10103) );
  AND2_X1 U12855 ( .A1(n10980), .A2(n10979), .ZN(n10104) );
  AND3_X1 U12856 ( .A1(n10136), .A2(n10135), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10105) );
  OAI211_X1 U12857 ( .C1(n9672), .C2(n17437), .A(n11127), .B(n11126), .ZN(
        n16091) );
  INV_X1 U12858 ( .A(n16091), .ZN(n18533) );
  AND2_X1 U12859 ( .A1(n9732), .A2(n17691), .ZN(n17555) );
  NAND2_X1 U12860 ( .A1(n15689), .A2(n13176), .ZN(n19465) );
  INV_X1 U12861 ( .A(n19465), .ZN(n13177) );
  INV_X1 U12862 ( .A(n13027), .ZN(n13002) );
  INV_X1 U12863 ( .A(n14327), .ZN(n10342) );
  INV_X1 U12864 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n16225) );
  NOR2_X1 U12865 ( .A1(n11877), .A2(n12006), .ZN(n12104) );
  INV_X1 U12866 ( .A(n12127), .ZN(n12567) );
  INV_X2 U12867 ( .A(n9659), .ZN(n10747) );
  INV_X1 U12868 ( .A(n10977), .ZN(n10970) );
  OR3_X1 U12869 ( .A1(n15857), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14830), .ZN(n10106) );
  OR3_X1 U12870 ( .A1(n15857), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n11658), .ZN(n10107) );
  OR2_X1 U12871 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10108) );
  INV_X1 U12872 ( .A(n15004), .ZN(n15032) );
  OR2_X1 U12873 ( .A1(n19212), .A2(n9730), .ZN(n16671) );
  OR2_X2 U12874 ( .A1(n10932), .A2(n10934), .ZN(n10109) );
  INV_X1 U12875 ( .A(n19538), .ZN(n11288) );
  INV_X1 U12876 ( .A(n17890), .ZN(n17929) );
  NOR2_X1 U12877 ( .A1(n17977), .A2(n18118), .ZN(n17890) );
  AND2_X1 U12878 ( .A1(n17835), .A2(n11715), .ZN(n10110) );
  OR2_X1 U12879 ( .A1(n12821), .A2(n13927), .ZN(n10111) );
  INV_X1 U12880 ( .A(n20813), .ZN(n20886) );
  NOR2_X1 U12881 ( .A1(n20769), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10112) );
  INV_X1 U12882 ( .A(n10310), .ZN(n10296) );
  AND2_X1 U12883 ( .A1(n9734), .A2(n10345), .ZN(n10113) );
  AND4_X1 U12884 ( .A1(n11790), .A2(n11789), .A3(n11788), .A4(n11787), .ZN(
        n10115) );
  AND2_X1 U12885 ( .A1(n13675), .A2(n12589), .ZN(n13291) );
  AND2_X1 U12886 ( .A1(n14162), .A2(n13545), .ZN(n11898) );
  NAND2_X1 U12887 ( .A1(n11879), .A2(n12589), .ZN(n11880) );
  OR2_X1 U12888 ( .A1(n10670), .A2(n11419), .ZN(n10300) );
  AND2_X1 U12889 ( .A1(n19538), .A2(n13338), .ZN(n10234) );
  INV_X1 U12890 ( .A(n12042), .ZN(n12003) );
  INV_X1 U12891 ( .A(n10272), .ZN(n10254) );
  MUX2_X1 U12892 ( .A(n11315), .B(n10248), .S(n10236), .Z(n10238) );
  OR2_X1 U12893 ( .A1(n12101), .A2(n12100), .ZN(n13279) );
  OR2_X1 U12894 ( .A1(n12076), .A2(n12075), .ZN(n13269) );
  OR2_X1 U12895 ( .A1(n12122), .A2(n12121), .ZN(n13287) );
  AND4_X1 U12896 ( .A1(n10552), .A2(n10551), .A3(n10550), .A4(n10549), .ZN(
        n10553) );
  OAI21_X1 U12897 ( .B1(n10416), .B2(n10415), .A(n10414), .ZN(n10579) );
  INV_X1 U12898 ( .A(n10267), .ZN(n11356) );
  INV_X1 U12899 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11056) );
  INV_X1 U12900 ( .A(n12594), .ZN(n12587) );
  INV_X1 U12901 ( .A(n14954), .ZN(n12373) );
  INV_X1 U12902 ( .A(n14068), .ZN(n12088) );
  INV_X1 U12903 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12057) );
  INV_X1 U12904 ( .A(n12129), .ZN(n12130) );
  OR2_X1 U12905 ( .A1(n13027), .A2(n13026), .ZN(n13028) );
  INV_X1 U12906 ( .A(n13156), .ZN(n13147) );
  INV_X1 U12907 ( .A(n14471), .ZN(n12856) );
  AOI22_X1 U12908 ( .A1(n9665), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14000), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10125) );
  NAND2_X1 U12909 ( .A1(n15712), .A2(n15710), .ZN(n15708) );
  INV_X1 U12910 ( .A(n10602), .ZN(n10557) );
  AND3_X1 U12911 ( .A1(n19538), .A2(n11315), .A3(n11350), .ZN(n10242) );
  NAND2_X1 U12912 ( .A1(n10253), .A2(n10252), .ZN(n10268) );
  AND2_X1 U12913 ( .A1(n11059), .A2(n18278), .ZN(n11054) );
  NOR2_X1 U12914 ( .A1(n11191), .A2(n11180), .ZN(n11167) );
  AOI21_X1 U12915 ( .B1(n12583), .B2(n12582), .A(n12577), .ZN(n12581) );
  INV_X1 U12916 ( .A(n14944), .ZN(n12395) );
  INV_X1 U12917 ( .A(n15031), .ZN(n12320) );
  INV_X1 U12918 ( .A(n13825), .ZN(n12030) );
  NAND2_X1 U12919 ( .A1(n12509), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11843) );
  NAND2_X1 U12920 ( .A1(n12423), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12424) );
  INV_X1 U12921 ( .A(n15041), .ZN(n12285) );
  INV_X1 U12922 ( .A(n12170), .ZN(n12139) );
  INV_X1 U12923 ( .A(n12104), .ZN(n12127) );
  OR2_X1 U12924 ( .A1(n13710), .A2(n13244), .ZN(n13245) );
  OR2_X1 U12925 ( .A1(n9674), .A2(n13313), .ZN(n15231) );
  AND2_X1 U12926 ( .A1(n12679), .A2(n12678), .ZN(n14557) );
  AOI21_X1 U12927 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20175), .A(
        n10623), .ZN(n10630) );
  AND2_X1 U12928 ( .A1(n14075), .A2(n13985), .ZN(n12823) );
  INV_X2 U12929 ( .A(n10670), .ZN(n11340) );
  INV_X1 U12930 ( .A(n15578), .ZN(n13049) );
  AND3_X1 U12931 ( .A1(n11622), .A2(n11621), .A3(n11620), .ZN(n15674) );
  INV_X1 U12932 ( .A(n11656), .ZN(n10617) );
  AND3_X1 U12933 ( .A1(n11612), .A2(n11611), .A3(n11610), .ZN(n14627) );
  AND2_X1 U12934 ( .A1(n15968), .A2(n14765), .ZN(n11377) );
  NAND2_X1 U12935 ( .A1(n10257), .A2(n13406), .ZN(n11344) );
  NAND2_X1 U12936 ( .A1(n12789), .A2(n20195), .ZN(n12813) );
  INV_X1 U12937 ( .A(n10340), .ZN(n10330) );
  AND2_X1 U12938 ( .A1(n11362), .A2(n11361), .ZN(n13996) );
  INV_X1 U12939 ( .A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17493) );
  OAI21_X1 U12940 ( .B1(n11718), .B2(n17692), .A(n11732), .ZN(n11719) );
  NOR2_X1 U12941 ( .A1(n17990), .A2(n11665), .ZN(n11061) );
  NOR2_X1 U12942 ( .A1(n11210), .A2(n17712), .ZN(n11040) );
  NOR2_X1 U12943 ( .A1(n17727), .A2(n18548), .ZN(n11238) );
  AOI211_X1 U12944 ( .C1(n17512), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n11125), .B(n11124), .ZN(n11126) );
  NAND2_X1 U12945 ( .A1(n13551), .A2(n11889), .ZN(n12630) );
  NAND2_X1 U12946 ( .A1(n11894), .A2(n13686), .ZN(n14091) );
  NAND2_X1 U12947 ( .A1(n12375), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12376) );
  INV_X1 U12948 ( .A(n12563), .ZN(n12534) );
  NAND2_X1 U12949 ( .A1(n12139), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12154) );
  NAND2_X1 U12950 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12059) );
  OAI211_X1 U12951 ( .C1(n12613), .C2(n20481), .A(n11943), .B(n11942), .ZN(
        n12021) );
  OR2_X1 U12952 ( .A1(n15034), .A2(n14991), .ZN(n12706) );
  AND2_X1 U12953 ( .A1(n12702), .A2(n12701), .ZN(n15034) );
  NAND2_X1 U12954 ( .A1(n12040), .A2(n12039), .ZN(n14098) );
  OR2_X1 U12955 ( .A1(n15489), .A2(n20880), .ZN(n14097) );
  OAI22_X1 U12956 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n13532), .B1(
        n10624), .B2(n10630), .ZN(n11309) );
  AND2_X1 U12957 ( .A1(n12996), .A2(n12995), .ZN(n13003) );
  INV_X1 U12958 ( .A(n14634), .ZN(n11616) );
  OR2_X1 U12959 ( .A1(n15992), .A2(n11376), .ZN(n15952) );
  AND3_X1 U12960 ( .A1(n11607), .A2(n11606), .A3(n11605), .ZN(n14434) );
  NAND2_X1 U12961 ( .A1(n10315), .A2(n10316), .ZN(n10314) );
  NAND2_X1 U12962 ( .A1(n14346), .A2(n12809), .ZN(n12800) );
  OR2_X2 U12963 ( .A1(n10351), .A2(n10330), .ZN(n19576) );
  OAI22_X1 U12964 ( .A1(n9997), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n19010), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11191) );
  INV_X1 U12965 ( .A(n11156), .ZN(n11128) );
  NAND2_X1 U12966 ( .A1(n17834), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11670) );
  NAND3_X1 U12967 ( .A1(n17876), .A2(n17882), .A3(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17864) );
  INV_X1 U12968 ( .A(n18056), .ZN(n18068) );
  NOR2_X1 U12969 ( .A1(n11223), .A2(n18106), .ZN(n11226) );
  AOI21_X1 U12970 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n19019), .A(
        n11176), .ZN(n11194) );
  INV_X1 U12971 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16321) );
  INV_X1 U12972 ( .A(n20347), .ZN(n14972) );
  NOR2_X1 U12973 ( .A1(n14163), .A2(n11941), .ZN(n12757) );
  NOR2_X1 U12974 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12537) );
  OR2_X1 U12975 ( .A1(n12376), .A2(n14945), .ZN(n12422) );
  NAND2_X1 U12976 ( .A1(n12315), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12351) );
  AND2_X1 U12977 ( .A1(n12184), .A2(n12183), .ZN(n14405) );
  OAI21_X1 U12978 ( .B1(n15131), .B2(n15133), .A(n10075), .ZN(n15153) );
  AND2_X1 U12979 ( .A1(n12695), .A2(n12694), .ZN(n15043) );
  AND2_X1 U12980 ( .A1(n13704), .A2(n20475), .ZN(n16404) );
  INV_X1 U12981 ( .A(n20466), .ZN(n13704) );
  OR2_X1 U12982 ( .A1(n20580), .A2(n20839), .ZN(n20588) );
  OR2_X1 U12983 ( .A1(n20580), .A2(n20579), .ZN(n20620) );
  OR2_X1 U12984 ( .A1(n20649), .A2(n20839), .ZN(n20670) );
  OR2_X1 U12985 ( .A1(n20885), .A2(n20616), .ZN(n14543) );
  OR3_X1 U12986 ( .A1(n20774), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n14105), 
        .ZN(n14149) );
  INV_X1 U12987 ( .A(n19432), .ZN(n19400) );
  OR2_X1 U12988 ( .A1(n11309), .A2(n10633), .ZN(n14021) );
  INV_X1 U12989 ( .A(n14305), .ZN(n19419) );
  OR2_X1 U12990 ( .A1(n13636), .A2(n13635), .ZN(n13637) );
  INV_X1 U12991 ( .A(n15575), .ZN(n15579) );
  AND4_X1 U12992 ( .A1(n11501), .A2(n11500), .A3(n11499), .A4(n11498), .ZN(
        n13888) );
  XNOR2_X1 U12993 ( .A(n11415), .B(n11414), .ZN(n13915) );
  INV_X1 U12994 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15813) );
  INV_X1 U12995 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19396) );
  OR2_X1 U12996 ( .A1(n15564), .A2(n15563), .ZN(n16509) );
  OR2_X1 U12997 ( .A1(n10883), .A2(n15932), .ZN(n15777) );
  OR2_X1 U12998 ( .A1(n15995), .A2(n11656), .ZN(n15944) );
  INV_X1 U12999 ( .A(n16710), .ZN(n16072) );
  INV_X1 U13000 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14308) );
  AND2_X1 U13001 ( .A1(n20178), .A2(n20190), .ZN(n20164) );
  INV_X1 U13002 ( .A(n10221), .ZN(n19522) );
  NOR2_X1 U13003 ( .A1(n19186), .A2(n17727), .ZN(n11252) );
  INV_X1 U13004 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17097) );
  INV_X1 U13005 ( .A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17471) );
  INV_X1 U13006 ( .A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17418) );
  NAND2_X1 U13007 ( .A1(n11671), .A2(n11670), .ZN(n11679) );
  AOI21_X1 U13008 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17890), .A(
        n18545), .ZN(n17941) );
  INV_X1 U13009 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n18008) );
  NOR2_X1 U13010 ( .A1(n11225), .A2(n11229), .ZN(n11231) );
  NAND2_X1 U13011 ( .A1(n18242), .A2(n11734), .ZN(n16199) );
  NAND2_X1 U13012 ( .A1(n17848), .A2(n18186), .ZN(n17847) );
  NOR2_X1 U13013 ( .A1(n18279), .A2(n18206), .ZN(n18231) );
  NAND2_X1 U13014 ( .A1(n19195), .A2(n16093), .ZN(n18469) );
  INV_X1 U13015 ( .A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16131) );
  INV_X1 U13016 ( .A(n14656), .ZN(n17726) );
  INV_X1 U13017 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19010) );
  INV_X1 U13018 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18976) );
  INV_X1 U13019 ( .A(n14086), .ZN(n13688) );
  AND2_X1 U13020 ( .A1(n16248), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14860) );
  OAI21_X1 U13021 ( .B1(n15016), .B2(n20351), .A(n12761), .ZN(n12762) );
  NOR2_X1 U13022 ( .A1(n14972), .A2(n14971), .ZN(n16342) );
  OR2_X1 U13023 ( .A1(n21025), .A2(n12635), .ZN(n20334) );
  INV_X1 U13024 ( .A(n20289), .ZN(n20310) );
  AND2_X1 U13025 ( .A1(n12757), .A2(n12755), .ZN(n20347) );
  INV_X1 U13026 ( .A(n14587), .ZN(n15044) );
  INV_X1 U13027 ( .A(n15048), .ZN(n15038) );
  AND2_X1 U13028 ( .A1(n15116), .A2(n15052), .ZN(n15053) );
  INV_X1 U13029 ( .A(n15084), .ZN(n15120) );
  OR2_X1 U13030 ( .A1(n14427), .A2(n14426), .ZN(n14555) );
  AND2_X1 U13031 ( .A1(n15116), .A2(n14092), .ZN(n15115) );
  INV_X2 U13032 ( .A(n13761), .ZN(n20413) );
  NOR2_X2 U13033 ( .A1(n20383), .A2(n14133), .ZN(n20398) );
  NAND2_X1 U13034 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n12282), .ZN(
        n12313) );
  NAND2_X1 U13035 ( .A1(n12190), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12218) );
  AND2_X1 U13036 ( .A1(n12123), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12134) );
  OR2_X1 U13037 ( .A1(n20422), .A2(n13325), .ZN(n15254) );
  INV_X1 U13038 ( .A(n20427), .ZN(n16355) );
  NOR2_X1 U13039 ( .A1(n15474), .A2(n15477), .ZN(n16428) );
  INV_X1 U13040 ( .A(n16404), .ZN(n20450) );
  INV_X1 U13041 ( .A(n20469), .ZN(n20440) );
  OR2_X1 U13042 ( .A1(n15489), .A2(n14232), .ZN(n20616) );
  INV_X1 U13043 ( .A(n20560), .ZN(n20553) );
  OAI21_X1 U13044 ( .B1(n20537), .B2(n20536), .A(n20535), .ZN(n20562) );
  INV_X1 U13045 ( .A(n20588), .ZN(n20611) );
  INV_X1 U13046 ( .A(n20620), .ZN(n20640) );
  INV_X1 U13047 ( .A(n20670), .ZN(n20699) );
  NOR2_X2 U13048 ( .A1(n20649), .A2(n20739), .ZN(n20698) );
  INV_X1 U13049 ( .A(n20811), .ZN(n20880) );
  NOR2_X2 U13050 ( .A1(n20649), .A2(n20579), .ZN(n20729) );
  INV_X1 U13051 ( .A(n20616), .ZN(n20704) );
  NOR2_X2 U13052 ( .A1(n20812), .A2(n20839), .ZN(n20834) );
  INV_X1 U13053 ( .A(n20812), .ZN(n20705) );
  INV_X1 U13054 ( .A(n20940), .ZN(n20926) );
  AND2_X1 U13055 ( .A1(n12747), .A2(n20954), .ZN(n16265) );
  INV_X1 U13056 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20954) );
  INV_X1 U13057 ( .A(n20987), .ZN(n20999) );
  NAND2_X1 U13058 ( .A1(n16553), .A2(n16554), .ZN(n16552) );
  INV_X1 U13059 ( .A(n19413), .ZN(n19432) );
  INV_X1 U13060 ( .A(n19434), .ZN(n19403) );
  OAI21_X1 U13061 ( .B1(n16481), .B2(n13835), .A(n13340), .ZN(n13341) );
  XNOR2_X1 U13062 ( .A(n13741), .B(n13745), .ZN(n13744) );
  NAND2_X1 U13063 ( .A1(n13175), .A2(n13336), .ZN(n19462) );
  INV_X1 U13064 ( .A(n16677), .ZN(n19501) );
  INV_X1 U13065 ( .A(n16668), .ZN(n19505) );
  INV_X1 U13066 ( .A(n15766), .ZN(n15914) );
  AND2_X1 U13067 ( .A1(n11368), .A2(n15964), .ZN(n15968) );
  INV_X1 U13068 ( .A(n20016), .ZN(n20170) );
  OAI21_X1 U13069 ( .B1(n19529), .B2(n19528), .A(n19527), .ZN(n19568) );
  NOR2_X1 U13070 ( .A1(n19811), .A2(n19719), .ZN(n19596) );
  AND2_X1 U13071 ( .A1(n20178), .A2(n19513), .ZN(n19573) );
  INV_X1 U13072 ( .A(n20164), .ZN(n19871) );
  NOR2_X1 U13073 ( .A1(n19719), .A2(n19940), .ZN(n19711) );
  AND2_X1 U13074 ( .A1(n19758), .A2(n19951), .ZN(n19745) );
  INV_X1 U13075 ( .A(n19803), .ZN(n19805) );
  INV_X1 U13076 ( .A(n19573), .ZN(n19811) );
  NOR2_X1 U13077 ( .A1(n19978), .A2(n19871), .ZN(n19902) );
  OAI21_X1 U13078 ( .B1(n19934), .B2(n20195), .A(n19913), .ZN(n19936) );
  INV_X1 U13079 ( .A(n20057), .ZN(n19965) );
  OAI21_X1 U13080 ( .B1(n19988), .B2(n19987), .A(n19986), .ZN(n20009) );
  INV_X1 U13081 ( .A(n19994), .ZN(n20030) );
  INV_X1 U13082 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19942) );
  INV_X1 U13083 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n20086) );
  NOR2_X1 U13084 ( .A1(n19116), .A2(n16872), .ZN(n16909) );
  INV_X1 U13085 ( .A(n16962), .ZN(n16953) );
  NOR2_X1 U13086 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16971), .ZN(n16964) );
  NOR2_X1 U13087 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16988), .ZN(n16972) );
  NOR2_X1 U13088 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17055), .ZN(n17038) );
  NOR2_X1 U13089 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17103), .ZN(n17087) );
  NOR2_X1 U13090 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17124), .ZN(n17109) );
  NOR2_X2 U13091 ( .A1(n19200), .A2(n19027), .ZN(n17165) );
  INV_X1 U13092 ( .A(n17221), .ZN(n17204) );
  NOR2_X1 U13093 ( .A1(n17774), .A2(n17630), .ZN(n17626) );
  OAI211_X1 U13094 ( .C1(n10946), .C2(n16131), .A(n11117), .B(n11116), .ZN(
        n17727) );
  NOR2_X1 U13095 ( .A1(n11679), .A2(n11678), .ZN(n11680) );
  INV_X1 U13096 ( .A(n18024), .ZN(n18036) );
  INV_X1 U13097 ( .A(n18093), .ZN(n18075) );
  INV_X1 U13098 ( .A(n18370), .ZN(n18004) );
  NOR2_X1 U13099 ( .A1(n11664), .A2(n16094), .ZN(n18168) );
  NOR2_X1 U13100 ( .A1(n18231), .A2(n18494), .ZN(n18255) );
  INV_X1 U13101 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18378) );
  INV_X1 U13102 ( .A(n18418), .ZN(n18399) );
  INV_X1 U13103 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18433) );
  INV_X1 U13104 ( .A(n18469), .ZN(n19000) );
  INV_X1 U13105 ( .A(n18492), .ZN(n18498) );
  NAND2_X1 U13106 ( .A1(n19039), .A2(n18515), .ZN(n18667) );
  CLKBUF_X1 U13107 ( .A(n18635), .Z(n18639) );
  INV_X1 U13108 ( .A(n18714), .ZN(n18701) );
  INV_X1 U13109 ( .A(n18737), .ZN(n18766) );
  INV_X1 U13110 ( .A(n18905), .ZN(n18890) );
  AND2_X1 U13111 ( .A1(n18879), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18908) );
  INV_X1 U13112 ( .A(n18593), .ZN(n18960) );
  INV_X1 U13113 ( .A(n11664), .ZN(n19025) );
  NOR2_X1 U13114 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13358), .ZN(n16836)
         );
  NAND2_X1 U13115 ( .A1(n13688), .A2(n14852), .ZN(n13660) );
  INV_X1 U13116 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21170) );
  INV_X1 U13117 ( .A(n12762), .ZN(n12763) );
  INV_X1 U13118 ( .A(n20287), .ZN(n16324) );
  INV_X1 U13119 ( .A(n20315), .ZN(n20342) );
  AND2_X1 U13120 ( .A1(n15118), .A2(n14700), .ZN(n14586) );
  INV_X1 U13121 ( .A(n20352), .ZN(n20375) );
  NOR2_X1 U13122 ( .A1(n13660), .A2(n13659), .ZN(n13795) );
  NAND2_X1 U13123 ( .A1(n15254), .A2(n13717), .ZN(n20427) );
  INV_X1 U13124 ( .A(n20422), .ZN(n20238) );
  NAND2_X1 U13125 ( .A1(n13703), .A2(n13697), .ZN(n20469) );
  NAND2_X1 U13126 ( .A1(n13703), .A2(n13695), .ZN(n20470) );
  NAND2_X1 U13127 ( .A1(n13703), .A2(n16217), .ZN(n20475) );
  INV_X1 U13128 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20733) );
  AOI211_X2 U13129 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20619), .A(n14394), 
        .B(n14393), .ZN(n20498) );
  OR2_X1 U13130 ( .A1(n20580), .A2(n20616), .ZN(n20511) );
  OR2_X1 U13131 ( .A1(n20580), .A2(n20739), .ZN(n20560) );
  AOI22_X1 U13132 ( .A1(n20531), .A2(n20536), .B1(n20771), .B2(n10112), .ZN(
        n20565) );
  AOI22_X1 U13133 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20574), .B1(n20576), 
        .B2(n20571), .ZN(n20615) );
  NAND2_X1 U13134 ( .A1(n20617), .A2(n20704), .ZN(n20669) );
  AOI22_X1 U13135 ( .A1(n20675), .A2(n20681), .B1(n20674), .B2(n10112), .ZN(
        n20703) );
  NAND2_X1 U13136 ( .A1(n20705), .A2(n20704), .ZN(n20763) );
  AOI22_X1 U13137 ( .A1(n20777), .A2(n20772), .B1(n20771), .B2(n20770), .ZN(
        n20804) );
  NAND2_X1 U13138 ( .A1(n20705), .A2(n14495), .ZN(n20838) );
  INV_X1 U13139 ( .A(n20923), .ZN(n20797) );
  AOI21_X1 U13140 ( .B1(n14231), .B2(n14499), .A(n20813), .ZN(n14273) );
  OR2_X1 U13141 ( .A1(n20885), .A2(n20839), .ZN(n20929) );
  INV_X1 U13142 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20942) );
  INV_X1 U13143 ( .A(n20945), .ZN(n21008) );
  AND2_X1 U13144 ( .A1(n20954), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n21031) );
  NOR2_X1 U13145 ( .A1(n14033), .A2(n19210), .ZN(n19208) );
  OR3_X1 U13146 ( .A1(n14188), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20215), 
        .ZN(n19422) );
  OR3_X1 U13147 ( .A1(n14188), .A2(n16472), .A3(n14176), .ZN(n19434) );
  INV_X1 U13148 ( .A(n13341), .ZN(n13342) );
  INV_X1 U13149 ( .A(n13835), .ZN(n15616) );
  AND2_X1 U13150 ( .A1(n13195), .A2(n13194), .ZN(n13196) );
  NAND2_X1 U13151 ( .A1(n15689), .A2(n13646), .ZN(n14356) );
  NOR2_X1 U13152 ( .A1(n19472), .A2(n19497), .ZN(n19484) );
  INV_X1 U13153 ( .A(n19472), .ZN(n19499) );
  INV_X1 U13154 ( .A(n14195), .ZN(n13534) );
  INV_X1 U13155 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16591) );
  INV_X1 U13156 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16619) );
  INV_X1 U13157 ( .A(n19504), .ZN(n16655) );
  NOR2_X1 U13158 ( .A1(n13231), .A2(n10084), .ZN(n13232) );
  INV_X1 U13159 ( .A(n16700), .ZN(n16717) );
  INV_X1 U13160 ( .A(n16721), .ZN(n16704) );
  INV_X1 U13161 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20182) );
  INV_X1 U13162 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13532) );
  INV_X1 U13163 ( .A(n19596), .ZN(n19572) );
  NAND2_X1 U13164 ( .A1(n19573), .A2(n19758), .ZN(n19628) );
  INV_X1 U13165 ( .A(n19687), .ZN(n19655) );
  INV_X1 U13166 ( .A(n19711), .ZN(n19718) );
  INV_X1 U13167 ( .A(n19745), .ZN(n19742) );
  INV_X1 U13168 ( .A(n19767), .ZN(n19778) );
  NAND2_X1 U13169 ( .A1(n19758), .A2(n19757), .ZN(n19803) );
  OR2_X1 U13170 ( .A1(n19978), .A2(n19811), .ZN(n19838) );
  INV_X1 U13171 ( .A(n19867), .ZN(n19864) );
  INV_X1 U13172 ( .A(n19902), .ZN(n19895) );
  INV_X1 U13173 ( .A(n20060), .ZN(n19933) );
  INV_X1 U13174 ( .A(n20054), .ZN(n19968) );
  OR2_X1 U13175 ( .A1(n19941), .A2(n19940), .ZN(n20013) );
  OR2_X1 U13176 ( .A1(n19941), .A2(n20020), .ZN(n20064) );
  INV_X1 U13177 ( .A(n20158), .ZN(n20085) );
  NAND2_X1 U13178 ( .A1(n19202), .A2(n17727), .ZN(n19200) );
  NAND2_X1 U13179 ( .A1(n19180), .A2(n19025), .ZN(n16856) );
  INV_X1 U13180 ( .A(n17192), .ZN(n17206) );
  INV_X1 U13181 ( .A(n17220), .ZN(n17209) );
  NOR2_X1 U13182 ( .A1(n17233), .A2(n17232), .ZN(n17262) );
  INV_X1 U13183 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17540) );
  INV_X1 U13184 ( .A(n17638), .ZN(n17648) );
  INV_X1 U13185 ( .A(n17722), .ZN(n17684) );
  AND2_X1 U13186 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17688), .ZN(n17682) );
  INV_X1 U13187 ( .A(n17718), .ZN(n17713) );
  INV_X1 U13188 ( .A(n17745), .ZN(n17763) );
  INV_X1 U13189 ( .A(n17914), .ZN(n17989) );
  INV_X1 U13190 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18392) );
  INV_X1 U13191 ( .A(n9729), .ZN(n18179) );
  INV_X1 U13192 ( .A(n18489), .ZN(n18495) );
  INV_X1 U13193 ( .A(n18413), .ZN(n18345) );
  NOR2_X1 U13194 ( .A1(n18347), .A2(n18346), .ZN(n18402) );
  OAI21_X2 U13195 ( .B1(n11202), .B2(n11201), .A(n19180), .ZN(n18494) );
  INV_X1 U13196 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19008) );
  INV_X1 U13197 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19018) );
  INV_X1 U13198 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n18579) );
  INV_X1 U13199 ( .A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n18746) );
  INV_X1 U13200 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n18749) );
  INV_X1 U13201 ( .A(n17176), .ZN(n19045) );
  NOR2_X1 U13202 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19189) );
  INV_X1 U13203 ( .A(n19135), .ZN(n19049) );
  INV_X1 U13204 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n19063) );
  NAND2_X1 U13205 ( .A1(n19063), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19194) );
  OAI21_X1 U13206 ( .B1(n12787), .B2(n15040), .A(n12786), .ZN(P1_U2842) );
  OAI211_X1 U13207 ( .C1(n15301), .C2(n20238), .A(n13334), .B(n9756), .ZN(
        P1_U2970) );
  INV_X1 U13208 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11458) );
  AND2_X4 U13209 ( .A1(n10368), .A2(n14006), .ZN(n13134) );
  AOI22_X1 U13210 ( .A1(n9737), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n13134), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10122) );
  INV_X2 U13211 ( .A(n10142), .ZN(n10372) );
  AOI22_X1 U13212 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10188), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10121) );
  INV_X1 U13213 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10118) );
  AOI22_X1 U13214 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10194), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10120) );
  INV_X2 U13215 ( .A(n13106), .ZN(n10358) );
  NAND4_X1 U13216 ( .A1(n10122), .A2(n10121), .A3(n10120), .A4(n10119), .ZN(
        n10123) );
  NAND2_X1 U13217 ( .A1(n10123), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10130) );
  AOI22_X1 U13218 ( .A1(n9737), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n13134), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10127) );
  AOI22_X1 U13219 ( .A1(n9721), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10194), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10126) );
  AOI22_X1 U13220 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10188), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10124) );
  NAND4_X1 U13221 ( .A1(n10127), .A2(n10126), .A3(n10125), .A4(n10124), .ZN(
        n10128) );
  NAND2_X1 U13222 ( .A1(n10128), .A2(n10359), .ZN(n10129) );
  AOI22_X1 U13223 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13134), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10134) );
  AOI22_X1 U13224 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10188), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10131) );
  AOI22_X1 U13225 ( .A1(n14000), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n10358), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U13226 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10194), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10132) );
  NAND4_X1 U13227 ( .A1(n10134), .A2(n10097), .A3(n10133), .A4(n10132), .ZN(
        n10140) );
  AOI22_X1 U13228 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13134), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10138) );
  AOI22_X1 U13229 ( .A1(n14000), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n13090), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10137) );
  AOI22_X1 U13230 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10188), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10135) );
  NAND3_X1 U13231 ( .A1(n10138), .A2(n10137), .A3(n10105), .ZN(n10139) );
  INV_X1 U13232 ( .A(n10225), .ZN(n10141) );
  AOI22_X1 U13233 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13134), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10144) );
  INV_X2 U13234 ( .A(n10142), .ZN(n12983) );
  AOI22_X1 U13235 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10188), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10143) );
  AND2_X1 U13236 ( .A1(n10144), .A2(n10143), .ZN(n10147) );
  AOI22_X1 U13237 ( .A1(n9686), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10194), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U13238 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n14000), .B1(
        n10358), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10145) );
  NAND3_X1 U13239 ( .A1(n10147), .A2(n10146), .A3(n10145), .ZN(n10148) );
  NAND2_X1 U13240 ( .A1(n10148), .A2(n10359), .ZN(n10155) );
  AOI22_X1 U13241 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n13134), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10152) );
  AOI22_X1 U13242 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10188), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U13243 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9668), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10150) );
  AOI22_X1 U13244 ( .A1(n14000), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10358), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10149) );
  NAND4_X1 U13245 ( .A1(n10152), .A2(n10151), .A3(n10150), .A4(n10149), .ZN(
        n10153) );
  AOI22_X1 U13246 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10194), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U13247 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10188), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U13248 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13134), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U13249 ( .A1(n14000), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9665), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10156) );
  NAND4_X1 U13250 ( .A1(n10159), .A2(n10158), .A3(n10157), .A4(n10156), .ZN(
        n10160) );
  NAND2_X1 U13251 ( .A1(n10160), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10167) );
  AOI22_X1 U13252 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n13134), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U13253 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n10188), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10163) );
  AOI22_X1 U13254 ( .A1(n9721), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n9668), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U13255 ( .A1(n14000), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13090), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10161) );
  NAND4_X1 U13256 ( .A1(n10164), .A2(n10163), .A3(n10162), .A4(n10161), .ZN(
        n10165) );
  NAND2_X1 U13257 ( .A1(n10165), .A2(n10359), .ZN(n10166) );
  NAND2_X1 U13258 ( .A1(n11352), .A2(n10094), .ZN(n10206) );
  AOI22_X1 U13259 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n13134), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10171) );
  AOI22_X1 U13260 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10188), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10170) );
  AOI22_X1 U13261 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10194), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10169) );
  AOI22_X1 U13262 ( .A1(n9665), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_7__5__SCAN_IN), .B2(n14000), .ZN(n10168) );
  NAND4_X1 U13263 ( .A1(n10171), .A2(n10170), .A3(n10169), .A4(n10168), .ZN(
        n10172) );
  NAND2_X1 U13264 ( .A1(n10172), .A2(n10359), .ZN(n10179) );
  AOI22_X1 U13265 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13134), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10176) );
  AOI22_X1 U13266 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10188), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10175) );
  AOI22_X1 U13267 ( .A1(n9665), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14000), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10173) );
  NAND4_X1 U13268 ( .A1(n10176), .A2(n10175), .A3(n10174), .A4(n10173), .ZN(
        n10177) );
  NAND2_X1 U13269 ( .A1(n10177), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10178) );
  AOI22_X1 U13270 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13134), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10183) );
  AOI22_X1 U13271 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10188), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10182) );
  AOI22_X1 U13272 ( .A1(n9721), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10194), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10181) );
  AOI22_X1 U13273 ( .A1(n14000), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9666), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U13274 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n13134), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U13275 ( .A1(n9721), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10194), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10186) );
  AOI22_X1 U13276 ( .A1(n14000), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9666), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U13277 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10188), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10184) );
  NAND2_X1 U13278 ( .A1(n11389), .A2(n10203), .ZN(n10202) );
  AOI22_X1 U13279 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n13134), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10192) );
  AOI22_X1 U13280 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10188), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10191) );
  AOI22_X1 U13281 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10194), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10190) );
  AOI22_X1 U13282 ( .A1(n10358), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_7__3__SCAN_IN), .B2(n14000), .ZN(n10189) );
  NAND4_X1 U13283 ( .A1(n10192), .A2(n10191), .A3(n10190), .A4(n10189), .ZN(
        n10193) );
  NAND2_X1 U13284 ( .A1(n10193), .A2(n10359), .ZN(n10201) );
  AOI22_X1 U13285 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13134), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10198) );
  AOI22_X1 U13286 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10188), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10197) );
  AOI22_X1 U13287 ( .A1(n9721), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10194), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U13288 ( .A1(n14000), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13090), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10195) );
  NAND4_X1 U13289 ( .A1(n10198), .A2(n10197), .A3(n10196), .A4(n10195), .ZN(
        n10199) );
  NAND2_X1 U13290 ( .A1(n10199), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10200) );
  NOR2_X2 U13291 ( .A1(n10206), .A2(n10205), .ZN(n11383) );
  AOI22_X1 U13292 ( .A1(n9686), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10194), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10210) );
  AOI22_X1 U13293 ( .A1(n14000), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10358), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10209) );
  AOI22_X1 U13294 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13134), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10208) );
  AOI22_X1 U13295 ( .A1(n10372), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10188), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10207) );
  NAND4_X1 U13296 ( .A1(n10210), .A2(n10209), .A3(n10208), .A4(n10207), .ZN(
        n10211) );
  NAND2_X1 U13297 ( .A1(n10211), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10218) );
  AOI22_X1 U13298 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10194), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10215) );
  AOI22_X1 U13299 ( .A1(n12983), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10188), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10214) );
  AOI22_X1 U13300 ( .A1(n9737), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n13134), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U13301 ( .A1(n14000), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n13090), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10212) );
  NAND4_X1 U13302 ( .A1(n10215), .A2(n10214), .A3(n10213), .A4(n10212), .ZN(
        n10216) );
  NAND2_X1 U13303 ( .A1(n10216), .A2(n10359), .ZN(n10217) );
  INV_X1 U13304 ( .A(n10271), .ZN(n10226) );
  NAND2_X1 U13305 ( .A1(n11383), .A2(n10226), .ZN(n10274) );
  AND2_X2 U13306 ( .A1(n10220), .A2(n10242), .ZN(n10244) );
  INV_X1 U13307 ( .A(n10256), .ZN(n10222) );
  NAND2_X1 U13308 ( .A1(n10222), .A2(n9730), .ZN(n13994) );
  AND2_X1 U13309 ( .A1(n11315), .A2(n10248), .ZN(n10223) );
  AND2_X2 U13310 ( .A1(n11390), .A2(n10236), .ZN(n13187) );
  NAND4_X1 U13311 ( .A1(n10223), .A2(n19543), .A3(n13187), .A4(n11288), .ZN(
        n10237) );
  INV_X1 U13312 ( .A(n10237), .ZN(n10224) );
  NAND3_X1 U13313 ( .A1(n13173), .A2(n19551), .A3(n13187), .ZN(n10227) );
  AND2_X2 U13314 ( .A1(n11314), .A2(n10227), .ZN(n10257) );
  NAND3_X1 U13315 ( .A1(n10274), .A2(n13994), .A3(n10257), .ZN(n10228) );
  NAND2_X1 U13316 ( .A1(n10228), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10284) );
  INV_X2 U13317 ( .A(n11390), .ZN(n19565) );
  AND2_X2 U13318 ( .A1(n10254), .A2(n10244), .ZN(n10298) );
  NAND2_X1 U13319 ( .A1(n10298), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10231) );
  NAND2_X1 U13320 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10230) );
  OAI211_X1 U13321 ( .C1(n9657), .C2(n14320), .A(n10231), .B(n10230), .ZN(
        n10232) );
  NAND2_X1 U13322 ( .A1(n10235), .A2(n10234), .ZN(n10239) );
  NAND2_X1 U13323 ( .A1(n11360), .A2(n10240), .ZN(n10241) );
  NAND2_X1 U13324 ( .A1(n10241), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10247) );
  INV_X1 U13325 ( .A(n13187), .ZN(n13192) );
  NOR2_X1 U13326 ( .A1(n13192), .A2(n9685), .ZN(n10243) );
  NAND2_X1 U13327 ( .A1(n10243), .A2(n10242), .ZN(n10642) );
  NAND2_X1 U13328 ( .A1(n11384), .A2(n20224), .ZN(n10246) );
  AND2_X2 U13329 ( .A1(n10247), .A2(n10246), .ZN(n10264) );
  XNOR2_X1 U13330 ( .A(n10248), .B(n13746), .ZN(n11322) );
  AOI21_X1 U13331 ( .B1(n10249), .B2(n11321), .A(n19565), .ZN(n10250) );
  OAI21_X1 U13332 ( .B1(n11322), .B2(n11321), .A(n10250), .ZN(n11348) );
  NAND2_X1 U13333 ( .A1(n11348), .A2(n11350), .ZN(n10253) );
  NAND2_X1 U13334 ( .A1(n10268), .A2(n10254), .ZN(n10255) );
  NAND2_X1 U13335 ( .A1(n10292), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10259) );
  NOR2_X1 U13336 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U13337 ( .A1(n11344), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n10260), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10258) );
  XNOR2_X1 U13338 ( .A(n10280), .B(n10279), .ZN(n10318) );
  INV_X1 U13339 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n11392) );
  INV_X1 U13340 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n14344) );
  NAND2_X1 U13341 ( .A1(n10298), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10263) );
  INV_X1 U13342 ( .A(n10260), .ZN(n13995) );
  NAND2_X1 U13343 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10261) );
  AND2_X1 U13344 ( .A1(n13995), .A2(n10261), .ZN(n10262) );
  OAI211_X1 U13345 ( .C1(n9657), .C2(n14344), .A(n10263), .B(n10262), .ZN(
        n10266) );
  INV_X1 U13346 ( .A(n10264), .ZN(n10265) );
  NOR2_X1 U13347 ( .A1(n10266), .A2(n10265), .ZN(n10270) );
  NAND3_X1 U13348 ( .A1(n10268), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10267), 
        .ZN(n10269) );
  OAI211_X1 U13349 ( .C1(n10284), .C2(n11392), .A(n10270), .B(n10269), .ZN(
        n10315) );
  NOR2_X1 U13350 ( .A1(n10272), .A2(n10271), .ZN(n10273) );
  OAI22_X1 U13351 ( .A1(n9692), .A2(n10273), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n9659), .ZN(n10278) );
  INV_X1 U13352 ( .A(n11345), .ZN(n10276) );
  NOR2_X1 U13353 ( .A1(n13995), .A2(n20202), .ZN(n10275) );
  AOI21_X1 U13354 ( .B1(n10276), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10275), 
        .ZN(n10277) );
  NAND2_X1 U13355 ( .A1(n10278), .A2(n10277), .ZN(n10316) );
  NAND2_X1 U13356 ( .A1(n10318), .A2(n10314), .ZN(n10283) );
  INV_X1 U13357 ( .A(n10279), .ZN(n10281) );
  NAND2_X1 U13358 ( .A1(n10281), .A2(n10280), .ZN(n10282) );
  INV_X1 U13359 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10290) );
  INV_X1 U13360 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10287) );
  NAND2_X1 U13361 ( .A1(n10298), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10286) );
  NAND2_X1 U13362 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10285) );
  INV_X1 U13363 ( .A(n10288), .ZN(n10289) );
  INV_X1 U13364 ( .A(n10291), .ZN(n10311) );
  NAND2_X1 U13365 ( .A1(n9692), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10294) );
  AOI21_X1 U13366 ( .B1(n20218), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10293) );
  NAND2_X1 U13367 ( .A1(n10291), .A2(n10310), .ZN(n10295) );
  NAND2_X1 U13368 ( .A1(n10296), .A2(n10311), .ZN(n10297) );
  INV_X1 U13369 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10301) );
  NAND2_X1 U13370 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10299) );
  OAI211_X1 U13371 ( .C1(n9657), .C2(n10301), .A(n10300), .B(n10299), .ZN(
        n10302) );
  INV_X1 U13372 ( .A(n10306), .ZN(n10305) );
  NOR2_X1 U13373 ( .A1(n13995), .A2(n20175), .ZN(n10303) );
  AOI21_X1 U13374 ( .B1(n9692), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n10303), .ZN(n10307) );
  INV_X1 U13375 ( .A(n10307), .ZN(n10304) );
  NAND2_X1 U13376 ( .A1(n10305), .A2(n10304), .ZN(n10308) );
  INV_X1 U13377 ( .A(n9734), .ZN(n10313) );
  XNOR2_X2 U13378 ( .A(n10309), .B(n10312), .ZN(n12788) );
  NAND2_X2 U13379 ( .A1(n10313), .A2(n12788), .ZN(n10329) );
  OR2_X1 U13380 ( .A1(n10316), .A2(n10315), .ZN(n10317) );
  AND2_X1 U13382 ( .A1(n14346), .A2(n10321), .ZN(n10345) );
  INV_X1 U13383 ( .A(n19749), .ZN(n10490) );
  INV_X1 U13384 ( .A(n10321), .ZN(n10319) );
  OR2_X2 U13385 ( .A1(n10329), .A2(n10330), .ZN(n19692) );
  INV_X1 U13386 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10320) );
  OAI22_X1 U13387 ( .A1(n11458), .A2(n10490), .B1(n19692), .B2(n10320), .ZN(
        n10325) );
  INV_X1 U13388 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12843) );
  OR2_X2 U13389 ( .A1(n9734), .A2(n12788), .ZN(n10351) );
  XNOR2_X2 U13390 ( .A(n10322), .B(n10321), .ZN(n14327) );
  NAND2_X1 U13391 ( .A1(n14327), .A2(n13467), .ZN(n10328) );
  OR2_X2 U13392 ( .A1(n10351), .A2(n10328), .ZN(n10492) );
  OR3_X2 U13393 ( .A1(n10341), .A2(n12788), .A3(n14327), .ZN(n10487) );
  INV_X1 U13394 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10323) );
  NOR2_X1 U13395 ( .A1(n10325), .A2(n10324), .ZN(n10339) );
  INV_X1 U13396 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10327) );
  OR2_X1 U13397 ( .A1(n14346), .A2(n14327), .ZN(n10326) );
  OR2_X2 U13398 ( .A1(n10329), .A2(n10326), .ZN(n19664) );
  OR2_X2 U13399 ( .A1(n10351), .A2(n10326), .ZN(n19525) );
  OAI22_X1 U13400 ( .A1(n10327), .A2(n19664), .B1(n19525), .B2(n19537), .ZN(
        n10332) );
  INV_X1 U13401 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11470) );
  INV_X1 U13402 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13014) );
  OAI22_X1 U13403 ( .A1(n11470), .A2(n19721), .B1(n19576), .B2(n13014), .ZN(
        n10331) );
  NOR2_X1 U13404 ( .A1(n10332), .A2(n10331), .ZN(n10338) );
  INV_X1 U13405 ( .A(n10341), .ZN(n10333) );
  NAND2_X1 U13406 ( .A1(n10333), .A2(n14327), .ZN(n10334) );
  INV_X1 U13407 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12845) );
  INV_X1 U13408 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12846) );
  NOR2_X1 U13409 ( .A1(n10336), .A2(n10335), .ZN(n10337) );
  NAND3_X1 U13410 ( .A1(n10339), .A2(n10338), .A3(n10337), .ZN(n10416) );
  INV_X1 U13411 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11457) );
  INV_X1 U13412 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13005) );
  OAI22_X1 U13413 ( .A1(n11457), .A2(n10480), .B1(n10486), .B2(n13005), .ZN(
        n10344) );
  INV_X1 U13414 ( .A(n10344), .ZN(n10349) );
  INV_X1 U13415 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11467) );
  INV_X1 U13416 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12844) );
  OAI22_X1 U13417 ( .A1(n11467), .A2(n19876), .B1(n10479), .B2(n12844), .ZN(
        n10347) );
  INV_X1 U13418 ( .A(n10347), .ZN(n10348) );
  NOR2_X2 U13419 ( .A1(n10351), .A2(n10350), .ZN(n19636) );
  INV_X1 U13420 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10355) );
  INV_X1 U13421 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10353) );
  OR2_X1 U13422 ( .A1(n20018), .A2(n10353), .ZN(n10354) );
  OAI211_X1 U13423 ( .C1(n19630), .C2(n10355), .A(n10354), .B(n15586), .ZN(
        n10356) );
  INV_X1 U13424 ( .A(n10356), .ZN(n10357) );
  AOI22_X1 U13425 ( .A1(n12960), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10367) );
  AOI22_X1 U13426 ( .A1(n12907), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12905), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10366) );
  INV_X1 U13427 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10362) );
  INV_X1 U13428 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10360) );
  OR2_X1 U13429 ( .A1(n12963), .A2(n10360), .ZN(n10361) );
  OAI21_X1 U13430 ( .B1(n12897), .B2(n10362), .A(n10361), .ZN(n10363) );
  INV_X1 U13431 ( .A(n10363), .ZN(n10365) );
  AOI22_X1 U13432 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12906), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10364) );
  NAND4_X1 U13433 ( .A1(n10367), .A2(n10366), .A3(n10365), .A4(n10364), .ZN(
        n10378) );
  AND2_X1 U13434 ( .A1(n10368), .A2(n12976), .ZN(n10460) );
  AOI22_X1 U13435 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10376) );
  NAND2_X1 U13436 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12977) );
  INV_X1 U13437 ( .A(n12977), .ZN(n10371) );
  AOI22_X1 U13438 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10375) );
  AND2_X1 U13439 ( .A1(n10016), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14039) );
  AOI22_X1 U13440 ( .A1(n10385), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10374) );
  AOI22_X1 U13441 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12904), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10373) );
  NAND4_X1 U13442 ( .A1(n10376), .A2(n10375), .A3(n10374), .A4(n10373), .ZN(
        n10377) );
  OR2_X1 U13443 ( .A1(n11395), .A2(n15586), .ZN(n13462) );
  INV_X1 U13444 ( .A(n13462), .ZN(n10394) );
  NAND2_X1 U13445 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10380) );
  NAND2_X1 U13446 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10379) );
  OAI211_X1 U13447 ( .C1(n12963), .C2(n11470), .A(n10380), .B(n10379), .ZN(
        n10382) );
  OAI22_X1 U13448 ( .A1(n12897), .A2(n12846), .B1(n12896), .B2(n11458), .ZN(
        n10381) );
  NOR2_X1 U13449 ( .A1(n10382), .A2(n10381), .ZN(n10393) );
  AOI22_X1 U13450 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10460), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U13451 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10384), .B1(
        n10385), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U13452 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10396), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10387) );
  NAND2_X1 U13453 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10386) );
  AND4_X1 U13454 ( .A1(n10389), .A2(n10388), .A3(n10387), .A4(n10386), .ZN(
        n10392) );
  AOI22_X1 U13455 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12905), .B1(
        n12904), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10391) );
  INV_X1 U13456 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19537) );
  AOI22_X1 U13457 ( .A1(n12907), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12906), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10390) );
  NAND4_X1 U13458 ( .A1(n10393), .A2(n10392), .A3(n10391), .A4(n10390), .ZN(
        n11402) );
  NAND2_X1 U13459 ( .A1(n10394), .A2(n11402), .ZN(n10582) );
  AOI22_X1 U13460 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10460), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10400) );
  AOI22_X1 U13461 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10384), .B1(
        n10385), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10399) );
  AOI22_X1 U13462 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10395), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10398) );
  NAND2_X1 U13463 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10397) );
  NAND4_X1 U13464 ( .A1(n10400), .A2(n10399), .A3(n10398), .A4(n10397), .ZN(
        n10406) );
  NAND2_X1 U13465 ( .A1(n12907), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10404) );
  NAND2_X1 U13466 ( .A1(n12905), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10403) );
  NAND2_X1 U13467 ( .A1(n12904), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10402) );
  NAND2_X1 U13468 ( .A1(n12906), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10401) );
  NAND4_X1 U13469 ( .A1(n10404), .A2(n10403), .A3(n10402), .A4(n10401), .ZN(
        n10405) );
  NOR2_X1 U13470 ( .A1(n10406), .A2(n10405), .ZN(n10413) );
  INV_X1 U13471 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10409) );
  NAND2_X1 U13472 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10408) );
  NAND2_X1 U13473 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10407) );
  OAI211_X1 U13474 ( .C1(n12963), .C2(n10409), .A(n10408), .B(n10407), .ZN(
        n10411) );
  INV_X1 U13475 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12864) );
  INV_X1 U13476 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11481) );
  OAI22_X1 U13477 ( .A1(n12897), .A2(n12864), .B1(n12896), .B2(n11481), .ZN(
        n10410) );
  NOR2_X1 U13478 ( .A1(n10411), .A2(n10410), .ZN(n10412) );
  NAND2_X1 U13479 ( .A1(n10582), .A2(n10643), .ZN(n10414) );
  INV_X1 U13480 ( .A(n10579), .ZN(n10459) );
  INV_X1 U13481 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12882) );
  NAND2_X1 U13482 ( .A1(n19749), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10418) );
  NAND2_X1 U13483 ( .A1(n19636), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10417) );
  NOR2_X1 U13484 ( .A1(n10419), .A2(n9730), .ZN(n10435) );
  INV_X1 U13485 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10439) );
  INV_X1 U13486 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12880) );
  OAI22_X1 U13487 ( .A1(n10439), .A2(n19525), .B1(n10492), .B2(n12880), .ZN(
        n10421) );
  INV_X1 U13488 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13060) );
  INV_X1 U13489 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11513) );
  NOR2_X1 U13490 ( .A1(n10421), .A2(n10420), .ZN(n10434) );
  INV_X1 U13491 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11512) );
  INV_X1 U13492 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10422) );
  OAI22_X1 U13493 ( .A1(n11512), .A2(n19876), .B1(n10480), .B2(n10422), .ZN(
        n10425) );
  INV_X1 U13494 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10423) );
  INV_X1 U13495 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13062) );
  OAI22_X1 U13496 ( .A1(n10423), .A2(n20018), .B1(n10479), .B2(n13062), .ZN(
        n10424) );
  INV_X1 U13497 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12881) );
  NOR2_X1 U13498 ( .A1(n10483), .A2(n12881), .ZN(n10426) );
  NOR2_X1 U13499 ( .A1(n10427), .A2(n10426), .ZN(n10433) );
  INV_X1 U13500 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10446) );
  INV_X1 U13501 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10428) );
  OAI22_X1 U13502 ( .A1(n10446), .A2(n19721), .B1(n19692), .B2(n10428), .ZN(
        n10431) );
  INV_X1 U13503 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10429) );
  INV_X1 U13504 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13054) );
  NOR2_X1 U13505 ( .A1(n10431), .A2(n10430), .ZN(n10432) );
  NAND4_X1 U13506 ( .A1(n10435), .A2(n10434), .A3(n10433), .A4(n10432), .ZN(
        n10457) );
  OAI22_X1 U13507 ( .A1(n13060), .A2(n12956), .B1(n12955), .B2(n11513), .ZN(
        n10438) );
  AOI22_X1 U13508 ( .A1(n12961), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12960), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10436) );
  OAI22_X1 U13509 ( .A1(n12953), .A2(n11512), .B1(n12951), .B2(n10439), .ZN(
        n10451) );
  AOI22_X1 U13510 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10460), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10443) );
  AOI22_X1 U13511 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10384), .B1(
        n10385), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10442) );
  AOI22_X1 U13512 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10395), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10441) );
  NAND2_X1 U13513 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10440) );
  AND4_X1 U13514 ( .A1(n10443), .A2(n10442), .A3(n10441), .A4(n10440), .ZN(
        n10449) );
  NAND2_X1 U13515 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10445) );
  NAND2_X1 U13516 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10444) );
  OAI211_X1 U13517 ( .C1(n12963), .C2(n10446), .A(n10445), .B(n10444), .ZN(
        n10447) );
  INV_X1 U13518 ( .A(n10447), .ZN(n10448) );
  INV_X1 U13519 ( .A(n11416), .ZN(n10455) );
  NAND2_X1 U13520 ( .A1(n10455), .A2(n9730), .ZN(n10456) );
  AOI22_X1 U13521 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10460), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10464) );
  AOI22_X1 U13522 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10384), .B1(
        n10385), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10463) );
  AOI22_X1 U13523 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10395), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U13524 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10461) );
  AND4_X1 U13525 ( .A1(n10464), .A2(n10463), .A3(n10462), .A4(n10461), .ZN(
        n10476) );
  INV_X1 U13526 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10465) );
  INV_X1 U13527 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12894) );
  OAI22_X1 U13528 ( .A1(n12963), .A2(n10465), .B1(n12956), .B2(n12894), .ZN(
        n10468) );
  INV_X1 U13529 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11529) );
  INV_X1 U13530 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10466) );
  OAI22_X1 U13531 ( .A1(n11529), .A2(n12896), .B1(n12955), .B2(n10466), .ZN(
        n10467) );
  NOR2_X1 U13532 ( .A1(n10468), .A2(n10467), .ZN(n10475) );
  AOI22_X1 U13533 ( .A1(n12907), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12906), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10474) );
  INV_X1 U13534 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10471) );
  NAND2_X1 U13535 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10470) );
  NAND2_X1 U13536 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10469) );
  OAI211_X1 U13537 ( .C1(n12897), .C2(n10471), .A(n10470), .B(n10469), .ZN(
        n10472) );
  INV_X1 U13538 ( .A(n10472), .ZN(n10473) );
  NAND4_X1 U13539 ( .A1(n10476), .A2(n10475), .A3(n10474), .A4(n10473), .ZN(
        n11420) );
  INV_X1 U13540 ( .A(n11420), .ZN(n10477) );
  INV_X1 U13541 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10478) );
  INV_X1 U13542 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13116) );
  OAI22_X1 U13543 ( .A1(n10478), .A2(n9653), .B1(n19876), .B2(n13116), .ZN(
        n10482) );
  INV_X1 U13544 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13117) );
  INV_X1 U13545 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11556) );
  OAI22_X1 U13546 ( .A1(n13117), .A2(n10479), .B1(n10480), .B2(n11556), .ZN(
        n10481) );
  OR2_X1 U13547 ( .A1(n10482), .A2(n10481), .ZN(n10485) );
  INV_X1 U13548 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12916) );
  NOR2_X1 U13549 ( .A1(n10483), .A2(n12916), .ZN(n10484) );
  NOR2_X1 U13550 ( .A1(n10485), .A2(n10484), .ZN(n10501) );
  INV_X1 U13551 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10504) );
  INV_X1 U13552 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13107) );
  OAI22_X1 U13553 ( .A1(n10504), .A2(n19721), .B1(n19576), .B2(n13107), .ZN(
        n10489) );
  INV_X1 U13554 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11549) );
  INV_X1 U13555 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13114) );
  OAI22_X1 U13556 ( .A1(n11549), .A2(n10486), .B1(n10487), .B2(n13114), .ZN(
        n10488) );
  NOR2_X1 U13557 ( .A1(n10489), .A2(n10488), .ZN(n10500) );
  INV_X1 U13558 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10491) );
  INV_X1 U13559 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11548) );
  OAI22_X1 U13560 ( .A1(n10491), .A2(n19664), .B1(n10490), .B2(n11548), .ZN(
        n10494) );
  INV_X1 U13561 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13105) );
  INV_X1 U13562 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13104) );
  OAI22_X1 U13563 ( .A1(n13105), .A2(n10492), .B1(n19525), .B2(n13104), .ZN(
        n10493) );
  NOR2_X1 U13564 ( .A1(n10494), .A2(n10493), .ZN(n10499) );
  INV_X1 U13565 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12917) );
  INV_X1 U13566 ( .A(n19692), .ZN(n19695) );
  NAND2_X1 U13567 ( .A1(n19695), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10496) );
  NAND2_X1 U13568 ( .A1(n19636), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10495) );
  OAI211_X1 U13569 ( .C1(n9750), .C2(n12917), .A(n10496), .B(n10495), .ZN(
        n10497) );
  INV_X1 U13570 ( .A(n10497), .ZN(n10498) );
  NAND4_X1 U13571 ( .A1(n10501), .A2(n10500), .A3(n10499), .A4(n10498), .ZN(
        n10517) );
  NAND2_X1 U13572 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10503) );
  NAND2_X1 U13573 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10502) );
  OAI211_X1 U13574 ( .C1(n12963), .C2(n10504), .A(n10503), .B(n10502), .ZN(
        n10506) );
  OAI22_X1 U13575 ( .A1(n12897), .A2(n12917), .B1(n12896), .B2(n11548), .ZN(
        n10505) );
  NOR2_X1 U13576 ( .A1(n10506), .A2(n10505), .ZN(n10514) );
  AOI22_X1 U13577 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10460), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10510) );
  AOI22_X1 U13578 ( .A1(n10385), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10509) );
  AOI22_X1 U13579 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10508) );
  NAND2_X1 U13580 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10507) );
  AND4_X1 U13581 ( .A1(n10510), .A2(n10509), .A3(n10508), .A4(n10507), .ZN(
        n10513) );
  AOI22_X1 U13582 ( .A1(n12905), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12904), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10512) );
  AOI22_X1 U13583 ( .A1(n12907), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12906), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10511) );
  NAND4_X1 U13584 ( .A1(n10514), .A2(n10513), .A3(n10512), .A4(n10511), .ZN(
        n11426) );
  INV_X1 U13585 ( .A(n11426), .ZN(n10515) );
  NAND2_X1 U13586 ( .A1(n10515), .A2(n9730), .ZN(n10516) );
  INV_X1 U13587 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10518) );
  INV_X1 U13588 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13127) );
  OAI22_X1 U13589 ( .A1(n10518), .A2(n20018), .B1(n10479), .B2(n13127), .ZN(
        n10521) );
  INV_X1 U13590 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10519) );
  INV_X1 U13591 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11574) );
  OAI22_X1 U13592 ( .A1(n10519), .A2(n19876), .B1(n10480), .B2(n11574), .ZN(
        n10520) );
  OR2_X1 U13593 ( .A1(n10521), .A2(n10520), .ZN(n10523) );
  INV_X1 U13594 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12934) );
  NOR2_X1 U13595 ( .A1(n10483), .A2(n12934), .ZN(n10522) );
  NOR2_X1 U13596 ( .A1(n10523), .A2(n10522), .ZN(n10537) );
  INV_X1 U13597 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13837) );
  INV_X1 U13598 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10524) );
  OAI22_X1 U13599 ( .A1(n13837), .A2(n19525), .B1(n10492), .B2(n10524), .ZN(
        n10527) );
  INV_X1 U13600 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10525) );
  INV_X1 U13601 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11573) );
  OAI22_X1 U13602 ( .A1(n10525), .A2(n10487), .B1(n10486), .B2(n11573), .ZN(
        n10526) );
  NOR2_X1 U13603 ( .A1(n10527), .A2(n10526), .ZN(n10536) );
  INV_X1 U13604 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10548) );
  INV_X1 U13605 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10528) );
  OAI22_X1 U13606 ( .A1(n10548), .A2(n19721), .B1(n19692), .B2(n10528), .ZN(
        n10530) );
  INV_X1 U13607 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11572) );
  INV_X1 U13608 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13131) );
  OAI22_X1 U13609 ( .A1(n11572), .A2(n19576), .B1(n19664), .B2(n13131), .ZN(
        n10529) );
  NOR2_X1 U13610 ( .A1(n10530), .A2(n10529), .ZN(n10535) );
  INV_X1 U13611 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12935) );
  NAND2_X1 U13612 ( .A1(n19749), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10532) );
  NAND2_X1 U13613 ( .A1(n19636), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10531) );
  OAI211_X1 U13614 ( .C1(n9750), .C2(n12935), .A(n10532), .B(n10531), .ZN(
        n10533) );
  INV_X1 U13615 ( .A(n10533), .ZN(n10534) );
  NAND4_X1 U13616 ( .A1(n10537), .A2(n10536), .A3(n10535), .A4(n10534), .ZN(
        n10556) );
  AOI22_X1 U13617 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10460), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10541) );
  AOI22_X1 U13618 ( .A1(n10385), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10540) );
  AOI22_X1 U13619 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10539) );
  NAND2_X1 U13620 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10538) );
  NAND4_X1 U13621 ( .A1(n10541), .A2(n10540), .A3(n10539), .A4(n10538), .ZN(
        n10547) );
  OR2_X1 U13622 ( .A1(n12897), .A2(n12935), .ZN(n10545) );
  NAND2_X1 U13623 ( .A1(n12906), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10544) );
  NAND2_X1 U13624 ( .A1(n12904), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n10543) );
  NAND2_X1 U13625 ( .A1(n12905), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10542) );
  NAND4_X1 U13626 ( .A1(n10545), .A2(n10544), .A3(n10543), .A4(n10542), .ZN(
        n10546) );
  NOR2_X1 U13627 ( .A1(n10547), .A2(n10546), .ZN(n10554) );
  AOI22_X1 U13628 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10552) );
  OR2_X1 U13629 ( .A1(n12963), .A2(n10548), .ZN(n10551) );
  NAND2_X1 U13630 ( .A1(n12907), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n10550) );
  NAND2_X1 U13631 ( .A1(n12960), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10549) );
  NAND2_X1 U13632 ( .A1(n9730), .A2(n11429), .ZN(n10555) );
  AOI22_X1 U13633 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10460), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U13634 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10384), .B1(
        n10385), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U13635 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10559) );
  NAND2_X1 U13636 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10558) );
  NAND2_X1 U13637 ( .A1(n12907), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10565) );
  NAND2_X1 U13638 ( .A1(n12904), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10564) );
  NAND2_X1 U13639 ( .A1(n12905), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10563) );
  NAND2_X1 U13640 ( .A1(n12906), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10562) );
  INV_X1 U13641 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12957) );
  INV_X1 U13642 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11591) );
  OAI22_X1 U13643 ( .A1(n12897), .A2(n12957), .B1(n12896), .B2(n11591), .ZN(
        n10566) );
  INV_X1 U13644 ( .A(n10566), .ZN(n10572) );
  INV_X1 U13645 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10569) );
  NAND2_X1 U13646 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10568) );
  NAND2_X1 U13647 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10567) );
  OAI211_X1 U13648 ( .C1(n12963), .C2(n10569), .A(n10568), .B(n10567), .ZN(
        n10570) );
  INV_X1 U13649 ( .A(n10570), .ZN(n10571) );
  NAND4_X2 U13650 ( .A1(n10574), .A2(n10573), .A3(n10572), .A4(n10571), .ZN(
        n14818) );
  NAND2_X1 U13651 ( .A1(n10575), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16640) );
  NAND2_X1 U13652 ( .A1(n14818), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10577) );
  NAND2_X1 U13653 ( .A1(n16640), .A2(n10612), .ZN(n10606) );
  NAND2_X1 U13654 ( .A1(n10579), .A2(n10580), .ZN(n10581) );
  XOR2_X1 U13655 ( .A(n10643), .B(n10582), .Z(n14756) );
  NAND2_X1 U13656 ( .A1(n13462), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13461) );
  XOR2_X1 U13657 ( .A(n11395), .B(n11402), .Z(n10583) );
  NOR2_X1 U13658 ( .A1(n13461), .A2(n10583), .ZN(n10585) );
  INV_X1 U13659 ( .A(n13461), .ZN(n10584) );
  XOR2_X1 U13660 ( .A(n10584), .B(n10583), .Z(n13477) );
  NOR2_X1 U13661 ( .A1(n14308), .A2(n13477), .ZN(n13476) );
  NOR2_X1 U13662 ( .A1(n10585), .A2(n13476), .ZN(n10586) );
  XOR2_X1 U13663 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10586), .Z(
        n14755) );
  NOR2_X1 U13664 ( .A1(n14756), .A2(n14755), .ZN(n14754) );
  NOR2_X1 U13665 ( .A1(n10586), .A2(n10290), .ZN(n10587) );
  OR2_X1 U13666 ( .A1(n14754), .A2(n10587), .ZN(n10588) );
  INV_X1 U13667 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14453) );
  XNOR2_X1 U13668 ( .A(n10588), .B(n14453), .ZN(n14377) );
  NAND2_X1 U13669 ( .A1(n10588), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10589) );
  NAND2_X1 U13670 ( .A1(n16086), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10594) );
  INV_X1 U13671 ( .A(n10590), .ZN(n10593) );
  NAND2_X1 U13672 ( .A1(n10591), .A2(n10477), .ZN(n10592) );
  NAND2_X1 U13673 ( .A1(n10593), .A2(n10592), .ZN(n16084) );
  NAND2_X1 U13674 ( .A1(n10594), .A2(n16084), .ZN(n10598) );
  INV_X1 U13675 ( .A(n16086), .ZN(n10596) );
  INV_X1 U13676 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10595) );
  NAND2_X1 U13677 ( .A1(n10596), .A2(n10595), .ZN(n10597) );
  INV_X1 U13678 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14462) );
  NAND2_X1 U13679 ( .A1(n10600), .A2(n14462), .ZN(n14444) );
  NAND2_X1 U13680 ( .A1(n10777), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14445) );
  XNOR2_X2 U13681 ( .A(n10601), .B(n10602), .ZN(n10808) );
  INV_X1 U13682 ( .A(n14445), .ZN(n14448) );
  NAND2_X1 U13683 ( .A1(n14448), .A2(n10602), .ZN(n10603) );
  INV_X1 U13684 ( .A(n10808), .ZN(n10604) );
  NAND3_X1 U13685 ( .A1(n10609), .A2(n15830), .A3(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10611) );
  NAND2_X1 U13686 ( .A1(n10605), .A2(n10604), .ZN(n15831) );
  NAND2_X1 U13687 ( .A1(n10609), .A2(n10608), .ZN(n10610) );
  INV_X1 U13688 ( .A(n10612), .ZN(n10614) );
  NAND2_X1 U13689 ( .A1(n16053), .A2(n10615), .ZN(n16035) );
  INV_X1 U13690 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16042) );
  NAND2_X1 U13691 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16004) );
  INV_X1 U13692 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16007) );
  NOR2_X1 U13693 ( .A1(n16004), .A2(n16007), .ZN(n11655) );
  AND2_X1 U13694 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15954) );
  AND2_X1 U13695 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10616) );
  NAND2_X1 U13696 ( .A1(n15954), .A2(n10616), .ZN(n11656) );
  NAND2_X1 U13697 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n13218) );
  INV_X1 U13698 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15906) );
  INV_X1 U13699 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15895) );
  INV_X1 U13700 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15884) );
  NAND2_X1 U13701 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15842) );
  INV_X1 U13702 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16273) );
  NOR2_X1 U13703 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n16273), .ZN(
        n10624) );
  NAND2_X1 U13704 ( .A1(n20193), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10619) );
  NAND2_X1 U13705 ( .A1(n14807), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10618) );
  NAND2_X1 U13706 ( .A1(n10619), .A2(n10618), .ZN(n11294) );
  NAND2_X1 U13707 ( .A1(n20182), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10626) );
  NAND2_X1 U13708 ( .A1(n10629), .A2(n10626), .ZN(n10621) );
  NAND2_X1 U13709 ( .A1(n14006), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10627) );
  INV_X1 U13710 ( .A(n10634), .ZN(n10625) );
  XNOR2_X1 U13711 ( .A(n11294), .B(n10625), .ZN(n11290) );
  NAND2_X1 U13712 ( .A1(n10627), .A2(n10626), .ZN(n10628) );
  XNOR2_X1 U13713 ( .A(n10629), .B(n10628), .ZN(n11299) );
  NAND3_X1 U13714 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10630), .A3(
        n13532), .ZN(n10647) );
  XNOR2_X1 U13715 ( .A(n10632), .B(n10631), .ZN(n10648) );
  NAND2_X1 U13716 ( .A1(n10647), .A2(n10648), .ZN(n11303) );
  NOR2_X1 U13717 ( .A1(n11299), .A2(n11303), .ZN(n10635) );
  AND2_X1 U13718 ( .A1(n11290), .A2(n10635), .ZN(n10633) );
  OAI21_X1 U13719 ( .B1(n20202), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n10634), .ZN(n11295) );
  INV_X1 U13720 ( .A(n11295), .ZN(n11291) );
  AOI21_X1 U13721 ( .B1(n11291), .B2(n10635), .A(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n10636) );
  NAND2_X1 U13722 ( .A1(n13408), .A2(n10636), .ZN(n10641) );
  NAND2_X1 U13723 ( .A1(n10637), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10638) );
  NAND2_X1 U13724 ( .A1(n10638), .A2(n13532), .ZN(n14028) );
  INV_X1 U13725 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n19213) );
  OAI21_X1 U13726 ( .B1(n10383), .B2(n14028), .A(n19213), .ZN(n10639) );
  AND2_X1 U13727 ( .A1(n10639), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n20199) );
  INV_X1 U13728 ( .A(n20199), .ZN(n10640) );
  OR2_X1 U13729 ( .A1(n10642), .A2(n9730), .ZN(n10652) );
  INV_X1 U13730 ( .A(n11299), .ZN(n10644) );
  INV_X1 U13731 ( .A(n10643), .ZN(n11409) );
  MUX2_X1 U13732 ( .A(n10644), .B(n11409), .S(n10646), .Z(n10759) );
  NOR2_X1 U13733 ( .A1(n11294), .A2(n11295), .ZN(n10645) );
  NOR2_X1 U13734 ( .A1(n10759), .A2(n10645), .ZN(n10650) );
  MUX2_X1 U13735 ( .A(n10647), .B(n11420), .S(n10646), .Z(n10765) );
  MUX2_X1 U13736 ( .A(n11416), .B(n10648), .S(n11336), .Z(n10762) );
  NAND2_X1 U13737 ( .A1(n10765), .A2(n10762), .ZN(n11289) );
  INV_X1 U13738 ( .A(n11309), .ZN(n10649) );
  OAI21_X1 U13739 ( .B1(n10650), .B2(n11289), .A(n10649), .ZN(n20205) );
  AND2_X1 U13740 ( .A1(n10221), .A2(n9730), .ZN(n11319) );
  INV_X1 U13741 ( .A(n11319), .ZN(n10651) );
  OR2_X1 U13742 ( .A1(n10642), .A2(n10651), .ZN(n11339) );
  OAI22_X1 U13743 ( .A1(n20208), .A2(n10652), .B1(n20205), .B2(n11339), .ZN(
        n11331) );
  AND2_X1 U13744 ( .A1(n14795), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14196) );
  NOR2_X1 U13745 ( .A1(n19522), .A2(n19210), .ZN(n10653) );
  INV_X1 U13746 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n16490) );
  NAND2_X1 U13747 ( .A1(n11340), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n10656) );
  NAND2_X1 U13748 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10655) );
  OAI211_X1 U13749 ( .C1(n10747), .C2(n16490), .A(n10656), .B(n10655), .ZN(
        n10657) );
  AOI21_X1 U13750 ( .B1(n10654), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n10657), .ZN(n10749) );
  INV_X1 U13751 ( .A(n10658), .ZN(n10659) );
  INV_X1 U13752 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14222) );
  OR2_X1 U13753 ( .A1(n10662), .A2(n10595), .ZN(n10664) );
  AOI22_X1 U13754 ( .A1(n11340), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10663) );
  OAI211_X1 U13755 ( .C1(n10747), .C2(n14222), .A(n10664), .B(n10663), .ZN(
        n13754) );
  NAND2_X1 U13756 ( .A1(n13755), .A2(n13754), .ZN(n14455) );
  OR2_X1 U13757 ( .A1(n10662), .A2(n14462), .ZN(n10669) );
  INV_X1 U13758 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n14790) );
  NAND2_X1 U13759 ( .A1(n11340), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n10666) );
  NAND2_X1 U13760 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10665) );
  OAI211_X1 U13761 ( .C1(n10747), .C2(n14790), .A(n10666), .B(n10665), .ZN(
        n10667) );
  INV_X1 U13762 ( .A(n10667), .ZN(n10668) );
  INV_X1 U13763 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n19412) );
  INV_X1 U13764 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14606) );
  OR2_X1 U13765 ( .A1(n10662), .A2(n14606), .ZN(n10672) );
  AOI22_X1 U13766 ( .A1(n11340), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10671) );
  OAI211_X1 U13767 ( .C1(n10747), .C2(n19412), .A(n10672), .B(n10671), .ZN(
        n14600) );
  NAND2_X1 U13768 ( .A1(n14457), .A2(n14600), .ZN(n13830) );
  INV_X1 U13769 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16708) );
  OR2_X1 U13770 ( .A1(n10662), .A2(n16708), .ZN(n10677) );
  INV_X1 U13771 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n19401) );
  NAND2_X1 U13772 ( .A1(n11340), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10674) );
  NAND2_X1 U13773 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10673) );
  OAI211_X1 U13774 ( .C1(n10747), .C2(n19401), .A(n10674), .B(n10673), .ZN(
        n10675) );
  INV_X1 U13775 ( .A(n10675), .ZN(n10676) );
  INV_X1 U13776 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10816) );
  OR2_X1 U13777 ( .A1(n10662), .A2(n10816), .ZN(n10683) );
  INV_X1 U13778 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n10680) );
  NAND2_X1 U13779 ( .A1(n11340), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10679) );
  NAND2_X1 U13780 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10678) );
  OAI211_X1 U13781 ( .C1(n10747), .C2(n10680), .A(n10679), .B(n10678), .ZN(
        n10681) );
  INV_X1 U13782 ( .A(n10681), .ZN(n10682) );
  NAND2_X1 U13783 ( .A1(n10683), .A2(n10682), .ZN(n13851) );
  INV_X1 U13784 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10826) );
  OR2_X1 U13785 ( .A1(n10662), .A2(n10826), .ZN(n10685) );
  AOI22_X1 U13786 ( .A1(n11340), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10684) );
  OAI211_X1 U13787 ( .C1(n10010), .C2(n10747), .A(n10685), .B(n10684), .ZN(
        n13907) );
  INV_X1 U13788 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10688) );
  INV_X1 U13789 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16694) );
  OR2_X1 U13790 ( .A1(n10662), .A2(n16694), .ZN(n10687) );
  AOI22_X1 U13791 ( .A1(n11340), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10686) );
  OAI211_X1 U13792 ( .C1(n10747), .C2(n10688), .A(n10687), .B(n10686), .ZN(
        n13931) );
  OR2_X1 U13793 ( .A1(n10662), .A2(n16042), .ZN(n10693) );
  INV_X1 U13794 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13948) );
  NAND2_X1 U13795 ( .A1(n11340), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n10690) );
  NAND2_X1 U13796 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10689) );
  OAI211_X1 U13797 ( .C1(n10747), .C2(n13948), .A(n10690), .B(n10689), .ZN(
        n10691) );
  INV_X1 U13798 ( .A(n10691), .ZN(n10692) );
  INV_X1 U13799 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16020) );
  OR2_X1 U13800 ( .A1(n10662), .A2(n16020), .ZN(n10698) );
  INV_X1 U13801 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n19359) );
  NAND2_X1 U13802 ( .A1(n11340), .A2(P2_REIP_REG_12__SCAN_IN), .ZN(n10695) );
  NAND2_X1 U13803 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10694) );
  OAI211_X1 U13804 ( .C1(n10747), .C2(n19359), .A(n10695), .B(n10694), .ZN(
        n10696) );
  INV_X1 U13805 ( .A(n10696), .ZN(n10697) );
  NAND2_X1 U13806 ( .A1(n10698), .A2(n10697), .ZN(n13989) );
  INV_X1 U13807 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10767) );
  INV_X1 U13808 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16605) );
  OR2_X1 U13809 ( .A1(n10662), .A2(n16605), .ZN(n10700) );
  AOI22_X1 U13810 ( .A1(n11340), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n10699) );
  OAI211_X1 U13811 ( .C1(n10767), .C2(n10747), .A(n10700), .B(n10699), .ZN(
        n14070) );
  INV_X1 U13812 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n10768) );
  OR2_X1 U13813 ( .A1(n10662), .A2(n16007), .ZN(n10702) );
  AOI22_X1 U13814 ( .A1(n11340), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n10701) );
  OAI211_X1 U13815 ( .C1(n10768), .C2(n10747), .A(n10702), .B(n10701), .ZN(
        n14300) );
  INV_X1 U13816 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15966) );
  OR2_X1 U13817 ( .A1(n10662), .A2(n15966), .ZN(n10707) );
  INV_X1 U13818 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n19316) );
  NAND2_X1 U13819 ( .A1(n11340), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10704) );
  NAND2_X1 U13820 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10703) );
  OAI211_X1 U13821 ( .C1(n10747), .C2(n19316), .A(n10704), .B(n10703), .ZN(
        n10705) );
  INV_X1 U13822 ( .A(n10705), .ZN(n10706) );
  NAND2_X1 U13823 ( .A1(n10707), .A2(n10706), .ZN(n14330) );
  NAND2_X1 U13824 ( .A1(n10708), .A2(n14330), .ZN(n14331) );
  INV_X1 U13825 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n14424) );
  NAND2_X1 U13826 ( .A1(n11340), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10710) );
  NAND2_X1 U13827 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10709) );
  OAI211_X1 U13828 ( .C1(n10747), .C2(n14424), .A(n10710), .B(n10709), .ZN(
        n10711) );
  AOI21_X1 U13829 ( .B1(n10654), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10711), .ZN(n14422) );
  INV_X1 U13830 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n19293) );
  NAND2_X1 U13831 ( .A1(n11340), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n10713) );
  NAND2_X1 U13832 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10712) );
  OAI211_X1 U13833 ( .C1(n10747), .C2(n19293), .A(n10713), .B(n10712), .ZN(
        n10714) );
  AOI21_X1 U13834 ( .B1(n10654), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10714), .ZN(n14473) );
  INV_X1 U13835 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n19277) );
  INV_X1 U13836 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15953) );
  OR2_X1 U13837 ( .A1(n10662), .A2(n15953), .ZN(n10716) );
  AOI22_X1 U13838 ( .A1(n11340), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10715) );
  OAI211_X1 U13839 ( .C1(n10747), .C2(n19277), .A(n10716), .B(n10715), .ZN(
        n14645) );
  INV_X1 U13840 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10719) );
  NAND2_X1 U13841 ( .A1(n11340), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n10718) );
  NAND2_X1 U13842 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10717) );
  OAI211_X1 U13843 ( .C1(n10747), .C2(n10719), .A(n10718), .B(n10717), .ZN(
        n10720) );
  AOI21_X1 U13844 ( .B1(n10654), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10720), .ZN(n14651) );
  INV_X1 U13845 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n19248) );
  NAND2_X1 U13846 ( .A1(n11340), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n10722) );
  NAND2_X1 U13847 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10721) );
  OAI211_X1 U13848 ( .C1(n10747), .C2(n19248), .A(n10722), .B(n10721), .ZN(
        n10723) );
  AOI21_X1 U13849 ( .B1(n10654), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n10723), .ZN(n15613) );
  INV_X1 U13850 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13224) );
  OR2_X1 U13851 ( .A1(n10662), .A2(n13224), .ZN(n10726) );
  INV_X1 U13852 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n20131) );
  INV_X1 U13853 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n14795) );
  INV_X1 U13854 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14670) );
  OAI22_X1 U13855 ( .A1(n10670), .A2(n20131), .B1(n14795), .B2(n14670), .ZN(
        n10724) );
  AOI21_X1 U13856 ( .B1(n9658), .B2(P2_EBX_REG_21__SCAN_IN), .A(n10724), .ZN(
        n10725) );
  NAND2_X1 U13857 ( .A1(n10726), .A2(n10725), .ZN(n13221) );
  INV_X1 U13858 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n10729) );
  INV_X1 U13859 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15905) );
  OR2_X1 U13860 ( .A1(n10662), .A2(n15905), .ZN(n10728) );
  AOI22_X1 U13861 ( .A1(n11340), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10727) );
  OAI211_X1 U13862 ( .C1(n10747), .C2(n10729), .A(n10728), .B(n10727), .ZN(
        n15603) );
  INV_X1 U13863 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n16558) );
  NAND2_X1 U13864 ( .A1(n11340), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n10731) );
  NAND2_X1 U13865 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10730) );
  OAI211_X1 U13866 ( .C1(n10747), .C2(n16558), .A(n10731), .B(n10730), .ZN(
        n10732) );
  AOI21_X1 U13867 ( .B1(n10654), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n10732), .ZN(n15597) );
  INV_X1 U13868 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10735) );
  NAND2_X1 U13869 ( .A1(n11340), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10734) );
  NAND2_X1 U13870 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10733) );
  OAI211_X1 U13871 ( .C1(n10747), .C2(n10735), .A(n10734), .B(n10733), .ZN(
        n10736) );
  AOI21_X1 U13872 ( .B1(n10654), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10736), .ZN(n15588) );
  INV_X1 U13873 ( .A(n15588), .ZN(n10737) );
  INV_X1 U13874 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n16531) );
  NAND2_X1 U13875 ( .A1(n11340), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n10739) );
  NAND2_X1 U13876 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10738) );
  OAI211_X1 U13877 ( .C1(n10747), .C2(n16531), .A(n10739), .B(n10738), .ZN(
        n10740) );
  AOI21_X1 U13878 ( .B1(n10654), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n10740), .ZN(n15581) );
  INV_X1 U13879 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n16518) );
  INV_X1 U13880 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15872) );
  OR2_X1 U13881 ( .A1(n10662), .A2(n15872), .ZN(n10742) );
  AOI22_X1 U13882 ( .A1(n11340), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n10741) );
  OAI211_X1 U13883 ( .C1(n10747), .C2(n16518), .A(n10742), .B(n10741), .ZN(
        n15571) );
  INV_X1 U13884 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n16502) );
  INV_X1 U13885 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15730) );
  OR2_X1 U13886 ( .A1(n10662), .A2(n15730), .ZN(n10744) );
  AOI22_X1 U13887 ( .A1(n11340), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n10743) );
  OAI211_X1 U13888 ( .C1(n10747), .C2(n16502), .A(n10744), .B(n10743), .ZN(
        n15562) );
  INV_X1 U13889 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n10774) );
  INV_X1 U13890 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11637) );
  OR2_X1 U13891 ( .A1(n10662), .A2(n11637), .ZN(n10746) );
  AOI22_X1 U13892 ( .A1(n11340), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n10745) );
  OAI211_X1 U13893 ( .C1(n10747), .C2(n10774), .A(n10746), .B(n10745), .ZN(
        n15509) );
  NAND2_X1 U13894 ( .A1(n14795), .A2(n20195), .ZN(n20165) );
  NAND2_X1 U13895 ( .A1(n20016), .A2(n20165), .ZN(n20194) );
  NAND2_X1 U13896 ( .A1(n20194), .A2(n20218), .ZN(n10750) );
  AND2_X1 U13897 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n20184) );
  INV_X1 U13898 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10756) );
  INV_X1 U13899 ( .A(n12809), .ZN(n10752) );
  NAND2_X1 U13900 ( .A1(n20226), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10751) );
  NAND2_X1 U13901 ( .A1(n10752), .A2(n10751), .ZN(n13460) );
  INV_X1 U13902 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16665) );
  NAND2_X1 U13903 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n14180), .ZN(
        n14179) );
  NOR2_X2 U13904 ( .A1(n16665), .A2(n14179), .ZN(n14182) );
  INV_X1 U13905 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15794) );
  INV_X1 U13906 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16533) );
  INV_X1 U13907 ( .A(n14678), .ZN(n10753) );
  AOI21_X1 U13908 ( .B1(n10756), .B2(n15533), .A(n10753), .ZN(n16470) );
  NAND2_X1 U13909 ( .A1(n16667), .A2(n16470), .ZN(n10755) );
  NOR2_X1 U13910 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n20165), .ZN(n10754) );
  NAND2_X1 U13911 ( .A1(n10754), .A2(n19942), .ZN(n19341) );
  NAND2_X1 U13912 ( .A1(n19500), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15840) );
  OAI211_X1 U13913 ( .C1(n16677), .C2(n10756), .A(n10755), .B(n15840), .ZN(
        n10757) );
  MUX2_X1 U13914 ( .A(n10759), .B(n10287), .S(n19551), .Z(n10792) );
  NOR2_X1 U13915 ( .A1(n14815), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10785) );
  INV_X1 U13916 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14320) );
  NAND2_X1 U13917 ( .A1(n10785), .A2(n14320), .ZN(n10761) );
  INV_X1 U13918 ( .A(n11402), .ZN(n10760) );
  NAND2_X1 U13919 ( .A1(n10761), .A2(n10093), .ZN(n10791) );
  NAND2_X1 U13920 ( .A1(n10792), .A2(n10791), .ZN(n10790) );
  MUX2_X1 U13921 ( .A(n10765), .B(n14222), .S(n19551), .Z(n10798) );
  MUX2_X1 U13922 ( .A(n14790), .B(n11426), .S(n14815), .Z(n10779) );
  MUX2_X1 U13923 ( .A(n11429), .B(P2_EBX_REG_6__SCAN_IN), .S(n19551), .Z(
        n10807) );
  NOR2_X2 U13924 ( .A1(n10778), .A2(n10807), .ZN(n10813) );
  MUX2_X1 U13925 ( .A(n19401), .B(n14818), .S(n14815), .Z(n10812) );
  NAND2_X1 U13926 ( .A1(n19551), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10810) );
  NAND2_X1 U13927 ( .A1(n19366), .A2(n13948), .ZN(n10830) );
  NAND2_X1 U13928 ( .A1(n19551), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10831) );
  NOR2_X1 U13929 ( .A1(n14815), .A2(n10767), .ZN(n10854) );
  NOR2_X1 U13930 ( .A1(n14815), .A2(n10768), .ZN(n10849) );
  NAND2_X1 U13931 ( .A1(n19551), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10846) );
  NOR2_X1 U13932 ( .A1(n14815), .A2(n14424), .ZN(n10769) );
  NOR2_X1 U13933 ( .A1(n14815), .A2(n19293), .ZN(n10841) );
  NOR2_X1 U13934 ( .A1(n14815), .A2(n19277), .ZN(n10861) );
  NAND2_X1 U13935 ( .A1(n19551), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10858) );
  NAND2_X1 U13936 ( .A1(n19551), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10888) );
  NAND2_X1 U13937 ( .A1(n10838), .A2(n10888), .ZN(n10887) );
  NOR2_X1 U13938 ( .A1(n14815), .A2(n16558), .ZN(n10895) );
  OR2_X2 U13939 ( .A1(n10887), .A2(n10895), .ZN(n10898) );
  INV_X1 U13940 ( .A(n10906), .ZN(n10772) );
  NOR2_X1 U13941 ( .A1(n10915), .A2(n10772), .ZN(n14816) );
  INV_X1 U13942 ( .A(n14816), .ZN(n10773) );
  NAND2_X1 U13943 ( .A1(n19551), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10914) );
  NOR2_X1 U13944 ( .A1(n14815), .A2(n10774), .ZN(n10911) );
  OR2_X2 U13945 ( .A1(n10919), .A2(n10911), .ZN(n11282) );
  INV_X1 U13946 ( .A(n11282), .ZN(n10775) );
  NAND2_X1 U13947 ( .A1(n19551), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n11280) );
  XNOR2_X1 U13948 ( .A(n10775), .B(n11280), .ZN(n10776) );
  INV_X1 U13949 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15843) );
  OAI21_X1 U13950 ( .B1(n10776), .B2(n10781), .A(n15843), .ZN(n11278) );
  INV_X1 U13951 ( .A(n10776), .ZN(n16492) );
  NAND3_X1 U13952 ( .A1(n16492), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14818), .ZN(n14809) );
  NAND2_X1 U13953 ( .A1(n10777), .A2(n10781), .ZN(n10780) );
  INV_X1 U13954 ( .A(n14818), .ZN(n10781) );
  INV_X1 U13955 ( .A(n10782), .ZN(n10799) );
  NAND2_X1 U13956 ( .A1(n10790), .A2(n10783), .ZN(n10784) );
  NAND2_X1 U13957 ( .A1(n10799), .A2(n10784), .ZN(n14288) );
  MUX2_X1 U13958 ( .A(n11395), .B(n11295), .S(n11336), .Z(n10786) );
  AOI21_X1 U13959 ( .B1(n10786), .B2(n14815), .A(n10785), .ZN(n14341) );
  NAND2_X1 U13960 ( .A1(n14341), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13474) );
  NAND2_X1 U13961 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), 
        .ZN(n10787) );
  NOR2_X1 U13962 ( .A1(n14815), .A2(n10787), .ZN(n10788) );
  OR2_X1 U13963 ( .A1(n10791), .A2(n10788), .ZN(n14318) );
  NOR2_X1 U13964 ( .A1(n13474), .A2(n14318), .ZN(n10789) );
  NAND2_X1 U13965 ( .A1(n13474), .A2(n14318), .ZN(n13473) );
  OAI21_X1 U13966 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10789), .A(
        n13473), .ZN(n14761) );
  OAI21_X1 U13967 ( .B1(n10792), .B2(n10791), .A(n10790), .ZN(n14743) );
  XNOR2_X1 U13968 ( .A(n14743), .B(n10290), .ZN(n14760) );
  OR2_X1 U13969 ( .A1(n14761), .A2(n14760), .ZN(n14778) );
  INV_X1 U13970 ( .A(n14743), .ZN(n10793) );
  NAND2_X1 U13971 ( .A1(n10793), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10794) );
  AND2_X1 U13972 ( .A1(n14778), .A2(n10794), .ZN(n14370) );
  NAND2_X1 U13973 ( .A1(n14368), .A2(n14370), .ZN(n10797) );
  NAND2_X1 U13974 ( .A1(n10797), .A2(n14369), .ZN(n16078) );
  NAND2_X1 U13975 ( .A1(n10799), .A2(n10000), .ZN(n10800) );
  NAND2_X1 U13976 ( .A1(n10801), .A2(n10800), .ZN(n14226) );
  XNOR2_X1 U13977 ( .A(n14226), .B(n10595), .ZN(n16079) );
  INV_X1 U13978 ( .A(n14226), .ZN(n10802) );
  NAND2_X1 U13979 ( .A1(n10802), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10803) );
  OAI21_X2 U13980 ( .B1(n16078), .B2(n16079), .A(n10803), .ZN(n14443) );
  NAND2_X1 U13981 ( .A1(n14442), .A2(n14443), .ZN(n10806) );
  NAND2_X1 U13982 ( .A1(n10804), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10805) );
  XNOR2_X1 U13983 ( .A(n10778), .B(n10807), .ZN(n19414) );
  XNOR2_X1 U13984 ( .A(n10809), .B(n14606), .ZN(n14593) );
  NAND2_X1 U13985 ( .A1(n10809), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15828) );
  OR2_X1 U13986 ( .A1(n10766), .A2(n10810), .ZN(n10811) );
  NAND2_X1 U13987 ( .A1(n10820), .A2(n10811), .ZN(n14214) );
  NOR2_X1 U13988 ( .A1(n14214), .A2(n10781), .ZN(n10815) );
  NAND2_X1 U13989 ( .A1(n10815), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16650) );
  NOR2_X1 U13990 ( .A1(n10813), .A2(n10812), .ZN(n10814) );
  OR2_X1 U13991 ( .A1(n10766), .A2(n10814), .ZN(n10818) );
  INV_X1 U13992 ( .A(n10818), .ZN(n19404) );
  NAND2_X1 U13993 ( .A1(n19404), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16647) );
  AND2_X1 U13994 ( .A1(n16650), .A2(n16647), .ZN(n16062) );
  AND2_X1 U13995 ( .A1(n15828), .A2(n16062), .ZN(n10822) );
  INV_X1 U13996 ( .A(n10815), .ZN(n10817) );
  NAND2_X1 U13997 ( .A1(n10817), .A2(n10816), .ZN(n16649) );
  NAND2_X1 U13998 ( .A1(n10818), .A2(n16708), .ZN(n16645) );
  AND2_X1 U13999 ( .A1(n16649), .A2(n16645), .ZN(n16063) );
  NAND2_X1 U14000 ( .A1(n19551), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10819) );
  XNOR2_X1 U14001 ( .A(n10820), .B(n10819), .ZN(n19379) );
  NAND2_X1 U14002 ( .A1(n19379), .A2(n14818), .ZN(n10827) );
  NAND2_X1 U14003 ( .A1(n10827), .A2(n10826), .ZN(n16065) );
  NAND2_X1 U14004 ( .A1(n16063), .A2(n16065), .ZN(n10821) );
  NAND3_X1 U14005 ( .A1(n10824), .A2(n19551), .A3(P2_EBX_REG_10__SCAN_IN), 
        .ZN(n10823) );
  OAI211_X1 U14006 ( .C1(n10824), .C2(P2_EBX_REG_10__SCAN_IN), .A(n10906), .B(
        n10823), .ZN(n14203) );
  OAI21_X1 U14007 ( .B1(n14203), .B2(n10781), .A(n16694), .ZN(n16624) );
  NAND2_X1 U14008 ( .A1(n14818), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10825) );
  OR2_X1 U14009 ( .A1(n14203), .A2(n10825), .ZN(n16623) );
  OR2_X1 U14010 ( .A1(n10827), .A2(n10826), .ZN(n16621) );
  AND2_X1 U14011 ( .A1(n16623), .A2(n16621), .ZN(n10828) );
  INV_X1 U14012 ( .A(n16037), .ZN(n10829) );
  INV_X1 U14013 ( .A(n10830), .ZN(n10832) );
  OR2_X1 U14014 ( .A1(n10832), .A2(n10831), .ZN(n10834) );
  AND2_X1 U14015 ( .A1(n10834), .A2(n10833), .ZN(n19356) );
  NAND2_X1 U14016 ( .A1(n19356), .A2(n14818), .ZN(n10857) );
  INV_X1 U14017 ( .A(n10857), .ZN(n10835) );
  AND3_X1 U14018 ( .A1(n10836), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n19551), .ZN(
        n10837) );
  OR2_X1 U14019 ( .A1(n10838), .A2(n10837), .ZN(n10870) );
  NAND3_X1 U14020 ( .A1(n10839), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n19551), 
        .ZN(n10840) );
  OAI211_X1 U14021 ( .C1(n10839), .C2(P2_EBX_REG_16__SCAN_IN), .A(n10840), .B(
        n10906), .ZN(n19304) );
  OR2_X1 U14022 ( .A1(n19304), .A2(n10781), .ZN(n10880) );
  XNOR2_X1 U14023 ( .A(n10880), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13207) );
  NAND2_X1 U14024 ( .A1(n10842), .A2(n10841), .ZN(n10843) );
  AND2_X1 U14025 ( .A1(n10862), .A2(n10843), .ZN(n19295) );
  NAND2_X1 U14026 ( .A1(n19295), .A2(n14818), .ZN(n10845) );
  INV_X1 U14027 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10844) );
  NAND2_X1 U14028 ( .A1(n10845), .A2(n10844), .ZN(n13210) );
  INV_X1 U14029 ( .A(n10846), .ZN(n10847) );
  XNOR2_X1 U14030 ( .A(n10852), .B(n10847), .ZN(n19318) );
  NAND2_X1 U14031 ( .A1(n19318), .A2(n14818), .ZN(n10848) );
  NAND2_X1 U14032 ( .A1(n10848), .A2(n15966), .ZN(n15988) );
  AND2_X1 U14033 ( .A1(n10850), .A2(n10849), .ZN(n10851) );
  OR2_X1 U14034 ( .A1(n10852), .A2(n10851), .ZN(n19329) );
  INV_X1 U14035 ( .A(n19329), .ZN(n10853) );
  NAND2_X1 U14036 ( .A1(n10853), .A2(n14818), .ZN(n10877) );
  INV_X1 U14037 ( .A(n10854), .ZN(n10855) );
  XNOR2_X1 U14038 ( .A(n10833), .B(n10855), .ZN(n19339) );
  NAND2_X1 U14039 ( .A1(n19339), .A2(n14818), .ZN(n10856) );
  NAND2_X1 U14040 ( .A1(n10856), .A2(n16605), .ZN(n13203) );
  NAND2_X1 U14041 ( .A1(n10857), .A2(n16020), .ZN(n16023) );
  NAND4_X1 U14042 ( .A1(n13215), .A2(n13207), .A3(n9755), .A4(n16023), .ZN(
        n10867) );
  NOR2_X1 U14043 ( .A1(n10863), .A2(n10858), .ZN(n10859) );
  OR2_X1 U14044 ( .A1(n10866), .A2(n10859), .ZN(n19264) );
  INV_X1 U14045 ( .A(n19264), .ZN(n10860) );
  NAND2_X1 U14046 ( .A1(n10860), .A2(n14818), .ZN(n10872) );
  INV_X1 U14047 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15929) );
  NAND2_X1 U14048 ( .A1(n10872), .A2(n15929), .ZN(n15790) );
  AND2_X1 U14049 ( .A1(n10862), .A2(n10861), .ZN(n10864) );
  OR2_X1 U14050 ( .A1(n10864), .A2(n10863), .ZN(n19280) );
  OAI21_X1 U14051 ( .B1(n19280), .B2(n10781), .A(n15953), .ZN(n15800) );
  NAND2_X1 U14052 ( .A1(n15790), .A2(n15800), .ZN(n15775) );
  NOR2_X1 U14053 ( .A1(n14815), .A2(n19248), .ZN(n10865) );
  XNOR2_X1 U14054 ( .A(n10866), .B(n10865), .ZN(n19246) );
  NAND2_X1 U14055 ( .A1(n19246), .A2(n14818), .ZN(n10883) );
  INV_X1 U14056 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15932) );
  AND2_X1 U14057 ( .A1(n10883), .A2(n15932), .ZN(n15778) );
  OR2_X1 U14058 ( .A1(n15775), .A2(n15778), .ZN(n13213) );
  NOR2_X1 U14059 ( .A1(n10867), .A2(n13213), .ZN(n10869) );
  OR2_X1 U14060 ( .A1(n19367), .A2(n10781), .ZN(n16038) );
  NAND2_X1 U14061 ( .A1(n10868), .A2(n16038), .ZN(n13199) );
  OAI211_X1 U14062 ( .C1(n13198), .C2(n16024), .A(n10869), .B(n13199), .ZN(
        n10886) );
  INV_X1 U14063 ( .A(n10870), .ZN(n19241) );
  AND2_X1 U14064 ( .A1(n14818), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10871) );
  NAND2_X1 U14065 ( .A1(n19241), .A2(n10871), .ZN(n13214) );
  INV_X1 U14066 ( .A(n10872), .ZN(n10873) );
  NAND2_X1 U14067 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15791) );
  NAND2_X1 U14068 ( .A1(n14818), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10874) );
  NOR2_X1 U14069 ( .A1(n19280), .A2(n10874), .ZN(n13211) );
  AND2_X1 U14070 ( .A1(n14818), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10875) );
  NAND2_X1 U14071 ( .A1(n19295), .A2(n10875), .ZN(n13209) );
  INV_X1 U14072 ( .A(n19339), .ZN(n10876) );
  OR3_X1 U14073 ( .A1(n10876), .A2(n10781), .A3(n16605), .ZN(n13202) );
  INV_X1 U14074 ( .A(n10877), .ZN(n10878) );
  NAND2_X1 U14075 ( .A1(n10878), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16016) );
  NAND3_X1 U14076 ( .A1(n13209), .A2(n13202), .A3(n16016), .ZN(n10879) );
  NOR2_X1 U14077 ( .A1(n13211), .A2(n10879), .ZN(n10882) );
  INV_X1 U14078 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15985) );
  OR2_X1 U14079 ( .A1(n10880), .A2(n15985), .ZN(n13208) );
  INV_X1 U14080 ( .A(n19318), .ZN(n10881) );
  AND4_X1 U14081 ( .A1(n15791), .A2(n10882), .A3(n13208), .A4(n15987), .ZN(
        n10884) );
  AND3_X1 U14082 ( .A1(n13214), .A2(n10884), .A3(n15777), .ZN(n10885) );
  NAND2_X1 U14083 ( .A1(n10886), .A2(n10885), .ZN(n15915) );
  INV_X1 U14084 ( .A(n10888), .ZN(n10889) );
  NAND2_X1 U14085 ( .A1(n10890), .A2(n10889), .ZN(n10891) );
  NAND2_X1 U14086 ( .A1(n10887), .A2(n10891), .ZN(n16207) );
  OR2_X1 U14087 ( .A1(n16207), .A2(n10781), .ZN(n10892) );
  NAND2_X1 U14088 ( .A1(n10892), .A2(n15905), .ZN(n15916) );
  NAND2_X1 U14089 ( .A1(n15915), .A2(n15916), .ZN(n10894) );
  INV_X1 U14090 ( .A(n10892), .ZN(n10893) );
  NAND2_X1 U14091 ( .A1(n10893), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15917) );
  INV_X1 U14092 ( .A(n10895), .ZN(n10896) );
  XNOR2_X1 U14093 ( .A(n10887), .B(n10896), .ZN(n16560) );
  NAND2_X1 U14094 ( .A1(n16560), .A2(n14818), .ZN(n10897) );
  XNOR2_X1 U14095 ( .A(n10897), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15771) );
  NAND3_X1 U14096 ( .A1(n10898), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n19551), 
        .ZN(n10899) );
  NAND2_X1 U14097 ( .A1(n10899), .A2(n10906), .ZN(n10900) );
  OR2_X1 U14098 ( .A1(n10900), .A2(n10904), .ZN(n16545) );
  NOR2_X1 U14099 ( .A1(n16545), .A2(n10781), .ZN(n10901) );
  AND2_X1 U14100 ( .A1(n10901), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15759) );
  INV_X1 U14101 ( .A(n10901), .ZN(n10902) );
  NAND2_X1 U14102 ( .A1(n10902), .A2(n15895), .ZN(n15760) );
  INV_X1 U14103 ( .A(n15734), .ZN(n10910) );
  NAND3_X1 U14104 ( .A1(n19551), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n10907), 
        .ZN(n10903) );
  NOR2_X1 U14105 ( .A1(n10904), .A2(n16531), .ZN(n10905) );
  NAND2_X1 U14106 ( .A1(n10919), .A2(n10911), .ZN(n10912) );
  NAND2_X1 U14107 ( .A1(n11282), .A2(n10912), .ZN(n15535) );
  INV_X1 U14108 ( .A(n10914), .ZN(n10917) );
  INV_X1 U14109 ( .A(n10915), .ZN(n10916) );
  NAND2_X1 U14110 ( .A1(n10917), .A2(n10916), .ZN(n10918) );
  NAND2_X1 U14111 ( .A1(n10919), .A2(n10918), .ZN(n16505) );
  NOR2_X2 U14112 ( .A1(n15712), .A2(n15710), .ZN(n15707) );
  INV_X1 U14113 ( .A(n10920), .ZN(n10921) );
  NAND2_X1 U14114 ( .A1(n10921), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10922) );
  INV_X1 U14115 ( .A(n15846), .ZN(n10924) );
  INV_X1 U14116 ( .A(n16671), .ZN(n10923) );
  NAND2_X1 U14117 ( .A1(n10924), .A2(n10923), .ZN(n10925) );
  NOR2_X2 U14118 ( .A1(n10934), .A2(n10927), .ZN(n17470) );
  NAND3_X1 U14119 ( .A1(n9997), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10933) );
  AOI22_X1 U14120 ( .A1(n16175), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10944) );
  NAND3_X1 U14121 ( .A1(n9715), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n18984), .ZN(n16111) );
  NOR3_X1 U14122 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n9716), .ZN(n10926) );
  NAND2_X2 U14123 ( .A1(n10926), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10978) );
  INV_X1 U14124 ( .A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10930) );
  INV_X4 U14125 ( .A(n11128), .ZN(n17456) );
  AOI22_X1 U14126 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10929) );
  NOR2_X2 U14127 ( .A1(n10927), .A2(n10931), .ZN(n11030) );
  INV_X2 U14128 ( .A(n11030), .ZN(n17256) );
  AOI22_X1 U14129 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17508), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10928) );
  OAI211_X1 U14130 ( .C1(n10978), .C2(n10930), .A(n10929), .B(n10928), .ZN(
        n10942) );
  AOI22_X1 U14131 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9670), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U14132 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17494), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U14133 ( .A1(n10981), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10938) );
  NAND2_X1 U14134 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10937) );
  NAND4_X1 U14135 ( .A1(n10940), .A2(n10939), .A3(n10938), .A4(n10937), .ZN(
        n10941) );
  AOI211_X1 U14136 ( .C1(n17512), .C2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n10942), .B(n10941), .ZN(n10943) );
  OAI211_X1 U14137 ( .C1(n10109), .C2(n17418), .A(n10944), .B(n10943), .ZN(
        n10945) );
  AOI22_X1 U14138 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10947) );
  OAI21_X1 U14139 ( .B1(n9672), .B2(n17540), .A(n10947), .ZN(n10958) );
  INV_X1 U14140 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17436) );
  AOI22_X1 U14141 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10956) );
  INV_X2 U14142 ( .A(n17472), .ZN(n10981) );
  INV_X1 U14143 ( .A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17332) );
  INV_X1 U14144 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16152) );
  OAI22_X1 U14145 ( .A1(n10949), .A2(n17332), .B1(n10978), .B2(n16152), .ZN(
        n10954) );
  INV_X2 U14146 ( .A(n10970), .ZN(n17520) );
  AOI22_X1 U14147 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10952) );
  AOI22_X1 U14148 ( .A1(n11030), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17494), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10951) );
  AOI22_X1 U14149 ( .A1(n17512), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10950) );
  NAND3_X1 U14150 ( .A1(n10952), .A2(n10951), .A3(n10950), .ZN(n10953) );
  AOI211_X1 U14151 ( .C1(n17339), .C2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A(
        n10954), .B(n10953), .ZN(n10955) );
  OAI211_X1 U14152 ( .C1(n17474), .C2(n17436), .A(n10956), .B(n10955), .ZN(
        n10957) );
  INV_X1 U14153 ( .A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17372) );
  AOI22_X1 U14154 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9671), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U14155 ( .A1(n11156), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10959) );
  OAI211_X1 U14156 ( .C1(n10978), .C2(n17372), .A(n10960), .B(n10959), .ZN(
        n10966) );
  AOI22_X1 U14157 ( .A1(n10981), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n10961), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10962) );
  OAI21_X1 U14158 ( .B1(n17455), .B2(n18579), .A(n10962), .ZN(n10964) );
  AOI22_X1 U14159 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17403), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10967) );
  AOI22_X1 U14160 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17494), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10971) );
  OAI21_X1 U14161 ( .B1(n17256), .B2(n18749), .A(n10971), .ZN(n10973) );
  AOI22_X1 U14162 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10980) );
  AOI22_X1 U14163 ( .A1(n17512), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17514), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10979) );
  INV_X1 U14164 ( .A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17355) );
  INV_X1 U14165 ( .A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n18582) );
  OAI22_X1 U14166 ( .A1(n11006), .A2(n17355), .B1(n17455), .B2(n18582), .ZN(
        n10983) );
  AND2_X1 U14167 ( .A1(n10981), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10982) );
  INV_X1 U14168 ( .A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U14169 ( .A1(n11030), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10987) );
  AOI22_X1 U14170 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9670), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10986) );
  NAND4_X1 U14171 ( .A1(n10104), .A2(n10988), .A3(n10987), .A4(n10986), .ZN(
        n10993) );
  AOI22_X1 U14172 ( .A1(n10961), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10989) );
  OAI21_X1 U14173 ( .B1(n10109), .B2(n17471), .A(n10989), .ZN(n10991) );
  NOR2_X2 U14174 ( .A1(n10993), .A2(n10992), .ZN(n17712) );
  AOI22_X1 U14175 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11003) );
  INV_X1 U14176 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n16099) );
  AOI22_X1 U14177 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10961), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10995) );
  AOI22_X1 U14178 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10994) );
  OAI211_X1 U14179 ( .C1(n10978), .C2(n16099), .A(n10995), .B(n10994), .ZN(
        n11001) );
  AOI22_X1 U14180 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17494), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U14181 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11030), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U14182 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10981), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10997) );
  NAND2_X1 U14183 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10996) );
  NAND4_X1 U14184 ( .A1(n10999), .A2(n10998), .A3(n10997), .A4(n10996), .ZN(
        n11000) );
  AOI211_X1 U14185 ( .C1(n17512), .C2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A(
        n11001), .B(n11000), .ZN(n11002) );
  NAND2_X1 U14186 ( .A1(n11040), .A2(n11205), .ZN(n11044) );
  AOI22_X1 U14187 ( .A1(n10981), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10961), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11014) );
  INV_X1 U14188 ( .A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n18589) );
  AOI22_X1 U14189 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U14190 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17495), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11004) );
  OAI211_X1 U14191 ( .C1(n17455), .C2(n18589), .A(n11005), .B(n11004), .ZN(
        n11012) );
  AOI22_X1 U14192 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11030), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11010) );
  AOI22_X1 U14193 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11009) );
  INV_X4 U14194 ( .A(n11006), .ZN(n17494) );
  AOI22_X1 U14195 ( .A1(n17494), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11008) );
  NAND2_X1 U14196 ( .A1(n17514), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11007) );
  NAND4_X1 U14197 ( .A1(n11010), .A2(n11009), .A3(n11008), .A4(n11007), .ZN(
        n11011) );
  OAI211_X1 U14198 ( .C1(n9672), .C2(n17537), .A(n11014), .B(n11013), .ZN(
        n11203) );
  INV_X1 U14199 ( .A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17248) );
  AOI22_X1 U14200 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n16175), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11015) );
  OAI21_X1 U14201 ( .B1(n10949), .B2(n17248), .A(n11015), .ZN(n11025) );
  INV_X1 U14202 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11023) );
  AOI22_X1 U14203 ( .A1(n17512), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17494), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11022) );
  INV_X1 U14204 ( .A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17402) );
  AOI22_X1 U14205 ( .A1(n10981), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17508), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11016) );
  OAI21_X1 U14206 ( .B1(n10970), .B2(n17402), .A(n11016), .ZN(n11020) );
  INV_X1 U14207 ( .A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17247) );
  AOI22_X1 U14208 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9671), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11018) );
  AOI22_X1 U14209 ( .A1(n17476), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11017) );
  OAI211_X1 U14210 ( .C1(n10978), .C2(n17247), .A(n11018), .B(n11017), .ZN(
        n11019) );
  AOI211_X1 U14211 ( .C1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .C2(n11129), .A(
        n11020), .B(n11019), .ZN(n11021) );
  OAI211_X1 U14212 ( .C1(n17474), .C2(n11023), .A(n11022), .B(n11021), .ZN(
        n11024) );
  INV_X1 U14213 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17958) );
  NAND2_X1 U14214 ( .A1(n18080), .A2(n17958), .ZN(n17957) );
  NOR2_X1 U14215 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17957), .ZN(
        n11026) );
  INV_X1 U14216 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17928) );
  NAND2_X1 U14217 ( .A1(n11026), .A2(n17928), .ZN(n17922) );
  INV_X1 U14218 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n18239) );
  INV_X1 U14219 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n18223) );
  NAND3_X1 U14220 ( .A1(n17900), .A2(n18239), .A3(n18223), .ZN(n11066) );
  AOI22_X1 U14221 ( .A1(n10981), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11038) );
  INV_X1 U14222 ( .A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n18576) );
  AOI22_X1 U14223 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10961), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U14224 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9670), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11028) );
  OAI211_X1 U14225 ( .C1(n17455), .C2(n18576), .A(n11029), .B(n11028), .ZN(
        n11036) );
  AOI22_X1 U14226 ( .A1(n11030), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11034) );
  AOI22_X1 U14227 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17495), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11033) );
  AOI22_X1 U14228 ( .A1(n17494), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17403), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11032) );
  NAND2_X1 U14229 ( .A1(n17514), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11031) );
  NAND4_X1 U14230 ( .A1(n11034), .A2(n11033), .A3(n11032), .A4(n11031), .ZN(
        n11035) );
  AOI211_X1 U14231 ( .C1(n17512), .C2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A(
        n11036), .B(n11035), .ZN(n11037) );
  NAND2_X1 U14232 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18175), .ZN(
        n18174) );
  INV_X1 U14233 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n19145) );
  XNOR2_X1 U14234 ( .A(n19145), .B(n17717), .ZN(n18167) );
  XNOR2_X1 U14235 ( .A(n11040), .B(n11205), .ZN(n11041) );
  NOR2_X1 U14236 ( .A1(n11042), .A2(n11041), .ZN(n11043) );
  INV_X1 U14237 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18465) );
  XNOR2_X1 U14238 ( .A(n11042), .B(n11041), .ZN(n18143) );
  NOR2_X1 U14239 ( .A1(n18465), .A2(n18143), .ZN(n18142) );
  XNOR2_X1 U14240 ( .A(n11044), .B(n17704), .ZN(n11045) );
  INV_X1 U14241 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18450) );
  NOR2_X1 U14242 ( .A1(n11046), .A2(n11045), .ZN(n11047) );
  XNOR2_X1 U14243 ( .A(n11048), .B(n11203), .ZN(n18123) );
  XOR2_X1 U14244 ( .A(n11049), .B(n17697), .Z(n11050) );
  XOR2_X1 U14245 ( .A(n18433), .B(n11050), .Z(n18110) );
  NOR2_X1 U14246 ( .A1(n18111), .A2(n18110), .ZN(n18109) );
  OAI21_X1 U14247 ( .B1(n11715), .B2(n17692), .A(n18080), .ZN(n11052) );
  INV_X1 U14248 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18423) );
  NAND2_X1 U14249 ( .A1(n11058), .A2(n11054), .ZN(n11255) );
  INV_X1 U14250 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18052) );
  INV_X1 U14251 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18362) );
  INV_X1 U14252 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18328) );
  NAND2_X1 U14253 ( .A1(n18014), .A2(n10101), .ZN(n11057) );
  NAND2_X1 U14254 ( .A1(n11057), .A2(n18080), .ZN(n11064) );
  INV_X1 U14255 ( .A(n11064), .ZN(n11060) );
  AOI21_X2 U14256 ( .B1(n11058), .B2(n11059), .A(n18278), .ZN(n18029) );
  NOR2_X1 U14257 ( .A1(n18392), .A2(n18378), .ZN(n18376) );
  NAND2_X1 U14258 ( .A1(n18376), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18363) );
  INV_X1 U14259 ( .A(n18363), .ZN(n18351) );
  NAND2_X1 U14260 ( .A1(n18351), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18352) );
  INV_X1 U14261 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18333) );
  NOR2_X1 U14262 ( .A1(n18352), .A2(n18333), .ZN(n18335) );
  NAND2_X1 U14263 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18335), .ZN(
        n18304) );
  INV_X1 U14264 ( .A(n18304), .ZN(n18314) );
  NAND2_X1 U14265 ( .A1(n18314), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11665) );
  NAND2_X1 U14266 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11261) );
  NAND2_X1 U14267 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17923) );
  INV_X1 U14268 ( .A(n17923), .ZN(n18259) );
  NAND3_X1 U14269 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n18259), .ZN(n11260) );
  OR2_X1 U14270 ( .A1(n11260), .A2(n18239), .ZN(n11258) );
  NOR2_X1 U14271 ( .A1(n11261), .A2(n11258), .ZN(n18218) );
  INV_X1 U14272 ( .A(n18218), .ZN(n18230) );
  NOR2_X1 U14273 ( .A1(n18230), .A2(n18223), .ZN(n17868) );
  INV_X1 U14274 ( .A(n17868), .ZN(n17878) );
  INV_X1 U14275 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18310) );
  OAI22_X1 U14276 ( .A1(n11061), .A2(n18310), .B1(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18080), .ZN(n11062) );
  INV_X1 U14277 ( .A(n11062), .ZN(n11063) );
  NAND2_X1 U14278 ( .A1(n11064), .A2(n11063), .ZN(n17965) );
  AOI21_X2 U14279 ( .B1(n11066), .B2(n11065), .A(n17935), .ZN(n17877) );
  INV_X1 U14280 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17881) );
  NOR2_X1 U14281 ( .A1(n9675), .A2(n11261), .ZN(n17920) );
  INV_X1 U14282 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11067) );
  NOR2_X1 U14283 ( .A1(n11068), .A2(n18066), .ZN(n17863) );
  AOI21_X2 U14284 ( .B1(n11069), .B2(n10100), .A(n17863), .ZN(n17848) );
  INV_X1 U14285 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n18186) );
  INV_X1 U14286 ( .A(n11069), .ZN(n11070) );
  NAND2_X2 U14287 ( .A1(n17847), .A2(n9753), .ZN(n11725) );
  INV_X1 U14288 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n18196) );
  INV_X1 U14289 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16200) );
  AOI22_X1 U14290 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n18066), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n11072), .ZN(n11077) );
  INV_X1 U14291 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19146) );
  NOR2_X1 U14292 ( .A1(n19146), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11071) );
  INV_X1 U14293 ( .A(n11071), .ZN(n11270) );
  INV_X1 U14294 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11726) );
  NOR2_X2 U14295 ( .A1(n11687), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11073) );
  INV_X1 U14296 ( .A(n11073), .ZN(n16255) );
  AOI221_X1 U14297 ( .B1(n18066), .B2(n19146), .C1(n18080), .C2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(n11071), .ZN(n11075) );
  INV_X1 U14298 ( .A(n11072), .ZN(n16256) );
  NAND2_X1 U14299 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n19146), .ZN(
        n11264) );
  OAI211_X1 U14300 ( .C1(n18066), .C2(n11073), .A(n16256), .B(n11264), .ZN(
        n11074) );
  AOI22_X1 U14301 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11079) );
  AOI22_X1 U14302 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9670), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11078) );
  OAI211_X1 U14303 ( .C1(n10978), .C2(n18749), .A(n11079), .B(n11078), .ZN(
        n11085) );
  AOI22_X1 U14304 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11083) );
  AOI22_X1 U14305 ( .A1(n16175), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17494), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11082) );
  AOI22_X1 U14306 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17508), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11081) );
  NAND2_X1 U14307 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11080) );
  NAND4_X1 U14308 ( .A1(n11083), .A2(n11082), .A3(n11081), .A4(n11080), .ZN(
        n11084) );
  INV_X1 U14309 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17358) );
  INV_X2 U14310 ( .A(n16118), .ZN(n17490) );
  AOI22_X1 U14311 ( .A1(n16175), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11088) );
  OAI21_X1 U14312 ( .B1(n10949), .B2(n17358), .A(n11088), .ZN(n11097) );
  AOI22_X1 U14313 ( .A1(n17403), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11095) );
  INV_X1 U14314 ( .A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17473) );
  AOI22_X1 U14315 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10981), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11089) );
  OAI21_X1 U14316 ( .B1(n9672), .B2(n17473), .A(n11089), .ZN(n11093) );
  INV_X1 U14317 ( .A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n18752) );
  AOI22_X1 U14318 ( .A1(n17494), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11091) );
  AOI22_X1 U14319 ( .A1(n17508), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11090) );
  OAI211_X1 U14320 ( .C1(n10978), .C2(n18752), .A(n11091), .B(n11090), .ZN(
        n11092) );
  AOI211_X1 U14321 ( .C1(n17512), .C2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A(
        n11093), .B(n11092), .ZN(n11094) );
  OAI211_X1 U14322 ( .C1(n10970), .C2(n17355), .A(n11095), .B(n11094), .ZN(
        n11096) );
  AOI211_X4 U14323 ( .C1(n17421), .C2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A(
        n11097), .B(n11096), .ZN(n18524) );
  NOR2_X1 U14324 ( .A1(n19186), .A2(n11186), .ZN(n11179) );
  AOI22_X1 U14325 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11107) );
  INV_X1 U14326 ( .A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n18764) );
  AOI22_X1 U14327 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17494), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11099) );
  AOI22_X1 U14328 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11098) );
  OAI211_X1 U14329 ( .C1(n10978), .C2(n18764), .A(n11099), .B(n11098), .ZN(
        n11105) );
  AOI22_X1 U14330 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11103) );
  AOI22_X1 U14331 ( .A1(n9671), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11102) );
  AOI22_X1 U14332 ( .A1(n16175), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11030), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11101) );
  NAND2_X1 U14333 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11100) );
  NAND4_X1 U14334 ( .A1(n11103), .A2(n11102), .A3(n11101), .A4(n11100), .ZN(
        n11104) );
  NAND2_X1 U14335 ( .A1(n11179), .A2(n11143), .ZN(n11200) );
  AOI22_X1 U14336 ( .A1(n17494), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11109) );
  AOI22_X1 U14337 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n16175), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11108) );
  OAI211_X1 U14338 ( .C1(n10978), .C2(n18746), .A(n11109), .B(n11108), .ZN(
        n11115) );
  AOI22_X1 U14339 ( .A1(n17508), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9670), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11113) );
  AOI22_X1 U14340 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U14341 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11111) );
  NAND2_X1 U14342 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11110) );
  NAND4_X1 U14343 ( .A1(n11113), .A2(n11112), .A3(n11111), .A4(n11110), .ZN(
        n11114) );
  NOR2_X1 U14344 ( .A1(n11186), .A2(n11252), .ZN(n11182) );
  INV_X1 U14345 ( .A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17437) );
  AOI22_X1 U14346 ( .A1(n17508), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17403), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11127) );
  INV_X1 U14347 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n18758) );
  AOI22_X1 U14348 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11119) );
  AOI22_X1 U14349 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17495), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11118) );
  OAI211_X1 U14350 ( .C1(n10978), .C2(n18758), .A(n11119), .B(n11118), .ZN(
        n11125) );
  AOI22_X1 U14351 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11123) );
  AOI22_X1 U14352 ( .A1(n17494), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11122) );
  AOI22_X1 U14353 ( .A1(n16175), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11121) );
  NAND2_X1 U14354 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11120) );
  NAND4_X1 U14355 ( .A1(n11123), .A2(n11122), .A3(n11121), .A4(n11120), .ZN(
        n11124) );
  INV_X1 U14356 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17313) );
  AOI22_X1 U14357 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17494), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11136) );
  INV_X1 U14358 ( .A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n18761) );
  OAI22_X1 U14359 ( .A1(n10978), .A2(n18761), .B1(n11128), .B2(n17537), .ZN(
        n11134) );
  AOI22_X1 U14360 ( .A1(n16175), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11132) );
  AOI22_X1 U14361 ( .A1(n9671), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11131) );
  AOI22_X1 U14362 ( .A1(n17512), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11130) );
  NAND3_X1 U14363 ( .A1(n11132), .A2(n11131), .A3(n11130), .ZN(n11133) );
  OAI211_X1 U14364 ( .C1(n10949), .C2(n17313), .A(n11136), .B(n11135), .ZN(
        n11137) );
  INV_X1 U14365 ( .A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17310) );
  AOI22_X1 U14366 ( .A1(n17508), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11138) );
  OAI21_X1 U14367 ( .B1(n10109), .B2(n17310), .A(n11138), .ZN(n11140) );
  AOI22_X1 U14368 ( .A1(n16175), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17476), .ZN(n11144) );
  OAI21_X1 U14369 ( .B1(n10949), .B2(n17412), .A(n11144), .ZN(n11154) );
  INV_X1 U14370 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17529) );
  AOI22_X1 U14371 ( .A1(n10981), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n9671), .ZN(n11152) );
  INV_X1 U14372 ( .A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11146) );
  AOI22_X1 U14373 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n9667), .B1(
        n17512), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11145) );
  OAI21_X1 U14374 ( .B1(n10970), .B2(n11146), .A(n11145), .ZN(n11150) );
  INV_X1 U14375 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n18770) );
  AOI22_X1 U14376 ( .A1(n17494), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17490), .ZN(n11148) );
  OAI211_X1 U14377 ( .C1(n18770), .C2(n10978), .A(n11148), .B(n11147), .ZN(
        n11149) );
  AOI211_X1 U14378 ( .C1(n11129), .C2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n11150), .B(n11149), .ZN(n11151) );
  OAI211_X1 U14379 ( .C1(n11128), .C2(n17529), .A(n11152), .B(n11151), .ZN(
        n11153) );
  AOI211_X4 U14380 ( .C1(n17420), .C2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A(
        n11154), .B(n11153), .ZN(n18548) );
  INV_X1 U14381 ( .A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16102) );
  OAI22_X1 U14382 ( .A1(n10949), .A2(n17452), .B1(n10948), .B2(n16102), .ZN(
        n11165) );
  AOI22_X1 U14383 ( .A1(n16175), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11164) );
  AOI22_X1 U14384 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11163) );
  AOI22_X1 U14385 ( .A1(n17514), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9670), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11155) );
  INV_X1 U14386 ( .A(n11155), .ZN(n11161) );
  AOI22_X1 U14387 ( .A1(n17508), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11159) );
  AOI22_X1 U14388 ( .A1(n17494), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11156), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11158) );
  AOI22_X1 U14389 ( .A1(n17512), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11157) );
  NAND3_X1 U14390 ( .A1(n11159), .A2(n11158), .A3(n11157), .ZN(n11160) );
  AOI211_X1 U14391 ( .C1(n17339), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n11161), .B(n11160), .ZN(n11162) );
  INV_X1 U14392 ( .A(n18529), .ZN(n11245) );
  AOI211_X1 U14393 ( .C1(n16091), .C2(n16278), .A(n11234), .B(n11254), .ZN(
        n11166) );
  NAND2_X1 U14394 ( .A1(n11182), .A2(n11166), .ZN(n11190) );
  NAND2_X1 U14395 ( .A1(n17567), .A2(n18524), .ZN(n11253) );
  INV_X1 U14396 ( .A(n11253), .ZN(n11242) );
  NAND2_X1 U14397 ( .A1(n19008), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11180) );
  XNOR2_X1 U14398 ( .A(n11180), .B(n11191), .ZN(n11177) );
  OAI22_X1 U14399 ( .A1(n10935), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n19015), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11172) );
  OAI22_X1 U14400 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19019), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11169), .ZN(n11174) );
  NOR2_X1 U14401 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n19019), .ZN(
        n11170) );
  NAND2_X1 U14402 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11169), .ZN(
        n11175) );
  AOI22_X1 U14403 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11174), .B1(
        n11170), .B2(n11175), .ZN(n11196) );
  NAND2_X1 U14404 ( .A1(n11173), .A2(n11172), .ZN(n11171) );
  OAI211_X1 U14405 ( .C1(n11173), .C2(n11172), .A(n11196), .B(n11171), .ZN(
        n11193) );
  AOI21_X1 U14406 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11175), .A(
        n11174), .ZN(n11176) );
  INV_X2 U14407 ( .A(n19194), .ZN(n19126) );
  NAND2_X2 U14408 ( .A1(n19126), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n19129) );
  OAI211_X1 U14409 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n19063), .B(n19129), .ZN(n19184) );
  OAI21_X1 U14410 ( .B1(n18524), .B2(n9725), .A(n19184), .ZN(n11178) );
  NAND2_X1 U14411 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n19187) );
  OAI21_X1 U14412 ( .B1(n11179), .B2(n11178), .A(n19187), .ZN(n16854) );
  NOR3_X1 U14413 ( .A1(n11242), .A2(n11181), .A3(n16854), .ZN(n11202) );
  OAI21_X1 U14414 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19008), .A(
        n11180), .ZN(n11192) );
  OAI21_X1 U14415 ( .B1(n11192), .B2(n11193), .A(n18970), .ZN(n11662) );
  NOR2_X1 U14416 ( .A1(n18538), .A2(n18542), .ZN(n11198) );
  AND4_X1 U14417 ( .A1(n18529), .A2(n18533), .A3(n11238), .A4(n11198), .ZN(
        n11246) );
  NAND2_X1 U14418 ( .A1(n11246), .A2(n11186), .ZN(n11237) );
  INV_X1 U14419 ( .A(n11198), .ZN(n11183) );
  NAND2_X1 U14420 ( .A1(n17691), .A2(n11183), .ZN(n11185) );
  INV_X1 U14421 ( .A(n11182), .ZN(n11184) );
  AOI22_X1 U14422 ( .A1(n11185), .A2(n16091), .B1(n11184), .B2(n11183), .ZN(
        n11188) );
  NAND2_X1 U14423 ( .A1(n18542), .A2(n16091), .ZN(n18982) );
  OAI211_X1 U14424 ( .C1(n19003), .C2(n18517), .A(n11235), .B(n18982), .ZN(
        n11187) );
  OAI211_X1 U14425 ( .C1(n11238), .C2(n11245), .A(n11188), .B(n11187), .ZN(
        n11243) );
  NOR2_X1 U14426 ( .A1(n18517), .A2(n9725), .ZN(n11251) );
  OAI21_X1 U14427 ( .B1(n18548), .B2(n19003), .A(n11251), .ZN(n11240) );
  INV_X1 U14428 ( .A(n11240), .ZN(n11189) );
  AOI211_X1 U14429 ( .C1(n11237), .C2(n11190), .A(n11243), .B(n11189), .ZN(
        n14659) );
  NOR2_X1 U14430 ( .A1(n11192), .A2(n11191), .ZN(n11197) );
  NAND2_X1 U14431 ( .A1(n11194), .A2(n11193), .ZN(n11195) );
  OAI211_X1 U14432 ( .C1(n16091), .C2(n11198), .A(n18524), .B(n18967), .ZN(
        n11199) );
  OAI211_X1 U14433 ( .C1(n11200), .C2(n11662), .A(n14659), .B(n11199), .ZN(
        n11201) );
  NAND2_X1 U14434 ( .A1(n19033), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19036) );
  NAND2_X1 U14435 ( .A1(n11732), .A2(n18429), .ZN(n18503) );
  NAND2_X1 U14436 ( .A1(n11700), .A2(n18399), .ZN(n11277) );
  NOR2_X1 U14437 ( .A1(n18196), .A2(n11726), .ZN(n16201) );
  NAND2_X1 U14438 ( .A1(n16201), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16258) );
  NAND4_X1 U14439 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11666) );
  NOR2_X1 U14440 ( .A1(n18230), .A2(n11666), .ZN(n11734) );
  NAND2_X1 U14441 ( .A1(n17712), .A2(n11207), .ZN(n11206) );
  NAND2_X1 U14442 ( .A1(n11205), .A2(n11206), .ZN(n11216) );
  NAND2_X1 U14443 ( .A1(n11204), .A2(n11203), .ZN(n11220) );
  NOR2_X1 U14444 ( .A1(n17697), .A2(n11220), .ZN(n11224) );
  NAND2_X1 U14445 ( .A1(n11224), .A2(n17692), .ZN(n11225) );
  INV_X1 U14446 ( .A(n11203), .ZN(n17701) );
  XNOR2_X1 U14447 ( .A(n17701), .B(n11204), .ZN(n11219) );
  INV_X1 U14448 ( .A(n11205), .ZN(n17708) );
  XNOR2_X1 U14449 ( .A(n11206), .B(n17708), .ZN(n11214) );
  AND2_X1 U14450 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11214), .ZN(
        n11215) );
  NOR2_X1 U14451 ( .A1(n11208), .A2(n11027), .ZN(n11213) );
  INV_X1 U14452 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19163) );
  NOR2_X1 U14453 ( .A1(n11210), .A2(n19163), .ZN(n11211) );
  INV_X1 U14454 ( .A(n18175), .ZN(n18164) );
  NAND3_X1 U14455 ( .A1(n18164), .A2(n11210), .A3(n19163), .ZN(n11209) );
  OAI221_X1 U14456 ( .B1(n11211), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n18164), .C2(n11210), .A(n11209), .ZN(n18157) );
  NOR2_X1 U14457 ( .A1(n18158), .A2(n18157), .ZN(n11212) );
  XOR2_X1 U14458 ( .A(n18465), .B(n11214), .Z(n18145) );
  NOR2_X1 U14459 ( .A1(n11217), .A2(n18450), .ZN(n11218) );
  XNOR2_X1 U14460 ( .A(n17704), .B(n11216), .ZN(n18136) );
  NOR2_X1 U14461 ( .A1(n18136), .A2(n18135), .ZN(n18134) );
  NOR2_X1 U14462 ( .A1(n11218), .A2(n18134), .ZN(n18121) );
  INV_X1 U14463 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18439) );
  XOR2_X1 U14464 ( .A(n18439), .B(n11219), .Z(n18120) );
  XNOR2_X1 U14465 ( .A(n17697), .B(n11220), .ZN(n11222) );
  NOR2_X1 U14466 ( .A1(n11221), .A2(n11222), .ZN(n11223) );
  XNOR2_X1 U14467 ( .A(n17692), .B(n11224), .ZN(n11227) );
  NAND2_X1 U14468 ( .A1(n11226), .A2(n11227), .ZN(n18094) );
  INV_X1 U14469 ( .A(n11225), .ZN(n11230) );
  OR2_X1 U14470 ( .A1(n11227), .A2(n11226), .ZN(n18095) );
  OAI21_X1 U14471 ( .B1(n11230), .B2(n11229), .A(n18095), .ZN(n11228) );
  NAND2_X1 U14472 ( .A1(n16738), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11232) );
  XOR2_X1 U14473 ( .A(n11232), .B(n19146), .Z(n11708) );
  NAND2_X1 U14474 ( .A1(n11234), .A2(n11233), .ZN(n16092) );
  NOR2_X1 U14475 ( .A1(n16092), .A2(n9725), .ZN(n11239) );
  INV_X1 U14476 ( .A(n11254), .ZN(n11236) );
  NAND4_X2 U14477 ( .A1(n11236), .A2(n18538), .A3(n11241), .A4(n17727), .ZN(
        n17765) );
  NAND2_X1 U14478 ( .A1(n11252), .A2(n16855), .ZN(n14655) );
  AOI21_X2 U14479 ( .B1(n11239), .B2(n11238), .A(n13364), .ZN(n11247) );
  OAI21_X1 U14480 ( .B1(n11242), .B2(n11241), .A(n11240), .ZN(n11244) );
  AOI21_X1 U14481 ( .B1(n11245), .B2(n11244), .A(n11243), .ZN(n11248) );
  NAND2_X1 U14482 ( .A1(n11246), .A2(n11248), .ZN(n13363) );
  NAND2_X1 U14483 ( .A1(n11247), .A2(n13363), .ZN(n18977) );
  NOR2_X1 U14484 ( .A1(n19186), .A2(n13364), .ZN(n11250) );
  INV_X1 U14485 ( .A(n11248), .ZN(n11249) );
  NOR2_X1 U14486 ( .A1(n11252), .A2(n11251), .ZN(n19195) );
  NAND2_X1 U14487 ( .A1(n18966), .A2(n18429), .ZN(n18492) );
  NAND2_X1 U14488 ( .A1(n11708), .A2(n18498), .ZN(n11276) );
  NAND2_X1 U14489 ( .A1(n16739), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11256) );
  XNOR2_X1 U14490 ( .A(n19146), .B(n11256), .ZN(n11709) );
  NOR2_X1 U14491 ( .A1(n17692), .A2(n18503), .ZN(n18413) );
  INV_X1 U14492 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n19125) );
  INV_X1 U14493 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n19147) );
  NAND2_X1 U14494 ( .A1(n19147), .A2(n19138), .ZN(n19150) );
  NOR2_X1 U14495 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n19150), .ZN(n19199) );
  NAND2_X2 U14496 ( .A1(n19199), .A2(n19039), .ZN(n18482) );
  NOR2_X1 U14497 ( .A1(n19125), .A2(n18482), .ZN(n11707) );
  NOR3_X1 U14498 ( .A1(n18278), .A2(n18433), .A3(n18423), .ZN(n18316) );
  NOR3_X1 U14499 ( .A1(n18465), .A2(n18450), .A3(n18439), .ZN(n18420) );
  INV_X1 U14500 ( .A(n18420), .ZN(n11257) );
  NAND2_X1 U14501 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18446) );
  NOR2_X1 U14502 ( .A1(n11257), .A2(n18446), .ZN(n18403) );
  NAND2_X1 U14503 ( .A1(n18316), .A2(n18403), .ZN(n18301) );
  NOR2_X1 U14504 ( .A1(n11665), .A2(n18301), .ZN(n18246) );
  NAND2_X1 U14505 ( .A1(n11734), .A2(n18246), .ZN(n11267) );
  INV_X1 U14506 ( .A(n11261), .ZN(n18286) );
  AOI21_X1 U14507 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18448) );
  NOR2_X1 U14508 ( .A1(n18448), .A2(n11257), .ZN(n18406) );
  NAND2_X1 U14509 ( .A1(n18406), .A2(n18316), .ZN(n18300) );
  NOR2_X1 U14510 ( .A1(n11665), .A2(n18300), .ZN(n11733) );
  NAND2_X1 U14511 ( .A1(n18286), .A2(n11733), .ZN(n18284) );
  NOR2_X1 U14512 ( .A1(n11258), .A2(n18284), .ZN(n18203) );
  INV_X1 U14513 ( .A(n18203), .ZN(n18224) );
  NOR2_X1 U14514 ( .A1(n11666), .A2(n18224), .ZN(n11265) );
  INV_X1 U14515 ( .A(n11265), .ZN(n11259) );
  OAI22_X1 U14516 ( .A1(n19004), .A2(n11267), .B1(n18469), .B2(n11259), .ZN(
        n11263) );
  OR2_X1 U14517 ( .A1(n19163), .A2(n18301), .ZN(n18373) );
  NOR2_X1 U14518 ( .A1(n11665), .A2(n18373), .ZN(n18299) );
  NOR2_X1 U14519 ( .A1(n11261), .A2(n11260), .ZN(n18247) );
  NAND2_X1 U14520 ( .A1(n18299), .A2(n18247), .ZN(n18249) );
  NOR3_X1 U14521 ( .A1(n18992), .A2(n11666), .A3(n18249), .ZN(n11262) );
  OAI211_X1 U14522 ( .C1(n11263), .C2(n11262), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n18429), .ZN(n16198) );
  NOR3_X1 U14523 ( .A1(n16198), .A2(n11264), .A3(n16258), .ZN(n11272) );
  INV_X1 U14524 ( .A(n18451), .ZN(n18407) );
  NAND2_X1 U14525 ( .A1(n18407), .A2(n18429), .ZN(n18483) );
  INV_X1 U14526 ( .A(n18483), .ZN(n11269) );
  NOR2_X1 U14527 ( .A1(n11265), .A2(n18469), .ZN(n18185) );
  AOI21_X1 U14528 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n18992), .ZN(n11266) );
  AOI211_X1 U14529 ( .C1(n18447), .C2(n11267), .A(n18185), .B(n11266), .ZN(
        n11722) );
  INV_X2 U14530 ( .A(n18482), .ZN(n18499) );
  NOR2_X2 U14531 ( .A1(n18499), .A2(n18429), .ZN(n18489) );
  OAI21_X1 U14532 ( .B1(n11722), .B2(n18494), .A(n18495), .ZN(n11268) );
  AOI21_X1 U14533 ( .B1(n11269), .B2(n16258), .A(n11268), .ZN(n16260) );
  OAI22_X1 U14534 ( .A1(n16260), .A2(n19146), .B1(n11270), .B2(n18483), .ZN(
        n11271) );
  NOR3_X1 U14535 ( .A1(n11707), .A2(n11272), .A3(n11271), .ZN(n11273) );
  OAI21_X1 U14536 ( .B1(n11709), .B2(n18345), .A(n11273), .ZN(n11274) );
  INV_X1 U14537 ( .A(n11274), .ZN(n11275) );
  NAND2_X1 U14538 ( .A1(n11277), .A2(n10098), .ZN(P3_U2831) );
  NAND2_X1 U14539 ( .A1(n14813), .A2(n14809), .ZN(n11287) );
  INV_X1 U14540 ( .A(n11280), .ZN(n11281) );
  OR2_X2 U14541 ( .A1(n11282), .A2(n11281), .ZN(n14814) );
  INV_X1 U14542 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n16478) );
  NOR2_X1 U14543 ( .A1(n14815), .A2(n16478), .ZN(n11283) );
  XNOR2_X1 U14544 ( .A(n14814), .B(n11283), .ZN(n11285) );
  INV_X1 U14545 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11284) );
  OAI21_X1 U14546 ( .B1(n11285), .B2(n10781), .A(n11284), .ZN(n14808) );
  INV_X1 U14547 ( .A(n11285), .ZN(n16480) );
  AND2_X1 U14548 ( .A1(n14818), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11286) );
  NAND2_X1 U14549 ( .A1(n16480), .A2(n11286), .ZN(n14810) );
  NAND2_X2 U14550 ( .A1(n20233), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n20147) );
  NOR2_X1 U14551 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n20094) );
  INV_X1 U14552 ( .A(n20094), .ZN(n20087) );
  NAND3_X1 U14553 ( .A1(n20086), .A2(n20147), .A3(n20087), .ZN(n20225) );
  NAND2_X1 U14554 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n20221) );
  NOR2_X1 U14555 ( .A1(n20225), .A2(n20215), .ZN(n14031) );
  NAND2_X1 U14556 ( .A1(n11288), .A2(n14031), .ZN(n11334) );
  NAND2_X1 U14557 ( .A1(n11289), .A2(n11336), .ZN(n11307) );
  OAI21_X1 U14558 ( .B1(n15586), .B2(n11291), .A(n11290), .ZN(n11292) );
  OAI21_X1 U14559 ( .B1(n11299), .B2(n15586), .A(n11292), .ZN(n11293) );
  NAND2_X1 U14560 ( .A1(n11293), .A2(n11354), .ZN(n11297) );
  OAI21_X1 U14561 ( .B1(n11295), .B2(n11294), .A(n10646), .ZN(n11296) );
  NAND2_X1 U14562 ( .A1(n11297), .A2(n11296), .ZN(n11302) );
  INV_X1 U14563 ( .A(n20224), .ZN(n11298) );
  NAND2_X1 U14564 ( .A1(n11298), .A2(n15586), .ZN(n11300) );
  MUX2_X1 U14565 ( .A(n11336), .B(n11300), .S(n11299), .Z(n11301) );
  NAND2_X1 U14566 ( .A1(n11302), .A2(n11301), .ZN(n11305) );
  INV_X1 U14567 ( .A(n11303), .ZN(n11304) );
  NAND2_X1 U14568 ( .A1(n11305), .A2(n11304), .ZN(n11306) );
  AOI21_X1 U14569 ( .B1(n11307), .B2(n11306), .A(n11309), .ZN(n11308) );
  MUX2_X1 U14570 ( .A(n11308), .B(n13532), .S(n20218), .Z(n11311) );
  OR2_X1 U14571 ( .A1(n14310), .A2(n9730), .ZN(n13536) );
  OAI21_X1 U14572 ( .B1(n11311), .B2(n10221), .A(n11321), .ZN(n11312) );
  INV_X1 U14573 ( .A(n11312), .ZN(n11313) );
  NAND2_X1 U14574 ( .A1(n13536), .A2(n11313), .ZN(n11333) );
  OAI21_X1 U14575 ( .B1(n13176), .B2(n11315), .A(n19538), .ZN(n11316) );
  NAND2_X1 U14576 ( .A1(n11314), .A2(n11316), .ZN(n11325) );
  NAND2_X1 U14577 ( .A1(n9730), .A2(n11321), .ZN(n11364) );
  NAND2_X1 U14578 ( .A1(n11364), .A2(n11354), .ZN(n11317) );
  NAND2_X1 U14579 ( .A1(n11317), .A2(n13338), .ZN(n11318) );
  AOI21_X1 U14580 ( .B1(n11318), .B2(n19538), .A(n10226), .ZN(n11324) );
  NAND2_X1 U14581 ( .A1(n11322), .A2(n13338), .ZN(n11320) );
  NAND2_X1 U14582 ( .A1(n11320), .A2(n11319), .ZN(n11349) );
  OR2_X1 U14583 ( .A1(n11322), .A2(n11321), .ZN(n11323) );
  NAND4_X1 U14584 ( .A1(n11325), .A2(n11324), .A3(n11349), .A4(n11323), .ZN(
        n11365) );
  INV_X1 U14585 ( .A(n11365), .ZN(n11327) );
  NAND3_X1 U14586 ( .A1(n13408), .A2(n10244), .A3(n14031), .ZN(n11326) );
  AND2_X1 U14587 ( .A1(n11327), .A2(n11326), .ZN(n13521) );
  MUX2_X1 U14588 ( .A(n10244), .B(n11288), .S(n9730), .Z(n11328) );
  NAND3_X1 U14589 ( .A1(n13408), .A2(n20221), .A3(n11328), .ZN(n11329) );
  NAND2_X1 U14590 ( .A1(n13521), .A2(n11329), .ZN(n11330) );
  NOR2_X1 U14591 ( .A1(n11331), .A2(n11330), .ZN(n11332) );
  OAI211_X1 U14592 ( .C1(n11334), .C2(n13536), .A(n11333), .B(n11332), .ZN(
        n11335) );
  NOR2_X1 U14593 ( .A1(n10642), .A2(n11336), .ZN(n20207) );
  AOI21_X1 U14594 ( .B1(n15718), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11338) );
  INV_X1 U14595 ( .A(n15842), .ZN(n11337) );
  AND2_X1 U14596 ( .A1(n11337), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15841) );
  NAND2_X1 U14597 ( .A1(n15841), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14830) );
  NOR2_X1 U14598 ( .A1(n11338), .A2(n14822), .ZN(n14683) );
  INV_X1 U14599 ( .A(n11339), .ZN(n20206) );
  NAND2_X1 U14600 ( .A1(n11340), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11342) );
  NAND2_X1 U14601 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11341) );
  OAI211_X1 U14602 ( .C1(n10747), .C2(n16478), .A(n11342), .B(n11341), .ZN(
        n11343) );
  AOI21_X1 U14603 ( .B1(n10654), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n11343), .ZN(n14834) );
  NAND2_X1 U14604 ( .A1(n11344), .A2(n9730), .ZN(n11346) );
  NAND2_X1 U14605 ( .A1(n11346), .A2(n11345), .ZN(n11347) );
  NAND2_X1 U14606 ( .A1(n11348), .A2(n15586), .ZN(n14037) );
  NAND2_X1 U14607 ( .A1(n14037), .A2(n11349), .ZN(n11351) );
  NAND2_X1 U14608 ( .A1(n11351), .A2(n11350), .ZN(n11362) );
  OAI22_X1 U14609 ( .A1(n11353), .A2(n11315), .B1(n19538), .B2(n11354), .ZN(
        n11355) );
  INV_X1 U14610 ( .A(n11355), .ZN(n11359) );
  OAI21_X1 U14611 ( .B1(n13172), .B2(n11356), .A(n11353), .ZN(n11357) );
  NAND2_X1 U14612 ( .A1(n11357), .A2(n10226), .ZN(n11358) );
  AND3_X1 U14613 ( .A1(n11360), .A2(n11359), .A3(n11358), .ZN(n11361) );
  NAND2_X1 U14614 ( .A1(n13996), .A2(n13997), .ZN(n11363) );
  NAND2_X1 U14615 ( .A1(n11388), .A2(n11363), .ZN(n11368) );
  INV_X1 U14616 ( .A(n13999), .ZN(n14022) );
  NAND2_X1 U14617 ( .A1(n11388), .A2(n14022), .ZN(n15964) );
  INV_X1 U14618 ( .A(n11388), .ZN(n11366) );
  NAND2_X1 U14619 ( .A1(n11366), .A2(n19341), .ZN(n14765) );
  INV_X1 U14620 ( .A(n11377), .ZN(n11374) );
  NAND2_X1 U14621 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16040) );
  NAND2_X1 U14622 ( .A1(n11374), .A2(n16040), .ZN(n11372) );
  NAND2_X1 U14623 ( .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n14596) );
  NOR2_X1 U14624 ( .A1(n14606), .A2(n14596), .ZN(n16070) );
  NOR2_X1 U14625 ( .A1(n10816), .A2(n16708), .ZN(n16707) );
  NOR2_X1 U14626 ( .A1(n11392), .A2(n14308), .ZN(n11369) );
  NOR2_X1 U14627 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n11369), .ZN(
        n14759) );
  INV_X1 U14628 ( .A(n14759), .ZN(n11367) );
  NAND4_X1 U14629 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n16070), .A3(
        n16707), .A4(n11367), .ZN(n11654) );
  INV_X1 U14630 ( .A(n11368), .ZN(n15967) );
  INV_X1 U14631 ( .A(n11369), .ZN(n14768) );
  NOR2_X1 U14632 ( .A1(n10290), .A2(n14768), .ZN(n14758) );
  INV_X1 U14633 ( .A(n14758), .ZN(n11652) );
  NAND2_X1 U14634 ( .A1(n15967), .A2(n11652), .ZN(n14767) );
  NAND2_X1 U14635 ( .A1(n14765), .A2(n14767), .ZN(n14372) );
  INV_X1 U14636 ( .A(n14372), .ZN(n11370) );
  NAND2_X1 U14637 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n11370), .ZN(
        n11371) );
  AOI21_X1 U14638 ( .B1(n14598), .B2(n11654), .A(n11371), .ZN(n16058) );
  NOR2_X1 U14639 ( .A1(n16058), .A2(n11377), .ZN(n16045) );
  INV_X1 U14640 ( .A(n16045), .ZN(n16693) );
  INV_X1 U14641 ( .A(n11655), .ZN(n11373) );
  NAND2_X1 U14642 ( .A1(n11374), .A2(n11373), .ZN(n11375) );
  NAND2_X1 U14643 ( .A1(n16028), .A2(n11375), .ZN(n15992) );
  NOR2_X1 U14644 ( .A1(n11377), .A2(n10617), .ZN(n11376) );
  INV_X1 U14645 ( .A(n13218), .ZN(n15928) );
  NOR2_X1 U14646 ( .A1(n11377), .A2(n15928), .ZN(n11378) );
  NOR2_X1 U14647 ( .A1(n15952), .A2(n11378), .ZN(n13225) );
  NAND2_X1 U14648 ( .A1(n14598), .A2(n13224), .ZN(n11379) );
  NAND2_X1 U14649 ( .A1(n13225), .A2(n11379), .ZN(n15923) );
  NOR2_X1 U14650 ( .A1(n15906), .A2(n15905), .ZN(n15904) );
  NOR2_X1 U14651 ( .A1(n15968), .A2(n15904), .ZN(n11380) );
  OR2_X1 U14652 ( .A1(n15923), .A2(n11380), .ZN(n15889) );
  NOR2_X1 U14653 ( .A1(n15968), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11381) );
  NOR2_X1 U14654 ( .A1(n15889), .A2(n11381), .ZN(n15878) );
  AND2_X1 U14655 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11657) );
  INV_X1 U14656 ( .A(n11657), .ZN(n15866) );
  NAND2_X1 U14657 ( .A1(n14598), .A2(n15866), .ZN(n11382) );
  AND2_X1 U14658 ( .A1(n15878), .A2(n11382), .ZN(n15839) );
  OAI21_X1 U14659 ( .B1(n15968), .B2(n15841), .A(n15839), .ZN(n14829) );
  NAND2_X1 U14660 ( .A1(n14829), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11650) );
  INV_X1 U14661 ( .A(n11384), .ZN(n11385) );
  AND2_X1 U14662 ( .A1(n11383), .A2(n11385), .ZN(n13335) );
  INV_X1 U14663 ( .A(n13335), .ZN(n14025) );
  NAND2_X1 U14664 ( .A1(n13406), .A2(n11314), .ZN(n14020) );
  NAND2_X1 U14665 ( .A1(n14020), .A2(n15586), .ZN(n11386) );
  NAND2_X1 U14666 ( .A1(n14025), .A2(n11386), .ZN(n11387) );
  INV_X1 U14667 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n19227) );
  NAND2_X1 U14668 ( .A1(n19565), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11391) );
  OAI211_X1 U14669 ( .C1(n9730), .C2(n11392), .A(n11391), .B(n20195), .ZN(
        n11393) );
  INV_X1 U14670 ( .A(n11393), .ZN(n11394) );
  OAI21_X1 U14671 ( .B1(n11632), .B2(n19227), .A(n11394), .ZN(n13609) );
  INV_X1 U14672 ( .A(n11395), .ZN(n11396) );
  NAND2_X1 U14673 ( .A1(n11396), .A2(n11602), .ZN(n11399) );
  MUX2_X1 U14674 ( .A(n13338), .B(n20202), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n11398) );
  NAND2_X1 U14675 ( .A1(n11397), .A2(n13176), .ZN(n11411) );
  NAND3_X1 U14676 ( .A1(n11399), .A2(n11398), .A3(n11411), .ZN(n13610) );
  INV_X1 U14677 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19495) );
  INV_X1 U14678 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n20102) );
  OR2_X1 U14679 ( .A1(n11632), .A2(n20102), .ZN(n11401) );
  NAND2_X1 U14680 ( .A1(n11397), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11400) );
  NOR2_X1 U14681 ( .A1(n13176), .A2(n19565), .ZN(n13646) );
  MUX2_X1 U14682 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n13646), .S(
        n20195), .Z(n11404) );
  AND2_X1 U14683 ( .A1(n11602), .A2(n11402), .ZN(n11403) );
  NOR2_X1 U14684 ( .A1(n11404), .A2(n11403), .ZN(n13628) );
  INV_X1 U14685 ( .A(n13628), .ZN(n11405) );
  NOR2_X1 U14686 ( .A1(n13612), .A2(n11406), .ZN(n11407) );
  NOR2_X2 U14687 ( .A1(n11408), .A2(n11407), .ZN(n11415) );
  NAND2_X1 U14688 ( .A1(n11602), .A2(n11409), .ZN(n11410) );
  OAI211_X1 U14689 ( .C1(n20195), .C2(n20182), .A(n11411), .B(n11410), .ZN(
        n11414) );
  INV_X1 U14690 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19493) );
  INV_X1 U14691 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n20104) );
  OR2_X1 U14692 ( .A1(n11632), .A2(n20104), .ZN(n11413) );
  NAND2_X1 U14693 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11412) );
  OAI211_X1 U14694 ( .C1(n19493), .C2(n11421), .A(n11413), .B(n11412), .ZN(
        n13914) );
  INV_X1 U14695 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n11419) );
  AOI22_X1 U14696 ( .A1(P2_EAX_REG_3__SCAN_IN), .A2(n14823), .B1(n11602), .B2(
        n11416), .ZN(n11418) );
  AOI22_X1 U14697 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11417) );
  OAI211_X1 U14698 ( .C1(n11419), .C2(n11632), .A(n11418), .B(n11417), .ZN(
        n13968) );
  INV_X1 U14699 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n14221) );
  OR2_X1 U14700 ( .A1(n11632), .A2(n14221), .ZN(n11425) );
  NAND2_X1 U14701 ( .A1(n11602), .A2(n11420), .ZN(n11424) );
  INV_X1 U14702 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n14276) );
  OR2_X1 U14703 ( .A1(n11421), .A2(n14276), .ZN(n11423) );
  NAND2_X1 U14704 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11422) );
  AOI22_X1 U14705 ( .A1(n14824), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n11638), 
        .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U14706 ( .A1(n14823), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n11602), .B2(
        n11426), .ZN(n11427) );
  NAND2_X1 U14707 ( .A1(n11428), .A2(n11427), .ZN(n14451) );
  NAND2_X1 U14708 ( .A1(n14452), .A2(n14451), .ZN(n14450) );
  INV_X1 U14709 ( .A(n11429), .ZN(n11430) );
  NAND2_X1 U14710 ( .A1(n11602), .A2(n11430), .ZN(n11431) );
  INV_X1 U14711 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19486) );
  INV_X1 U14712 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n20109) );
  OR2_X1 U14713 ( .A1(n11632), .A2(n20109), .ZN(n11433) );
  NAND2_X1 U14714 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11432) );
  OAI211_X1 U14715 ( .C1(n19486), .C2(n11421), .A(n11433), .B(n11432), .ZN(
        n13668) );
  NAND2_X1 U14716 ( .A1(n13670), .A2(n13668), .ZN(n11435) );
  NAND2_X1 U14717 ( .A1(n11602), .A2(n14818), .ZN(n11434) );
  NAND2_X2 U14718 ( .A1(n11435), .A2(n11434), .ZN(n13667) );
  INV_X1 U14719 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19483) );
  INV_X1 U14720 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n20111) );
  OR2_X1 U14721 ( .A1(n11632), .A2(n20111), .ZN(n11437) );
  NAND2_X1 U14722 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11436) );
  OAI211_X1 U14723 ( .C1(n19483), .C2(n11421), .A(n11437), .B(n11436), .ZN(
        n13666) );
  INV_X1 U14724 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n11438) );
  OR2_X1 U14725 ( .A1(n11632), .A2(n11438), .ZN(n11456) );
  INV_X1 U14726 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11441) );
  NAND2_X1 U14727 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11440) );
  NAND2_X1 U14728 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11439) );
  OAI211_X1 U14729 ( .C1(n12963), .C2(n11441), .A(n11440), .B(n11439), .ZN(
        n11444) );
  INV_X1 U14730 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11442) );
  INV_X1 U14731 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12826) );
  OAI22_X1 U14732 ( .A1(n12897), .A2(n11442), .B1(n12896), .B2(n12826), .ZN(
        n11443) );
  NOR2_X1 U14733 ( .A1(n11444), .A2(n11443), .ZN(n11452) );
  AOI22_X1 U14734 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10460), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11448) );
  AOI22_X1 U14735 ( .A1(n10385), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11447) );
  AOI22_X1 U14736 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11446) );
  NAND2_X1 U14737 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11445) );
  AND4_X1 U14738 ( .A1(n11448), .A2(n11447), .A3(n11446), .A4(n11445), .ZN(
        n11451) );
  AOI22_X1 U14739 ( .A1(n12905), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12904), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U14740 ( .A1(n12907), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12906), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11449) );
  NAND4_X1 U14741 ( .A1(n11452), .A2(n11451), .A3(n11450), .A4(n11449), .ZN(
        n13849) );
  NAND2_X1 U14742 ( .A1(n11602), .A2(n13849), .ZN(n11455) );
  NAND2_X1 U14743 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11454) );
  INV_X1 U14744 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n13423) );
  OR2_X1 U14745 ( .A1(n11421), .A2(n13423), .ZN(n11453) );
  OAI22_X1 U14746 ( .A1(n12963), .A2(n11458), .B1(n12956), .B2(n11457), .ZN(
        n11460) );
  OAI22_X1 U14747 ( .A1(n13014), .A2(n12951), .B1(n12955), .B2(n12844), .ZN(
        n11459) );
  OR2_X1 U14748 ( .A1(n11460), .A2(n11459), .ZN(n11466) );
  AOI22_X1 U14749 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10385), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U14750 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10460), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U14751 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10384), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11462) );
  NAND2_X1 U14752 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11461) );
  NAND4_X1 U14753 ( .A1(n11464), .A2(n11463), .A3(n11462), .A4(n11461), .ZN(
        n11465) );
  NOR2_X1 U14754 ( .A1(n11466), .A2(n11465), .ZN(n11474) );
  OAI22_X1 U14755 ( .A1(n11467), .A2(n12897), .B1(n12953), .B2(n13005), .ZN(
        n11472) );
  NAND2_X1 U14756 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11469) );
  NAND2_X1 U14757 ( .A1(n12960), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11468) );
  OAI211_X1 U14758 ( .C1(n10099), .C2(n11470), .A(n11469), .B(n11468), .ZN(
        n11471) );
  NOR2_X1 U14759 ( .A1(n11472), .A2(n11471), .ZN(n11473) );
  INV_X1 U14760 ( .A(n11602), .ZN(n11477) );
  AOI22_X1 U14761 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n14823), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n11476) );
  NAND2_X1 U14762 ( .A1(n14824), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n11475) );
  OAI211_X1 U14763 ( .C1(n13909), .C2(n11477), .A(n11476), .B(n11475), .ZN(
        n13760) );
  INV_X1 U14764 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n11478) );
  OR2_X1 U14765 ( .A1(n11632), .A2(n11478), .ZN(n11501) );
  NAND2_X1 U14766 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11480) );
  NAND2_X1 U14767 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11479) );
  OAI211_X1 U14768 ( .C1(n12963), .C2(n11481), .A(n11480), .B(n11479), .ZN(
        n11485) );
  INV_X1 U14769 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11483) );
  INV_X1 U14770 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11482) );
  OAI22_X1 U14771 ( .A1(n12897), .A2(n11483), .B1(n12896), .B2(n11482), .ZN(
        n11484) );
  NOR2_X1 U14772 ( .A1(n11485), .A2(n11484), .ZN(n11497) );
  AOI22_X1 U14773 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10460), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U14774 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10385), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U14775 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10395), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11487) );
  NAND2_X1 U14776 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11486) );
  AND4_X1 U14777 ( .A1(n11489), .A2(n11488), .A3(n11487), .A4(n11486), .ZN(
        n11496) );
  INV_X1 U14778 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11491) );
  INV_X1 U14779 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11490) );
  OAI22_X1 U14780 ( .A1(n12953), .A2(n11491), .B1(n12951), .B2(n11490), .ZN(
        n11494) );
  INV_X1 U14781 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11492) );
  INV_X1 U14782 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13037) );
  OAI22_X1 U14783 ( .A1(n11492), .A2(n12956), .B1(n12955), .B2(n13037), .ZN(
        n11493) );
  NOR2_X1 U14784 ( .A1(n11494), .A2(n11493), .ZN(n11495) );
  AND3_X1 U14785 ( .A1(n11497), .A2(n11496), .A3(n11495), .ZN(n13927) );
  INV_X1 U14786 ( .A(n13927), .ZN(n13929) );
  NAND2_X1 U14787 ( .A1(n11602), .A2(n13929), .ZN(n11500) );
  NAND2_X1 U14788 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11499) );
  INV_X1 U14789 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n13520) );
  OR2_X1 U14790 ( .A1(n11421), .A2(n13520), .ZN(n11498) );
  INV_X1 U14791 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n13514) );
  NAND2_X1 U14792 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11522) );
  AOI22_X1 U14793 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10385), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14794 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10460), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14795 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10384), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11503) );
  NAND2_X1 U14796 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11502) );
  NAND4_X1 U14797 ( .A1(n11505), .A2(n11504), .A3(n11503), .A4(n11502), .ZN(
        n11511) );
  NAND2_X1 U14798 ( .A1(n12960), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11509) );
  NAND2_X1 U14799 ( .A1(n12905), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11508) );
  NAND2_X1 U14800 ( .A1(n12906), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11507) );
  NAND2_X1 U14801 ( .A1(n12904), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11506) );
  NAND4_X1 U14802 ( .A1(n11509), .A2(n11508), .A3(n11507), .A4(n11506), .ZN(
        n11510) );
  NOR2_X1 U14803 ( .A1(n11511), .A2(n11510), .ZN(n11520) );
  OAI22_X1 U14804 ( .A1(n11513), .A2(n12953), .B1(n12897), .B2(n11512), .ZN(
        n11518) );
  INV_X1 U14805 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11516) );
  NAND2_X1 U14806 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11515) );
  NAND2_X1 U14807 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11514) );
  OAI211_X1 U14808 ( .C1(n12963), .C2(n11516), .A(n11515), .B(n11514), .ZN(
        n11517) );
  NOR2_X1 U14809 ( .A1(n11518), .A2(n11517), .ZN(n11519) );
  AND2_X1 U14810 ( .A1(n11520), .A2(n11519), .ZN(n12821) );
  INV_X1 U14811 ( .A(n12821), .ZN(n13940) );
  NAND2_X1 U14812 ( .A1(n11602), .A2(n13940), .ZN(n11521) );
  OAI211_X1 U14813 ( .C1(n11421), .C2(n13514), .A(n11522), .B(n11521), .ZN(
        n11525) );
  INV_X1 U14814 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n11523) );
  NOR2_X1 U14815 ( .A1(n11632), .A2(n11523), .ZN(n11524) );
  INV_X1 U14816 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n11526) );
  OR2_X1 U14817 ( .A1(n11632), .A2(n11526), .ZN(n11545) );
  NAND2_X1 U14818 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11528) );
  NAND2_X1 U14819 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11527) );
  OAI211_X1 U14820 ( .C1(n12963), .C2(n11529), .A(n11528), .B(n11527), .ZN(
        n11532) );
  INV_X1 U14821 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11530) );
  OAI22_X1 U14822 ( .A1(n12897), .A2(n11530), .B1(n12896), .B2(n12894), .ZN(
        n11531) );
  NOR2_X1 U14823 ( .A1(n11532), .A2(n11531), .ZN(n11540) );
  AOI22_X1 U14824 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10460), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14825 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10385), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14826 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10395), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11534) );
  NAND2_X1 U14827 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11533) );
  AND4_X1 U14828 ( .A1(n11536), .A2(n11535), .A3(n11534), .A4(n11533), .ZN(
        n11539) );
  AOI22_X1 U14829 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12905), .B1(
        n12904), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11538) );
  AOI22_X1 U14830 ( .A1(n12907), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12906), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11537) );
  NAND4_X1 U14831 ( .A1(n11540), .A2(n11539), .A3(n11538), .A4(n11537), .ZN(
        n13986) );
  NAND2_X1 U14832 ( .A1(n11602), .A2(n13986), .ZN(n11544) );
  NAND2_X1 U14833 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11543) );
  INV_X1 U14834 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n11541) );
  OR2_X1 U14835 ( .A1(n11421), .A2(n11541), .ZN(n11542) );
  INV_X1 U14836 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n13426) );
  NAND2_X1 U14837 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11563) );
  NAND2_X1 U14838 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11547) );
  NAND2_X1 U14839 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11546) );
  OAI211_X1 U14840 ( .C1(n12963), .C2(n11548), .A(n11547), .B(n11546), .ZN(
        n11551) );
  OAI22_X1 U14841 ( .A1(n12953), .A2(n11549), .B1(n12951), .B2(n13107), .ZN(
        n11550) );
  NOR2_X1 U14842 ( .A1(n11551), .A2(n11550), .ZN(n11561) );
  AOI22_X1 U14843 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10385), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14844 ( .A1(n10460), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U14845 ( .A1(n10384), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11553) );
  NAND2_X1 U14846 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11552) );
  AND4_X1 U14847 ( .A1(n11555), .A2(n11554), .A3(n11553), .A4(n11552), .ZN(
        n11560) );
  OAI22_X1 U14848 ( .A1(n12897), .A2(n13116), .B1(n12955), .B2(n13117), .ZN(
        n11558) );
  OAI22_X1 U14849 ( .A1(n12896), .A2(n13114), .B1(n12956), .B2(n11556), .ZN(
        n11557) );
  NOR2_X1 U14850 ( .A1(n11558), .A2(n11557), .ZN(n11559) );
  NAND3_X1 U14851 ( .A1(n11561), .A2(n11560), .A3(n11559), .ZN(n14075) );
  NAND2_X1 U14852 ( .A1(n11602), .A2(n14075), .ZN(n11562) );
  OAI211_X1 U14853 ( .C1(n11421), .C2(n13426), .A(n11563), .B(n11562), .ZN(
        n11566) );
  INV_X1 U14854 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n11564) );
  NOR2_X1 U14855 ( .A1(n11632), .A2(n11564), .ZN(n11565) );
  INV_X1 U14856 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n11567) );
  OR2_X1 U14857 ( .A1(n11632), .A2(n11567), .ZN(n11588) );
  AOI22_X1 U14858 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10460), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U14859 ( .A1(n10385), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14860 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11569) );
  NAND2_X1 U14861 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11568) );
  NAND4_X1 U14862 ( .A1(n11571), .A2(n11570), .A3(n11569), .A4(n11568), .ZN(
        n11577) );
  OAI22_X1 U14863 ( .A1(n12953), .A2(n11573), .B1(n12951), .B2(n11572), .ZN(
        n11576) );
  OAI22_X1 U14864 ( .A1(n12956), .A2(n11574), .B1(n12955), .B2(n13127), .ZN(
        n11575) );
  OR3_X1 U14865 ( .A1(n11577), .A2(n11576), .A3(n11575), .ZN(n11583) );
  AOI22_X1 U14866 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11581) );
  NAND2_X1 U14867 ( .A1(n12961), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11580) );
  NAND2_X1 U14868 ( .A1(n12960), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11579) );
  INV_X1 U14869 ( .A(n12963), .ZN(n12939) );
  NAND2_X1 U14870 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11578) );
  NAND4_X1 U14871 ( .A1(n11581), .A2(n11580), .A3(n11579), .A4(n11578), .ZN(
        n11582) );
  NAND2_X1 U14872 ( .A1(n11602), .A2(n9744), .ZN(n11587) );
  NAND2_X1 U14873 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11586) );
  INV_X1 U14874 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n11584) );
  OR2_X1 U14875 ( .A1(n11421), .A2(n11584), .ZN(n11585) );
  NAND2_X1 U14876 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11590) );
  NAND2_X1 U14877 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11589) );
  OAI211_X1 U14878 ( .C1(n12963), .C2(n11591), .A(n11590), .B(n11589), .ZN(
        n11593) );
  INV_X1 U14879 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12966) );
  INV_X1 U14880 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12962) );
  OAI22_X1 U14881 ( .A1(n12897), .A2(n12966), .B1(n12896), .B2(n12962), .ZN(
        n11592) );
  NOR2_X1 U14882 ( .A1(n11593), .A2(n11592), .ZN(n11601) );
  AOI22_X1 U14883 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10460), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14884 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10385), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U14885 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11595) );
  NAND2_X1 U14886 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11594) );
  AND4_X1 U14887 ( .A1(n11597), .A2(n11596), .A3(n11595), .A4(n11594), .ZN(
        n11600) );
  AOI22_X1 U14888 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n12905), .B1(
        n12904), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U14889 ( .A1(n12907), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12906), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11598) );
  NAND4_X1 U14890 ( .A1(n11601), .A2(n11600), .A3(n11599), .A4(n11598), .ZN(
        n14336) );
  AOI22_X1 U14891 ( .A1(n14824), .A2(P2_REIP_REG_15__SCAN_IN), .B1(n11602), 
        .B2(n14336), .ZN(n11604) );
  AOI22_X1 U14892 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n11638), .B1(
        n14823), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n11603) );
  NAND2_X1 U14893 ( .A1(n11604), .A2(n11603), .ZN(n14354) );
  INV_X1 U14894 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15977) );
  OR2_X1 U14895 ( .A1(n11632), .A2(n15977), .ZN(n11607) );
  NAND2_X1 U14896 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11606) );
  INV_X1 U14897 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n13490) );
  OR2_X1 U14898 ( .A1(n11421), .A2(n13490), .ZN(n11605) );
  INV_X1 U14899 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13731) );
  INV_X1 U14900 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n20123) );
  OR2_X1 U14901 ( .A1(n11632), .A2(n20123), .ZN(n11609) );
  NAND2_X1 U14902 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11608) );
  OAI211_X1 U14903 ( .C1(n13731), .C2(n11421), .A(n11609), .B(n11608), .ZN(
        n15971) );
  INV_X1 U14904 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n20125) );
  OR2_X1 U14905 ( .A1(n11632), .A2(n20125), .ZN(n11612) );
  NAND2_X1 U14906 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11611) );
  INV_X1 U14907 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13485) );
  OR2_X1 U14908 ( .A1(n11421), .A2(n13485), .ZN(n11610) );
  INV_X1 U14909 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n20127) );
  OR2_X1 U14910 ( .A1(n11632), .A2(n20127), .ZN(n11615) );
  NAND2_X1 U14911 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11614) );
  INV_X1 U14912 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14638) );
  OR2_X1 U14913 ( .A1(n11421), .A2(n14638), .ZN(n11613) );
  INV_X1 U14914 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13418) );
  INV_X1 U14915 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n20129) );
  OR2_X1 U14916 ( .A1(n11632), .A2(n20129), .ZN(n11618) );
  NAND2_X1 U14917 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11617) );
  OAI211_X1 U14918 ( .C1(n11421), .C2(n13418), .A(n11618), .B(n11617), .ZN(
        n15686) );
  AND2_X2 U14919 ( .A1(n14636), .A2(n15686), .ZN(n15688) );
  INV_X1 U14920 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15680) );
  OAI222_X1 U14921 ( .A1(n11632), .A2(n20131), .B1(n11421), .B2(n15680), .C1(
        n13224), .C2(n9683), .ZN(n13216) );
  NAND2_X2 U14922 ( .A1(n15688), .A2(n13216), .ZN(n15673) );
  INV_X1 U14923 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n11619) );
  OR2_X1 U14924 ( .A1(n11632), .A2(n11619), .ZN(n11622) );
  NAND2_X1 U14925 ( .A1(n9735), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11621) );
  INV_X1 U14926 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n13506) );
  OR2_X1 U14927 ( .A1(n11421), .A2(n13506), .ZN(n11620) );
  INV_X1 U14928 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15666) );
  INV_X1 U14929 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n20134) );
  OR2_X1 U14930 ( .A1(n11632), .A2(n20134), .ZN(n11624) );
  NAND2_X1 U14931 ( .A1(n11638), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11623) );
  OAI211_X1 U14932 ( .C1(n15666), .C2(n11421), .A(n11624), .B(n11623), .ZN(
        n15668) );
  INV_X1 U14933 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n20136) );
  OR2_X1 U14934 ( .A1(n11632), .A2(n20136), .ZN(n11627) );
  NAND2_X1 U14935 ( .A1(n9735), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11626) );
  INV_X1 U14936 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13509) );
  OR2_X1 U14937 ( .A1(n11421), .A2(n13509), .ZN(n11625) );
  INV_X1 U14938 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15653) );
  INV_X1 U14939 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n20138) );
  OR2_X1 U14940 ( .A1(n11632), .A2(n20138), .ZN(n11629) );
  NAND2_X1 U14941 ( .A1(n9735), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11628) );
  OAI211_X1 U14942 ( .C1(n15653), .C2(n11421), .A(n11629), .B(n11628), .ZN(
        n15651) );
  INV_X1 U14943 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n20140) );
  OR2_X1 U14944 ( .A1(n11632), .A2(n20140), .ZN(n11631) );
  NAND2_X1 U14945 ( .A1(n14823), .A2(P2_EAX_REG_26__SCAN_IN), .ZN(n11630) );
  OAI211_X1 U14946 ( .C1(n9683), .C2(n15872), .A(n11631), .B(n11630), .ZN(
        n15642) );
  AOI22_X1 U14947 ( .A1(n9735), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n14823), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n11634) );
  INV_X1 U14948 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n20143) );
  OR2_X1 U14949 ( .A1(n11632), .A2(n20143), .ZN(n11633) );
  AND2_X1 U14950 ( .A1(n11634), .A2(n11633), .ZN(n15633) );
  INV_X1 U14951 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n15720) );
  OR2_X1 U14952 ( .A1(n11632), .A2(n15720), .ZN(n11636) );
  NAND2_X1 U14953 ( .A1(n14823), .A2(P2_EAX_REG_28__SCAN_IN), .ZN(n11635) );
  OAI211_X1 U14954 ( .C1(n9683), .C2(n11637), .A(n11636), .B(n11635), .ZN(
        n15537) );
  AOI22_X1 U14955 ( .A1(n9735), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n14823), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n11640) );
  INV_X1 U14956 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20145) );
  OR2_X1 U14957 ( .A1(n11632), .A2(n20145), .ZN(n11639) );
  AND2_X1 U14958 ( .A1(n11640), .A2(n11639), .ZN(n15620) );
  AOI22_X1 U14959 ( .A1(n9735), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n14823), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n11642) );
  INV_X1 U14960 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n20148) );
  OR2_X1 U14961 ( .A1(n11632), .A2(n20148), .ZN(n11641) );
  AND2_X1 U14962 ( .A1(n11642), .A2(n11641), .ZN(n11645) );
  INV_X1 U14963 ( .A(n11645), .ZN(n11643) );
  NAND2_X1 U14964 ( .A1(n11646), .A2(n11645), .ZN(n11647) );
  INV_X1 U14965 ( .A(n13189), .ZN(n11648) );
  INV_X2 U14966 ( .A(n19341), .ZN(n19500) );
  INV_X1 U14967 ( .A(n19500), .ZN(n19395) );
  NOR2_X1 U14968 ( .A1(n19395), .A2(n20148), .ZN(n14676) );
  OAI211_X1 U14969 ( .C1(n16481), .C2(n16716), .A(n11650), .B(n11649), .ZN(
        n11651) );
  INV_X1 U14970 ( .A(n11651), .ZN(n11659) );
  NAND2_X1 U14971 ( .A1(n15964), .A2(n11652), .ZN(n11653) );
  NAND2_X1 U14972 ( .A1(n14598), .A2(n11653), .ZN(n14454) );
  NOR2_X1 U14973 ( .A1(n14454), .A2(n11654), .ZN(n16057) );
  NAND2_X1 U14974 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16057), .ZN(
        n16695) );
  NAND2_X1 U14975 ( .A1(n16680), .A2(n11655), .ZN(n15995) );
  NOR3_X1 U14976 ( .A1(n15944), .A2(n13224), .A3(n13218), .ZN(n15903) );
  AND3_X1 U14977 ( .A1(n15903), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15904), .ZN(n15885) );
  NAND2_X1 U14978 ( .A1(n15885), .A2(n11657), .ZN(n15857) );
  INV_X1 U14979 ( .A(n15841), .ZN(n11658) );
  NAND2_X1 U14980 ( .A1(n11659), .A2(n10107), .ZN(n11660) );
  AOI21_X1 U14981 ( .B1(n14683), .B2(n16700), .A(n11660), .ZN(n11661) );
  OAI21_X1 U14982 ( .B1(n14685), .B2(n16704), .A(n11661), .ZN(P2_U3016) );
  AOI22_X1 U14983 ( .A1(n18066), .A2(n11726), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18080), .ZN(n11728) );
  INV_X1 U14984 ( .A(n11662), .ZN(n18971) );
  NAND2_X1 U14985 ( .A1(n19180), .A2(n9725), .ZN(n16094) );
  AOI211_X1 U14986 ( .C1(n11663), .C2(n11728), .A(n11717), .B(n18093), .ZN(
        n11683) );
  NOR2_X2 U14988 ( .A1(n18078), .A2(n11665), .ZN(n17914) );
  INV_X1 U14989 ( .A(n17841), .ZN(n11681) );
  NAND2_X1 U14990 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n11726), .ZN(
        n11735) );
  NOR2_X1 U14991 ( .A1(n18090), .A2(n18150), .ZN(n17934) );
  INV_X1 U14992 ( .A(n17934), .ZN(n11667) );
  AOI22_X1 U14993 ( .A1(n18090), .A2(n16199), .B1(n18150), .B2(n18190), .ZN(
        n17849) );
  NAND2_X1 U14994 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17849), .ZN(
        n17840) );
  NAND3_X1 U14995 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n11667), .A3(
        n17840), .ZN(n11671) );
  NAND2_X1 U14996 ( .A1(n19039), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17977) );
  INV_X1 U14997 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n19029) );
  NAND2_X1 U14998 ( .A1(n19029), .A2(n19138), .ZN(n16852) );
  AND2_X1 U14999 ( .A1(n19150), .A2(n16852), .ZN(n19179) );
  INV_X1 U15000 ( .A(n17977), .ZN(n18019) );
  NAND2_X1 U15001 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17857) );
  INV_X1 U15002 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n18169) );
  NAND2_X1 U15003 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n18083) );
  NOR3_X1 U15004 ( .A1(n18083), .A2(n17097), .A3(n18058), .ZN(n17064) );
  NAND2_X1 U15005 ( .A1(n18082), .A2(n17064), .ZN(n18006) );
  NAND2_X1 U15006 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n18021) );
  NOR2_X1 U15007 ( .A1(n18021), .A2(n18008), .ZN(n13360) );
  NAND2_X1 U15008 ( .A1(n17979), .A2(n13360), .ZN(n17975) );
  NAND2_X1 U15009 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17982) );
  NAND2_X1 U15010 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17942) );
  INV_X1 U15011 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17918) );
  INV_X1 U15012 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n13399) );
  NOR2_X1 U15013 ( .A1(n17918), .A2(n13399), .ZN(n13382) );
  INV_X1 U15014 ( .A(n13382), .ZN(n17908) );
  NAND2_X1 U15015 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17887), .ZN(
        n11668) );
  NOR2_X1 U15016 ( .A1(n18169), .A2(n11668), .ZN(n13388) );
  INV_X1 U15017 ( .A(n13388), .ZN(n13387) );
  OR2_X1 U15018 ( .A1(n17857), .A2(n13387), .ZN(n13380) );
  INV_X1 U15019 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n19185) );
  NOR2_X1 U15020 ( .A1(n19147), .A2(n19185), .ZN(n17976) );
  INV_X1 U15021 ( .A(n17976), .ZN(n18081) );
  OAI21_X1 U15022 ( .B1(n11672), .B2(n18081), .A(n18176), .ZN(n11669) );
  AOI21_X1 U15023 ( .B1(n18019), .B2(n13380), .A(n11669), .ZN(n17854) );
  OAI21_X1 U15024 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17929), .A(
        n17854), .ZN(n17834) );
  INV_X1 U15025 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17838) );
  NOR2_X1 U15026 ( .A1(n16876), .A2(n17838), .ZN(n16875) );
  NAND2_X1 U15027 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n11676) );
  INV_X1 U15028 ( .A(n11676), .ZN(n11673) );
  OAI21_X1 U15029 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16875), .A(
        n11693), .ZN(n16874) );
  NAND2_X1 U15030 ( .A1(n18349), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n11739) );
  NAND2_X1 U15031 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18504) );
  INV_X1 U15032 ( .A(n18504), .ZN(n11674) );
  NAND2_X1 U15033 ( .A1(n18976), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n19149) );
  OAI21_X1 U15034 ( .B1(n19189), .B2(n11674), .A(n19149), .ZN(n18515) );
  NAND3_X1 U15035 ( .A1(n19029), .A2(n19138), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18876) );
  NOR2_X4 U15036 ( .A1(n18667), .A2(n18876), .ZN(n18545) );
  INV_X1 U15037 ( .A(n11672), .ZN(n11675) );
  NOR2_X1 U15038 ( .A1(n17941), .A2(n11675), .ZN(n17839) );
  OAI211_X1 U15039 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17839), .B(n11676), .ZN(n11677) );
  OAI211_X1 U15040 ( .C1(n18024), .C2(n16874), .A(n11739), .B(n11677), .ZN(
        n11678) );
  OR2_X1 U15041 ( .A1(n11683), .A2(n11682), .ZN(P3_U2802) );
  INV_X1 U15042 ( .A(n16199), .ZN(n18188) );
  NAND2_X1 U15043 ( .A1(n18188), .A2(n16201), .ZN(n11718) );
  AOI211_X1 U15044 ( .C1(n16200), .C2(n11718), .A(n16739), .B(n18027), .ZN(
        n11684) );
  INV_X1 U15045 ( .A(n11684), .ZN(n11699) );
  INV_X1 U15046 ( .A(n18190), .ZN(n16196) );
  NAND2_X1 U15047 ( .A1(n16201), .A2(n16196), .ZN(n11723) );
  AOI211_X1 U15048 ( .C1(n16200), .C2(n11723), .A(n16738), .B(n18180), .ZN(
        n11685) );
  INV_X1 U15049 ( .A(n11685), .ZN(n11698) );
  INV_X1 U15050 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16901) );
  NAND3_X1 U15051 ( .A1(n11672), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11691) );
  NOR2_X1 U15052 ( .A1(n16901), .A2(n11691), .ZN(n11702) );
  INV_X1 U15053 ( .A(n11702), .ZN(n11689) );
  AOI22_X1 U15054 ( .A1(n18019), .A2(n11693), .B1(n18545), .B2(n11689), .ZN(
        n11690) );
  NAND2_X1 U15055 ( .A1(n11690), .A2(n18176), .ZN(n11703) );
  OAI21_X1 U15056 ( .B1(n18741), .B2(n11691), .A(n16901), .ZN(n11692) );
  AOI22_X1 U15057 ( .A1(n18349), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n11703), 
        .B2(n11692), .ZN(n11695) );
  NOR2_X1 U15058 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17929), .ZN(
        n11704) );
  AOI21_X1 U15059 ( .B1(n16901), .B2(n11693), .A(n16733), .ZN(n16900) );
  OAI21_X1 U15060 ( .B1(n11704), .B2(n18036), .A(n16900), .ZN(n11694) );
  OAI211_X1 U15061 ( .C1(n16204), .C2(n18093), .A(n11695), .B(n11694), .ZN(
        n11696) );
  INV_X1 U15062 ( .A(n11696), .ZN(n11697) );
  NAND3_X1 U15063 ( .A1(n11699), .A2(n11698), .A3(n11697), .ZN(P3_U2801) );
  NAND2_X1 U15064 ( .A1(n11700), .A2(n18075), .ZN(n11714) );
  NAND2_X1 U15065 ( .A1(n16733), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11701) );
  INV_X1 U15066 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16885) );
  INV_X1 U15067 ( .A(n17941), .ZN(n17980) );
  NAND2_X1 U15068 ( .A1(n11702), .A2(n17980), .ZN(n16736) );
  XNOR2_X1 U15069 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n11705) );
  NOR2_X1 U15070 ( .A1(n11704), .A2(n11703), .ZN(n16735) );
  OAI22_X1 U15071 ( .A1(n16736), .A2(n11705), .B1(n16735), .B2(n16885), .ZN(
        n11706) );
  AOI211_X1 U15072 ( .C1(n18036), .C2(n9724), .A(n11707), .B(n11706), .ZN(
        n11712) );
  NOR2_X1 U15073 ( .A1(n11709), .A2(n18027), .ZN(n11710) );
  NAND2_X1 U15074 ( .A1(n11714), .A2(n11713), .ZN(P3_U2799) );
  OAI21_X1 U15075 ( .B1(n11717), .B2(n10110), .A(n17692), .ZN(n11721) );
  INV_X1 U15076 ( .A(n11719), .ZN(n11720) );
  NAND2_X1 U15077 ( .A1(n18469), .A2(n19004), .ZN(n18303) );
  OAI21_X1 U15078 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n18386), .A(
        n11722), .ZN(n16193) );
  NOR2_X1 U15079 ( .A1(n18499), .A2(n11726), .ZN(n11731) );
  NOR4_X1 U15080 ( .A1(n18080), .A2(n18196), .A3(n11725), .A4(n18503), .ZN(
        n11727) );
  AND3_X1 U15081 ( .A1(n11728), .A2(n18399), .A3(n17836), .ZN(n11729) );
  INV_X1 U15082 ( .A(n11732), .ZN(n18972) );
  NOR2_X1 U15083 ( .A1(n17692), .A2(n18972), .ZN(n18371) );
  INV_X1 U15084 ( .A(n18371), .ZN(n18354) );
  OAI22_X1 U15085 ( .A1(n18240), .A2(n18312), .B1(n18313), .B2(n18354), .ZN(
        n18279) );
  INV_X1 U15086 ( .A(n11733), .ZN(n18244) );
  INV_X1 U15087 ( .A(n18246), .ZN(n18183) );
  AOI21_X1 U15088 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n19002), .A(
        n18977), .ZN(n18467) );
  OAI22_X1 U15089 ( .A1(n18469), .A2(n18244), .B1(n18183), .B2(n18467), .ZN(
        n18206) );
  NAND2_X1 U15090 ( .A1(n11734), .A2(n18255), .ZN(n18182) );
  INV_X1 U15091 ( .A(n18182), .ZN(n11737) );
  INV_X1 U15092 ( .A(n11735), .ZN(n11736) );
  NAND2_X1 U15093 ( .A1(n11737), .A2(n11736), .ZN(n11738) );
  NOR2_X4 U15094 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13875) );
  AOI22_X1 U15095 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11796), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11748) );
  AND2_X2 U15096 ( .A1(n13859), .A2(n13875), .ZN(n12549) );
  AOI22_X1 U15097 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9661), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11747) );
  AND2_X4 U15098 ( .A1(n11750), .A2(n11749), .ZN(n12450) );
  AOI22_X1 U15099 ( .A1(n12450), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11746) );
  AOI22_X1 U15100 ( .A1(n9723), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11745) );
  AND2_X2 U15101 ( .A1(n13859), .A2(n11751), .ZN(n12378) );
  AOI22_X1 U15102 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11804), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11756) );
  AND2_X2 U15103 ( .A1(n11749), .A2(n13859), .ZN(n11859) );
  AOI22_X1 U15104 ( .A1(n11866), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11859), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11755) );
  AOI22_X1 U15105 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11754) );
  AOI22_X1 U15106 ( .A1(n11774), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11753) );
  AOI22_X1 U15107 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11859), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11761) );
  AOI22_X1 U15108 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11804), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11760) );
  AOI22_X1 U15109 ( .A1(n9723), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9662), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U15110 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9719), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U15111 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12450), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11765) );
  AOI22_X1 U15112 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U15113 ( .A1(n11866), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11823), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U15114 ( .A1(n11774), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11762) );
  INV_X1 U15115 ( .A(n13321), .ZN(n11834) );
  NAND2_X1 U15116 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11769) );
  NAND2_X1 U15117 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11768) );
  NAND2_X1 U15118 ( .A1(n11861), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11767) );
  NAND2_X1 U15119 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11766) );
  NAND2_X1 U15120 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11773) );
  NAND2_X1 U15121 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11772) );
  NAND2_X1 U15122 ( .A1(n12450), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11771) );
  NAND2_X1 U15123 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11770) );
  NAND2_X1 U15124 ( .A1(n11774), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11778) );
  NAND2_X1 U15125 ( .A1(n11866), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11777) );
  NAND2_X1 U15126 ( .A1(n11796), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11776) );
  NAND2_X1 U15127 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11775) );
  NAND2_X1 U15128 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11782) );
  NAND2_X1 U15129 ( .A1(n11823), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11781) );
  NAND2_X1 U15130 ( .A1(n12509), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11780) );
  NAND2_X1 U15131 ( .A1(n12542), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11779) );
  AOI22_X1 U15132 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11790) );
  AOI22_X1 U15133 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11804), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11789) );
  AOI22_X1 U15134 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11796), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U15135 ( .A1(n11861), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U15136 ( .A1(n12509), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U15137 ( .A1(n11774), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12549), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U15138 ( .A1(n12450), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12527), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U15139 ( .A1(n9722), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9662), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11800) );
  AOI22_X1 U15140 ( .A1(n11774), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12549), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U15141 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11859), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U15142 ( .A1(n9719), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(n9661), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U15143 ( .A1(n9726), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11802) );
  AOI22_X1 U15144 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11801) );
  NAND2_X1 U15145 ( .A1(n11802), .A2(n11801), .ZN(n11808) );
  AOI22_X1 U15146 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12450), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11806) );
  AOI22_X1 U15147 ( .A1(n11866), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11804), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11805) );
  NAND2_X1 U15148 ( .A1(n11806), .A2(n11805), .ZN(n11807) );
  NAND2_X1 U15149 ( .A1(n11774), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11814) );
  NAND2_X1 U15150 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11813) );
  NAND2_X1 U15151 ( .A1(n9662), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11812) );
  NAND2_X1 U15152 ( .A1(n9723), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11811) );
  NAND2_X1 U15153 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11818) );
  NAND2_X1 U15154 ( .A1(n12450), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11817) );
  NAND2_X1 U15155 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11816) );
  NAND2_X1 U15156 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11815) );
  NAND2_X1 U15157 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11822) );
  NAND2_X1 U15158 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11821) );
  NAND2_X1 U15159 ( .A1(n11866), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11820) );
  NAND2_X1 U15160 ( .A1(n11861), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11819) );
  NAND2_X1 U15161 ( .A1(n11796), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11828) );
  NAND2_X1 U15162 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11827) );
  NAND2_X1 U15163 ( .A1(n11823), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11826) );
  NAND2_X1 U15164 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11825) );
  NOR2_X1 U15165 ( .A1(n11879), .A2(n9698), .ZN(n11833) );
  NAND2_X1 U15166 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11838) );
  NAND2_X1 U15167 ( .A1(n12450), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11837) );
  NAND2_X1 U15168 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11836) );
  NAND2_X1 U15169 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11835) );
  NAND2_X1 U15170 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11842) );
  NAND2_X1 U15171 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11841) );
  NAND2_X1 U15172 ( .A1(n11866), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11840) );
  NAND2_X1 U15173 ( .A1(n11861), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11839) );
  NAND2_X1 U15174 ( .A1(n11774), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11846) );
  NAND2_X1 U15175 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11845) );
  NAND2_X1 U15176 ( .A1(n12542), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11844) );
  NAND2_X1 U15177 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11850) );
  NAND2_X1 U15178 ( .A1(n9661), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11848) );
  NAND2_X1 U15179 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11847) );
  XNOR2_X1 U15180 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12746) );
  NAND2_X1 U15181 ( .A1(n12450), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11858) );
  NAND2_X1 U15182 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11857) );
  NAND2_X1 U15183 ( .A1(n11804), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11856) );
  NAND2_X1 U15184 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11855) );
  NAND2_X1 U15185 ( .A1(n11859), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11865) );
  NAND2_X1 U15186 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11864) );
  NAND2_X1 U15187 ( .A1(n11861), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11863) );
  NAND2_X1 U15188 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11862) );
  NAND2_X1 U15189 ( .A1(n11774), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11870) );
  NAND2_X1 U15190 ( .A1(n11866), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11869) );
  NAND2_X1 U15191 ( .A1(n11796), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11868) );
  NAND2_X1 U15192 ( .A1(n11824), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11867) );
  NAND2_X1 U15193 ( .A1(n11823), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11873) );
  NAND2_X1 U15194 ( .A1(n9723), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11872) );
  NAND2_X1 U15195 ( .A1(n12542), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11871) );
  NAND3_X1 U15196 ( .A1(n13865), .A2(n9660), .A3(n14148), .ZN(n13552) );
  NAND2_X1 U15197 ( .A1(n11877), .A2(n11879), .ZN(n13686) );
  NAND2_X1 U15198 ( .A1(n9717), .A2(n11876), .ZN(n11896) );
  NAND2_X1 U15199 ( .A1(n12636), .A2(n11879), .ZN(n11878) );
  INV_X1 U15200 ( .A(n11877), .ZN(n15052) );
  NAND2_X1 U15201 ( .A1(n11882), .A2(n11881), .ZN(n11883) );
  NAND2_X1 U15202 ( .A1(n11885), .A2(n11941), .ZN(n11886) );
  INV_X2 U15203 ( .A(n13675), .ZN(n14133) );
  NAND2_X1 U15204 ( .A1(n13551), .A2(n14857), .ZN(n11887) );
  NOR2_X1 U15205 ( .A1(n13658), .A2(n14106), .ZN(n11893) );
  NAND2_X1 U15206 ( .A1(n11885), .A2(n12739), .ZN(n12771) );
  NAND2_X1 U15207 ( .A1(n13678), .A2(n11889), .ZN(n11892) );
  NAND2_X1 U15208 ( .A1(n12771), .A2(n11892), .ZN(n13550) );
  NAND2_X1 U15209 ( .A1(n14148), .A2(n11879), .ZN(n12777) );
  AND2_X1 U15210 ( .A1(n12777), .A2(n14106), .ZN(n11895) );
  INV_X1 U15211 ( .A(n14093), .ZN(n11894) );
  NAND2_X1 U15212 ( .A1(n11895), .A2(n14091), .ZN(n13543) );
  NAND2_X1 U15213 ( .A1(n13543), .A2(n11897), .ZN(n11899) );
  NAND2_X1 U15214 ( .A1(n11941), .A2(n13675), .ZN(n14162) );
  INV_X1 U15215 ( .A(n13865), .ZN(n13545) );
  NAND3_X1 U15216 ( .A1(n11915), .A2(n11899), .A3(n11898), .ZN(n11902) );
  NAND2_X1 U15217 ( .A1(n11979), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11905) );
  NAND2_X1 U15218 ( .A1(n15498), .A2(n21023), .ZN(n13324) );
  MUX2_X1 U15219 ( .A(n13324), .B(n16248), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11904) );
  NAND2_X1 U15220 ( .A1(n11900), .A2(n9660), .ZN(n13549) );
  AND2_X1 U15221 ( .A1(n11906), .A2(n11891), .ZN(n11909) );
  INV_X1 U15222 ( .A(n9660), .ZN(n14160) );
  INV_X2 U15223 ( .A(n12739), .ZN(n12637) );
  NAND2_X1 U15224 ( .A1(n14160), .A2(n12637), .ZN(n14847) );
  AND2_X1 U15225 ( .A1(n12777), .A2(n11877), .ZN(n12775) );
  INV_X1 U15226 ( .A(n12775), .ZN(n11907) );
  INV_X1 U15227 ( .A(n13658), .ZN(n21019) );
  NAND2_X1 U15228 ( .A1(n11907), .A2(n21019), .ZN(n11908) );
  OAI21_X1 U15229 ( .B1(n11909), .B2(n14847), .A(n11908), .ZN(n11912) );
  NAND2_X1 U15230 ( .A1(n13865), .A2(n11910), .ZN(n12773) );
  NAND4_X1 U15231 ( .A1(n12773), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n15498), 
        .A4(n14162), .ZN(n11911) );
  NOR2_X1 U15232 ( .A1(n11912), .A2(n11911), .ZN(n11914) );
  NAND3_X1 U15233 ( .A1(n13543), .A2(n13675), .A3(n11897), .ZN(n11913) );
  NAND4_X1 U15234 ( .A1(n13549), .A2(n11915), .A3(n11914), .A4(n11913), .ZN(
        n11966) );
  INV_X1 U15235 ( .A(n11966), .ZN(n11916) );
  XNOR2_X2 U15236 ( .A(n11967), .B(n11916), .ZN(n12024) );
  NAND2_X1 U15237 ( .A1(n12024), .A2(n21023), .ZN(n11940) );
  AOI22_X1 U15238 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11920) );
  AOI22_X1 U15239 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U15240 ( .A1(n12450), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11918) );
  AOI22_X1 U15241 ( .A1(n11796), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11917) );
  NAND4_X1 U15242 ( .A1(n11920), .A2(n11919), .A3(n11918), .A4(n11917), .ZN(
        n11926) );
  AOI22_X1 U15243 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11924) );
  AOI22_X1 U15244 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12549), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11923) );
  AOI22_X1 U15245 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9661), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11922) );
  AOI22_X1 U15246 ( .A1(n9723), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9662), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11921) );
  NAND4_X1 U15247 ( .A1(n11924), .A2(n11923), .A3(n11922), .A4(n11921), .ZN(
        n11925) );
  INV_X1 U15248 ( .A(n13300), .ZN(n11927) );
  NOR2_X1 U15249 ( .A1(n11927), .A2(n12041), .ZN(n11944) );
  NOR2_X1 U15250 ( .A1(n12041), .A2(n13300), .ZN(n11946) );
  AOI22_X1 U15251 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11931) );
  AOI22_X1 U15252 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11930) );
  AOI22_X1 U15253 ( .A1(n12509), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11929) );
  AOI22_X1 U15254 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11823), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11928) );
  NAND4_X1 U15255 ( .A1(n11931), .A2(n11930), .A3(n11929), .A4(n11928), .ZN(
        n11937) );
  AOI22_X1 U15256 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11935) );
  AOI22_X1 U15257 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U15258 ( .A1(n11866), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9719), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U15259 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11932) );
  NAND4_X1 U15260 ( .A1(n11935), .A2(n11934), .A3(n11933), .A4(n11932), .ZN(
        n11936) );
  MUX2_X1 U15261 ( .A(n11944), .B(n11946), .S(n13238), .Z(n11938) );
  NAND2_X2 U15262 ( .A1(n11940), .A2(n11939), .ZN(n12022) );
  INV_X1 U15263 ( .A(n12619), .ZN(n12613) );
  INV_X1 U15264 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20481) );
  AOI21_X1 U15265 ( .B1(n14106), .B2(n13300), .A(n21023), .ZN(n11943) );
  NAND2_X1 U15266 ( .A1(n11941), .A2(n13238), .ZN(n11942) );
  NAND2_X1 U15267 ( .A1(n12022), .A2(n12021), .ZN(n11945) );
  INV_X1 U15268 ( .A(n11944), .ZN(n13296) );
  INV_X1 U15269 ( .A(n11946), .ZN(n11960) );
  NAND2_X1 U15270 ( .A1(n12619), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11959) );
  AOI22_X1 U15271 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U15272 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12450), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U15274 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U15275 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11947) );
  NAND4_X1 U15276 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n11956) );
  AOI22_X1 U15277 ( .A1(n12527), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U15278 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9661), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U15279 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9866), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U15280 ( .A1(n9723), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9662), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11951) );
  NAND4_X1 U15281 ( .A1(n11954), .A2(n11953), .A3(n11952), .A4(n11951), .ZN(
        n11955) );
  INV_X1 U15282 ( .A(n13239), .ZN(n11957) );
  OR2_X1 U15283 ( .A1(n12042), .A2(n11957), .ZN(n11958) );
  NAND2_X1 U15285 ( .A1(n11979), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11963) );
  NAND2_X1 U15286 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11982) );
  OAI21_X1 U15287 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11982), .ZN(n20769) );
  OR2_X1 U15288 ( .A1(n16248), .A2(n20532), .ZN(n11976) );
  OAI21_X1 U15289 ( .B1(n13324), .B2(n20769), .A(n11976), .ZN(n11961) );
  INV_X1 U15290 ( .A(n11961), .ZN(n11962) );
  NAND2_X1 U15291 ( .A1(n11963), .A2(n11962), .ZN(n11965) );
  NAND2_X1 U15292 ( .A1(n11967), .A2(n11966), .ZN(n11968) );
  NAND2_X1 U15293 ( .A1(n14099), .A2(n11968), .ZN(n20503) );
  NAND2_X1 U15294 ( .A1(n11990), .A2(n20503), .ZN(n14391) );
  INV_X1 U15295 ( .A(n12041), .ZN(n11969) );
  NAND2_X1 U15296 ( .A1(n11969), .A2(n13239), .ZN(n11970) );
  INV_X1 U15298 ( .A(n11973), .ZN(n11974) );
  NAND2_X1 U15300 ( .A1(n11976), .A2(n11742), .ZN(n11977) );
  NAND2_X1 U15301 ( .A1(n11978), .A2(n11977), .ZN(n11988) );
  NAND2_X1 U15302 ( .A1(n11990), .A2(n11988), .ZN(n11986) );
  NOR2_X1 U15303 ( .A1(n16248), .A2(n16225), .ZN(n11980) );
  INV_X1 U15304 ( .A(n13324), .ZN(n11984) );
  INV_X1 U15305 ( .A(n11982), .ZN(n11981) );
  NAND2_X1 U15306 ( .A1(n11981), .A2(n16225), .ZN(n20569) );
  NAND2_X1 U15307 ( .A1(n11982), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11983) );
  NAND2_X1 U15308 ( .A1(n20569), .A2(n11983), .ZN(n14396) );
  NAND2_X1 U15309 ( .A1(n11984), .A2(n14396), .ZN(n11987) );
  NAND2_X1 U15310 ( .A1(n11989), .A2(n11987), .ZN(n11985) );
  NAND4_X1 U15311 ( .A1(n11990), .A2(n11989), .A3(n11988), .A4(n11987), .ZN(
        n11991) );
  AOI22_X1 U15312 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11995) );
  AOI22_X1 U15313 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U15314 ( .A1(n9726), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U15315 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11992) );
  NAND4_X1 U15316 ( .A1(n11995), .A2(n11994), .A3(n11993), .A4(n11992), .ZN(
        n12001) );
  AOI22_X1 U15317 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12507), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11999) );
  AOI22_X1 U15318 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U15319 ( .A1(n9722), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9662), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11997) );
  INV_X1 U15320 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n20487) );
  AOI22_X1 U15321 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11996) );
  NAND4_X1 U15322 ( .A1(n11999), .A2(n11998), .A3(n11997), .A4(n11996), .ZN(
        n12000) );
  AOI22_X1 U15323 ( .A1(n12003), .A2(n12002), .B1(n12619), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12004) );
  INV_X2 U15324 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n12006) );
  INV_X1 U15325 ( .A(n13686), .ZN(n14094) );
  NAND2_X1 U15326 ( .A1(n14094), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12082) );
  XNOR2_X1 U15327 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14164) );
  AOI21_X1 U15328 ( .B1(n12537), .B2(n14164), .A(n12566), .ZN(n12008) );
  NAND2_X1 U15329 ( .A1(n12567), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n12007) );
  OAI211_X1 U15330 ( .C1(n12082), .C2(n11740), .A(n12008), .B(n12007), .ZN(
        n12009) );
  INV_X1 U15331 ( .A(n12009), .ZN(n12010) );
  NAND2_X1 U15332 ( .A1(n12566), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12032) );
  INV_X1 U15333 ( .A(n13824), .ZN(n12031) );
  INV_X1 U15334 ( .A(n12011), .ZN(n12012) );
  NAND2_X2 U15335 ( .A1(n12015), .A2(n12014), .ZN(n15489) );
  NAND2_X1 U15336 ( .A1(n15489), .A2(n12247), .ZN(n12020) );
  AOI22_X1 U15337 ( .A1(n12567), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n12006), .ZN(n12018) );
  INV_X1 U15338 ( .A(n12082), .ZN(n12016) );
  NAND2_X1 U15339 ( .A1(n12016), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12017) );
  AND2_X1 U15340 ( .A1(n12018), .A2(n12017), .ZN(n12019) );
  NAND2_X1 U15341 ( .A1(n12020), .A2(n12019), .ZN(n13650) );
  XNOR2_X2 U15342 ( .A(n12022), .B(n12021), .ZN(n13236) );
  NAND2_X1 U15343 ( .A1(n13236), .A2(n11910), .ZN(n12023) );
  NAND2_X1 U15344 ( .A1(n12023), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13712) );
  NAND2_X1 U15345 ( .A1(n12006), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12026) );
  NAND2_X1 U15346 ( .A1(n12104), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12025) );
  OAI211_X1 U15347 ( .C1(n12082), .C2(n11741), .A(n12026), .B(n12025), .ZN(
        n12027) );
  AOI21_X1 U15348 ( .B1(n12024), .B2(n12247), .A(n12027), .ZN(n12028) );
  OR2_X1 U15349 ( .A1(n13712), .A2(n12028), .ZN(n13713) );
  INV_X1 U15350 ( .A(n12028), .ZN(n13714) );
  OR2_X1 U15351 ( .A1(n13714), .A2(n12631), .ZN(n12029) );
  NAND2_X1 U15352 ( .A1(n13713), .A2(n12029), .ZN(n13649) );
  NAND2_X1 U15353 ( .A1(n13650), .A2(n13649), .ZN(n13825) );
  NAND2_X1 U15354 ( .A1(n12031), .A2(n12030), .ZN(n13826) );
  INV_X1 U15355 ( .A(n12033), .ZN(n12035) );
  NAND2_X1 U15356 ( .A1(n12035), .A2(n12034), .ZN(n12055) );
  NAND2_X1 U15357 ( .A1(n11979), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12040) );
  NAND3_X1 U15358 ( .A1(n20768), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20676) );
  INV_X1 U15359 ( .A(n20676), .ZN(n14109) );
  NAND2_X1 U15360 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14109), .ZN(
        n14107) );
  NAND2_X1 U15361 ( .A1(n20768), .A2(n14107), .ZN(n12037) );
  NOR3_X1 U15362 ( .A1(n20768), .A2(n16225), .A3(n20532), .ZN(n20887) );
  NAND2_X1 U15363 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20887), .ZN(
        n20875) );
  NAND2_X1 U15364 ( .A1(n12037), .A2(n20875), .ZN(n14497) );
  OAI22_X1 U15365 ( .A1(n13324), .A2(n14497), .B1(n16248), .B2(n20768), .ZN(
        n12038) );
  INV_X1 U15366 ( .A(n12038), .ZN(n12039) );
  NAND2_X1 U15367 ( .A1(n13856), .A2(n21023), .ZN(n12054) );
  AOI22_X1 U15368 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U15369 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U15370 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12044) );
  AOI22_X1 U15371 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12043) );
  NAND4_X1 U15372 ( .A1(n12046), .A2(n12045), .A3(n12044), .A4(n12043), .ZN(
        n12052) );
  AOI22_X1 U15373 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12549), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15374 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15375 ( .A1(n12509), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12048) );
  AOI22_X1 U15376 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12047) );
  NAND4_X1 U15377 ( .A1(n12050), .A2(n12049), .A3(n12048), .A4(n12047), .ZN(
        n12051) );
  AOI22_X1 U15378 ( .A1(n12596), .A2(n13270), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12619), .ZN(n12053) );
  NAND2_X1 U15379 ( .A1(n12055), .A2(n13954), .ZN(n12056) );
  NAND2_X1 U15380 ( .A1(n12079), .A2(n12056), .ZN(n13254) );
  INV_X1 U15381 ( .A(n12247), .ZN(n12264) );
  INV_X1 U15382 ( .A(n12059), .ZN(n12058) );
  INV_X1 U15383 ( .A(n12084), .ZN(n12062) );
  INV_X1 U15384 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12060) );
  NAND2_X1 U15385 ( .A1(n12060), .A2(n12059), .ZN(n12061) );
  NAND2_X1 U15386 ( .A1(n12062), .A2(n12061), .ZN(n20322) );
  AOI22_X1 U15387 ( .A1(n20322), .A2(n12560), .B1(n12566), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12064) );
  NAND2_X1 U15388 ( .A1(n12567), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12063) );
  OAI211_X1 U15389 ( .C1(n12082), .C2(n12057), .A(n12064), .B(n12063), .ZN(
        n12065) );
  INV_X1 U15390 ( .A(n12065), .ZN(n12066) );
  OAI21_X2 U15391 ( .B1(n13254), .B2(n12264), .A(n12066), .ZN(n13902) );
  NAND2_X1 U15392 ( .A1(n13901), .A2(n13902), .ZN(n14067) );
  INV_X1 U15393 ( .A(n14067), .ZN(n12089) );
  AOI22_X1 U15394 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12396), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U15395 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15396 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12383), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15397 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12067) );
  NAND4_X1 U15398 ( .A1(n12070), .A2(n12069), .A3(n12068), .A4(n12067), .ZN(
        n12076) );
  AOI22_X1 U15399 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12235), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12074) );
  AOI22_X1 U15400 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12073) );
  AOI22_X1 U15401 ( .A1(n9723), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U15402 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12071) );
  NAND4_X1 U15403 ( .A1(n12074), .A2(n12073), .A3(n12072), .A4(n12071), .ZN(
        n12075) );
  NAND2_X1 U15404 ( .A1(n12596), .A2(n13269), .ZN(n12078) );
  NAND2_X1 U15405 ( .A1(n12619), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12077) );
  NAND2_X1 U15406 ( .A1(n12078), .A2(n12077), .ZN(n12090) );
  XNOR2_X1 U15407 ( .A(n12079), .B(n12090), .ZN(n13260) );
  NAND2_X1 U15408 ( .A1(n12006), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12081) );
  NAND2_X1 U15409 ( .A1(n12567), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12080) );
  OAI211_X1 U15410 ( .C1(n12082), .C2(n16459), .A(n12081), .B(n12080), .ZN(
        n12083) );
  NAND2_X1 U15411 ( .A1(n12083), .A2(n12631), .ZN(n12086) );
  OAI21_X1 U15412 ( .B1(n12084), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n12105), .ZN(n20426) );
  NAND2_X1 U15413 ( .A1(n20426), .A2(n12560), .ZN(n12085) );
  NAND2_X1 U15414 ( .A1(n12086), .A2(n12085), .ZN(n12087) );
  AOI21_X1 U15415 ( .B1(n13260), .B2(n12247), .A(n12087), .ZN(n14068) );
  NAND2_X1 U15416 ( .A1(n12089), .A2(n12088), .ZN(n13980) );
  NAND2_X1 U15417 ( .A1(n12091), .A2(n12090), .ZN(n12111) );
  AOI22_X1 U15418 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12095) );
  AOI22_X1 U15419 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12094) );
  AOI22_X1 U15420 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U15421 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12092) );
  NAND4_X1 U15422 ( .A1(n12095), .A2(n12094), .A3(n12093), .A4(n12092), .ZN(
        n12101) );
  AOI22_X1 U15423 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12507), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12099) );
  AOI22_X1 U15424 ( .A1(n9722), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12097) );
  INV_X1 U15425 ( .A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n20493) );
  AOI22_X1 U15426 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12096) );
  NAND4_X1 U15427 ( .A1(n12099), .A2(n12098), .A3(n12097), .A4(n12096), .ZN(
        n12100) );
  NAND2_X1 U15428 ( .A1(n12596), .A2(n13279), .ZN(n12103) );
  NAND2_X1 U15429 ( .A1(n12619), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12102) );
  NAND2_X1 U15430 ( .A1(n12103), .A2(n12102), .ZN(n12112) );
  XNOR2_X1 U15431 ( .A(n12111), .B(n12112), .ZN(n13267) );
  INV_X1 U15432 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n14095) );
  AND2_X1 U15433 ( .A1(n12105), .A2(n12107), .ZN(n12106) );
  OR2_X1 U15434 ( .A1(n12106), .A2(n12123), .ZN(n20293) );
  INV_X1 U15435 ( .A(n12566), .ZN(n12171) );
  NOR2_X1 U15436 ( .A1(n12171), .A2(n12107), .ZN(n12108) );
  AOI21_X1 U15437 ( .B1(n20293), .B2(n12560), .A(n12108), .ZN(n12109) );
  OAI21_X1 U15438 ( .B1(n12127), .B2(n14095), .A(n12109), .ZN(n12110) );
  AOI21_X1 U15439 ( .B1(n13267), .B2(n12247), .A(n12110), .ZN(n13981) );
  INV_X1 U15440 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20363) );
  AOI22_X1 U15441 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12116) );
  AOI22_X1 U15442 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12115) );
  AOI22_X1 U15443 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12114) );
  AOI22_X1 U15444 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9866), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12113) );
  NAND4_X1 U15445 ( .A1(n12116), .A2(n12115), .A3(n12114), .A4(n12113), .ZN(
        n12122) );
  AOI22_X1 U15446 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12120) );
  AOI22_X1 U15447 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12507), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15448 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12118) );
  AOI22_X1 U15449 ( .A1(n9723), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9662), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12117) );
  NAND4_X1 U15450 ( .A1(n12120), .A2(n12119), .A3(n12118), .A4(n12117), .ZN(
        n12121) );
  AOI22_X1 U15451 ( .A1(n12596), .A2(n13287), .B1(n12619), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12129) );
  NAND2_X1 U15452 ( .A1(n12128), .A2(n12129), .ZN(n13278) );
  NAND2_X1 U15453 ( .A1(n13278), .A2(n12247), .ZN(n12126) );
  NOR2_X1 U15454 ( .A1(n12123), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12124) );
  OR2_X1 U15455 ( .A1(n12134), .A2(n12124), .ZN(n20281) );
  AOI22_X1 U15456 ( .A1(n20281), .A2(n12560), .B1(n12566), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12125) );
  NAND2_X1 U15457 ( .A1(n13979), .A2(n14281), .ZN(n14280) );
  INV_X1 U15458 ( .A(n14280), .ZN(n12188) );
  NAND2_X1 U15459 ( .A1(n12596), .A2(n13300), .ZN(n12132) );
  NAND2_X1 U15460 ( .A1(n12619), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12131) );
  NAND2_X1 U15461 ( .A1(n12132), .A2(n12131), .ZN(n12133) );
  INV_X1 U15462 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12137) );
  OR2_X1 U15463 ( .A1(n12134), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12135) );
  NAND2_X1 U15464 ( .A1(n12135), .A2(n12170), .ZN(n20269) );
  AOI22_X1 U15465 ( .A1(n20269), .A2(n12560), .B1(n12566), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12136) );
  OAI21_X1 U15466 ( .B1(n12127), .B2(n12137), .A(n12136), .ZN(n12138) );
  AOI21_X1 U15467 ( .B1(n13292), .B2(n12247), .A(n12138), .ZN(n14357) );
  INV_X1 U15468 ( .A(n14357), .ZN(n12187) );
  XNOR2_X1 U15469 ( .A(n12189), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15280) );
  AOI22_X1 U15470 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12143) );
  BUF_X1 U15471 ( .A(n11803), .Z(n12407) );
  AOI22_X1 U15472 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12142) );
  AOI22_X1 U15473 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15474 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12140) );
  NAND4_X1 U15475 ( .A1(n12143), .A2(n12142), .A3(n12141), .A4(n12140), .ZN(
        n12149) );
  AOI22_X1 U15476 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12147) );
  AOI22_X1 U15477 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15478 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9866), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U15479 ( .A1(n9722), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12144) );
  NAND4_X1 U15480 ( .A1(n12147), .A2(n12146), .A3(n12145), .A4(n12144), .ZN(
        n12148) );
  NOR2_X1 U15481 ( .A1(n12149), .A2(n12148), .ZN(n12152) );
  NAND2_X1 U15482 ( .A1(n12567), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12151) );
  NAND2_X1 U15483 ( .A1(n12566), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12150) );
  OAI211_X1 U15484 ( .C1(n12264), .C2(n12152), .A(n12151), .B(n12150), .ZN(
        n12153) );
  AOI21_X1 U15485 ( .B1(n15280), .B2(n12560), .A(n12153), .ZN(n14556) );
  XOR2_X1 U15486 ( .A(n20260), .B(n12154), .Z(n20258) );
  INV_X1 U15487 ( .A(n20258), .ZN(n12169) );
  AOI22_X1 U15488 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15489 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U15490 ( .A1(n12509), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U15491 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12155) );
  NAND4_X1 U15492 ( .A1(n12158), .A2(n12157), .A3(n12156), .A4(n12155), .ZN(
        n12164) );
  AOI22_X1 U15493 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15494 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U15495 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9866), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U15496 ( .A1(n12467), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12159) );
  NAND4_X1 U15497 ( .A1(n12162), .A2(n12161), .A3(n12160), .A4(n12159), .ZN(
        n12163) );
  NOR2_X1 U15498 ( .A1(n12164), .A2(n12163), .ZN(n12167) );
  NAND2_X1 U15499 ( .A1(n12567), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12166) );
  NAND2_X1 U15500 ( .A1(n12566), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12165) );
  OAI211_X1 U15501 ( .C1(n12264), .C2(n12167), .A(n12166), .B(n12165), .ZN(
        n12168) );
  AOI21_X1 U15502 ( .B1(n12169), .B2(n12560), .A(n12168), .ZN(n14426) );
  OR2_X1 U15503 ( .A1(n14556), .A2(n14426), .ZN(n12185) );
  XNOR2_X1 U15504 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12170), .ZN(
        n14482) );
  INV_X1 U15505 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n14480) );
  OAI22_X1 U15506 ( .A1(n12631), .A2(n14482), .B1(n12171), .B2(n14480), .ZN(
        n12172) );
  AOI21_X1 U15507 ( .B1(n12567), .B2(P1_EAX_REG_8__SCAN_IN), .A(n12172), .ZN(
        n12184) );
  AOI22_X1 U15508 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U15509 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12175) );
  AOI22_X1 U15510 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9866), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12174) );
  AOI22_X1 U15511 ( .A1(n9723), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n9662), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12173) );
  NAND4_X1 U15512 ( .A1(n12176), .A2(n12175), .A3(n12174), .A4(n12173), .ZN(
        n12182) );
  AOI22_X1 U15513 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11803), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15514 ( .A1(n12450), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15515 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15516 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12177) );
  NAND4_X1 U15517 ( .A1(n12180), .A2(n12179), .A3(n12178), .A4(n12177), .ZN(
        n12181) );
  OAI21_X1 U15518 ( .B1(n12182), .B2(n12181), .A(n12247), .ZN(n12183) );
  NOR2_X1 U15519 ( .A1(n12185), .A2(n14405), .ZN(n12186) );
  NAND2_X1 U15520 ( .A1(n12567), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n12192) );
  OAI21_X1 U15521 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12190), .A(
        n12218), .ZN(n16367) );
  AOI22_X1 U15522 ( .A1(n12537), .A2(n16367), .B1(n12566), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12191) );
  NAND2_X1 U15523 ( .A1(n12192), .A2(n12191), .ZN(n14487) );
  AOI22_X1 U15524 ( .A1(n12450), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U15525 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15526 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12507), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15527 ( .A1(n9722), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(n9662), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12193) );
  NAND4_X1 U15528 ( .A1(n12196), .A2(n12195), .A3(n12194), .A4(n12193), .ZN(
        n12202) );
  AOI22_X1 U15529 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12200) );
  AOI22_X1 U15530 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15531 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9866), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15532 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12197) );
  NAND4_X1 U15533 ( .A1(n12200), .A2(n12199), .A3(n12198), .A4(n12197), .ZN(
        n12201) );
  OR2_X1 U15534 ( .A1(n12202), .A2(n12201), .ZN(n12203) );
  NAND2_X1 U15535 ( .A1(n12247), .A2(n12203), .ZN(n14549) );
  INV_X1 U15536 ( .A(n14549), .ZN(n12204) );
  INV_X1 U15537 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14530) );
  AOI22_X1 U15538 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15539 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12507), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15540 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9866), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15541 ( .A1(n9723), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9662), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12205) );
  NAND4_X1 U15542 ( .A1(n12208), .A2(n12207), .A3(n12206), .A4(n12205), .ZN(
        n12214) );
  AOI22_X1 U15543 ( .A1(n12450), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15544 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U15545 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15546 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12209) );
  NAND4_X1 U15547 ( .A1(n12212), .A2(n12211), .A3(n12210), .A4(n12209), .ZN(
        n12213) );
  OAI21_X1 U15548 ( .B1(n12214), .B2(n12213), .A(n12247), .ZN(n12217) );
  INV_X1 U15549 ( .A(n12234), .ZN(n12215) );
  XNOR2_X1 U15550 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12215), .ZN(
        n16317) );
  AOI22_X1 U15551 ( .A1(n12537), .A2(n16317), .B1(n12566), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12216) );
  OAI211_X1 U15552 ( .C1(n12127), .C2(n14530), .A(n12217), .B(n12216), .ZN(
        n14524) );
  INV_X1 U15553 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14491) );
  INV_X1 U15554 ( .A(n12218), .ZN(n12219) );
  XNOR2_X1 U15555 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12219), .ZN(
        n16331) );
  AOI22_X1 U15556 ( .A1(n12537), .A2(n16331), .B1(n12566), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U15557 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12235), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15558 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15559 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12383), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15560 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12220) );
  NAND4_X1 U15561 ( .A1(n12223), .A2(n12222), .A3(n12221), .A4(n12220), .ZN(
        n12230) );
  AOI22_X1 U15562 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12548), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15563 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15564 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12526), .B1(
        n9866), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15565 ( .A1(n9723), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(n9662), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12225) );
  NAND4_X1 U15566 ( .A1(n12228), .A2(n12227), .A3(n12226), .A4(n12225), .ZN(
        n12229) );
  OR2_X1 U15567 ( .A1(n12230), .A2(n12229), .ZN(n12231) );
  NAND2_X1 U15568 ( .A1(n12247), .A2(n12231), .ZN(n12232) );
  OAI211_X1 U15569 ( .C1(n12127), .C2(n14491), .A(n12233), .B(n12232), .ZN(
        n14489) );
  XOR2_X1 U15570 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n12250), .Z(
        n16354) );
  AOI22_X1 U15571 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12383), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U15572 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12407), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12238) );
  AOI22_X1 U15573 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U15574 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12236) );
  NAND4_X1 U15575 ( .A1(n12239), .A2(n12238), .A3(n12237), .A4(n12236), .ZN(
        n12245) );
  AOI22_X1 U15576 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12243) );
  AOI22_X1 U15577 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12242) );
  AOI22_X1 U15578 ( .A1(n9722), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U15579 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12240) );
  NAND4_X1 U15580 ( .A1(n12243), .A2(n12242), .A3(n12241), .A4(n12240), .ZN(
        n12244) );
  OR2_X1 U15581 ( .A1(n12245), .A2(n12244), .ZN(n12246) );
  AOI22_X1 U15582 ( .A1(n12247), .A2(n12246), .B1(n12566), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12249) );
  NAND2_X1 U15583 ( .A1(n12567), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12248) );
  OAI211_X1 U15584 ( .C1(n16354), .C2(n12631), .A(n12249), .B(n12248), .ZN(
        n14571) );
  XNOR2_X1 U15585 ( .A(n12281), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16306) );
  AOI22_X1 U15586 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U15587 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15588 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15589 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12251) );
  NAND4_X1 U15590 ( .A1(n12254), .A2(n12253), .A3(n12252), .A4(n12251), .ZN(
        n12260) );
  AOI22_X1 U15591 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12258) );
  AOI22_X1 U15592 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12257) );
  AOI22_X1 U15593 ( .A1(n9722), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9662), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12255) );
  NAND4_X1 U15594 ( .A1(n12258), .A2(n12257), .A3(n12256), .A4(n12255), .ZN(
        n12259) );
  NOR2_X1 U15595 ( .A1(n12260), .A2(n12259), .ZN(n12263) );
  NAND2_X1 U15596 ( .A1(n12567), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12262) );
  NAND2_X1 U15597 ( .A1(n12566), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12261) );
  OAI211_X1 U15598 ( .C1(n12264), .C2(n12263), .A(n12262), .B(n12261), .ZN(
        n12265) );
  INV_X1 U15599 ( .A(n12265), .ZN(n12266) );
  OAI21_X1 U15600 ( .B1(n16306), .B2(n12631), .A(n12266), .ZN(n14584) );
  NAND2_X1 U15601 ( .A1(n14572), .A2(n14584), .ZN(n14583) );
  AOI22_X1 U15602 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12270) );
  AOI22_X1 U15603 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12269) );
  AOI22_X1 U15604 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12268) );
  AOI22_X1 U15605 ( .A1(n12508), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12267) );
  NAND4_X1 U15606 ( .A1(n12270), .A2(n12269), .A3(n12268), .A4(n12267), .ZN(
        n12276) );
  AOI22_X1 U15607 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15608 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12507), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15609 ( .A1(n9723), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12271) );
  NAND4_X1 U15610 ( .A1(n12274), .A2(n12273), .A3(n12272), .A4(n12271), .ZN(
        n12275) );
  NOR2_X1 U15611 ( .A1(n12276), .A2(n12275), .ZN(n12280) );
  NAND2_X1 U15612 ( .A1(n12006), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12277) );
  NAND2_X1 U15613 ( .A1(n12631), .A2(n12277), .ZN(n12278) );
  AOI21_X1 U15614 ( .B1(n12567), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12278), .ZN(
        n12279) );
  OAI21_X1 U15615 ( .B1(n12563), .B2(n12280), .A(n12279), .ZN(n12284) );
  OAI21_X1 U15616 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12282), .A(
        n12313), .ZN(n16353) );
  OR2_X1 U15617 ( .A1(n16353), .A2(n12631), .ZN(n12283) );
  NAND2_X1 U15618 ( .A1(n12284), .A2(n12283), .ZN(n15041) );
  AOI22_X1 U15619 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15620 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12288) );
  AOI22_X1 U15621 ( .A1(n9722), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n9662), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12287) );
  NAND4_X1 U15622 ( .A1(n12289), .A2(n12288), .A3(n12287), .A4(n12286), .ZN(
        n12295) );
  AOI22_X1 U15623 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15624 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U15625 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U15626 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12290) );
  NAND4_X1 U15627 ( .A1(n12293), .A2(n12292), .A3(n12291), .A4(n12290), .ZN(
        n12294) );
  OR2_X1 U15628 ( .A1(n12295), .A2(n12294), .ZN(n12298) );
  INV_X1 U15629 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n15107) );
  INV_X1 U15630 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15010) );
  XNOR2_X1 U15631 ( .A(n12313), .B(n15010), .ZN(n15240) );
  AOI22_X1 U15632 ( .A1(n15240), .A2(n12560), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n12566), .ZN(n12296) );
  OAI21_X1 U15633 ( .B1(n12127), .B2(n15107), .A(n12296), .ZN(n12297) );
  AOI21_X1 U15634 ( .B1(n12534), .B2(n12298), .A(n12297), .ZN(n15005) );
  AOI22_X1 U15635 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U15636 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12301) );
  AOI22_X1 U15637 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12300) );
  AOI22_X1 U15638 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12299) );
  NAND4_X1 U15639 ( .A1(n12302), .A2(n12301), .A3(n12300), .A4(n12299), .ZN(
        n12308) );
  AOI22_X1 U15640 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12306) );
  AOI22_X1 U15641 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12507), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12305) );
  AOI22_X1 U15642 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9866), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U15643 ( .A1(n9722), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12303) );
  NAND4_X1 U15644 ( .A1(n12306), .A2(n12305), .A3(n12304), .A4(n12303), .ZN(
        n12307) );
  NOR2_X1 U15645 ( .A1(n12308), .A2(n12307), .ZN(n12312) );
  OAI21_X1 U15646 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n21170), .A(
        n12006), .ZN(n12309) );
  INV_X1 U15647 ( .A(n12309), .ZN(n12310) );
  AOI21_X1 U15648 ( .B1(n12567), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12310), .ZN(
        n12311) );
  OAI21_X1 U15649 ( .B1(n12563), .B2(n12312), .A(n12311), .ZN(n12319) );
  INV_X1 U15650 ( .A(n12315), .ZN(n12316) );
  INV_X1 U15651 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15226) );
  NAND2_X1 U15652 ( .A1(n12316), .A2(n15226), .ZN(n12317) );
  AND2_X1 U15653 ( .A1(n12351), .A2(n12317), .ZN(n16281) );
  NAND2_X1 U15654 ( .A1(n16281), .A2(n12560), .ZN(n12318) );
  NAND2_X1 U15655 ( .A1(n12319), .A2(n12318), .ZN(n15031) );
  AOI22_X1 U15656 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12324) );
  AOI22_X1 U15657 ( .A1(n12450), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12323) );
  AOI22_X1 U15658 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12322) );
  AOI22_X1 U15659 ( .A1(n12508), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12321) );
  NAND4_X1 U15660 ( .A1(n12324), .A2(n12323), .A3(n12322), .A4(n12321), .ZN(
        n12330) );
  AOI22_X1 U15661 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U15662 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12507), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15663 ( .A1(n12509), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9662), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12325) );
  NAND4_X1 U15664 ( .A1(n12328), .A2(n12327), .A3(n12326), .A4(n12325), .ZN(
        n12329) );
  NOR2_X1 U15665 ( .A1(n12330), .A2(n12329), .ZN(n12334) );
  NAND2_X1 U15666 ( .A1(n12006), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12331) );
  NAND2_X1 U15667 ( .A1(n12631), .A2(n12331), .ZN(n12332) );
  AOI21_X1 U15668 ( .B1(n12104), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12332), .ZN(
        n12333) );
  OAI21_X1 U15669 ( .B1(n12563), .B2(n12334), .A(n12333), .ZN(n12336) );
  XNOR2_X1 U15670 ( .A(n12351), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15222) );
  NAND2_X1 U15671 ( .A1(n15222), .A2(n12560), .ZN(n12335) );
  NAND2_X1 U15672 ( .A1(n14986), .A2(n14987), .ZN(n14968) );
  AOI22_X1 U15673 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12340) );
  AOI22_X1 U15674 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12224), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U15675 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12507), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12338) );
  AOI22_X1 U15676 ( .A1(n9723), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n9662), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12337) );
  NAND4_X1 U15677 ( .A1(n12340), .A2(n12339), .A3(n12338), .A4(n12337), .ZN(
        n12346) );
  AOI22_X1 U15678 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12383), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12344) );
  AOI22_X1 U15679 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12343) );
  AOI22_X1 U15680 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12342) );
  AOI22_X1 U15681 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12341) );
  NAND4_X1 U15682 ( .A1(n12344), .A2(n12343), .A3(n12342), .A4(n12341), .ZN(
        n12345) );
  NOR2_X1 U15683 ( .A1(n12346), .A2(n12345), .ZN(n12350) );
  NAND2_X1 U15684 ( .A1(n12006), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12347) );
  NAND2_X1 U15685 ( .A1(n12631), .A2(n12347), .ZN(n12348) );
  AOI21_X1 U15686 ( .B1(n12104), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12348), .ZN(
        n12349) );
  OAI21_X1 U15687 ( .B1(n12563), .B2(n12350), .A(n12349), .ZN(n12356) );
  NAND2_X1 U15688 ( .A1(n12353), .A2(n14978), .ZN(n12354) );
  NAND2_X1 U15689 ( .A1(n12374), .A2(n12354), .ZN(n15209) );
  NAND2_X1 U15690 ( .A1(n12356), .A2(n12355), .ZN(n14970) );
  NOR2_X2 U15691 ( .A1(n14968), .A2(n14970), .ZN(n14953) );
  AOI22_X1 U15692 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15693 ( .A1(n12407), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12359) );
  AOI22_X1 U15694 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15695 ( .A1(n12508), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12357) );
  NAND4_X1 U15696 ( .A1(n12360), .A2(n12359), .A3(n12358), .A4(n12357), .ZN(
        n12366) );
  AOI22_X1 U15697 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12364) );
  AOI22_X1 U15698 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12507), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U15699 ( .A1(n12509), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9662), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12361) );
  NAND4_X1 U15700 ( .A1(n12364), .A2(n12363), .A3(n12362), .A4(n12361), .ZN(
        n12365) );
  NOR2_X1 U15701 ( .A1(n12366), .A2(n12365), .ZN(n12370) );
  NAND2_X1 U15702 ( .A1(n12006), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12367) );
  NAND2_X1 U15703 ( .A1(n12631), .A2(n12367), .ZN(n12368) );
  AOI21_X1 U15704 ( .B1(n12104), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12368), .ZN(
        n12369) );
  OAI21_X1 U15705 ( .B1(n12563), .B2(n12370), .A(n12369), .ZN(n12372) );
  XNOR2_X1 U15706 ( .A(n12374), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15202) );
  NAND2_X1 U15707 ( .A1(n15202), .A2(n12560), .ZN(n12371) );
  NAND2_X1 U15708 ( .A1(n12372), .A2(n12371), .ZN(n14954) );
  INV_X1 U15709 ( .A(n12376), .ZN(n12377) );
  INV_X1 U15710 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14945) );
  OAI21_X1 U15711 ( .B1(n12377), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n12422), .ZN(n15190) );
  INV_X1 U15712 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n12393) );
  AOI22_X1 U15713 ( .A1(n12450), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U15714 ( .A1(n12378), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15715 ( .A1(n9722), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12380) );
  NAND4_X1 U15716 ( .A1(n12382), .A2(n12381), .A3(n12380), .A4(n12379), .ZN(
        n12390) );
  AOI22_X1 U15717 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12407), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12388) );
  AOI22_X1 U15718 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12387) );
  AOI22_X1 U15719 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U15720 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12385) );
  NAND4_X1 U15721 ( .A1(n12388), .A2(n12387), .A3(n12386), .A4(n12385), .ZN(
        n12389) );
  OAI21_X1 U15722 ( .B1(n12390), .B2(n12389), .A(n12534), .ZN(n12392) );
  AOI21_X1 U15723 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12006), .A(
        n12537), .ZN(n12391) );
  OAI211_X1 U15724 ( .C1(n12127), .C2(n12393), .A(n12392), .B(n12391), .ZN(
        n12394) );
  OAI21_X1 U15725 ( .B1(n12631), .B2(n15190), .A(n12394), .ZN(n14944) );
  AOI22_X1 U15726 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12407), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12400) );
  AOI22_X1 U15727 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15728 ( .A1(n12508), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12397) );
  NAND4_X1 U15729 ( .A1(n12400), .A2(n12399), .A3(n12398), .A4(n12397), .ZN(
        n12406) );
  AOI22_X1 U15730 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12404) );
  AOI22_X1 U15731 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12384), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U15732 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12402) );
  AOI22_X1 U15733 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12509), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12401) );
  NAND4_X1 U15734 ( .A1(n12404), .A2(n12403), .A3(n12402), .A4(n12401), .ZN(
        n12405) );
  NOR2_X1 U15735 ( .A1(n12406), .A2(n12405), .ZN(n12427) );
  AOI22_X1 U15736 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12407), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12411) );
  AOI22_X1 U15737 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U15738 ( .A1(n11774), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9662), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12409) );
  AOI22_X1 U15739 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12408) );
  NAND4_X1 U15740 ( .A1(n12411), .A2(n12410), .A3(n12409), .A4(n12408), .ZN(
        n12417) );
  AOI22_X1 U15741 ( .A1(n12450), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U15742 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11804), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U15743 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n9722), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U15744 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12412) );
  NAND4_X1 U15745 ( .A1(n12415), .A2(n12414), .A3(n12413), .A4(n12412), .ZN(
        n12416) );
  NOR2_X1 U15746 ( .A1(n12417), .A2(n12416), .ZN(n12426) );
  XOR2_X1 U15747 ( .A(n12427), .B(n12426), .Z(n12418) );
  NAND2_X1 U15748 ( .A1(n12418), .A2(n12534), .ZN(n12421) );
  INV_X1 U15749 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15180) );
  AOI21_X1 U15750 ( .B1(n15180), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12419) );
  AOI21_X1 U15751 ( .B1(n12104), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12419), .ZN(
        n12420) );
  XNOR2_X1 U15752 ( .A(n12422), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15184) );
  AOI22_X1 U15753 ( .A1(n12421), .A2(n12420), .B1(n12537), .B2(n15184), .ZN(
        n14930) );
  INV_X1 U15754 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n14921) );
  NAND2_X1 U15755 ( .A1(n12424), .A2(n14921), .ZN(n12425) );
  NAND2_X1 U15756 ( .A1(n12461), .A2(n12425), .ZN(n15175) );
  NOR2_X1 U15757 ( .A1(n12427), .A2(n12426), .ZN(n12445) );
  AOI22_X1 U15758 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12431) );
  AOI22_X1 U15759 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12430) );
  AOI22_X1 U15760 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11804), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12429) );
  AOI22_X1 U15761 ( .A1(n12383), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12428) );
  NAND4_X1 U15762 ( .A1(n12431), .A2(n12430), .A3(n12429), .A4(n12428), .ZN(
        n12438) );
  AOI22_X1 U15763 ( .A1(n11774), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12507), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12436) );
  INV_X1 U15764 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n20484) );
  AOI22_X1 U15765 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12435) );
  AOI22_X1 U15766 ( .A1(n12509), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n9662), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12434) );
  AOI22_X1 U15767 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12432), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12433) );
  NAND4_X1 U15768 ( .A1(n12436), .A2(n12435), .A3(n12434), .A4(n12433), .ZN(
        n12437) );
  OR2_X1 U15769 ( .A1(n12438), .A2(n12437), .ZN(n12444) );
  XNOR2_X1 U15770 ( .A(n12445), .B(n12444), .ZN(n12441) );
  AOI21_X1 U15771 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n12006), .A(
        n12560), .ZN(n12440) );
  NAND2_X1 U15772 ( .A1(n12567), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n12439) );
  OAI211_X1 U15773 ( .C1(n12441), .C2(n12563), .A(n12440), .B(n12439), .ZN(
        n12442) );
  OAI21_X1 U15774 ( .B1(n12631), .B2(n15175), .A(n12442), .ZN(n14918) );
  INV_X1 U15775 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15165) );
  NOR2_X1 U15776 ( .A1(n15165), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12443) );
  AOI211_X1 U15777 ( .C1(n12567), .C2(P1_EAX_REG_25__SCAN_IN), .A(n12560), .B(
        n12443), .ZN(n12460) );
  NAND2_X1 U15778 ( .A1(n12445), .A2(n12444), .ZN(n12465) );
  AOI22_X1 U15779 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12449) );
  AOI22_X1 U15780 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12507), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U15781 ( .A1(n11774), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12447) );
  AOI22_X1 U15782 ( .A1(n12508), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12446) );
  NAND4_X1 U15783 ( .A1(n12449), .A2(n12448), .A3(n12447), .A4(n12446), .ZN(
        n12456) );
  AOI22_X1 U15784 ( .A1(n12450), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U15785 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11804), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U15786 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9722), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12452) );
  NAND4_X1 U15787 ( .A1(n12454), .A2(n12453), .A3(n12452), .A4(n12451), .ZN(
        n12455) );
  NOR2_X1 U15788 ( .A1(n12456), .A2(n12455), .ZN(n12466) );
  XOR2_X1 U15789 ( .A(n12465), .B(n12466), .Z(n12457) );
  NAND2_X1 U15790 ( .A1(n12457), .A2(n12534), .ZN(n12459) );
  INV_X1 U15791 ( .A(n12461), .ZN(n12458) );
  XOR2_X1 U15792 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B(n12458), .Z(
        n15169) );
  AOI22_X1 U15793 ( .A1(n12460), .A2(n12459), .B1(n15169), .B2(n12560), .ZN(
        n14906) );
  INV_X1 U15794 ( .A(n12462), .ZN(n12463) );
  INV_X1 U15795 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14896) );
  NAND2_X1 U15796 ( .A1(n12463), .A2(n14896), .ZN(n12464) );
  NAND2_X1 U15797 ( .A1(n12498), .A2(n12464), .ZN(n15156) );
  NOR2_X1 U15798 ( .A1(n12466), .A2(n12465), .ZN(n12483) );
  AOI22_X1 U15799 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12471) );
  AOI22_X1 U15800 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12470) );
  AOI22_X1 U15801 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11804), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12469) );
  AOI22_X1 U15802 ( .A1(n11866), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12468) );
  NAND4_X1 U15803 ( .A1(n12471), .A2(n12470), .A3(n12469), .A4(n12468), .ZN(
        n12477) );
  AOI22_X1 U15804 ( .A1(n11774), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12507), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U15805 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12474) );
  AOI22_X1 U15806 ( .A1(n12509), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12473) );
  AOI22_X1 U15807 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12472) );
  NAND4_X1 U15808 ( .A1(n12475), .A2(n12474), .A3(n12473), .A4(n12472), .ZN(
        n12476) );
  OR2_X1 U15809 ( .A1(n12477), .A2(n12476), .ZN(n12482) );
  XNOR2_X1 U15810 ( .A(n12483), .B(n12482), .ZN(n12480) );
  AOI21_X1 U15811 ( .B1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n12006), .A(
        n12560), .ZN(n12479) );
  NAND2_X1 U15812 ( .A1(n12567), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n12478) );
  OAI211_X1 U15813 ( .C1(n12480), .C2(n12563), .A(n12479), .B(n12478), .ZN(
        n12481) );
  OAI21_X1 U15814 ( .B1(n12631), .B2(n15156), .A(n12481), .ZN(n14895) );
  NAND2_X1 U15815 ( .A1(n12483), .A2(n12482), .ZN(n12501) );
  AOI22_X1 U15816 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12526), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12487) );
  AOI22_X1 U15817 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12384), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12486) );
  AOI22_X1 U15818 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12432), .B1(
        n9662), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12485) );
  NAND4_X1 U15819 ( .A1(n12487), .A2(n12486), .A3(n12485), .A4(n12484), .ZN(
        n12493) );
  AOI22_X1 U15820 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12548), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12491) );
  AOI22_X1 U15821 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12507), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12490) );
  AOI22_X1 U15822 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12543), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12489) );
  AOI22_X1 U15823 ( .A1(n11774), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9723), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12488) );
  NAND4_X1 U15824 ( .A1(n12491), .A2(n12490), .A3(n12489), .A4(n12488), .ZN(
        n12492) );
  NOR2_X1 U15825 ( .A1(n12493), .A2(n12492), .ZN(n12502) );
  XOR2_X1 U15826 ( .A(n12501), .B(n12502), .Z(n12494) );
  NAND2_X1 U15827 ( .A1(n12494), .A2(n12534), .ZN(n12497) );
  INV_X1 U15828 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15143) );
  NOR2_X1 U15829 ( .A1(n15143), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12495) );
  AOI211_X1 U15830 ( .C1(n12104), .C2(P1_EAX_REG_27__SCAN_IN), .A(n12560), .B(
        n12495), .ZN(n12496) );
  XNOR2_X1 U15831 ( .A(n12498), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15145) );
  AOI22_X1 U15832 ( .A1(n12497), .A2(n12496), .B1(n12537), .B2(n15145), .ZN(
        n14882) );
  INV_X1 U15833 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14873) );
  NAND2_X1 U15834 ( .A1(n12499), .A2(n14873), .ZN(n12500) );
  NAND2_X1 U15835 ( .A1(n12540), .A2(n12500), .ZN(n15139) );
  NOR2_X1 U15836 ( .A1(n12502), .A2(n12501), .ZN(n12521) );
  AOI22_X1 U15837 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12506) );
  AOI22_X1 U15838 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12505) );
  AOI22_X1 U15839 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11804), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12504) );
  AOI22_X1 U15840 ( .A1(n11866), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12503) );
  NAND4_X1 U15841 ( .A1(n12506), .A2(n12505), .A3(n12504), .A4(n12503), .ZN(
        n12515) );
  AOI22_X1 U15842 ( .A1(n11774), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12507), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12513) );
  AOI22_X1 U15843 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12512) );
  AOI22_X1 U15844 ( .A1(n9722), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12511) );
  AOI22_X1 U15845 ( .A1(n11860), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12510) );
  NAND4_X1 U15846 ( .A1(n12513), .A2(n12512), .A3(n12511), .A4(n12510), .ZN(
        n12514) );
  OR2_X1 U15847 ( .A1(n12515), .A2(n12514), .ZN(n12520) );
  XNOR2_X1 U15848 ( .A(n12521), .B(n12520), .ZN(n12518) );
  AOI21_X1 U15849 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n12006), .A(
        n12560), .ZN(n12517) );
  NAND2_X1 U15850 ( .A1(n12567), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n12516) );
  OAI211_X1 U15851 ( .C1(n12518), .C2(n12563), .A(n12517), .B(n12516), .ZN(
        n12519) );
  OAI21_X1 U15852 ( .B1(n12631), .B2(n15139), .A(n12519), .ZN(n14870) );
  NAND2_X1 U15853 ( .A1(n12521), .A2(n12520), .ZN(n12556) );
  AOI22_X1 U15854 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12548), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12525) );
  AOI22_X1 U15855 ( .A1(n11866), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11804), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12524) );
  AOI22_X1 U15856 ( .A1(n12508), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12523) );
  AOI22_X1 U15857 ( .A1(n12507), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12522) );
  NAND4_X1 U15858 ( .A1(n12525), .A2(n12524), .A3(n12523), .A4(n12522), .ZN(
        n12533) );
  AOI22_X1 U15859 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12526), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12531) );
  AOI22_X1 U15860 ( .A1(n12235), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12543), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12530) );
  AOI22_X1 U15861 ( .A1(n12224), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U15862 ( .A1(n9866), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(n9722), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12528) );
  NAND4_X1 U15863 ( .A1(n12531), .A2(n12530), .A3(n12529), .A4(n12528), .ZN(
        n12532) );
  NOR2_X1 U15864 ( .A1(n12533), .A2(n12532), .ZN(n12557) );
  XOR2_X1 U15865 ( .A(n12556), .B(n12557), .Z(n12535) );
  NAND2_X1 U15866 ( .A1(n12535), .A2(n12534), .ZN(n12539) );
  INV_X1 U15867 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n13328) );
  NOR2_X1 U15868 ( .A1(n13328), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12536) );
  AOI211_X1 U15869 ( .C1(n12104), .C2(P1_EAX_REG_29__SCAN_IN), .A(n12560), .B(
        n12536), .ZN(n12538) );
  XNOR2_X1 U15870 ( .A(n12540), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14692) );
  AOI22_X1 U15871 ( .A1(n12539), .A2(n12538), .B1(n12537), .B2(n14692), .ZN(
        n13331) );
  INV_X1 U15872 ( .A(n12540), .ZN(n12541) );
  NAND2_X1 U15873 ( .A1(n12541), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12569) );
  XOR2_X1 U15874 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B(n12569), .Z(
        n15127) );
  AOI22_X1 U15875 ( .A1(n12396), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11860), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12547) );
  AOI22_X1 U15876 ( .A1(n11803), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11866), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12546) );
  AOI22_X1 U15877 ( .A1(n12509), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12542), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12545) );
  AOI22_X1 U15878 ( .A1(n12543), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12544) );
  NAND4_X1 U15879 ( .A1(n12547), .A2(n12546), .A3(n12545), .A4(n12544), .ZN(
        n12555) );
  AOI22_X1 U15880 ( .A1(n12548), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12224), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12553) );
  AOI22_X1 U15881 ( .A1(n12384), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11861), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12552) );
  AOI22_X1 U15882 ( .A1(n12549), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12508), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12551) );
  AOI22_X1 U15883 ( .A1(n12526), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9866), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12550) );
  NAND4_X1 U15884 ( .A1(n12553), .A2(n12552), .A3(n12551), .A4(n12550), .ZN(
        n12554) );
  NOR2_X1 U15885 ( .A1(n12555), .A2(n12554), .ZN(n12559) );
  NOR2_X1 U15886 ( .A1(n12557), .A2(n12556), .ZN(n12558) );
  XOR2_X1 U15887 ( .A(n12559), .B(n12558), .Z(n12564) );
  AOI21_X1 U15888 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n12006), .A(
        n12560), .ZN(n12562) );
  NAND2_X1 U15889 ( .A1(n12567), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n12561) );
  OAI211_X1 U15890 ( .C1(n12564), .C2(n12563), .A(n12562), .B(n12561), .ZN(
        n12565) );
  OAI21_X1 U15891 ( .B1(n15127), .B2(n12631), .A(n12565), .ZN(n12767) );
  AOI22_X1 U15892 ( .A1(n12567), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12566), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12568) );
  INV_X1 U15893 ( .A(n12569), .ZN(n12570) );
  NAND2_X1 U15894 ( .A1(n12570), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12571) );
  INV_X1 U15895 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12758) );
  XNOR2_X1 U15896 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12586) );
  NAND2_X1 U15897 ( .A1(n20733), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12594) );
  NAND2_X1 U15898 ( .A1(n12586), .A2(n12587), .ZN(n12574) );
  NAND2_X1 U15899 ( .A1(n20532), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12573) );
  NAND2_X1 U15900 ( .A1(n12574), .A2(n12573), .ZN(n12585) );
  MUX2_X1 U15901 ( .A(n16225), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12584) );
  NAND2_X1 U15902 ( .A1(n12585), .A2(n12584), .ZN(n12576) );
  NAND2_X1 U15903 ( .A1(n16225), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12575) );
  XNOR2_X1 U15904 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12582) );
  NOR2_X1 U15905 ( .A1(n12057), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12577) );
  INV_X1 U15906 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n12578) );
  NAND2_X1 U15907 ( .A1(n12578), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12579) );
  XNOR2_X1 U15908 ( .A(n12583), .B(n12582), .ZN(n12614) );
  XNOR2_X1 U15909 ( .A(n12585), .B(n12584), .ZN(n12608) );
  XNOR2_X1 U15910 ( .A(n12587), .B(n12586), .ZN(n12601) );
  NOR4_X1 U15911 ( .A1(n12617), .A2(n12614), .A3(n12608), .A4(n12601), .ZN(
        n12588) );
  OR2_X1 U15912 ( .A1(n12591), .A2(n12588), .ZN(n14853) );
  NAND2_X1 U15913 ( .A1(n12572), .A2(n13576), .ZN(n13468) );
  INV_X1 U15914 ( .A(n14860), .ZN(n14081) );
  INV_X1 U15915 ( .A(n12591), .ZN(n12590) );
  NAND2_X1 U15916 ( .A1(n12591), .A2(n12596), .ZN(n12627) );
  NAND2_X1 U15917 ( .A1(n12603), .A2(n13675), .ZN(n12624) );
  NAND2_X1 U15918 ( .A1(n12619), .A2(n12617), .ZN(n12623) );
  INV_X1 U15919 ( .A(n12603), .ZN(n12592) );
  NOR2_X1 U15920 ( .A1(n12601), .A2(n12592), .ZN(n12600) );
  NAND2_X1 U15921 ( .A1(n14148), .A2(n11889), .ZN(n12593) );
  NAND2_X1 U15922 ( .A1(n12593), .A2(n14133), .ZN(n12609) );
  OAI21_X1 U15923 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20733), .A(
        n12594), .ZN(n12597) );
  INV_X1 U15924 ( .A(n12597), .ZN(n12595) );
  OAI211_X1 U15925 ( .C1(n11941), .C2(n13323), .A(n12609), .B(n12595), .ZN(
        n12599) );
  INV_X1 U15926 ( .A(n12596), .ZN(n12610) );
  OAI21_X1 U15927 ( .B1(n12610), .B2(n12597), .A(n12615), .ZN(n12598) );
  NAND2_X1 U15928 ( .A1(n12599), .A2(n12598), .ZN(n12602) );
  NAND2_X1 U15929 ( .A1(n12600), .A2(n12602), .ZN(n12607) );
  OAI211_X1 U15930 ( .C1(n12603), .C2(n12602), .A(n12601), .B(n12624), .ZN(
        n12606) );
  NAND2_X1 U15931 ( .A1(n12619), .A2(n12608), .ZN(n12604) );
  OAI211_X1 U15932 ( .C1(n12610), .C2(n12608), .A(n12604), .B(n12609), .ZN(
        n12605) );
  NAND3_X1 U15933 ( .A1(n12607), .A2(n12606), .A3(n12605), .ZN(n12612) );
  AOI22_X1 U15934 ( .A1(n12613), .A2(n12614), .B1(n12612), .B2(n12611), .ZN(
        n12621) );
  INV_X1 U15935 ( .A(n12614), .ZN(n12616) );
  NOR2_X1 U15936 ( .A1(n12616), .A2(n12615), .ZN(n12620) );
  INV_X1 U15937 ( .A(n12617), .ZN(n12618) );
  OAI22_X1 U15938 ( .A1(n12621), .A2(n12620), .B1(n12619), .B2(n12618), .ZN(
        n12622) );
  OAI21_X1 U15939 ( .B1(n12624), .B2(n12623), .A(n12622), .ZN(n12625) );
  AOI21_X1 U15940 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21023), .A(
        n12625), .ZN(n12626) );
  NAND2_X1 U15941 ( .A1(n12627), .A2(n12626), .ZN(n12628) );
  INV_X1 U15942 ( .A(n12630), .ZN(n14852) );
  NAND2_X1 U15943 ( .A1(n12006), .A2(n20942), .ZN(n21022) );
  NOR2_X1 U15944 ( .A1(n20774), .A2(n21022), .ZN(n16464) );
  INV_X1 U15945 ( .A(n16464), .ZN(n16253) );
  NAND2_X1 U15946 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21023), .ZN(n12632) );
  OAI21_X1 U15947 ( .B1(n12632), .B2(n12631), .A(n20432), .ZN(n12633) );
  INV_X1 U15948 ( .A(n12633), .ZN(n12634) );
  OAI21_X1 U15949 ( .B1(n16253), .B2(n21023), .A(n12634), .ZN(n12635) );
  NAND2_X1 U15950 ( .A1(n20334), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14165) );
  NAND2_X1 U15951 ( .A1(n15054), .A2(n20287), .ZN(n12764) );
  NAND2_X1 U15952 ( .A1(n12636), .A2(n11889), .ZN(n12650) );
  INV_X1 U15953 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20451) );
  NAND2_X1 U15954 ( .A1(n12650), .A2(n20451), .ZN(n12639) );
  INV_X1 U15955 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n20341) );
  NAND2_X1 U15956 ( .A1(n14857), .A2(n20341), .ZN(n12638) );
  NAND3_X1 U15957 ( .A1(n12639), .A2(n12637), .A3(n12638), .ZN(n12640) );
  INV_X1 U15958 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13814) );
  NAND2_X1 U15959 ( .A1(n12637), .A2(n13814), .ZN(n12642) );
  INV_X1 U15960 ( .A(n12650), .ZN(n12645) );
  NAND2_X1 U15961 ( .A1(n12650), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12641) );
  OR2_X1 U15962 ( .A1(n20350), .A2(n14084), .ZN(n12644) );
  INV_X1 U15963 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20464) );
  NAND2_X1 U15964 ( .A1(n12650), .A2(n20464), .ZN(n12648) );
  INV_X1 U15965 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n12646) );
  NAND2_X1 U15966 ( .A1(n14857), .A2(n12646), .ZN(n12647) );
  NAND3_X1 U15967 ( .A1(n12648), .A2(n12637), .A3(n12647), .ZN(n12649) );
  OAI21_X1 U15968 ( .B1(n12738), .B2(P1_EBX_REG_2__SCAN_IN), .A(n12649), .ZN(
        n13827) );
  MUX2_X1 U15969 ( .A(n12727), .B(n12637), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12652) );
  INV_X1 U15970 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20447) );
  NAND2_X1 U15971 ( .A1(n13811), .A2(n20447), .ZN(n12651) );
  NAND2_X1 U15972 ( .A1(n12652), .A2(n12651), .ZN(n13903) );
  MUX2_X1 U15973 ( .A(n12738), .B(n12650), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n12655) );
  NAND2_X1 U15974 ( .A1(n12645), .A2(n14084), .ZN(n12683) );
  NAND2_X1 U15975 ( .A1(n14084), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12653) );
  AND2_X1 U15976 ( .A1(n12683), .A2(n12653), .ZN(n12654) );
  NAND2_X1 U15977 ( .A1(n12655), .A2(n12654), .ZN(n14062) );
  INV_X1 U15978 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16447) );
  INV_X1 U15979 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20297) );
  NAND2_X1 U15980 ( .A1(n14857), .A2(n20297), .ZN(n12656) );
  OAI211_X1 U15981 ( .C1(n12739), .C2(n16447), .A(n12656), .B(n12650), .ZN(
        n12657) );
  OAI21_X1 U15982 ( .B1(n12727), .B2(P1_EBX_REG_5__SCAN_IN), .A(n12657), .ZN(
        n13983) );
  MUX2_X1 U15983 ( .A(n12738), .B(n12650), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n12662) );
  NAND2_X1 U15984 ( .A1(n14084), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12660) );
  AND2_X1 U15985 ( .A1(n12683), .A2(n12660), .ZN(n12661) );
  NAND2_X1 U15986 ( .A1(n12662), .A2(n12661), .ZN(n14283) );
  INV_X1 U15987 ( .A(n14283), .ZN(n12663) );
  INV_X1 U15988 ( .A(n12727), .ZN(n12664) );
  INV_X1 U15989 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n20272) );
  NAND2_X1 U15990 ( .A1(n12664), .A2(n20272), .ZN(n12667) );
  INV_X1 U15991 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16439) );
  NAND2_X1 U15992 ( .A1(n14857), .A2(n20272), .ZN(n12665) );
  OAI211_X1 U15993 ( .C1(n12739), .C2(n16439), .A(n12665), .B(n12650), .ZN(
        n12666) );
  MUX2_X1 U15994 ( .A(n12738), .B(n12650), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n12670) );
  NAND2_X1 U15995 ( .A1(n14084), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12668) );
  AND2_X1 U15996 ( .A1(n12683), .A2(n12668), .ZN(n12669) );
  NAND2_X1 U15997 ( .A1(n12670), .A2(n12669), .ZN(n14408) );
  INV_X1 U15998 ( .A(n14408), .ZN(n12671) );
  INV_X1 U15999 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16420) );
  INV_X1 U16000 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n12672) );
  NAND2_X1 U16001 ( .A1(n14857), .A2(n12672), .ZN(n12673) );
  OAI211_X1 U16002 ( .C1(n12739), .C2(n16420), .A(n12673), .B(n12650), .ZN(
        n12674) );
  OAI21_X1 U16003 ( .B1(n12727), .B2(P1_EBX_REG_9__SCAN_IN), .A(n12674), .ZN(
        n14430) );
  INV_X1 U16004 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14561) );
  NAND2_X1 U16005 ( .A1(n12730), .A2(n14561), .ZN(n12679) );
  INV_X1 U16006 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12675) );
  NAND2_X1 U16007 ( .A1(n12650), .A2(n12675), .ZN(n12677) );
  NAND2_X1 U16008 ( .A1(n14857), .A2(n14561), .ZN(n12676) );
  NAND3_X1 U16009 ( .A1(n12677), .A2(n12637), .A3(n12676), .ZN(n12678) );
  MUX2_X1 U16010 ( .A(n12727), .B(n12637), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12681) );
  INV_X1 U16011 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16395) );
  NAND2_X1 U16012 ( .A1(n16395), .A2(n13811), .ZN(n12680) );
  MUX2_X1 U16013 ( .A(n12738), .B(n12650), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n12685) );
  NAND2_X1 U16014 ( .A1(n14084), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12682) );
  AND2_X1 U16015 ( .A1(n12683), .A2(n12682), .ZN(n12684) );
  NAND2_X1 U16016 ( .A1(n12685), .A2(n12684), .ZN(n14493) );
  INV_X1 U16017 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15413) );
  INV_X1 U16018 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14537) );
  NAND2_X1 U16019 ( .A1(n14857), .A2(n14537), .ZN(n12686) );
  OAI211_X1 U16020 ( .C1(n12739), .C2(n15413), .A(n12686), .B(n12650), .ZN(
        n12687) );
  OAI21_X1 U16021 ( .B1(n12727), .B2(P1_EBX_REG_13__SCAN_IN), .A(n12687), .ZN(
        n14534) );
  MUX2_X1 U16022 ( .A(n12738), .B(n12650), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n12689) );
  NAND2_X1 U16023 ( .A1(n14084), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12688) );
  NAND2_X1 U16024 ( .A1(n12689), .A2(n12688), .ZN(n14576) );
  MUX2_X1 U16025 ( .A(n12727), .B(n12637), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12691) );
  INV_X1 U16026 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16393) );
  NAND2_X1 U16027 ( .A1(n13811), .A2(n16393), .ZN(n12690) );
  NAND2_X1 U16028 ( .A1(n12691), .A2(n12690), .ZN(n14588) );
  INV_X1 U16029 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n16291) );
  NAND2_X1 U16030 ( .A1(n12730), .A2(n16291), .ZN(n12695) );
  INV_X1 U16031 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15439) );
  NAND2_X1 U16032 ( .A1(n12650), .A2(n15439), .ZN(n12693) );
  NAND2_X1 U16033 ( .A1(n14857), .A2(n16291), .ZN(n12692) );
  NAND3_X1 U16034 ( .A1(n12693), .A2(n12637), .A3(n12692), .ZN(n12694) );
  MUX2_X1 U16035 ( .A(n12727), .B(n12637), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12697) );
  OAI21_X1 U16036 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n12769), .A(
        n12697), .ZN(n15007) );
  INV_X1 U16037 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n12698) );
  NAND2_X1 U16038 ( .A1(n12730), .A2(n12698), .ZN(n12702) );
  INV_X1 U16039 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15419) );
  NAND2_X1 U16040 ( .A1(n12650), .A2(n15419), .ZN(n12700) );
  NAND2_X1 U16041 ( .A1(n14857), .A2(n12698), .ZN(n12699) );
  NAND3_X1 U16042 ( .A1(n12700), .A2(n12637), .A3(n12699), .ZN(n12701) );
  INV_X1 U16043 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15401) );
  INV_X1 U16044 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n12703) );
  NAND2_X1 U16045 ( .A1(n14857), .A2(n12703), .ZN(n12704) );
  OAI211_X1 U16046 ( .C1(n12739), .C2(n15401), .A(n12704), .B(n12650), .ZN(
        n12705) );
  OAI21_X1 U16047 ( .B1(n12727), .B2(P1_EBX_REG_19__SCAN_IN), .A(n12705), .ZN(
        n14991) );
  MUX2_X1 U16048 ( .A(n12738), .B(n12650), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n12708) );
  NAND2_X1 U16049 ( .A1(n14084), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12707) );
  NAND2_X1 U16050 ( .A1(n12708), .A2(n12707), .ZN(n14956) );
  INV_X1 U16051 ( .A(n14956), .ZN(n14977) );
  MUX2_X1 U16052 ( .A(n12727), .B(n12637), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n12710) );
  INV_X1 U16053 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n13316) );
  NAND2_X1 U16054 ( .A1(n13811), .A2(n13316), .ZN(n12709) );
  NAND2_X1 U16055 ( .A1(n12710), .A2(n12709), .ZN(n14959) );
  MUX2_X1 U16056 ( .A(n12727), .B(n12637), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12712) );
  INV_X1 U16057 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15343) );
  NAND2_X1 U16058 ( .A1(n13811), .A2(n15343), .ZN(n12711) );
  AND2_X1 U16059 ( .A1(n12712), .A2(n12711), .ZN(n14932) );
  INV_X1 U16060 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15370) );
  NAND2_X1 U16061 ( .A1(n12650), .A2(n15370), .ZN(n12714) );
  INV_X1 U16062 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15026) );
  NAND2_X1 U16063 ( .A1(n14857), .A2(n15026), .ZN(n12713) );
  NAND3_X1 U16064 ( .A1(n12714), .A2(n12637), .A3(n12713), .ZN(n12715) );
  OAI21_X1 U16065 ( .B1(n12738), .B2(P1_EBX_REG_22__SCAN_IN), .A(n12715), .ZN(
        n14943) );
  NAND2_X1 U16066 ( .A1(n14932), .A2(n14943), .ZN(n12716) );
  INV_X1 U16067 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n12717) );
  NAND2_X1 U16068 ( .A1(n12730), .A2(n12717), .ZN(n12721) );
  INV_X1 U16069 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15346) );
  NAND2_X1 U16070 ( .A1(n12650), .A2(n15346), .ZN(n12719) );
  NAND2_X1 U16071 ( .A1(n14857), .A2(n12717), .ZN(n12718) );
  NAND3_X1 U16072 ( .A1(n12719), .A2(n12637), .A3(n12718), .ZN(n12720) );
  MUX2_X1 U16073 ( .A(n12727), .B(n12637), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12723) );
  INV_X1 U16074 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15324) );
  NAND2_X1 U16075 ( .A1(n13811), .A2(n15324), .ZN(n12722) );
  AND2_X1 U16076 ( .A1(n12723), .A2(n12722), .ZN(n14913) );
  INV_X1 U16077 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15322) );
  NAND2_X1 U16078 ( .A1(n12650), .A2(n15322), .ZN(n12725) );
  INV_X1 U16079 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15019) );
  NAND2_X1 U16080 ( .A1(n14857), .A2(n15019), .ZN(n12724) );
  NAND3_X1 U16081 ( .A1(n12725), .A2(n12637), .A3(n12724), .ZN(n12726) );
  OAI21_X1 U16082 ( .B1(n12738), .B2(P1_EBX_REG_26__SCAN_IN), .A(n12726), .ZN(
        n14892) );
  MUX2_X1 U16083 ( .A(n12727), .B(n12637), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12729) );
  INV_X1 U16084 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15316) );
  NAND2_X1 U16085 ( .A1(n13811), .A2(n15316), .ZN(n12728) );
  NAND2_X1 U16086 ( .A1(n12729), .A2(n12728), .ZN(n14884) );
  INV_X1 U16087 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n12731) );
  NAND2_X1 U16088 ( .A1(n12730), .A2(n12731), .ZN(n12735) );
  INV_X1 U16089 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15306) );
  NAND2_X1 U16090 ( .A1(n12650), .A2(n15306), .ZN(n12733) );
  NAND2_X1 U16091 ( .A1(n14857), .A2(n12731), .ZN(n12732) );
  NAND3_X1 U16092 ( .A1(n12733), .A2(n12637), .A3(n12732), .ZN(n12734) );
  AND2_X1 U16093 ( .A1(n12735), .A2(n12734), .ZN(n14872) );
  OR2_X1 U16094 ( .A1(n12769), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12737) );
  INV_X1 U16095 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14704) );
  NAND2_X1 U16096 ( .A1(n14857), .A2(n14704), .ZN(n12736) );
  NAND2_X1 U16097 ( .A1(n12737), .A2(n12736), .ZN(n12780) );
  OAI22_X1 U16098 ( .A1(n12780), .A2(n12739), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n12738), .ZN(n14687) );
  INV_X1 U16099 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15288) );
  NOR2_X1 U16100 ( .A1(n14857), .A2(n15288), .ZN(n12740) );
  AOI21_X1 U16101 ( .B1(n12769), .B2(P1_EBX_REG_30__SCAN_IN), .A(n12740), .ZN(
        n12783) );
  AOI22_X1 U16102 ( .A1(n12769), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n14084), .ZN(n12743) );
  NAND2_X1 U16103 ( .A1(n13675), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12753) );
  NAND2_X1 U16104 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21027) );
  AND2_X1 U16105 ( .A1(n21027), .A2(n21170), .ZN(n16243) );
  NOR2_X1 U16106 ( .A1(n12753), .A2(n16243), .ZN(n12745) );
  INV_X1 U16107 ( .A(n12746), .ZN(n12747) );
  INV_X1 U16108 ( .A(n16265), .ZN(n13674) );
  NAND2_X1 U16109 ( .A1(n14133), .A2(n13674), .ZN(n13685) );
  AND2_X1 U16110 ( .A1(n13685), .A2(n16243), .ZN(n12755) );
  NAND4_X1 U16111 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_4__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n20275)
         );
  NAND4_X1 U16112 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n20256)
         );
  NOR2_X1 U16113 ( .A1(n20275), .A2(n20256), .ZN(n14406) );
  NAND3_X1 U16114 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(n14406), .ZN(n14971) );
  NAND4_X1 U16115 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_11__SCAN_IN), .ZN(n14989) );
  NAND3_X1 U16116 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .ZN(n14974) );
  NOR3_X1 U16117 ( .A1(n14971), .A2(n14989), .A3(n14974), .ZN(n12749) );
  NAND2_X1 U16118 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n14976) );
  INV_X1 U16119 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15207) );
  NOR2_X1 U16120 ( .A1(n14976), .A2(n15207), .ZN(n12748) );
  AND2_X1 U16121 ( .A1(n12749), .A2(n12748), .ZN(n14946) );
  AND2_X1 U16122 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n12750) );
  NAND2_X1 U16123 ( .A1(n14946), .A2(n12750), .ZN(n14936) );
  INV_X1 U16124 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n21093) );
  OR2_X1 U16125 ( .A1(n14936), .A2(n21093), .ZN(n14922) );
  NAND2_X1 U16126 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n12751) );
  NOR2_X1 U16127 ( .A1(n14922), .A2(n12751), .ZN(n14897) );
  NAND2_X1 U16128 ( .A1(n14897), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14885) );
  INV_X1 U16129 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n21199) );
  INV_X1 U16130 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n21038) );
  NOR3_X1 U16131 ( .A1(n14885), .A2(n21199), .A3(n21038), .ZN(n14874) );
  INV_X1 U16132 ( .A(n14874), .ZN(n14690) );
  INV_X1 U16133 ( .A(n20334), .ZN(n20276) );
  AOI21_X1 U16134 ( .B1(n20347), .B2(n14690), .A(n20276), .ZN(n14878) );
  INV_X1 U16135 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n21096) );
  INV_X1 U16136 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n21108) );
  OAI21_X1 U16137 ( .B1(n21096), .B2(n21108), .A(n20347), .ZN(n12752) );
  NAND2_X1 U16138 ( .A1(n14878), .A2(n12752), .ZN(n14862) );
  INV_X1 U16139 ( .A(n12753), .ZN(n12754) );
  NOR2_X1 U16140 ( .A1(n12755), .A2(n12754), .ZN(n12756) );
  NAND2_X1 U16141 ( .A1(n12757), .A2(n12756), .ZN(n20340) );
  INV_X1 U16142 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15015) );
  OAI22_X1 U16143 ( .A1(n20340), .A2(n15015), .B1(n12758), .B2(n20335), .ZN(
        n12760) );
  NAND3_X1 U16144 ( .A1(n20347), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n14874), 
        .ZN(n14864) );
  NOR3_X1 U16145 ( .A1(n14864), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n21108), 
        .ZN(n12759) );
  AOI211_X1 U16146 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14862), .A(n12760), 
        .B(n12759), .ZN(n12761) );
  NAND2_X1 U16147 ( .A1(n12764), .A2(n12763), .ZN(P1_U2809) );
  INV_X1 U16148 ( .A(n15129), .ZN(n12787) );
  NOR2_X1 U16149 ( .A1(n11885), .A2(n14162), .ZN(n12768) );
  AOI21_X1 U16150 ( .B1(n12769), .B2(n13321), .A(n12768), .ZN(n13555) );
  MUX2_X1 U16151 ( .A(n12771), .B(n12770), .S(n11889), .Z(n12772) );
  NAND3_X1 U16152 ( .A1(n13555), .A2(n12773), .A3(n12772), .ZN(n13699) );
  NAND2_X1 U16153 ( .A1(n9717), .A2(n14106), .ZN(n12774) );
  NAND3_X1 U16154 ( .A1(n13546), .A2(n9717), .A3(n9669), .ZN(n12776) );
  INV_X1 U16155 ( .A(n12777), .ZN(n12778) );
  NAND4_X1 U16156 ( .A1(n12778), .A2(n14106), .A3(n15052), .A4(n13865), .ZN(
        n14080) );
  OAI22_X1 U16157 ( .A1(n14850), .A2(n13682), .B1(n14084), .B2(n14080), .ZN(
        n12779) );
  OAI22_X1 U16158 ( .A1(n14689), .A2(n12637), .B1(n12781), .B2(n12780), .ZN(
        n12782) );
  INV_X1 U16159 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n12784) );
  OAI22_X1 U16160 ( .A1(n15285), .A2(n15048), .B1(n12784), .B2(n15047), .ZN(
        n12785) );
  INV_X1 U16161 ( .A(n12785), .ZN(n12786) );
  NAND2_X1 U16162 ( .A1(n12788), .A2(n12809), .ZN(n12794) );
  NAND2_X1 U16163 ( .A1(n13746), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12789) );
  NOR2_X1 U16164 ( .A1(n20182), .A2(n20193), .ZN(n19979) );
  INV_X1 U16165 ( .A(n12810), .ZN(n12791) );
  NAND2_X1 U16166 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19872) );
  NAND2_X1 U16167 ( .A1(n19872), .A2(n20182), .ZN(n12790) );
  NAND2_X1 U16168 ( .A1(n12791), .A2(n12790), .ZN(n19663) );
  NOR2_X1 U16169 ( .A1(n19663), .A2(n20016), .ZN(n12792) );
  AOI21_X1 U16170 ( .B1(n12813), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12792), .ZN(n12793) );
  NAND2_X1 U16171 ( .A1(n13750), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12803) );
  NAND2_X1 U16172 ( .A1(n12813), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12796) );
  XNOR2_X1 U16173 ( .A(n20202), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19662) );
  NAND2_X1 U16174 ( .A1(n19662), .A2(n20170), .ZN(n19841) );
  NAND2_X1 U16175 ( .A1(n12796), .A2(n19841), .ZN(n12797) );
  NOR2_X1 U16176 ( .A1(n20016), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12798) );
  AOI21_X1 U16177 ( .B1(n12813), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12798), .ZN(n12799) );
  NAND2_X1 U16178 ( .A1(n13750), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12801) );
  NAND2_X1 U16179 ( .A1(n13622), .A2(n12801), .ZN(n12802) );
  NAND2_X1 U16180 ( .A1(n13640), .A2(n13641), .ZN(n12807) );
  INV_X1 U16181 ( .A(n12803), .ZN(n12804) );
  NAND2_X1 U16182 ( .A1(n12805), .A2(n12804), .ZN(n12806) );
  NAND2_X1 U16183 ( .A1(n9734), .A2(n12809), .ZN(n12815) );
  OAI21_X1 U16184 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n12810), .A(
        n20170), .ZN(n12811) );
  NOR2_X1 U16185 ( .A1(n12811), .A2(n20067), .ZN(n12812) );
  AOI21_X1 U16186 ( .B1(n12813), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12812), .ZN(n12814) );
  AND2_X1 U16187 ( .A1(n13741), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12819) );
  INV_X1 U16188 ( .A(n13741), .ZN(n12817) );
  NAND2_X1 U16189 ( .A1(n13750), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n13745) );
  NAND3_X1 U16190 ( .A1(n15586), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12816) );
  NAND2_X1 U16191 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12820) );
  NOR2_X1 U16192 ( .A1(n10111), .A2(n13909), .ZN(n13937) );
  AND2_X1 U16193 ( .A1(n13986), .A2(n13937), .ZN(n12822) );
  NAND2_X1 U16194 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12825) );
  NAND2_X1 U16195 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12824) );
  OAI211_X1 U16196 ( .C1(n12963), .C2(n12826), .A(n12825), .B(n12824), .ZN(
        n12830) );
  INV_X1 U16197 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12828) );
  INV_X1 U16198 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12827) );
  OAI22_X1 U16199 ( .A1(n12897), .A2(n12828), .B1(n12896), .B2(n12827), .ZN(
        n12829) );
  NOR2_X1 U16200 ( .A1(n12830), .A2(n12829), .ZN(n12838) );
  INV_X1 U16201 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19532) );
  AOI22_X1 U16202 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10460), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U16203 ( .A1(n10385), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U16204 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12832) );
  NAND2_X1 U16205 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12831) );
  AND4_X1 U16206 ( .A1(n12834), .A2(n12833), .A3(n12832), .A4(n12831), .ZN(
        n12837) );
  AOI22_X1 U16207 ( .A1(n12905), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12904), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12836) );
  AOI22_X1 U16208 ( .A1(n12907), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12906), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12835) );
  NAND4_X1 U16209 ( .A1(n12838), .A2(n12837), .A3(n12836), .A4(n12835), .ZN(
        n14421) );
  INV_X1 U16210 ( .A(n14420), .ZN(n12857) );
  AOI22_X1 U16211 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10460), .B1(
        n10383), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12842) );
  AOI22_X1 U16212 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10384), .B1(
        n10385), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12841) );
  AOI22_X1 U16213 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10396), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12840) );
  NAND2_X1 U16214 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12839) );
  NAND4_X1 U16215 ( .A1(n12842), .A2(n12841), .A3(n12840), .A4(n12839), .ZN(
        n12849) );
  OAI22_X1 U16216 ( .A1(n12953), .A2(n12844), .B1(n12951), .B2(n12843), .ZN(
        n12848) );
  OAI22_X1 U16217 ( .A1(n12846), .A2(n12956), .B1(n12955), .B2(n12845), .ZN(
        n12847) );
  OR3_X1 U16218 ( .A1(n12849), .A2(n12848), .A3(n12847), .ZN(n12855) );
  AOI22_X1 U16219 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12853) );
  NAND2_X1 U16220 ( .A1(n12961), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12852) );
  NAND2_X1 U16221 ( .A1(n12960), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12851) );
  NAND2_X1 U16222 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12850) );
  NAND4_X1 U16223 ( .A1(n12853), .A2(n12852), .A3(n12851), .A4(n12850), .ZN(
        n12854) );
  NOR2_X1 U16224 ( .A1(n12855), .A2(n12854), .ZN(n14471) );
  NAND2_X1 U16225 ( .A1(n12857), .A2(n12856), .ZN(n14470) );
  INV_X1 U16226 ( .A(n14470), .ZN(n12875) );
  AOI22_X1 U16227 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10383), .B1(
        n10460), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12861) );
  AOI22_X1 U16228 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10385), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12860) );
  AOI22_X1 U16229 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10396), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12859) );
  NAND2_X1 U16230 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12858) );
  NAND4_X1 U16231 ( .A1(n12861), .A2(n12860), .A3(n12859), .A4(n12858), .ZN(
        n12867) );
  INV_X1 U16232 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12862) );
  OAI22_X1 U16233 ( .A1(n12953), .A2(n13037), .B1(n12951), .B2(n12862), .ZN(
        n12866) );
  INV_X1 U16234 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12863) );
  OAI22_X1 U16235 ( .A1(n12864), .A2(n12956), .B1(n12955), .B2(n12863), .ZN(
        n12865) );
  OR3_X1 U16236 ( .A1(n12867), .A2(n12866), .A3(n12865), .ZN(n12873) );
  AOI22_X1 U16237 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12871) );
  NAND2_X1 U16238 ( .A1(n12961), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n12870) );
  NAND2_X1 U16239 ( .A1(n12960), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12869) );
  NAND2_X1 U16240 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12868) );
  NAND4_X1 U16241 ( .A1(n12871), .A2(n12870), .A3(n12869), .A4(n12868), .ZN(
        n12872) );
  NOR2_X1 U16242 ( .A1(n12873), .A2(n12872), .ZN(n14624) );
  INV_X1 U16243 ( .A(n14624), .ZN(n12874) );
  AOI22_X1 U16244 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10383), .B1(
        n10460), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12879) );
  AOI22_X1 U16245 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10385), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12878) );
  AOI22_X1 U16246 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10395), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12877) );
  NAND2_X1 U16247 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12876) );
  NAND4_X1 U16248 ( .A1(n12879), .A2(n12878), .A3(n12877), .A4(n12876), .ZN(
        n12885) );
  OAI22_X1 U16249 ( .A1(n12953), .A2(n13062), .B1(n12951), .B2(n12880), .ZN(
        n12884) );
  OAI22_X1 U16250 ( .A1(n12882), .A2(n12956), .B1(n12955), .B2(n12881), .ZN(
        n12883) );
  OR3_X1 U16251 ( .A1(n12885), .A2(n12884), .A3(n12883), .ZN(n12891) );
  AOI22_X1 U16252 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12889) );
  NAND2_X1 U16253 ( .A1(n12961), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n12888) );
  NAND2_X1 U16254 ( .A1(n12960), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12887) );
  NAND2_X1 U16255 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12886) );
  NAND4_X1 U16256 ( .A1(n12889), .A2(n12888), .A3(n12887), .A4(n12886), .ZN(
        n12890) );
  NOR2_X1 U16257 ( .A1(n12891), .A2(n12890), .ZN(n14642) );
  NAND2_X1 U16258 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12893) );
  NAND2_X1 U16259 ( .A1(n12965), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12892) );
  OAI211_X1 U16260 ( .C1(n12963), .C2(n12894), .A(n12893), .B(n12892), .ZN(
        n12899) );
  INV_X1 U16261 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12895) );
  OAI22_X1 U16262 ( .A1(n12897), .A2(n10466), .B1(n12896), .B2(n12895), .ZN(
        n12898) );
  NOR2_X1 U16263 ( .A1(n12899), .A2(n12898), .ZN(n12911) );
  AOI22_X1 U16264 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n10383), .B1(
        n10460), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12903) );
  AOI22_X1 U16265 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10385), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12902) );
  AOI22_X1 U16266 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10396), .B1(
        n10395), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12901) );
  NAND2_X1 U16267 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12900) );
  AND4_X1 U16268 ( .A1(n12903), .A2(n12902), .A3(n12901), .A4(n12900), .ZN(
        n12910) );
  AOI22_X1 U16269 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12905), .B1(
        n12904), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12909) );
  AOI22_X1 U16270 ( .A1(n12907), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12906), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12908) );
  NAND4_X1 U16271 ( .A1(n12911), .A2(n12910), .A3(n12909), .A4(n12908), .ZN(
        n15612) );
  AOI22_X1 U16272 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10460), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12915) );
  AOI22_X1 U16273 ( .A1(n10385), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12914) );
  AOI22_X1 U16274 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12913) );
  NAND2_X1 U16275 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12912) );
  NAND4_X1 U16276 ( .A1(n12915), .A2(n12914), .A3(n12913), .A4(n12912), .ZN(
        n12920) );
  OAI22_X1 U16277 ( .A1(n12953), .A2(n13117), .B1(n12951), .B2(n13105), .ZN(
        n12919) );
  OAI22_X1 U16278 ( .A1(n12956), .A2(n12917), .B1(n12955), .B2(n12916), .ZN(
        n12918) );
  OR3_X1 U16279 ( .A1(n12920), .A2(n12919), .A3(n12918), .ZN(n12926) );
  AOI22_X1 U16280 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12924) );
  NAND2_X1 U16281 ( .A1(n12961), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n12923) );
  NAND2_X1 U16282 ( .A1(n12960), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12922) );
  NAND2_X1 U16283 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12921) );
  NAND4_X1 U16284 ( .A1(n12924), .A2(n12923), .A3(n12922), .A4(n12921), .ZN(
        n12925) );
  NOR2_X1 U16285 ( .A1(n12926), .A2(n12925), .ZN(n15608) );
  INV_X1 U16286 ( .A(n15608), .ZN(n12927) );
  NAND2_X1 U16287 ( .A1(n12928), .A2(n12927), .ZN(n15600) );
  AOI22_X1 U16288 ( .A1(n10383), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10460), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12933) );
  AOI22_X1 U16289 ( .A1(n10385), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12932) );
  AOI22_X1 U16290 ( .A1(n10395), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12931) );
  NAND2_X1 U16291 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12930) );
  NAND4_X1 U16292 ( .A1(n12933), .A2(n12932), .A3(n12931), .A4(n12930), .ZN(
        n12938) );
  OAI22_X1 U16293 ( .A1(n12953), .A2(n13127), .B1(n12951), .B2(n10524), .ZN(
        n12937) );
  OAI22_X1 U16294 ( .A1(n12956), .A2(n12935), .B1(n12955), .B2(n12934), .ZN(
        n12936) );
  OR3_X1 U16295 ( .A1(n12938), .A2(n12937), .A3(n12936), .ZN(n12945) );
  AOI22_X1 U16296 ( .A1(n12964), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12965), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12943) );
  NAND2_X1 U16297 ( .A1(n12961), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n12942) );
  NAND2_X1 U16298 ( .A1(n12960), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12941) );
  NAND2_X1 U16299 ( .A1(n12939), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12940) );
  NAND4_X1 U16300 ( .A1(n12943), .A2(n12942), .A3(n12941), .A4(n12940), .ZN(
        n12944) );
  NOR2_X1 U16301 ( .A1(n12945), .A2(n12944), .ZN(n15601) );
  AOI22_X1 U16302 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10383), .B1(
        n10460), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12949) );
  AOI22_X1 U16303 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10385), .B1(
        n10384), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12948) );
  AOI22_X1 U16304 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10395), .B1(
        n10396), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12947) );
  NAND2_X1 U16305 ( .A1(n12929), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12946) );
  AND4_X1 U16306 ( .A1(n12949), .A2(n12948), .A3(n12947), .A4(n12946), .ZN(
        n12975) );
  INV_X1 U16307 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12952) );
  INV_X1 U16308 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12950) );
  OAI22_X1 U16309 ( .A1(n12953), .A2(n12952), .B1(n12951), .B2(n12950), .ZN(
        n12959) );
  INV_X1 U16310 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12954) );
  OAI22_X1 U16311 ( .A1(n12957), .A2(n12956), .B1(n12955), .B2(n12954), .ZN(
        n12958) );
  NOR2_X1 U16312 ( .A1(n12959), .A2(n12958), .ZN(n12974) );
  AOI22_X1 U16313 ( .A1(n12961), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12960), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12973) );
  NOR2_X1 U16314 ( .A1(n12963), .A2(n12962), .ZN(n12971) );
  INV_X1 U16315 ( .A(n12964), .ZN(n12969) );
  INV_X1 U16316 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12968) );
  INV_X1 U16317 ( .A(n12965), .ZN(n12967) );
  OAI22_X1 U16318 ( .A1(n12969), .A2(n12968), .B1(n12967), .B2(n12966), .ZN(
        n12970) );
  NOR2_X1 U16319 ( .A1(n12971), .A2(n12970), .ZN(n12972) );
  NAND4_X1 U16320 ( .A1(n12975), .A2(n12974), .A3(n12973), .A4(n12972), .ZN(
        n12997) );
  INV_X1 U16321 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12980) );
  INV_X1 U16322 ( .A(n12976), .ZN(n12978) );
  NAND2_X1 U16323 ( .A1(n12978), .A2(n12977), .ZN(n13154) );
  INV_X1 U16324 ( .A(n10188), .ZN(n13132) );
  INV_X1 U16325 ( .A(n13132), .ZN(n13163) );
  NAND2_X1 U16326 ( .A1(n13163), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12979) );
  OAI211_X1 U16327 ( .C1(n13128), .C2(n12980), .A(n13154), .B(n12979), .ZN(
        n12981) );
  INV_X1 U16328 ( .A(n12981), .ZN(n12987) );
  AOI22_X1 U16329 ( .A1(n9686), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n13150), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12986) );
  AOI22_X1 U16330 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13090), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12985) );
  INV_X1 U16331 ( .A(n12983), .ZN(n13156) );
  AOI22_X1 U16332 ( .A1(n13147), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12984) );
  NAND4_X1 U16333 ( .A1(n12987), .A2(n12986), .A3(n12985), .A4(n12984), .ZN(
        n12996) );
  INV_X1 U16334 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12989) );
  INV_X1 U16335 ( .A(n13154), .ZN(n13113) );
  NAND2_X1 U16336 ( .A1(n13163), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12988) );
  OAI211_X1 U16337 ( .C1(n13128), .C2(n12989), .A(n13113), .B(n12988), .ZN(
        n12990) );
  INV_X1 U16338 ( .A(n12990), .ZN(n12994) );
  AOI22_X1 U16339 ( .A1(n9686), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13150), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12993) );
  AOI22_X1 U16340 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9665), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12992) );
  AOI22_X1 U16341 ( .A1(n13147), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12991) );
  NAND4_X1 U16342 ( .A1(n12994), .A2(n12993), .A3(n12992), .A4(n12991), .ZN(
        n12995) );
  AND2_X1 U16343 ( .A1(n12997), .A2(n13003), .ZN(n13023) );
  NAND2_X1 U16344 ( .A1(n13023), .A2(n15586), .ZN(n13001) );
  INV_X1 U16345 ( .A(n12997), .ZN(n12999) );
  NAND2_X1 U16346 ( .A1(n15586), .A2(n13003), .ZN(n12998) );
  NAND2_X1 U16347 ( .A1(n12999), .A2(n12998), .ZN(n13000) );
  NAND2_X1 U16348 ( .A1(n13001), .A2(n13000), .ZN(n13027) );
  XNOR2_X1 U16349 ( .A(n13004), .B(n13002), .ZN(n15593) );
  NAND2_X1 U16350 ( .A1(n9730), .A2(n13003), .ZN(n15594) );
  AOI22_X1 U16351 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n13162), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13012) );
  AOI22_X1 U16352 ( .A1(n13147), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13011) );
  AOI22_X1 U16353 ( .A1(n14000), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9665), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13010) );
  OR2_X1 U16354 ( .A1(n13132), .A2(n13005), .ZN(n13006) );
  OAI211_X1 U16355 ( .C1(n13007), .C2(n12845), .A(n13113), .B(n13006), .ZN(
        n13008) );
  INV_X1 U16356 ( .A(n13008), .ZN(n13009) );
  NAND4_X1 U16357 ( .A1(n13012), .A2(n13011), .A3(n13010), .A4(n13009), .ZN(
        n13021) );
  INV_X1 U16358 ( .A(n13091), .ZN(n13159) );
  OR2_X1 U16359 ( .A1(n13156), .A2(n19537), .ZN(n13013) );
  OAI211_X1 U16360 ( .C1(n13159), .C2(n13014), .A(n13154), .B(n13013), .ZN(
        n13015) );
  INV_X1 U16361 ( .A(n13015), .ZN(n13019) );
  AOI22_X1 U16362 ( .A1(n9686), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n13150), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13018) );
  AOI22_X1 U16363 ( .A1(n13162), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9665), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13017) );
  AOI22_X1 U16364 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13163), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13016) );
  NAND4_X1 U16365 ( .A1(n13019), .A2(n13018), .A3(n13017), .A4(n13016), .ZN(
        n13020) );
  NAND2_X1 U16366 ( .A1(n13021), .A2(n13020), .ZN(n15585) );
  INV_X1 U16367 ( .A(n15585), .ZN(n13024) );
  INV_X1 U16368 ( .A(n13023), .ZN(n13022) );
  OR2_X1 U16369 ( .A1(n13022), .A2(n15585), .ZN(n13045) );
  OAI211_X1 U16370 ( .C1(n13023), .C2(n13024), .A(n13750), .B(n13045), .ZN(
        n15584) );
  INV_X1 U16371 ( .A(n15594), .ZN(n13025) );
  NAND2_X1 U16372 ( .A1(n13025), .A2(n13024), .ZN(n13026) );
  INV_X1 U16373 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13030) );
  NAND2_X1 U16374 ( .A1(n13163), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n13029) );
  OAI211_X1 U16375 ( .C1(n13128), .C2(n13030), .A(n13154), .B(n13029), .ZN(
        n13031) );
  INV_X1 U16376 ( .A(n13031), .ZN(n13035) );
  AOI22_X1 U16377 ( .A1(n9686), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13150), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13034) );
  AOI22_X1 U16378 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10358), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13033) );
  AOI22_X1 U16379 ( .A1(n13147), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13032) );
  NAND4_X1 U16380 ( .A1(n13035), .A2(n13034), .A3(n13033), .A4(n13032), .ZN(
        n13044) );
  NAND2_X1 U16381 ( .A1(n13163), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n13036) );
  OAI211_X1 U16382 ( .C1(n13128), .C2(n13037), .A(n13113), .B(n13036), .ZN(
        n13038) );
  INV_X1 U16383 ( .A(n13038), .ZN(n13042) );
  AOI22_X1 U16384 ( .A1(n9686), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13150), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13041) );
  AOI22_X1 U16385 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9665), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13040) );
  AOI22_X1 U16386 ( .A1(n13147), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13039) );
  NAND4_X1 U16387 ( .A1(n13042), .A2(n13041), .A3(n13040), .A4(n13039), .ZN(
        n13043) );
  NAND2_X1 U16388 ( .A1(n13044), .A2(n13043), .ZN(n13047) );
  OR2_X1 U16389 ( .A1(n13045), .A2(n13047), .ZN(n13073) );
  NAND2_X1 U16390 ( .A1(n13045), .A2(n13047), .ZN(n13046) );
  NAND3_X1 U16391 ( .A1(n13073), .A2(n13750), .A3(n13046), .ZN(n13050) );
  INV_X1 U16392 ( .A(n13047), .ZN(n13048) );
  NAND2_X1 U16393 ( .A1(n9730), .A2(n13048), .ZN(n15578) );
  NAND2_X1 U16394 ( .A1(n15575), .A2(n13049), .ZN(n15576) );
  INV_X1 U16395 ( .A(n13050), .ZN(n13051) );
  NAND2_X1 U16396 ( .A1(n13052), .A2(n13051), .ZN(n13053) );
  INV_X1 U16397 ( .A(n13073), .ZN(n13070) );
  AOI22_X1 U16398 ( .A1(n9686), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n9737), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13059) );
  OAI21_X1 U16399 ( .B1(n13132), .B2(n13054), .A(n13154), .ZN(n13055) );
  AOI21_X1 U16400 ( .B1(n13162), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n13055), .ZN(n13058) );
  AOI22_X1 U16401 ( .A1(n13147), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13057) );
  AOI22_X1 U16402 ( .A1(n14000), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n13090), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13056) );
  NAND4_X1 U16403 ( .A1(n13059), .A2(n13058), .A3(n13057), .A4(n13056), .ZN(
        n13069) );
  OR2_X1 U16404 ( .A1(n13156), .A2(n13060), .ZN(n13061) );
  OAI211_X1 U16405 ( .C1(n13128), .C2(n13062), .A(n13113), .B(n13061), .ZN(
        n13063) );
  INV_X1 U16406 ( .A(n13063), .ZN(n13067) );
  AOI22_X1 U16407 ( .A1(n9686), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13150), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13066) );
  AOI22_X1 U16408 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10358), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13065) );
  AOI22_X1 U16409 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13163), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13064) );
  NAND4_X1 U16410 ( .A1(n13067), .A2(n13066), .A3(n13065), .A4(n13064), .ZN(
        n13068) );
  AND2_X1 U16411 ( .A1(n13069), .A2(n13068), .ZN(n13071) );
  NAND2_X1 U16412 ( .A1(n13070), .A2(n13071), .ZN(n13079) );
  INV_X1 U16413 ( .A(n13071), .ZN(n13076) );
  INV_X1 U16414 ( .A(n13750), .ZN(n13072) );
  AOI21_X1 U16415 ( .B1(n13073), .B2(n13076), .A(n13072), .ZN(n13074) );
  NAND2_X1 U16416 ( .A1(n13079), .A2(n13074), .ZN(n13078) );
  INV_X1 U16417 ( .A(n13078), .ZN(n13075) );
  NOR2_X1 U16418 ( .A1(n15586), .A2(n13076), .ZN(n15568) );
  INV_X1 U16419 ( .A(n13079), .ZN(n13098) );
  INV_X1 U16420 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13081) );
  NAND2_X1 U16421 ( .A1(n13163), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n13080) );
  OAI211_X1 U16422 ( .C1(n13128), .C2(n13081), .A(n13154), .B(n13080), .ZN(
        n13082) );
  INV_X1 U16423 ( .A(n13082), .ZN(n13086) );
  AOI22_X1 U16424 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n13150), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13085) );
  AOI22_X1 U16425 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10358), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13084) );
  AOI22_X1 U16426 ( .A1(n13147), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13083) );
  NAND4_X1 U16427 ( .A1(n13086), .A2(n13085), .A3(n13084), .A4(n13083), .ZN(
        n13097) );
  INV_X1 U16428 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13088) );
  NAND2_X1 U16429 ( .A1(n13163), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n13087) );
  OAI211_X1 U16430 ( .C1(n13128), .C2(n13088), .A(n13113), .B(n13087), .ZN(
        n13089) );
  INV_X1 U16431 ( .A(n13089), .ZN(n13095) );
  AOI22_X1 U16432 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13150), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13094) );
  AOI22_X1 U16433 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9665), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13093) );
  AOI22_X1 U16434 ( .A1(n13147), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13092) );
  NAND4_X1 U16435 ( .A1(n13095), .A2(n13094), .A3(n13093), .A4(n13092), .ZN(
        n13096) );
  AND2_X1 U16436 ( .A1(n13097), .A2(n13096), .ZN(n13100) );
  NAND2_X1 U16437 ( .A1(n13098), .A2(n13100), .ZN(n15550) );
  OAI211_X1 U16438 ( .C1(n13098), .C2(n13100), .A(n13750), .B(n15550), .ZN(
        n13102) );
  INV_X1 U16439 ( .A(n13102), .ZN(n13099) );
  NAND2_X1 U16440 ( .A1(n9730), .A2(n13100), .ZN(n15558) );
  INV_X1 U16441 ( .A(n13101), .ZN(n13103) );
  NOR2_X2 U16442 ( .A1(n13103), .A2(n13102), .ZN(n15552) );
  OAI21_X1 U16443 ( .B1(n13156), .B2(n13104), .A(n13154), .ZN(n13109) );
  OAI22_X1 U16444 ( .A1(n13159), .A2(n13107), .B1(n13106), .B2(n13105), .ZN(
        n13108) );
  AOI211_X1 U16445 ( .C1(n13162), .C2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n13109), .B(n13108), .ZN(n13112) );
  AOI22_X1 U16446 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13163), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13111) );
  AOI22_X1 U16447 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n13150), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13110) );
  NAND3_X1 U16448 ( .A1(n13112), .A2(n13111), .A3(n13110), .ZN(n13124) );
  OAI21_X1 U16449 ( .B1(n13156), .B2(n13114), .A(n13113), .ZN(n13119) );
  OAI22_X1 U16450 ( .A1(n13128), .A2(n13117), .B1(n13115), .B2(n13116), .ZN(
        n13118) );
  AOI211_X1 U16451 ( .C1(n9737), .C2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A(
        n13119), .B(n13118), .ZN(n13122) );
  AOI22_X1 U16452 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13163), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13121) );
  AOI22_X1 U16453 ( .A1(n9686), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10358), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13120) );
  NAND3_X1 U16454 ( .A1(n13122), .A2(n13121), .A3(n13120), .ZN(n13123) );
  AND2_X1 U16455 ( .A1(n13124), .A2(n13123), .ZN(n13142) );
  AOI22_X1 U16456 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9665), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13126) );
  AOI21_X1 U16457 ( .B1(n13163), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A(
        n13154), .ZN(n13125) );
  OAI211_X1 U16458 ( .C1(n13128), .C2(n13127), .A(n13126), .B(n13125), .ZN(
        n13141) );
  AOI22_X1 U16459 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n13150), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13130) );
  AOI22_X1 U16460 ( .A1(n13147), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13129) );
  NAND2_X1 U16461 ( .A1(n13130), .A2(n13129), .ZN(n13140) );
  OAI21_X1 U16462 ( .B1(n13132), .B2(n13131), .A(n13154), .ZN(n13133) );
  AOI21_X1 U16463 ( .B1(n13162), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n13133), .ZN(n13138) );
  AOI22_X1 U16464 ( .A1(n13147), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13137) );
  AOI22_X1 U16465 ( .A1(n9686), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13150), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13136) );
  AOI22_X1 U16466 ( .A1(n13091), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13090), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13135) );
  NAND4_X1 U16467 ( .A1(n13138), .A2(n13137), .A3(n13136), .A4(n13135), .ZN(
        n13139) );
  OAI21_X1 U16468 ( .B1(n13141), .B2(n13140), .A(n13139), .ZN(n13144) );
  INV_X1 U16469 ( .A(n13142), .ZN(n15553) );
  NOR3_X1 U16470 ( .A1(n15550), .A2(n9730), .A3(n15553), .ZN(n13143) );
  XOR2_X1 U16471 ( .A(n13144), .B(n13143), .Z(n15547) );
  INV_X1 U16472 ( .A(n13143), .ZN(n13145) );
  AOI22_X1 U16473 ( .A1(n12982), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13162), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13149) );
  AOI22_X1 U16474 ( .A1(n13147), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13146), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13148) );
  NAND2_X1 U16475 ( .A1(n13149), .A2(n13148), .ZN(n13169) );
  INV_X1 U16476 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13153) );
  AOI22_X1 U16477 ( .A1(n13150), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10358), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13152) );
  AOI21_X1 U16478 ( .B1(n13163), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n13154), .ZN(n13151) );
  OAI211_X1 U16479 ( .C1(n13159), .C2(n13153), .A(n13152), .B(n13151), .ZN(
        n13168) );
  INV_X1 U16480 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13155) );
  OAI21_X1 U16481 ( .B1(n13156), .B2(n13155), .A(n13154), .ZN(n13161) );
  INV_X1 U16482 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13158) );
  INV_X1 U16483 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13157) );
  OAI22_X1 U16484 ( .A1(n13159), .A2(n13158), .B1(n13115), .B2(n13157), .ZN(
        n13160) );
  AOI211_X1 U16485 ( .C1(n13162), .C2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n13161), .B(n13160), .ZN(n13166) );
  AOI22_X1 U16486 ( .A1(n13146), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13163), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13165) );
  AOI22_X1 U16487 ( .A1(n9686), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n9665), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13164) );
  NAND3_X1 U16488 ( .A1(n13166), .A2(n13165), .A3(n13164), .ZN(n13167) );
  OAI21_X1 U16489 ( .B1(n13169), .B2(n13168), .A(n13167), .ZN(n13170) );
  NAND2_X1 U16490 ( .A1(n11353), .A2(n20221), .ZN(n14030) );
  NAND2_X1 U16491 ( .A1(n13408), .A2(n14020), .ZN(n14033) );
  OAI22_X1 U16492 ( .A1(n14310), .A2(n13999), .B1(n14030), .B2(n14033), .ZN(
        n13524) );
  AND2_X1 U16493 ( .A1(n13173), .A2(n13172), .ZN(n13174) );
  NAND2_X1 U16494 ( .A1(n13339), .A2(n13177), .ZN(n13197) );
  NOR4_X1 U16495 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n13181) );
  NOR4_X1 U16496 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n13180) );
  NOR4_X1 U16497 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n13179) );
  NOR4_X1 U16498 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n13178) );
  NAND4_X1 U16499 ( .A1(n13181), .A2(n13180), .A3(n13179), .A4(n13178), .ZN(
        n13186) );
  NOR4_X1 U16500 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n13184) );
  NOR4_X1 U16501 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n13183) );
  NOR4_X1 U16502 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n13182) );
  INV_X1 U16503 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n20106) );
  NAND4_X1 U16504 ( .A1(n13184), .A2(n13183), .A3(n13182), .A4(n20106), .ZN(
        n13185) );
  NAND2_X1 U16505 ( .A1(n13187), .A2(n13498), .ZN(n13188) );
  OR2_X1 U16506 ( .A1(n19462), .A2(n13338), .ZN(n15675) );
  INV_X1 U16507 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13190) );
  OAI22_X1 U16508 ( .A1(n15675), .A2(n13189), .B1(n15689), .B2(n13190), .ZN(
        n13191) );
  AOI21_X1 U16509 ( .B1(n19450), .B2(BUF2_REG_30__SCAN_IN), .A(n13191), .ZN(
        n13195) );
  NOR3_X2 U16510 ( .A1(n19462), .A2(n19519), .A3(n13192), .ZN(n19451) );
  NAND2_X1 U16511 ( .A1(n19551), .A2(n13338), .ZN(n13193) );
  INV_X1 U16512 ( .A(n15690), .ZN(n16572) );
  MUX2_X1 U16513 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n19519), .Z(n19455) );
  AOI22_X1 U16514 ( .A1(n19451), .A2(BUF1_REG_30__SCAN_IN), .B1(n16572), .B2(
        n19455), .ZN(n13194) );
  NAND2_X1 U16515 ( .A1(n13197), .A2(n13196), .ZN(P2_U2889) );
  NAND2_X1 U16516 ( .A1(n13199), .A2(n13198), .ZN(n16022) );
  INV_X1 U16517 ( .A(n16024), .ZN(n13200) );
  NAND2_X1 U16518 ( .A1(n16022), .A2(n13200), .ZN(n13201) );
  NAND2_X1 U16519 ( .A1(n13201), .A2(n16023), .ZN(n16599) );
  AND2_X1 U16520 ( .A1(n13203), .A2(n13202), .ZN(n16601) );
  INV_X1 U16521 ( .A(n15989), .ZN(n13205) );
  NAND2_X1 U16522 ( .A1(n13205), .A2(n15987), .ZN(n13206) );
  INV_X1 U16523 ( .A(n13207), .ZN(n15819) );
  NAND2_X1 U16524 ( .A1(n15810), .A2(n13210), .ZN(n15799) );
  INV_X1 U16525 ( .A(n13211), .ZN(n15801) );
  INV_X1 U16526 ( .A(n15791), .ZN(n13212) );
  OAI21_X1 U16527 ( .B1(n15688), .B2(n13216), .A(n15673), .ZN(n13217) );
  INV_X1 U16528 ( .A(n13217), .ZN(n19242) );
  NOR3_X1 U16529 ( .A1(n15944), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n13218), .ZN(n13227) );
  NAND2_X1 U16530 ( .A1(n19500), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n14668) );
  NOR2_X1 U16531 ( .A1(n13220), .A2(n13221), .ZN(n13222) );
  OR2_X1 U16532 ( .A1(n13219), .A2(n13222), .ZN(n15610) );
  INV_X1 U16533 ( .A(n15610), .ZN(n19240) );
  NAND2_X1 U16534 ( .A1(n19240), .A2(n16699), .ZN(n13223) );
  OAI211_X1 U16535 ( .C1(n13225), .C2(n13224), .A(n14668), .B(n13223), .ZN(
        n13226) );
  AOI211_X1 U16536 ( .C1(n19242), .C2(n16710), .A(n13227), .B(n13226), .ZN(
        n13228) );
  INV_X1 U16537 ( .A(n13228), .ZN(n13231) );
  NOR2_X1 U16538 ( .A1(n15783), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n14671) );
  OAI21_X1 U16539 ( .B1(n14675), .B2(n16704), .A(n13232), .ZN(P2_U3025) );
  INV_X1 U16540 ( .A(n13291), .ZN(n13235) );
  NAND2_X1 U16541 ( .A1(n11941), .A2(n11891), .ZN(n13247) );
  OAI21_X1 U16542 ( .B1(n13658), .B2(n13238), .A(n13247), .ZN(n13233) );
  INV_X1 U16543 ( .A(n13233), .ZN(n13234) );
  NAND2_X1 U16544 ( .A1(n13239), .A2(n13238), .ZN(n13256) );
  OAI21_X1 U16545 ( .B1(n13239), .B2(n13238), .A(n13256), .ZN(n13240) );
  OAI211_X1 U16546 ( .C1(n13240), .C2(n13658), .A(n12770), .B(n12589), .ZN(
        n13241) );
  INV_X1 U16547 ( .A(n13241), .ZN(n13242) );
  INV_X1 U16548 ( .A(n13243), .ZN(n13244) );
  NAND2_X1 U16549 ( .A1(n13246), .A2(n13291), .ZN(n13251) );
  XNOR2_X1 U16550 ( .A(n13256), .B(n13255), .ZN(n13249) );
  INV_X1 U16551 ( .A(n13247), .ZN(n13248) );
  AOI21_X1 U16552 ( .B1(n13249), .B2(n21019), .A(n13248), .ZN(n13250) );
  NAND2_X1 U16553 ( .A1(n13251), .A2(n13250), .ZN(n13896) );
  NAND2_X1 U16554 ( .A1(n13252), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13253) );
  NAND2_X1 U16555 ( .A1(n13256), .A2(n13255), .ZN(n13272) );
  XNOR2_X1 U16556 ( .A(n13272), .B(n13270), .ZN(n13257) );
  OAI22_X1 U16557 ( .A1(n13254), .A2(n13235), .B1(n13658), .B2(n13257), .ZN(
        n13961) );
  NAND2_X1 U16558 ( .A1(n13962), .A2(n13961), .ZN(n13960) );
  NAND2_X1 U16559 ( .A1(n13258), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13259) );
  NAND2_X1 U16560 ( .A1(n13960), .A2(n13259), .ZN(n20418) );
  NAND2_X1 U16561 ( .A1(n13260), .A2(n13291), .ZN(n13264) );
  NAND2_X1 U16562 ( .A1(n13272), .A2(n13270), .ZN(n13261) );
  XNOR2_X1 U16563 ( .A(n13261), .B(n13269), .ZN(n13262) );
  NAND2_X1 U16564 ( .A1(n13262), .A2(n21019), .ZN(n13263) );
  NAND2_X1 U16565 ( .A1(n13264), .A2(n13263), .ZN(n13265) );
  INV_X1 U16566 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20438) );
  XNOR2_X1 U16567 ( .A(n13265), .B(n20438), .ZN(n20417) );
  NAND2_X1 U16568 ( .A1(n13265), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13266) );
  INV_X1 U16569 ( .A(n13267), .ZN(n13268) );
  OR2_X1 U16570 ( .A1(n13268), .A2(n13235), .ZN(n13275) );
  AND2_X1 U16571 ( .A1(n13270), .A2(n13269), .ZN(n13271) );
  NAND2_X1 U16572 ( .A1(n13272), .A2(n13271), .ZN(n13281) );
  XNOR2_X1 U16573 ( .A(n13281), .B(n13279), .ZN(n13273) );
  NAND2_X1 U16574 ( .A1(n13273), .A2(n21019), .ZN(n13274) );
  NAND2_X1 U16575 ( .A1(n13275), .A2(n13274), .ZN(n13276) );
  XNOR2_X1 U16576 ( .A(n13276), .B(n16447), .ZN(n16380) );
  NAND2_X1 U16577 ( .A1(n13276), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13277) );
  NAND3_X1 U16578 ( .A1(n13298), .A2(n13278), .A3(n13291), .ZN(n13284) );
  INV_X1 U16579 ( .A(n13279), .ZN(n13280) );
  OR2_X1 U16580 ( .A1(n13281), .A2(n13280), .ZN(n13286) );
  XNOR2_X1 U16581 ( .A(n13286), .B(n13287), .ZN(n13282) );
  NAND2_X1 U16582 ( .A1(n13282), .A2(n21019), .ZN(n13283) );
  NAND2_X1 U16583 ( .A1(n13284), .A2(n13283), .ZN(n16375) );
  OR2_X1 U16584 ( .A1(n16375), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13285) );
  INV_X1 U16585 ( .A(n13286), .ZN(n13288) );
  NAND2_X1 U16586 ( .A1(n13288), .A2(n13287), .ZN(n13299) );
  XNOR2_X1 U16587 ( .A(n13299), .B(n13300), .ZN(n13289) );
  AND2_X1 U16588 ( .A1(n13289), .A2(n21019), .ZN(n13290) );
  AOI21_X1 U16589 ( .B1(n13292), .B2(n13291), .A(n13290), .ZN(n13293) );
  NAND2_X1 U16590 ( .A1(n13293), .A2(n16439), .ZN(n16370) );
  NAND2_X1 U16591 ( .A1(n16368), .A2(n16370), .ZN(n13295) );
  INV_X1 U16592 ( .A(n13293), .ZN(n13294) );
  NAND2_X1 U16593 ( .A1(n13294), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16369) );
  NOR2_X1 U16594 ( .A1(n13296), .A2(n13235), .ZN(n13297) );
  INV_X1 U16595 ( .A(n13299), .ZN(n13301) );
  NAND3_X1 U16596 ( .A1(n13301), .A2(n21019), .A3(n13300), .ZN(n13302) );
  NAND2_X1 U16597 ( .A1(n15449), .A2(n13302), .ZN(n14477) );
  OR2_X1 U16598 ( .A1(n14477), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13303) );
  NAND2_X1 U16599 ( .A1(n14477), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13304) );
  NAND2_X1 U16600 ( .A1(n9674), .A2(n16420), .ZN(n13305) );
  NAND2_X1 U16601 ( .A1(n9673), .A2(n15413), .ZN(n13306) );
  INV_X1 U16602 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15481) );
  NAND2_X1 U16603 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13307) );
  NAND2_X1 U16604 ( .A1(n15449), .A2(n13307), .ZN(n15444) );
  INV_X1 U16605 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15456) );
  NAND2_X1 U16606 ( .A1(n15449), .A2(n15456), .ZN(n13308) );
  AND2_X1 U16607 ( .A1(n15444), .A2(n13308), .ZN(n13309) );
  NAND2_X1 U16608 ( .A1(n15445), .A2(n13309), .ZN(n15244) );
  OR2_X1 U16609 ( .A1(n9674), .A2(n15456), .ZN(n13310) );
  AND2_X1 U16610 ( .A1(n15447), .A2(n13310), .ZN(n13314) );
  AND2_X1 U16611 ( .A1(n13314), .A2(n15248), .ZN(n15232) );
  OR2_X1 U16612 ( .A1(n9674), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15236) );
  NAND2_X1 U16613 ( .A1(n9674), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13311) );
  NAND2_X1 U16614 ( .A1(n15236), .A2(n13311), .ZN(n15435) );
  NAND2_X1 U16615 ( .A1(n15449), .A2(n16393), .ZN(n15433) );
  NAND2_X1 U16616 ( .A1(n15435), .A2(n15433), .ZN(n13312) );
  NOR3_X1 U16617 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13313) );
  NAND2_X1 U16618 ( .A1(n13314), .A2(n15231), .ZN(n15245) );
  XNOR2_X1 U16619 ( .A(n9673), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15224) );
  NAND3_X1 U16620 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14728) );
  INV_X1 U16621 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15368) );
  NAND4_X1 U16622 ( .A1(n13316), .A2(n15419), .A3(n15368), .A4(n15401), .ZN(
        n13317) );
  AND2_X1 U16623 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15325) );
  NAND2_X1 U16624 ( .A1(n15325), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15132) );
  NAND2_X1 U16625 ( .A1(n15131), .A2(n15132), .ZN(n13319) );
  NAND2_X1 U16626 ( .A1(n13318), .A2(n15449), .ZN(n15160) );
  NAND3_X1 U16627 ( .A1(n13319), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15160), .ZN(n15147) );
  NAND3_X1 U16628 ( .A1(n15343), .A2(n15324), .A3(n15346), .ZN(n15133) );
  AND2_X1 U16629 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15293) );
  MUX2_X1 U16630 ( .A(n14707), .B(n9768), .S(n9674), .Z(n13320) );
  XNOR2_X1 U16631 ( .A(n13320), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15301) );
  AOI21_X1 U16632 ( .B1(n11897), .B2(n11941), .A(n13321), .ZN(n13322) );
  NAND2_X1 U16633 ( .A1(n13546), .A2(n13322), .ZN(n13572) );
  OR2_X1 U16634 ( .A1(n13572), .A2(n13323), .ZN(n13693) );
  NOR2_X2 U16635 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20811) );
  NAND2_X1 U16636 ( .A1(n20880), .A2(n13324), .ZN(n21026) );
  AND2_X1 U16637 ( .A1(n21026), .A2(n21023), .ZN(n13325) );
  NAND2_X1 U16638 ( .A1(n21023), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13327) );
  NAND2_X1 U16639 ( .A1(n21170), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13326) );
  NAND2_X1 U16640 ( .A1(n13327), .A2(n13326), .ZN(n13717) );
  OR2_X1 U16641 ( .A1(n20432), .A2(n21096), .ZN(n15295) );
  OAI21_X1 U16642 ( .B1(n15254), .B2(n13328), .A(n15295), .ZN(n13329) );
  AOI21_X1 U16643 ( .B1(n16355), .B2(n14692), .A(n13329), .ZN(n13334) );
  NAND3_X1 U16644 ( .A1(n21023), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16462) );
  INV_X1 U16645 ( .A(n16462), .ZN(n13333) );
  AND2_X2 U16646 ( .A1(n13333), .A2(n20811), .ZN(n16364) );
  INV_X1 U16647 ( .A(n16364), .ZN(n15258) );
  NAND2_X1 U16648 ( .A1(n14310), .A2(n13335), .ZN(n13522) );
  NAND2_X1 U16649 ( .A1(n13522), .A2(n13997), .ZN(n13337) );
  NAND2_X1 U16650 ( .A1(n13339), .A2(n14786), .ZN(n13343) );
  NAND2_X1 U16651 ( .A1(n13835), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13340) );
  NAND2_X1 U16652 ( .A1(n13343), .A2(n13342), .ZN(P2_U2857) );
  NOR2_X1 U16653 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13345) );
  NOR4_X1 U16654 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13344) );
  NAND4_X1 U16655 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13345), .A4(n13344), .ZN(n13358) );
  NOR4_X1 U16656 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13349) );
  NOR4_X1 U16657 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n13348) );
  NOR4_X1 U16658 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13347) );
  NOR4_X1 U16659 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n13346) );
  AND4_X1 U16660 ( .A1(n13349), .A2(n13348), .A3(n13347), .A4(n13346), .ZN(
        n13354) );
  NOR4_X1 U16661 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13352) );
  NOR4_X1 U16662 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13351) );
  NOR4_X1 U16663 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13350) );
  INV_X1 U16664 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20964) );
  AND4_X1 U16665 ( .A1(n13352), .A2(n13351), .A3(n13350), .A4(n20964), .ZN(
        n13353) );
  NAND2_X1 U16666 ( .A1(n13354), .A2(n13353), .ZN(n13355) );
  INV_X1 U16667 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n21092) );
  NOR3_X1 U16668 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        n21092), .ZN(n13357) );
  NOR4_X1 U16669 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(P1_BE_N_REG_2__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n13356)
         );
  NAND4_X1 U16670 ( .A1(n14699), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13357), .A4(
        n13356), .ZN(U214) );
  NOR2_X1 U16671 ( .A1(n13498), .A2(n13358), .ZN(n16747) );
  NAND2_X1 U16672 ( .A1(n16747), .A2(U214), .ZN(U212) );
  INV_X1 U16673 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n13366) );
  NAND2_X1 U16674 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n13359), .ZN(
        n17905) );
  NOR2_X1 U16675 ( .A1(n13366), .A2(n17905), .ZN(n13385) );
  AOI21_X1 U16676 ( .B1(n13366), .B2(n17905), .A(n13385), .ZN(n17933) );
  INV_X1 U16677 ( .A(n13360), .ZN(n17981) );
  NOR2_X1 U16678 ( .A1(n18169), .A2(n18006), .ZN(n17084) );
  NAND2_X1 U16679 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n17084), .ZN(
        n18018) );
  NOR2_X1 U16680 ( .A1(n17981), .A2(n18018), .ZN(n17978) );
  NAND2_X1 U16681 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17978), .ZN(
        n17028) );
  NOR2_X1 U16682 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17028), .ZN(
        n17005) );
  NOR2_X1 U16683 ( .A1(n18169), .A2(n13361), .ZN(n17940) );
  NAND2_X1 U16684 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17940), .ZN(
        n16993) );
  INV_X1 U16685 ( .A(n16993), .ZN(n16983) );
  NOR3_X1 U16686 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(P3_STATEBS16_REG_SCAN_IN), .ZN(n19048) );
  NAND2_X1 U16687 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n19048), .ZN(n17176) );
  AOI211_X1 U16688 ( .C1(n17933), .C2(n13362), .A(n13386), .B(n17176), .ZN(
        n13374) );
  NOR3_X1 U16689 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17188) );
  INV_X1 U16690 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17527) );
  NAND2_X1 U16691 ( .A1(n17188), .A2(n17527), .ZN(n17185) );
  NOR2_X1 U16692 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17185), .ZN(n17166) );
  NAND2_X1 U16693 ( .A1(n17166), .A2(n17532), .ZN(n17151) );
  INV_X1 U16694 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17126) );
  NAND2_X1 U16695 ( .A1(n17134), .A2(n17126), .ZN(n17124) );
  INV_X1 U16696 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17104) );
  NAND2_X1 U16697 ( .A1(n17109), .A2(n17104), .ZN(n17103) );
  INV_X1 U16698 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17083) );
  NAND2_X1 U16699 ( .A1(n17087), .A2(n17083), .ZN(n17080) );
  INV_X1 U16700 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n17395) );
  NAND2_X1 U16701 ( .A1(n17061), .A2(n17395), .ZN(n17055) );
  INV_X1 U16702 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n17397) );
  NAND2_X1 U16703 ( .A1(n17038), .A2(n17397), .ZN(n17034) );
  INV_X1 U16704 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17013) );
  NAND2_X1 U16705 ( .A1(n17019), .A2(n17013), .ZN(n17011) );
  INV_X1 U16706 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16989) );
  NAND2_X1 U16707 ( .A1(n16996), .A2(n16989), .ZN(n16988) );
  NAND2_X1 U16708 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n9725), .ZN(n13365) );
  AOI211_X4 U16709 ( .C1(n19185), .C2(n19187), .A(n19200), .B(n13365), .ZN(
        n17219) );
  AOI211_X1 U16710 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16988), .A(n16972), .B(
        n17216), .ZN(n13373) );
  INV_X1 U16711 ( .A(n19033), .ZN(n19041) );
  NOR2_X2 U16712 ( .A1(n19138), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n19042) );
  INV_X1 U16713 ( .A(n19042), .ZN(n18795) );
  NOR2_X1 U16714 ( .A1(n18499), .A2(n19045), .ZN(n17172) );
  INV_X1 U16715 ( .A(n19187), .ZN(n19182) );
  AOI211_X1 U16716 ( .C1(n19186), .C2(n19184), .A(n19182), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n13367) );
  AOI211_X4 U16717 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n9725), .A(n13367), .B(
        n19200), .ZN(n17220) );
  INV_X1 U16718 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17226) );
  OAI22_X1 U16719 ( .A1(n13366), .A2(n17206), .B1(n17209), .B2(n17226), .ZN(
        n13372) );
  NAND2_X1 U16720 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n13368) );
  NAND3_X1 U16721 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16981) );
  INV_X1 U16722 ( .A(n13367), .ZN(n19027) );
  INV_X1 U16723 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n19093) );
  INV_X1 U16724 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n19088) );
  INV_X1 U16725 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n19084) );
  INV_X1 U16726 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n19080) );
  INV_X1 U16727 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n19072) );
  NAND3_X1 U16728 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n17164) );
  NOR2_X1 U16729 ( .A1(n19072), .A2(n17164), .ZN(n17145) );
  NAND2_X1 U16730 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n17145), .ZN(n17122) );
  INV_X1 U16731 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n19078) );
  INV_X1 U16732 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n19076) );
  NOR2_X1 U16733 ( .A1(n19078), .A2(n19076), .ZN(n17123) );
  INV_X1 U16734 ( .A(n17123), .ZN(n17114) );
  NOR3_X1 U16735 ( .A1(n19080), .A2(n17122), .A3(n17114), .ZN(n17089) );
  NAND2_X1 U16736 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n17089), .ZN(n17091) );
  NOR2_X1 U16737 ( .A1(n19084), .A2(n17091), .ZN(n17073) );
  NAND2_X1 U16738 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n17073), .ZN(n17067) );
  NOR2_X1 U16739 ( .A1(n19088), .A2(n17067), .ZN(n17056) );
  NAND2_X1 U16740 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n17056), .ZN(n17040) );
  INV_X1 U16741 ( .A(n17033), .ZN(n17021) );
  NOR2_X1 U16742 ( .A1(n16981), .A2(n17021), .ZN(n17000) );
  INV_X1 U16743 ( .A(n17000), .ZN(n16982) );
  NOR2_X1 U16744 ( .A1(n13368), .A2(n16982), .ZN(n13370) );
  NOR2_X1 U16745 ( .A1(n19093), .A2(n17040), .ZN(n16980) );
  INV_X1 U16746 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n19104) );
  NOR3_X1 U16747 ( .A1(n19104), .A2(n16981), .A3(n13368), .ZN(n13400) );
  NAND2_X1 U16748 ( .A1(n16980), .A2(n13400), .ZN(n13376) );
  AOI21_X1 U16749 ( .B1(n17165), .B2(n13376), .A(n17204), .ZN(n16978) );
  INV_X1 U16750 ( .A(n16978), .ZN(n13369) );
  MUX2_X1 U16751 ( .A(n13370), .B(n13369), .S(P3_REIP_REG_20__SCAN_IN), .Z(
        n13371) );
  OR4_X1 U16752 ( .A1(n13374), .A2(n13373), .A3(n13372), .A4(n13371), .ZN(
        P3_U2651) );
  INV_X1 U16753 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16952) );
  INV_X1 U16754 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16974) );
  NAND2_X1 U16755 ( .A1(n16972), .A2(n16974), .ZN(n16971) );
  INV_X1 U16756 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16963) );
  NAND2_X1 U16757 ( .A1(n16964), .A2(n16963), .ZN(n16962) );
  NAND2_X1 U16758 ( .A1(n16952), .A2(n16953), .ZN(n16936) );
  INV_X1 U16759 ( .A(n16936), .ZN(n16935) );
  INV_X1 U16760 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n17228) );
  NAND2_X1 U16761 ( .A1(n16935), .A2(n17228), .ZN(n13375) );
  NOR2_X1 U16762 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n13375), .ZN(n16927) );
  AOI211_X1 U16763 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n13375), .A(n16927), .B(
        n17216), .ZN(n13396) );
  INV_X1 U16764 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n19116) );
  INV_X1 U16765 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n19112) );
  INV_X1 U16766 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n19107) );
  INV_X1 U16767 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n19108) );
  NOR3_X1 U16768 ( .A1(n19107), .A2(n19108), .A3(n13376), .ZN(n16958) );
  NAND2_X1 U16769 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16958), .ZN(n13377) );
  NOR3_X1 U16770 ( .A1(n19112), .A2(n17210), .A3(n13377), .ZN(n16931) );
  NAND2_X1 U16771 ( .A1(P3_REIP_REG_25__SCAN_IN), .A2(n16931), .ZN(n16872) );
  NOR2_X1 U16772 ( .A1(n17165), .A2(n17204), .ZN(n17010) );
  INV_X1 U16773 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n19114) );
  NOR3_X1 U16774 ( .A1(n19116), .A2(n19114), .A3(n19112), .ZN(n13378) );
  INV_X1 U16775 ( .A(n13377), .ZN(n16949) );
  OAI21_X1 U16776 ( .B1(n17210), .B2(n16949), .A(n17221), .ZN(n16932) );
  INV_X1 U16777 ( .A(n16932), .ZN(n16967) );
  OAI21_X1 U16778 ( .B1(n17010), .B2(n13378), .A(n16967), .ZN(n16879) );
  INV_X1 U16779 ( .A(n16879), .ZN(n16922) );
  AOI21_X1 U16780 ( .B1(n19116), .B2(n16872), .A(n16922), .ZN(n13395) );
  INV_X1 U16781 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13392) );
  AOI21_X1 U16782 ( .B1(n13392), .B2(n13380), .A(n13379), .ZN(n17846) );
  INV_X1 U16783 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17874) );
  NOR2_X1 U16784 ( .A1(n17874), .A2(n13387), .ZN(n13381) );
  OAI21_X1 U16785 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n13381), .A(
        n13380), .ZN(n17860) );
  INV_X1 U16786 ( .A(n17860), .ZN(n16938) );
  INV_X1 U16787 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17893) );
  NAND2_X1 U16788 ( .A1(n13382), .A2(n13385), .ZN(n17891) );
  AOI21_X1 U16789 ( .B1(n17893), .B2(n17891), .A(n13388), .ZN(n17885) );
  NAND2_X1 U16790 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n13385), .ZN(
        n13384) );
  INV_X1 U16791 ( .A(n17891), .ZN(n13383) );
  AOI21_X1 U16792 ( .B1(n13399), .B2(n13384), .A(n13383), .ZN(n17906) );
  OAI21_X1 U16793 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n13385), .A(
        n13384), .ZN(n17915) );
  INV_X1 U16794 ( .A(n17915), .ZN(n16970) );
  NOR2_X1 U16795 ( .A1(n17906), .A2(n13398), .ZN(n13397) );
  NOR2_X1 U16796 ( .A1(n13397), .A2(n17175), .ZN(n16957) );
  NOR2_X1 U16797 ( .A1(n17885), .A2(n16957), .ZN(n16956) );
  NOR2_X1 U16798 ( .A1(n16956), .A2(n17175), .ZN(n16946) );
  INV_X1 U16799 ( .A(n16946), .ZN(n13390) );
  OAI22_X1 U16800 ( .A1(n17874), .A2(n13388), .B1(n13387), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17870) );
  INV_X1 U16801 ( .A(n17870), .ZN(n13389) );
  NAND2_X1 U16802 ( .A1(n13390), .A2(n13389), .ZN(n16944) );
  AOI211_X1 U16803 ( .C1(n17846), .C2(n13391), .A(n16877), .B(n17176), .ZN(
        n13394) );
  INV_X1 U16804 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17280) );
  OAI22_X1 U16805 ( .A1(n13392), .A2(n17206), .B1(n17209), .B2(n17280), .ZN(
        n13393) );
  OR4_X1 U16806 ( .A1(n13396), .A2(n13395), .A3(n13394), .A4(n13393), .ZN(
        P3_U2645) );
  AOI211_X1 U16807 ( .C1(n17906), .C2(n13398), .A(n13397), .B(n17176), .ZN(
        n13405) );
  AOI211_X1 U16808 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16971), .A(n16964), .B(
        n17216), .ZN(n13404) );
  INV_X1 U16809 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16096) );
  OAI22_X1 U16810 ( .A1(n13399), .A2(n17206), .B1(n17209), .B2(n16096), .ZN(
        n13403) );
  NAND2_X1 U16811 ( .A1(n13400), .A2(n17033), .ZN(n16979) );
  XOR2_X1 U16812 ( .A(P3_REIP_REG_22__SCAN_IN), .B(n19107), .Z(n13401) );
  OAI22_X1 U16813 ( .A1(n16979), .A2(n13401), .B1(n19108), .B2(n16978), .ZN(
        n13402) );
  OR4_X1 U16814 ( .A1(n13405), .A2(n13404), .A3(n13403), .A4(n13402), .ZN(
        P3_U2649) );
  NOR2_X1 U16815 ( .A1(n11314), .A2(n19210), .ZN(n13533) );
  NAND2_X1 U16816 ( .A1(n13408), .A2(n13533), .ZN(n14752) );
  INV_X1 U16817 ( .A(n14752), .ZN(n13411) );
  INV_X1 U16818 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13410) );
  NOR2_X1 U16819 ( .A1(n13406), .A2(n19210), .ZN(n13407) );
  INV_X1 U16820 ( .A(n14191), .ZN(n13415) );
  NOR2_X1 U16821 ( .A1(n20016), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13412) );
  INV_X1 U16822 ( .A(n13412), .ZN(n13409) );
  OAI211_X1 U16823 ( .C1(n13411), .C2(n13410), .A(n13415), .B(n13409), .ZN(
        P2_U2814) );
  INV_X1 U16824 ( .A(n11353), .ZN(n13414) );
  INV_X1 U16825 ( .A(n19208), .ZN(n20213) );
  OAI21_X1 U16826 ( .B1(n13412), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n20213), 
        .ZN(n13413) );
  OAI21_X1 U16827 ( .B1(n13414), .B2(n20213), .A(n13413), .ZN(P2_U3612) );
  NOR3_X2 U16828 ( .A1(n13415), .A2(n9730), .A3(n20215), .ZN(n13500) );
  AOI22_X1 U16829 ( .A1(n19521), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19519), .ZN(n19547) );
  INV_X1 U16830 ( .A(n19547), .ZN(n13416) );
  NAND2_X1 U16831 ( .A1(n13500), .A2(n13416), .ZN(n13497) );
  NAND2_X1 U16832 ( .A1(n13483), .A2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13417) );
  OAI211_X1 U16833 ( .C1(n13534), .C2(n13418), .A(n13497), .B(n13417), .ZN(
        P2_U2956) );
  AOI22_X1 U16834 ( .A1(n19521), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19519), .ZN(n19559) );
  INV_X1 U16835 ( .A(n19559), .ZN(n13419) );
  NAND2_X1 U16836 ( .A1(n13500), .A2(n13419), .ZN(n13505) );
  NAND2_X1 U16837 ( .A1(n13483), .A2(P2_LWORD_REG_6__SCAN_IN), .ZN(n13420) );
  OAI211_X1 U16838 ( .C1(n13534), .C2(n19486), .A(n13505), .B(n13420), .ZN(
        P2_U2973) );
  AOI22_X1 U16839 ( .A1(n19521), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n13498), .ZN(n15661) );
  INV_X1 U16840 ( .A(n15661), .ZN(n13421) );
  NAND2_X1 U16841 ( .A1(n13500), .A2(n13421), .ZN(n13508) );
  NAND2_X1 U16842 ( .A1(n13483), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13422) );
  OAI211_X1 U16843 ( .C1(n13423), .C2(n13534), .A(n13508), .B(n13422), .ZN(
        P2_U2975) );
  AOI22_X1 U16844 ( .A1(n19521), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n19519), .ZN(n15622) );
  INV_X1 U16845 ( .A(n15622), .ZN(n13424) );
  NAND2_X1 U16846 ( .A1(n13500), .A2(n13424), .ZN(n13492) );
  NAND2_X1 U16847 ( .A1(n13483), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13425) );
  OAI211_X1 U16848 ( .C1(n13534), .C2(n13426), .A(n13492), .B(n13425), .ZN(
        P2_U2980) );
  NAND2_X1 U16849 ( .A1(n13500), .A2(n19455), .ZN(n13511) );
  NAND2_X1 U16850 ( .A1(n13483), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13427) );
  OAI211_X1 U16851 ( .C1(n13190), .C2(n13534), .A(n13511), .B(n13427), .ZN(
        P2_U2966) );
  INV_X1 U16852 ( .A(n13483), .ZN(n13456) );
  INV_X1 U16853 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13429) );
  INV_X1 U16854 ( .A(n13500), .ZN(n13454) );
  INV_X1 U16855 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16796) );
  INV_X1 U16856 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18537) );
  OAI22_X1 U16857 ( .A1(n13498), .A2(n16796), .B1(n18537), .B2(n19521), .ZN(
        n19463) );
  INV_X1 U16858 ( .A(n19463), .ZN(n19552) );
  NOR2_X1 U16859 ( .A1(n13454), .A2(n19552), .ZN(n13439) );
  AOI21_X1 U16860 ( .B1(n14195), .B2(P2_EAX_REG_21__SCAN_IN), .A(n13439), .ZN(
        n13428) );
  OAI21_X1 U16861 ( .B1(n13456), .B2(n13429), .A(n13428), .ZN(P2_U2957) );
  INV_X1 U16862 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n13431) );
  OAI22_X1 U16863 ( .A1(n13498), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19521), .ZN(n19533) );
  NOR2_X1 U16864 ( .A1(n13454), .A2(n19533), .ZN(n13450) );
  AOI21_X1 U16865 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n14195), .A(n13450), .ZN(
        n13430) );
  OAI21_X1 U16866 ( .B1(n13456), .B2(n13431), .A(n13430), .ZN(P2_U2968) );
  INV_X1 U16867 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n13433) );
  AOI22_X1 U16868 ( .A1(n19521), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19519), .ZN(n19544) );
  NOR2_X1 U16869 ( .A1(n13454), .A2(n19544), .ZN(n13434) );
  AOI21_X1 U16870 ( .B1(P2_EAX_REG_3__SCAN_IN), .B2(n14195), .A(n13434), .ZN(
        n13432) );
  OAI21_X1 U16871 ( .B1(n13456), .B2(n13433), .A(n13432), .ZN(P2_U2970) );
  INV_X1 U16872 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n13436) );
  AOI21_X1 U16873 ( .B1(n14195), .B2(P2_EAX_REG_19__SCAN_IN), .A(n13434), .ZN(
        n13435) );
  OAI21_X1 U16874 ( .B1(n13456), .B2(n13436), .A(n13435), .ZN(P2_U2955) );
  INV_X1 U16875 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n13438) );
  AOI22_X1 U16876 ( .A1(n19521), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n19519), .ZN(n19567) );
  NOR2_X1 U16877 ( .A1(n13454), .A2(n19567), .ZN(n13444) );
  AOI21_X1 U16878 ( .B1(n14195), .B2(P2_EAX_REG_23__SCAN_IN), .A(n13444), .ZN(
        n13437) );
  OAI21_X1 U16879 ( .B1(n13456), .B2(n13438), .A(n13437), .ZN(P2_U2959) );
  INV_X1 U16880 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n13441) );
  AOI21_X1 U16881 ( .B1(P2_EAX_REG_5__SCAN_IN), .B2(n14195), .A(n13439), .ZN(
        n13440) );
  OAI21_X1 U16882 ( .B1(n13456), .B2(n13441), .A(n13440), .ZN(P2_U2972) );
  INV_X1 U16883 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n13443) );
  AOI22_X1 U16884 ( .A1(n19521), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n13498), .ZN(n15654) );
  NOR2_X1 U16885 ( .A1(n13454), .A2(n15654), .ZN(n13447) );
  AOI21_X1 U16886 ( .B1(n14195), .B2(P2_EAX_REG_9__SCAN_IN), .A(n13447), .ZN(
        n13442) );
  OAI21_X1 U16887 ( .B1(n13456), .B2(n13443), .A(n13442), .ZN(P2_U2976) );
  INV_X1 U16888 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n13446) );
  AOI21_X1 U16889 ( .B1(n14195), .B2(P2_EAX_REG_7__SCAN_IN), .A(n13444), .ZN(
        n13445) );
  OAI21_X1 U16890 ( .B1(n13456), .B2(n13446), .A(n13445), .ZN(P2_U2974) );
  INV_X1 U16891 ( .A(P2_UWORD_REG_9__SCAN_IN), .ZN(n13449) );
  AOI21_X1 U16892 ( .B1(n14195), .B2(P2_EAX_REG_25__SCAN_IN), .A(n13447), .ZN(
        n13448) );
  OAI21_X1 U16893 ( .B1(n13456), .B2(n13449), .A(n13448), .ZN(P2_U2961) );
  INV_X1 U16894 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n13452) );
  AOI21_X1 U16895 ( .B1(P2_EAX_REG_17__SCAN_IN), .B2(n14195), .A(n13450), .ZN(
        n13451) );
  OAI21_X1 U16896 ( .B1(n13456), .B2(n13452), .A(n13451), .ZN(P2_U2953) );
  INV_X1 U16897 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13455) );
  AOI22_X1 U16898 ( .A1(n19521), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n19519), .ZN(n14355) );
  INV_X1 U16899 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13453) );
  OAI222_X1 U16900 ( .A1(n13456), .A2(n13455), .B1(n13454), .B2(n14355), .C1(
        n13534), .C2(n13453), .ZN(P2_U2982) );
  INV_X1 U16901 ( .A(n13457), .ZN(n13459) );
  INV_X1 U16902 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n13458) );
  AND2_X1 U16903 ( .A1(n20811), .A2(n20942), .ZN(n14410) );
  INV_X1 U16904 ( .A(n14410), .ZN(n14846) );
  OAI211_X1 U16905 ( .C1(n13459), .C2(n13458), .A(n13660), .B(n14846), .ZN(
        P1_U2801) );
  OR2_X1 U16906 ( .A1(n19501), .A2(n13460), .ZN(n13465) );
  OAI21_X1 U16907 ( .B1(n14341), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13474), .ZN(n13615) );
  NOR2_X1 U16908 ( .A1(n16671), .A2(n13615), .ZN(n13464) );
  OAI21_X1 U16909 ( .B1(n13462), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13461), .ZN(n13614) );
  OR2_X1 U16910 ( .A1(n19395), .A2(n19227), .ZN(n13613) );
  OAI21_X1 U16911 ( .B1(n16668), .B2(n13614), .A(n13613), .ZN(n13463) );
  AOI211_X1 U16912 ( .C1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .C2(n13465), .A(
        n13464), .B(n13463), .ZN(n13466) );
  OAI21_X1 U16913 ( .B1(n13467), .B2(n16655), .A(n13466), .ZN(P2_U3014) );
  NAND2_X1 U16914 ( .A1(n13468), .A2(n12630), .ZN(n13470) );
  NAND2_X1 U16915 ( .A1(n14851), .A2(n14160), .ZN(n13469) );
  NAND2_X1 U16916 ( .A1(n13470), .A2(n13469), .ZN(n14859) );
  NOR2_X1 U16917 ( .A1(n14859), .A2(n14081), .ZN(n13472) );
  INV_X1 U16918 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21194) );
  NAND2_X1 U16919 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14410), .ZN(n13471) );
  OAI21_X1 U16920 ( .B1(n13472), .B2(n21194), .A(n13471), .ZN(P1_U2803) );
  OAI21_X1 U16921 ( .B1(n14318), .B2(n13474), .A(n13473), .ZN(n13475) );
  XOR2_X1 U16922 ( .A(n13475), .B(n14308), .Z(n13633) );
  AOI21_X1 U16923 ( .B1(n14308), .B2(n13477), .A(n13476), .ZN(n13625) );
  INV_X1 U16924 ( .A(n13625), .ZN(n13480) );
  AOI22_X1 U16925 ( .A1(n19501), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19500), .ZN(n13479) );
  INV_X1 U16926 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14319) );
  NAND2_X1 U16927 ( .A1(n16667), .A2(n14319), .ZN(n13478) );
  OAI211_X1 U16928 ( .C1(n16668), .C2(n13480), .A(n13479), .B(n13478), .ZN(
        n13481) );
  AOI21_X1 U16929 ( .B1(n10923), .B2(n13633), .A(n13481), .ZN(n13482) );
  OAI21_X1 U16930 ( .B1(n10342), .B2(n16655), .A(n13482), .ZN(P2_U3013) );
  AOI22_X1 U16931 ( .A1(n19521), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19519), .ZN(n19540) );
  INV_X1 U16932 ( .A(n19540), .ZN(n13922) );
  NAND2_X1 U16933 ( .A1(n13500), .A2(n13922), .ZN(n13503) );
  NAND2_X1 U16934 ( .A1(n13517), .A2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13484) );
  OAI211_X1 U16935 ( .C1(n13534), .C2(n13485), .A(n13503), .B(n13484), .ZN(
        P2_U2954) );
  INV_X1 U16936 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13487) );
  AOI22_X1 U16937 ( .A1(n19521), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13498), .ZN(n19523) );
  INV_X1 U16938 ( .A(n19523), .ZN(n13653) );
  NAND2_X1 U16939 ( .A1(n13500), .A2(n13653), .ZN(n13489) );
  NAND2_X1 U16940 ( .A1(n13517), .A2(P2_LWORD_REG_0__SCAN_IN), .ZN(n13486) );
  OAI211_X1 U16941 ( .C1(n13487), .C2(n13534), .A(n13489), .B(n13486), .ZN(
        P2_U2967) );
  NAND2_X1 U16942 ( .A1(n13517), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13488) );
  OAI211_X1 U16943 ( .C1(n13534), .C2(n13490), .A(n13489), .B(n13488), .ZN(
        P2_U2952) );
  INV_X1 U16944 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15621) );
  NAND2_X1 U16945 ( .A1(n13517), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13491) );
  OAI211_X1 U16946 ( .C1(n13534), .C2(n15621), .A(n13492), .B(n13491), .ZN(
        P2_U2965) );
  INV_X1 U16947 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n13728) );
  INV_X1 U16948 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16783) );
  INV_X1 U16949 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17670) );
  MUX2_X1 U16950 ( .A(n16783), .B(n17670), .S(n19519), .Z(n15627) );
  INV_X1 U16951 ( .A(n15627), .ZN(n19459) );
  NAND2_X1 U16952 ( .A1(n13500), .A2(n19459), .ZN(n13516) );
  NAND2_X1 U16953 ( .A1(n13517), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13493) );
  OAI211_X1 U16954 ( .C1(n13728), .C2(n13534), .A(n13516), .B(n13493), .ZN(
        P2_U2964) );
  INV_X1 U16955 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15635) );
  AOI22_X1 U16956 ( .A1(n19521), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n13498), .ZN(n15636) );
  INV_X1 U16957 ( .A(n15636), .ZN(n13494) );
  NAND2_X1 U16958 ( .A1(n13500), .A2(n13494), .ZN(n13513) );
  NAND2_X1 U16959 ( .A1(n13517), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13495) );
  OAI211_X1 U16960 ( .C1(n13534), .C2(n15635), .A(n13513), .B(n13495), .ZN(
        P2_U2963) );
  NAND2_X1 U16961 ( .A1(n13517), .A2(P2_LWORD_REG_4__SCAN_IN), .ZN(n13496) );
  OAI211_X1 U16962 ( .C1(n13534), .C2(n14276), .A(n13497), .B(n13496), .ZN(
        P2_U2971) );
  INV_X1 U16963 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n15644) );
  AOI22_X1 U16964 ( .A1(n19521), .A2(BUF1_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n13498), .ZN(n15645) );
  INV_X1 U16965 ( .A(n15645), .ZN(n13499) );
  NAND2_X1 U16966 ( .A1(n13500), .A2(n13499), .ZN(n13519) );
  NAND2_X1 U16967 ( .A1(n13517), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13501) );
  OAI211_X1 U16968 ( .C1(n13534), .C2(n15644), .A(n13519), .B(n13501), .ZN(
        P2_U2962) );
  NAND2_X1 U16969 ( .A1(n13517), .A2(P2_LWORD_REG_2__SCAN_IN), .ZN(n13502) );
  OAI211_X1 U16970 ( .C1(n13534), .C2(n19493), .A(n13503), .B(n13502), .ZN(
        P2_U2969) );
  NAND2_X1 U16971 ( .A1(n13517), .A2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13504) );
  OAI211_X1 U16972 ( .C1(n13534), .C2(n13506), .A(n13505), .B(n13504), .ZN(
        P2_U2958) );
  NAND2_X1 U16973 ( .A1(n13517), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13507) );
  OAI211_X1 U16974 ( .C1(n13534), .C2(n13509), .A(n13508), .B(n13507), .ZN(
        P2_U2960) );
  NAND2_X1 U16975 ( .A1(n13517), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n13510) );
  OAI211_X1 U16976 ( .C1(n11584), .C2(n13534), .A(n13511), .B(n13510), .ZN(
        P2_U2981) );
  NAND2_X1 U16977 ( .A1(n13517), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13512) );
  OAI211_X1 U16978 ( .C1(n13534), .C2(n13514), .A(n13513), .B(n13512), .ZN(
        P2_U2978) );
  NAND2_X1 U16979 ( .A1(n13517), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13515) );
  OAI211_X1 U16980 ( .C1(n11541), .C2(n13534), .A(n13516), .B(n13515), .ZN(
        P2_U2979) );
  NAND2_X1 U16981 ( .A1(n13517), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13518) );
  OAI211_X1 U16982 ( .C1(n13520), .C2(n13534), .A(n13519), .B(n13518), .ZN(
        P2_U2977) );
  NAND2_X1 U16983 ( .A1(n13522), .A2(n13521), .ZN(n13523) );
  NOR2_X1 U16984 ( .A1(n13524), .A2(n13523), .ZN(n13528) );
  INV_X1 U16985 ( .A(n13536), .ZN(n13526) );
  INV_X1 U16986 ( .A(n14031), .ZN(n13993) );
  NOR2_X1 U16987 ( .A1(n11314), .A2(n13993), .ZN(n13525) );
  NAND2_X1 U16988 ( .A1(n13526), .A2(n13525), .ZN(n13527) );
  NAND2_X1 U16989 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n16270) );
  NOR2_X1 U16990 ( .A1(n20218), .A2(n16270), .ZN(n16272) );
  INV_X1 U16991 ( .A(n16272), .ZN(n16726) );
  OAI22_X1 U16992 ( .A1(n14046), .A2(n19210), .B1(n19213), .B2(n16726), .ZN(
        n13529) );
  AOI21_X1 U16993 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20218), .A(n13529), 
        .ZN(n14314) );
  NOR2_X1 U16994 ( .A1(n11314), .A2(n15586), .ZN(n14029) );
  INV_X1 U16995 ( .A(n20165), .ZN(n13530) );
  NAND4_X1 U16996 ( .A1(n20162), .A2(n14029), .A3(n14028), .A4(n13530), .ZN(
        n13531) );
  OAI21_X1 U16997 ( .B1(n20162), .B2(n13532), .A(n13531), .ZN(P2_U3595) );
  INV_X1 U16998 ( .A(n13533), .ZN(n13535) );
  OAI21_X1 U16999 ( .B1(n13536), .B2(n13535), .A(n13534), .ZN(n13537) );
  INV_X1 U17000 ( .A(n20225), .ZN(n20219) );
  AND2_X1 U17001 ( .A1(n13537), .A2(n20219), .ZN(n19472) );
  NAND2_X1 U17002 ( .A1(n19472), .A2(n20224), .ZN(n13739) );
  INV_X1 U17003 ( .A(n13737), .ZN(n20214) );
  AOI22_X1 U17004 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n19484), .B1(n19497), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13538) );
  OAI21_X1 U17005 ( .B1(n13190), .B2(n13739), .A(n13538), .ZN(P2_U2921) );
  AOI22_X1 U17006 ( .A1(n19497), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13539) );
  OAI21_X1 U17007 ( .B1(n15653), .B2(n13739), .A(n13539), .ZN(P2_U2926) );
  AOI22_X1 U17008 ( .A1(n19497), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13540) );
  OAI21_X1 U17009 ( .B1(n15666), .B2(n13739), .A(n13540), .ZN(P2_U2928) );
  AOI22_X1 U17010 ( .A1(n13737), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13541) );
  OAI21_X1 U17011 ( .B1(n15635), .B2(n13739), .A(n13541), .ZN(P2_U2924) );
  OAI21_X1 U17012 ( .B1(n9717), .B2(n11941), .A(n13658), .ZN(n13544) );
  NAND2_X1 U17013 ( .A1(n13544), .A2(n13543), .ZN(n13574) );
  NAND2_X1 U17014 ( .A1(n13546), .A2(n13545), .ZN(n13547) );
  NAND2_X1 U17015 ( .A1(n13547), .A2(n13675), .ZN(n13548) );
  NAND3_X1 U17016 ( .A1(n13549), .A2(n13574), .A3(n13548), .ZN(n13700) );
  INV_X1 U17017 ( .A(n13550), .ZN(n13554) );
  INV_X1 U17018 ( .A(n13551), .ZN(n13553) );
  NAND4_X1 U17019 ( .A1(n13555), .A2(n13554), .A3(n13553), .A4(n13552), .ZN(
        n13556) );
  NOR2_X1 U17020 ( .A1(n13700), .A2(n13556), .ZN(n13558) );
  AND2_X1 U17021 ( .A1(n13558), .A2(n13557), .ZN(n15495) );
  NAND2_X1 U17022 ( .A1(n14850), .A2(n14088), .ZN(n13863) );
  XNOR2_X1 U17023 ( .A(n13559), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13561) );
  AND2_X1 U17024 ( .A1(n12572), .A2(n13675), .ZN(n16217) );
  XNOR2_X1 U17025 ( .A(n11740), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13560) );
  AOI22_X1 U17026 ( .A1(n13863), .A2(n13561), .B1(n16217), .B2(n13560), .ZN(
        n13563) );
  INV_X1 U17027 ( .A(n13561), .ZN(n13564) );
  NAND3_X1 U17028 ( .A1(n15495), .A2(n13865), .A3(n13564), .ZN(n13562) );
  OAI211_X1 U17029 ( .C1(n13542), .C2(n15495), .A(n13563), .B(n13562), .ZN(
        n13855) );
  OAI22_X1 U17030 ( .A1(n14709), .A2(n20451), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15501) );
  INV_X1 U17031 ( .A(n15501), .ZN(n13565) );
  INV_X1 U17032 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20455) );
  NOR2_X1 U17033 ( .A1(n20942), .A2(n20455), .ZN(n15500) );
  AOI222_X1 U17034 ( .A1(n13855), .A2(n15498), .B1(n13565), .B2(n15500), .C1(
        n13882), .C2(n13564), .ZN(n13582) );
  NAND2_X1 U17035 ( .A1(n16217), .A2(n16265), .ZN(n13567) );
  OR2_X1 U17036 ( .A1(n12630), .A2(n13675), .ZN(n13696) );
  INV_X1 U17037 ( .A(n13696), .ZN(n13566) );
  NAND2_X1 U17038 ( .A1(n13566), .A2(n16265), .ZN(n16240) );
  NAND2_X1 U17039 ( .A1(n13567), .A2(n16240), .ZN(n13584) );
  OR2_X1 U17040 ( .A1(n13584), .A2(n13551), .ZN(n13570) );
  INV_X1 U17041 ( .A(n21027), .ZN(n21018) );
  AOI21_X1 U17042 ( .B1(n14084), .B2(n13674), .A(n21018), .ZN(n13569) );
  INV_X1 U17043 ( .A(n14088), .ZN(n13568) );
  AOI21_X1 U17044 ( .B1(n13570), .B2(n13569), .A(n13568), .ZN(n13571) );
  MUX2_X1 U17045 ( .A(n13571), .B(n14850), .S(n14851), .Z(n13580) );
  INV_X1 U17046 ( .A(n13572), .ZN(n13573) );
  OR2_X1 U17047 ( .A1(n12572), .A2(n13573), .ZN(n13575) );
  NAND2_X1 U17048 ( .A1(n13575), .A2(n13574), .ZN(n13684) );
  INV_X1 U17049 ( .A(n13684), .ZN(n13577) );
  NAND2_X1 U17050 ( .A1(n13576), .A2(n21027), .ZN(n13676) );
  OR2_X1 U17051 ( .A1(n13557), .A2(n13676), .ZN(n14083) );
  OAI211_X1 U17052 ( .C1(n14162), .C2(n13678), .A(n13577), .B(n14083), .ZN(
        n13578) );
  INV_X1 U17053 ( .A(n13578), .ZN(n13579) );
  NAND2_X1 U17054 ( .A1(n13877), .A2(n14860), .ZN(n16455) );
  NAND2_X1 U17055 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16467) );
  NOR2_X1 U17056 ( .A1(n21023), .A2(n16467), .ZN(n13881) );
  NAND2_X1 U17057 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13881), .ZN(n13581) );
  OAI211_X1 U17058 ( .C1(P1_STATE2_REG_0__SCAN_IN), .C2(n20774), .A(n16455), 
        .B(n13581), .ZN(n16460) );
  MUX2_X1 U17059 ( .A(n11740), .B(n13582), .S(n16460), .Z(n13583) );
  INV_X1 U17060 ( .A(n13583), .ZN(P1_U3472) );
  INV_X1 U17061 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13586) );
  NAND2_X1 U17062 ( .A1(n20352), .A2(n11889), .ZN(n13822) );
  NOR2_X1 U17063 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16467), .ZN(n20373) );
  NOR2_X4 U17064 ( .A1(n20352), .A2(n21028), .ZN(n16268) );
  AOI22_X1 U17065 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13585) );
  OAI21_X1 U17066 ( .B1(n13586), .B2(n13822), .A(n13585), .ZN(P1_U2912) );
  INV_X1 U17067 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13588) );
  AOI22_X1 U17068 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13587) );
  OAI21_X1 U17069 ( .B1(n13588), .B2(n13822), .A(n13587), .ZN(P1_U2909) );
  INV_X1 U17070 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13590) );
  AOI22_X1 U17071 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13589) );
  OAI21_X1 U17072 ( .B1(n13590), .B2(n13822), .A(n13589), .ZN(P1_U2913) );
  INV_X1 U17073 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13592) );
  AOI22_X1 U17074 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13591) );
  OAI21_X1 U17075 ( .B1(n13592), .B2(n13822), .A(n13591), .ZN(P1_U2907) );
  INV_X1 U17076 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13594) );
  AOI22_X1 U17077 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13593) );
  OAI21_X1 U17078 ( .B1(n13594), .B2(n13822), .A(n13593), .ZN(P1_U2917) );
  INV_X1 U17079 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13596) );
  AOI22_X1 U17080 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13595) );
  OAI21_X1 U17081 ( .B1(n13596), .B2(n13822), .A(n13595), .ZN(P1_U2908) );
  INV_X1 U17082 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13598) );
  AOI22_X1 U17083 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13597) );
  OAI21_X1 U17084 ( .B1(n13598), .B2(n13822), .A(n13597), .ZN(P1_U2915) );
  AOI22_X1 U17085 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13599) );
  OAI21_X1 U17086 ( .B1(n15092), .B2(n13822), .A(n13599), .ZN(P1_U2916) );
  AOI22_X1 U17087 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13600) );
  OAI21_X1 U17088 ( .B1(n12393), .B2(n13822), .A(n13600), .ZN(P1_U2914) );
  INV_X1 U17089 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n13602) );
  AOI22_X1 U17090 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13601) );
  OAI21_X1 U17091 ( .B1(n13602), .B2(n13822), .A(n13601), .ZN(P1_U2911) );
  INV_X1 U17092 ( .A(n16460), .ZN(n13606) );
  AOI21_X1 U17093 ( .B1(n16217), .B2(n15498), .A(n13606), .ZN(n13608) );
  INV_X1 U17094 ( .A(n15495), .ZN(n13871) );
  NOR2_X1 U17095 ( .A1(n11897), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13603) );
  AOI21_X1 U17096 ( .B1(n12024), .B2(n13871), .A(n13603), .ZN(n16219) );
  INV_X1 U17097 ( .A(n16219), .ZN(n13605) );
  OAI22_X1 U17098 ( .A1(n20942), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16251), .ZN(n13604) );
  AOI21_X1 U17099 ( .B1(n13605), .B2(n15498), .A(n13604), .ZN(n13607) );
  OAI22_X1 U17100 ( .A1(n13608), .A2(n11741), .B1(n13607), .B2(n13606), .ZN(
        P1_U3474) );
  NOR2_X1 U17101 ( .A1(n13610), .A2(n13609), .ZN(n13611) );
  NOR2_X1 U17102 ( .A1(n13612), .A2(n13611), .ZN(n14340) );
  INV_X1 U17103 ( .A(n14340), .ZN(n13656) );
  OAI21_X1 U17104 ( .B1(n16072), .B2(n13656), .A(n13613), .ZN(n13617) );
  OAI22_X1 U17105 ( .A1(n16704), .A2(n13615), .B1(n16717), .B2(n13614), .ZN(
        n13616) );
  AOI211_X1 U17106 ( .C1(n14346), .C2(n16699), .A(n13617), .B(n13616), .ZN(
        n13619) );
  MUX2_X1 U17107 ( .A(n15968), .B(n14765), .S(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Z(n13618) );
  NAND2_X1 U17108 ( .A1(n13619), .A2(n13618), .ZN(P2_U3046) );
  INV_X1 U17109 ( .A(n13835), .ZN(n14791) );
  NAND2_X1 U17110 ( .A1(n20195), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19206) );
  NOR2_X1 U17111 ( .A1(n13746), .A2(n19206), .ZN(n13620) );
  OAI21_X1 U17112 ( .B1(n9730), .B2(n19532), .A(n13620), .ZN(n13621) );
  NAND2_X1 U17113 ( .A1(n19779), .A2(n14786), .ZN(n13624) );
  NAND2_X1 U17114 ( .A1(n14346), .A2(n15616), .ZN(n13623) );
  OAI211_X1 U17115 ( .C1(n14791), .C2(n14344), .A(n13624), .B(n13623), .ZN(
        P2_U2887) );
  NAND2_X1 U17116 ( .A1(n16700), .A2(n13625), .ZN(n13626) );
  OAI21_X1 U17117 ( .B1(n20102), .B2(n19341), .A(n13626), .ZN(n13632) );
  OAI211_X1 U17118 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n14598), .B(n14768), .ZN(n13630) );
  XNOR2_X1 U17119 ( .A(n13627), .B(n13628), .ZN(n14325) );
  INV_X1 U17120 ( .A(n14325), .ZN(n20186) );
  NAND2_X1 U17121 ( .A1(n16710), .A2(n20186), .ZN(n13629) );
  OAI211_X1 U17122 ( .C1(n14765), .C2(n14308), .A(n13630), .B(n13629), .ZN(
        n13631) );
  AOI211_X1 U17123 ( .C1(n16721), .C2(n13633), .A(n13632), .B(n13631), .ZN(
        n13634) );
  OAI21_X1 U17124 ( .B1(n10342), .B2(n16716), .A(n13634), .ZN(P2_U3045) );
  MUX2_X1 U17125 ( .A(n14320), .B(n10342), .S(n15616), .Z(n13639) );
  OAI21_X1 U17126 ( .B1(n19513), .B2(n15618), .A(n13639), .ZN(P2_U2886) );
  MUX2_X1 U17127 ( .A(n10287), .B(n10352), .S(n15616), .Z(n13642) );
  OAI21_X1 U17128 ( .B1(n20178), .B2(n15618), .A(n13642), .ZN(P2_U2885) );
  XNOR2_X1 U17129 ( .A(n20190), .B(n14325), .ZN(n13644) );
  NAND2_X1 U17130 ( .A1(n19779), .A2(n14340), .ZN(n13643) );
  NAND2_X1 U17131 ( .A1(n13644), .A2(n13643), .ZN(n13917) );
  OAI21_X1 U17132 ( .B1(n13644), .B2(n13643), .A(n13917), .ZN(n13645) );
  NAND2_X1 U17133 ( .A1(n13645), .A2(n13177), .ZN(n13648) );
  INV_X1 U17134 ( .A(n19533), .ZN(n16571) );
  AOI22_X1 U17135 ( .A1(n19464), .A2(n16571), .B1(P2_EAX_REG_1__SCAN_IN), .B2(
        n19462), .ZN(n13647) );
  OAI211_X1 U17136 ( .C1(n14325), .C2(n15675), .A(n13648), .B(n13647), .ZN(
        P2_U2918) );
  OR2_X1 U17137 ( .A1(n13650), .A2(n13649), .ZN(n13651) );
  NAND2_X1 U17138 ( .A1(n13825), .A2(n13651), .ZN(n20343) );
  XNOR2_X1 U17139 ( .A(n20350), .B(n14084), .ZN(n13707) );
  AOI22_X1 U17140 ( .A1(n15038), .A2(n13707), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n15037), .ZN(n13652) );
  OAI21_X1 U17141 ( .B1(n20343), .B2(n15040), .A(n13652), .ZN(P1_U2871) );
  AOI21_X1 U17142 ( .B1(n20197), .B2(n13177), .A(n19449), .ZN(n13657) );
  AOI22_X1 U17143 ( .A1(n19464), .A2(n13653), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19462), .ZN(n13655) );
  NAND3_X1 U17144 ( .A1(n19779), .A2(n13177), .A3(n13656), .ZN(n13654) );
  OAI211_X1 U17145 ( .C1(n13657), .C2(n13656), .A(n13655), .B(n13654), .ZN(
        P2_U2919) );
  AND2_X1 U17146 ( .A1(n13658), .A2(n21018), .ZN(n13659) );
  OR2_X1 U17147 ( .A1(n20383), .A2(n9669), .ZN(n13761) );
  INV_X1 U17148 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13665) );
  INV_X1 U17149 ( .A(n20398), .ZN(n13664) );
  INV_X1 U17150 ( .A(DATAI_15_), .ZN(n13661) );
  NOR2_X1 U17151 ( .A1(n14699), .A2(n13661), .ZN(n13662) );
  AOI21_X1 U17152 ( .B1(n14699), .B2(BUF1_REG_15__SCAN_IN), .A(n13662), .ZN(
        n14585) );
  INV_X1 U17153 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13663) );
  OAI222_X1 U17154 ( .A1(n13761), .A2(n13665), .B1(n13664), .B2(n14585), .C1(
        n13663), .C2(n13795), .ZN(P1_U2967) );
  XNOR2_X1 U17155 ( .A(n13667), .B(n13666), .ZN(n19406) );
  OAI222_X1 U17156 ( .A1(n14356), .A2(n19567), .B1(n19406), .B2(n19471), .C1(
        n19483), .C2(n15689), .ZN(P2_U2912) );
  INV_X1 U17157 ( .A(n13668), .ZN(n13669) );
  XNOR2_X1 U17158 ( .A(n13670), .B(n13669), .ZN(n14599) );
  INV_X1 U17159 ( .A(n14599), .ZN(n19424) );
  OAI222_X1 U17160 ( .A1(n14356), .A2(n19559), .B1(n19424), .B2(n19471), .C1(
        n19486), .C2(n15689), .ZN(P2_U2913) );
  OR2_X1 U17161 ( .A1(n13671), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13846) );
  NAND2_X1 U17162 ( .A1(n13673), .A2(n9669), .ZN(n13681) );
  NAND2_X1 U17163 ( .A1(n13675), .A2(n13674), .ZN(n13679) );
  INV_X1 U17164 ( .A(n13676), .ZN(n13677) );
  NAND3_X1 U17165 ( .A1(n13679), .A2(n13678), .A3(n13677), .ZN(n13680) );
  OAI21_X1 U17166 ( .B1(n13682), .B2(n13681), .A(n13680), .ZN(n13683) );
  OAI21_X1 U17167 ( .B1(n13684), .B2(n13683), .A(n14860), .ZN(n13691) );
  NAND2_X1 U17168 ( .A1(n13551), .A2(n21027), .ZN(n14085) );
  INV_X1 U17169 ( .A(n13685), .ZN(n13687) );
  OAI211_X1 U17170 ( .C1(n14085), .C2(n13687), .A(n11889), .B(n13686), .ZN(
        n13689) );
  NAND3_X1 U17171 ( .A1(n13689), .A2(n13688), .A3(n12770), .ZN(n13690) );
  INV_X1 U17172 ( .A(n13692), .ZN(n13694) );
  AND2_X1 U17173 ( .A1(n14088), .A2(n13693), .ZN(n14849) );
  OAI211_X1 U17174 ( .C1(n14106), .C2(n10116), .A(n13694), .B(n14849), .ZN(
        n13695) );
  NAND3_X1 U17175 ( .A1(n13846), .A2(n13672), .A3(n20452), .ZN(n13709) );
  OAI21_X1 U17176 ( .B1(n10116), .B2(n9698), .A(n13696), .ZN(n13697) );
  INV_X1 U17177 ( .A(n14850), .ZN(n13698) );
  OR2_X1 U17178 ( .A1(n13700), .A2(n13699), .ZN(n13701) );
  OR2_X1 U17179 ( .A1(n13703), .A2(n20473), .ZN(n15411) );
  OAI21_X1 U17180 ( .B1(n13704), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n15411), .ZN(n20449) );
  AOI21_X1 U17181 ( .B1(n20467), .B2(n20455), .A(n20449), .ZN(n20476) );
  INV_X1 U17182 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n13702) );
  OR2_X1 U17183 ( .A1(n20432), .A2(n13702), .ZN(n13843) );
  OAI21_X1 U17184 ( .B1(n20476), .B2(n20451), .A(n13843), .ZN(n13706) );
  NAND2_X1 U17185 ( .A1(n16404), .A2(n20428), .ZN(n16425) );
  INV_X1 U17186 ( .A(n16425), .ZN(n14718) );
  NOR3_X1 U17187 ( .A1(n14718), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n14725), .ZN(n13705) );
  AOI211_X1 U17188 ( .C1(n20440), .C2(n13707), .A(n13706), .B(n13705), .ZN(
        n13708) );
  NAND2_X1 U17189 ( .A1(n13709), .A2(n13708), .ZN(P1_U3030) );
  OAI21_X1 U17190 ( .B1(n13711), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13710), .ZN(n20471) );
  INV_X1 U17191 ( .A(n13712), .ZN(n13715) );
  OAI21_X1 U17192 ( .B1(n13715), .B2(n13714), .A(n13713), .ZN(n14364) );
  INV_X1 U17193 ( .A(n14364), .ZN(n13716) );
  NAND2_X1 U17194 ( .A1(n13716), .A2(n16364), .ZN(n13720) );
  OR2_X1 U17195 ( .A1(n20416), .A2(n13717), .ZN(n13718) );
  AOI22_X1 U17196 ( .A1(n13718), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n20473), .B2(P1_REIP_REG_0__SCAN_IN), .ZN(n13719) );
  OAI211_X1 U17197 ( .C1(n20238), .C2(n20471), .A(n13720), .B(n13719), .ZN(
        P1_U2999) );
  AOI21_X1 U17198 ( .B1(n13723), .B2(n13722), .A(n13721), .ZN(n16709) );
  INV_X1 U17199 ( .A(n16709), .ZN(n13724) );
  OAI222_X1 U17200 ( .A1(n14356), .A2(n15661), .B1(n13724), .B2(n19471), .C1(
        n13423), .C2(n15689), .ZN(P2_U2911) );
  AOI22_X1 U17201 ( .A1(n19497), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13725) );
  OAI21_X1 U17202 ( .B1(n15644), .B2(n13739), .A(n13725), .ZN(P2_U2925) );
  AOI22_X1 U17203 ( .A1(n19497), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13726) );
  OAI21_X1 U17204 ( .B1(n13509), .B2(n13739), .A(n13726), .ZN(P2_U2927) );
  AOI22_X1 U17205 ( .A1(n13737), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13727) );
  OAI21_X1 U17206 ( .B1(n13728), .B2(n13739), .A(n13727), .ZN(P2_U2923) );
  AOI22_X1 U17207 ( .A1(n13737), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13729) );
  OAI21_X1 U17208 ( .B1(n13490), .B2(n13739), .A(n13729), .ZN(P2_U2935) );
  AOI22_X1 U17209 ( .A1(n13737), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13730) );
  OAI21_X1 U17210 ( .B1(n13731), .B2(n13739), .A(n13730), .ZN(P2_U2934) );
  AOI22_X1 U17211 ( .A1(n13737), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13732) );
  OAI21_X1 U17212 ( .B1(n13485), .B2(n13739), .A(n13732), .ZN(P2_U2933) );
  AOI22_X1 U17213 ( .A1(n13737), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13733) );
  OAI21_X1 U17214 ( .B1(n14638), .B2(n13739), .A(n13733), .ZN(P2_U2932) );
  AOI22_X1 U17215 ( .A1(n13737), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13734) );
  OAI21_X1 U17216 ( .B1(n13418), .B2(n13739), .A(n13734), .ZN(P2_U2931) );
  AOI22_X1 U17217 ( .A1(n13737), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13735) );
  OAI21_X1 U17218 ( .B1(n15680), .B2(n13739), .A(n13735), .ZN(P2_U2930) );
  AOI22_X1 U17219 ( .A1(n13737), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13736) );
  OAI21_X1 U17220 ( .B1(n13506), .B2(n13739), .A(n13736), .ZN(P2_U2929) );
  AOI22_X1 U17221 ( .A1(n13737), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13738) );
  OAI21_X1 U17222 ( .B1(n15621), .B2(n13739), .A(n13738), .ZN(P2_U2922) );
  NOR2_X1 U17223 ( .A1(n15616), .A2(n10301), .ZN(n13742) );
  AOI21_X1 U17224 ( .B1(n9734), .B2(n15616), .A(n13742), .ZN(n13743) );
  OAI21_X1 U17225 ( .B1(n20167), .B2(n15618), .A(n13743), .ZN(P2_U2884) );
  NAND2_X1 U17226 ( .A1(n13744), .A2(n13740), .ZN(n13749) );
  INV_X1 U17227 ( .A(n13745), .ZN(n13747) );
  AOI22_X1 U17228 ( .A1(n13741), .A2(n13747), .B1(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13746), .ZN(n13748) );
  NAND2_X1 U17229 ( .A1(n13749), .A2(n13748), .ZN(n13752) );
  AND2_X1 U17230 ( .A1(n13750), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13751) );
  NAND2_X1 U17231 ( .A1(n13752), .A2(n13751), .ZN(n14785) );
  OR2_X1 U17232 ( .A1(n13752), .A2(n13751), .ZN(n13753) );
  NAND2_X1 U17233 ( .A1(n14785), .A2(n13753), .ZN(n19466) );
  OR2_X1 U17234 ( .A1(n13755), .A2(n13754), .ZN(n13756) );
  AND2_X1 U17235 ( .A1(n14455), .A2(n13756), .ZN(n19503) );
  NOR2_X1 U17236 ( .A1(n14791), .A2(n14222), .ZN(n13757) );
  AOI21_X1 U17237 ( .B1(n19503), .B2(n15616), .A(n13757), .ZN(n13758) );
  OAI21_X1 U17238 ( .B1(n19466), .B2(n15618), .A(n13758), .ZN(P2_U2883) );
  OAI21_X1 U17239 ( .B1(n13760), .B2(n13721), .A(n13759), .ZN(n19391) );
  INV_X1 U17240 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19480) );
  OAI222_X1 U17241 ( .A1(n14356), .A2(n15654), .B1(n19391), .B2(n19471), .C1(
        n19480), .C2(n15689), .ZN(P2_U2910) );
  AOI22_X1 U17242 ( .A1(n20413), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20412), .ZN(n13765) );
  INV_X1 U17243 ( .A(n14699), .ZN(n14104) );
  NAND2_X1 U17244 ( .A1(n14104), .A2(DATAI_5_), .ZN(n13763) );
  NAND2_X1 U17245 ( .A1(n14699), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13762) );
  AND2_X1 U17246 ( .A1(n13763), .A2(n13762), .ZN(n15088) );
  INV_X1 U17247 ( .A(n15088), .ZN(n13764) );
  NAND2_X1 U17248 ( .A1(n20398), .A2(n13764), .ZN(n13800) );
  NAND2_X1 U17249 ( .A1(n13765), .A2(n13800), .ZN(P1_U2957) );
  AOI22_X1 U17250 ( .A1(n20413), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20412), .ZN(n13769) );
  NAND2_X1 U17251 ( .A1(n14104), .A2(DATAI_1_), .ZN(n13767) );
  NAND2_X1 U17252 ( .A1(n14699), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13766) );
  AND2_X1 U17253 ( .A1(n13767), .A2(n13766), .ZN(n15108) );
  INV_X1 U17254 ( .A(n15108), .ZN(n13768) );
  NAND2_X1 U17255 ( .A1(n20398), .A2(n13768), .ZN(n13806) );
  NAND2_X1 U17256 ( .A1(n13769), .A2(n13806), .ZN(P1_U2953) );
  AOI22_X1 U17257 ( .A1(n20413), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20412), .ZN(n13773) );
  NAND2_X1 U17258 ( .A1(n14104), .A2(DATAI_2_), .ZN(n13771) );
  NAND2_X1 U17259 ( .A1(n14699), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13770) );
  AND2_X1 U17260 ( .A1(n13771), .A2(n13770), .ZN(n15103) );
  INV_X1 U17261 ( .A(n15103), .ZN(n13772) );
  NAND2_X1 U17262 ( .A1(n20398), .A2(n13772), .ZN(n13798) );
  NAND2_X1 U17263 ( .A1(n13773), .A2(n13798), .ZN(P1_U2954) );
  AOI22_X1 U17264 ( .A1(n20413), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20412), .ZN(n13777) );
  NAND2_X1 U17265 ( .A1(n14104), .A2(DATAI_3_), .ZN(n13775) );
  NAND2_X1 U17266 ( .A1(n14699), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13774) );
  AND2_X1 U17267 ( .A1(n13775), .A2(n13774), .ZN(n15098) );
  INV_X1 U17268 ( .A(n15098), .ZN(n13776) );
  NAND2_X1 U17269 ( .A1(n20398), .A2(n13776), .ZN(n13802) );
  NAND2_X1 U17270 ( .A1(n13777), .A2(n13802), .ZN(P1_U2955) );
  AOI22_X1 U17271 ( .A1(n20413), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20412), .ZN(n13780) );
  INV_X1 U17272 ( .A(DATAI_6_), .ZN(n13779) );
  NAND2_X1 U17273 ( .A1(n14699), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13778) );
  OAI21_X1 U17274 ( .B1(n14699), .B2(n13779), .A(n13778), .ZN(n15081) );
  NAND2_X1 U17275 ( .A1(n20398), .A2(n15081), .ZN(n13789) );
  NAND2_X1 U17276 ( .A1(n13780), .A2(n13789), .ZN(P1_U2958) );
  AOI22_X1 U17277 ( .A1(n20413), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20412), .ZN(n13784) );
  NAND2_X1 U17278 ( .A1(n14104), .A2(DATAI_4_), .ZN(n13782) );
  NAND2_X1 U17279 ( .A1(n14699), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13781) );
  AND2_X1 U17280 ( .A1(n13782), .A2(n13781), .ZN(n15093) );
  INV_X1 U17281 ( .A(n15093), .ZN(n13783) );
  NAND2_X1 U17282 ( .A1(n20398), .A2(n13783), .ZN(n13796) );
  NAND2_X1 U17283 ( .A1(n13784), .A2(n13796), .ZN(P1_U2956) );
  AOI22_X1 U17284 ( .A1(n20413), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20412), .ZN(n13788) );
  NAND2_X1 U17285 ( .A1(n14104), .A2(DATAI_0_), .ZN(n13786) );
  NAND2_X1 U17286 ( .A1(n14699), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13785) );
  AND2_X1 U17287 ( .A1(n13786), .A2(n13785), .ZN(n15117) );
  INV_X1 U17288 ( .A(n15117), .ZN(n13787) );
  NAND2_X1 U17289 ( .A1(n20398), .A2(n13787), .ZN(n13804) );
  NAND2_X1 U17290 ( .A1(n13788), .A2(n13804), .ZN(P1_U2952) );
  AOI22_X1 U17291 ( .A1(n20413), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20412), .ZN(n13790) );
  NAND2_X1 U17292 ( .A1(n13790), .A2(n13789), .ZN(P1_U2943) );
  AOI22_X1 U17293 ( .A1(n20413), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20412), .ZN(n13794) );
  INV_X1 U17294 ( .A(DATAI_7_), .ZN(n13792) );
  INV_X1 U17295 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n13791) );
  MUX2_X1 U17296 ( .A(n13792), .B(n13791), .S(n14699), .Z(n15076) );
  INV_X1 U17297 ( .A(n15076), .ZN(n13793) );
  NAND2_X1 U17298 ( .A1(n20398), .A2(n13793), .ZN(n13808) );
  NAND2_X1 U17299 ( .A1(n13794), .A2(n13808), .ZN(P1_U2944) );
  INV_X1 U17300 ( .A(n13795), .ZN(n20412) );
  AOI22_X1 U17301 ( .A1(n20413), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20412), .ZN(n13797) );
  NAND2_X1 U17302 ( .A1(n13797), .A2(n13796), .ZN(P1_U2941) );
  AOI22_X1 U17303 ( .A1(n20413), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20412), .ZN(n13799) );
  NAND2_X1 U17304 ( .A1(n13799), .A2(n13798), .ZN(P1_U2939) );
  AOI22_X1 U17305 ( .A1(n20413), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20412), .ZN(n13801) );
  NAND2_X1 U17306 ( .A1(n13801), .A2(n13800), .ZN(P1_U2942) );
  AOI22_X1 U17307 ( .A1(n20413), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20412), .ZN(n13803) );
  NAND2_X1 U17308 ( .A1(n13803), .A2(n13802), .ZN(P1_U2940) );
  AOI22_X1 U17309 ( .A1(n20413), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20412), .ZN(n13805) );
  NAND2_X1 U17310 ( .A1(n13805), .A2(n13804), .ZN(P1_U2937) );
  AOI22_X1 U17311 ( .A1(n20413), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20412), .ZN(n13807) );
  NAND2_X1 U17312 ( .A1(n13807), .A2(n13806), .ZN(P1_U2938) );
  AOI22_X1 U17313 ( .A1(n20413), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20412), .ZN(n13809) );
  NAND2_X1 U17314 ( .A1(n13809), .A2(n13808), .ZN(P1_U2959) );
  INV_X1 U17315 ( .A(n13810), .ZN(n13813) );
  NAND2_X1 U17316 ( .A1(n13811), .A2(n20455), .ZN(n13812) );
  NAND2_X1 U17317 ( .A1(n13813), .A2(n13812), .ZN(n20468) );
  OAI222_X1 U17318 ( .A1(n20468), .A2(n15048), .B1(n13814), .B2(n15047), .C1(
        n14364), .C2(n15040), .ZN(P1_U2872) );
  INV_X1 U17319 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13816) );
  AOI22_X1 U17320 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20373), .B1(n16268), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13815) );
  OAI21_X1 U17321 ( .B1(n13816), .B2(n13822), .A(n13815), .ZN(P1_U2920) );
  AOI22_X1 U17322 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20373), .B1(n16268), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13817) );
  OAI21_X1 U17323 ( .B1(n15107), .B2(n13822), .A(n13817), .ZN(P1_U2919) );
  INV_X1 U17324 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n15102) );
  AOI22_X1 U17325 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20373), .B1(n16268), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13818) );
  OAI21_X1 U17326 ( .B1(n15102), .B2(n13822), .A(n13818), .ZN(P1_U2918) );
  INV_X1 U17327 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n13820) );
  AOI22_X1 U17328 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13819) );
  OAI21_X1 U17329 ( .B1(n13820), .B2(n13822), .A(n13819), .ZN(P1_U2910) );
  INV_X1 U17330 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n13823) );
  AOI22_X1 U17331 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n21028), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n16268), .ZN(n13821) );
  OAI21_X1 U17332 ( .B1(n13823), .B2(n13822), .A(n13821), .ZN(P1_U2906) );
  OAI21_X1 U17333 ( .B1(n12031), .B2(n12030), .A(n13826), .ZN(n14175) );
  OAI21_X1 U17334 ( .B1(n13828), .B2(n13827), .A(n13904), .ZN(n20460) );
  INV_X1 U17335 ( .A(n20460), .ZN(n14170) );
  AOI22_X1 U17336 ( .A1(n15038), .A2(n14170), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n15037), .ZN(n13829) );
  OAI21_X1 U17337 ( .B1(n14175), .B2(n15040), .A(n13829), .ZN(P1_U2870) );
  NAND2_X1 U17338 ( .A1(n13831), .A2(n13830), .ZN(n13834) );
  INV_X1 U17339 ( .A(n13832), .ZN(n13833) );
  NAND2_X1 U17340 ( .A1(n13834), .A2(n13833), .ZN(n19405) );
  NOR2_X1 U17341 ( .A1(n13836), .A2(n13837), .ZN(n13840) );
  INV_X1 U17342 ( .A(n13838), .ZN(n13839) );
  OAI211_X1 U17343 ( .C1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .C2(n13840), .A(
        n13839), .B(n14786), .ZN(n13842) );
  NAND2_X1 U17344 ( .A1(n13835), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n13841) );
  OAI211_X1 U17345 ( .C1(n19405), .C2(n13835), .A(n13842), .B(n13841), .ZN(
        P2_U2880) );
  INV_X1 U17346 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20337) );
  OAI21_X1 U17347 ( .B1(n15254), .B2(n20337), .A(n13843), .ZN(n13845) );
  NOR2_X1 U17348 ( .A1(n20343), .A2(n15258), .ZN(n13844) );
  AOI211_X1 U17349 ( .C1(n16355), .C2(n20337), .A(n13845), .B(n13844), .ZN(
        n13848) );
  NAND3_X1 U17350 ( .A1(n13846), .A2(n13672), .A3(n20422), .ZN(n13847) );
  NAND2_X1 U17351 ( .A1(n13848), .A2(n13847), .ZN(P1_U2998) );
  NAND2_X1 U17352 ( .A1(n13838), .A2(n13849), .ZN(n13910) );
  OAI211_X1 U17353 ( .C1(n13838), .C2(n13849), .A(n13910), .B(n14786), .ZN(
        n13854) );
  NOR2_X1 U17354 ( .A1(n13851), .A2(n13832), .ZN(n13852) );
  OR2_X1 U17355 ( .A1(n13850), .A2(n13852), .ZN(n16715) );
  INV_X1 U17356 ( .A(n16715), .ZN(n14211) );
  NAND2_X1 U17357 ( .A1(n14791), .A2(n14211), .ZN(n13853) );
  OAI211_X1 U17358 ( .C1(n14791), .C2(n10680), .A(n13854), .B(n13853), .ZN(
        P2_U2879) );
  MUX2_X1 U17359 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13855), .S(
        n13877), .Z(n16226) );
  NOR2_X1 U17360 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20942), .ZN(n13878) );
  AOI22_X1 U17361 ( .A1(n16226), .A2(n20942), .B1(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n13878), .ZN(n13874) );
  INV_X1 U17362 ( .A(n16217), .ZN(n13869) );
  XNOR2_X1 U17363 ( .A(n13857), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13868) );
  INV_X1 U17364 ( .A(n13858), .ZN(n13862) );
  INV_X1 U17365 ( .A(n13859), .ZN(n13860) );
  MUX2_X1 U17366 ( .A(n13860), .B(n10066), .S(n13559), .Z(n13861) );
  NAND3_X1 U17367 ( .A1(n13863), .A2(n13862), .A3(n13861), .ZN(n13867) );
  AOI21_X1 U17368 ( .B1(n13559), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13864) );
  NOR2_X1 U17369 ( .A1(n12432), .A2(n13864), .ZN(n15504) );
  NAND3_X1 U17370 ( .A1(n15495), .A2(n13865), .A3(n15504), .ZN(n13866) );
  OAI211_X1 U17371 ( .C1(n13869), .C2(n13868), .A(n13867), .B(n13866), .ZN(
        n13870) );
  AOI21_X1 U17372 ( .B1(n13856), .B2(n13871), .A(n13870), .ZN(n15506) );
  INV_X1 U17373 ( .A(n15506), .ZN(n13872) );
  MUX2_X1 U17374 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13872), .S(
        n13877), .Z(n16229) );
  AOI22_X1 U17375 ( .A1(n13878), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n20942), .B2(n16229), .ZN(n13873) );
  OR2_X1 U17376 ( .A1(n13874), .A2(n13873), .ZN(n16231) );
  INV_X1 U17377 ( .A(n14098), .ZN(n14233) );
  XNOR2_X1 U17378 ( .A(n13876), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n20308) );
  OAI21_X1 U17379 ( .B1(n20308), .B2(n13557), .A(n13877), .ZN(n13880) );
  INV_X1 U17380 ( .A(n13877), .ZN(n16220) );
  AOI21_X1 U17381 ( .B1(n16220), .B2(n16459), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n13879) );
  AOI22_X1 U17382 ( .A1(n13880), .A2(n13879), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13878), .ZN(n16238) );
  OAI21_X1 U17383 ( .B1(n16231), .B2(n13875), .A(n16238), .ZN(n13884) );
  OAI21_X1 U17384 ( .B1(n13884), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13881), .ZN(
        n13883) );
  NAND2_X1 U17385 ( .A1(n13883), .A2(n14500), .ZN(n20478) );
  NOR2_X1 U17386 ( .A1(n13884), .A2(n16467), .ZN(n16246) );
  INV_X1 U17387 ( .A(n12024), .ZN(n13885) );
  AND2_X1 U17388 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20774), .ZN(n15493) );
  OAI22_X1 U17389 ( .A1(n13236), .A2(n20880), .B1(n13885), .B2(n15493), .ZN(
        n13886) );
  OAI21_X1 U17390 ( .B1(n16246), .B2(n13886), .A(n20478), .ZN(n13887) );
  OAI21_X1 U17391 ( .B1(n20478), .B2(n20733), .A(n13887), .ZN(P1_U3478) );
  NAND2_X1 U17392 ( .A1(n13888), .A2(n13759), .ZN(n13891) );
  INV_X1 U17393 ( .A(n13889), .ZN(n13890) );
  NAND2_X1 U17394 ( .A1(n13891), .A2(n13890), .ZN(n16691) );
  OAI222_X1 U17395 ( .A1(n14356), .A2(n15645), .B1(n16691), .B2(n19471), .C1(
        n13520), .C2(n15689), .ZN(P2_U2909) );
  INV_X1 U17396 ( .A(n14175), .ZN(n13895) );
  NOR2_X1 U17397 ( .A1(n20427), .A2(n14164), .ZN(n13894) );
  INV_X1 U17398 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14167) );
  INV_X1 U17399 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13892) );
  OAI22_X1 U17400 ( .A1(n15254), .A2(n14167), .B1(n20432), .B2(n13892), .ZN(
        n13893) );
  AOI211_X1 U17401 ( .C1(n13895), .C2(n16364), .A(n13894), .B(n13893), .ZN(
        n13900) );
  OR2_X1 U17402 ( .A1(n13897), .A2(n13896), .ZN(n20453) );
  NAND3_X1 U17403 ( .A1(n20453), .A2(n13898), .A3(n20422), .ZN(n13899) );
  NAND2_X1 U17404 ( .A1(n13900), .A2(n13899), .ZN(P1_U2997) );
  XNOR2_X1 U17405 ( .A(n13902), .B(n13901), .ZN(n20327) );
  AOI21_X1 U17406 ( .B1(n13904), .B2(n13903), .A(n14063), .ZN(n20441) );
  AOI22_X1 U17407 ( .A1(n20441), .A2(n15038), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n15037), .ZN(n13905) );
  OAI21_X1 U17408 ( .B1(n20327), .B2(n15040), .A(n13905), .ZN(P1_U2869) );
  NOR2_X1 U17409 ( .A1(n13850), .A2(n13907), .ZN(n13908) );
  OR2_X1 U17410 ( .A1(n13906), .A2(n13908), .ZN(n16055) );
  INV_X1 U17411 ( .A(n13910), .ZN(n13938) );
  INV_X1 U17412 ( .A(n13909), .ZN(n13911) );
  OR2_X1 U17413 ( .A1(n13910), .A2(n13909), .ZN(n13928) );
  OAI211_X1 U17414 ( .C1(n13938), .C2(n13911), .A(n14786), .B(n13928), .ZN(
        n13913) );
  NAND2_X1 U17415 ( .A1(n13835), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n13912) );
  OAI211_X1 U17416 ( .C1(n16055), .C2(n13835), .A(n13913), .B(n13912), .ZN(
        P2_U2878) );
  NAND2_X1 U17417 ( .A1(n13915), .A2(n13914), .ZN(n13916) );
  AND2_X1 U17418 ( .A1(n13916), .A2(n9895), .ZN(n14753) );
  XOR2_X1 U17419 ( .A(n14753), .B(n20178), .Z(n13920) );
  NAND2_X1 U17420 ( .A1(n19513), .A2(n14325), .ZN(n13918) );
  NAND2_X1 U17421 ( .A1(n13918), .A2(n13917), .ZN(n13919) );
  NAND2_X1 U17422 ( .A1(n13920), .A2(n13919), .ZN(n13971) );
  OAI21_X1 U17423 ( .B1(n13920), .B2(n13919), .A(n13971), .ZN(n13921) );
  NAND2_X1 U17424 ( .A1(n13921), .A2(n13177), .ZN(n13924) );
  AOI22_X1 U17425 ( .A1(n19464), .A2(n13922), .B1(n19462), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13923) );
  OAI211_X1 U17426 ( .C1(n14753), .C2(n15675), .A(n13924), .B(n13923), .ZN(
        P2_U2917) );
  OAI21_X1 U17427 ( .B1(n13926), .B2(n13889), .A(n13925), .ZN(n19378) );
  OAI222_X1 U17428 ( .A1(n14356), .A2(n15636), .B1(n19378), .B2(n19471), .C1(
        n13514), .C2(n15689), .ZN(P2_U2908) );
  INV_X1 U17429 ( .A(n13928), .ZN(n13930) );
  OR2_X1 U17430 ( .A1(n13928), .A2(n13927), .ZN(n13936) );
  OAI211_X1 U17431 ( .C1(n13930), .C2(n13929), .A(n14786), .B(n13936), .ZN(
        n13935) );
  OR2_X1 U17432 ( .A1(n13906), .A2(n13931), .ZN(n13933) );
  AND2_X1 U17433 ( .A1(n13933), .A2(n13932), .ZN(n16698) );
  NAND2_X1 U17434 ( .A1(n16698), .A2(n15616), .ZN(n13934) );
  OAI211_X1 U17435 ( .C1(n14791), .C2(n10688), .A(n13935), .B(n13934), .ZN(
        P2_U2877) );
  INV_X1 U17436 ( .A(n13936), .ZN(n13941) );
  AND2_X1 U17437 ( .A1(n13938), .A2(n13937), .ZN(n13987) );
  INV_X1 U17438 ( .A(n13987), .ZN(n13939) );
  OAI211_X1 U17439 ( .C1(n13941), .C2(n13940), .A(n13939), .B(n14786), .ZN(
        n13947) );
  NAND2_X1 U17440 ( .A1(n13942), .A2(n13932), .ZN(n13945) );
  INV_X1 U17441 ( .A(n13943), .ZN(n13944) );
  AND2_X1 U17442 ( .A1(n13945), .A2(n13944), .ZN(n19374) );
  NAND2_X1 U17443 ( .A1(n14791), .A2(n19374), .ZN(n13946) );
  OAI211_X1 U17444 ( .C1(n14791), .C2(n13948), .A(n13947), .B(n13946), .ZN(
        P2_U2876) );
  INV_X1 U17445 ( .A(n13954), .ZN(n13950) );
  INV_X1 U17446 ( .A(n20885), .ZN(n13952) );
  INV_X1 U17447 ( .A(n15489), .ZN(n13951) );
  AOI21_X1 U17448 ( .B1(n13952), .B2(n13951), .A(n20705), .ZN(n13956) );
  NOR2_X1 U17449 ( .A1(n20880), .A2(n21170), .ZN(n13953) );
  INV_X1 U17450 ( .A(n13953), .ZN(n13955) );
  NAND2_X1 U17451 ( .A1(n15489), .A2(n13953), .ZN(n20884) );
  OAI22_X1 U17452 ( .A1(n13956), .A2(n13955), .B1(n20884), .B2(n20649), .ZN(
        n14230) );
  NAND2_X1 U17453 ( .A1(n20811), .A2(n21170), .ZN(n20766) );
  INV_X1 U17454 ( .A(n13856), .ZN(n13957) );
  OAI22_X1 U17455 ( .A1(n13254), .A2(n20766), .B1(n13957), .B2(n15493), .ZN(
        n13958) );
  OAI21_X1 U17456 ( .B1(n14230), .B2(n13958), .A(n20478), .ZN(n13959) );
  OAI21_X1 U17457 ( .B1(n20478), .B2(n20768), .A(n13959), .ZN(P1_U3475) );
  OAI21_X1 U17458 ( .B1(n13962), .B2(n13961), .A(n13960), .ZN(n13963) );
  INV_X1 U17459 ( .A(n13963), .ZN(n20444) );
  NAND2_X1 U17460 ( .A1(n20444), .A2(n20422), .ZN(n13967) );
  INV_X1 U17461 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n13964) );
  NOR2_X1 U17462 ( .A1(n20432), .A2(n13964), .ZN(n20439) );
  NOR2_X1 U17463 ( .A1(n20427), .A2(n20322), .ZN(n13965) );
  AOI211_X1 U17464 ( .C1(n20416), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n20439), .B(n13965), .ZN(n13966) );
  OAI211_X1 U17465 ( .C1(n15258), .C2(n20327), .A(n13967), .B(n13966), .ZN(
        P1_U2996) );
  OR2_X1 U17466 ( .A1(n9799), .A2(n13968), .ZN(n13970) );
  NAND2_X1 U17467 ( .A1(n13970), .A2(n13969), .ZN(n20168) );
  XOR2_X1 U17468 ( .A(n20168), .B(n20167), .Z(n13974) );
  NAND2_X1 U17469 ( .A1(n20178), .A2(n14753), .ZN(n13972) );
  NAND2_X1 U17470 ( .A1(n13972), .A2(n13971), .ZN(n13973) );
  NAND2_X1 U17471 ( .A1(n13974), .A2(n13973), .ZN(n14274) );
  OAI21_X1 U17472 ( .B1(n13974), .B2(n13973), .A(n14274), .ZN(n13975) );
  NAND2_X1 U17473 ( .A1(n13975), .A2(n13177), .ZN(n13978) );
  INV_X1 U17474 ( .A(n19544), .ZN(n13976) );
  AOI22_X1 U17475 ( .A1(n19464), .A2(n13976), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19462), .ZN(n13977) );
  OAI211_X1 U17476 ( .C1(n20168), .C2(n15675), .A(n13978), .B(n13977), .ZN(
        P2_U2916) );
  AND2_X1 U17477 ( .A1(n13980), .A2(n13981), .ZN(n13982) );
  OR2_X1 U17478 ( .A1(n13979), .A2(n13982), .ZN(n16382) );
  AOI21_X1 U17479 ( .B1(n13983), .B2(n14065), .A(n9863), .ZN(n20294) );
  AOI22_X1 U17480 ( .A1(n20294), .A2(n15038), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n15037), .ZN(n13984) );
  OAI21_X1 U17481 ( .B1(n16382), .B2(n15040), .A(n13984), .ZN(P1_U2867) );
  NAND2_X1 U17482 ( .A1(n13838), .A2(n13985), .ZN(n14073) );
  OAI211_X1 U17483 ( .C1(n13987), .C2(n13986), .A(n14073), .B(n14786), .ZN(
        n13992) );
  NOR2_X1 U17484 ( .A1(n13989), .A2(n13943), .ZN(n13990) );
  NAND2_X1 U17485 ( .A1(n14791), .A2(n10090), .ZN(n13991) );
  OAI211_X1 U17486 ( .C1(n14791), .C2(n19359), .A(n13992), .B(n13991), .ZN(
        P2_U2875) );
  NOR2_X1 U17487 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13993), .ZN(n14192) );
  INV_X1 U17488 ( .A(n13994), .ZN(n14061) );
  NAND2_X1 U17489 ( .A1(n13995), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n20217) );
  INV_X1 U17490 ( .A(n13996), .ZN(n14045) );
  NOR2_X1 U17491 ( .A1(n10370), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14008) );
  NAND2_X1 U17492 ( .A1(n11345), .A2(n13997), .ZN(n13998) );
  NAND2_X1 U17493 ( .A1(n13998), .A2(n13115), .ZN(n14014) );
  NAND2_X1 U17494 ( .A1(n14025), .A2(n13999), .ZN(n14011) );
  OAI21_X1 U17495 ( .B1(n14000), .B2(n14008), .A(n14011), .ZN(n14004) );
  INV_X1 U17496 ( .A(n10637), .ZN(n14001) );
  NAND2_X1 U17497 ( .A1(n11344), .A2(n14001), .ZN(n14012) );
  NOR2_X1 U17498 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14002) );
  OR2_X1 U17499 ( .A1(n14012), .A2(n14002), .ZN(n14003) );
  OAI211_X1 U17500 ( .C1(n14008), .C2(n14014), .A(n14004), .B(n14003), .ZN(
        n14005) );
  AOI21_X1 U17501 ( .B1(n12788), .B2(n14045), .A(n14005), .ZN(n14311) );
  INV_X1 U17502 ( .A(n14046), .ZN(n14019) );
  AND2_X1 U17503 ( .A1(n14046), .A2(n14006), .ZN(n14007) );
  AOI21_X1 U17504 ( .B1(n14311), .B2(n14019), .A(n14007), .ZN(n14059) );
  NAND2_X1 U17505 ( .A1(n9734), .A2(n14045), .ZN(n14018) );
  INV_X1 U17506 ( .A(n14008), .ZN(n14013) );
  NAND2_X1 U17507 ( .A1(n11344), .A2(n10637), .ZN(n14009) );
  NAND2_X1 U17508 ( .A1(n14009), .A2(n13115), .ZN(n14010) );
  AOI21_X1 U17509 ( .B1(n14011), .B2(n14013), .A(n14010), .ZN(n14016) );
  AND3_X1 U17510 ( .A1(n14014), .A2(n14013), .A3(n14012), .ZN(n14015) );
  MUX2_X1 U17511 ( .A(n14016), .B(n14015), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n14017) );
  NAND2_X1 U17512 ( .A1(n14018), .A2(n14017), .ZN(n20159) );
  MUX2_X1 U17513 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20159), .S(
        n14019), .Z(n14058) );
  NAND2_X1 U17514 ( .A1(n14046), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14036) );
  NAND2_X1 U17515 ( .A1(n14021), .A2(n14020), .ZN(n14024) );
  NAND2_X1 U17516 ( .A1(n14310), .A2(n14022), .ZN(n14023) );
  OAI211_X1 U17517 ( .C1(n14310), .C2(n14025), .A(n14024), .B(n14023), .ZN(
        n14026) );
  INV_X1 U17518 ( .A(n14026), .ZN(n20210) );
  INV_X1 U17519 ( .A(n10642), .ZN(n14027) );
  AOI22_X1 U17520 ( .A1(n14029), .A2(n14028), .B1(n14027), .B2(n10221), .ZN(
        n14035) );
  INV_X1 U17521 ( .A(n14030), .ZN(n14032) );
  NOR3_X1 U17522 ( .A1(n14033), .A2(n14032), .A3(n14031), .ZN(n19211) );
  OAI21_X1 U17523 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n19211), .ZN(n14034) );
  NAND4_X1 U17524 ( .A1(n14036), .A2(n20210), .A3(n14035), .A4(n14034), .ZN(
        n14057) );
  NOR2_X1 U17525 ( .A1(n14059), .A2(n20182), .ZN(n14050) );
  INV_X1 U17526 ( .A(n11383), .ZN(n14038) );
  NAND2_X1 U17527 ( .A1(n14038), .A2(n14037), .ZN(n14043) );
  OAI21_X1 U17528 ( .B1(n14039), .B2(n10368), .A(n14043), .ZN(n14041) );
  NAND2_X1 U17529 ( .A1(n11344), .A2(n14807), .ZN(n14040) );
  NAND2_X1 U17530 ( .A1(n14041), .A2(n14040), .ZN(n14042) );
  AOI21_X1 U17531 ( .B1(n14327), .B2(n14045), .A(n14042), .ZN(n14803) );
  MUX2_X1 U17532 ( .A(n14043), .B(n11344), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n14044) );
  AOI21_X1 U17533 ( .B1(n14346), .B2(n14045), .A(n14044), .ZN(n14796) );
  OAI211_X1 U17534 ( .C1(n14803), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n14796), .ZN(n14048) );
  AOI21_X1 U17535 ( .B1(n14803), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n14046), .ZN(n14047) );
  NAND2_X1 U17536 ( .A1(n14048), .A2(n14047), .ZN(n14052) );
  INV_X1 U17537 ( .A(n14059), .ZN(n14049) );
  OAI22_X1 U17538 ( .A1(n14050), .A2(n14052), .B1(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n14049), .ZN(n14051) );
  OAI21_X1 U17539 ( .B1(n14051), .B2(n14058), .A(n20175), .ZN(n14055) );
  INV_X1 U17540 ( .A(n14052), .ZN(n14053) );
  NAND3_X1 U17541 ( .A1(n14058), .A2(n14053), .A3(n20182), .ZN(n14054) );
  AOI21_X1 U17542 ( .B1(n14055), .B2(n14054), .A(
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n14056) );
  AOI211_X1 U17543 ( .C1(n14059), .C2(n14058), .A(n14057), .B(n14056), .ZN(
        n16732) );
  AOI21_X1 U17544 ( .B1(n16732), .B2(n14795), .A(n20218), .ZN(n14060) );
  AOI211_X1 U17545 ( .C1(n14192), .C2(n14061), .A(n20217), .B(n14060), .ZN(
        n16729) );
  NOR2_X1 U17546 ( .A1(n16729), .A2(n20218), .ZN(n20077) );
  OAI21_X1 U17547 ( .B1(n20077), .B2(n20195), .A(n16726), .ZN(P2_U3593) );
  OR2_X1 U17548 ( .A1(n14063), .A2(n14062), .ZN(n14064) );
  NAND2_X1 U17549 ( .A1(n14065), .A2(n14064), .ZN(n20433) );
  INV_X1 U17550 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n14069) );
  INV_X1 U17551 ( .A(n13980), .ZN(n14066) );
  AOI21_X1 U17552 ( .B1(n14068), .B2(n14067), .A(n14066), .ZN(n20421) );
  INV_X1 U17553 ( .A(n20421), .ZN(n14096) );
  OAI222_X1 U17554 ( .A1(n20433), .A2(n15048), .B1(n14069), .B2(n15047), .C1(
        n14096), .C2(n15040), .ZN(P1_U2868) );
  INV_X1 U17555 ( .A(n14070), .ZN(n14072) );
  INV_X1 U17556 ( .A(n13988), .ZN(n14071) );
  AOI21_X1 U17557 ( .B1(n14072), .B2(n14071), .A(n14301), .ZN(n19347) );
  INV_X1 U17558 ( .A(n19347), .ZN(n14079) );
  INV_X1 U17559 ( .A(n14073), .ZN(n14076) );
  OAI211_X1 U17560 ( .C1(n14076), .C2(n14075), .A(n14786), .B(n14074), .ZN(
        n14078) );
  NAND2_X1 U17561 ( .A1(n13835), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n14077) );
  OAI211_X1 U17562 ( .C1(n14079), .C2(n13835), .A(n14078), .B(n14077), .ZN(
        P2_U2874) );
  OR2_X1 U17563 ( .A1(n14080), .A2(n14160), .ZN(n14082) );
  OR2_X1 U17564 ( .A1(n14085), .A2(n14084), .ZN(n14087) );
  INV_X1 U17565 ( .A(n14091), .ZN(n14092) );
  NAND2_X1 U17566 ( .A1(n15116), .A2(n14093), .ZN(n15118) );
  OAI222_X1 U17567 ( .A1(n16382), .A2(n15113), .B1(n15088), .B2(n14586), .C1(
        n14095), .C2(n15116), .ZN(P1_U2899) );
  INV_X1 U17568 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20372) );
  OAI222_X1 U17569 ( .A1(n20343), .A2(n15113), .B1(n15108), .B2(n14586), .C1(
        n15116), .C2(n20372), .ZN(P1_U2903) );
  INV_X1 U17570 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20376) );
  OAI222_X1 U17571 ( .A1(n14364), .A2(n15113), .B1(n15117), .B2(n14586), .C1(
        n15116), .C2(n20376), .ZN(P1_U2904) );
  INV_X1 U17572 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20366) );
  OAI222_X1 U17573 ( .A1(n14096), .A2(n15113), .B1(n15093), .B2(n14586), .C1(
        n15116), .C2(n20366), .ZN(P1_U2900) );
  INV_X1 U17574 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20368) );
  OAI222_X1 U17575 ( .A1(n20327), .A2(n15113), .B1(n15098), .B2(n14586), .C1(
        n15116), .C2(n20368), .ZN(P1_U2901) );
  INV_X1 U17576 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20370) );
  OAI222_X1 U17577 ( .A1(n14175), .A2(n15113), .B1(n15103), .B2(n14586), .C1(
        n15116), .C2(n20370), .ZN(P1_U2902) );
  OAI21_X1 U17578 ( .B1(n20774), .B2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n14117), .ZN(n20813) );
  AOI21_X1 U17579 ( .B1(n20649), .B2(n20811), .A(n20810), .ZN(n14102) );
  OR2_X1 U17580 ( .A1(n13542), .A2(n14098), .ZN(n20673) );
  INV_X1 U17581 ( .A(n14099), .ZN(n14100) );
  NAND2_X1 U17582 ( .A1(n14100), .A2(n12024), .ZN(n20876) );
  OR2_X1 U17583 ( .A1(n20673), .A2(n20876), .ZN(n14101) );
  NAND2_X1 U17584 ( .A1(n14101), .A2(n14107), .ZN(n14108) );
  NOR2_X1 U17585 ( .A1(n14102), .A2(n14108), .ZN(n14103) );
  AOI211_X2 U17586 ( .C1(n20676), .C2(n20880), .A(n20813), .B(n14103), .ZN(
        n14156) );
  INV_X1 U17587 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14115) );
  INV_X1 U17588 ( .A(DATAI_20_), .ZN(n21171) );
  INV_X1 U17589 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16768) );
  OAI22_X1 U17590 ( .A1(n21171), .A2(n14146), .B1(n16768), .B2(n14147), .ZN(
        n20913) );
  INV_X1 U17591 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16753) );
  INV_X1 U17592 ( .A(DATAI_28_), .ZN(n21138) );
  OAI22_X1 U17593 ( .A1(n16753), .A2(n14147), .B1(n21138), .B2(n14146), .ZN(
        n20859) );
  INV_X1 U17594 ( .A(n20859), .ZN(n20916) );
  NOR2_X2 U17595 ( .A1(n14149), .A2(n14106), .ZN(n20912) );
  INV_X1 U17596 ( .A(n14107), .ZN(n14151) );
  NAND2_X1 U17597 ( .A1(n14108), .A2(n20811), .ZN(n14111) );
  NAND2_X1 U17598 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n14109), .ZN(n14110) );
  NAND2_X1 U17599 ( .A1(n14111), .A2(n14110), .ZN(n14150) );
  AOI22_X1 U17600 ( .A1(n20912), .A2(n14151), .B1(n20911), .B2(n14150), .ZN(
        n14112) );
  OAI21_X1 U17601 ( .B1(n20916), .B2(n20670), .A(n14112), .ZN(n14113) );
  AOI21_X1 U17602 ( .B1(n20913), .B2(n20729), .A(n14113), .ZN(n14114) );
  OAI21_X1 U17603 ( .B1(n14156), .B2(n14115), .A(n14114), .ZN(P1_U3093) );
  INV_X1 U17604 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14121) );
  INV_X1 U17605 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16765) );
  INV_X1 U17606 ( .A(DATAI_22_), .ZN(n21035) );
  OAI22_X1 U17607 ( .A1(n16765), .A2(n14147), .B1(n21035), .B2(n14146), .ZN(
        n20925) );
  INV_X1 U17608 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n19556) );
  INV_X1 U17609 ( .A(DATAI_30_), .ZN(n14116) );
  OAI22_X1 U17610 ( .A1(n19556), .A2(n14147), .B1(n14116), .B2(n14146), .ZN(
        n20865) );
  INV_X1 U17611 ( .A(n20865), .ZN(n20930) );
  NOR2_X2 U17612 ( .A1(n14149), .A2(n11910), .ZN(n20924) );
  AOI22_X1 U17613 ( .A1(n20924), .A2(n14151), .B1(n20923), .B2(n14150), .ZN(
        n14118) );
  OAI21_X1 U17614 ( .B1(n20930), .B2(n20670), .A(n14118), .ZN(n14119) );
  AOI21_X1 U17615 ( .B1(n20925), .B2(n20729), .A(n14119), .ZN(n14120) );
  OAI21_X1 U17616 ( .B1(n14156), .B2(n14121), .A(n14120), .ZN(P1_U3095) );
  INV_X1 U17617 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14126) );
  INV_X1 U17618 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16763) );
  INV_X1 U17619 ( .A(DATAI_23_), .ZN(n14122) );
  OAI22_X1 U17620 ( .A1(n16763), .A2(n14147), .B1(n14122), .B2(n14146), .ZN(
        n20799) );
  INV_X1 U17621 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16748) );
  INV_X1 U17622 ( .A(DATAI_31_), .ZN(n21140) );
  INV_X1 U17623 ( .A(n20935), .ZN(n20764) );
  NOR2_X2 U17624 ( .A1(n14149), .A2(n15052), .ZN(n20934) );
  AOI22_X1 U17625 ( .A1(n20934), .A2(n14151), .B1(n20932), .B2(n14150), .ZN(
        n14123) );
  OAI21_X1 U17626 ( .B1(n20764), .B2(n20670), .A(n14123), .ZN(n14124) );
  AOI21_X1 U17627 ( .B1(n20799), .B2(n20729), .A(n14124), .ZN(n14125) );
  OAI21_X1 U17628 ( .B1(n14156), .B2(n14126), .A(n14125), .ZN(P1_U3096) );
  INV_X1 U17629 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14131) );
  INV_X1 U17630 ( .A(DATAI_16_), .ZN(n21187) );
  INV_X1 U17631 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16776) );
  OAI22_X1 U17632 ( .A1(n21187), .A2(n14146), .B1(n16776), .B2(n14147), .ZN(
        n20889) );
  INV_X1 U17633 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16761) );
  INV_X1 U17634 ( .A(DATAI_24_), .ZN(n14127) );
  OAI22_X1 U17635 ( .A1(n16761), .A2(n14147), .B1(n14127), .B2(n14146), .ZN(
        n20849) );
  INV_X1 U17636 ( .A(n20849), .ZN(n20892) );
  NOR2_X2 U17637 ( .A1(n14149), .A2(n11941), .ZN(n20883) );
  AOI22_X1 U17638 ( .A1(n20883), .A2(n14151), .B1(n20882), .B2(n14150), .ZN(
        n14128) );
  OAI21_X1 U17639 ( .B1(n20892), .B2(n20670), .A(n14128), .ZN(n14129) );
  AOI21_X1 U17640 ( .B1(n20889), .B2(n20729), .A(n14129), .ZN(n14130) );
  OAI21_X1 U17641 ( .B1(n14156), .B2(n14131), .A(n14130), .ZN(P1_U3089) );
  INV_X1 U17642 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14137) );
  INV_X1 U17643 ( .A(DATAI_17_), .ZN(n21036) );
  INV_X1 U17644 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16774) );
  OAI22_X1 U17645 ( .A1(n21036), .A2(n14146), .B1(n16774), .B2(n14147), .ZN(
        n20781) );
  INV_X1 U17646 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16759) );
  INV_X1 U17647 ( .A(DATAI_25_), .ZN(n14132) );
  OAI22_X2 U17648 ( .A1(n16759), .A2(n14147), .B1(n14132), .B2(n14146), .ZN(
        n20895) );
  INV_X1 U17649 ( .A(n20895), .ZN(n20744) );
  NOR2_X2 U17650 ( .A1(n14149), .A2(n14133), .ZN(n20894) );
  AOI22_X1 U17651 ( .A1(n20894), .A2(n14151), .B1(n20893), .B2(n14150), .ZN(
        n14134) );
  OAI21_X1 U17652 ( .B1(n20744), .B2(n20670), .A(n14134), .ZN(n14135) );
  AOI21_X1 U17653 ( .B1(n20781), .B2(n20729), .A(n14135), .ZN(n14136) );
  OAI21_X1 U17654 ( .B1(n14156), .B2(n14137), .A(n14136), .ZN(P1_U3090) );
  INV_X1 U17655 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14141) );
  INV_X1 U17656 ( .A(DATAI_18_), .ZN(n21198) );
  INV_X1 U17657 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16772) );
  OAI22_X1 U17658 ( .A1(n21198), .A2(n14146), .B1(n16772), .B2(n14147), .ZN(
        n20784) );
  INV_X1 U17659 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16757) );
  INV_X1 U17660 ( .A(DATAI_26_), .ZN(n21177) );
  INV_X1 U17661 ( .A(n20901), .ZN(n20747) );
  NOR2_X2 U17662 ( .A1(n14149), .A2(n12770), .ZN(n20900) );
  AOI22_X1 U17663 ( .A1(n20900), .A2(n14151), .B1(n20899), .B2(n14150), .ZN(
        n14138) );
  OAI21_X1 U17664 ( .B1(n20747), .B2(n20670), .A(n14138), .ZN(n14139) );
  AOI21_X1 U17665 ( .B1(n20784), .B2(n20729), .A(n14139), .ZN(n14140) );
  OAI21_X1 U17666 ( .B1(n14156), .B2(n14141), .A(n14140), .ZN(P1_U3091) );
  INV_X1 U17667 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14145) );
  INV_X1 U17668 ( .A(DATAI_19_), .ZN(n21042) );
  INV_X1 U17669 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16770) );
  OAI22_X1 U17670 ( .A1(n21042), .A2(n14146), .B1(n16770), .B2(n14147), .ZN(
        n20787) );
  INV_X1 U17671 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16755) );
  INV_X1 U17672 ( .A(DATAI_27_), .ZN(n21209) );
  OAI22_X2 U17673 ( .A1(n16755), .A2(n14147), .B1(n21209), .B2(n14146), .ZN(
        n20907) );
  INV_X1 U17674 ( .A(n20907), .ZN(n20750) );
  NOR2_X2 U17675 ( .A1(n14149), .A2(n12636), .ZN(n20906) );
  AOI22_X1 U17676 ( .A1(n20906), .A2(n14151), .B1(n20905), .B2(n14150), .ZN(
        n14142) );
  OAI21_X1 U17677 ( .B1(n20750), .B2(n20670), .A(n14142), .ZN(n14143) );
  AOI21_X1 U17678 ( .B1(n20787), .B2(n20729), .A(n14143), .ZN(n14144) );
  OAI21_X1 U17679 ( .B1(n14156), .B2(n14145), .A(n14144), .ZN(P1_U3092) );
  INV_X1 U17680 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14155) );
  INV_X1 U17681 ( .A(DATAI_21_), .ZN(n21193) );
  INV_X1 U17682 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n19550) );
  OAI22_X1 U17683 ( .A1(n21193), .A2(n14146), .B1(n19550), .B2(n14147), .ZN(
        n20792) );
  INV_X1 U17684 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16751) );
  INV_X1 U17685 ( .A(DATAI_29_), .ZN(n21201) );
  OAI22_X2 U17686 ( .A1(n16751), .A2(n14147), .B1(n21201), .B2(n14146), .ZN(
        n20919) );
  INV_X1 U17687 ( .A(n20919), .ZN(n20755) );
  NOR2_X2 U17688 ( .A1(n14149), .A2(n14148), .ZN(n20918) );
  AOI22_X1 U17689 ( .A1(n20918), .A2(n14151), .B1(n20917), .B2(n14150), .ZN(
        n14152) );
  OAI21_X1 U17690 ( .B1(n20755), .B2(n20670), .A(n14152), .ZN(n14153) );
  AOI21_X1 U17691 ( .B1(n20792), .B2(n20729), .A(n14153), .ZN(n14154) );
  OAI21_X1 U17692 ( .B1(n14156), .B2(n14155), .A(n14154), .ZN(P1_U3094) );
  OAI21_X1 U17693 ( .B1(n14159), .B2(n14157), .A(n14158), .ZN(n19352) );
  OAI222_X1 U17694 ( .A1(n14356), .A2(n15622), .B1(n19352), .B2(n19471), .C1(
        n13426), .C2(n15689), .ZN(P2_U2906) );
  NOR2_X1 U17695 ( .A1(n14163), .A2(n14160), .ZN(n14161) );
  OR2_X1 U17696 ( .A1(n20287), .A2(n14161), .ZN(n20315) );
  INV_X1 U17697 ( .A(n13542), .ZN(n14390) );
  NOR2_X1 U17698 ( .A1(n14163), .A2(n14162), .ZN(n20346) );
  AOI21_X1 U17699 ( .B1(n20347), .B2(n13702), .A(n20276), .ZN(n20326) );
  INV_X1 U17700 ( .A(n14164), .ZN(n14169) );
  INV_X1 U17701 ( .A(n14165), .ZN(n14166) );
  NAND2_X1 U17702 ( .A1(n20347), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20333) );
  OAI22_X1 U17703 ( .A1(n20335), .A2(n14167), .B1(P1_REIP_REG_2__SCAN_IN), 
        .B2(n20333), .ZN(n14168) );
  AOI21_X1 U17704 ( .B1(n14169), .B2(n20338), .A(n14168), .ZN(n14172) );
  AOI22_X1 U17705 ( .A1(n20321), .A2(P1_EBX_REG_2__SCAN_IN), .B1(n20320), .B2(
        n14170), .ZN(n14171) );
  OAI211_X1 U17706 ( .C1(n20326), .C2(n13892), .A(n14172), .B(n14171), .ZN(
        n14173) );
  AOI21_X1 U17707 ( .B1(n14390), .B2(n20346), .A(n14173), .ZN(n14174) );
  OAI21_X1 U17708 ( .B1(n14175), .B2(n20342), .A(n14174), .ZN(P1_U2838) );
  NAND2_X1 U17709 ( .A1(n19208), .A2(n10646), .ZN(n14188) );
  INV_X1 U17710 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16472) );
  AND2_X1 U17711 ( .A1(n20226), .A2(n20221), .ZN(n14176) );
  INV_X1 U17712 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14838) );
  INV_X1 U17713 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14677) );
  NOR2_X2 U17714 ( .A1(n14678), .A2(n14677), .ZN(n14177) );
  XNOR2_X1 U17715 ( .A(n14177), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n15698) );
  AOI21_X1 U17716 ( .B1(n19381), .B2(n14183), .A(n14185), .ZN(n19386) );
  AOI21_X1 U17717 ( .B1(n19396), .B2(n14181), .A(n14184), .ZN(n19394) );
  AOI21_X1 U17718 ( .B1(n16665), .B2(n14179), .A(n14182), .ZN(n19440) );
  AOI21_X1 U17719 ( .B1(n16678), .B2(n14178), .A(n14180), .ZN(n16666) );
  OAI22_X1 U17720 ( .A1(n20218), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n14309) );
  OAI22_X1 U17721 ( .A1(n20218), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n14319), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14307) );
  AND2_X1 U17722 ( .A1(n14309), .A2(n14307), .ZN(n14306) );
  OAI21_X1 U17723 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n14178), .ZN(n14773) );
  NAND2_X1 U17724 ( .A1(n14306), .A2(n14773), .ZN(n14286) );
  NOR2_X1 U17725 ( .A1(n16666), .A2(n14286), .ZN(n14215) );
  OAI21_X1 U17726 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n14180), .A(
        n14179), .ZN(n19509) );
  NAND2_X1 U17727 ( .A1(n14215), .A2(n19509), .ZN(n19438) );
  NOR2_X1 U17728 ( .A1(n19440), .A2(n19438), .ZN(n19418) );
  OAI21_X1 U17729 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n14182), .A(
        n14181), .ZN(n19421) );
  NAND2_X1 U17730 ( .A1(n19418), .A2(n19421), .ZN(n19392) );
  NOR2_X1 U17731 ( .A1(n19394), .A2(n19392), .ZN(n14204) );
  OAI21_X1 U17732 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n14184), .A(
        n14183), .ZN(n16659) );
  NAND2_X1 U17733 ( .A1(n14204), .A2(n16659), .ZN(n19383) );
  NOR2_X1 U17734 ( .A1(n19386), .A2(n19383), .ZN(n15514) );
  NOR2_X1 U17735 ( .A1(n19419), .A2(n15514), .ZN(n14186) );
  OAI21_X1 U17736 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n14185), .A(
        n15513), .ZN(n16632) );
  XNOR2_X1 U17737 ( .A(n14186), .B(n16632), .ZN(n14187) );
  NAND4_X1 U17738 ( .A1(n20218), .A2(n19942), .A3(n20226), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19411) );
  NAND2_X1 U17739 ( .A1(n14187), .A2(n19443), .ZN(n14202) );
  OAI21_X1 U17740 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n20215), .A(n16472), 
        .ZN(n14189) );
  INV_X1 U17741 ( .A(n14189), .ZN(n14190) );
  AND2_X1 U17742 ( .A1(n14191), .A2(n14190), .ZN(n14194) );
  INV_X1 U17743 ( .A(n14192), .ZN(n14193) );
  OAI21_X1 U17744 ( .B1(n14195), .B2(n14194), .A(n14193), .ZN(n19413) );
  AND2_X1 U17745 ( .A1(n19942), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20079) );
  NAND2_X1 U17746 ( .A1(n14196), .A2(n20079), .ZN(n16725) );
  NAND2_X1 U17747 ( .A1(n16725), .A2(n19341), .ZN(n14197) );
  OR3_X2 U17748 ( .A1(n19208), .A2(n19443), .A3(n14197), .ZN(n19417) );
  INV_X1 U17749 ( .A(n19417), .ZN(n19437) );
  AOI22_X1 U17750 ( .A1(n19432), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19437), .ZN(n14199) );
  AOI21_X1 U17751 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19431), .A(
        n19500), .ZN(n14198) );
  OAI211_X1 U17752 ( .C1(n19447), .C2(n16691), .A(n14199), .B(n14198), .ZN(
        n14200) );
  AOI21_X1 U17753 ( .B1(n16698), .B2(n19441), .A(n14200), .ZN(n14201) );
  OAI211_X1 U17754 ( .C1(n19434), .C2(n14203), .A(n14202), .B(n14201), .ZN(
        P2_U2845) );
  NOR2_X1 U17755 ( .A1(n19419), .A2(n14204), .ZN(n14205) );
  XNOR2_X1 U17756 ( .A(n14205), .B(n16659), .ZN(n14206) );
  NAND2_X1 U17757 ( .A1(n14206), .A2(n19443), .ZN(n14213) );
  OAI21_X1 U17758 ( .B1(n11438), .B2(n19417), .A(n19395), .ZN(n14207) );
  AOI21_X1 U17759 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19431), .A(
        n14207), .ZN(n14209) );
  NAND2_X1 U17760 ( .A1(n19361), .A2(n16709), .ZN(n14208) );
  OAI211_X1 U17761 ( .C1(n19413), .C2(n10680), .A(n14209), .B(n14208), .ZN(
        n14210) );
  AOI21_X1 U17762 ( .B1(n14211), .B2(n19441), .A(n14210), .ZN(n14212) );
  OAI211_X1 U17763 ( .C1(n19434), .C2(n14214), .A(n14213), .B(n14212), .ZN(
        P2_U2847) );
  NOR2_X1 U17764 ( .A1(n19419), .A2(n14215), .ZN(n14216) );
  XNOR2_X1 U17765 ( .A(n19509), .B(n14216), .ZN(n14217) );
  NAND2_X1 U17766 ( .A1(n14217), .A2(n19443), .ZN(n14229) );
  INV_X1 U17767 ( .A(n13969), .ZN(n14218) );
  XNOR2_X1 U17768 ( .A(n14219), .B(n14218), .ZN(n16083) );
  INV_X1 U17769 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n14220) );
  OAI21_X1 U17770 ( .B1(n19397), .B2(n14220), .A(n19341), .ZN(n14224) );
  OAI22_X1 U17771 ( .A1(n19400), .A2(n14222), .B1(n14221), .B2(n19417), .ZN(
        n14223) );
  AOI211_X1 U17772 ( .C1(n16083), .C2(n19361), .A(n14224), .B(n14223), .ZN(
        n14225) );
  OAI21_X1 U17773 ( .B1(n14226), .B2(n19434), .A(n14225), .ZN(n14227) );
  AOI21_X1 U17774 ( .B1(n19503), .B2(n19441), .A(n14227), .ZN(n14228) );
  OAI211_X1 U17775 ( .C1(n14752), .C2(n19466), .A(n14229), .B(n14228), .ZN(
        P2_U2851) );
  NAND3_X1 U17776 ( .A1(n14230), .A2(n13949), .A3(n20810), .ZN(n14231) );
  OR3_X1 U17777 ( .A1(n16225), .A2(n20768), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14499) );
  INV_X1 U17778 ( .A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14242) );
  NOR2_X1 U17779 ( .A1(n20733), .A2(n14499), .ZN(n14268) );
  OR2_X1 U17780 ( .A1(n13542), .A2(n14233), .ZN(n20840) );
  INV_X1 U17781 ( .A(n14268), .ZN(n14234) );
  OAI21_X1 U17782 ( .B1(n20840), .B2(n20503), .A(n14234), .ZN(n14235) );
  NAND2_X1 U17783 ( .A1(n14235), .A2(n20811), .ZN(n14238) );
  INV_X1 U17784 ( .A(n14499), .ZN(n14236) );
  NAND2_X1 U17785 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n14236), .ZN(n14237) );
  NAND2_X1 U17786 ( .A1(n14238), .A2(n14237), .ZN(n14267) );
  AOI22_X1 U17787 ( .A1(n20900), .A2(n14268), .B1(n20899), .B2(n14267), .ZN(
        n14239) );
  OAI21_X1 U17788 ( .B1(n20747), .B2(n14543), .A(n14239), .ZN(n14240) );
  AOI21_X1 U17789 ( .B1(n20871), .B2(n20784), .A(n14240), .ZN(n14241) );
  OAI21_X1 U17790 ( .B1(n14273), .B2(n14242), .A(n14241), .ZN(P1_U3139) );
  INV_X1 U17791 ( .A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14246) );
  AOI22_X1 U17792 ( .A1(n20894), .A2(n14268), .B1(n20893), .B2(n14267), .ZN(
        n14243) );
  OAI21_X1 U17793 ( .B1(n20744), .B2(n14543), .A(n14243), .ZN(n14244) );
  AOI21_X1 U17794 ( .B1(n20871), .B2(n20781), .A(n14244), .ZN(n14245) );
  OAI21_X1 U17795 ( .B1(n14273), .B2(n14246), .A(n14245), .ZN(P1_U3138) );
  INV_X1 U17796 ( .A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14250) );
  AOI22_X1 U17797 ( .A1(n20883), .A2(n14268), .B1(n20882), .B2(n14267), .ZN(
        n14247) );
  OAI21_X1 U17798 ( .B1(n20892), .B2(n14543), .A(n14247), .ZN(n14248) );
  AOI21_X1 U17799 ( .B1(n20871), .B2(n20889), .A(n14248), .ZN(n14249) );
  OAI21_X1 U17800 ( .B1(n14273), .B2(n14250), .A(n14249), .ZN(P1_U3137) );
  INV_X1 U17801 ( .A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14254) );
  AOI22_X1 U17802 ( .A1(n20934), .A2(n14268), .B1(n20932), .B2(n14267), .ZN(
        n14251) );
  OAI21_X1 U17803 ( .B1(n20764), .B2(n14543), .A(n14251), .ZN(n14252) );
  AOI21_X1 U17804 ( .B1(n20871), .B2(n20799), .A(n14252), .ZN(n14253) );
  OAI21_X1 U17805 ( .B1(n14273), .B2(n14254), .A(n14253), .ZN(P1_U3144) );
  INV_X1 U17806 ( .A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14258) );
  AOI22_X1 U17807 ( .A1(n20924), .A2(n14268), .B1(n20923), .B2(n14267), .ZN(
        n14255) );
  OAI21_X1 U17808 ( .B1(n20930), .B2(n14543), .A(n14255), .ZN(n14256) );
  AOI21_X1 U17809 ( .B1(n20871), .B2(n20925), .A(n14256), .ZN(n14257) );
  OAI21_X1 U17810 ( .B1(n14273), .B2(n14258), .A(n14257), .ZN(P1_U3143) );
  INV_X1 U17811 ( .A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14262) );
  AOI22_X1 U17812 ( .A1(n20918), .A2(n14268), .B1(n20917), .B2(n14267), .ZN(
        n14259) );
  OAI21_X1 U17813 ( .B1(n20755), .B2(n14543), .A(n14259), .ZN(n14260) );
  AOI21_X1 U17814 ( .B1(n20871), .B2(n20792), .A(n14260), .ZN(n14261) );
  OAI21_X1 U17815 ( .B1(n14273), .B2(n14262), .A(n14261), .ZN(P1_U3142) );
  INV_X1 U17816 ( .A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14266) );
  AOI22_X1 U17817 ( .A1(n20912), .A2(n14268), .B1(n20911), .B2(n14267), .ZN(
        n14263) );
  OAI21_X1 U17818 ( .B1(n20916), .B2(n14543), .A(n14263), .ZN(n14264) );
  AOI21_X1 U17819 ( .B1(n20913), .B2(n20871), .A(n14264), .ZN(n14265) );
  OAI21_X1 U17820 ( .B1(n14273), .B2(n14266), .A(n14265), .ZN(P1_U3141) );
  INV_X1 U17821 ( .A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14272) );
  AOI22_X1 U17822 ( .A1(n20906), .A2(n14268), .B1(n20905), .B2(n14267), .ZN(
        n14269) );
  OAI21_X1 U17823 ( .B1(n20750), .B2(n14543), .A(n14269), .ZN(n14270) );
  AOI21_X1 U17824 ( .B1(n20871), .B2(n20787), .A(n14270), .ZN(n14271) );
  OAI21_X1 U17825 ( .B1(n14273), .B2(n14272), .A(n14271), .ZN(P1_U3140) );
  NAND2_X1 U17826 ( .A1(n20167), .A2(n20168), .ZN(n14275) );
  AOI21_X1 U17827 ( .B1(n14275), .B2(n14274), .A(n16083), .ZN(n19467) );
  XNOR2_X1 U17828 ( .A(n19467), .B(n19466), .ZN(n14279) );
  OAI22_X1 U17829 ( .A1(n14356), .A2(n19547), .B1(n15689), .B2(n14276), .ZN(
        n14277) );
  AOI21_X1 U17830 ( .B1(n19449), .B2(n16083), .A(n14277), .ZN(n14278) );
  OAI21_X1 U17831 ( .B1(n14279), .B2(n19465), .A(n14278), .ZN(P2_U2915) );
  OR2_X1 U17832 ( .A1(n13979), .A2(n14281), .ZN(n14282) );
  AND2_X1 U17833 ( .A1(n14280), .A2(n14282), .ZN(n20288) );
  INV_X1 U17834 ( .A(n20288), .ZN(n14297) );
  XNOR2_X1 U17835 ( .A(n14284), .B(n14283), .ZN(n20282) );
  AOI22_X1 U17836 ( .A1(n20282), .A2(n15038), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n15037), .ZN(n14285) );
  OAI21_X1 U17837 ( .B1(n14297), .B2(n15040), .A(n14285), .ZN(P1_U2866) );
  NAND2_X1 U17838 ( .A1(n19384), .A2(n14286), .ZN(n14287) );
  XNOR2_X1 U17839 ( .A(n16666), .B(n14287), .ZN(n14294) );
  OAI22_X1 U17840 ( .A1(n19417), .A2(n11419), .B1(n19397), .B2(n16678), .ZN(
        n14290) );
  NOR2_X1 U17841 ( .A1(n19434), .A2(n14288), .ZN(n14289) );
  AOI211_X1 U17842 ( .C1(n19432), .C2(P2_EBX_REG_3__SCAN_IN), .A(n14290), .B(
        n14289), .ZN(n14292) );
  NAND2_X1 U17843 ( .A1(n9734), .A2(n19441), .ZN(n14291) );
  OAI211_X1 U17844 ( .C1(n20168), .C2(n19447), .A(n14292), .B(n14291), .ZN(
        n14293) );
  AOI21_X1 U17845 ( .B1(n14294), .B2(n19443), .A(n14293), .ZN(n14295) );
  OAI21_X1 U17846 ( .B1(n20167), .B2(n14752), .A(n14295), .ZN(P2_U2852) );
  INV_X1 U17847 ( .A(n15081), .ZN(n14296) );
  OAI222_X1 U17848 ( .A1(n14297), .A2(n15113), .B1(n14296), .B2(n14586), .C1(
        n20363), .C2(n15116), .ZN(P1_U2898) );
  INV_X1 U17849 ( .A(n14074), .ZN(n14299) );
  OAI211_X1 U17850 ( .C1(n14299), .C2(n9744), .A(n10031), .B(n14786), .ZN(
        n14304) );
  OR2_X1 U17851 ( .A1(n14301), .A2(n14300), .ZN(n14302) );
  AND2_X1 U17852 ( .A1(n14302), .A2(n14333), .ZN(n19332) );
  NAND2_X1 U17853 ( .A1(n19332), .A2(n15616), .ZN(n14303) );
  OAI211_X1 U17854 ( .C1(n14791), .C2(n10768), .A(n14304), .B(n14303), .ZN(
        P2_U2873) );
  NOR2_X1 U17855 ( .A1(n19419), .A2(n14306), .ZN(n14741) );
  OAI21_X1 U17856 ( .B1(n14309), .B2(n14307), .A(n14741), .ZN(n14316) );
  OAI21_X1 U17857 ( .B1(n19384), .B2(n14308), .A(n14316), .ZN(n14802) );
  INV_X1 U17858 ( .A(n14309), .ZN(n14351) );
  AOI22_X1 U17859 ( .A1(n19419), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n14351), .B2(n19384), .ZN(n14793) );
  NOR2_X1 U17860 ( .A1(n14793), .A2(n14795), .ZN(n14800) );
  OAI22_X1 U17861 ( .A1(n20178), .A2(n20161), .B1(n20165), .B2(n14311), .ZN(
        n14312) );
  AOI21_X1 U17862 ( .B1(n14802), .B2(n14800), .A(n14312), .ZN(n14315) );
  NAND2_X1 U17863 ( .A1(n14314), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14313) );
  OAI21_X1 U17864 ( .B1(n14315), .B2(n14314), .A(n14313), .ZN(P2_U3599) );
  NOR2_X1 U17865 ( .A1(n19384), .A2(n19411), .ZN(n19349) );
  INV_X1 U17866 ( .A(n19349), .ZN(n19259) );
  OAI22_X1 U17867 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19259), .B1(
        n14316), .B2(n19411), .ZN(n14317) );
  INV_X1 U17868 ( .A(n14317), .ZN(n14329) );
  INV_X1 U17869 ( .A(n14318), .ZN(n14323) );
  OAI22_X1 U17870 ( .A1(n19417), .A2(n20102), .B1(n19397), .B2(n14319), .ZN(
        n14322) );
  NOR2_X1 U17871 ( .A1(n19400), .A2(n14320), .ZN(n14321) );
  AOI211_X1 U17872 ( .C1(n14323), .C2(n19403), .A(n14322), .B(n14321), .ZN(
        n14324) );
  OAI21_X1 U17873 ( .B1(n19447), .B2(n14325), .A(n14324), .ZN(n14326) );
  AOI21_X1 U17874 ( .B1(n14327), .B2(n19441), .A(n14326), .ZN(n14328) );
  OAI211_X1 U17875 ( .C1(n19513), .C2(n14752), .A(n14329), .B(n14328), .ZN(
        P2_U2854) );
  INV_X1 U17876 ( .A(n14330), .ZN(n14334) );
  INV_X1 U17877 ( .A(n14331), .ZN(n14332) );
  AOI21_X1 U17878 ( .B1(n14334), .B2(n14333), .A(n14332), .ZN(n19322) );
  INV_X1 U17879 ( .A(n19322), .ZN(n14339) );
  OAI211_X1 U17880 ( .C1(n14298), .C2(n14336), .A(n10030), .B(n14786), .ZN(
        n14338) );
  NAND2_X1 U17881 ( .A1(n13835), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n14337) );
  OAI211_X1 U17882 ( .C1(n14339), .C2(n13835), .A(n14338), .B(n14337), .ZN(
        P2_U2872) );
  NOR2_X1 U17883 ( .A1(n19411), .A2(n19419), .ZN(n19235) );
  AOI22_X1 U17884 ( .A1(n19437), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19361), 
        .B2(n14340), .ZN(n14343) );
  NAND2_X1 U17885 ( .A1(n19403), .A2(n14341), .ZN(n14342) );
  OAI211_X1 U17886 ( .C1(n19400), .C2(n14344), .A(n14343), .B(n14342), .ZN(
        n14345) );
  AOI21_X1 U17887 ( .B1(n14346), .B2(n19441), .A(n14345), .ZN(n14347) );
  OAI21_X1 U17888 ( .B1(n20197), .B2(n14752), .A(n14347), .ZN(n14350) );
  OAI21_X1 U17889 ( .B1(n19431), .B2(n19349), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14348) );
  INV_X1 U17890 ( .A(n14348), .ZN(n14349) );
  AOI211_X1 U17891 ( .C1(n19235), .C2(n14351), .A(n14350), .B(n14349), .ZN(
        n14352) );
  INV_X1 U17892 ( .A(n14352), .ZN(P2_U2855) );
  OAI21_X1 U17893 ( .B1(n14353), .B2(n14354), .A(n9777), .ZN(n19326) );
  OAI222_X1 U17894 ( .A1(n14356), .A2(n14355), .B1(n19326), .B2(n19471), .C1(
        n13453), .C2(n15689), .ZN(P2_U2904) );
  OR2_X1 U17895 ( .A1(n14280), .A2(n14357), .ZN(n14404) );
  NAND2_X1 U17896 ( .A1(n14280), .A2(n14357), .ZN(n14358) );
  INV_X1 U17897 ( .A(n20278), .ZN(n14359) );
  OAI222_X1 U17898 ( .A1(n14359), .A2(n15113), .B1(n15076), .B2(n14586), .C1(
        n15116), .C2(n12137), .ZN(P1_U2897) );
  NOR2_X1 U17899 ( .A1(n20347), .A2(n20276), .ZN(n20312) );
  INV_X1 U17900 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n14363) );
  INV_X1 U17901 ( .A(n20468), .ZN(n14360) );
  AOI22_X1 U17902 ( .A1(n20321), .A2(P1_EBX_REG_0__SCAN_IN), .B1(n20320), .B2(
        n14360), .ZN(n14362) );
  OAI21_X1 U17903 ( .B1(n20338), .B2(n20323), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14361) );
  OAI211_X1 U17904 ( .C1(n20312), .C2(n14363), .A(n14362), .B(n14361), .ZN(
        n14366) );
  NOR2_X1 U17905 ( .A1(n14364), .A2(n20342), .ZN(n14365) );
  AOI211_X1 U17906 ( .C1(n20346), .C2(n12024), .A(n14366), .B(n14365), .ZN(
        n14367) );
  INV_X1 U17907 ( .A(n14367), .ZN(P1_U2840) );
  NAND2_X1 U17908 ( .A1(n14369), .A2(n14368), .ZN(n14371) );
  XNOR2_X1 U17909 ( .A(n14371), .B(n14370), .ZN(n16672) );
  INV_X1 U17910 ( .A(n15964), .ZN(n14757) );
  AOI21_X1 U17911 ( .B1(n14757), .B2(n14759), .A(n14372), .ZN(n14460) );
  INV_X1 U17912 ( .A(n14460), .ZN(n14374) );
  NOR2_X1 U17913 ( .A1(n14454), .A2(n14759), .ZN(n14373) );
  MUX2_X1 U17914 ( .A(n14374), .B(n14373), .S(n14453), .Z(n14375) );
  AOI21_X1 U17915 ( .B1(n19500), .B2(P2_REIP_REG_3__SCAN_IN), .A(n14375), .ZN(
        n14376) );
  OAI21_X1 U17916 ( .B1(n20168), .B2(n16072), .A(n14376), .ZN(n14380) );
  INV_X1 U17917 ( .A(n14378), .ZN(n16669) );
  NOR3_X1 U17918 ( .A1(n16670), .A2(n16669), .A3(n16717), .ZN(n14379) );
  AOI211_X1 U17919 ( .C1(n16699), .C2(n9734), .A(n14380), .B(n14379), .ZN(
        n14381) );
  OAI21_X1 U17920 ( .B1(n16672), .B2(n16704), .A(n14381), .ZN(P2_U3043) );
  INV_X1 U17921 ( .A(n15040), .ZN(n15050) );
  OR2_X1 U17922 ( .A1(n14383), .A2(n14382), .ZN(n14384) );
  NAND2_X1 U17923 ( .A1(n14407), .A2(n14384), .ZN(n20268) );
  OAI22_X1 U17924 ( .A1(n20268), .A2(n15048), .B1(n20272), .B2(n15047), .ZN(
        n14385) );
  AOI21_X1 U17925 ( .B1(n20278), .B2(n15050), .A(n14385), .ZN(n14386) );
  INV_X1 U17926 ( .A(n14386), .ZN(P1_U2865) );
  NAND2_X1 U17927 ( .A1(n14497), .A2(n20769), .ZN(n20619) );
  NOR3_X1 U17928 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20508) );
  INV_X1 U17929 ( .A(n20508), .ZN(n20505) );
  NOR2_X1 U17930 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20505), .ZN(
        n20497) );
  INV_X1 U17931 ( .A(n14396), .ZN(n14387) );
  NOR2_X1 U17932 ( .A1(n14387), .A2(n12006), .ZN(n20674) );
  OAI21_X1 U17933 ( .B1(n20497), .B2(n20774), .A(n20773), .ZN(n14394) );
  OAI21_X1 U17934 ( .B1(n20526), .B2(n20926), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n14389) );
  NAND2_X1 U17935 ( .A1(n14389), .A2(n20811), .ZN(n14398) );
  OR2_X1 U17936 ( .A1(n13856), .A2(n14390), .ZN(n20568) );
  INV_X1 U17937 ( .A(n14392), .ZN(n20841) );
  NOR2_X1 U17938 ( .A1(n20568), .A2(n20841), .ZN(n14395) );
  NOR2_X1 U17939 ( .A1(n14398), .A2(n14395), .ZN(n14393) );
  INV_X1 U17940 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n14402) );
  INV_X1 U17941 ( .A(n14395), .ZN(n14397) );
  NOR2_X1 U17942 ( .A1(n14396), .A2(n12006), .ZN(n20771) );
  INV_X1 U17943 ( .A(n20771), .ZN(n20708) );
  OAI22_X1 U17944 ( .A1(n14398), .A2(n14397), .B1(n20619), .B2(n20708), .ZN(
        n20499) );
  AOI22_X1 U17945 ( .A1(n20526), .A2(n20913), .B1(n20912), .B2(n20497), .ZN(
        n14399) );
  OAI21_X1 U17946 ( .B1(n20940), .B2(n20916), .A(n14399), .ZN(n14400) );
  AOI21_X1 U17947 ( .B1(n20499), .B2(n20911), .A(n14400), .ZN(n14401) );
  OAI21_X1 U17948 ( .B1(n20498), .B2(n14402), .A(n14401), .ZN(P1_U3037) );
  INV_X1 U17949 ( .A(n14427), .ZN(n14403) );
  AOI21_X1 U17950 ( .B1(n14405), .B2(n14404), .A(n14403), .ZN(n14483) );
  INV_X1 U17951 ( .A(n14483), .ZN(n14419) );
  OAI21_X1 U17952 ( .B1(n14972), .B2(n14406), .A(n20334), .ZN(n20263) );
  INV_X1 U17953 ( .A(n14407), .ZN(n14409) );
  OAI21_X1 U17954 ( .B1(n14409), .B2(n14408), .A(n14431), .ZN(n16429) );
  AOI22_X1 U17955 ( .A1(n20321), .A2(P1_EBX_REG_8__SCAN_IN), .B1(n20338), .B2(
        n14482), .ZN(n14414) );
  NAND2_X1 U17956 ( .A1(n20334), .A2(n14410), .ZN(n20289) );
  NAND3_X1 U17957 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n14411) );
  NOR2_X1 U17958 ( .A1(n14972), .A2(n20275), .ZN(n20301) );
  INV_X1 U17959 ( .A(n20301), .ZN(n20255) );
  NOR3_X1 U17960 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n14411), .A3(n20255), .ZN(
        n14412) );
  AOI211_X1 U17961 ( .C1(n20323), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n20310), .B(n14412), .ZN(n14413) );
  OAI211_X1 U17962 ( .C1(n20351), .C2(n16429), .A(n14414), .B(n14413), .ZN(
        n14415) );
  AOI21_X1 U17963 ( .B1(P1_REIP_REG_8__SCAN_IN), .B2(n20263), .A(n14415), .ZN(
        n14416) );
  OAI21_X1 U17964 ( .B1(n14419), .B2(n16324), .A(n14416), .ZN(P1_U2832) );
  INV_X1 U17965 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14417) );
  OAI222_X1 U17966 ( .A1(n14419), .A2(n15040), .B1(n15047), .B2(n14417), .C1(
        n16429), .C2(n15048), .ZN(P1_U2864) );
  INV_X1 U17967 ( .A(DATAI_8_), .ZN(n21202) );
  INV_X1 U17968 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16790) );
  MUX2_X1 U17969 ( .A(n21202), .B(n16790), .S(n14699), .Z(n20377) );
  INV_X1 U17970 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14418) );
  OAI222_X1 U17971 ( .A1(n14419), .A2(n15113), .B1(n20377), .B2(n14586), .C1(
        n14418), .C2(n15116), .ZN(P1_U2896) );
  OAI21_X1 U17972 ( .B1(n14335), .B2(n14421), .A(n14420), .ZN(n14440) );
  NAND2_X1 U17973 ( .A1(n14331), .A2(n14422), .ZN(n14423) );
  NAND2_X1 U17974 ( .A1(n14472), .A2(n14423), .ZN(n15978) );
  MUX2_X1 U17975 ( .A(n14424), .B(n15978), .S(n15616), .Z(n14425) );
  OAI21_X1 U17976 ( .B1(n14440), .B2(n15618), .A(n14425), .ZN(P2_U2871) );
  NAND2_X1 U17977 ( .A1(n14427), .A2(n14426), .ZN(n14428) );
  NAND2_X1 U17978 ( .A1(n14555), .A2(n14428), .ZN(n20262) );
  INV_X1 U17979 ( .A(n14558), .ZN(n14429) );
  AOI21_X1 U17980 ( .B1(n14431), .B2(n14430), .A(n14429), .ZN(n20257) );
  AOI22_X1 U17981 ( .A1(n20257), .A2(n15038), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n15037), .ZN(n14432) );
  OAI21_X1 U17982 ( .B1(n20262), .B2(n15040), .A(n14432), .ZN(P1_U2863) );
  AND2_X1 U17983 ( .A1(n9777), .A2(n14434), .ZN(n14435) );
  NOR2_X1 U17984 ( .A1(n14433), .A2(n14435), .ZN(n19310) );
  OAI22_X1 U17985 ( .A1(n19523), .A2(n15690), .B1(n15689), .B2(n13490), .ZN(
        n14438) );
  INV_X1 U17986 ( .A(n19451), .ZN(n15693) );
  INV_X1 U17987 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n14436) );
  OAI22_X1 U17988 ( .A1(n15693), .A2(n16776), .B1(n15692), .B2(n14436), .ZN(
        n14437) );
  AOI211_X1 U17989 ( .C1(n19310), .C2(n19449), .A(n14438), .B(n14437), .ZN(
        n14439) );
  OAI21_X1 U17990 ( .B1(n19465), .B2(n14440), .A(n14439), .ZN(P2_U2903) );
  INV_X1 U17991 ( .A(DATAI_9_), .ZN(n21168) );
  INV_X1 U17992 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16788) );
  MUX2_X1 U17993 ( .A(n21168), .B(n16788), .S(n14699), .Z(n20380) );
  INV_X1 U17994 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n14441) );
  OAI222_X1 U17995 ( .A1(n20262), .A2(n15113), .B1(n20380), .B2(n14586), .C1(
        n14441), .C2(n15116), .ZN(P1_U2895) );
  XNOR2_X1 U17996 ( .A(n14442), .B(n14443), .ZN(n16661) );
  AND2_X1 U17997 ( .A1(n14445), .A2(n14444), .ZN(n14446) );
  OAI22_X1 U17998 ( .A1(n14449), .A2(n14448), .B1(n14447), .B2(n14446), .ZN(
        n16660) );
  INV_X1 U17999 ( .A(n16660), .ZN(n14468) );
  OAI21_X1 U18000 ( .B1(n14452), .B2(n14451), .A(n14450), .ZN(n19470) );
  NOR3_X1 U18001 ( .A1(n14759), .A2(n14454), .A3(n14453), .ZN(n16082) );
  OAI211_X1 U18002 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n16082), .B(n14596), .ZN(n14466) );
  NAND2_X1 U18003 ( .A1(n14456), .A2(n14455), .ZN(n14459) );
  INV_X1 U18004 ( .A(n14457), .ZN(n14458) );
  AND2_X1 U18005 ( .A1(n14459), .A2(n14458), .ZN(n19442) );
  INV_X1 U18006 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n14463) );
  OAI21_X1 U18007 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15968), .A(
        n14460), .ZN(n16081) );
  INV_X1 U18008 ( .A(n16081), .ZN(n14461) );
  OAI22_X1 U18009 ( .A1(n19395), .A2(n14463), .B1(n14462), .B2(n14461), .ZN(
        n14464) );
  AOI21_X1 U18010 ( .B1(n16699), .B2(n19442), .A(n14464), .ZN(n14465) );
  OAI211_X1 U18011 ( .C1(n19470), .C2(n16072), .A(n14466), .B(n14465), .ZN(
        n14467) );
  AOI21_X1 U18012 ( .B1(n14468), .B2(n16700), .A(n14467), .ZN(n14469) );
  OAI21_X1 U18013 ( .B1(n16704), .B2(n16661), .A(n14469), .ZN(P2_U3041) );
  AOI21_X1 U18014 ( .B1(n14471), .B2(n14420), .A(n12875), .ZN(n16574) );
  NAND2_X1 U18015 ( .A1(n16574), .A2(n14786), .ZN(n14475) );
  AOI21_X1 U18016 ( .B1(n14473), .B2(n14472), .A(n14646), .ZN(n19296) );
  NAND2_X1 U18017 ( .A1(n19296), .A2(n15616), .ZN(n14474) );
  OAI211_X1 U18018 ( .C1(n14791), .C2(n19293), .A(n14475), .B(n14474), .ZN(
        P2_U2870) );
  XOR2_X1 U18019 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n14477), .Z(
        n14478) );
  XNOR2_X1 U18020 ( .A(n14476), .B(n14478), .ZN(n16427) );
  INV_X1 U18021 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n14479) );
  OAI22_X1 U18022 ( .A1(n15254), .A2(n14480), .B1(n20432), .B2(n14479), .ZN(
        n14481) );
  AOI21_X1 U18023 ( .B1(n16355), .B2(n14482), .A(n14481), .ZN(n14485) );
  NAND2_X1 U18024 ( .A1(n14483), .A2(n16364), .ZN(n14484) );
  OAI211_X1 U18025 ( .C1(n16427), .C2(n20238), .A(n14485), .B(n14484), .ZN(
        P1_U2991) );
  OAI21_X1 U18026 ( .B1(n14486), .B2(n14487), .A(n14488), .ZN(n14548) );
  OAI21_X1 U18027 ( .B1(n14548), .B2(n14549), .A(n14488), .ZN(n14490) );
  NAND2_X1 U18028 ( .A1(n14490), .A2(n14489), .ZN(n14527) );
  OAI21_X1 U18029 ( .B1(n14490), .B2(n14489), .A(n14527), .ZN(n15272) );
  INV_X1 U18030 ( .A(DATAI_12_), .ZN(n21071) );
  MUX2_X1 U18031 ( .A(n21071), .B(n16783), .S(n14699), .Z(n20390) );
  OAI222_X1 U18032 ( .A1(n15272), .A2(n15113), .B1(n20390), .B2(n14586), .C1(
        n14491), .C2(n15116), .ZN(P1_U2892) );
  INV_X1 U18033 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n14494) );
  OAI21_X1 U18034 ( .B1(n14492), .B2(n14493), .A(n14535), .ZN(n16333) );
  OAI222_X1 U18035 ( .A1(n15272), .A2(n15040), .B1(n14494), .B2(n15047), .C1(
        n16333), .C2(n15048), .ZN(P1_U2860) );
  INV_X1 U18036 ( .A(n20579), .ZN(n14495) );
  NAND2_X1 U18037 ( .A1(n20838), .A2(n14543), .ZN(n14496) );
  AOI21_X1 U18038 ( .B1(n14496), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20880), 
        .ZN(n14504) );
  NOR2_X1 U18039 ( .A1(n20840), .A2(n20841), .ZN(n14501) );
  INV_X1 U18040 ( .A(n14497), .ZN(n14498) );
  AND2_X1 U18041 ( .A1(n14498), .A2(n20769), .ZN(n20706) );
  INV_X1 U18042 ( .A(n20925), .ZN(n20868) );
  NOR2_X1 U18043 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14499), .ZN(
        n14541) );
  INV_X1 U18044 ( .A(n14501), .ZN(n14503) );
  NOR2_X1 U18045 ( .A1(n20706), .A2(n12006), .ZN(n14502) );
  AOI21_X1 U18046 ( .B1(n14504), .B2(n14503), .A(n14502), .ZN(n14505) );
  OAI211_X1 U18047 ( .C1(n14541), .C2(n20774), .A(n20847), .B(n14505), .ZN(
        n14540) );
  AOI22_X1 U18048 ( .A1(n20924), .A2(n14541), .B1(
        P1_INSTQUEUE_REG_12__6__SCAN_IN), .B2(n14540), .ZN(n14506) );
  OAI21_X1 U18049 ( .B1(n14543), .B2(n20868), .A(n14506), .ZN(n14507) );
  AOI21_X1 U18050 ( .B1(n14545), .B2(n20865), .A(n14507), .ZN(n14508) );
  OAI21_X1 U18051 ( .B1(n14547), .B2(n20797), .A(n14508), .ZN(P1_U3135) );
  INV_X1 U18052 ( .A(n20784), .ZN(n20904) );
  AOI22_X1 U18053 ( .A1(n20900), .A2(n14541), .B1(
        P1_INSTQUEUE_REG_12__2__SCAN_IN), .B2(n14540), .ZN(n14509) );
  OAI21_X1 U18054 ( .B1(n14543), .B2(n20904), .A(n14509), .ZN(n14510) );
  AOI21_X1 U18055 ( .B1(n14545), .B2(n20901), .A(n14510), .ZN(n14511) );
  OAI21_X1 U18056 ( .B1(n14547), .B2(n9679), .A(n14511), .ZN(P1_U3131) );
  INV_X1 U18057 ( .A(n20799), .ZN(n20941) );
  AOI22_X1 U18058 ( .A1(n20934), .A2(n14541), .B1(
        P1_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n14540), .ZN(n14512) );
  OAI21_X1 U18059 ( .B1(n14543), .B2(n20941), .A(n14512), .ZN(n14513) );
  AOI21_X1 U18060 ( .B1(n14545), .B2(n20935), .A(n14513), .ZN(n14514) );
  OAI21_X1 U18061 ( .B1(n14547), .B2(n9681), .A(n14514), .ZN(P1_U3136) );
  INV_X1 U18062 ( .A(n20787), .ZN(n20910) );
  AOI22_X1 U18063 ( .A1(n20906), .A2(n14541), .B1(
        P1_INSTQUEUE_REG_12__3__SCAN_IN), .B2(n14540), .ZN(n14515) );
  OAI21_X1 U18064 ( .B1(n14543), .B2(n20910), .A(n14515), .ZN(n14516) );
  AOI21_X1 U18065 ( .B1(n14545), .B2(n20907), .A(n14516), .ZN(n14517) );
  OAI21_X1 U18066 ( .B1(n14547), .B2(n9676), .A(n14517), .ZN(P1_U3132) );
  INV_X1 U18067 ( .A(n20792), .ZN(n20922) );
  AOI22_X1 U18068 ( .A1(n20918), .A2(n14541), .B1(
        P1_INSTQUEUE_REG_12__5__SCAN_IN), .B2(n14540), .ZN(n14518) );
  OAI21_X1 U18069 ( .B1(n14543), .B2(n20922), .A(n14518), .ZN(n14519) );
  AOI21_X1 U18070 ( .B1(n14545), .B2(n20919), .A(n14519), .ZN(n14520) );
  OAI21_X1 U18071 ( .B1(n14547), .B2(n9682), .A(n14520), .ZN(P1_U3134) );
  INV_X1 U18072 ( .A(n20781), .ZN(n20898) );
  AOI22_X1 U18073 ( .A1(n20894), .A2(n14541), .B1(
        P1_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n14540), .ZN(n14521) );
  OAI21_X1 U18074 ( .B1(n14543), .B2(n20898), .A(n14521), .ZN(n14522) );
  AOI21_X1 U18075 ( .B1(n14545), .B2(n20895), .A(n14522), .ZN(n14523) );
  OAI21_X1 U18076 ( .B1(n14547), .B2(n9678), .A(n14523), .ZN(P1_U3130) );
  INV_X1 U18077 ( .A(n14524), .ZN(n14526) );
  AOI21_X1 U18078 ( .B1(n14527), .B2(n14526), .A(n14525), .ZN(n15267) );
  INV_X1 U18079 ( .A(n15267), .ZN(n16325) );
  INV_X1 U18080 ( .A(DATAI_13_), .ZN(n14529) );
  INV_X1 U18081 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14528) );
  MUX2_X1 U18082 ( .A(n14529), .B(n14528), .S(n14699), .Z(n20393) );
  OAI222_X1 U18083 ( .A1(n16325), .A2(n15113), .B1(n20393), .B2(n14586), .C1(
        n14530), .C2(n15116), .ZN(P1_U2891) );
  INV_X1 U18084 ( .A(n20913), .ZN(n20862) );
  AOI22_X1 U18085 ( .A1(n20912), .A2(n14541), .B1(
        P1_INSTQUEUE_REG_12__4__SCAN_IN), .B2(n14540), .ZN(n14531) );
  OAI21_X1 U18086 ( .B1(n20862), .B2(n14543), .A(n14531), .ZN(n14532) );
  AOI21_X1 U18087 ( .B1(n14545), .B2(n20859), .A(n14532), .ZN(n14533) );
  OAI21_X1 U18088 ( .B1(n14547), .B2(n9677), .A(n14533), .ZN(P1_U3133) );
  AND2_X1 U18089 ( .A1(n14535), .A2(n14534), .ZN(n14536) );
  OR2_X1 U18090 ( .A1(n9789), .A2(n14536), .ZN(n16320) );
  OAI22_X1 U18091 ( .A1(n16320), .A2(n15048), .B1(n14537), .B2(n15047), .ZN(
        n14538) );
  AOI21_X1 U18092 ( .B1(n15267), .B2(n15050), .A(n14538), .ZN(n14539) );
  INV_X1 U18093 ( .A(n14539), .ZN(P1_U2859) );
  INV_X1 U18094 ( .A(n20889), .ZN(n20852) );
  AOI22_X1 U18095 ( .A1(n20883), .A2(n14541), .B1(
        P1_INSTQUEUE_REG_12__0__SCAN_IN), .B2(n14540), .ZN(n14542) );
  OAI21_X1 U18096 ( .B1(n20852), .B2(n14543), .A(n14542), .ZN(n14544) );
  AOI21_X1 U18097 ( .B1(n14545), .B2(n20849), .A(n14544), .ZN(n14546) );
  OAI21_X1 U18098 ( .B1(n14547), .B2(n9680), .A(n14546), .ZN(P1_U3129) );
  XOR2_X1 U18099 ( .A(n14549), .B(n14548), .Z(n16363) );
  INV_X1 U18100 ( .A(n16363), .ZN(n14554) );
  INV_X1 U18101 ( .A(n14551), .ZN(n14560) );
  AOI21_X1 U18102 ( .B1(n9881), .B2(n14560), .A(n14492), .ZN(n16396) );
  AOI22_X1 U18103 ( .A1(n16396), .A2(n15038), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n15037), .ZN(n14552) );
  OAI21_X1 U18104 ( .B1(n14554), .B2(n15040), .A(n14552), .ZN(P1_U2861) );
  INV_X1 U18105 ( .A(DATAI_11_), .ZN(n21129) );
  INV_X1 U18106 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n16785) );
  MUX2_X1 U18107 ( .A(n21129), .B(n16785), .S(n14699), .Z(n20387) );
  INV_X1 U18108 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14553) );
  OAI222_X1 U18109 ( .A1(n14554), .A2(n15113), .B1(n20387), .B2(n14586), .C1(
        n14553), .C2(n15116), .ZN(P1_U2893) );
  AOI21_X1 U18110 ( .B1(n14556), .B2(n14555), .A(n14486), .ZN(n15282) );
  NAND2_X1 U18111 ( .A1(n14558), .A2(n14557), .ZN(n14559) );
  NAND2_X1 U18112 ( .A1(n14560), .A2(n14559), .ZN(n16409) );
  OAI22_X1 U18113 ( .A1(n16409), .A2(n15048), .B1(n14561), .B2(n15047), .ZN(
        n14562) );
  AOI21_X1 U18114 ( .B1(n15282), .B2(n15050), .A(n14562), .ZN(n14563) );
  INV_X1 U18115 ( .A(n14563), .ZN(P1_U2862) );
  INV_X1 U18116 ( .A(n15282), .ZN(n14582) );
  INV_X1 U18117 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n16414) );
  NOR3_X1 U18118 ( .A1(n16414), .A2(n20256), .A3(n20255), .ZN(n14569) );
  INV_X1 U18119 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20972) );
  INV_X1 U18120 ( .A(n14971), .ZN(n14564) );
  OAI21_X1 U18121 ( .B1(n14564), .B2(n14972), .A(n20334), .ZN(n16345) );
  AOI21_X1 U18122 ( .B1(n20323), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20310), .ZN(n14567) );
  INV_X1 U18123 ( .A(n15280), .ZN(n14565) );
  AOI22_X1 U18124 ( .A1(n20321), .A2(P1_EBX_REG_10__SCAN_IN), .B1(n14565), 
        .B2(n20338), .ZN(n14566) );
  OAI211_X1 U18125 ( .C1(n20351), .C2(n16409), .A(n14567), .B(n14566), .ZN(
        n14568) );
  AOI221_X1 U18126 ( .B1(n14569), .B2(n20972), .C1(n16345), .C2(
        P1_REIP_REG_10__SCAN_IN), .A(n14568), .ZN(n14570) );
  OAI21_X1 U18127 ( .B1(n14582), .B2(n16324), .A(n14570), .ZN(P1_U2830) );
  INV_X1 U18128 ( .A(n14571), .ZN(n14574) );
  INV_X1 U18129 ( .A(n14525), .ZN(n14573) );
  AOI21_X1 U18130 ( .B1(n14574), .B2(n14573), .A(n14572), .ZN(n16356) );
  INV_X1 U18131 ( .A(n16356), .ZN(n14578) );
  INV_X1 U18132 ( .A(DATAI_14_), .ZN(n21217) );
  INV_X1 U18133 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n16780) );
  MUX2_X1 U18134 ( .A(n21217), .B(n16780), .S(n14699), .Z(n20396) );
  INV_X1 U18135 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14575) );
  OAI222_X1 U18136 ( .A1(n14578), .A2(n15113), .B1(n20396), .B2(n14586), .C1(
        n14575), .C2(n15116), .ZN(P1_U2890) );
  INV_X1 U18137 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14577) );
  OAI21_X1 U18138 ( .B1(n9789), .B2(n14576), .A(n14589), .ZN(n15452) );
  OAI222_X1 U18139 ( .A1(n14578), .A2(n15040), .B1(n14577), .B2(n15047), .C1(
        n15452), .C2(n15048), .ZN(P1_U2858) );
  INV_X1 U18140 ( .A(DATAI_10_), .ZN(n14580) );
  INV_X1 U18141 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n14579) );
  MUX2_X1 U18142 ( .A(n14580), .B(n14579), .S(n14699), .Z(n20384) );
  INV_X1 U18143 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14581) );
  OAI222_X1 U18144 ( .A1(n14582), .A2(n15113), .B1(n20384), .B2(n14586), .C1(
        n14581), .C2(n15116), .ZN(P1_U2894) );
  OAI21_X1 U18145 ( .B1(n14572), .B2(n14584), .A(n14583), .ZN(n16303) );
  OAI222_X1 U18146 ( .A1(n16303), .A2(n15113), .B1(n14586), .B2(n14585), .C1(
        n15116), .C2(n13665), .ZN(P1_U2889) );
  NAND2_X1 U18147 ( .A1(n14589), .A2(n14588), .ZN(n14590) );
  NAND2_X1 U18148 ( .A1(n15044), .A2(n14590), .ZN(n16299) );
  INV_X1 U18149 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14591) );
  OAI222_X1 U18150 ( .A1(n16299), .A2(n15048), .B1(n14591), .B2(n15047), .C1(
        n16303), .C2(n15040), .ZN(P1_U2857) );
  XNOR2_X1 U18151 ( .A(n15830), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n14616) );
  INV_X1 U18152 ( .A(n14593), .ZN(n14594) );
  XNOR2_X1 U18153 ( .A(n14592), .B(n14594), .ZN(n14614) );
  INV_X1 U18154 ( .A(n16082), .ZN(n14595) );
  NOR3_X1 U18155 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n14596), .A3(
        n14595), .ZN(n14608) );
  INV_X1 U18156 ( .A(n16070), .ZN(n14597) );
  AOI21_X1 U18157 ( .B1(n14598), .B2(n14597), .A(n16081), .ZN(n16724) );
  NAND2_X1 U18158 ( .A1(n14599), .A2(n16710), .ZN(n14605) );
  OR2_X1 U18159 ( .A1(n14600), .A2(n14457), .ZN(n14601) );
  NAND2_X1 U18160 ( .A1(n14601), .A2(n13830), .ZN(n19423) );
  INV_X1 U18161 ( .A(n19423), .ZN(n14603) );
  NOR2_X1 U18162 ( .A1(n20109), .A2(n19395), .ZN(n14602) );
  AOI21_X1 U18163 ( .B1(n16699), .B2(n14603), .A(n14602), .ZN(n14604) );
  OAI211_X1 U18164 ( .C1(n16724), .C2(n14606), .A(n14605), .B(n14604), .ZN(
        n14607) );
  OR2_X1 U18165 ( .A1(n14608), .A2(n14607), .ZN(n14609) );
  AOI21_X1 U18166 ( .B1(n14614), .B2(n16721), .A(n14609), .ZN(n14610) );
  OAI21_X1 U18167 ( .B1(n14616), .B2(n16717), .A(n14610), .ZN(P2_U3040) );
  OAI22_X1 U18168 ( .A1(n20109), .A2(n19395), .B1(n19510), .B2(n19421), .ZN(
        n14613) );
  INV_X1 U18169 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n14611) );
  OAI22_X1 U18170 ( .A1(n16655), .A2(n19423), .B1(n16677), .B2(n14611), .ZN(
        n14612) );
  AOI211_X1 U18171 ( .C1(n14614), .C2(n10923), .A(n14613), .B(n14612), .ZN(
        n14615) );
  OAI21_X1 U18172 ( .B1(n14616), .B2(n16668), .A(n14615), .ZN(P2_U3008) );
  MUX2_X1 U18173 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n16420), .S(n9673), .Z(n14618) );
  XNOR2_X1 U18174 ( .A(n14617), .B(n14618), .ZN(n16418) );
  AOI22_X1 U18175 ( .A1(n20416), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(
        n20473), .B2(P1_REIP_REG_9__SCAN_IN), .ZN(n14620) );
  NAND2_X1 U18176 ( .A1(n16355), .A2(n20258), .ZN(n14619) );
  OAI211_X1 U18177 ( .C1(n20262), .C2(n15258), .A(n14620), .B(n14619), .ZN(
        n14621) );
  AOI21_X1 U18178 ( .B1(n16418), .B2(n20422), .A(n14621), .ZN(n14622) );
  INV_X1 U18179 ( .A(n14622), .ZN(P1_U2990) );
  NAND2_X1 U18180 ( .A1(n14470), .A2(n14624), .ZN(n14625) );
  NAND2_X1 U18181 ( .A1(n14623), .A2(n14625), .ZN(n14649) );
  INV_X1 U18182 ( .A(n14626), .ZN(n14635) );
  NAND2_X1 U18183 ( .A1(n14628), .A2(n14627), .ZN(n14629) );
  NAND2_X1 U18184 ( .A1(n14635), .A2(n14629), .ZN(n15957) );
  INV_X1 U18185 ( .A(n15957), .ZN(n19284) );
  OAI22_X1 U18186 ( .A1(n19540), .A2(n15690), .B1(n15689), .B2(n13485), .ZN(
        n14632) );
  INV_X1 U18187 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n14630) );
  OAI22_X1 U18188 ( .A1(n15693), .A2(n16772), .B1(n15692), .B2(n14630), .ZN(
        n14631) );
  AOI211_X1 U18189 ( .C1(n19284), .C2(n19449), .A(n14632), .B(n14631), .ZN(
        n14633) );
  OAI21_X1 U18190 ( .B1(n19465), .B2(n14649), .A(n14633), .ZN(P2_U2901) );
  AND2_X1 U18191 ( .A1(n14635), .A2(n14634), .ZN(n14637) );
  OR2_X1 U18192 ( .A1(n14637), .A2(n14636), .ZN(n19273) );
  NOR2_X1 U18193 ( .A1(n15692), .A2(n18527), .ZN(n14640) );
  OAI22_X1 U18194 ( .A1(n19544), .A2(n15690), .B1(n15689), .B2(n14638), .ZN(
        n14639) );
  AOI211_X1 U18195 ( .C1(BUF1_REG_19__SCAN_IN), .C2(n19451), .A(n14640), .B(
        n14639), .ZN(n14644) );
  AOI21_X1 U18196 ( .B1(n14642), .B2(n14623), .A(n14641), .ZN(n14650) );
  NAND2_X1 U18197 ( .A1(n14650), .A2(n13177), .ZN(n14643) );
  OAI211_X1 U18198 ( .C1(n19273), .C2(n15675), .A(n14644), .B(n14643), .ZN(
        P2_U2900) );
  OAI21_X1 U18199 ( .B1(n14646), .B2(n14645), .A(n9774), .ZN(n19282) );
  NOR2_X1 U18200 ( .A1(n19282), .A2(n13835), .ZN(n14647) );
  AOI21_X1 U18201 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n13835), .A(n14647), .ZN(
        n14648) );
  OAI21_X1 U18202 ( .B1(n14649), .B2(n15618), .A(n14648), .ZN(P2_U2869) );
  NAND2_X1 U18203 ( .A1(n14650), .A2(n14786), .ZN(n14654) );
  NAND2_X1 U18204 ( .A1(n9774), .A2(n14651), .ZN(n14652) );
  NAND2_X1 U18205 ( .A1(n9748), .A2(n14652), .ZN(n15940) );
  INV_X1 U18206 ( .A(n15940), .ZN(n19269) );
  NAND2_X1 U18207 ( .A1(n19269), .A2(n15616), .ZN(n14653) );
  OAI211_X1 U18208 ( .C1(n15616), .C2(n10719), .A(n14654), .B(n14653), .ZN(
        P2_U2868) );
  AOI21_X1 U18209 ( .B1(n18984), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14663) );
  OR2_X1 U18210 ( .A1(n14657), .A2(n14663), .ZN(n18974) );
  NOR2_X1 U18211 ( .A1(n19150), .A2(n18974), .ZN(n14662) );
  OR2_X1 U18212 ( .A1(n9725), .A2(n17765), .ZN(n19028) );
  AOI21_X1 U18213 ( .B1(n14655), .B2(n19028), .A(n19184), .ZN(n14656) );
  NAND2_X1 U18214 ( .A1(n18970), .A2(n19187), .ZN(n14660) );
  AOI221_X2 U18215 ( .B1(n19186), .B2(n14657), .C1(n17765), .C2(n14657), .A(
        n14660), .ZN(n16277) );
  AOI21_X1 U18216 ( .B1(n16093), .B2(n18967), .A(n16277), .ZN(n14658) );
  OAI211_X1 U18217 ( .C1(n17726), .C2(n14660), .A(n14659), .B(n14658), .ZN(
        n19001) );
  NOR2_X1 U18218 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n19138), .ZN(n18516) );
  INV_X1 U18219 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18506) );
  NOR3_X1 U18220 ( .A1(n19147), .A2(n19039), .A3(n19029), .ZN(n19046) );
  INV_X1 U18221 ( .A(n19046), .ZN(n19136) );
  NOR2_X1 U18222 ( .A1(n18506), .A2(n19136), .ZN(n14661) );
  MUX2_X1 U18223 ( .A(n14662), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19166), .Z(P3_U3284) );
  NAND2_X1 U18224 ( .A1(n14663), .A2(n17474), .ZN(n18505) );
  NOR2_X1 U18225 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18505), .ZN(n14664) );
  OAI21_X1 U18226 ( .B1(n14664), .B2(n19136), .A(n18667), .ZN(n18511) );
  INV_X1 U18227 ( .A(n18511), .ZN(n14665) );
  NOR2_X1 U18228 ( .A1(n19179), .A2(n17976), .ZN(n16190) );
  AOI21_X1 U18229 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n16190), .ZN(n16191) );
  NOR2_X1 U18230 ( .A1(n14665), .A2(n16191), .ZN(n14667) );
  INV_X1 U18231 ( .A(n18876), .ZN(n18773) );
  NOR2_X1 U18232 ( .A1(n19138), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18552) );
  INV_X1 U18233 ( .A(n18552), .ZN(n18692) );
  NAND2_X1 U18234 ( .A1(n18692), .A2(n18511), .ZN(n16189) );
  OR2_X1 U18235 ( .A1(n18773), .A2(n16189), .ZN(n14666) );
  MUX2_X1 U18236 ( .A(n14667), .B(n14666), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  AOI21_X1 U18237 ( .B1(n14670), .B2(n15522), .A(n15524), .ZN(n19245) );
  NAND2_X1 U18238 ( .A1(n16667), .A2(n19245), .ZN(n14669) );
  OAI211_X1 U18239 ( .C1(n16677), .C2(n14670), .A(n14669), .B(n14668), .ZN(
        n14673) );
  NOR3_X1 U18240 ( .A1(n14671), .A2(n13229), .A3(n16668), .ZN(n14672) );
  AOI211_X1 U18241 ( .C1(n19504), .C2(n19240), .A(n14673), .B(n14672), .ZN(
        n14674) );
  OAI21_X1 U18242 ( .B1(n14675), .B2(n16671), .A(n14674), .ZN(P2_U2993) );
  AOI21_X1 U18243 ( .B1(n19501), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14676), .ZN(n14681) );
  XNOR2_X1 U18244 ( .A(n14678), .B(n14677), .ZN(n16485) );
  INV_X1 U18245 ( .A(n16485), .ZN(n14679) );
  NAND2_X1 U18246 ( .A1(n16667), .A2(n14679), .ZN(n14680) );
  OAI211_X1 U18247 ( .C1(n16481), .C2(n16655), .A(n14681), .B(n14680), .ZN(
        n14682) );
  AOI21_X1 U18248 ( .B1(n14683), .B2(n19505), .A(n14682), .ZN(n14684) );
  OAI21_X1 U18249 ( .B1(n14685), .B2(n16671), .A(n14684), .ZN(P2_U2984) );
  NOR2_X1 U18250 ( .A1(n14871), .A2(n14687), .ZN(n14688) );
  OR2_X1 U18251 ( .A1(n14689), .A2(n14688), .ZN(n14703) );
  INV_X1 U18252 ( .A(n14703), .ZN(n15299) );
  NOR3_X1 U18253 ( .A1(n14972), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n14690), 
        .ZN(n14691) );
  AOI21_X1 U18254 ( .B1(P1_EBX_REG_29__SCAN_IN), .B2(n20321), .A(n14691), .ZN(
        n14694) );
  AOI22_X1 U18255 ( .A1(n20338), .A2(n14692), .B1(
        P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20323), .ZN(n14693) );
  OAI211_X1 U18256 ( .C1(n14878), .C2(n21096), .A(n14694), .B(n14693), .ZN(
        n14695) );
  AOI21_X1 U18257 ( .B1(n15299), .B2(n20320), .A(n14695), .ZN(n14696) );
  OAI21_X1 U18258 ( .B1(n14686), .B2(n16324), .A(n14696), .ZN(P1_U2811) );
  INV_X1 U18259 ( .A(n14700), .ZN(n14697) );
  NAND2_X1 U18260 ( .A1(n14697), .A2(n14699), .ZN(n15084) );
  OAI22_X1 U18261 ( .A1(n15118), .A2(n20393), .B1(n13592), .B2(n15116), .ZN(
        n14698) );
  AOI21_X1 U18262 ( .B1(n15120), .B2(BUF1_REG_29__SCAN_IN), .A(n14698), .ZN(
        n14702) );
  NOR2_X2 U18263 ( .A1(n14700), .A2(n14699), .ZN(n15110) );
  NAND2_X1 U18264 ( .A1(n15110), .A2(DATAI_29_), .ZN(n14701) );
  OAI211_X1 U18265 ( .C1(n14686), .C2(n15113), .A(n14702), .B(n14701), .ZN(
        P1_U2875) );
  OAI222_X1 U18266 ( .A1(n15040), .A2(n14686), .B1(n14704), .B2(n15047), .C1(
        n14703), .C2(n15048), .ZN(P1_U2843) );
  NAND2_X1 U18267 ( .A1(n15449), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14705) );
  NOR2_X1 U18268 ( .A1(n9674), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14706) );
  XNOR2_X1 U18269 ( .A(n14710), .B(n14709), .ZN(n14740) );
  NOR2_X1 U18270 ( .A1(n15016), .A2(n20469), .ZN(n14733) );
  INV_X1 U18271 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15296) );
  INV_X1 U18272 ( .A(n15132), .ZN(n15323) );
  NAND4_X1 U18273 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15416) );
  NOR2_X1 U18274 ( .A1(n15416), .A2(n15419), .ZN(n14729) );
  AND2_X1 U18275 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14729), .ZN(
        n15366) );
  INV_X1 U18276 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16434) );
  INV_X1 U18277 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16426) );
  NOR3_X1 U18278 ( .A1(n16434), .A2(n16439), .A3(n16426), .ZN(n16402) );
  NAND3_X1 U18279 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16402), .ZN(n15475) );
  NOR2_X1 U18280 ( .A1(n16395), .A2(n15475), .ZN(n15485) );
  AND2_X1 U18281 ( .A1(n15485), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14714) );
  INV_X1 U18282 ( .A(n14714), .ZN(n14712) );
  NAND2_X1 U18283 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16423) );
  NAND2_X1 U18284 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20456) );
  NOR2_X1 U18285 ( .A1(n16423), .A2(n20456), .ZN(n14711) );
  AND2_X1 U18286 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14711), .ZN(
        n16403) );
  INV_X1 U18287 ( .A(n16403), .ZN(n15476) );
  NOR2_X1 U18288 ( .A1(n14712), .A2(n15476), .ZN(n15465) );
  AOI21_X1 U18289 ( .B1(n15366), .B2(n15465), .A(n16404), .ZN(n14716) );
  INV_X1 U18290 ( .A(n16423), .ZN(n20430) );
  OAI21_X1 U18291 ( .B1(n20455), .B2(n20451), .A(n20464), .ZN(n20454) );
  NAND3_X1 U18292 ( .A1(n20430), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        n20454), .ZN(n15477) );
  INV_X1 U18293 ( .A(n15477), .ZN(n14713) );
  AND2_X1 U18294 ( .A1(n14714), .A2(n14713), .ZN(n15457) );
  AOI21_X1 U18295 ( .B1(n15366), .B2(n15457), .A(n20428), .ZN(n14715) );
  NOR3_X1 U18296 ( .A1(n14716), .A2(n14715), .A3(n20449), .ZN(n15402) );
  NOR2_X1 U18297 ( .A1(n15401), .A2(n15368), .ZN(n15388) );
  INV_X1 U18298 ( .A(n20449), .ZN(n14717) );
  AOI22_X1 U18299 ( .A1(n15402), .A2(n15388), .B1(n14718), .B2(n14717), .ZN(
        n15382) );
  AOI21_X1 U18300 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(n14718), .ZN(n14719) );
  OR2_X1 U18301 ( .A1(n15382), .A2(n14719), .ZN(n15354) );
  AOI21_X1 U18302 ( .B1(n20467), .B2(n15343), .A(n15354), .ZN(n15345) );
  INV_X1 U18303 ( .A(n15325), .ZN(n14720) );
  AOI22_X1 U18304 ( .A1(n20467), .A2(n15346), .B1(n20466), .B2(n14720), .ZN(
        n14721) );
  OAI211_X1 U18305 ( .C1(n15323), .C2(n20475), .A(n15345), .B(n14721), .ZN(
        n15337) );
  INV_X1 U18306 ( .A(n15293), .ZN(n15303) );
  NAND2_X1 U18307 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15302) );
  NOR3_X1 U18308 ( .A1(n15337), .A2(n15303), .A3(n15302), .ZN(n14722) );
  NOR2_X1 U18309 ( .A1(n15337), .A2(n16425), .ZN(n14723) );
  NOR2_X1 U18310 ( .A1(n14722), .A2(n14723), .ZN(n15292) );
  AOI211_X1 U18311 ( .C1(n15296), .C2(n16425), .A(n15288), .B(n15292), .ZN(
        n15286) );
  NOR3_X1 U18312 ( .A1(n15286), .A2(n14723), .A3(n14709), .ZN(n14732) );
  INV_X1 U18313 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n21185) );
  NOR2_X1 U18314 ( .A1(n20432), .A2(n21185), .ZN(n14735) );
  INV_X1 U18315 ( .A(n15457), .ZN(n14724) );
  OR2_X1 U18316 ( .A1(n20428), .A2(n14724), .ZN(n15363) );
  NAND2_X1 U18317 ( .A1(n15465), .A2(n15479), .ZN(n14726) );
  NAND2_X1 U18318 ( .A1(n15363), .A2(n14726), .ZN(n14727) );
  NAND2_X1 U18319 ( .A1(n14727), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15424) );
  INV_X1 U18320 ( .A(n14728), .ZN(n15371) );
  NAND3_X1 U18321 ( .A1(n14729), .A2(n15371), .A3(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14730) );
  NOR3_X1 U18322 ( .A1(n15357), .A2(n15132), .A3(n15322), .ZN(n15317) );
  NAND3_X1 U18323 ( .A1(n15317), .A2(n15293), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15287) );
  NOR3_X1 U18324 ( .A1(n15287), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15288), .ZN(n14731) );
  OAI21_X1 U18325 ( .B1(n14740), .B2(n20470), .A(n14734), .ZN(P1_U3000) );
  AOI21_X1 U18326 ( .B1(n20416), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14735), .ZN(n14736) );
  OAI21_X1 U18327 ( .B1(n14737), .B2(n20427), .A(n14736), .ZN(n14738) );
  AOI21_X1 U18328 ( .B1(n15054), .B2(n16364), .A(n14738), .ZN(n14739) );
  OAI21_X1 U18329 ( .B1(n14740), .B2(n20238), .A(n14739), .ZN(P1_U2968) );
  XNOR2_X1 U18330 ( .A(n14741), .B(n14773), .ZN(n14742) );
  NAND2_X1 U18331 ( .A1(n14742), .A2(n19443), .ZN(n14751) );
  NOR2_X1 U18332 ( .A1(n14753), .A2(n19447), .ZN(n14748) );
  NOR2_X1 U18333 ( .A1(n19434), .A2(n14743), .ZN(n14747) );
  NOR2_X1 U18334 ( .A1(n19400), .A2(n10287), .ZN(n14746) );
  INV_X1 U18335 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14744) );
  OAI22_X1 U18336 ( .A1(n19417), .A2(n20104), .B1(n19397), .B2(n14744), .ZN(
        n14745) );
  OR4_X1 U18337 ( .A1(n14748), .A2(n14747), .A3(n14746), .A4(n14745), .ZN(
        n14749) );
  AOI21_X1 U18338 ( .B1(n12788), .B2(n19441), .A(n14749), .ZN(n14750) );
  OAI211_X1 U18339 ( .C1(n20178), .C2(n14752), .A(n14751), .B(n14750), .ZN(
        P2_U2853) );
  INV_X1 U18340 ( .A(n14753), .ZN(n20180) );
  AOI21_X1 U18341 ( .B1(n14756), .B2(n14755), .A(n14754), .ZN(n14781) );
  NAND2_X1 U18342 ( .A1(n14781), .A2(n16700), .ZN(n14764) );
  OAI21_X1 U18343 ( .B1(n14759), .B2(n14758), .A(n14757), .ZN(n14763) );
  NAND2_X1 U18344 ( .A1(n19500), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n14775) );
  NAND2_X1 U18345 ( .A1(n14761), .A2(n14760), .ZN(n14777) );
  NAND3_X1 U18346 ( .A1(n16721), .A2(n14778), .A3(n14777), .ZN(n14762) );
  NAND4_X1 U18347 ( .A1(n14764), .A2(n14763), .A3(n14775), .A4(n14762), .ZN(
        n14771) );
  INV_X1 U18348 ( .A(n14765), .ZN(n14766) );
  AOI21_X1 U18349 ( .B1(n15967), .B2(n14768), .A(n14766), .ZN(n14769) );
  OAI22_X1 U18350 ( .A1(n14769), .A2(n10290), .B1(n14768), .B2(n14767), .ZN(
        n14770) );
  AOI211_X1 U18351 ( .C1(n20180), .C2(n16710), .A(n14771), .B(n14770), .ZN(
        n14772) );
  OAI21_X1 U18352 ( .B1(n10352), .B2(n16716), .A(n14772), .ZN(P2_U3044) );
  INV_X1 U18353 ( .A(n14773), .ZN(n14774) );
  NAND2_X1 U18354 ( .A1(n16667), .A2(n14774), .ZN(n14776) );
  OAI211_X1 U18355 ( .C1(n14744), .C2(n16677), .A(n14776), .B(n14775), .ZN(
        n14780) );
  AND3_X1 U18356 ( .A1(n14778), .A2(n10923), .A3(n14777), .ZN(n14779) );
  AOI211_X1 U18357 ( .C1(n14781), .C2(n19505), .A(n14780), .B(n14779), .ZN(
        n14782) );
  OAI21_X1 U18358 ( .B1(n10352), .B2(n16655), .A(n14782), .ZN(P2_U3012) );
  XOR2_X1 U18359 ( .A(n13836), .B(P2_INSTQUEUE_REG_0__6__SCAN_IN), .Z(n14784)
         );
  MUX2_X1 U18360 ( .A(n19412), .B(n19423), .S(n15616), .Z(n14783) );
  OAI21_X1 U18361 ( .B1(n14784), .B2(n15618), .A(n14783), .ZN(P2_U2881) );
  INV_X1 U18362 ( .A(n14785), .ZN(n14787) );
  OAI211_X1 U18363 ( .C1(n14787), .C2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n14786), .B(n13836), .ZN(n14789) );
  NAND2_X1 U18364 ( .A1(n14791), .A2(n19442), .ZN(n14788) );
  OAI211_X1 U18365 ( .C1(n14791), .C2(n14790), .A(n14789), .B(n14788), .ZN(
        P2_U2882) );
  NOR2_X1 U18366 ( .A1(n14792), .A2(n20161), .ZN(n14798) );
  INV_X1 U18367 ( .A(n14793), .ZN(n14794) );
  OAI22_X1 U18368 ( .A1(n14796), .A2(n20165), .B1(n14795), .B2(n14794), .ZN(
        n14797) );
  OAI21_X1 U18369 ( .B1(n14798), .B2(n14797), .A(n20162), .ZN(n14799) );
  OAI21_X1 U18370 ( .B1(n20162), .B2(n10016), .A(n14799), .ZN(P2_U3601) );
  INV_X1 U18371 ( .A(n14800), .ZN(n14801) );
  NOR2_X1 U18372 ( .A1(n14802), .A2(n14801), .ZN(n14805) );
  OAI22_X1 U18373 ( .A1(n19513), .A2(n20161), .B1(n20165), .B2(n14803), .ZN(
        n14804) );
  OAI21_X1 U18374 ( .B1(n14805), .B2(n14804), .A(n20162), .ZN(n14806) );
  OAI21_X1 U18375 ( .B1(n20162), .B2(n14807), .A(n14806), .ZN(P2_U3600) );
  INV_X1 U18376 ( .A(n14808), .ZN(n14812) );
  NOR2_X1 U18377 ( .A1(n14814), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14817) );
  MUX2_X1 U18378 ( .A(n14817), .B(n14816), .S(n14815), .Z(n16471) );
  NAND2_X1 U18379 ( .A1(n16471), .A2(n14818), .ZN(n14819) );
  XNOR2_X1 U18380 ( .A(n14819), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14820) );
  XNOR2_X1 U18381 ( .A(n14821), .B(n14820), .ZN(n15706) );
  AOI222_X1 U18382 ( .A1(n14824), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n9735), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n14823), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n14825) );
  INV_X1 U18383 ( .A(n14825), .ZN(n14826) );
  INV_X1 U18384 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n20150) );
  NOR2_X1 U18385 ( .A1(n19395), .A2(n20150), .ZN(n15700) );
  NOR2_X1 U18386 ( .A1(n15968), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14828) );
  OAI21_X1 U18387 ( .B1(n14829), .B2(n14828), .A(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14831) );
  AND2_X1 U18388 ( .A1(n14831), .A2(n10106), .ZN(n14832) );
  AOI22_X1 U18389 ( .A1(n11340), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14837) );
  NAND2_X1 U18390 ( .A1(n9658), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14836) );
  OAI211_X1 U18391 ( .C1(n10662), .C2(n14838), .A(n14837), .B(n14836), .ZN(
        n14839) );
  XNOR2_X1 U18392 ( .A(n14840), .B(n14839), .ZN(n15702) );
  OAI21_X1 U18393 ( .B1(n15706), .B2(n16704), .A(n14844), .ZN(P2_U3015) );
  INV_X1 U18394 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n14845) );
  NAND2_X1 U18395 ( .A1(n14846), .A2(n14845), .ZN(n14848) );
  MUX2_X1 U18396 ( .A(n14848), .B(n14847), .S(n21025), .Z(P1_U3487) );
  MUX2_X1 U18397 ( .A(n14850), .B(n14849), .S(n14851), .Z(n14855) );
  AOI22_X1 U18398 ( .A1(n12572), .A2(n14853), .B1(n14852), .B2(n14851), .ZN(
        n14854) );
  NAND2_X1 U18399 ( .A1(n14855), .A2(n14854), .ZN(n16233) );
  OR3_X1 U18400 ( .A1(n14857), .A2(n9660), .A3(n16265), .ZN(n21020) );
  AND2_X1 U18401 ( .A1(n21020), .A2(n21027), .ZN(n14858) );
  OR2_X1 U18402 ( .A1(n14859), .A2(n14858), .ZN(n16232) );
  AND2_X1 U18403 ( .A1(n16232), .A2(n14860), .ZN(n20239) );
  MUX2_X1 U18404 ( .A(P1_MORE_REG_SCAN_IN), .B(n16233), .S(n20239), .Z(
        P1_U3484) );
  NAND2_X1 U18405 ( .A1(n15129), .A2(n20287), .ZN(n14868) );
  INV_X1 U18406 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14861) );
  OAI22_X1 U18407 ( .A1(n20306), .A2(n15127), .B1(n14861), .B2(n20335), .ZN(
        n14866) );
  INV_X1 U18408 ( .A(n14862), .ZN(n14863) );
  AOI21_X1 U18409 ( .B1(n21108), .B2(n14864), .A(n14863), .ZN(n14865) );
  AOI211_X1 U18410 ( .C1(n20321), .C2(P1_EBX_REG_30__SCAN_IN), .A(n14866), .B(
        n14865), .ZN(n14867) );
  OAI211_X1 U18411 ( .C1(n20351), .C2(n15285), .A(n14868), .B(n14867), .ZN(
        P1_U2810) );
  AOI21_X1 U18412 ( .B1(n14870), .B2(n14869), .A(n13330), .ZN(n15141) );
  INV_X1 U18413 ( .A(n15141), .ZN(n15063) );
  AOI21_X1 U18414 ( .B1(n14872), .B2(n14883), .A(n14871), .ZN(n15308) );
  OAI22_X1 U18415 ( .A1(n20306), .A2(n15139), .B1(n14873), .B2(n20335), .ZN(
        n14876) );
  NOR4_X1 U18416 ( .A1(n14972), .A2(n14874), .A3(n21199), .A4(n14885), .ZN(
        n14875) );
  AOI211_X1 U18417 ( .C1(P1_EBX_REG_28__SCAN_IN), .C2(n20321), .A(n14876), .B(
        n14875), .ZN(n14877) );
  OAI21_X1 U18418 ( .B1(n14878), .B2(n21038), .A(n14877), .ZN(n14879) );
  AOI21_X1 U18419 ( .B1(n15308), .B2(n20320), .A(n14879), .ZN(n14880) );
  OAI21_X1 U18420 ( .B1(n15063), .B2(n16324), .A(n14880), .ZN(P1_U2812) );
  OAI21_X1 U18421 ( .B1(n14881), .B2(n14882), .A(n14869), .ZN(n15151) );
  AOI21_X1 U18422 ( .B1(n14884), .B2(n14891), .A(n9887), .ZN(n15311) );
  AOI21_X1 U18423 ( .B1(n20347), .B2(n14885), .A(n20276), .ZN(n14899) );
  NOR3_X1 U18424 ( .A1(n14972), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14885), 
        .ZN(n14886) );
  AOI21_X1 U18425 ( .B1(P1_EBX_REG_27__SCAN_IN), .B2(n20321), .A(n14886), .ZN(
        n14888) );
  AOI22_X1 U18426 ( .A1(n20338), .A2(n15145), .B1(
        P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20323), .ZN(n14887) );
  OAI211_X1 U18427 ( .C1(n14899), .C2(n21199), .A(n14888), .B(n14887), .ZN(
        n14889) );
  AOI21_X1 U18428 ( .B1(n15311), .B2(n20320), .A(n14889), .ZN(n14890) );
  OAI21_X1 U18429 ( .B1(n15151), .B2(n16324), .A(n14890), .ZN(P1_U2813) );
  OAI21_X1 U18430 ( .B1(n14911), .B2(n14892), .A(n14891), .ZN(n15321) );
  AOI21_X1 U18432 ( .B1(n14895), .B2(n14894), .A(n14881), .ZN(n15158) );
  NAND2_X1 U18433 ( .A1(n15158), .A2(n20287), .ZN(n14903) );
  OAI22_X1 U18434 ( .A1(n20306), .A2(n15156), .B1(n14896), .B2(n20335), .ZN(
        n14901) );
  AOI21_X1 U18435 ( .B1(n20347), .B2(n14897), .A(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14898) );
  NOR2_X1 U18436 ( .A1(n14899), .A2(n14898), .ZN(n14900) );
  AOI211_X1 U18437 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n20321), .A(n14901), .B(
        n14900), .ZN(n14902) );
  OAI211_X1 U18438 ( .C1(n20351), .C2(n15321), .A(n14903), .B(n14902), .ZN(
        P1_U2814) );
  OAI21_X1 U18439 ( .B1(n14905), .B2(n14906), .A(n14894), .ZN(n15166) );
  INV_X1 U18440 ( .A(n14922), .ZN(n14907) );
  OAI21_X1 U18441 ( .B1(n14972), .B2(n14907), .A(n20334), .ZN(n14937) );
  INV_X1 U18442 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15021) );
  OAI21_X1 U18443 ( .B1(n14922), .B2(P1_REIP_REG_25__SCAN_IN), .A(
        P1_REIP_REG_24__SCAN_IN), .ZN(n14908) );
  OAI211_X1 U18444 ( .C1(P1_REIP_REG_24__SCAN_IN), .C2(P1_REIP_REG_25__SCAN_IN), .A(n20347), .B(n14908), .ZN(n14910) );
  AOI22_X1 U18445 ( .A1(n20338), .A2(n15169), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20323), .ZN(n14909) );
  OAI211_X1 U18446 ( .C1(n15021), .C2(n20340), .A(n14910), .B(n14909), .ZN(
        n14915) );
  INV_X1 U18447 ( .A(n14911), .ZN(n14912) );
  OAI21_X1 U18448 ( .B1(n14913), .B2(n14919), .A(n14912), .ZN(n15338) );
  NOR2_X1 U18449 ( .A1(n15338), .A2(n20351), .ZN(n14914) );
  AOI211_X1 U18450 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n14937), .A(n14915), 
        .B(n14914), .ZN(n14916) );
  OAI21_X1 U18451 ( .B1(n15166), .B2(n16324), .A(n14916), .ZN(P1_U2815) );
  AOI21_X1 U18452 ( .B1(n14918), .B2(n14917), .A(n14905), .ZN(n15177) );
  INV_X1 U18453 ( .A(n15177), .ZN(n15023) );
  AOI21_X1 U18454 ( .B1(n14920), .B2(n14933), .A(n14919), .ZN(n15351) );
  INV_X1 U18455 ( .A(n14937), .ZN(n14926) );
  INV_X1 U18456 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n21047) );
  OAI22_X1 U18457 ( .A1(n20306), .A2(n15175), .B1(n14921), .B2(n20335), .ZN(
        n14924) );
  NOR3_X1 U18458 ( .A1(n14972), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n14922), 
        .ZN(n14923) );
  AOI211_X1 U18459 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n20321), .A(n14924), .B(
        n14923), .ZN(n14925) );
  OAI21_X1 U18460 ( .B1(n14926), .B2(n21047), .A(n14925), .ZN(n14927) );
  AOI21_X1 U18461 ( .B1(n15351), .B2(n20320), .A(n14927), .ZN(n14928) );
  OAI21_X1 U18462 ( .B1(n15023), .B2(n16324), .A(n14928), .ZN(P1_U2816) );
  OAI21_X1 U18463 ( .B1(n14929), .B2(n14930), .A(n14917), .ZN(n15181) );
  INV_X1 U18464 ( .A(n14931), .ZN(n14957) );
  AOI21_X1 U18465 ( .B1(n14957), .B2(n14943), .A(n14932), .ZN(n14935) );
  INV_X1 U18466 ( .A(n14933), .ZN(n14934) );
  NOR2_X1 U18467 ( .A1(n14935), .A2(n14934), .ZN(n15359) );
  INV_X1 U18468 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15025) );
  NOR2_X1 U18469 ( .A1(n14972), .A2(n14936), .ZN(n14938) );
  OAI21_X1 U18470 ( .B1(n14938), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14937), 
        .ZN(n14940) );
  AOI22_X1 U18471 ( .A1(n20338), .A2(n15184), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20323), .ZN(n14939) );
  OAI211_X1 U18472 ( .C1(n20340), .C2(n15025), .A(n14940), .B(n14939), .ZN(
        n14941) );
  AOI21_X1 U18473 ( .B1(n15359), .B2(n20320), .A(n14941), .ZN(n14942) );
  OAI21_X1 U18474 ( .B1(n15181), .B2(n16324), .A(n14942), .ZN(P1_U2817) );
  XNOR2_X1 U18475 ( .A(n14957), .B(n14943), .ZN(n15362) );
  AOI21_X1 U18476 ( .B1(n14944), .B2(n9757), .A(n14929), .ZN(n15192) );
  NAND2_X1 U18477 ( .A1(n15192), .A2(n20287), .ZN(n14952) );
  OAI21_X1 U18478 ( .B1(n14972), .B2(n14946), .A(n20334), .ZN(n14983) );
  OAI22_X1 U18479 ( .A1(n20306), .A2(n15190), .B1(n14945), .B2(n20335), .ZN(
        n14950) );
  INV_X1 U18480 ( .A(n14946), .ZN(n14960) );
  OAI21_X1 U18481 ( .B1(n14960), .B2(P1_REIP_REG_22__SCAN_IN), .A(
        P1_REIP_REG_21__SCAN_IN), .ZN(n14947) );
  OAI211_X1 U18482 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(P1_REIP_REG_22__SCAN_IN), .A(n20347), .B(n14947), .ZN(n14948) );
  OAI21_X1 U18483 ( .B1(n15026), .B2(n20340), .A(n14948), .ZN(n14949) );
  AOI211_X1 U18484 ( .C1(n14983), .C2(P1_REIP_REG_22__SCAN_IN), .A(n14950), 
        .B(n14949), .ZN(n14951) );
  OAI211_X1 U18485 ( .C1(n15362), .C2(n20351), .A(n14952), .B(n14951), .ZN(
        P1_U2818) );
  NAND2_X1 U18486 ( .A1(n14969), .A2(n14954), .ZN(n14955) );
  NAND2_X1 U18487 ( .A1(n9757), .A2(n14955), .ZN(n15199) );
  NAND2_X1 U18488 ( .A1(n14993), .A2(n14956), .ZN(n14958) );
  AOI21_X1 U18489 ( .B1(n14959), .B2(n14958), .A(n14957), .ZN(n15383) );
  INV_X1 U18490 ( .A(n14983), .ZN(n14965) );
  INV_X1 U18491 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n14964) );
  NOR3_X1 U18492 ( .A1(n14972), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n14960), 
        .ZN(n14961) );
  AOI21_X1 U18493 ( .B1(P1_EBX_REG_21__SCAN_IN), .B2(n20321), .A(n14961), .ZN(
        n14963) );
  AOI22_X1 U18494 ( .A1(n20338), .A2(n15202), .B1(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20323), .ZN(n14962) );
  OAI211_X1 U18495 ( .C1(n14965), .C2(n14964), .A(n14963), .B(n14962), .ZN(
        n14966) );
  AOI21_X1 U18496 ( .B1(n15383), .B2(n20320), .A(n14966), .ZN(n14967) );
  OAI21_X1 U18497 ( .B1(n15199), .B2(n16324), .A(n14967), .ZN(P1_U2819) );
  AOI21_X1 U18498 ( .B1(n14970), .B2(n14968), .A(n14953), .ZN(n15211) );
  INV_X1 U18499 ( .A(n15211), .ZN(n15097) );
  NAND3_X1 U18500 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .ZN(n14973) );
  INV_X1 U18501 ( .A(n16342), .ZN(n16319) );
  NOR2_X1 U18502 ( .A1(n14973), .A2(n16319), .ZN(n16308) );
  NAND2_X1 U18503 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n16308), .ZN(n16302) );
  INV_X1 U18504 ( .A(n16302), .ZN(n14975) );
  INV_X1 U18505 ( .A(n14974), .ZN(n14990) );
  NAND2_X1 U18506 ( .A1(n14975), .A2(n14990), .ZN(n16290) );
  OAI21_X1 U18507 ( .B1(n14976), .B2(n16290), .A(n15207), .ZN(n14984) );
  XNOR2_X1 U18508 ( .A(n14993), .B(n14977), .ZN(n15395) );
  INV_X1 U18509 ( .A(n15395), .ZN(n14981) );
  OAI22_X1 U18510 ( .A1(n20306), .A2(n15209), .B1(n14978), .B2(n20335), .ZN(
        n14979) );
  AOI21_X1 U18511 ( .B1(n20321), .B2(P1_EBX_REG_20__SCAN_IN), .A(n14979), .ZN(
        n14980) );
  OAI21_X1 U18512 ( .B1(n14981), .B2(n20351), .A(n14980), .ZN(n14982) );
  AOI21_X1 U18513 ( .B1(n14984), .B2(n14983), .A(n14982), .ZN(n14985) );
  OAI21_X1 U18514 ( .B1(n15097), .B2(n16324), .A(n14985), .ZN(P1_U2820) );
  XNOR2_X1 U18515 ( .A(P1_REIP_REG_18__SCAN_IN), .B(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15002) );
  OAI21_X1 U18516 ( .B1(n14986), .B2(n14987), .A(n14968), .ZN(n15219) );
  INV_X1 U18517 ( .A(n15219), .ZN(n14988) );
  NAND2_X1 U18518 ( .A1(n14988), .A2(n20287), .ZN(n15001) );
  AOI21_X1 U18519 ( .B1(n20347), .B2(n14989), .A(n16345), .ZN(n16316) );
  OAI21_X1 U18520 ( .B1(n14990), .B2(n20312), .A(n16316), .ZN(n16280) );
  OAI21_X1 U18521 ( .B1(n15035), .B2(n15034), .A(n14991), .ZN(n14992) );
  INV_X1 U18522 ( .A(n14992), .ZN(n14994) );
  OR2_X1 U18523 ( .A1(n14994), .A2(n14993), .ZN(n15029) );
  NOR2_X1 U18524 ( .A1(n20340), .A2(n12703), .ZN(n14997) );
  INV_X1 U18525 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15218) );
  NAND2_X1 U18526 ( .A1(n20338), .A2(n15222), .ZN(n14995) );
  OAI211_X1 U18527 ( .C1(n20335), .C2(n15218), .A(n14995), .B(n20289), .ZN(
        n14996) );
  NOR2_X1 U18528 ( .A1(n14997), .A2(n14996), .ZN(n14998) );
  OAI21_X1 U18529 ( .B1(n15029), .B2(n20351), .A(n14998), .ZN(n14999) );
  AOI21_X1 U18530 ( .B1(n16280), .B2(P1_REIP_REG_19__SCAN_IN), .A(n14999), 
        .ZN(n15000) );
  OAI211_X1 U18531 ( .C1(n16290), .C2(n15002), .A(n15001), .B(n15000), .ZN(
        P1_U2821) );
  AOI21_X1 U18532 ( .B1(n15005), .B2(n15003), .A(n15004), .ZN(n15242) );
  INV_X1 U18533 ( .A(n15242), .ZN(n15114) );
  INV_X1 U18534 ( .A(n15035), .ZN(n15006) );
  AOI21_X1 U18535 ( .B1(n15007), .B2(n15046), .A(n15006), .ZN(n15430) );
  INV_X1 U18536 ( .A(n15240), .ZN(n15008) );
  AOI22_X1 U18537 ( .A1(n15008), .A2(n20338), .B1(n20321), .B2(
        P1_EBX_REG_17__SCAN_IN), .ZN(n15009) );
  OAI211_X1 U18538 ( .C1(n20335), .C2(n15010), .A(n15009), .B(n20289), .ZN(
        n15011) );
  AOI21_X1 U18539 ( .B1(n15430), .B2(n20320), .A(n15011), .ZN(n15014) );
  NAND2_X1 U18540 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n16294) );
  NOR2_X1 U18541 ( .A1(n16302), .A2(n16294), .ZN(n15012) );
  OAI21_X1 U18542 ( .B1(n15012), .B2(P1_REIP_REG_17__SCAN_IN), .A(n16280), 
        .ZN(n15013) );
  OAI211_X1 U18543 ( .C1(n15114), .C2(n16324), .A(n15014), .B(n15013), .ZN(
        P1_U2823) );
  OAI22_X1 U18544 ( .A1(n15016), .A2(n15048), .B1(n15047), .B2(n15015), .ZN(
        P1_U2841) );
  AOI22_X1 U18545 ( .A1(n15308), .A2(n15038), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n15037), .ZN(n15017) );
  OAI21_X1 U18546 ( .B1(n15063), .B2(n15040), .A(n15017), .ZN(P1_U2844) );
  AOI22_X1 U18547 ( .A1(n15311), .A2(n15038), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n15037), .ZN(n15018) );
  OAI21_X1 U18548 ( .B1(n15151), .B2(n15040), .A(n15018), .ZN(P1_U2845) );
  INV_X1 U18549 ( .A(n15158), .ZN(n15020) );
  OAI222_X1 U18550 ( .A1(n15040), .A2(n15020), .B1(n15019), .B2(n15047), .C1(
        n15321), .C2(n15048), .ZN(P1_U2846) );
  OAI222_X1 U18551 ( .A1(n15040), .A2(n15166), .B1(n15021), .B2(n15047), .C1(
        n15338), .C2(n15048), .ZN(P1_U2847) );
  AOI22_X1 U18552 ( .A1(n15351), .A2(n15038), .B1(P1_EBX_REG_24__SCAN_IN), 
        .B2(n15037), .ZN(n15022) );
  OAI21_X1 U18553 ( .B1(n15023), .B2(n15040), .A(n15022), .ZN(P1_U2848) );
  INV_X1 U18554 ( .A(n15359), .ZN(n15024) );
  OAI222_X1 U18555 ( .A1(n15040), .A2(n15181), .B1(n15025), .B2(n15047), .C1(
        n15024), .C2(n15048), .ZN(P1_U2849) );
  INV_X1 U18556 ( .A(n15192), .ZN(n15087) );
  OAI222_X1 U18557 ( .A1(n15087), .A2(n15040), .B1(n15026), .B2(n15047), .C1(
        n15048), .C2(n15362), .ZN(P1_U2850) );
  AOI22_X1 U18558 ( .A1(n15383), .A2(n15038), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n15037), .ZN(n15027) );
  OAI21_X1 U18559 ( .B1(n15199), .B2(n15040), .A(n15027), .ZN(P1_U2851) );
  AOI22_X1 U18560 ( .A1(n15395), .A2(n15038), .B1(P1_EBX_REG_20__SCAN_IN), 
        .B2(n15037), .ZN(n15028) );
  OAI21_X1 U18561 ( .B1(n15097), .B2(n15040), .A(n15028), .ZN(P1_U2852) );
  INV_X1 U18562 ( .A(n15029), .ZN(n15404) );
  AOI22_X1 U18563 ( .A1(n15404), .A2(n15038), .B1(P1_EBX_REG_19__SCAN_IN), 
        .B2(n15037), .ZN(n15030) );
  OAI21_X1 U18564 ( .B1(n15219), .B2(n15040), .A(n15030), .ZN(P1_U2853) );
  AND2_X1 U18565 ( .A1(n15032), .A2(n15031), .ZN(n15033) );
  OR2_X1 U18566 ( .A1(n15033), .A2(n14986), .ZN(n16286) );
  XNOR2_X1 U18567 ( .A(n15035), .B(n15034), .ZN(n16285) );
  INV_X1 U18568 ( .A(n16285), .ZN(n15421) );
  AOI22_X1 U18569 ( .A1(n15421), .A2(n15038), .B1(P1_EBX_REG_18__SCAN_IN), 
        .B2(n15037), .ZN(n15036) );
  OAI21_X1 U18570 ( .B1(n16286), .B2(n15040), .A(n15036), .ZN(P1_U2854) );
  AOI22_X1 U18571 ( .A1(n15430), .A2(n15038), .B1(P1_EBX_REG_17__SCAN_IN), 
        .B2(n15037), .ZN(n15039) );
  OAI21_X1 U18572 ( .B1(n15114), .B2(n15040), .A(n15039), .ZN(P1_U2855) );
  NAND2_X1 U18573 ( .A1(n14583), .A2(n15041), .ZN(n15042) );
  AND2_X1 U18574 ( .A1(n15003), .A2(n15042), .ZN(n16349) );
  NAND2_X1 U18575 ( .A1(n15044), .A2(n15043), .ZN(n15045) );
  NAND2_X1 U18576 ( .A1(n15046), .A2(n15045), .ZN(n16292) );
  OAI22_X1 U18577 ( .A1(n16292), .A2(n15048), .B1(n16291), .B2(n15047), .ZN(
        n15049) );
  AOI21_X1 U18578 ( .B1(n16349), .B2(n15050), .A(n15049), .ZN(n15051) );
  INV_X1 U18579 ( .A(n15051), .ZN(P1_U2856) );
  AOI22_X1 U18580 ( .A1(n15110), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15080), .ZN(n15055) );
  OAI211_X1 U18581 ( .C1(n15084), .C2(n16748), .A(n15056), .B(n15055), .ZN(
        P1_U2873) );
  INV_X1 U18582 ( .A(n15110), .ZN(n15123) );
  NAND2_X1 U18583 ( .A1(n15129), .A2(n15115), .ZN(n15059) );
  OAI22_X1 U18584 ( .A1(n15118), .A2(n20396), .B1(n13823), .B2(n15116), .ZN(
        n15057) );
  AOI21_X1 U18585 ( .B1(n15120), .B2(BUF1_REG_30__SCAN_IN), .A(n15057), .ZN(
        n15058) );
  OAI211_X1 U18586 ( .C1(n15123), .C2(n14116), .A(n15059), .B(n15058), .ZN(
        P1_U2874) );
  OAI22_X1 U18587 ( .A1(n15118), .A2(n20390), .B1(n13596), .B2(n15116), .ZN(
        n15060) );
  AOI21_X1 U18588 ( .B1(n15120), .B2(BUF1_REG_28__SCAN_IN), .A(n15060), .ZN(
        n15062) );
  NAND2_X1 U18589 ( .A1(n15110), .A2(DATAI_28_), .ZN(n15061) );
  OAI211_X1 U18590 ( .C1(n15063), .C2(n15113), .A(n15062), .B(n15061), .ZN(
        P1_U2876) );
  OAI22_X1 U18591 ( .A1(n15118), .A2(n20387), .B1(n13588), .B2(n15116), .ZN(
        n15064) );
  AOI21_X1 U18592 ( .B1(n15120), .B2(BUF1_REG_27__SCAN_IN), .A(n15064), .ZN(
        n15066) );
  NAND2_X1 U18593 ( .A1(n15110), .A2(DATAI_27_), .ZN(n15065) );
  OAI211_X1 U18594 ( .C1(n15151), .C2(n15113), .A(n15066), .B(n15065), .ZN(
        P1_U2877) );
  NAND2_X1 U18595 ( .A1(n15158), .A2(n15115), .ZN(n15069) );
  OAI22_X1 U18596 ( .A1(n15118), .A2(n20384), .B1(n13820), .B2(n15116), .ZN(
        n15067) );
  AOI21_X1 U18597 ( .B1(n15120), .B2(BUF1_REG_26__SCAN_IN), .A(n15067), .ZN(
        n15068) );
  OAI211_X1 U18598 ( .C1(n15123), .C2(n21177), .A(n15069), .B(n15068), .ZN(
        P1_U2878) );
  OAI22_X1 U18599 ( .A1(n15118), .A2(n20380), .B1(n13602), .B2(n15116), .ZN(
        n15070) );
  AOI21_X1 U18600 ( .B1(n15120), .B2(BUF1_REG_25__SCAN_IN), .A(n15070), .ZN(
        n15072) );
  NAND2_X1 U18601 ( .A1(n15110), .A2(DATAI_25_), .ZN(n15071) );
  OAI211_X1 U18602 ( .C1(n15166), .C2(n15113), .A(n15072), .B(n15071), .ZN(
        P1_U2879) );
  NAND2_X1 U18603 ( .A1(n15177), .A2(n15115), .ZN(n15075) );
  OAI22_X1 U18604 ( .A1(n15118), .A2(n20377), .B1(n13586), .B2(n15116), .ZN(
        n15073) );
  AOI21_X1 U18605 ( .B1(n15120), .B2(BUF1_REG_24__SCAN_IN), .A(n15073), .ZN(
        n15074) );
  OAI211_X1 U18606 ( .C1(n15123), .C2(n14127), .A(n15075), .B(n15074), .ZN(
        P1_U2880) );
  OAI22_X1 U18607 ( .A1(n15118), .A2(n15076), .B1(n13590), .B2(n15116), .ZN(
        n15077) );
  AOI21_X1 U18608 ( .B1(n15120), .B2(BUF1_REG_23__SCAN_IN), .A(n15077), .ZN(
        n15079) );
  NAND2_X1 U18609 ( .A1(n15110), .A2(DATAI_23_), .ZN(n15078) );
  OAI211_X1 U18610 ( .C1(n15181), .C2(n15113), .A(n15079), .B(n15078), .ZN(
        P1_U2881) );
  INV_X1 U18611 ( .A(n15118), .ZN(n15082) );
  AOI22_X1 U18612 ( .A1(n15082), .A2(n15081), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n15080), .ZN(n15083) );
  OAI21_X1 U18613 ( .B1(n15084), .B2(n16765), .A(n15083), .ZN(n15085) );
  AOI21_X1 U18614 ( .B1(n15110), .B2(DATAI_22_), .A(n15085), .ZN(n15086) );
  OAI21_X1 U18615 ( .B1(n15087), .B2(n15113), .A(n15086), .ZN(P1_U2882) );
  OAI22_X1 U18616 ( .A1(n15118), .A2(n15088), .B1(n13598), .B2(n15116), .ZN(
        n15089) );
  AOI21_X1 U18617 ( .B1(n15120), .B2(BUF1_REG_21__SCAN_IN), .A(n15089), .ZN(
        n15091) );
  NAND2_X1 U18618 ( .A1(n15110), .A2(DATAI_21_), .ZN(n15090) );
  OAI211_X1 U18619 ( .C1(n15199), .C2(n15113), .A(n15091), .B(n15090), .ZN(
        P1_U2883) );
  INV_X1 U18620 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n15092) );
  OAI22_X1 U18621 ( .A1(n15118), .A2(n15093), .B1(n15092), .B2(n15116), .ZN(
        n15094) );
  AOI21_X1 U18622 ( .B1(n15120), .B2(BUF1_REG_20__SCAN_IN), .A(n15094), .ZN(
        n15096) );
  NAND2_X1 U18623 ( .A1(n15110), .A2(DATAI_20_), .ZN(n15095) );
  OAI211_X1 U18624 ( .C1(n15097), .C2(n15113), .A(n15096), .B(n15095), .ZN(
        P1_U2884) );
  OAI22_X1 U18625 ( .A1(n15118), .A2(n15098), .B1(n13594), .B2(n15116), .ZN(
        n15099) );
  AOI21_X1 U18626 ( .B1(n15120), .B2(BUF1_REG_19__SCAN_IN), .A(n15099), .ZN(
        n15101) );
  NAND2_X1 U18627 ( .A1(n15110), .A2(DATAI_19_), .ZN(n15100) );
  OAI211_X1 U18628 ( .C1(n15219), .C2(n15113), .A(n15101), .B(n15100), .ZN(
        P1_U2885) );
  OAI22_X1 U18629 ( .A1(n15118), .A2(n15103), .B1(n15102), .B2(n15116), .ZN(
        n15104) );
  AOI21_X1 U18630 ( .B1(n15120), .B2(BUF1_REG_18__SCAN_IN), .A(n15104), .ZN(
        n15106) );
  NAND2_X1 U18631 ( .A1(n15110), .A2(DATAI_18_), .ZN(n15105) );
  OAI211_X1 U18632 ( .C1(n16286), .C2(n15113), .A(n15106), .B(n15105), .ZN(
        P1_U2886) );
  OAI22_X1 U18633 ( .A1(n15118), .A2(n15108), .B1(n15107), .B2(n15116), .ZN(
        n15109) );
  AOI21_X1 U18634 ( .B1(n15120), .B2(BUF1_REG_17__SCAN_IN), .A(n15109), .ZN(
        n15112) );
  NAND2_X1 U18635 ( .A1(n15110), .A2(DATAI_17_), .ZN(n15111) );
  OAI211_X1 U18636 ( .C1(n15114), .C2(n15113), .A(n15112), .B(n15111), .ZN(
        P1_U2887) );
  NAND2_X1 U18637 ( .A1(n16349), .A2(n15115), .ZN(n15122) );
  OAI22_X1 U18638 ( .A1(n15118), .A2(n15117), .B1(n13816), .B2(n15116), .ZN(
        n15119) );
  AOI21_X1 U18639 ( .B1(n15120), .B2(BUF1_REG_16__SCAN_IN), .A(n15119), .ZN(
        n15121) );
  OAI211_X1 U18640 ( .C1(n15123), .C2(n21187), .A(n15122), .B(n15121), .ZN(
        P1_U2888) );
  INV_X1 U18641 ( .A(n15124), .ZN(n15125) );
  AOI21_X1 U18642 ( .B1(n15125), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n9769), .ZN(n15291) );
  NOR2_X1 U18643 ( .A1(n20432), .A2(n21108), .ZN(n15290) );
  AOI21_X1 U18644 ( .B1(n20416), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15290), .ZN(n15126) );
  OAI21_X1 U18645 ( .B1(n15127), .B2(n20427), .A(n15126), .ZN(n15128) );
  AOI21_X1 U18646 ( .B1(n15129), .B2(n16364), .A(n15128), .ZN(n15130) );
  OAI21_X1 U18647 ( .B1(n15291), .B2(n20238), .A(n15130), .ZN(P1_U2969) );
  NAND2_X1 U18648 ( .A1(n9674), .A2(n15132), .ZN(n15152) );
  NAND2_X1 U18649 ( .A1(n15131), .A2(n15152), .ZN(n15136) );
  OAI21_X1 U18650 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15133), .A(
        n15136), .ZN(n15135) );
  MUX2_X1 U18651 ( .A(n15316), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n9673), .Z(n15134) );
  OAI211_X1 U18652 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15136), .A(
        n15135), .B(n15134), .ZN(n15137) );
  XNOR2_X1 U18653 ( .A(n15137), .B(n15306), .ZN(n15310) );
  OR2_X1 U18654 ( .A1(n20432), .A2(n21038), .ZN(n15305) );
  NAND2_X1 U18655 ( .A1(n20416), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15138) );
  OAI211_X1 U18656 ( .C1(n20427), .C2(n15139), .A(n15305), .B(n15138), .ZN(
        n15140) );
  AOI21_X1 U18657 ( .B1(n15141), .B2(n16364), .A(n15140), .ZN(n15142) );
  OAI21_X1 U18658 ( .B1(n20238), .B2(n15310), .A(n15142), .ZN(P1_U2971) );
  NOR2_X1 U18659 ( .A1(n20432), .A2(n21199), .ZN(n15315) );
  NOR2_X1 U18660 ( .A1(n15254), .A2(n15143), .ZN(n15144) );
  AOI211_X1 U18661 ( .C1(n16355), .C2(n15145), .A(n15315), .B(n15144), .ZN(
        n15150) );
  MUX2_X1 U18662 ( .A(n15147), .B(n15146), .S(n10075), .Z(n15148) );
  XNOR2_X1 U18663 ( .A(n15148), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15312) );
  NAND2_X1 U18664 ( .A1(n15312), .A2(n20422), .ZN(n15149) );
  OAI211_X1 U18665 ( .C1(n15151), .C2(n15258), .A(n15150), .B(n15149), .ZN(
        P1_U2972) );
  OAI211_X1 U18666 ( .C1(n10075), .C2(n15131), .A(n15153), .B(n15152), .ZN(
        n15154) );
  XNOR2_X1 U18667 ( .A(n15154), .B(n15322), .ZN(n15333) );
  NAND2_X1 U18668 ( .A1(n20473), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n15327) );
  NAND2_X1 U18669 ( .A1(n20416), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15155) );
  OAI211_X1 U18670 ( .C1(n20427), .C2(n15156), .A(n15327), .B(n15155), .ZN(
        n15157) );
  AOI21_X1 U18671 ( .B1(n15158), .B2(n16364), .A(n15157), .ZN(n15159) );
  OAI21_X1 U18672 ( .B1(n20238), .B2(n15333), .A(n15159), .ZN(P1_U2973) );
  NAND2_X1 U18673 ( .A1(n15171), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15163) );
  INV_X1 U18674 ( .A(n15131), .ZN(n15161) );
  NAND3_X1 U18675 ( .A1(n15161), .A2(n15343), .A3(n15346), .ZN(n15162) );
  MUX2_X1 U18676 ( .A(n15163), .B(n15162), .S(n10075), .Z(n15164) );
  XNOR2_X1 U18677 ( .A(n15164), .B(n15324), .ZN(n15342) );
  NAND2_X1 U18678 ( .A1(n20473), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15334) );
  OAI21_X1 U18679 ( .B1(n15254), .B2(n15165), .A(n15334), .ZN(n15168) );
  NOR2_X1 U18680 ( .A1(n15166), .A2(n15258), .ZN(n15167) );
  AOI211_X1 U18681 ( .C1(n16355), .C2(n15169), .A(n15168), .B(n15167), .ZN(
        n15170) );
  OAI21_X1 U18682 ( .B1(n20238), .B2(n15342), .A(n15170), .ZN(P1_U2974) );
  NOR2_X1 U18683 ( .A1(n15171), .A2(n15131), .ZN(n15172) );
  MUX2_X1 U18684 ( .A(n15172), .B(n15171), .S(n9674), .Z(n15173) );
  XNOR2_X1 U18685 ( .A(n15173), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15353) );
  OR2_X1 U18686 ( .A1(n20432), .A2(n21047), .ZN(n15347) );
  NAND2_X1 U18687 ( .A1(n20416), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15174) );
  OAI211_X1 U18688 ( .C1(n20427), .C2(n15175), .A(n15347), .B(n15174), .ZN(
        n15176) );
  AOI21_X1 U18689 ( .B1(n15177), .B2(n16364), .A(n15176), .ZN(n15178) );
  OAI21_X1 U18690 ( .B1(n20238), .B2(n15353), .A(n15178), .ZN(P1_U2975) );
  XNOR2_X1 U18691 ( .A(n9673), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15179) );
  XNOR2_X1 U18692 ( .A(n15131), .B(n15179), .ZN(n15361) );
  OR2_X1 U18693 ( .A1(n20432), .A2(n21093), .ZN(n15355) );
  OAI21_X1 U18694 ( .B1(n15254), .B2(n15180), .A(n15355), .ZN(n15183) );
  NOR2_X1 U18695 ( .A1(n15181), .A2(n15258), .ZN(n15182) );
  AOI211_X1 U18696 ( .C1(n16355), .C2(n15184), .A(n15183), .B(n15182), .ZN(
        n15185) );
  OAI21_X1 U18697 ( .B1(n15361), .B2(n20238), .A(n15185), .ZN(P1_U2976) );
  NAND2_X1 U18698 ( .A1(n15187), .A2(n9699), .ZN(n15188) );
  XNOR2_X1 U18699 ( .A(n15188), .B(n15370), .ZN(n15378) );
  NAND2_X1 U18700 ( .A1(n20473), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n15373) );
  NAND2_X1 U18701 ( .A1(n20416), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15189) );
  OAI211_X1 U18702 ( .C1(n20427), .C2(n15190), .A(n15373), .B(n15189), .ZN(
        n15191) );
  AOI21_X1 U18703 ( .B1(n15192), .B2(n16364), .A(n15191), .ZN(n15193) );
  OAI21_X1 U18704 ( .B1(n20238), .B2(n15378), .A(n15193), .ZN(P1_U2977) );
  OAI21_X1 U18705 ( .B1(n15449), .B2(n15419), .A(n15194), .ZN(n15216) );
  NAND2_X1 U18706 ( .A1(n10075), .A2(n15401), .ZN(n15214) );
  NAND2_X1 U18707 ( .A1(n9673), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15213) );
  OAI22_X1 U18708 ( .A1(n15216), .A2(n15214), .B1(n15194), .B2(n15213), .ZN(
        n15205) );
  NAND2_X1 U18709 ( .A1(n15205), .A2(n15368), .ZN(n15204) );
  INV_X1 U18710 ( .A(n15213), .ZN(n15195) );
  NAND2_X1 U18711 ( .A1(n15195), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15196) );
  OAI22_X1 U18712 ( .A1(n15204), .A2(n9673), .B1(n15194), .B2(n15196), .ZN(
        n15197) );
  XNOR2_X1 U18713 ( .A(n15197), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15386) );
  INV_X1 U18714 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15198) );
  NAND2_X1 U18715 ( .A1(n20473), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15379) );
  OAI21_X1 U18716 ( .B1(n15254), .B2(n15198), .A(n15379), .ZN(n15201) );
  NOR2_X1 U18717 ( .A1(n15199), .A2(n15258), .ZN(n15200) );
  AOI211_X1 U18718 ( .C1(n16355), .C2(n15202), .A(n15201), .B(n15200), .ZN(
        n15203) );
  OAI21_X1 U18719 ( .B1(n15386), .B2(n20238), .A(n15203), .ZN(P1_U2978) );
  OAI21_X1 U18720 ( .B1(n15205), .B2(n15368), .A(n15204), .ZN(n15206) );
  INV_X1 U18721 ( .A(n15206), .ZN(n15397) );
  OR2_X1 U18722 ( .A1(n20432), .A2(n15207), .ZN(n15387) );
  NAND2_X1 U18723 ( .A1(n20416), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15208) );
  OAI211_X1 U18724 ( .C1(n20427), .C2(n15209), .A(n15387), .B(n15208), .ZN(
        n15210) );
  AOI21_X1 U18725 ( .B1(n15211), .B2(n16364), .A(n15210), .ZN(n15212) );
  OAI21_X1 U18726 ( .B1(n15397), .B2(n20238), .A(n15212), .ZN(P1_U2979) );
  NAND2_X1 U18727 ( .A1(n15214), .A2(n15213), .ZN(n15215) );
  XNOR2_X1 U18728 ( .A(n15216), .B(n15215), .ZN(n15406) );
  INV_X1 U18729 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n15217) );
  OR2_X1 U18730 ( .A1(n20432), .A2(n15217), .ZN(n15399) );
  OAI21_X1 U18731 ( .B1(n15254), .B2(n15218), .A(n15399), .ZN(n15221) );
  NOR2_X1 U18732 ( .A1(n15219), .A2(n15258), .ZN(n15220) );
  AOI211_X1 U18733 ( .C1(n16355), .C2(n15222), .A(n15221), .B(n15220), .ZN(
        n15223) );
  OAI21_X1 U18734 ( .B1(n20238), .B2(n15406), .A(n15223), .ZN(P1_U2980) );
  OAI21_X1 U18735 ( .B1(n9700), .B2(n15224), .A(n15194), .ZN(n15423) );
  OR2_X1 U18736 ( .A1(n20432), .A2(n20985), .ZN(n15418) );
  OAI21_X1 U18737 ( .B1(n15254), .B2(n15226), .A(n15418), .ZN(n15228) );
  NOR2_X1 U18738 ( .A1(n16286), .A2(n15258), .ZN(n15227) );
  AOI211_X1 U18739 ( .C1(n16355), .C2(n16281), .A(n15228), .B(n15227), .ZN(
        n15229) );
  OAI21_X1 U18740 ( .B1(n20238), .B2(n15423), .A(n15229), .ZN(P1_U2981) );
  NAND2_X1 U18741 ( .A1(n15230), .A2(n15231), .ZN(n15446) );
  INV_X1 U18742 ( .A(n15232), .ZN(n15234) );
  OAI21_X1 U18743 ( .B1(n15446), .B2(n15234), .A(n15233), .ZN(n15235) );
  MUX2_X1 U18744 ( .A(n10075), .B(n15236), .S(n15235), .Z(n15237) );
  XOR2_X1 U18745 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B(n15237), .Z(
        n15432) );
  INV_X1 U18746 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n15238) );
  NOR2_X1 U18747 ( .A1(n20432), .A2(n15238), .ZN(n15429) );
  AOI21_X1 U18748 ( .B1(n20416), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15429), .ZN(n15239) );
  OAI21_X1 U18749 ( .B1(n15240), .B2(n20427), .A(n15239), .ZN(n15241) );
  AOI21_X1 U18750 ( .B1(n15242), .B2(n16364), .A(n15241), .ZN(n15243) );
  OAI21_X1 U18751 ( .B1(n15432), .B2(n20238), .A(n15243), .ZN(P1_U2982) );
  INV_X1 U18752 ( .A(n15230), .ZN(n15247) );
  INV_X1 U18753 ( .A(n15244), .ZN(n15246) );
  AOI21_X1 U18754 ( .B1(n15247), .B2(n15246), .A(n15245), .ZN(n15251) );
  NAND2_X1 U18755 ( .A1(n15251), .A2(n15248), .ZN(n15434) );
  INV_X1 U18756 ( .A(n15433), .ZN(n15252) );
  NOR2_X1 U18757 ( .A1(n15249), .A2(n15252), .ZN(n15250) );
  OAI22_X1 U18758 ( .A1(n15434), .A2(n15252), .B1(n15251), .B2(n15250), .ZN(
        n16390) );
  NAND2_X1 U18759 ( .A1(n16390), .A2(n20422), .ZN(n15257) );
  INV_X1 U18760 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n15253) );
  NOR2_X1 U18761 ( .A1(n20432), .A2(n15253), .ZN(n16386) );
  NOR2_X1 U18762 ( .A1(n15254), .A2(n16301), .ZN(n15255) );
  AOI211_X1 U18763 ( .C1(n16355), .C2(n16306), .A(n16386), .B(n15255), .ZN(
        n15256) );
  OAI211_X1 U18764 ( .C1(n15258), .C2(n16303), .A(n15257), .B(n15256), .ZN(
        P1_U2984) );
  INV_X1 U18765 ( .A(n15444), .ZN(n15260) );
  OAI21_X1 U18766 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n10075), .ZN(n15259) );
  OAI21_X1 U18767 ( .B1(n15230), .B2(n15260), .A(n15259), .ZN(n15271) );
  INV_X1 U18768 ( .A(n15262), .ZN(n15261) );
  OAI21_X1 U18769 ( .B1(n15449), .B2(n15481), .A(n15261), .ZN(n15270) );
  NOR2_X1 U18770 ( .A1(n15271), .A2(n15270), .ZN(n15269) );
  NOR2_X1 U18771 ( .A1(n15269), .A2(n15262), .ZN(n15263) );
  XOR2_X1 U18772 ( .A(n15264), .B(n15263), .Z(n15473) );
  INV_X1 U18773 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20977) );
  NOR2_X1 U18774 ( .A1(n20432), .A2(n20977), .ZN(n15464) );
  AOI21_X1 U18775 ( .B1(n20416), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n15464), .ZN(n15265) );
  OAI21_X1 U18776 ( .B1(n16317), .B2(n20427), .A(n15265), .ZN(n15266) );
  AOI21_X1 U18777 ( .B1(n15267), .B2(n16364), .A(n15266), .ZN(n15268) );
  OAI21_X1 U18778 ( .B1(n15473), .B2(n20238), .A(n15268), .ZN(P1_U2986) );
  AOI21_X1 U18779 ( .B1(n15271), .B2(n15270), .A(n15269), .ZN(n15488) );
  INV_X1 U18780 ( .A(n15272), .ZN(n16336) );
  NAND2_X1 U18781 ( .A1(n20416), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15274) );
  INV_X1 U18782 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15273) );
  OR2_X1 U18783 ( .A1(n20432), .A2(n15273), .ZN(n15480) );
  OAI211_X1 U18784 ( .C1(n20427), .C2(n16331), .A(n15274), .B(n15480), .ZN(
        n15275) );
  AOI21_X1 U18785 ( .B1(n16336), .B2(n16364), .A(n15275), .ZN(n15276) );
  OAI21_X1 U18786 ( .B1(n15488), .B2(n20238), .A(n15276), .ZN(P1_U2987) );
  MUX2_X1 U18787 ( .A(n15277), .B(n15230), .S(n15449), .Z(n15278) );
  XOR2_X1 U18788 ( .A(n12675), .B(n15278), .Z(n16411) );
  INV_X1 U18789 ( .A(n16411), .ZN(n15284) );
  AOI22_X1 U18790 ( .A1(n20416), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20473), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n15279) );
  OAI21_X1 U18791 ( .B1(n15280), .B2(n20427), .A(n15279), .ZN(n15281) );
  AOI21_X1 U18792 ( .B1(n15282), .B2(n16364), .A(n15281), .ZN(n15283) );
  OAI21_X1 U18793 ( .B1(n15284), .B2(n20238), .A(n15283), .ZN(P1_U2989) );
  AOI21_X1 U18794 ( .B1(n15288), .B2(n15287), .A(n15286), .ZN(n15289) );
  INV_X1 U18795 ( .A(n15292), .ZN(n15297) );
  NAND3_X1 U18796 ( .A1(n15317), .A2(n15293), .A3(n15296), .ZN(n15294) );
  OAI211_X1 U18797 ( .C1(n15297), .C2(n15296), .A(n15295), .B(n15294), .ZN(
        n15298) );
  AOI21_X1 U18798 ( .B1(n15299), .B2(n20440), .A(n15298), .ZN(n15300) );
  OAI21_X1 U18799 ( .B1(n15301), .B2(n20470), .A(n15300), .ZN(P1_U3002) );
  AOI21_X1 U18800 ( .B1(n16425), .B2(n15302), .A(n15337), .ZN(n15313) );
  NAND3_X1 U18801 ( .A1(n15317), .A2(n10108), .A3(n15303), .ZN(n15304) );
  OAI211_X1 U18802 ( .C1(n15313), .C2(n15306), .A(n15305), .B(n15304), .ZN(
        n15307) );
  AOI21_X1 U18803 ( .B1(n15308), .B2(n20440), .A(n15307), .ZN(n15309) );
  OAI21_X1 U18804 ( .B1(n15310), .B2(n20470), .A(n15309), .ZN(P1_U3003) );
  INV_X1 U18805 ( .A(n15311), .ZN(n15320) );
  NAND2_X1 U18806 ( .A1(n15312), .A2(n20452), .ZN(n15319) );
  NOR2_X1 U18807 ( .A1(n15313), .A2(n15316), .ZN(n15314) );
  AOI211_X1 U18808 ( .C1(n15317), .C2(n15316), .A(n15315), .B(n15314), .ZN(
        n15318) );
  OAI211_X1 U18809 ( .C1(n20469), .C2(n15320), .A(n15319), .B(n15318), .ZN(
        P1_U3004) );
  INV_X1 U18810 ( .A(n15321), .ZN(n15331) );
  NAND2_X1 U18811 ( .A1(n15323), .A2(n15322), .ZN(n15329) );
  NAND2_X1 U18812 ( .A1(n15325), .A2(n15324), .ZN(n15326) );
  NOR2_X1 U18813 ( .A1(n15357), .A2(n15326), .ZN(n15335) );
  OAI21_X1 U18814 ( .B1(n15337), .B2(n15335), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15328) );
  OAI211_X1 U18815 ( .C1(n15357), .C2(n15329), .A(n15328), .B(n15327), .ZN(
        n15330) );
  AOI21_X1 U18816 ( .B1(n15331), .B2(n20440), .A(n15330), .ZN(n15332) );
  OAI21_X1 U18817 ( .B1(n15333), .B2(n20470), .A(n15332), .ZN(P1_U3005) );
  INV_X1 U18818 ( .A(n15334), .ZN(n15336) );
  AOI211_X1 U18819 ( .C1(n15337), .C2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15336), .B(n15335), .ZN(n15341) );
  INV_X1 U18820 ( .A(n15338), .ZN(n15339) );
  NAND2_X1 U18821 ( .A1(n15339), .A2(n20440), .ZN(n15340) );
  OAI211_X1 U18822 ( .C1(n15342), .C2(n20470), .A(n15341), .B(n15340), .ZN(
        P1_U3006) );
  NAND2_X1 U18823 ( .A1(n15343), .A2(n15479), .ZN(n15344) );
  AOI21_X1 U18824 ( .B1(n15345), .B2(n15344), .A(n15346), .ZN(n15350) );
  NAND2_X1 U18825 ( .A1(n15346), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15348) );
  OAI21_X1 U18826 ( .B1(n15357), .B2(n15348), .A(n15347), .ZN(n15349) );
  AOI211_X1 U18827 ( .C1(n15351), .C2(n20440), .A(n15350), .B(n15349), .ZN(
        n15352) );
  OAI21_X1 U18828 ( .B1(n15353), .B2(n20470), .A(n15352), .ZN(P1_U3007) );
  NAND2_X1 U18829 ( .A1(n15354), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15356) );
  OAI211_X1 U18830 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n15357), .A(
        n15356), .B(n15355), .ZN(n15358) );
  AOI21_X1 U18831 ( .B1(n15359), .B2(n20440), .A(n15358), .ZN(n15360) );
  OAI21_X1 U18832 ( .B1(n15361), .B2(n20470), .A(n15360), .ZN(P1_U3008) );
  INV_X1 U18833 ( .A(n15362), .ZN(n15376) );
  AND2_X1 U18834 ( .A1(n15465), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n15407) );
  NAND2_X1 U18835 ( .A1(n20466), .A2(n15407), .ZN(n15364) );
  NAND2_X1 U18836 ( .A1(n15364), .A2(n15363), .ZN(n15414) );
  INV_X1 U18837 ( .A(n15465), .ZN(n15365) );
  NOR2_X1 U18838 ( .A1(n20475), .A2(n15365), .ZN(n15367) );
  OAI21_X1 U18839 ( .B1(n15414), .B2(n15367), .A(n15366), .ZN(n15369) );
  NOR4_X1 U18840 ( .A1(n15369), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15401), .A4(n15368), .ZN(n15380) );
  OAI21_X1 U18841 ( .B1(n15382), .B2(n15380), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15374) );
  INV_X1 U18842 ( .A(n15369), .ZN(n15398) );
  NAND3_X1 U18843 ( .A1(n15398), .A2(n15371), .A3(n15370), .ZN(n15372) );
  NAND3_X1 U18844 ( .A1(n15374), .A2(n15373), .A3(n15372), .ZN(n15375) );
  AOI21_X1 U18845 ( .B1(n15376), .B2(n20440), .A(n15375), .ZN(n15377) );
  OAI21_X1 U18846 ( .B1(n15378), .B2(n20470), .A(n15377), .ZN(P1_U3009) );
  INV_X1 U18847 ( .A(n15379), .ZN(n15381) );
  AOI211_X1 U18848 ( .C1(n15382), .C2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15381), .B(n15380), .ZN(n15385) );
  NAND2_X1 U18849 ( .A1(n15383), .A2(n20440), .ZN(n15384) );
  OAI211_X1 U18850 ( .C1(n15386), .C2(n20470), .A(n15385), .B(n15384), .ZN(
        P1_U3010) );
  INV_X1 U18851 ( .A(n15387), .ZN(n15394) );
  INV_X1 U18852 ( .A(n20475), .ZN(n15390) );
  INV_X1 U18853 ( .A(n15388), .ZN(n15389) );
  OAI21_X1 U18854 ( .B1(n15414), .B2(n15390), .A(n15389), .ZN(n15392) );
  AOI21_X1 U18855 ( .B1(n15398), .B2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15391) );
  AOI21_X1 U18856 ( .B1(n15402), .B2(n15392), .A(n15391), .ZN(n15393) );
  AOI211_X1 U18857 ( .C1(n15395), .C2(n20440), .A(n15394), .B(n15393), .ZN(
        n15396) );
  OAI21_X1 U18858 ( .B1(n15397), .B2(n20470), .A(n15396), .ZN(P1_U3011) );
  NAND2_X1 U18859 ( .A1(n15398), .A2(n15401), .ZN(n15400) );
  OAI211_X1 U18860 ( .C1(n15402), .C2(n15401), .A(n15400), .B(n15399), .ZN(
        n15403) );
  AOI21_X1 U18861 ( .B1(n15404), .B2(n20440), .A(n15403), .ZN(n15405) );
  OAI21_X1 U18862 ( .B1(n15406), .B2(n20470), .A(n15405), .ZN(P1_U3012) );
  INV_X1 U18863 ( .A(n15407), .ZN(n15408) );
  NAND2_X1 U18864 ( .A1(n20466), .A2(n15408), .ZN(n15412) );
  AND2_X1 U18865 ( .A1(n15465), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15409) );
  OR2_X1 U18866 ( .A1(n20475), .A2(n15409), .ZN(n15463) );
  OR2_X1 U18867 ( .A1(n20428), .A2(n15457), .ZN(n15410) );
  NAND4_X1 U18868 ( .A1(n15412), .A2(n15463), .A3(n15411), .A4(n15410), .ZN(
        n15462) );
  INV_X1 U18869 ( .A(n15462), .ZN(n15415) );
  NAND2_X1 U18870 ( .A1(n15414), .A2(n15413), .ZN(n15467) );
  NAND2_X1 U18871 ( .A1(n15415), .A2(n15467), .ZN(n15453) );
  AOI21_X1 U18872 ( .B1(n16425), .B2(n15416), .A(n15453), .ZN(n15425) );
  OR3_X1 U18873 ( .A1(n15424), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15416), .ZN(n15417) );
  OAI211_X1 U18874 ( .C1(n15425), .C2(n15419), .A(n15418), .B(n15417), .ZN(
        n15420) );
  AOI21_X1 U18875 ( .B1(n15421), .B2(n20440), .A(n15420), .ZN(n15422) );
  OAI21_X1 U18876 ( .B1(n15423), .B2(n20470), .A(n15422), .ZN(P1_U3013) );
  INV_X1 U18877 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15427) );
  NOR2_X1 U18878 ( .A1(n15424), .A2(n15456), .ZN(n15437) );
  NAND3_X1 U18879 ( .A1(n15437), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15426) );
  AOI21_X1 U18880 ( .B1(n15427), .B2(n15426), .A(n15425), .ZN(n15428) );
  AOI211_X1 U18881 ( .C1(n15430), .C2(n20440), .A(n15429), .B(n15428), .ZN(
        n15431) );
  OAI21_X1 U18882 ( .B1(n15432), .B2(n20470), .A(n15431), .ZN(P1_U3014) );
  NAND2_X1 U18883 ( .A1(n15434), .A2(n15433), .ZN(n15436) );
  XNOR2_X1 U18884 ( .A(n15436), .B(n15435), .ZN(n16350) );
  NAND2_X1 U18885 ( .A1(n16350), .A2(n20452), .ZN(n15443) );
  AOI21_X1 U18886 ( .B1(n15456), .B2(n16425), .A(n15453), .ZN(n16394) );
  NAND2_X1 U18887 ( .A1(n15437), .A2(n16393), .ZN(n16388) );
  NAND2_X1 U18888 ( .A1(n15437), .A2(n15439), .ZN(n15438) );
  OAI211_X1 U18889 ( .C1(n16394), .C2(n15439), .A(n16388), .B(n15438), .ZN(
        n15441) );
  NAND2_X1 U18890 ( .A1(n16393), .A2(n15439), .ZN(n15440) );
  AOI22_X1 U18891 ( .A1(n15441), .A2(n15440), .B1(n20473), .B2(
        P1_REIP_REG_16__SCAN_IN), .ZN(n15442) );
  OAI211_X1 U18892 ( .C1(n20469), .C2(n16292), .A(n15443), .B(n15442), .ZN(
        P1_U3015) );
  NAND3_X1 U18893 ( .A1(n15446), .A2(n15445), .A3(n15444), .ZN(n15448) );
  NAND2_X1 U18894 ( .A1(n15448), .A2(n15447), .ZN(n15451) );
  XNOR2_X1 U18895 ( .A(n15449), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15450) );
  XNOR2_X1 U18896 ( .A(n15451), .B(n15450), .ZN(n16359) );
  INV_X1 U18897 ( .A(n15452), .ZN(n16309) );
  INV_X1 U18898 ( .A(n15453), .ZN(n15455) );
  INV_X1 U18899 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n15454) );
  OAI22_X1 U18900 ( .A1(n15455), .A2(n15456), .B1(n20432), .B2(n15454), .ZN(
        n15460) );
  NAND2_X1 U18901 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n15479), .ZN(
        n20465) );
  NAND2_X1 U18902 ( .A1(n16424), .A2(n20428), .ZN(n16446) );
  NAND3_X1 U18903 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15457), .A3(
        n15456), .ZN(n15458) );
  NOR2_X1 U18904 ( .A1(n15474), .A2(n15458), .ZN(n15459) );
  AOI211_X1 U18905 ( .C1(n20440), .C2(n16309), .A(n15460), .B(n15459), .ZN(
        n15461) );
  OAI21_X1 U18906 ( .B1(n16359), .B2(n20470), .A(n15461), .ZN(P1_U3017) );
  INV_X1 U18907 ( .A(n16320), .ZN(n15471) );
  NAND2_X1 U18908 ( .A1(n15462), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15469) );
  INV_X1 U18909 ( .A(n15463), .ZN(n15466) );
  AOI21_X1 U18910 ( .B1(n15466), .B2(n15465), .A(n15464), .ZN(n15468) );
  NAND3_X1 U18911 ( .A1(n15469), .A2(n15468), .A3(n15467), .ZN(n15470) );
  AOI21_X1 U18912 ( .B1(n15471), .B2(n20440), .A(n15470), .ZN(n15472) );
  OAI21_X1 U18913 ( .B1(n15473), .B2(n20470), .A(n15472), .ZN(P1_U3018) );
  INV_X1 U18914 ( .A(n16428), .ZN(n16445) );
  NOR2_X1 U18915 ( .A1(n16445), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15486) );
  NOR2_X1 U18916 ( .A1(n16333), .A2(n20469), .ZN(n15484) );
  OAI21_X1 U18917 ( .B1(n15476), .B2(n15475), .A(n20450), .ZN(n15478) );
  AOI21_X1 U18918 ( .B1(n20467), .B2(n15477), .A(n20449), .ZN(n16405) );
  OAI211_X1 U18919 ( .C1(n15485), .C2(n20428), .A(n15478), .B(n16405), .ZN(
        n16397) );
  AOI21_X1 U18920 ( .B1(n15479), .B2(n16395), .A(n16397), .ZN(n15482) );
  OAI21_X1 U18921 ( .B1(n15482), .B2(n15481), .A(n15480), .ZN(n15483) );
  AOI211_X1 U18922 ( .C1(n15486), .C2(n15485), .A(n15484), .B(n15483), .ZN(
        n15487) );
  OAI21_X1 U18923 ( .B1(n15488), .B2(n20470), .A(n15487), .ZN(P1_U3019) );
  OAI21_X1 U18924 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15489), .A(n20810), 
        .ZN(n15490) );
  OAI21_X1 U18925 ( .B1(n15493), .B2(n14392), .A(n15490), .ZN(n15491) );
  MUX2_X1 U18926 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15491), .S(
        n20478), .Z(P1_U3477) );
  INV_X1 U18927 ( .A(n20810), .ZN(n20566) );
  MUX2_X1 U18928 ( .A(n20884), .B(n20566), .S(n13949), .Z(n15492) );
  OAI21_X1 U18929 ( .B1(n15493), .B2(n13542), .A(n15492), .ZN(n15494) );
  MUX2_X1 U18930 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15494), .S(
        n20478), .Z(P1_U3476) );
  NOR3_X1 U18931 ( .A1(n11897), .A2(n13875), .A3(n13559), .ZN(n15497) );
  NOR2_X1 U18932 ( .A1(n14392), .A2(n15495), .ZN(n15496) );
  AOI211_X1 U18933 ( .C1(n16217), .C2(n11742), .A(n15497), .B(n15496), .ZN(
        n16221) );
  INV_X1 U18934 ( .A(n15498), .ZN(n16454) );
  NOR3_X1 U18935 ( .A1(n13875), .A2(n13559), .A3(n16251), .ZN(n15499) );
  AOI21_X1 U18936 ( .B1(n15501), .B2(n15500), .A(n15499), .ZN(n15502) );
  OAI21_X1 U18937 ( .B1(n16221), .B2(n16454), .A(n15502), .ZN(n15503) );
  MUX2_X1 U18938 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15503), .S(
        n16460), .Z(P1_U3473) );
  INV_X1 U18939 ( .A(n15504), .ZN(n15505) );
  OAI22_X1 U18940 ( .A1(n15506), .A2(n16454), .B1(n16251), .B2(n15505), .ZN(
        n15507) );
  MUX2_X1 U18941 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n15507), .S(
        n16460), .Z(P1_U3469) );
  OAI21_X1 U18942 ( .B1(n15564), .B2(n15509), .A(n15508), .ZN(n15850) );
  NOR2_X1 U18943 ( .A1(n15527), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15510) );
  OR2_X1 U18944 ( .A1(n15529), .A2(n15510), .ZN(n16526) );
  AOI21_X1 U18945 ( .B1(n15794), .B2(n15511), .A(n15523), .ZN(n19267) );
  AOI21_X1 U18946 ( .B1(n15519), .B2(n15813), .A(n15521), .ZN(n19290) );
  AOI21_X1 U18947 ( .B1(n16591), .B2(n15517), .A(n15520), .ZN(n19321) );
  AOI21_X1 U18948 ( .B1(n15512), .B2(n15515), .A(n15518), .ZN(n19348) );
  AOI21_X1 U18949 ( .B1(n16619), .B2(n15513), .A(n15516), .ZN(n19373) );
  NAND2_X1 U18950 ( .A1(n15514), .A2(n16632), .ZN(n19371) );
  NOR2_X1 U18951 ( .A1(n19373), .A2(n19371), .ZN(n19353) );
  OAI21_X1 U18952 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n15516), .A(
        n15515), .ZN(n19354) );
  NAND2_X1 U18953 ( .A1(n19353), .A2(n19354), .ZN(n19338) );
  NOR2_X1 U18954 ( .A1(n19348), .A2(n19338), .ZN(n19337) );
  OAI21_X1 U18955 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n15518), .A(
        n15517), .ZN(n19327) );
  NAND2_X1 U18956 ( .A1(n19337), .A2(n19327), .ZN(n19319) );
  NOR2_X1 U18957 ( .A1(n19321), .A2(n19319), .ZN(n19301) );
  OAI21_X1 U18958 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n15520), .A(
        n15519), .ZN(n19302) );
  NAND2_X1 U18959 ( .A1(n19301), .A2(n19302), .ZN(n19288) );
  NOR2_X1 U18960 ( .A1(n19290), .A2(n19288), .ZN(n19274) );
  OAI21_X1 U18961 ( .B1(n15521), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15511), .ZN(n19275) );
  NAND2_X1 U18962 ( .A1(n19274), .A2(n19275), .ZN(n19266) );
  NOR2_X1 U18963 ( .A1(n19267), .A2(n19266), .ZN(n19256) );
  OAI21_X1 U18964 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n15523), .A(
        n15522), .ZN(n19260) );
  NAND2_X1 U18965 ( .A1(n19256), .A2(n19260), .ZN(n19237) );
  OAI21_X1 U18966 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n15524), .A(
        n15525), .ZN(n16585) );
  AOI21_X1 U18967 ( .B1(n15525), .B2(n9812), .A(n15526), .ZN(n15768) );
  INV_X1 U18968 ( .A(n15768), .ZN(n16566) );
  NAND2_X1 U18969 ( .A1(n14305), .A2(n16564), .ZN(n16553) );
  OAI21_X1 U18970 ( .B1(n15526), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15528), .ZN(n16554) );
  AOI21_X1 U18971 ( .B1(n16533), .B2(n15528), .A(n15527), .ZN(n15752) );
  INV_X1 U18972 ( .A(n15752), .ZN(n16540) );
  INV_X1 U18973 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16504) );
  INV_X1 U18974 ( .A(n15529), .ZN(n15530) );
  AOI21_X1 U18975 ( .B1(n16504), .B2(n15530), .A(n15531), .ZN(n15728) );
  INV_X1 U18976 ( .A(n15728), .ZN(n16513) );
  NAND2_X1 U18977 ( .A1(n19384), .A2(n16511), .ZN(n15534) );
  OR2_X1 U18978 ( .A1(n15531), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15532) );
  NAND2_X1 U18979 ( .A1(n15533), .A2(n15532), .ZN(n15721) );
  OAI211_X1 U18980 ( .C1(n15534), .C2(n15721), .A(n19443), .B(n16469), .ZN(
        n15545) );
  INV_X1 U18981 ( .A(n15535), .ZN(n15543) );
  OR2_X1 U18982 ( .A1(n15536), .A2(n15537), .ZN(n15538) );
  INV_X1 U18983 ( .A(n15848), .ZN(n15540) );
  INV_X1 U18984 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15539) );
  OAI22_X1 U18985 ( .A1(n15540), .A2(n19447), .B1(n15539), .B2(n19397), .ZN(
        n15542) );
  OAI22_X1 U18986 ( .A1(n19413), .A2(n10774), .B1(n15720), .B2(n19417), .ZN(
        n15541) );
  AOI211_X1 U18987 ( .C1(n15543), .C2(n19403), .A(n15542), .B(n15541), .ZN(
        n15544) );
  OAI211_X1 U18988 ( .C1(n15850), .C2(n19422), .A(n15545), .B(n15544), .ZN(
        P2_U2827) );
  INV_X1 U18989 ( .A(n15702), .ZN(n16475) );
  MUX2_X1 U18990 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n16475), .S(n15616), .Z(
        P2_U2856) );
  XNOR2_X1 U18991 ( .A(n15546), .B(n15547), .ZN(n15626) );
  NAND2_X1 U18992 ( .A1(n13835), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15549) );
  NAND2_X1 U18993 ( .A1(n16494), .A2(n15616), .ZN(n15548) );
  OAI211_X1 U18994 ( .C1(n15626), .C2(n15618), .A(n15549), .B(n15548), .ZN(
        P2_U2858) );
  INV_X1 U18995 ( .A(n15550), .ZN(n15551) );
  NOR2_X1 U18996 ( .A1(n15552), .A2(n15551), .ZN(n15554) );
  XNOR2_X1 U18997 ( .A(n15554), .B(n15553), .ZN(n15631) );
  NOR2_X1 U18998 ( .A1(n15850), .A2(n13835), .ZN(n15555) );
  AOI21_X1 U18999 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n13835), .A(n15555), .ZN(
        n15556) );
  OAI21_X1 U19000 ( .B1(n15631), .B2(n15618), .A(n15556), .ZN(P2_U2859) );
  AOI21_X1 U19001 ( .B1(n15559), .B2(n15558), .A(n15557), .ZN(n15560) );
  INV_X1 U19002 ( .A(n15560), .ZN(n15640) );
  NOR2_X1 U19003 ( .A1(n15561), .A2(n15562), .ZN(n15563) );
  NOR2_X1 U19004 ( .A1(n16509), .A2(n13835), .ZN(n15565) );
  AOI21_X1 U19005 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n13835), .A(n15565), .ZN(
        n15566) );
  OAI21_X1 U19006 ( .B1(n15640), .B2(n15618), .A(n15566), .ZN(P2_U2860) );
  OAI21_X1 U19007 ( .B1(n15569), .B2(n15568), .A(n15567), .ZN(n15649) );
  NOR2_X1 U19008 ( .A1(n15570), .A2(n15571), .ZN(n15572) );
  OR2_X1 U19009 ( .A1(n15561), .A2(n15572), .ZN(n16522) );
  NOR2_X1 U19010 ( .A1(n16522), .A2(n13835), .ZN(n15573) );
  AOI21_X1 U19011 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n13835), .A(n15573), .ZN(
        n15574) );
  OAI21_X1 U19012 ( .B1(n15649), .B2(n15618), .A(n15574), .ZN(P2_U2861) );
  INV_X1 U19013 ( .A(n15576), .ZN(n15577) );
  AOI21_X1 U19014 ( .B1(n15579), .B2(n15578), .A(n15577), .ZN(n15580) );
  INV_X1 U19015 ( .A(n15580), .ZN(n15658) );
  AOI21_X1 U19016 ( .B1(n15581), .B2(n9740), .A(n15570), .ZN(n16537) );
  INV_X1 U19017 ( .A(n16537), .ZN(n15881) );
  NOR2_X1 U19018 ( .A1(n15881), .A2(n13835), .ZN(n15582) );
  AOI21_X1 U19019 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n13835), .A(n15582), .ZN(
        n15583) );
  OAI21_X1 U19020 ( .B1(n15658), .B2(n15618), .A(n15583), .ZN(P2_U2862) );
  OAI21_X1 U19021 ( .B1(n15586), .B2(n15585), .A(n15584), .ZN(n15587) );
  XOR2_X1 U19022 ( .A(n15587), .B(n9779), .Z(n15665) );
  NAND2_X1 U19023 ( .A1(n9788), .A2(n15588), .ZN(n15589) );
  NAND2_X1 U19024 ( .A1(n9740), .A2(n15589), .ZN(n16549) );
  NOR2_X1 U19025 ( .A1(n16549), .A2(n13835), .ZN(n15590) );
  AOI21_X1 U19026 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n13835), .A(n15590), .ZN(
        n15591) );
  OAI21_X1 U19027 ( .B1(n15665), .B2(n15618), .A(n15591), .ZN(P2_U2863) );
  AOI21_X1 U19028 ( .B1(n15594), .B2(n15593), .A(n15592), .ZN(n15595) );
  INV_X1 U19029 ( .A(n15595), .ZN(n15672) );
  NAND2_X1 U19030 ( .A1(n13835), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n15599) );
  XOR2_X1 U19031 ( .A(n15597), .B(n15596), .Z(n16563) );
  NAND2_X1 U19032 ( .A1(n16563), .A2(n15616), .ZN(n15598) );
  OAI211_X1 U19033 ( .C1(n15672), .C2(n15618), .A(n15599), .B(n15598), .ZN(
        P2_U2864) );
  AOI21_X1 U19034 ( .B1(n15601), .B2(n15600), .A(n13004), .ZN(n15602) );
  INV_X1 U19035 ( .A(n15602), .ZN(n15679) );
  OR2_X1 U19036 ( .A1(n13219), .A2(n15603), .ZN(n15604) );
  NAND2_X1 U19037 ( .A1(n15596), .A2(n15604), .ZN(n16578) );
  NOR2_X1 U19038 ( .A1(n16578), .A2(n13835), .ZN(n15605) );
  AOI21_X1 U19039 ( .B1(P2_EBX_REG_22__SCAN_IN), .B2(n13835), .A(n15605), .ZN(
        n15606) );
  OAI21_X1 U19040 ( .B1(n15679), .B2(n15618), .A(n15606), .ZN(P2_U2865) );
  NAND2_X1 U19041 ( .A1(n15607), .A2(n15608), .ZN(n15609) );
  NAND2_X1 U19042 ( .A1(n15600), .A2(n15609), .ZN(n15685) );
  MUX2_X1 U19043 ( .A(n15610), .B(n10011), .S(n13835), .Z(n15611) );
  OAI21_X1 U19044 ( .B1(n15685), .B2(n15618), .A(n15611), .ZN(P2_U2866) );
  OAI21_X1 U19045 ( .B1(n14641), .B2(n15612), .A(n15607), .ZN(n15697) );
  AND2_X1 U19046 ( .A1(n9748), .A2(n15613), .ZN(n15614) );
  NOR2_X1 U19047 ( .A1(n13220), .A2(n15614), .ZN(n19250) );
  NOR2_X1 U19048 ( .A1(n15616), .A2(n19248), .ZN(n15615) );
  AOI21_X1 U19049 ( .B1(n19250), .B2(n15616), .A(n15615), .ZN(n15617) );
  OAI21_X1 U19050 ( .B1(n15697), .B2(n15618), .A(n15617), .ZN(P2_U2867) );
  XOR2_X1 U19051 ( .A(n15620), .B(n15619), .Z(n16493) );
  AOI22_X1 U19052 ( .A1(n19451), .A2(BUF1_REG_29__SCAN_IN), .B1(n19449), .B2(
        n16493), .ZN(n15625) );
  OAI22_X1 U19053 ( .A1(n15622), .A2(n15690), .B1(n15689), .B2(n15621), .ZN(
        n15623) );
  AOI21_X1 U19054 ( .B1(n19450), .B2(BUF2_REG_29__SCAN_IN), .A(n15623), .ZN(
        n15624) );
  OAI211_X1 U19055 ( .C1(n15626), .C2(n19465), .A(n15625), .B(n15624), .ZN(
        P2_U2890) );
  AOI22_X1 U19056 ( .A1(n19451), .A2(BUF1_REG_28__SCAN_IN), .B1(n19449), .B2(
        n15848), .ZN(n15630) );
  OAI22_X1 U19057 ( .A1(n15627), .A2(n15690), .B1(n15689), .B2(n13728), .ZN(
        n15628) );
  AOI21_X1 U19058 ( .B1(n19450), .B2(BUF2_REG_28__SCAN_IN), .A(n15628), .ZN(
        n15629) );
  OAI211_X1 U19059 ( .C1(n15631), .C2(n19465), .A(n15630), .B(n15629), .ZN(
        P2_U2891) );
  AND2_X1 U19060 ( .A1(n15632), .A2(n15633), .ZN(n15634) );
  NOR2_X1 U19061 ( .A1(n15536), .A2(n15634), .ZN(n16507) );
  AOI22_X1 U19062 ( .A1(n19451), .A2(BUF1_REG_27__SCAN_IN), .B1(n19449), .B2(
        n16507), .ZN(n15639) );
  OAI22_X1 U19063 ( .A1(n15636), .A2(n15690), .B1(n15689), .B2(n15635), .ZN(
        n15637) );
  AOI21_X1 U19064 ( .B1(n19450), .B2(BUF2_REG_27__SCAN_IN), .A(n15637), .ZN(
        n15638) );
  OAI211_X1 U19065 ( .C1(n15640), .C2(n19465), .A(n15639), .B(n15638), .ZN(
        P2_U2892) );
  OAI21_X1 U19066 ( .B1(n15641), .B2(n15642), .A(n15632), .ZN(n16521) );
  INV_X1 U19067 ( .A(n16521), .ZN(n15643) );
  AOI22_X1 U19068 ( .A1(n19451), .A2(BUF1_REG_26__SCAN_IN), .B1(n19449), .B2(
        n15643), .ZN(n15648) );
  OAI22_X1 U19069 ( .A1(n15645), .A2(n15690), .B1(n15689), .B2(n15644), .ZN(
        n15646) );
  AOI21_X1 U19070 ( .B1(n19450), .B2(BUF2_REG_26__SCAN_IN), .A(n15646), .ZN(
        n15647) );
  OAI211_X1 U19071 ( .C1(n15649), .C2(n19465), .A(n15648), .B(n15647), .ZN(
        P2_U2893) );
  NOR2_X1 U19072 ( .A1(n15651), .A2(n15650), .ZN(n15652) );
  NOR2_X1 U19073 ( .A1(n15652), .A2(n15641), .ZN(n16536) );
  AOI22_X1 U19074 ( .A1(n19451), .A2(BUF1_REG_25__SCAN_IN), .B1(n19449), .B2(
        n16536), .ZN(n15657) );
  OAI22_X1 U19075 ( .A1(n15654), .A2(n15690), .B1(n15689), .B2(n15653), .ZN(
        n15655) );
  AOI21_X1 U19076 ( .B1(n19450), .B2(BUF2_REG_25__SCAN_IN), .A(n15655), .ZN(
        n15656) );
  OAI211_X1 U19077 ( .C1(n15658), .C2(n19465), .A(n15657), .B(n15656), .ZN(
        P2_U2894) );
  XNOR2_X1 U19078 ( .A(n15659), .B(n9741), .ZN(n16557) );
  INV_X1 U19079 ( .A(n16557), .ZN(n15660) );
  AOI22_X1 U19080 ( .A1(n19451), .A2(BUF1_REG_24__SCAN_IN), .B1(n19449), .B2(
        n15660), .ZN(n15664) );
  OAI22_X1 U19081 ( .A1(n15661), .A2(n15690), .B1(n15689), .B2(n13509), .ZN(
        n15662) );
  AOI21_X1 U19082 ( .B1(n19450), .B2(BUF2_REG_24__SCAN_IN), .A(n15662), .ZN(
        n15663) );
  OAI211_X1 U19083 ( .C1(n15665), .C2(n19465), .A(n15664), .B(n15663), .ZN(
        P2_U2895) );
  OAI22_X1 U19084 ( .A1(n19567), .A2(n15690), .B1(n15689), .B2(n15666), .ZN(
        n15670) );
  OAI21_X1 U19085 ( .B1(n15668), .B2(n15667), .A(n9741), .ZN(n16561) );
  OAI22_X1 U19086 ( .A1(n15693), .A2(n16763), .B1(n15675), .B2(n16561), .ZN(
        n15669) );
  AOI211_X1 U19087 ( .C1(n19450), .C2(BUF2_REG_23__SCAN_IN), .A(n15670), .B(
        n15669), .ZN(n15671) );
  OAI21_X1 U19088 ( .B1(n15672), .B2(n19465), .A(n15671), .ZN(P2_U2896) );
  OAI22_X1 U19089 ( .A1(n19559), .A2(n15690), .B1(n15689), .B2(n13506), .ZN(
        n15677) );
  AOI21_X1 U19090 ( .B1(n15674), .B2(n15673), .A(n15667), .ZN(n15919) );
  INV_X1 U19091 ( .A(n15919), .ZN(n16205) );
  OAI22_X1 U19092 ( .A1(n15693), .A2(n16765), .B1(n15675), .B2(n16205), .ZN(
        n15676) );
  AOI211_X1 U19093 ( .C1(n19450), .C2(BUF2_REG_22__SCAN_IN), .A(n15677), .B(
        n15676), .ZN(n15678) );
  OAI21_X1 U19094 ( .B1(n15679), .B2(n19465), .A(n15678), .ZN(P2_U2897) );
  OAI22_X1 U19095 ( .A1(n19552), .A2(n15690), .B1(n15689), .B2(n15680), .ZN(
        n15683) );
  INV_X1 U19096 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15681) );
  OAI22_X1 U19097 ( .A1(n15693), .A2(n19550), .B1(n15692), .B2(n15681), .ZN(
        n15682) );
  AOI211_X1 U19098 ( .C1(n19242), .C2(n19449), .A(n15683), .B(n15682), .ZN(
        n15684) );
  OAI21_X1 U19099 ( .B1(n19465), .B2(n15685), .A(n15684), .ZN(P2_U2898) );
  NOR2_X1 U19100 ( .A1(n14636), .A2(n15686), .ZN(n15687) );
  OAI22_X1 U19101 ( .A1(n15690), .A2(n19547), .B1(n15689), .B2(n13418), .ZN(
        n15695) );
  INV_X1 U19102 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n15691) );
  OAI22_X1 U19103 ( .A1(n15693), .A2(n16768), .B1(n15692), .B2(n15691), .ZN(
        n15694) );
  AOI211_X1 U19104 ( .C1(n9778), .C2(n19449), .A(n15695), .B(n15694), .ZN(
        n15696) );
  OAI21_X1 U19105 ( .B1(n19465), .B2(n15697), .A(n15696), .ZN(P2_U2899) );
  NOR2_X1 U19106 ( .A1(n19510), .A2(n15698), .ZN(n15699) );
  AOI211_X1 U19107 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n19501), .A(
        n15700), .B(n15699), .ZN(n15701) );
  OAI21_X1 U19108 ( .B1(n15702), .B2(n16655), .A(n15701), .ZN(n15703) );
  AOI21_X1 U19109 ( .B1(n15704), .B2(n19505), .A(n15703), .ZN(n15705) );
  OAI21_X1 U19110 ( .B1(n15706), .B2(n16671), .A(n15705), .ZN(P2_U2983) );
  INV_X1 U19111 ( .A(n15707), .ZN(n15709) );
  NOR2_X1 U19112 ( .A1(n15731), .A2(n15730), .ZN(n15729) );
  AOI21_X1 U19113 ( .B1(n15712), .B2(n15711), .A(n15710), .ZN(n15713) );
  XNOR2_X1 U19114 ( .A(n15714), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15715) );
  XNOR2_X1 U19115 ( .A(n15716), .B(n15715), .ZN(n15854) );
  AOI21_X1 U19116 ( .B1(n15738), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15719) );
  NOR2_X1 U19117 ( .A1(n15719), .A2(n15718), .ZN(n15853) );
  NOR2_X1 U19118 ( .A1(n19395), .A2(n15720), .ZN(n15847) );
  NOR2_X1 U19119 ( .A1(n19510), .A2(n15721), .ZN(n15722) );
  AOI211_X1 U19120 ( .C1(n19501), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15847), .B(n15722), .ZN(n15723) );
  OAI21_X1 U19121 ( .B1(n15850), .B2(n16655), .A(n15723), .ZN(n15724) );
  AOI21_X1 U19122 ( .B1(n15853), .B2(n19505), .A(n15724), .ZN(n15725) );
  OAI21_X1 U19123 ( .B1(n15854), .B2(n16671), .A(n15725), .ZN(P2_U2986) );
  XNOR2_X1 U19124 ( .A(n15738), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15865) );
  NAND2_X1 U19125 ( .A1(n19500), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15856) );
  OAI21_X1 U19126 ( .B1(n16677), .B2(n16504), .A(n15856), .ZN(n15727) );
  NOR2_X1 U19127 ( .A1(n16509), .A2(n16655), .ZN(n15726) );
  AOI211_X1 U19128 ( .C1(n16667), .C2(n15728), .A(n15727), .B(n15726), .ZN(
        n15733) );
  INV_X1 U19129 ( .A(n15729), .ZN(n15862) );
  NAND2_X1 U19130 ( .A1(n15731), .A2(n15730), .ZN(n15861) );
  NAND3_X1 U19131 ( .A1(n15862), .A2(n10923), .A3(n15861), .ZN(n15732) );
  OAI211_X1 U19132 ( .C1(n15865), .C2(n16668), .A(n15733), .B(n15732), .ZN(
        P2_U2987) );
  AOI21_X1 U19133 ( .B1(n15735), .B2(n15747), .A(n15746), .ZN(n15736) );
  XOR2_X1 U19134 ( .A(n15737), .B(n15736), .Z(n15876) );
  INV_X1 U19135 ( .A(n15751), .ZN(n15739) );
  AOI21_X1 U19136 ( .B1(n15872), .B2(n15739), .A(n15738), .ZN(n15874) );
  INV_X1 U19137 ( .A(n16526), .ZN(n15742) );
  INV_X1 U19138 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n15740) );
  OR2_X1 U19139 ( .A1(n19395), .A2(n20140), .ZN(n15867) );
  OAI21_X1 U19140 ( .B1(n16677), .B2(n15740), .A(n15867), .ZN(n15741) );
  AOI21_X1 U19141 ( .B1(n16667), .B2(n15742), .A(n15741), .ZN(n15743) );
  OAI21_X1 U19142 ( .B1(n16522), .B2(n16655), .A(n15743), .ZN(n15744) );
  AOI21_X1 U19143 ( .B1(n15874), .B2(n19505), .A(n15744), .ZN(n15745) );
  OAI21_X1 U19144 ( .B1(n16671), .B2(n15876), .A(n15745), .ZN(P2_U2988) );
  INV_X1 U19145 ( .A(n15746), .ZN(n15748) );
  NAND2_X1 U19146 ( .A1(n15748), .A2(n15747), .ZN(n15749) );
  XNOR2_X1 U19147 ( .A(n15735), .B(n15749), .ZN(n15888) );
  AOI21_X1 U19148 ( .B1(n15884), .B2(n15750), .A(n15751), .ZN(n15877) );
  NAND2_X1 U19149 ( .A1(n15877), .A2(n19505), .ZN(n15756) );
  NAND2_X1 U19150 ( .A1(n16667), .A2(n15752), .ZN(n15753) );
  NAND2_X1 U19151 ( .A1(n19500), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15880) );
  OAI211_X1 U19152 ( .C1(n16677), .C2(n16533), .A(n15753), .B(n15880), .ZN(
        n15754) );
  AOI21_X1 U19153 ( .B1(n16537), .B2(n19504), .A(n15754), .ZN(n15755) );
  OAI211_X1 U19154 ( .C1(n15888), .C2(n16671), .A(n15756), .B(n15755), .ZN(
        P2_U2989) );
  INV_X1 U19155 ( .A(n15767), .ZN(n15757) );
  OAI21_X1 U19156 ( .B1(n15757), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15750), .ZN(n15900) );
  NAND2_X1 U19157 ( .A1(n9915), .A2(n15760), .ZN(n15761) );
  XNOR2_X1 U19158 ( .A(n15758), .B(n15761), .ZN(n15898) );
  NOR2_X1 U19159 ( .A1(n19395), .A2(n20136), .ZN(n15891) );
  NOR2_X1 U19160 ( .A1(n19510), .A2(n16554), .ZN(n15762) );
  AOI211_X1 U19161 ( .C1(n19501), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15891), .B(n15762), .ZN(n15763) );
  OAI21_X1 U19162 ( .B1(n16549), .B2(n16655), .A(n15763), .ZN(n15764) );
  AOI21_X1 U19163 ( .B1(n15898), .B2(n10923), .A(n15764), .ZN(n15765) );
  OAI21_X1 U19164 ( .B1(n15900), .B2(n16668), .A(n15765), .ZN(P2_U2990) );
  OAI21_X1 U19165 ( .B1(n15766), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15767), .ZN(n15913) );
  NAND2_X1 U19166 ( .A1(n16667), .A2(n15768), .ZN(n15769) );
  NAND2_X1 U19167 ( .A1(n19500), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15901) );
  OAI211_X1 U19168 ( .C1(n16677), .C2(n9812), .A(n15769), .B(n15901), .ZN(
        n15770) );
  AOI21_X1 U19169 ( .B1(n16563), .B2(n19504), .A(n15770), .ZN(n15774) );
  OR2_X1 U19170 ( .A1(n15772), .A2(n15771), .ZN(n15910) );
  NAND3_X1 U19171 ( .A1(n15910), .A2(n15909), .A3(n10923), .ZN(n15773) );
  OAI211_X1 U19172 ( .C1(n15913), .C2(n16668), .A(n15774), .B(n15773), .ZN(
        P2_U2991) );
  INV_X1 U19173 ( .A(n15777), .ZN(n15779) );
  NOR2_X1 U19174 ( .A1(n15779), .A2(n15778), .ZN(n15780) );
  XNOR2_X1 U19175 ( .A(n15781), .B(n15780), .ZN(n15939) );
  INV_X1 U19176 ( .A(n15782), .ZN(n15803) );
  AOI21_X1 U19177 ( .B1(n15803), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15784) );
  NOR2_X1 U19178 ( .A1(n15784), .A2(n15783), .ZN(n15936) );
  NAND2_X1 U19179 ( .A1(n19250), .A2(n19504), .ZN(n15786) );
  NOR2_X1 U19180 ( .A1(n19395), .A2(n20129), .ZN(n15930) );
  AOI21_X1 U19181 ( .B1(n19501), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15930), .ZN(n15785) );
  OAI211_X1 U19182 ( .C1(n19260), .C2(n19510), .A(n15786), .B(n15785), .ZN(
        n15787) );
  AOI21_X1 U19183 ( .B1(n15936), .B2(n19505), .A(n15787), .ZN(n15788) );
  OAI21_X1 U19184 ( .B1(n15939), .B2(n16671), .A(n15788), .ZN(P2_U2994) );
  NAND2_X1 U19185 ( .A1(n15789), .A2(n15800), .ZN(n15793) );
  NAND2_X1 U19186 ( .A1(n15791), .A2(n15790), .ZN(n15792) );
  XNOR2_X1 U19187 ( .A(n15793), .B(n15792), .ZN(n15949) );
  XNOR2_X1 U19188 ( .A(n15782), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15947) );
  NOR2_X1 U19189 ( .A1(n19395), .A2(n20127), .ZN(n15942) );
  NOR2_X1 U19190 ( .A1(n16677), .A2(n15794), .ZN(n15795) );
  AOI211_X1 U19191 ( .C1(n19267), .C2(n16667), .A(n15942), .B(n15795), .ZN(
        n15796) );
  OAI21_X1 U19192 ( .B1(n16655), .B2(n15940), .A(n15796), .ZN(n15797) );
  AOI21_X1 U19193 ( .B1(n15947), .B2(n19505), .A(n15797), .ZN(n15798) );
  OAI21_X1 U19194 ( .B1(n15949), .B2(n16671), .A(n15798), .ZN(P2_U2995) );
  NAND2_X1 U19195 ( .A1(n15801), .A2(n15800), .ZN(n15802) );
  XNOR2_X1 U19196 ( .A(n15799), .B(n15802), .ZN(n15961) );
  AOI21_X1 U19197 ( .B1(n15963), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15804) );
  NOR2_X1 U19198 ( .A1(n15804), .A2(n15803), .ZN(n15959) );
  NOR2_X1 U19199 ( .A1(n19395), .A2(n20125), .ZN(n15951) );
  NOR2_X1 U19200 ( .A1(n19275), .A2(n19510), .ZN(n15805) );
  AOI211_X1 U19201 ( .C1(n19501), .C2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15951), .B(n15805), .ZN(n15806) );
  OAI21_X1 U19202 ( .B1(n16655), .B2(n19282), .A(n15806), .ZN(n15807) );
  AOI21_X1 U19203 ( .B1(n15959), .B2(n19505), .A(n15807), .ZN(n15808) );
  OAI21_X1 U19204 ( .B1(n15961), .B2(n16671), .A(n15808), .ZN(P2_U2996) );
  XNOR2_X1 U19205 ( .A(n15963), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15817) );
  OAI21_X1 U19206 ( .B1(n15809), .B2(n15811), .A(n15810), .ZN(n15962) );
  NAND2_X1 U19207 ( .A1(n15962), .A2(n10923), .ZN(n15816) );
  NAND2_X1 U19208 ( .A1(n19290), .A2(n16667), .ZN(n15812) );
  NAND2_X1 U19209 ( .A1(n19500), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15973) );
  OAI211_X1 U19210 ( .C1(n16677), .C2(n15813), .A(n15812), .B(n15973), .ZN(
        n15814) );
  AOI21_X1 U19211 ( .B1(n19504), .B2(n19296), .A(n15814), .ZN(n15815) );
  OAI211_X1 U19212 ( .C1(n16668), .C2(n15817), .A(n15816), .B(n15815), .ZN(
        P2_U2997) );
  XNOR2_X1 U19213 ( .A(n15996), .B(n15985), .ZN(n15826) );
  AND2_X1 U19214 ( .A1(n15820), .A2(n15819), .ZN(n15821) );
  NOR2_X1 U19215 ( .A1(n15818), .A2(n15821), .ZN(n15982) );
  NAND2_X1 U19216 ( .A1(n15982), .A2(n10923), .ZN(n15825) );
  INV_X1 U19217 ( .A(n15978), .ZN(n19309) );
  NOR2_X1 U19218 ( .A1(n15977), .A2(n19395), .ZN(n15823) );
  OAI22_X1 U19219 ( .A1(n16677), .A2(n9809), .B1(n19510), .B2(n19302), .ZN(
        n15822) );
  AOI211_X1 U19220 ( .C1(n19504), .C2(n19309), .A(n15823), .B(n15822), .ZN(
        n15824) );
  OAI211_X1 U19221 ( .C1(n16668), .C2(n15826), .A(n15825), .B(n15824), .ZN(
        P2_U2998) );
  NAND2_X1 U19222 ( .A1(n16647), .A2(n16645), .ZN(n15829) );
  NAND2_X1 U19223 ( .A1(n15827), .A2(n15828), .ZN(n16646) );
  XOR2_X1 U19224 ( .A(n15829), .B(n16646), .Z(n16077) );
  NAND2_X1 U19225 ( .A1(n15830), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15832) );
  NAND2_X1 U19226 ( .A1(n15832), .A2(n15831), .ZN(n16639) );
  XOR2_X1 U19227 ( .A(n16638), .B(n16639), .Z(n16075) );
  OAI22_X1 U19228 ( .A1(n16677), .A2(n19396), .B1(n20111), .B2(n19395), .ZN(
        n15833) );
  AOI21_X1 U19229 ( .B1(n16667), .B2(n19394), .A(n15833), .ZN(n15834) );
  OAI21_X1 U19230 ( .B1(n16655), .B2(n19405), .A(n15834), .ZN(n15835) );
  AOI21_X1 U19231 ( .B1(n16075), .B2(n19505), .A(n15835), .ZN(n15836) );
  OAI21_X1 U19232 ( .B1(n16077), .B2(n16671), .A(n15836), .ZN(P2_U3007) );
  INV_X1 U19233 ( .A(n15837), .ZN(n15838) );
  NAND2_X1 U19234 ( .A1(n15838), .A2(n16700), .ZN(n15845) );
  INV_X1 U19235 ( .A(n15839), .ZN(n15860) );
  AOI211_X1 U19236 ( .C1(n15843), .C2(n15842), .A(n15841), .B(n15857), .ZN(
        n15844) );
  XNOR2_X1 U19237 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15852) );
  OAI21_X1 U19238 ( .B1(n15850), .B2(n16716), .A(n15849), .ZN(n15851) );
  NAND2_X1 U19239 ( .A1(n16710), .A2(n16507), .ZN(n15855) );
  OAI211_X1 U19240 ( .C1(n16509), .C2(n16716), .A(n15856), .B(n15855), .ZN(
        n15859) );
  NOR2_X1 U19241 ( .A1(n15857), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15858) );
  AOI211_X1 U19242 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15860), .A(
        n15859), .B(n15858), .ZN(n15864) );
  NAND3_X1 U19243 ( .A1(n15862), .A2(n16721), .A3(n15861), .ZN(n15863) );
  OAI211_X1 U19244 ( .C1(n15865), .C2(n16717), .A(n15864), .B(n15863), .ZN(
        P2_U3019) );
  OAI211_X1 U19245 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n15885), .B(n15866), .ZN(
        n15871) );
  INV_X1 U19246 ( .A(n16522), .ZN(n15869) );
  OAI21_X1 U19247 ( .B1(n16072), .B2(n16521), .A(n15867), .ZN(n15868) );
  AOI21_X1 U19248 ( .B1(n15869), .B2(n16699), .A(n15868), .ZN(n15870) );
  OAI211_X1 U19249 ( .C1(n15878), .C2(n15872), .A(n15871), .B(n15870), .ZN(
        n15873) );
  AOI21_X1 U19250 ( .B1(n15874), .B2(n16700), .A(n15873), .ZN(n15875) );
  OAI21_X1 U19251 ( .B1(n16704), .B2(n15876), .A(n15875), .ZN(P2_U3020) );
  NAND2_X1 U19252 ( .A1(n15877), .A2(n16700), .ZN(n15887) );
  NOR2_X1 U19253 ( .A1(n15878), .A2(n15884), .ZN(n15883) );
  NAND2_X1 U19254 ( .A1(n16710), .A2(n16536), .ZN(n15879) );
  OAI211_X1 U19255 ( .C1(n15881), .C2(n16716), .A(n15880), .B(n15879), .ZN(
        n15882) );
  AOI211_X1 U19256 ( .C1(n15885), .C2(n15884), .A(n15883), .B(n15882), .ZN(
        n15886) );
  OAI211_X1 U19257 ( .C1(n15888), .C2(n16704), .A(n15887), .B(n15886), .ZN(
        P2_U3021) );
  INV_X1 U19258 ( .A(n15889), .ZN(n15896) );
  NAND3_X1 U19259 ( .A1(n15903), .A2(n15904), .A3(n15895), .ZN(n15894) );
  INV_X1 U19260 ( .A(n16549), .ZN(n15892) );
  NOR2_X1 U19261 ( .A1(n16072), .A2(n16557), .ZN(n15890) );
  AOI211_X1 U19262 ( .C1(n15892), .C2(n16699), .A(n15891), .B(n15890), .ZN(
        n15893) );
  OAI211_X1 U19263 ( .C1(n15896), .C2(n15895), .A(n15894), .B(n15893), .ZN(
        n15897) );
  AOI21_X1 U19264 ( .B1(n15898), .B2(n16721), .A(n15897), .ZN(n15899) );
  OAI21_X1 U19265 ( .B1(n15900), .B2(n16717), .A(n15899), .ZN(P2_U3022) );
  NAND2_X1 U19266 ( .A1(n16563), .A2(n16699), .ZN(n15902) );
  OAI211_X1 U19267 ( .C1(n16072), .C2(n16561), .A(n15902), .B(n15901), .ZN(
        n15908) );
  INV_X1 U19268 ( .A(n15903), .ZN(n15925) );
  AOI211_X1 U19269 ( .C1(n15906), .C2(n15905), .A(n15904), .B(n15925), .ZN(
        n15907) );
  AOI211_X1 U19270 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n15923), .A(
        n15908), .B(n15907), .ZN(n15912) );
  NAND3_X1 U19271 ( .A1(n15910), .A2(n15909), .A3(n16721), .ZN(n15911) );
  OAI211_X1 U19272 ( .C1(n15913), .C2(n16717), .A(n15912), .B(n15911), .ZN(
        P2_U3023) );
  OAI21_X1 U19273 ( .B1(n13229), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15914), .ZN(n16579) );
  NAND2_X1 U19274 ( .A1(n15917), .A2(n15916), .ZN(n15918) );
  XNOR2_X1 U19275 ( .A(n9687), .B(n15918), .ZN(n16582) );
  NAND2_X1 U19276 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19500), .ZN(n15921) );
  NAND2_X1 U19277 ( .A1(n16710), .A2(n15919), .ZN(n15920) );
  OAI211_X1 U19278 ( .C1(n16578), .C2(n16716), .A(n15921), .B(n15920), .ZN(
        n15922) );
  AOI21_X1 U19279 ( .B1(n15923), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15922), .ZN(n15924) );
  OAI21_X1 U19280 ( .B1(n15925), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15924), .ZN(n15926) );
  AOI21_X1 U19281 ( .B1(n16582), .B2(n16721), .A(n15926), .ZN(n15927) );
  OAI21_X1 U19282 ( .B1(n16579), .B2(n16717), .A(n15927), .ZN(P2_U3024) );
  AOI211_X1 U19283 ( .C1(n15932), .C2(n15929), .A(n15928), .B(n15944), .ZN(
        n15935) );
  INV_X1 U19284 ( .A(n15952), .ZN(n15933) );
  AOI21_X1 U19285 ( .B1(n19250), .B2(n16699), .A(n15930), .ZN(n15931) );
  OAI21_X1 U19286 ( .B1(n15933), .B2(n15932), .A(n15931), .ZN(n15934) );
  AOI211_X1 U19287 ( .C1(n9778), .C2(n16710), .A(n15935), .B(n15934), .ZN(
        n15938) );
  NAND2_X1 U19288 ( .A1(n15936), .A2(n16700), .ZN(n15937) );
  OAI211_X1 U19289 ( .C1(n15939), .C2(n16704), .A(n15938), .B(n15937), .ZN(
        P2_U3026) );
  NOR2_X1 U19290 ( .A1(n19273), .A2(n16072), .ZN(n15946) );
  NOR2_X1 U19291 ( .A1(n15940), .A2(n16716), .ZN(n15941) );
  AOI211_X1 U19292 ( .C1(n15952), .C2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15942), .B(n15941), .ZN(n15943) );
  OAI21_X1 U19293 ( .B1(n15944), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15943), .ZN(n15945) );
  AOI211_X1 U19294 ( .C1(n15947), .C2(n16700), .A(n15946), .B(n15945), .ZN(
        n15948) );
  OAI21_X1 U19295 ( .B1(n15949), .B2(n16704), .A(n15948), .ZN(P2_U3027) );
  NOR2_X1 U19296 ( .A1(n19282), .A2(n16716), .ZN(n15950) );
  AOI211_X1 U19297 ( .C1(n15952), .C2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15951), .B(n15950), .ZN(n15956) );
  INV_X1 U19298 ( .A(n15995), .ZN(n15969) );
  NAND4_X1 U19299 ( .A1(n15969), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15954), .A4(n15953), .ZN(n15955) );
  OAI211_X1 U19300 ( .C1(n15957), .C2(n16072), .A(n15956), .B(n15955), .ZN(
        n15958) );
  AOI21_X1 U19301 ( .B1(n15959), .B2(n16700), .A(n15958), .ZN(n15960) );
  OAI21_X1 U19302 ( .B1(n15961), .B2(n16704), .A(n15960), .ZN(P2_U3028) );
  INV_X1 U19303 ( .A(n15962), .ZN(n15976) );
  AOI21_X1 U19304 ( .B1(n16717), .B2(n15964), .A(n15963), .ZN(n15965) );
  INV_X1 U19305 ( .A(n15996), .ZN(n15970) );
  AOI22_X1 U19306 ( .A1(n15970), .A2(n16700), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15969), .ZN(n15979) );
  NOR3_X1 U19307 ( .A1(n15979), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15985), .ZN(n15975) );
  XNOR2_X1 U19308 ( .A(n14433), .B(n15971), .ZN(n16573) );
  NAND2_X1 U19309 ( .A1(n19296), .A2(n16699), .ZN(n15972) );
  OAI211_X1 U19310 ( .C1(n16573), .C2(n16072), .A(n15973), .B(n15972), .ZN(
        n15974) );
  OAI22_X1 U19311 ( .A1(n16716), .A2(n15978), .B1(n15977), .B2(n19341), .ZN(
        n15981) );
  NOR2_X1 U19312 ( .A1(n15979), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15980) );
  AOI211_X1 U19313 ( .C1(n16710), .C2(n19310), .A(n15981), .B(n15980), .ZN(
        n15984) );
  NAND2_X1 U19314 ( .A1(n15982), .A2(n16721), .ZN(n15983) );
  OAI211_X1 U19315 ( .C1(n15986), .C2(n15985), .A(n15984), .B(n15983), .ZN(
        P2_U3030) );
  NAND2_X1 U19316 ( .A1(n15988), .A2(n15987), .ZN(n15990) );
  XOR2_X1 U19317 ( .A(n15990), .B(n15989), .Z(n16587) );
  INV_X1 U19318 ( .A(n19326), .ZN(n16000) );
  INV_X1 U19319 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n20120) );
  NOR2_X1 U19320 ( .A1(n20120), .A2(n19395), .ZN(n15991) );
  AOI21_X1 U19321 ( .B1(n16699), .B2(n19322), .A(n15991), .ZN(n15994) );
  NAND2_X1 U19322 ( .A1(n15992), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15993) );
  OAI211_X1 U19323 ( .C1(n15995), .C2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15994), .B(n15993), .ZN(n15999) );
  OAI21_X1 U19324 ( .B1(n15997), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15996), .ZN(n16586) );
  NOR2_X1 U19325 ( .A1(n16586), .A2(n16717), .ZN(n15998) );
  AOI211_X1 U19326 ( .C1(n16710), .C2(n16000), .A(n15999), .B(n15998), .ZN(
        n16001) );
  OAI21_X1 U19327 ( .B1(n16587), .B2(n16704), .A(n16001), .ZN(P2_U3031) );
  INV_X1 U19328 ( .A(n16004), .ZN(n16008) );
  NAND2_X1 U19329 ( .A1(n16003), .A2(n16008), .ZN(n16602) );
  NAND2_X1 U19330 ( .A1(n16602), .A2(n16007), .ZN(n16006) );
  NAND2_X1 U19331 ( .A1(n16006), .A2(n16005), .ZN(n16595) );
  INV_X1 U19332 ( .A(n16680), .ZN(n16029) );
  OAI21_X1 U19333 ( .B1(n16029), .B2(n16008), .A(n16028), .ZN(n16679) );
  INV_X1 U19334 ( .A(n19332), .ZN(n16012) );
  NAND3_X1 U19335 ( .A1(n16680), .A2(n16008), .A3(n16007), .ZN(n16011) );
  AOI21_X1 U19336 ( .B1(n16009), .B2(n14158), .A(n14353), .ZN(n19454) );
  AOI22_X1 U19337 ( .A1(n16710), .A2(n19454), .B1(n19500), .B2(
        P2_REIP_REG_14__SCAN_IN), .ZN(n16010) );
  OAI211_X1 U19338 ( .C1(n16012), .C2(n16716), .A(n16011), .B(n16010), .ZN(
        n16013) );
  AOI21_X1 U19339 ( .B1(n16679), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n16013), .ZN(n16019) );
  AND2_X1 U19340 ( .A1(n16016), .A2(n16015), .ZN(n16017) );
  XNOR2_X1 U19341 ( .A(n16014), .B(n16017), .ZN(n16592) );
  NAND2_X1 U19342 ( .A1(n16592), .A2(n16721), .ZN(n16018) );
  OAI211_X1 U19343 ( .C1(n16595), .C2(n16717), .A(n16019), .B(n16018), .ZN(
        P2_U3032) );
  XNOR2_X1 U19344 ( .A(n16003), .B(n16020), .ZN(n16611) );
  NAND2_X1 U19345 ( .A1(n16611), .A2(n16700), .ZN(n16034) );
  AOI21_X1 U19346 ( .B1(n16021), .B2(n13925), .A(n14157), .ZN(n19458) );
  AOI22_X1 U19347 ( .A1(n16699), .A2(n10090), .B1(n16710), .B2(n19458), .ZN(
        n16033) );
  INV_X1 U19348 ( .A(n16023), .ZN(n16025) );
  NOR2_X1 U19349 ( .A1(n16025), .A2(n16024), .ZN(n16026) );
  XNOR2_X1 U19350 ( .A(n16022), .B(n16026), .ZN(n16610) );
  NAND2_X1 U19351 ( .A1(n16610), .A2(n16721), .ZN(n16032) );
  NAND2_X1 U19352 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19500), .ZN(n16027) );
  OAI221_X1 U19353 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16029), 
        .C1(n16020), .C2(n16028), .A(n16027), .ZN(n16030) );
  INV_X1 U19354 ( .A(n16030), .ZN(n16031) );
  NAND4_X1 U19355 ( .A1(n16034), .A2(n16033), .A3(n16032), .A4(n16031), .ZN(
        P2_U3034) );
  INV_X1 U19356 ( .A(n16035), .ZN(n16627) );
  INV_X1 U19357 ( .A(n16003), .ZN(n16036) );
  OAI21_X1 U19358 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16627), .A(
        n16036), .ZN(n16615) );
  XNOR2_X1 U19359 ( .A(n16038), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n16039) );
  XNOR2_X1 U19360 ( .A(n9702), .B(n16039), .ZN(n16614) );
  NOR2_X1 U19361 ( .A1(n11523), .A2(n19395), .ZN(n16044) );
  INV_X1 U19362 ( .A(n16040), .ZN(n16041) );
  AOI211_X1 U19363 ( .C1(n16694), .C2(n16042), .A(n16041), .B(n16695), .ZN(
        n16043) );
  AOI211_X1 U19364 ( .C1(n16045), .C2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n16044), .B(n16043), .ZN(n16048) );
  INV_X1 U19365 ( .A(n19378), .ZN(n16046) );
  AOI22_X1 U19366 ( .A1(n16699), .A2(n19374), .B1(n16710), .B2(n16046), .ZN(
        n16047) );
  OAI211_X1 U19367 ( .C1(n16614), .C2(n16704), .A(n16048), .B(n16047), .ZN(
        n16049) );
  INV_X1 U19368 ( .A(n16049), .ZN(n16050) );
  OAI21_X1 U19369 ( .B1(n16615), .B2(n16717), .A(n16050), .ZN(P2_U3035) );
  AND2_X1 U19370 ( .A1(n16053), .A2(n16051), .ZN(n16054) );
  NAND2_X1 U19371 ( .A1(n16053), .A2(n16052), .ZN(n16628) );
  OAI21_X1 U19372 ( .B1(n16054), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n16628), .ZN(n16634) );
  INV_X1 U19373 ( .A(n16055), .ZN(n19387) );
  INV_X1 U19374 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n16056) );
  OAI22_X1 U19375 ( .A1(n16072), .A2(n19391), .B1(n19395), .B2(n16056), .ZN(
        n16061) );
  NOR2_X1 U19376 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16057), .ZN(
        n16059) );
  NOR2_X1 U19377 ( .A1(n16059), .A2(n16058), .ZN(n16060) );
  AOI211_X1 U19378 ( .C1(n16699), .C2(n19387), .A(n16061), .B(n16060), .ZN(
        n16069) );
  INV_X1 U19379 ( .A(n16062), .ZN(n16064) );
  OAI21_X1 U19380 ( .B1(n16646), .B2(n16064), .A(n16063), .ZN(n16067) );
  NAND2_X1 U19381 ( .A1(n16621), .A2(n16065), .ZN(n16066) );
  XNOR2_X1 U19382 ( .A(n16067), .B(n16066), .ZN(n16633) );
  OR2_X1 U19383 ( .A1(n16633), .A2(n16704), .ZN(n16068) );
  OAI211_X1 U19384 ( .C1(n16634), .C2(n16717), .A(n16069), .B(n16068), .ZN(
        P2_U3037) );
  NAND2_X1 U19385 ( .A1(n16070), .A2(n16082), .ZN(n16706) );
  NAND2_X1 U19386 ( .A1(P2_REIP_REG_7__SCAN_IN), .A2(n19500), .ZN(n16071) );
  OAI221_X1 U19387 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16706), .C1(
        n16708), .C2(n16724), .A(n16071), .ZN(n16074) );
  OAI22_X1 U19388 ( .A1(n19406), .A2(n16072), .B1(n16716), .B2(n19405), .ZN(
        n16073) );
  AOI211_X1 U19389 ( .C1(n16075), .C2(n16700), .A(n16074), .B(n16073), .ZN(
        n16076) );
  OAI21_X1 U19390 ( .B1(n16077), .B2(n16704), .A(n16076), .ZN(P2_U3039) );
  XOR2_X1 U19391 ( .A(n16079), .B(n16078), .Z(n19502) );
  NAND2_X1 U19392 ( .A1(n19502), .A2(n16721), .ZN(n16090) );
  NOR2_X1 U19393 ( .A1(n14221), .A2(n19395), .ZN(n16080) );
  AOI221_X1 U19394 ( .B1(n16082), .B2(n10595), .C1(n16081), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n16080), .ZN(n16089) );
  AOI22_X1 U19395 ( .A1(n19503), .A2(n16699), .B1(n16710), .B2(n16083), .ZN(
        n16088) );
  XNOR2_X1 U19396 ( .A(n16084), .B(n10595), .ZN(n16085) );
  XNOR2_X1 U19397 ( .A(n16086), .B(n16085), .ZN(n19506) );
  NAND2_X1 U19398 ( .A1(n19506), .A2(n16700), .ZN(n16087) );
  NAND4_X1 U19399 ( .A1(n16090), .A2(n16089), .A3(n16088), .A4(n16087), .ZN(
        P2_U3042) );
  INV_X1 U19400 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n17365) );
  INV_X1 U19401 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17400) );
  INV_X1 U19402 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17396) );
  INV_X1 U19403 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n16186) );
  INV_X1 U19404 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17489) );
  INV_X1 U19405 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17121) );
  INV_X1 U19406 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17528) );
  NAND3_X1 U19407 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17543) );
  NOR4_X1 U19408 ( .A1(n17126), .A2(n17528), .A3(n17532), .A4(n17543), .ZN(
        n16095) );
  NAND4_X1 U19409 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17557), .A4(n16095), .ZN(n17507) );
  NAND2_X1 U19410 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17526), .ZN(n17486) );
  NAND2_X1 U19411 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17370), .ZN(n17369) );
  INV_X1 U19412 ( .A(n17275), .ZN(n17270) );
  NAND2_X1 U19413 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n17270), .ZN(n16174) );
  AND2_X1 U19414 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17269) );
  NAND2_X1 U19415 ( .A1(n18548), .A2(n9732), .ZN(n17559) );
  INV_X2 U19416 ( .A(n17555), .ZN(n17551) );
  AOI22_X1 U19417 ( .A1(n17508), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17494), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n16097) );
  OAI21_X1 U19418 ( .B1(n10949), .B2(n17544), .A(n16097), .ZN(n16108) );
  INV_X1 U19419 ( .A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n18755) );
  AOI22_X1 U19420 ( .A1(n16175), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n16106) );
  AOI22_X1 U19421 ( .A1(n17512), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16098) );
  OAI21_X1 U19422 ( .B1(n10109), .B2(n16099), .A(n16098), .ZN(n16104) );
  AOI22_X1 U19423 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n16101) );
  AOI22_X1 U19424 ( .A1(n9671), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16100) );
  OAI211_X1 U19425 ( .C1(n10978), .C2(n16102), .A(n16101), .B(n16100), .ZN(
        n16103) );
  AOI211_X1 U19426 ( .C1(n11129), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n16104), .B(n16103), .ZN(n16105) );
  OAI211_X1 U19427 ( .C1(n17472), .C2(n18755), .A(n16106), .B(n16105), .ZN(
        n16107) );
  AOI211_X1 U19428 ( .C1(n17421), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n16108), .B(n16107), .ZN(n17277) );
  AOI22_X1 U19429 ( .A1(n17508), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16109) );
  OAI21_X1 U19430 ( .B1(n10109), .B2(n17372), .A(n16109), .ZN(n16120) );
  AOI22_X1 U19431 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16117) );
  AOI22_X1 U19432 ( .A1(n17494), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n16110) );
  OAI21_X1 U19433 ( .B1(n17472), .B2(n18749), .A(n16110), .ZN(n16115) );
  AOI22_X1 U19434 ( .A1(n16175), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9671), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n16113) );
  AOI22_X1 U19435 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n16112) );
  OAI211_X1 U19436 ( .C1(n17460), .C2(n18579), .A(n16113), .B(n16112), .ZN(
        n16114) );
  AOI211_X1 U19437 ( .C1(n17514), .C2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n16115), .B(n16114), .ZN(n16116) );
  OAI211_X1 U19438 ( .C1(n16118), .C2(n17492), .A(n16117), .B(n16116), .ZN(
        n16119) );
  AOI211_X1 U19439 ( .C1(n17421), .C2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A(
        n16120), .B(n16119), .ZN(n17287) );
  AOI22_X1 U19440 ( .A1(n17403), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17514), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16130) );
  AOI22_X1 U19441 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17495), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16122) );
  AOI22_X1 U19442 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16121) );
  OAI211_X1 U19443 ( .C1(n17460), .C2(n18576), .A(n16122), .B(n16121), .ZN(
        n16128) );
  AOI22_X1 U19444 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n16175), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n16126) );
  AOI22_X1 U19445 ( .A1(n9670), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16125) );
  AOI22_X1 U19446 ( .A1(n17508), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n16124) );
  NAND2_X1 U19447 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n16123) );
  NAND4_X1 U19448 ( .A1(n16126), .A2(n16125), .A3(n16124), .A4(n16123), .ZN(
        n16127) );
  AOI211_X1 U19449 ( .C1(n11129), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n16128), .B(n16127), .ZN(n16129) );
  OAI211_X1 U19450 ( .C1(n11006), .C2(n16131), .A(n16130), .B(n16129), .ZN(
        n17292) );
  AOI22_X1 U19451 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17512), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16141) );
  AOI22_X1 U19452 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n16175), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16133) );
  AOI22_X1 U19453 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17508), .ZN(n16132) );
  OAI211_X1 U19454 ( .C1(n10978), .C2(n17412), .A(n16133), .B(n16132), .ZN(
        n16139) );
  AOI22_X1 U19455 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n17476), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n9670), .ZN(n16137) );
  AOI22_X1 U19456 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17520), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n17494), .ZN(n16136) );
  AOI22_X1 U19457 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n17490), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16135) );
  NAND2_X1 U19458 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17339), .ZN(
        n16134) );
  NAND4_X1 U19459 ( .A1(n16137), .A2(n16136), .A3(n16135), .A4(n16134), .ZN(
        n16138) );
  AOI211_X1 U19460 ( .C1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .C2(n11129), .A(
        n16139), .B(n16138), .ZN(n16140) );
  OAI211_X1 U19461 ( .C1(n17474), .C2(n17529), .A(n16141), .B(n16140), .ZN(
        n17293) );
  NAND2_X1 U19462 ( .A1(n17292), .A2(n17293), .ZN(n17291) );
  NOR2_X1 U19463 ( .A1(n17287), .A2(n17291), .ZN(n17284) );
  AOI22_X1 U19464 ( .A1(n17512), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9671), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16151) );
  AOI22_X1 U19465 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n16143) );
  AOI22_X1 U19466 ( .A1(n11030), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16142) );
  OAI211_X1 U19467 ( .C1(n10978), .C2(n17353), .A(n16143), .B(n16142), .ZN(
        n16149) );
  AOI22_X1 U19468 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n16175), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16147) );
  AOI22_X1 U19469 ( .A1(n17494), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16146) );
  AOI22_X1 U19470 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16145) );
  NAND2_X1 U19471 ( .A1(n17403), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n16144) );
  NAND4_X1 U19472 ( .A1(n16147), .A2(n16146), .A3(n16145), .A4(n16144), .ZN(
        n16148) );
  AOI211_X1 U19473 ( .C1(n11129), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n16149), .B(n16148), .ZN(n16150) );
  OAI211_X1 U19474 ( .C1(n17472), .C2(n18752), .A(n16151), .B(n16150), .ZN(
        n17283) );
  NAND2_X1 U19475 ( .A1(n17284), .A2(n17283), .ZN(n17282) );
  NOR2_X1 U19476 ( .A1(n17277), .A2(n17282), .ZN(n17276) );
  AOI22_X1 U19477 ( .A1(n16175), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16162) );
  AOI22_X1 U19478 ( .A1(n17494), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n16161) );
  AOI22_X1 U19479 ( .A1(n17512), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16160) );
  OAI22_X1 U19480 ( .A1(n10109), .A2(n16152), .B1(n10978), .B2(n17332), .ZN(
        n16158) );
  AOI22_X1 U19481 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16156) );
  AOI22_X1 U19482 ( .A1(n17508), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9670), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16155) );
  AOI22_X1 U19483 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17495), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16154) );
  NAND2_X1 U19484 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n16153) );
  NAND4_X1 U19485 ( .A1(n16156), .A2(n16155), .A3(n16154), .A4(n16153), .ZN(
        n16157) );
  AOI211_X1 U19486 ( .C1(n17339), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n16158), .B(n16157), .ZN(n16159) );
  NAND4_X1 U19487 ( .A1(n16162), .A2(n16161), .A3(n16160), .A4(n16159), .ZN(
        n17273) );
  NAND2_X1 U19488 ( .A1(n17276), .A2(n17273), .ZN(n17272) );
  INV_X1 U19489 ( .A(n17272), .ZN(n17263) );
  AOI22_X1 U19490 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16172) );
  AOI22_X1 U19491 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17495), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16164) );
  AOI22_X1 U19492 ( .A1(n16175), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n16163) );
  OAI211_X1 U19493 ( .C1(n17460), .C2(n18589), .A(n16164), .B(n16163), .ZN(
        n16170) );
  AOI22_X1 U19494 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17508), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16168) );
  AOI22_X1 U19495 ( .A1(n17494), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9670), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16167) );
  AOI22_X1 U19496 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17403), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16166) );
  NAND2_X1 U19497 ( .A1(n17514), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n16165) );
  NAND4_X1 U19498 ( .A1(n16168), .A2(n16167), .A3(n16166), .A4(n16165), .ZN(
        n16169) );
  AOI211_X1 U19499 ( .C1(n11129), .C2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A(
        n16170), .B(n16169), .ZN(n16171) );
  OAI211_X1 U19500 ( .C1(n17472), .C2(n18761), .A(n16172), .B(n16171), .ZN(
        n17264) );
  XOR2_X1 U19501 ( .A(n17263), .B(n17264), .Z(n17577) );
  AOI22_X1 U19502 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17267), .B1(n17555), 
        .B2(n17577), .ZN(n16173) );
  OAI21_X1 U19503 ( .B1(P3_EBX_REG_28__SCAN_IN), .B2(n16174), .A(n16173), .ZN(
        P3_U2675) );
  AOI22_X1 U19504 ( .A1(n10981), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17514), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16185) );
  AOI22_X1 U19505 ( .A1(n16175), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16177) );
  AOI22_X1 U19506 ( .A1(n11030), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9670), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16176) );
  OAI211_X1 U19507 ( .C1(n17460), .C2(n17537), .A(n16177), .B(n16176), .ZN(
        n16183) );
  AOI22_X1 U19508 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16181) );
  AOI22_X1 U19509 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16180) );
  AOI22_X1 U19510 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17494), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16179) );
  NAND2_X1 U19511 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n16178) );
  NAND4_X1 U19512 ( .A1(n16181), .A2(n16180), .A3(n16179), .A4(n16178), .ZN(
        n16182) );
  AOI211_X1 U19513 ( .C1(n11129), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n16183), .B(n16182), .ZN(n16184) );
  OAI211_X1 U19514 ( .C1(n10946), .C2(n18761), .A(n16185), .B(n16184), .ZN(
        n17663) );
  INV_X1 U19515 ( .A(n17663), .ZN(n16188) );
  NOR3_X1 U19516 ( .A1(n17691), .A2(n16186), .A3(n17467), .ZN(n17447) );
  NAND2_X1 U19517 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17447), .ZN(n17434) );
  OAI211_X1 U19518 ( .C1(n17447), .C2(P3_EBX_REG_13__SCAN_IN), .A(n17551), .B(
        n17434), .ZN(n16187) );
  OAI21_X1 U19519 ( .B1(n16188), .B2(n17551), .A(n16187), .ZN(P3_U2690) );
  NOR2_X1 U19520 ( .A1(n19010), .A2(n19015), .ZN(n18691) );
  INV_X1 U19521 ( .A(n18691), .ZN(n18512) );
  AOI221_X1 U19522 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18512), .C1(n16190), 
        .C2(n18512), .A(n16189), .ZN(n18510) );
  NOR2_X1 U19523 ( .A1(n16191), .A2(n19010), .ZN(n16192) );
  OAI21_X1 U19524 ( .B1(n16192), .B2(n18773), .A(n18511), .ZN(n18508) );
  AOI22_X1 U19525 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18510), .B1(
        n18508), .B2(n19015), .ZN(P3_U2865) );
  OAI22_X1 U19526 ( .A1(n16738), .A2(n18492), .B1(n16739), .B2(n18345), .ZN(
        n16261) );
  AOI211_X1 U19527 ( .C1(n18429), .C2(n16193), .A(n18489), .B(n16261), .ZN(
        n16194) );
  OAI21_X1 U19528 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18483), .A(
        n16194), .ZN(n16195) );
  AOI22_X1 U19529 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n16195), .B1(
        n18499), .B2(P3_REIP_REG_29__SCAN_IN), .ZN(n16203) );
  NAND2_X1 U19530 ( .A1(n16196), .A2(n18498), .ZN(n16197) );
  OAI211_X1 U19531 ( .C1(n18345), .C2(n16199), .A(n16198), .B(n16197), .ZN(
        n16259) );
  NAND3_X1 U19532 ( .A1(n16201), .A2(n16200), .A3(n16259), .ZN(n16202) );
  OAI211_X1 U19533 ( .C1(n16204), .C2(n18418), .A(n16203), .B(n16202), .ZN(
        P3_U2833) );
  OAI22_X1 U19534 ( .A1(n16578), .A2(n19422), .B1(n16205), .B2(n19447), .ZN(
        n16206) );
  INV_X1 U19535 ( .A(n16206), .ZN(n16216) );
  INV_X1 U19536 ( .A(n16207), .ZN(n16214) );
  AOI22_X1 U19537 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19437), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19431), .ZN(n16208) );
  OAI21_X1 U19538 ( .B1(n19413), .B2(n10729), .A(n16208), .ZN(n16213) );
  OAI211_X1 U19539 ( .C1(n16210), .C2(n16585), .A(n19443), .B(n16209), .ZN(
        n16211) );
  INV_X1 U19540 ( .A(n16211), .ZN(n16212) );
  AOI211_X1 U19541 ( .C1(n16214), .C2(n19403), .A(n16213), .B(n16212), .ZN(
        n16215) );
  NAND2_X1 U19542 ( .A1(n16216), .A2(n16215), .ZN(P2_U2833) );
  INV_X1 U19543 ( .A(n16226), .ZN(n16228) );
  AOI21_X1 U19544 ( .B1(n16217), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n20733), .ZN(n16218) );
  AND2_X1 U19545 ( .A1(n16219), .A2(n16218), .ZN(n16222) );
  OAI22_X1 U19546 ( .A1(n16221), .A2(n16220), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n16222), .ZN(n16224) );
  NAND2_X1 U19547 ( .A1(n16222), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n16223) );
  OAI211_X1 U19548 ( .C1(n16226), .C2(n16225), .A(n16224), .B(n16223), .ZN(
        n16227) );
  OAI21_X1 U19549 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16228), .A(
        n16227), .ZN(n16230) );
  AOI222_X1 U19550 ( .A1(n16230), .A2(n20768), .B1(n16230), .B2(n16229), .C1(
        n20768), .C2(n16229), .ZN(n16239) );
  INV_X1 U19551 ( .A(n16231), .ZN(n16236) );
  INV_X1 U19552 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n21106) );
  INV_X1 U19553 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n21212) );
  AOI21_X1 U19554 ( .B1(n21106), .B2(n21212), .A(n16232), .ZN(n16234) );
  NOR4_X1 U19555 ( .A1(n16236), .A2(n16235), .A3(n16234), .A4(n16233), .ZN(
        n16237) );
  OAI211_X1 U19556 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n16239), .A(
        n16238), .B(n16237), .ZN(n16247) );
  INV_X1 U19557 ( .A(n16240), .ZN(n16244) );
  NOR3_X1 U19558 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n12006), .A3(n21027), 
        .ZN(n16241) );
  NOR2_X1 U19559 ( .A1(n16248), .A2(n16241), .ZN(n16242) );
  AOI21_X1 U19560 ( .B1(n16244), .B2(n16243), .A(n16242), .ZN(n16463) );
  INV_X1 U19561 ( .A(n16463), .ZN(n16245) );
  AOI221_X1 U19562 ( .B1(n21023), .B2(n20942), .C1(n16247), .C2(n20942), .A(
        n16245), .ZN(n16249) );
  NOR2_X1 U19563 ( .A1(n16249), .A2(n21023), .ZN(n16468) );
  OAI21_X1 U19564 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21027), .A(n16468), 
        .ZN(n16466) );
  AOI211_X1 U19565 ( .C1(n16248), .C2(n16247), .A(n16246), .B(n16466), .ZN(
        n16254) );
  INV_X1 U19566 ( .A(n16249), .ZN(n16250) );
  OAI21_X1 U19567 ( .B1(n16251), .B2(n21022), .A(n16250), .ZN(n16252) );
  AOI22_X1 U19568 ( .A1(n16254), .A2(n16253), .B1(n21023), .B2(n16252), .ZN(
        P1_U3161) );
  NAND2_X1 U19569 ( .A1(n16256), .A2(n16255), .ZN(n16257) );
  XNOR2_X1 U19570 ( .A(n16257), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16744) );
  NOR2_X1 U19571 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16258), .ZN(
        n16740) );
  AOI22_X1 U19572 ( .A1(n18349), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n16740), 
        .B2(n16259), .ZN(n16264) );
  INV_X1 U19573 ( .A(n16260), .ZN(n16262) );
  OAI21_X1 U19574 ( .B1(n16262), .B2(n16261), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16263) );
  OAI211_X1 U19575 ( .C1(n16744), .C2(n18418), .A(n16264), .B(n16263), .ZN(
        P3_U2832) );
  INV_X1 U19576 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20960) );
  NAND2_X1 U19577 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20960), .ZN(n20955) );
  INV_X1 U19578 ( .A(HOLD), .ZN(n20946) );
  INV_X1 U19579 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21176) );
  NOR2_X1 U19580 ( .A1(n20954), .A2(n21176), .ZN(n20948) );
  AOI221_X1 U19581 ( .B1(n20960), .B2(n20948), .C1(n20946), .C2(n20948), .A(
        n16265), .ZN(n16267) );
  NAND2_X1 U19582 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21018), .ZN(n16266) );
  OAI211_X1 U19583 ( .C1(n20955), .C2(n20946), .A(n16267), .B(n16266), .ZN(
        P1_U3195) );
  AND2_X1 U19584 ( .A1(n16268), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  OAI221_X1 U19585 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n20226), .C1(n20218), 
        .C2(n20215), .A(n19942), .ZN(n20084) );
  NAND2_X1 U19586 ( .A1(n14795), .A2(n19942), .ZN(n19205) );
  AND3_X1 U19587 ( .A1(n20084), .A2(n19205), .A3(n16726), .ZN(P2_U3178) );
  OAI21_X1 U19588 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n20218), .ZN(n16269) );
  INV_X1 U19589 ( .A(n16269), .ZN(n20220) );
  NAND2_X1 U19590 ( .A1(n16270), .A2(n20220), .ZN(n16271) );
  AOI221_X1 U19591 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16272), .C1(n20208), .C2(
        n16272), .A(n20022), .ZN(n20203) );
  INV_X1 U19592 ( .A(n20203), .ZN(n20200) );
  NOR2_X1 U19593 ( .A1(n16273), .A2(n20200), .ZN(P2_U3047) );
  NOR3_X1 U19594 ( .A1(n16275), .A2(n17727), .A3(n9725), .ZN(n16276) );
  NAND2_X1 U19595 ( .A1(n18548), .A2(n17690), .ZN(n17653) );
  INV_X1 U19596 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17797) );
  NAND2_X1 U19597 ( .A1(n17691), .A2(n17690), .ZN(n17722) );
  AOI22_X1 U19598 ( .A1(n17719), .A2(BUF2_REG_0__SCAN_IN), .B1(n17718), .B2(
        n18175), .ZN(n16279) );
  OAI221_X1 U19599 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17653), .C1(n17797), 
        .C2(n17690), .A(n16279), .ZN(P3_U2735) );
  INV_X1 U19600 ( .A(n16280), .ZN(n16283) );
  AOI22_X1 U19601 ( .A1(n20321), .A2(P1_EBX_REG_18__SCAN_IN), .B1(n20338), 
        .B2(n16281), .ZN(n16282) );
  OAI21_X1 U19602 ( .B1(n16283), .B2(n20985), .A(n16282), .ZN(n16284) );
  AOI211_X1 U19603 ( .C1(n20323), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20310), .B(n16284), .ZN(n16289) );
  OAI22_X1 U19604 ( .A1(n16286), .A2(n16324), .B1(n16285), .B2(n20351), .ZN(
        n16287) );
  INV_X1 U19605 ( .A(n16287), .ZN(n16288) );
  OAI211_X1 U19606 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n16290), .A(n16289), 
        .B(n16288), .ZN(P1_U2822) );
  OAI22_X1 U19607 ( .A1(n16292), .A2(n20351), .B1(n16291), .B2(n20340), .ZN(
        n16293) );
  AOI211_X1 U19608 ( .C1(n20323), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20310), .B(n16293), .ZN(n16298) );
  INV_X1 U19609 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20981) );
  OAI21_X1 U19610 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n16294), .ZN(n16295) );
  OAI22_X1 U19611 ( .A1(n16316), .A2(n20981), .B1(n16302), .B2(n16295), .ZN(
        n16296) );
  AOI21_X1 U19612 ( .B1(n16349), .B2(n20287), .A(n16296), .ZN(n16297) );
  OAI211_X1 U19613 ( .C1(n16353), .C2(n20306), .A(n16298), .B(n16297), .ZN(
        P1_U2824) );
  INV_X1 U19614 ( .A(n16299), .ZN(n16387) );
  AOI22_X1 U19615 ( .A1(n16387), .A2(n20320), .B1(n20321), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n16300) );
  OAI211_X1 U19616 ( .C1(n20335), .C2(n16301), .A(n16300), .B(n20289), .ZN(
        n16305) );
  OAI22_X1 U19617 ( .A1(n16303), .A2(n16324), .B1(P1_REIP_REG_15__SCAN_IN), 
        .B2(n16302), .ZN(n16304) );
  AOI211_X1 U19618 ( .C1(n16306), .C2(n20338), .A(n16305), .B(n16304), .ZN(
        n16307) );
  OAI21_X1 U19619 ( .B1(n16316), .B2(n15253), .A(n16307), .ZN(P1_U2825) );
  NOR2_X1 U19620 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(n16308), .ZN(n16315) );
  AOI22_X1 U19621 ( .A1(n20321), .A2(P1_EBX_REG_14__SCAN_IN), .B1(n20338), 
        .B2(n16354), .ZN(n16314) );
  INV_X1 U19622 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16311) );
  NAND2_X1 U19623 ( .A1(n16309), .A2(n20320), .ZN(n16310) );
  OAI211_X1 U19624 ( .C1(n16311), .C2(n20335), .A(n16310), .B(n20289), .ZN(
        n16312) );
  AOI21_X1 U19625 ( .B1(n16356), .B2(n20287), .A(n16312), .ZN(n16313) );
  OAI211_X1 U19626 ( .C1(n16316), .C2(n16315), .A(n16314), .B(n16313), .ZN(
        P1_U2826) );
  INV_X1 U19627 ( .A(n16317), .ZN(n16318) );
  AOI22_X1 U19628 ( .A1(n20321), .A2(P1_EBX_REG_13__SCAN_IN), .B1(n20338), 
        .B2(n16318), .ZN(n16330) );
  NAND2_X1 U19629 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n16322) );
  NOR3_X1 U19630 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n16322), .A3(n16319), 
        .ZN(n16328) );
  OAI22_X1 U19631 ( .A1(n16321), .A2(n20335), .B1(n20351), .B2(n16320), .ZN(
        n16327) );
  AND2_X1 U19632 ( .A1(n20347), .A2(n16322), .ZN(n16323) );
  NOR2_X1 U19633 ( .A1(n16345), .A2(n16323), .ZN(n16340) );
  OAI22_X1 U19634 ( .A1(n16325), .A2(n16324), .B1(n16340), .B2(n20977), .ZN(
        n16326) );
  NOR4_X1 U19635 ( .A1(n20310), .A2(n16328), .A3(n16327), .A4(n16326), .ZN(
        n16329) );
  NAND2_X1 U19636 ( .A1(n16330), .A2(n16329), .ZN(P1_U2827) );
  AOI21_X1 U19637 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n16342), .A(
        P1_REIP_REG_12__SCAN_IN), .ZN(n16339) );
  INV_X1 U19638 ( .A(n16331), .ZN(n16332) );
  AOI22_X1 U19639 ( .A1(n20321), .A2(P1_EBX_REG_12__SCAN_IN), .B1(n20338), 
        .B2(n16332), .ZN(n16338) );
  OAI22_X1 U19640 ( .A1(n16334), .A2(n20335), .B1(n20351), .B2(n16333), .ZN(
        n16335) );
  AOI211_X1 U19641 ( .C1(n16336), .C2(n20287), .A(n20310), .B(n16335), .ZN(
        n16337) );
  OAI211_X1 U19642 ( .C1(n16340), .C2(n16339), .A(n16338), .B(n16337), .ZN(
        P1_U2828) );
  INV_X1 U19643 ( .A(n16367), .ZN(n16341) );
  AOI22_X1 U19644 ( .A1(n20321), .A2(P1_EBX_REG_11__SCAN_IN), .B1(n16341), 
        .B2(n20338), .ZN(n16348) );
  INV_X1 U19645 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20974) );
  AOI22_X1 U19646 ( .A1(n20974), .A2(n16342), .B1(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n20323), .ZN(n16343) );
  INV_X1 U19647 ( .A(n16343), .ZN(n16344) );
  AOI211_X1 U19648 ( .C1(n16396), .C2(n20320), .A(n20310), .B(n16344), .ZN(
        n16347) );
  AOI22_X1 U19649 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n16345), .B1(n20287), 
        .B2(n16363), .ZN(n16346) );
  NAND3_X1 U19650 ( .A1(n16348), .A2(n16347), .A3(n16346), .ZN(P1_U2829) );
  AOI22_X1 U19651 ( .A1(n20416), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n20473), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n16352) );
  AOI22_X1 U19652 ( .A1(n16350), .A2(n20422), .B1(n16364), .B2(n16349), .ZN(
        n16351) );
  OAI211_X1 U19653 ( .C1(n20427), .C2(n16353), .A(n16352), .B(n16351), .ZN(
        P1_U2983) );
  AOI22_X1 U19654 ( .A1(n20416), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20473), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16358) );
  AOI22_X1 U19655 ( .A1(n16356), .A2(n16364), .B1(n16355), .B2(n16354), .ZN(
        n16357) );
  OAI211_X1 U19656 ( .C1(n16359), .C2(n20238), .A(n16358), .B(n16357), .ZN(
        P1_U2985) );
  AOI22_X1 U19657 ( .A1(n20416), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n20473), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16366) );
  NOR2_X1 U19658 ( .A1(n15277), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16361) );
  NOR2_X1 U19659 ( .A1(n15230), .A2(n12675), .ZN(n16360) );
  MUX2_X1 U19660 ( .A(n16361), .B(n16360), .S(n9674), .Z(n16362) );
  XOR2_X1 U19661 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n16362), .Z(
        n16398) );
  AOI22_X1 U19662 ( .A1(n20422), .A2(n16398), .B1(n16364), .B2(n16363), .ZN(
        n16365) );
  OAI211_X1 U19663 ( .C1(n20427), .C2(n16367), .A(n16366), .B(n16365), .ZN(
        P1_U2988) );
  AOI22_X1 U19664 ( .A1(n20416), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20473), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16373) );
  NAND2_X1 U19665 ( .A1(n16370), .A2(n16369), .ZN(n16371) );
  XNOR2_X1 U19666 ( .A(n16368), .B(n16371), .ZN(n16436) );
  AOI22_X1 U19667 ( .A1(n16436), .A2(n20422), .B1(n16364), .B2(n20278), .ZN(
        n16372) );
  OAI211_X1 U19668 ( .C1(n20427), .C2(n20269), .A(n16373), .B(n16372), .ZN(
        P1_U2992) );
  AOI22_X1 U19669 ( .A1(n20416), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20473), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16378) );
  XNOR2_X1 U19670 ( .A(n16375), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16376) );
  XNOR2_X1 U19671 ( .A(n16374), .B(n16376), .ZN(n16442) );
  AOI22_X1 U19672 ( .A1(n16442), .A2(n20422), .B1(n16364), .B2(n20288), .ZN(
        n16377) );
  OAI211_X1 U19673 ( .C1(n20427), .C2(n20281), .A(n16378), .B(n16377), .ZN(
        P1_U2993) );
  AOI22_X1 U19674 ( .A1(n20416), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20473), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n16385) );
  OAI21_X1 U19675 ( .B1(n16381), .B2(n16380), .A(n16379), .ZN(n16449) );
  INV_X1 U19676 ( .A(n16449), .ZN(n16383) );
  INV_X1 U19677 ( .A(n16382), .ZN(n20299) );
  AOI22_X1 U19678 ( .A1(n16383), .A2(n20422), .B1(n16364), .B2(n20299), .ZN(
        n16384) );
  OAI211_X1 U19679 ( .C1(n20427), .C2(n20293), .A(n16385), .B(n16384), .ZN(
        P1_U2994) );
  AOI21_X1 U19680 ( .B1(n16387), .B2(n20440), .A(n16386), .ZN(n16392) );
  INV_X1 U19681 ( .A(n16388), .ZN(n16389) );
  AOI21_X1 U19682 ( .B1(n16390), .B2(n20452), .A(n16389), .ZN(n16391) );
  OAI211_X1 U19683 ( .C1(n16394), .C2(n16393), .A(n16392), .B(n16391), .ZN(
        P1_U3016) );
  NAND2_X1 U19684 ( .A1(n16402), .A2(n16428), .ZN(n16413) );
  NAND3_X1 U19685 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16395), .ZN(n16401) );
  AOI22_X1 U19686 ( .A1(n16396), .A2(n20440), .B1(n20473), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16400) );
  AOI22_X1 U19687 ( .A1(n16398), .A2(n20452), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16397), .ZN(n16399) );
  OAI211_X1 U19688 ( .C1(n16413), .C2(n16401), .A(n16400), .B(n16399), .ZN(
        P1_U3020) );
  OAI21_X1 U19689 ( .B1(n16404), .B2(n16403), .A(n16402), .ZN(n16406) );
  INV_X1 U19690 ( .A(n16405), .ZN(n16422) );
  AOI21_X1 U19691 ( .B1(n16425), .B2(n16406), .A(n16422), .ZN(n16421) );
  AOI221_X1 U19692 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n12675), .C2(n16420), .A(
        n16413), .ZN(n16407) );
  AOI21_X1 U19693 ( .B1(n20473), .B2(P1_REIP_REG_10__SCAN_IN), .A(n16407), 
        .ZN(n16408) );
  OAI21_X1 U19694 ( .B1(n16409), .B2(n20469), .A(n16408), .ZN(n16410) );
  AOI21_X1 U19695 ( .B1(n16411), .B2(n20452), .A(n16410), .ZN(n16412) );
  OAI21_X1 U19696 ( .B1(n16421), .B2(n12675), .A(n16412), .ZN(P1_U3021) );
  NOR2_X1 U19697 ( .A1(n16413), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16417) );
  INV_X1 U19698 ( .A(n20257), .ZN(n16415) );
  OAI22_X1 U19699 ( .A1(n16415), .A2(n20469), .B1(n16414), .B2(n20432), .ZN(
        n16416) );
  AOI211_X1 U19700 ( .C1(n16418), .C2(n20452), .A(n16417), .B(n16416), .ZN(
        n16419) );
  OAI21_X1 U19701 ( .B1(n16421), .B2(n16420), .A(n16419), .ZN(P1_U3022) );
  NAND2_X1 U19702 ( .A1(n20430), .A2(n16447), .ZN(n16453) );
  AOI221_X1 U19703 ( .B1(n20456), .B2(n20450), .C1(n16423), .C2(n20450), .A(
        n16422), .ZN(n16448) );
  OAI21_X1 U19704 ( .B1(n16424), .B2(n16453), .A(n16448), .ZN(n16441) );
  AOI21_X1 U19705 ( .B1(n16426), .B2(n16425), .A(n16441), .ZN(n16438) );
  INV_X1 U19706 ( .A(n16427), .ZN(n16432) );
  NAND2_X1 U19707 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16428), .ZN(
        n16440) );
  AOI221_X1 U19708 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16434), .C2(n16439), .A(
        n16440), .ZN(n16431) );
  OAI22_X1 U19709 ( .A1(n16429), .A2(n20469), .B1(n14479), .B2(n20432), .ZN(
        n16430) );
  AOI211_X1 U19710 ( .C1(n16432), .C2(n20452), .A(n16431), .B(n16430), .ZN(
        n16433) );
  OAI21_X1 U19711 ( .B1(n16438), .B2(n16434), .A(n16433), .ZN(P1_U3023) );
  INV_X1 U19712 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20270) );
  OAI22_X1 U19713 ( .A1(n20268), .A2(n20469), .B1(n20270), .B2(n20432), .ZN(
        n16435) );
  AOI21_X1 U19714 ( .B1(n16436), .B2(n20452), .A(n16435), .ZN(n16437) );
  OAI221_X1 U19715 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16440), .C1(
        n16439), .C2(n16438), .A(n16437), .ZN(P1_U3024) );
  AOI22_X1 U19716 ( .A1(n20282), .A2(n20440), .B1(n20473), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16444) );
  AOI22_X1 U19717 ( .A1(n16442), .A2(n20452), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16441), .ZN(n16443) );
  OAI211_X1 U19718 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16445), .A(
        n16444), .B(n16443), .ZN(P1_U3025) );
  NAND2_X1 U19719 ( .A1(n20454), .A2(n16446), .ZN(n20442) );
  AOI22_X1 U19720 ( .A1(n20294), .A2(n20440), .B1(n20473), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16452) );
  OAI22_X1 U19721 ( .A1(n16449), .A2(n20470), .B1(n16448), .B2(n16447), .ZN(
        n16450) );
  INV_X1 U19722 ( .A(n16450), .ZN(n16451) );
  OAI211_X1 U19723 ( .C1(n16453), .C2(n20442), .A(n16452), .B(n16451), .ZN(
        P1_U3026) );
  INV_X1 U19724 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16459) );
  INV_X1 U19725 ( .A(n20308), .ZN(n16457) );
  NOR3_X1 U19726 ( .A1(n13557), .A2(n16455), .A3(n16454), .ZN(n16456) );
  NAND2_X1 U19727 ( .A1(n16457), .A2(n16456), .ZN(n16458) );
  OAI21_X1 U19728 ( .B1(n16460), .B2(n16459), .A(n16458), .ZN(P1_U3468) );
  NAND4_X1 U19729 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n12006), .A4(n21027), .ZN(n16461) );
  AND2_X1 U19730 ( .A1(n16462), .A2(n16461), .ZN(n20943) );
  AOI21_X1 U19731 ( .B1(n20943), .B2(n16467), .A(n16463), .ZN(n16465) );
  AOI211_X1 U19732 ( .C1(n20942), .C2(n16466), .A(n16465), .B(n16464), .ZN(
        P1_U3162) );
  OAI22_X1 U19733 ( .A1(n16468), .A2(n20774), .B1(n21023), .B2(n16467), .ZN(
        P1_U3466) );
  INV_X1 U19734 ( .A(n19235), .ZN(n19336) );
  INV_X1 U19735 ( .A(n16470), .ZN(n16497) );
  INV_X1 U19736 ( .A(n16471), .ZN(n16473) );
  OAI222_X1 U19737 ( .A1(n19417), .A2(n20150), .B1(n19434), .B2(n16473), .C1(
        n19400), .C2(n16472), .ZN(n16474) );
  AOI21_X1 U19738 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19431), .A(
        n16474), .ZN(n16477) );
  AOI22_X1 U19739 ( .A1(n16475), .A2(n19441), .B1(n19361), .B2(n19448), .ZN(
        n16476) );
  OAI211_X1 U19740 ( .C1(n19336), .C2(n16483), .A(n16477), .B(n16476), .ZN(
        P2_U2824) );
  OAI22_X1 U19741 ( .A1(n19413), .A2(n16478), .B1(n20148), .B2(n19417), .ZN(
        n16479) );
  INV_X1 U19742 ( .A(n16479), .ZN(n16489) );
  AOI22_X1 U19743 ( .A1(n16480), .A2(n19403), .B1(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n19431), .ZN(n16488) );
  OAI22_X1 U19744 ( .A1(n16481), .A2(n19422), .B1(n19447), .B2(n13189), .ZN(
        n16482) );
  INV_X1 U19745 ( .A(n16482), .ZN(n16487) );
  OAI211_X1 U19746 ( .C1(n16485), .C2(n16484), .A(n19443), .B(n16483), .ZN(
        n16486) );
  NAND4_X1 U19747 ( .A1(n16489), .A2(n16488), .A3(n16487), .A4(n16486), .ZN(
        P2_U2825) );
  OAI22_X1 U19748 ( .A1(n19413), .A2(n16490), .B1(n20145), .B2(n19417), .ZN(
        n16491) );
  INV_X1 U19749 ( .A(n16491), .ZN(n16501) );
  AOI22_X1 U19750 ( .A1(n16492), .A2(n19403), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19431), .ZN(n16500) );
  AOI22_X1 U19751 ( .A1(n16494), .A2(n19441), .B1(n19361), .B2(n16493), .ZN(
        n16499) );
  OAI211_X1 U19752 ( .C1(n16497), .C2(n16496), .A(n19443), .B(n16495), .ZN(
        n16498) );
  NAND4_X1 U19753 ( .A1(n16501), .A2(n16500), .A3(n16499), .A4(n16498), .ZN(
        P2_U2826) );
  OAI22_X1 U19754 ( .A1(n19400), .A2(n16502), .B1(n20143), .B2(n19417), .ZN(
        n16503) );
  INV_X1 U19755 ( .A(n16503), .ZN(n16517) );
  OAI22_X1 U19756 ( .A1(n16505), .A2(n19434), .B1(n19397), .B2(n16504), .ZN(
        n16506) );
  INV_X1 U19757 ( .A(n16506), .ZN(n16516) );
  INV_X1 U19758 ( .A(n16507), .ZN(n16508) );
  OAI22_X1 U19759 ( .A1(n16509), .A2(n19422), .B1(n16508), .B2(n19447), .ZN(
        n16510) );
  INV_X1 U19760 ( .A(n16510), .ZN(n16515) );
  OAI211_X1 U19761 ( .C1(n16513), .C2(n16512), .A(n19443), .B(n16511), .ZN(
        n16514) );
  NAND4_X1 U19762 ( .A1(n16517), .A2(n16516), .A3(n16515), .A4(n16514), .ZN(
        P2_U2828) );
  OAI22_X1 U19763 ( .A1(n19413), .A2(n16518), .B1(n20140), .B2(n19417), .ZN(
        n16519) );
  INV_X1 U19764 ( .A(n16519), .ZN(n16530) );
  AOI22_X1 U19765 ( .A1(n16520), .A2(n19403), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19431), .ZN(n16529) );
  OAI22_X1 U19766 ( .A1(n16522), .A2(n19422), .B1(n16521), .B2(n19447), .ZN(
        n16523) );
  INV_X1 U19767 ( .A(n16523), .ZN(n16528) );
  OAI211_X1 U19768 ( .C1(n16526), .C2(n16525), .A(n19443), .B(n16524), .ZN(
        n16527) );
  NAND4_X1 U19769 ( .A1(n16530), .A2(n16529), .A3(n16528), .A4(n16527), .ZN(
        P2_U2829) );
  OAI22_X1 U19770 ( .A1(n19413), .A2(n16531), .B1(n20138), .B2(n19417), .ZN(
        n16532) );
  INV_X1 U19771 ( .A(n16532), .ZN(n16544) );
  OAI22_X1 U19772 ( .A1(n16534), .A2(n19434), .B1(n19397), .B2(n16533), .ZN(
        n16535) );
  INV_X1 U19773 ( .A(n16535), .ZN(n16543) );
  AOI22_X1 U19774 ( .A1(n16537), .A2(n19441), .B1(n16536), .B2(n19361), .ZN(
        n16542) );
  OAI211_X1 U19775 ( .C1(n16540), .C2(n16539), .A(n19443), .B(n16538), .ZN(
        n16541) );
  NAND4_X1 U19776 ( .A1(n16544), .A2(n16543), .A3(n16542), .A4(n16541), .ZN(
        P2_U2830) );
  INV_X1 U19777 ( .A(n16545), .ZN(n16551) );
  INV_X1 U19778 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16546) );
  OAI22_X1 U19779 ( .A1(n19417), .A2(n20136), .B1(n19397), .B2(n16546), .ZN(
        n16547) );
  AOI21_X1 U19780 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n19432), .A(n16547), .ZN(
        n16548) );
  OAI21_X1 U19781 ( .B1(n16549), .B2(n19422), .A(n16548), .ZN(n16550) );
  AOI21_X1 U19782 ( .B1(n16551), .B2(n19403), .A(n16550), .ZN(n16556) );
  OAI211_X1 U19783 ( .C1(n16554), .C2(n16553), .A(n19443), .B(n16552), .ZN(
        n16555) );
  OAI211_X1 U19784 ( .C1(n19447), .C2(n16557), .A(n16556), .B(n16555), .ZN(
        P2_U2831) );
  OAI22_X1 U19785 ( .A1(n19400), .A2(n16558), .B1(n20134), .B2(n19417), .ZN(
        n16559) );
  INV_X1 U19786 ( .A(n16559), .ZN(n16570) );
  AOI22_X1 U19787 ( .A1(n16560), .A2(n19403), .B1(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19431), .ZN(n16569) );
  INV_X1 U19788 ( .A(n16561), .ZN(n16562) );
  AOI22_X1 U19789 ( .A1(n16563), .A2(n19441), .B1(n19361), .B2(n16562), .ZN(
        n16568) );
  OAI211_X1 U19790 ( .C1(n16566), .C2(n16565), .A(n19443), .B(n16564), .ZN(
        n16567) );
  NAND4_X1 U19791 ( .A1(n16570), .A2(n16569), .A3(n16568), .A4(n16567), .ZN(
        P2_U2832) );
  AOI22_X1 U19792 ( .A1(n16572), .A2(n16571), .B1(P2_EAX_REG_17__SCAN_IN), 
        .B2(n19462), .ZN(n16577) );
  AOI22_X1 U19793 ( .A1(n19450), .A2(BUF2_REG_17__SCAN_IN), .B1(n19451), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n16576) );
  INV_X1 U19794 ( .A(n16573), .ZN(n19297) );
  AOI22_X1 U19795 ( .A1(n19297), .A2(n19449), .B1(n13177), .B2(n16574), .ZN(
        n16575) );
  NAND3_X1 U19796 ( .A1(n16577), .A2(n16576), .A3(n16575), .ZN(P2_U2902) );
  AOI22_X1 U19797 ( .A1(n19501), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19500), .ZN(n16584) );
  INV_X1 U19798 ( .A(n16578), .ZN(n16581) );
  INV_X1 U19799 ( .A(n16579), .ZN(n16580) );
  AOI222_X1 U19800 ( .A1(n16582), .A2(n10923), .B1(n19504), .B2(n16581), .C1(
        n19505), .C2(n16580), .ZN(n16583) );
  OAI211_X1 U19801 ( .C1(n19510), .C2(n16585), .A(n16584), .B(n16583), .ZN(
        P2_U2992) );
  AOI22_X1 U19802 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19500), .B1(n16667), 
        .B2(n19321), .ZN(n16590) );
  OAI22_X1 U19803 ( .A1(n16587), .A2(n16671), .B1(n16668), .B2(n16586), .ZN(
        n16588) );
  AOI21_X1 U19804 ( .B1(n19504), .B2(n19322), .A(n16588), .ZN(n16589) );
  OAI211_X1 U19805 ( .C1(n16677), .C2(n16591), .A(n16590), .B(n16589), .ZN(
        P2_U2999) );
  AOI22_X1 U19806 ( .A1(n19501), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19500), .ZN(n16598) );
  NAND2_X1 U19807 ( .A1(n19332), .A2(n19504), .ZN(n16594) );
  NAND2_X1 U19808 ( .A1(n16592), .A2(n10923), .ZN(n16593) );
  OAI211_X1 U19809 ( .C1(n16595), .C2(n16668), .A(n16594), .B(n16593), .ZN(
        n16596) );
  INV_X1 U19810 ( .A(n16596), .ZN(n16597) );
  OAI211_X1 U19811 ( .C1(n19510), .C2(n19327), .A(n16598), .B(n16597), .ZN(
        P2_U3000) );
  AOI22_X1 U19812 ( .A1(n19501), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n16667), .B2(n19348), .ZN(n16609) );
  OAI21_X1 U19813 ( .B1(n16599), .B2(n16601), .A(n16600), .ZN(n16687) );
  AOI22_X1 U19814 ( .A1(n16687), .A2(n10923), .B1(n19504), .B2(n19347), .ZN(
        n16608) );
  NAND2_X1 U19815 ( .A1(n16003), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16604) );
  INV_X1 U19816 ( .A(n16602), .ZN(n16603) );
  AOI21_X1 U19817 ( .B1(n16605), .B2(n16604), .A(n16603), .ZN(n16688) );
  NAND2_X1 U19818 ( .A1(n16688), .A2(n19505), .ZN(n16607) );
  NOR2_X1 U19819 ( .A1(n19395), .A2(n11564), .ZN(n16681) );
  INV_X1 U19820 ( .A(n16681), .ZN(n16606) );
  NAND4_X1 U19821 ( .A1(n16609), .A2(n16608), .A3(n16607), .A4(n16606), .ZN(
        P2_U3001) );
  AOI22_X1 U19822 ( .A1(n19501), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19500), .ZN(n16613) );
  AOI222_X1 U19823 ( .A1(n16611), .A2(n19505), .B1(n10923), .B2(n16610), .C1(
        n19504), .C2(n10090), .ZN(n16612) );
  OAI211_X1 U19824 ( .C1(n19510), .C2(n19354), .A(n16613), .B(n16612), .ZN(
        P2_U3002) );
  AOI22_X1 U19825 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19500), .B1(n16667), 
        .B2(n19373), .ZN(n16618) );
  OAI22_X1 U19826 ( .A1(n16615), .A2(n16668), .B1(n16614), .B2(n16671), .ZN(
        n16616) );
  AOI21_X1 U19827 ( .B1(n19504), .B2(n19374), .A(n16616), .ZN(n16617) );
  OAI211_X1 U19828 ( .C1(n16677), .C2(n16619), .A(n16618), .B(n16617), .ZN(
        P2_U3003) );
  AOI22_X1 U19829 ( .A1(n19501), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19500), .ZN(n16631) );
  INV_X1 U19830 ( .A(n16621), .ZN(n16622) );
  NOR2_X1 U19831 ( .A1(n16620), .A2(n16622), .ZN(n16626) );
  NAND2_X1 U19832 ( .A1(n16624), .A2(n16623), .ZN(n16625) );
  XNOR2_X1 U19833 ( .A(n16626), .B(n16625), .ZN(n16705) );
  INV_X1 U19834 ( .A(n16705), .ZN(n16629) );
  AOI21_X1 U19835 ( .B1(n16694), .B2(n16628), .A(n16627), .ZN(n16701) );
  AOI222_X1 U19836 ( .A1(n16629), .A2(n10923), .B1(n19504), .B2(n16698), .C1(
        n19505), .C2(n16701), .ZN(n16630) );
  OAI211_X1 U19837 ( .C1(n19510), .C2(n16632), .A(n16631), .B(n16630), .ZN(
        P2_U3004) );
  AOI22_X1 U19838 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19500), .B1(n16667), 
        .B2(n19386), .ZN(n16637) );
  OAI22_X1 U19839 ( .A1(n16634), .A2(n16668), .B1(n16671), .B2(n16633), .ZN(
        n16635) );
  AOI21_X1 U19840 ( .B1(n19504), .B2(n19387), .A(n16635), .ZN(n16636) );
  OAI211_X1 U19841 ( .C1(n16677), .C2(n19381), .A(n16637), .B(n16636), .ZN(
        P2_U3005) );
  AOI22_X1 U19842 ( .A1(n19501), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19500), .ZN(n16658) );
  NAND2_X1 U19843 ( .A1(n16639), .A2(n16638), .ZN(n16641) );
  NAND2_X1 U19844 ( .A1(n16641), .A2(n16640), .ZN(n16644) );
  INV_X1 U19845 ( .A(n16642), .ZN(n16643) );
  XNOR2_X1 U19846 ( .A(n16644), .B(n16643), .ZN(n16714) );
  NAND2_X1 U19847 ( .A1(n16714), .A2(n19505), .ZN(n16654) );
  NAND2_X1 U19848 ( .A1(n16646), .A2(n16645), .ZN(n16648) );
  NAND2_X1 U19849 ( .A1(n16648), .A2(n16647), .ZN(n16652) );
  NAND2_X1 U19850 ( .A1(n16650), .A2(n16649), .ZN(n16651) );
  XNOR2_X1 U19851 ( .A(n16652), .B(n16651), .ZN(n16720) );
  NAND2_X1 U19852 ( .A1(n16720), .A2(n10923), .ZN(n16653) );
  OAI211_X1 U19853 ( .C1(n16655), .C2(n16715), .A(n16654), .B(n16653), .ZN(
        n16656) );
  INV_X1 U19854 ( .A(n16656), .ZN(n16657) );
  OAI211_X1 U19855 ( .C1(n19510), .C2(n16659), .A(n16658), .B(n16657), .ZN(
        P2_U3006) );
  AOI22_X1 U19856 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19500), .B1(n16667), 
        .B2(n19440), .ZN(n16664) );
  OAI22_X1 U19857 ( .A1(n16661), .A2(n16671), .B1(n16660), .B2(n16668), .ZN(
        n16662) );
  AOI21_X1 U19858 ( .B1(n19504), .B2(n19442), .A(n16662), .ZN(n16663) );
  OAI211_X1 U19859 ( .C1(n16677), .C2(n16665), .A(n16664), .B(n16663), .ZN(
        P2_U3009) );
  AOI22_X1 U19860 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19500), .B1(n16667), 
        .B2(n16666), .ZN(n16676) );
  NOR3_X1 U19861 ( .A1(n16670), .A2(n16669), .A3(n16668), .ZN(n16674) );
  NOR2_X1 U19862 ( .A1(n16672), .A2(n16671), .ZN(n16673) );
  AOI211_X1 U19863 ( .C1(n19504), .C2(n9734), .A(n16674), .B(n16673), .ZN(
        n16675) );
  OAI211_X1 U19864 ( .C1(n16678), .C2(n16677), .A(n16676), .B(n16675), .ZN(
        P2_U3011) );
  INV_X1 U19865 ( .A(n16679), .ZN(n16685) );
  AOI21_X1 U19866 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n16680), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16684) );
  INV_X1 U19867 ( .A(n19352), .ZN(n16682) );
  AOI21_X1 U19868 ( .B1(n16710), .B2(n16682), .A(n16681), .ZN(n16683) );
  OAI21_X1 U19869 ( .B1(n16685), .B2(n16684), .A(n16683), .ZN(n16686) );
  AOI21_X1 U19870 ( .B1(n16687), .B2(n16721), .A(n16686), .ZN(n16690) );
  AOI22_X1 U19871 ( .A1(n16688), .A2(n16700), .B1(n16699), .B2(n19347), .ZN(
        n16689) );
  NAND2_X1 U19872 ( .A1(n16690), .A2(n16689), .ZN(P2_U3033) );
  INV_X1 U19873 ( .A(n16691), .ZN(n16697) );
  NAND2_X1 U19874 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19500), .ZN(n16692) );
  OAI221_X1 U19875 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16695), 
        .C1(n16694), .C2(n16693), .A(n16692), .ZN(n16696) );
  AOI21_X1 U19876 ( .B1(n16697), .B2(n16710), .A(n16696), .ZN(n16703) );
  AOI22_X1 U19877 ( .A1(n16701), .A2(n16700), .B1(n16699), .B2(n16698), .ZN(
        n16702) );
  OAI211_X1 U19878 ( .C1(n16705), .C2(n16704), .A(n16703), .B(n16702), .ZN(
        P2_U3036) );
  AOI211_X1 U19879 ( .C1(n10816), .C2(n16708), .A(n16707), .B(n16706), .ZN(
        n16713) );
  NAND2_X1 U19880 ( .A1(n16710), .A2(n16709), .ZN(n16711) );
  OAI21_X1 U19881 ( .B1(n11438), .B2(n19341), .A(n16711), .ZN(n16712) );
  NOR2_X1 U19882 ( .A1(n16713), .A2(n16712), .ZN(n16723) );
  INV_X1 U19883 ( .A(n16714), .ZN(n16718) );
  OAI22_X1 U19884 ( .A1(n16718), .A2(n16717), .B1(n16716), .B2(n16715), .ZN(
        n16719) );
  AOI21_X1 U19885 ( .B1(n16721), .B2(n16720), .A(n16719), .ZN(n16722) );
  OAI211_X1 U19886 ( .C1(n16724), .C2(n10816), .A(n16723), .B(n16722), .ZN(
        P2_U3038) );
  INV_X1 U19887 ( .A(n16725), .ZN(n16728) );
  NAND2_X1 U19888 ( .A1(n20215), .A2(n19942), .ZN(n20078) );
  OAI22_X1 U19889 ( .A1(n20208), .A2(n16726), .B1(n20078), .B2(n20218), .ZN(
        n16727) );
  AOI211_X1 U19890 ( .C1(n16729), .C2(P2_STATE2_REG_0__SCAN_IN), .A(n16728), 
        .B(n16727), .ZN(n16731) );
  NAND2_X1 U19891 ( .A1(n16729), .A2(n20215), .ZN(n20083) );
  OAI211_X1 U19892 ( .C1(n19205), .C2(n20161), .A(n20218), .B(n20083), .ZN(
        n16730) );
  OAI211_X1 U19893 ( .C1(n16732), .C2(n19210), .A(n16731), .B(n16730), .ZN(
        P2_U3176) );
  INV_X1 U19894 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16889) );
  XNOR2_X1 U19895 ( .A(n16889), .B(n16733), .ZN(n16888) );
  NAND2_X1 U19896 ( .A1(n18499), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16734) );
  OAI221_X1 U19897 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16736), .C1(
        n16889), .C2(n16735), .A(n16734), .ZN(n16737) );
  AOI21_X1 U19898 ( .B1(n18036), .B2(n16888), .A(n16737), .ZN(n16743) );
  OAI22_X1 U19899 ( .A1(n16739), .A2(n18027), .B1(n16738), .B2(n18180), .ZN(
        n16741) );
  AOI22_X1 U19900 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16741), .B1(
        n17841), .B2(n16740), .ZN(n16742) );
  OAI211_X1 U19901 ( .C1(n16744), .C2(n18093), .A(n16743), .B(n16742), .ZN(
        P3_U2800) );
  NOR3_X1 U19902 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16746) );
  NOR4_X1 U19903 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16745) );
  INV_X2 U19904 ( .A(n16842), .ZN(U215) );
  NAND4_X1 U19905 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16746), .A3(n16745), .A4(
        U215), .ZN(U213) );
  INV_X1 U19906 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16844) );
  INV_X2 U19907 ( .A(U214), .ZN(n16805) );
  INV_X1 U19908 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16845) );
  OAI222_X1 U19909 ( .A1(U212), .A2(n16844), .B1(n16807), .B2(n16748), .C1(
        U214), .C2(n16845), .ZN(U216) );
  AOI22_X1 U19910 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16791), .ZN(n16749) );
  OAI21_X1 U19911 ( .B1(n19556), .B2(n16807), .A(n16749), .ZN(U217) );
  AOI22_X1 U19912 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16791), .ZN(n16750) );
  OAI21_X1 U19913 ( .B1(n16751), .B2(n16807), .A(n16750), .ZN(U218) );
  AOI22_X1 U19914 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16791), .ZN(n16752) );
  OAI21_X1 U19915 ( .B1(n16753), .B2(n16807), .A(n16752), .ZN(U219) );
  AOI22_X1 U19916 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16791), .ZN(n16754) );
  OAI21_X1 U19917 ( .B1(n16755), .B2(n16807), .A(n16754), .ZN(U220) );
  AOI22_X1 U19918 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16791), .ZN(n16756) );
  OAI21_X1 U19919 ( .B1(n16757), .B2(n16807), .A(n16756), .ZN(U221) );
  AOI22_X1 U19920 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16791), .ZN(n16758) );
  OAI21_X1 U19921 ( .B1(n16759), .B2(n16807), .A(n16758), .ZN(U222) );
  AOI22_X1 U19922 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16791), .ZN(n16760) );
  OAI21_X1 U19923 ( .B1(n16761), .B2(n16807), .A(n16760), .ZN(U223) );
  AOI22_X1 U19924 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16791), .ZN(n16762) );
  OAI21_X1 U19925 ( .B1(n16763), .B2(n16807), .A(n16762), .ZN(U224) );
  AOI22_X1 U19926 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16791), .ZN(n16764) );
  OAI21_X1 U19927 ( .B1(n16765), .B2(n16807), .A(n16764), .ZN(U225) );
  AOI22_X1 U19928 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16791), .ZN(n16766) );
  OAI21_X1 U19929 ( .B1(n19550), .B2(n16807), .A(n16766), .ZN(U226) );
  AOI22_X1 U19930 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16791), .ZN(n16767) );
  OAI21_X1 U19931 ( .B1(n16768), .B2(n16807), .A(n16767), .ZN(U227) );
  AOI22_X1 U19932 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16791), .ZN(n16769) );
  OAI21_X1 U19933 ( .B1(n16770), .B2(n16807), .A(n16769), .ZN(U228) );
  AOI22_X1 U19934 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16791), .ZN(n16771) );
  OAI21_X1 U19935 ( .B1(n16772), .B2(n16807), .A(n16771), .ZN(U229) );
  AOI22_X1 U19936 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16791), .ZN(n16773) );
  OAI21_X1 U19937 ( .B1(n16774), .B2(n16807), .A(n16773), .ZN(U230) );
  AOI22_X1 U19938 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16791), .ZN(n16775) );
  OAI21_X1 U19939 ( .B1(n16776), .B2(n16807), .A(n16775), .ZN(U231) );
  INV_X1 U19940 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n16778) );
  AOI22_X1 U19941 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16791), .ZN(n16777) );
  OAI21_X1 U19942 ( .B1(n16778), .B2(n16807), .A(n16777), .ZN(U232) );
  AOI22_X1 U19943 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n16791), .ZN(n16779) );
  OAI21_X1 U19944 ( .B1(n16780), .B2(n16807), .A(n16779), .ZN(U233) );
  AOI22_X1 U19945 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16791), .ZN(n16781) );
  OAI21_X1 U19946 ( .B1(n14528), .B2(n16807), .A(n16781), .ZN(U234) );
  AOI22_X1 U19947 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16791), .ZN(n16782) );
  OAI21_X1 U19948 ( .B1(n16783), .B2(n16807), .A(n16782), .ZN(U235) );
  AOI22_X1 U19949 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16791), .ZN(n16784) );
  OAI21_X1 U19950 ( .B1(n16785), .B2(n16807), .A(n16784), .ZN(U236) );
  AOI22_X1 U19951 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16791), .ZN(n16786) );
  OAI21_X1 U19952 ( .B1(n14579), .B2(n16807), .A(n16786), .ZN(U237) );
  AOI22_X1 U19953 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16791), .ZN(n16787) );
  OAI21_X1 U19954 ( .B1(n16788), .B2(n16807), .A(n16787), .ZN(U238) );
  AOI22_X1 U19955 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16791), .ZN(n16789) );
  OAI21_X1 U19956 ( .B1(n16790), .B2(n16807), .A(n16789), .ZN(U239) );
  AOI22_X1 U19957 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16791), .ZN(n16792) );
  OAI21_X1 U19958 ( .B1(n13791), .B2(n16807), .A(n16792), .ZN(U240) );
  INV_X1 U19959 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16794) );
  AOI22_X1 U19960 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n16791), .ZN(n16793) );
  OAI21_X1 U19961 ( .B1(n16794), .B2(n16807), .A(n16793), .ZN(U241) );
  AOI22_X1 U19962 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16791), .ZN(n16795) );
  OAI21_X1 U19963 ( .B1(n16796), .B2(n16807), .A(n16795), .ZN(U242) );
  INV_X1 U19964 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16798) );
  AOI22_X1 U19965 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16791), .ZN(n16797) );
  OAI21_X1 U19966 ( .B1(n16798), .B2(n16807), .A(n16797), .ZN(U243) );
  INV_X1 U19967 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16800) );
  AOI22_X1 U19968 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16791), .ZN(n16799) );
  OAI21_X1 U19969 ( .B1(n16800), .B2(n16807), .A(n16799), .ZN(U244) );
  INV_X1 U19970 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16802) );
  AOI22_X1 U19971 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16791), .ZN(n16801) );
  OAI21_X1 U19972 ( .B1(n16802), .B2(n16807), .A(n16801), .ZN(U245) );
  INV_X1 U19973 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n16804) );
  AOI22_X1 U19974 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16791), .ZN(n16803) );
  OAI21_X1 U19975 ( .B1(n16804), .B2(n16807), .A(n16803), .ZN(U246) );
  INV_X1 U19976 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16808) );
  AOI22_X1 U19977 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16805), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16791), .ZN(n16806) );
  OAI21_X1 U19978 ( .B1(n16808), .B2(n16807), .A(n16806), .ZN(U247) );
  OAI22_X1 U19979 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16842), .ZN(n16809) );
  INV_X1 U19980 ( .A(n16809), .ZN(U251) );
  OAI22_X1 U19981 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16842), .ZN(n16810) );
  INV_X1 U19982 ( .A(n16810), .ZN(U252) );
  OAI22_X1 U19983 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16842), .ZN(n16811) );
  INV_X1 U19984 ( .A(n16811), .ZN(U253) );
  OAI22_X1 U19985 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16842), .ZN(n16812) );
  INV_X1 U19986 ( .A(n16812), .ZN(U254) );
  OAI22_X1 U19987 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16842), .ZN(n16813) );
  INV_X1 U19988 ( .A(n16813), .ZN(U255) );
  OAI22_X1 U19989 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16842), .ZN(n16814) );
  INV_X1 U19990 ( .A(n16814), .ZN(U256) );
  OAI22_X1 U19991 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16842), .ZN(n16815) );
  INV_X1 U19992 ( .A(n16815), .ZN(U257) );
  OAI22_X1 U19993 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16842), .ZN(n16816) );
  INV_X1 U19994 ( .A(n16816), .ZN(U258) );
  OAI22_X1 U19995 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16842), .ZN(n16817) );
  INV_X1 U19996 ( .A(n16817), .ZN(U259) );
  OAI22_X1 U19997 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16836), .ZN(n16818) );
  INV_X1 U19998 ( .A(n16818), .ZN(U260) );
  OAI22_X1 U19999 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16836), .ZN(n16819) );
  INV_X1 U20000 ( .A(n16819), .ZN(U261) );
  OAI22_X1 U20001 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16842), .ZN(n16820) );
  INV_X1 U20002 ( .A(n16820), .ZN(U262) );
  OAI22_X1 U20003 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16842), .ZN(n16821) );
  INV_X1 U20004 ( .A(n16821), .ZN(U263) );
  OAI22_X1 U20005 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16842), .ZN(n16822) );
  INV_X1 U20006 ( .A(n16822), .ZN(U264) );
  OAI22_X1 U20007 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16842), .ZN(n16823) );
  INV_X1 U20008 ( .A(n16823), .ZN(U265) );
  OAI22_X1 U20009 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16836), .ZN(n16824) );
  INV_X1 U20010 ( .A(n16824), .ZN(U266) );
  OAI22_X1 U20011 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16836), .ZN(n16825) );
  INV_X1 U20012 ( .A(n16825), .ZN(U267) );
  OAI22_X1 U20013 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16836), .ZN(n16826) );
  INV_X1 U20014 ( .A(n16826), .ZN(U268) );
  OAI22_X1 U20015 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16836), .ZN(n16827) );
  INV_X1 U20016 ( .A(n16827), .ZN(U269) );
  OAI22_X1 U20017 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16836), .ZN(n16828) );
  INV_X1 U20018 ( .A(n16828), .ZN(U270) );
  OAI22_X1 U20019 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16836), .ZN(n16829) );
  INV_X1 U20020 ( .A(n16829), .ZN(U271) );
  OAI22_X1 U20021 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16842), .ZN(n16830) );
  INV_X1 U20022 ( .A(n16830), .ZN(U272) );
  OAI22_X1 U20023 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16842), .ZN(n16831) );
  INV_X1 U20024 ( .A(n16831), .ZN(U273) );
  OAI22_X1 U20025 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16836), .ZN(n16832) );
  INV_X1 U20026 ( .A(n16832), .ZN(U274) );
  OAI22_X1 U20027 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16842), .ZN(n16833) );
  INV_X1 U20028 ( .A(n16833), .ZN(U275) );
  OAI22_X1 U20029 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16842), .ZN(n16834) );
  INV_X1 U20030 ( .A(n16834), .ZN(U276) );
  OAI22_X1 U20031 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16842), .ZN(n16835) );
  INV_X1 U20032 ( .A(n16835), .ZN(U277) );
  OAI22_X1 U20033 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16836), .ZN(n16837) );
  INV_X1 U20034 ( .A(n16837), .ZN(U278) );
  OAI22_X1 U20035 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16842), .ZN(n16838) );
  INV_X1 U20036 ( .A(n16838), .ZN(U279) );
  OAI22_X1 U20037 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16842), .ZN(n16839) );
  INV_X1 U20038 ( .A(n16839), .ZN(U280) );
  OAI22_X1 U20039 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16842), .ZN(n16841) );
  INV_X1 U20040 ( .A(n16841), .ZN(U281) );
  INV_X1 U20041 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n17566) );
  AOI22_X1 U20042 ( .A1(n16842), .A2(n16844), .B1(n17566), .B2(U215), .ZN(U282) );
  INV_X1 U20043 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16843) );
  AOI222_X1 U20044 ( .A1(n16845), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16844), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16843), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16846) );
  INV_X2 U20045 ( .A(n16848), .ZN(n16847) );
  INV_X1 U20046 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19085) );
  INV_X1 U20047 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n20115) );
  AOI22_X1 U20048 ( .A1(n16847), .A2(n19085), .B1(n20115), .B2(n16848), .ZN(
        U347) );
  INV_X1 U20049 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19083) );
  INV_X1 U20050 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20114) );
  AOI22_X1 U20051 ( .A1(n16847), .A2(n19083), .B1(n20114), .B2(n16848), .ZN(
        U348) );
  INV_X1 U20052 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19081) );
  INV_X1 U20053 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n20113) );
  AOI22_X1 U20054 ( .A1(n16847), .A2(n19081), .B1(n20113), .B2(n16848), .ZN(
        U349) );
  INV_X1 U20055 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19079) );
  INV_X1 U20056 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n20112) );
  AOI22_X1 U20057 ( .A1(n16847), .A2(n19079), .B1(n20112), .B2(n16848), .ZN(
        U350) );
  INV_X1 U20058 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19077) );
  INV_X1 U20059 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20110) );
  AOI22_X1 U20060 ( .A1(n16847), .A2(n19077), .B1(n20110), .B2(n16848), .ZN(
        U351) );
  INV_X1 U20061 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n19074) );
  INV_X1 U20062 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n20108) );
  AOI22_X1 U20063 ( .A1(n16847), .A2(n19074), .B1(n20108), .B2(n16848), .ZN(
        U352) );
  INV_X1 U20064 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n19073) );
  INV_X1 U20065 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n20107) );
  AOI22_X1 U20066 ( .A1(n16847), .A2(n19073), .B1(n20107), .B2(n16848), .ZN(
        U353) );
  INV_X1 U20067 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n19071) );
  AOI22_X1 U20068 ( .A1(n16847), .A2(n19071), .B1(n20106), .B2(n16848), .ZN(
        U354) );
  INV_X1 U20069 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19123) );
  INV_X1 U20070 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n20146) );
  AOI22_X1 U20071 ( .A1(n16847), .A2(n19123), .B1(n20146), .B2(n16848), .ZN(
        U356) );
  INV_X1 U20072 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19120) );
  INV_X1 U20073 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n20144) );
  AOI22_X1 U20074 ( .A1(n16847), .A2(n19120), .B1(n20144), .B2(n16848), .ZN(
        U357) );
  INV_X1 U20075 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19119) );
  INV_X1 U20076 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n20142) );
  AOI22_X1 U20077 ( .A1(n16847), .A2(n19119), .B1(n20142), .B2(n16848), .ZN(
        U358) );
  INV_X1 U20078 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19117) );
  INV_X1 U20079 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n20141) );
  AOI22_X1 U20080 ( .A1(n16847), .A2(n19117), .B1(n20141), .B2(n16848), .ZN(
        U359) );
  INV_X1 U20081 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19115) );
  INV_X1 U20082 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n20139) );
  AOI22_X1 U20083 ( .A1(n16847), .A2(n19115), .B1(n20139), .B2(n16848), .ZN(
        U360) );
  INV_X1 U20084 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19113) );
  INV_X1 U20085 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n20137) );
  AOI22_X1 U20086 ( .A1(n16847), .A2(n19113), .B1(n20137), .B2(n16848), .ZN(
        U361) );
  INV_X1 U20087 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19110) );
  INV_X1 U20088 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n20135) );
  AOI22_X1 U20089 ( .A1(n16847), .A2(n19110), .B1(n20135), .B2(n16848), .ZN(
        U362) );
  INV_X1 U20090 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19109) );
  INV_X1 U20091 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n20133) );
  AOI22_X1 U20092 ( .A1(n16847), .A2(n19109), .B1(n20133), .B2(n16848), .ZN(
        U363) );
  INV_X1 U20093 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19106) );
  INV_X1 U20094 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n20132) );
  AOI22_X1 U20095 ( .A1(n16847), .A2(n19106), .B1(n20132), .B2(n16848), .ZN(
        U364) );
  INV_X1 U20096 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n19069) );
  INV_X1 U20097 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20105) );
  AOI22_X1 U20098 ( .A1(n16847), .A2(n19069), .B1(n20105), .B2(n16848), .ZN(
        U365) );
  INV_X1 U20099 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n19105) );
  INV_X1 U20100 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n20130) );
  AOI22_X1 U20101 ( .A1(n16847), .A2(n19105), .B1(n20130), .B2(n16848), .ZN(
        U366) );
  INV_X1 U20102 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n19103) );
  INV_X1 U20103 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n20128) );
  AOI22_X1 U20104 ( .A1(n16847), .A2(n19103), .B1(n20128), .B2(n16848), .ZN(
        U367) );
  INV_X1 U20105 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19101) );
  INV_X1 U20106 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n20126) );
  AOI22_X1 U20107 ( .A1(n16847), .A2(n19101), .B1(n20126), .B2(n16848), .ZN(
        U368) );
  INV_X1 U20108 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19098) );
  INV_X1 U20109 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n20124) );
  AOI22_X1 U20110 ( .A1(n16847), .A2(n19098), .B1(n20124), .B2(n16848), .ZN(
        U369) );
  INV_X1 U20111 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19097) );
  INV_X1 U20112 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n20122) );
  AOI22_X1 U20113 ( .A1(n16847), .A2(n19097), .B1(n20122), .B2(n16848), .ZN(
        U370) );
  INV_X1 U20114 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19095) );
  INV_X1 U20115 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n20121) );
  AOI22_X1 U20116 ( .A1(n16847), .A2(n19095), .B1(n20121), .B2(n16848), .ZN(
        U371) );
  INV_X1 U20117 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19092) );
  INV_X1 U20118 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n20119) );
  AOI22_X1 U20119 ( .A1(n16847), .A2(n19092), .B1(n20119), .B2(n16848), .ZN(
        U372) );
  INV_X1 U20120 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19091) );
  INV_X1 U20121 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n20118) );
  AOI22_X1 U20122 ( .A1(n16847), .A2(n19091), .B1(n20118), .B2(n16848), .ZN(
        U373) );
  INV_X1 U20123 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19089) );
  INV_X1 U20124 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n20117) );
  AOI22_X1 U20125 ( .A1(n16847), .A2(n19089), .B1(n20117), .B2(n16848), .ZN(
        U374) );
  INV_X1 U20126 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19087) );
  INV_X1 U20127 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n20116) );
  AOI22_X1 U20128 ( .A1(n16847), .A2(n19087), .B1(n20116), .B2(n16848), .ZN(
        U375) );
  INV_X1 U20129 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n19066) );
  INV_X1 U20130 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n20103) );
  AOI22_X1 U20131 ( .A1(n16847), .A2(n19066), .B1(n20103), .B2(n16848), .ZN(
        U376) );
  INV_X1 U20132 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n19065) );
  NAND2_X1 U20133 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n19065), .ZN(n19056) );
  AOI22_X1 U20134 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n19056), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n19063), .ZN(n19135) );
  AOI21_X1 U20135 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n19135), .ZN(n16849) );
  INV_X1 U20136 ( .A(n16849), .ZN(P3_U2633) );
  INV_X1 U20137 ( .A(n16855), .ZN(n16850) );
  OAI21_X1 U20138 ( .B1(n16850), .B2(n17764), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16851) );
  OAI21_X1 U20139 ( .B1(n16852), .B2(n19041), .A(n16851), .ZN(P3_U2634) );
  AOI21_X1 U20140 ( .B1(n19063), .B2(n19065), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16853) );
  AOI22_X1 U20141 ( .A1(n19126), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16853), 
        .B2(n19194), .ZN(P3_U2635) );
  NOR2_X1 U20142 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n19050) );
  OAI21_X1 U20143 ( .B1(n19050), .B2(BS16), .A(n19135), .ZN(n19133) );
  OAI21_X1 U20144 ( .B1(n19135), .B2(n19185), .A(n19133), .ZN(P3_U2636) );
  AND3_X1 U20145 ( .A1(n16855), .A2(n18970), .A3(n16854), .ZN(n18973) );
  NOR2_X1 U20146 ( .A1(n18973), .A2(n19036), .ZN(n19177) );
  OAI21_X1 U20147 ( .B1(n19177), .B2(n18506), .A(n16856), .ZN(P3_U2637) );
  NOR4_X1 U20148 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16860) );
  NOR4_X1 U20149 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16859) );
  NOR4_X1 U20150 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16858) );
  NOR4_X1 U20151 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16857) );
  NAND4_X1 U20152 ( .A1(n16860), .A2(n16859), .A3(n16858), .A4(n16857), .ZN(
        n16866) );
  NOR4_X1 U20153 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_5__SCAN_IN), .A3(P3_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n16864) );
  AOI211_X1 U20154 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_2__SCAN_IN), .B(
        P3_DATAWIDTH_REG_3__SCAN_IN), .ZN(n16863) );
  NOR4_X1 U20155 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16862) );
  NOR4_X1 U20156 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16861) );
  NAND4_X1 U20157 ( .A1(n16864), .A2(n16863), .A3(n16862), .A4(n16861), .ZN(
        n16865) );
  NOR2_X1 U20158 ( .A1(n16866), .A2(n16865), .ZN(n19167) );
  INV_X1 U20159 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16868) );
  INV_X1 U20160 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19134) );
  NAND2_X1 U20161 ( .A1(n19167), .A2(n19134), .ZN(n19168) );
  NOR3_X1 U20162 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A3(n19168), .ZN(n16869) );
  INV_X1 U20163 ( .A(n16869), .ZN(n16867) );
  NAND2_X1 U20164 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n19167), .ZN(n19171) );
  OAI211_X1 U20165 ( .C1(n19167), .C2(n16868), .A(n16867), .B(n19171), .ZN(
        P3_U2638) );
  NOR2_X1 U20166 ( .A1(n16869), .A2(n19171), .ZN(n16871) );
  NOR2_X1 U20167 ( .A1(P3_BYTEENABLE_REG_3__SCAN_IN), .A2(n19167), .ZN(n16870)
         );
  AOI211_X1 U20168 ( .C1(n19167), .C2(P3_DATAWIDTH_REG_1__SCAN_IN), .A(n16871), 
        .B(n16870), .ZN(P3_U2639) );
  INV_X1 U20169 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n19128) );
  NAND4_X1 U20170 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16909), .ZN(n16881) );
  NOR3_X1 U20171 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n19128), .A3(n16881), 
        .ZN(n16873) );
  AOI21_X1 U20172 ( .B1(n17220), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16873), .ZN(
        n16884) );
  INV_X1 U20173 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16926) );
  NAND2_X1 U20174 ( .A1(n16927), .A2(n16926), .ZN(n16925) );
  NOR2_X1 U20175 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16925), .ZN(n16910) );
  INV_X1 U20176 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n17268) );
  NAND2_X1 U20177 ( .A1(n16910), .A2(n17268), .ZN(n16886) );
  NOR2_X1 U20178 ( .A1(n17216), .A2(n16886), .ZN(n16893) );
  INV_X1 U20179 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17233) );
  INV_X1 U20180 ( .A(n16874), .ZN(n16913) );
  AOI21_X1 U20181 ( .B1(n16876), .B2(n17838), .A(n16875), .ZN(n17833) );
  NOR2_X1 U20182 ( .A1(n16877), .A2(n17175), .ZN(n16921) );
  NOR2_X1 U20183 ( .A1(n17833), .A2(n16921), .ZN(n16920) );
  NOR2_X1 U20184 ( .A1(n16920), .A2(n17175), .ZN(n16912) );
  NOR2_X1 U20185 ( .A1(n16913), .A2(n16912), .ZN(n16911) );
  OR2_X1 U20186 ( .A1(n16911), .A2(n17175), .ZN(n16896) );
  INV_X1 U20187 ( .A(n16900), .ZN(n16878) );
  NAND2_X1 U20188 ( .A1(n16896), .A2(n16878), .ZN(n16897) );
  NAND3_X1 U20189 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16880) );
  INV_X1 U20190 ( .A(n17010), .ZN(n17218) );
  AOI21_X1 U20191 ( .B1(n16880), .B2(n17218), .A(n16879), .ZN(n16902) );
  NOR2_X1 U20192 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16881), .ZN(n16891) );
  INV_X1 U20193 ( .A(n16891), .ZN(n16882) );
  AOI21_X1 U20194 ( .B1(n16902), .B2(n16882), .A(n19125), .ZN(n16883) );
  NAND2_X1 U20195 ( .A1(n17219), .A2(n16886), .ZN(n16907) );
  XOR2_X1 U20196 ( .A(n16888), .B(n16887), .Z(n16892) );
  OAI22_X1 U20197 ( .A1(n16902), .A2(n19128), .B1(n16889), .B2(n17206), .ZN(
        n16890) );
  AOI211_X1 U20198 ( .C1(n16892), .C2(n19045), .A(n16891), .B(n16890), .ZN(
        n16895) );
  OAI21_X1 U20199 ( .B1(n17220), .B2(n16893), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16894) );
  OAI211_X1 U20200 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16907), .A(n16895), .B(
        n16894), .ZN(P3_U2641) );
  NOR2_X1 U20201 ( .A1(n16910), .A2(n17268), .ZN(n16908) );
  INV_X1 U20202 ( .A(n16896), .ZN(n16899) );
  INV_X1 U20203 ( .A(n16897), .ZN(n16898) );
  AOI211_X1 U20204 ( .C1(n16900), .C2(n16899), .A(n16898), .B(n17176), .ZN(
        n16904) );
  INV_X1 U20205 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n19122) );
  OAI22_X1 U20206 ( .A1(n16902), .A2(n19122), .B1(n16901), .B2(n17206), .ZN(
        n16903) );
  AOI211_X1 U20207 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n17220), .A(n16904), .B(
        n16903), .ZN(n16906) );
  NAND4_X1 U20208 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16909), .A4(n19122), .ZN(n16905) );
  OAI211_X1 U20209 ( .C1(n16908), .C2(n16907), .A(n16906), .B(n16905), .ZN(
        P3_U2642) );
  NAND2_X1 U20210 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16909), .ZN(n16919) );
  AOI22_X1 U20211 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17192), .B1(
        n17220), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16918) );
  INV_X1 U20212 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n19118) );
  NAND2_X1 U20213 ( .A1(n16909), .A2(n19118), .ZN(n16929) );
  NAND2_X1 U20214 ( .A1(n16922), .A2(n16929), .ZN(n16916) );
  AOI211_X1 U20215 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16925), .A(n16910), .B(
        n17216), .ZN(n16915) );
  AOI211_X1 U20216 ( .C1(n16913), .C2(n16912), .A(n16911), .B(n17176), .ZN(
        n16914) );
  AOI211_X1 U20217 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16916), .A(n16915), 
        .B(n16914), .ZN(n16917) );
  OAI211_X1 U20218 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16919), .A(n16918), 
        .B(n16917), .ZN(P3_U2643) );
  AOI211_X1 U20219 ( .C1(n17833), .C2(n16921), .A(n16920), .B(n17176), .ZN(
        n16924) );
  OAI22_X1 U20220 ( .A1(n16922), .A2(n19118), .B1(n17838), .B2(n17206), .ZN(
        n16923) );
  AOI211_X1 U20221 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n17220), .A(n16924), .B(
        n16923), .ZN(n16930) );
  OAI211_X1 U20222 ( .C1(n16927), .C2(n16926), .A(n17219), .B(n16925), .ZN(
        n16928) );
  NAND3_X1 U20223 ( .A1(n16930), .A2(n16929), .A3(n16928), .ZN(P3_U2644) );
  INV_X1 U20224 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n16943) );
  INV_X1 U20225 ( .A(n16931), .ZN(n16934) );
  NOR2_X1 U20226 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n17210), .ZN(n16950) );
  NOR2_X1 U20227 ( .A1(n16932), .A2(n16950), .ZN(n16933) );
  MUX2_X1 U20228 ( .A(n16934), .B(n16933), .S(P3_REIP_REG_25__SCAN_IN), .Z(
        n16942) );
  NOR2_X1 U20229 ( .A1(n16935), .A2(n17216), .ZN(n16951) );
  OAI21_X1 U20230 ( .B1(n17216), .B2(n16936), .A(n17209), .ZN(n16940) );
  AOI211_X1 U20231 ( .C1(n16938), .C2(n16937), .A(n9784), .B(n17176), .ZN(
        n16939) );
  AOI221_X1 U20232 ( .B1(n16951), .B2(n17228), .C1(n16940), .C2(
        P3_EBX_REG_25__SCAN_IN), .A(n16939), .ZN(n16941) );
  OAI211_X1 U20233 ( .C1(n16943), .C2(n17206), .A(n16942), .B(n16941), .ZN(
        P3_U2646) );
  INV_X1 U20234 ( .A(n16944), .ZN(n16945) );
  AOI211_X1 U20235 ( .C1(n17870), .C2(n16946), .A(n16945), .B(n17176), .ZN(
        n16948) );
  OAI22_X1 U20236 ( .A1(n17874), .A2(n17206), .B1(n17209), .B2(n16952), .ZN(
        n16947) );
  AOI211_X1 U20237 ( .C1(n16950), .C2(n16949), .A(n16948), .B(n16947), .ZN(
        n16955) );
  OAI21_X1 U20238 ( .B1(n16953), .B2(n16952), .A(n16951), .ZN(n16954) );
  OAI211_X1 U20239 ( .C1(n16967), .C2(n19112), .A(n16955), .B(n16954), .ZN(
        P3_U2647) );
  INV_X1 U20240 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n19111) );
  AOI211_X1 U20241 ( .C1(n17885), .C2(n16957), .A(n16956), .B(n17176), .ZN(
        n16961) );
  NAND2_X1 U20242 ( .A1(n17165), .A2(n16958), .ZN(n16959) );
  OAI22_X1 U20243 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(n16959), .B1(n16963), 
        .B2(n17209), .ZN(n16960) );
  AOI211_X1 U20244 ( .C1(n17192), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16961), .B(n16960), .ZN(n16966) );
  OAI211_X1 U20245 ( .C1(n16964), .C2(n16963), .A(n17219), .B(n16962), .ZN(
        n16965) );
  OAI211_X1 U20246 ( .C1(n16967), .C2(n19111), .A(n16966), .B(n16965), .ZN(
        P3_U2648) );
  AOI211_X1 U20247 ( .C1(n16970), .C2(n16969), .A(n16968), .B(n17176), .ZN(
        n16976) );
  OAI211_X1 U20248 ( .C1(n16972), .C2(n16974), .A(n17219), .B(n16971), .ZN(
        n16973) );
  OAI21_X1 U20249 ( .B1(n16974), .B2(n17209), .A(n16973), .ZN(n16975) );
  AOI211_X1 U20250 ( .C1(n17192), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16976), .B(n16975), .ZN(n16977) );
  OAI221_X1 U20251 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16979), .C1(n19107), 
        .C2(n16978), .A(n16977), .ZN(P3_U2650) );
  AOI22_X1 U20252 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17192), .B1(
        n17220), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n16992) );
  NAND2_X1 U20253 ( .A1(n16980), .A2(n17221), .ZN(n17041) );
  NOR2_X1 U20254 ( .A1(n16981), .A2(n17041), .ZN(n17009) );
  AOI21_X1 U20255 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n17009), .A(n17010), 
        .ZN(n16999) );
  INV_X1 U20256 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n19100) );
  NOR3_X1 U20257 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n19100), .A3(n16982), 
        .ZN(n16987) );
  OAI21_X1 U20258 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16983), .A(
        n17905), .ZN(n17944) );
  INV_X1 U20259 ( .A(n17944), .ZN(n16985) );
  AOI221_X1 U20260 ( .B1(n16985), .B2(n16984), .C1(n17944), .C2(n16995), .A(
        n17176), .ZN(n16986) );
  AOI211_X1 U20261 ( .C1(n16999), .C2(P3_REIP_REG_19__SCAN_IN), .A(n16987), 
        .B(n16986), .ZN(n16991) );
  OAI211_X1 U20262 ( .C1(n16996), .C2(n16989), .A(n17219), .B(n16988), .ZN(
        n16990) );
  NAND4_X1 U20263 ( .A1(n16992), .A2(n16991), .A3(n18482), .A4(n16990), .ZN(
        P3_U2652) );
  AOI21_X1 U20264 ( .B1(n17220), .B2(P3_EBX_REG_18__SCAN_IN), .A(n18349), .ZN(
        n17003) );
  OAI21_X1 U20265 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17940), .A(
        n16993), .ZN(n17952) );
  NOR2_X1 U20266 ( .A1(n17176), .A2(n17205), .ZN(n17138) );
  INV_X1 U20267 ( .A(n17138), .ZN(n17202) );
  INV_X1 U20268 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17955) );
  OAI221_X1 U20269 ( .B1(n17952), .B2(n17005), .C1(n17952), .C2(n17955), .A(
        n19045), .ZN(n16994) );
  AOI22_X1 U20270 ( .A1(n16995), .A2(n17952), .B1(n17202), .B2(n16994), .ZN(
        n16998) );
  AOI211_X1 U20271 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n17011), .A(n16996), .B(
        n17216), .ZN(n16997) );
  AOI211_X1 U20272 ( .C1(n17192), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16998), .B(n16997), .ZN(n17002) );
  OAI21_X1 U20273 ( .B1(P3_REIP_REG_18__SCAN_IN), .B2(n17000), .A(n16999), 
        .ZN(n17001) );
  NAND3_X1 U20274 ( .A1(n17003), .A2(n17002), .A3(n17001), .ZN(P3_U2653) );
  INV_X1 U20275 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17004) );
  AND2_X1 U20276 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17963), .ZN(
        n17007) );
  AOI21_X1 U20277 ( .B1(n17004), .B2(n17028), .A(n17007), .ZN(n17023) );
  INV_X1 U20278 ( .A(n17023), .ZN(n17985) );
  AOI21_X1 U20279 ( .B1(n17005), .B2(n17985), .A(n17175), .ZN(n17008) );
  INV_X1 U20280 ( .A(n17940), .ZN(n17006) );
  OAI21_X1 U20281 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17007), .A(
        n17006), .ZN(n17966) );
  XOR2_X1 U20282 ( .A(n17008), .B(n17966), .Z(n17018) );
  INV_X1 U20283 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n19099) );
  NOR3_X1 U20284 ( .A1(n17010), .A2(n17009), .A3(n19099), .ZN(n17015) );
  OAI211_X1 U20285 ( .C1(n17019), .C2(n17013), .A(n17219), .B(n17011), .ZN(
        n17012) );
  OAI211_X1 U20286 ( .C1(n17209), .C2(n17013), .A(n18482), .B(n17012), .ZN(
        n17014) );
  AOI211_X1 U20287 ( .C1(n17192), .C2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n17015), .B(n17014), .ZN(n17017) );
  NAND4_X1 U20288 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(n17033), .A4(n19099), .ZN(n17016) );
  OAI211_X1 U20289 ( .C1(n17018), .C2(n17176), .A(n17017), .B(n17016), .ZN(
        P3_U2654) );
  AOI211_X1 U20290 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n17034), .A(n17019), .B(
        n17216), .ZN(n17020) );
  AOI211_X1 U20291 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n17192), .A(
        n18349), .B(n17020), .ZN(n17027) );
  AND2_X1 U20292 ( .A1(n17218), .A2(n17041), .ZN(n17043) );
  INV_X1 U20293 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n19096) );
  INV_X1 U20294 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n19094) );
  AOI221_X1 U20295 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n19096), .C2(n19094), .A(n17021), .ZN(n17025) );
  AOI221_X1 U20296 ( .B1(n17030), .B2(n17023), .C1(n17022), .C2(n17985), .A(
        n17176), .ZN(n17024) );
  AOI211_X1 U20297 ( .C1(n17043), .C2(P3_REIP_REG_16__SCAN_IN), .A(n17025), 
        .B(n17024), .ZN(n17026) );
  OAI211_X1 U20298 ( .C1(n17209), .C2(n17400), .A(n17027), .B(n17026), .ZN(
        P3_U2655) );
  OAI21_X1 U20299 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17978), .A(
        n17028), .ZN(n17999) );
  AOI21_X1 U20300 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17202), .A(
        n17999), .ZN(n17029) );
  INV_X1 U20301 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n17208) );
  OAI21_X1 U20302 ( .B1(n17175), .B2(n17208), .A(n19045), .ZN(n17051) );
  INV_X1 U20303 ( .A(n17051), .ZN(n17212) );
  AOI22_X1 U20304 ( .A1(n17220), .A2(P3_EBX_REG_15__SCAN_IN), .B1(n17029), 
        .B2(n17212), .ZN(n17037) );
  INV_X1 U20305 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17995) );
  NAND3_X1 U20306 ( .A1(n17030), .A2(n19045), .A3(n17999), .ZN(n17031) );
  OAI211_X1 U20307 ( .C1(n17995), .C2(n17206), .A(n18482), .B(n17031), .ZN(
        n17032) );
  AOI221_X1 U20308 ( .B1(n17043), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n17033), 
        .C2(n19094), .A(n17032), .ZN(n17036) );
  OAI211_X1 U20309 ( .C1(n17038), .C2(n17397), .A(n17219), .B(n17034), .ZN(
        n17035) );
  NAND3_X1 U20310 ( .A1(n17037), .A2(n17036), .A3(n17035), .ZN(P3_U2656) );
  AOI211_X1 U20311 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n17055), .A(n17038), .B(
        n17216), .ZN(n17039) );
  AOI21_X1 U20312 ( .B1(n17192), .B2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n17039), .ZN(n17047) );
  NOR2_X1 U20313 ( .A1(n17210), .A2(n17040), .ZN(n17042) );
  AOI22_X1 U20314 ( .A1(n17220), .A2(P3_EBX_REG_14__SCAN_IN), .B1(n17042), 
        .B2(n17041), .ZN(n17046) );
  OR2_X1 U20315 ( .A1(n18021), .A2(n18018), .ZN(n17048) );
  AOI21_X1 U20316 ( .B1(n18008), .B2(n17048), .A(n17978), .ZN(n18010) );
  OAI21_X1 U20317 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17048), .A(
        n17205), .ZN(n17049) );
  XNOR2_X1 U20318 ( .A(n18010), .B(n17049), .ZN(n17044) );
  AOI22_X1 U20319 ( .A1(n19045), .A2(n17044), .B1(P3_REIP_REG_14__SCAN_IN), 
        .B2(n17043), .ZN(n17045) );
  NAND4_X1 U20320 ( .A1(n17047), .A2(n17046), .A3(n17045), .A4(n18482), .ZN(
        P3_U2657) );
  AOI22_X1 U20321 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17192), .B1(
        n17220), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n17060) );
  AOI21_X1 U20322 ( .B1(n17165), .B2(n17067), .A(n17204), .ZN(n17077) );
  NAND2_X1 U20323 ( .A1(n17165), .A2(n19088), .ZN(n17066) );
  INV_X1 U20324 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n19090) );
  AOI21_X1 U20325 ( .B1(n17077), .B2(n17066), .A(n19090), .ZN(n17054) );
  INV_X1 U20326 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17068) );
  NOR2_X1 U20327 ( .A1(n17068), .A2(n18018), .ZN(n17063) );
  OAI21_X1 U20328 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17063), .A(
        n17048), .ZN(n18023) );
  INV_X1 U20329 ( .A(n18023), .ZN(n17050) );
  NOR3_X1 U20330 ( .A1(n17050), .A2(n17176), .A3(n17049), .ZN(n17053) );
  AOI211_X1 U20331 ( .C1(n9724), .C2(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n17051), .B(n18023), .ZN(n17052) );
  NOR4_X1 U20332 ( .A1(n18499), .A2(n17054), .A3(n17053), .A4(n17052), .ZN(
        n17059) );
  OAI211_X1 U20333 ( .C1(n17061), .C2(n17395), .A(n17219), .B(n17055), .ZN(
        n17058) );
  NAND3_X1 U20334 ( .A1(n17165), .A2(n17056), .A3(n19090), .ZN(n17057) );
  NAND4_X1 U20335 ( .A1(n17060), .A2(n17059), .A3(n17058), .A4(n17057), .ZN(
        P3_U2658) );
  AOI211_X1 U20336 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17080), .A(n17061), .B(
        n17216), .ZN(n17062) );
  AOI21_X1 U20337 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17220), .A(n17062), .ZN(
        n17072) );
  AOI21_X1 U20338 ( .B1(n17068), .B2(n18018), .A(n17063), .ZN(n18035) );
  NAND2_X1 U20339 ( .A1(n17208), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17085) );
  INV_X1 U20340 ( .A(n17085), .ZN(n17199) );
  NAND3_X1 U20341 ( .A1(n18082), .A2(n17064), .A3(n17199), .ZN(n17074) );
  OAI21_X1 U20342 ( .B1(n18045), .B2(n17074), .A(n9724), .ZN(n17065) );
  XNOR2_X1 U20343 ( .A(n18035), .B(n17065), .ZN(n17070) );
  OAI22_X1 U20344 ( .A1(n17068), .A2(n17206), .B1(n17067), .B2(n17066), .ZN(
        n17069) );
  AOI211_X1 U20345 ( .C1(n19045), .C2(n17070), .A(n18349), .B(n17069), .ZN(
        n17071) );
  OAI211_X1 U20346 ( .C1(n19088), .C2(n17077), .A(n17072), .B(n17071), .ZN(
        P3_U2659) );
  AOI21_X1 U20347 ( .B1(n17165), .B2(n17073), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n17078) );
  OAI21_X1 U20348 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17084), .A(
        n18018), .ZN(n18046) );
  NAND2_X1 U20349 ( .A1(n9724), .A2(n17074), .ZN(n17075) );
  XNOR2_X1 U20350 ( .A(n18046), .B(n17075), .ZN(n17076) );
  OAI22_X1 U20351 ( .A1(n17078), .A2(n17077), .B1(n17176), .B2(n17076), .ZN(
        n17079) );
  AOI211_X1 U20352 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n17192), .A(
        n18349), .B(n17079), .ZN(n17082) );
  OAI211_X1 U20353 ( .C1(n17087), .C2(n17083), .A(n17219), .B(n17080), .ZN(
        n17081) );
  OAI211_X1 U20354 ( .C1(n17083), .C2(n17209), .A(n17082), .B(n17081), .ZN(
        P3_U2660) );
  INV_X1 U20355 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17154) );
  NAND3_X1 U20356 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17155), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17156) );
  NOR2_X1 U20357 ( .A1(n17154), .A2(n17156), .ZN(n17146) );
  NAND2_X1 U20358 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17146), .ZN(
        n17135) );
  NOR2_X1 U20359 ( .A1(n18083), .A2(n17135), .ZN(n17111) );
  NAND2_X1 U20360 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17111), .ZN(
        n17099) );
  AOI21_X1 U20361 ( .B1(n18058), .B2(n17099), .A(n17084), .ZN(n18063) );
  INV_X1 U20362 ( .A(n18082), .ZN(n18097) );
  OAI21_X1 U20363 ( .B1(n18097), .B2(n17085), .A(n9724), .ZN(n17130) );
  INV_X1 U20364 ( .A(n17130), .ZN(n17136) );
  AOI21_X1 U20365 ( .B1(n9724), .B2(n18083), .A(n17136), .ZN(n17100) );
  OAI21_X1 U20366 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17175), .A(
        n17100), .ZN(n17086) );
  XNOR2_X1 U20367 ( .A(n18063), .B(n17086), .ZN(n17096) );
  AOI211_X1 U20368 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17103), .A(n17087), .B(
        n17216), .ZN(n17088) );
  AOI211_X1 U20369 ( .C1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n17192), .A(
        n18349), .B(n17088), .ZN(n17095) );
  OAI21_X1 U20370 ( .B1(n17210), .B2(n17089), .A(n17221), .ZN(n17115) );
  INV_X1 U20371 ( .A(n17115), .ZN(n17090) );
  INV_X1 U20372 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n19082) );
  NAND3_X1 U20373 ( .A1(n17165), .A2(n17089), .A3(n19082), .ZN(n17107) );
  AOI21_X1 U20374 ( .B1(n17090), .B2(n17107), .A(n19084), .ZN(n17093) );
  NOR3_X1 U20375 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n17210), .A3(n17091), 
        .ZN(n17092) );
  AOI211_X1 U20376 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n17220), .A(n17093), .B(
        n17092), .ZN(n17094) );
  OAI211_X1 U20377 ( .C1(n17176), .C2(n17096), .A(n17095), .B(n17094), .ZN(
        P3_U2661) );
  OAI22_X1 U20378 ( .A1(n17097), .A2(n17206), .B1(n17209), .B2(n17104), .ZN(
        n17098) );
  AOI211_X1 U20379 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n17115), .A(n18349), .B(
        n17098), .ZN(n17108) );
  OAI21_X1 U20380 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17111), .A(
        n17099), .ZN(n18073) );
  INV_X1 U20381 ( .A(n18073), .ZN(n17102) );
  INV_X1 U20382 ( .A(n17100), .ZN(n17101) );
  OAI221_X1 U20383 ( .B1(n17102), .B2(n17101), .C1(n18073), .C2(n17100), .A(
        n19045), .ZN(n17106) );
  OAI211_X1 U20384 ( .C1(n17109), .C2(n17104), .A(n17219), .B(n17103), .ZN(
        n17105) );
  NAND4_X1 U20385 ( .A1(n17108), .A2(n17107), .A3(n17106), .A4(n17105), .ZN(
        P3_U2662) );
  AOI211_X1 U20386 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17124), .A(n17109), .B(
        n17216), .ZN(n17110) );
  AOI211_X1 U20387 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17192), .A(
        n18349), .B(n17110), .ZN(n17120) );
  INV_X1 U20388 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n18098) );
  NOR3_X1 U20389 ( .A1(n18169), .A2(n18097), .A3(n18098), .ZN(n17129) );
  INV_X1 U20390 ( .A(n17111), .ZN(n17112) );
  OAI21_X1 U20391 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17129), .A(
        n17112), .ZN(n18086) );
  AOI21_X1 U20392 ( .B1(n17129), .B2(n17208), .A(n17175), .ZN(n17113) );
  XNOR2_X1 U20393 ( .A(n18086), .B(n17113), .ZN(n17118) );
  NAND3_X1 U20394 ( .A1(n17165), .A2(P3_REIP_REG_5__SCAN_IN), .A3(n17145), 
        .ZN(n17144) );
  NOR2_X1 U20395 ( .A1(n17114), .A2(n17144), .ZN(n17116) );
  MUX2_X1 U20396 ( .A(n17116), .B(n17115), .S(P3_REIP_REG_8__SCAN_IN), .Z(
        n17117) );
  AOI21_X1 U20397 ( .B1(n17118), .B2(n19045), .A(n17117), .ZN(n17119) );
  OAI211_X1 U20398 ( .C1(n17209), .C2(n17121), .A(n17120), .B(n17119), .ZN(
        P3_U2663) );
  AOI21_X1 U20399 ( .B1(n17165), .B2(n17122), .A(n17204), .ZN(n17149) );
  AOI211_X1 U20400 ( .C1(n19078), .C2(n19076), .A(n17123), .B(n17144), .ZN(
        n17128) );
  OAI211_X1 U20401 ( .C1(n17134), .C2(n17126), .A(n17219), .B(n17124), .ZN(
        n17125) );
  OAI211_X1 U20402 ( .C1(n17209), .C2(n17126), .A(n18482), .B(n17125), .ZN(
        n17127) );
  AOI211_X1 U20403 ( .C1(n17192), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n17128), .B(n17127), .ZN(n17133) );
  AOI21_X1 U20404 ( .B1(n18098), .B2(n17135), .A(n17129), .ZN(n18103) );
  INV_X1 U20405 ( .A(n18103), .ZN(n17131) );
  OAI221_X1 U20406 ( .B1(n18103), .B2(n17136), .C1(n17131), .C2(n17130), .A(
        n19045), .ZN(n17132) );
  OAI211_X1 U20407 ( .C1(n17149), .C2(n19078), .A(n17133), .B(n17132), .ZN(
        P3_U2664) );
  AOI211_X1 U20408 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n17151), .A(n17134), .B(
        n17216), .ZN(n17142) );
  OAI21_X1 U20409 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17146), .A(
        n17135), .ZN(n18114) );
  NAND3_X1 U20410 ( .A1(n19045), .A2(n17136), .A3(n18114), .ZN(n17137) );
  OAI211_X1 U20411 ( .C1(n18113), .C2(n17206), .A(n18482), .B(n17137), .ZN(
        n17141) );
  OAI21_X1 U20412 ( .B1(n17138), .B2(n18113), .A(n17212), .ZN(n17139) );
  OAI22_X1 U20413 ( .A1(n17209), .A2(n17528), .B1(n18114), .B2(n17139), .ZN(
        n17140) );
  NOR3_X1 U20414 ( .A1(n17142), .A2(n17141), .A3(n17140), .ZN(n17143) );
  OAI221_X1 U20415 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n17144), .C1(n19076), 
        .C2(n17149), .A(n17143), .ZN(P3_U2665) );
  AOI21_X1 U20416 ( .B1(n17165), .B2(n17145), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n17148) );
  AOI21_X1 U20417 ( .B1(n17154), .B2(n17156), .A(n17146), .ZN(n18125) );
  OAI21_X1 U20418 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17156), .A(
        n9724), .ZN(n17158) );
  XOR2_X1 U20419 ( .A(n18125), .B(n17158), .Z(n17147) );
  OAI22_X1 U20420 ( .A1(n17149), .A2(n17148), .B1(n17176), .B2(n17147), .ZN(
        n17150) );
  AOI211_X1 U20421 ( .C1(n17220), .C2(P3_EBX_REG_5__SCAN_IN), .A(n18349), .B(
        n17150), .ZN(n17153) );
  OAI211_X1 U20422 ( .C1(n17166), .C2(n17532), .A(n17219), .B(n17151), .ZN(
        n17152) );
  OAI211_X1 U20423 ( .C1(n17206), .C2(n17154), .A(n17153), .B(n17152), .ZN(
        P3_U2666) );
  NOR2_X1 U20424 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18132), .ZN(
        n17161) );
  NAND2_X1 U20425 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17155), .ZN(
        n17173) );
  INV_X1 U20426 ( .A(n17173), .ZN(n17157) );
  OAI21_X1 U20427 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17157), .A(
        n17156), .ZN(n18141) );
  INV_X1 U20428 ( .A(n18141), .ZN(n17159) );
  OAI221_X1 U20429 ( .B1(n17159), .B2(n17158), .C1(n18141), .C2(n17205), .A(
        n18482), .ZN(n17160) );
  AOI21_X1 U20430 ( .B1(n17161), .B2(n17199), .A(n17160), .ZN(n17171) );
  NAND2_X1 U20431 ( .A1(n18517), .A2(n19202), .ZN(n17191) );
  AOI22_X1 U20432 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17192), .B1(
        n17220), .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n17162) );
  OAI221_X1 U20433 ( .B1(n9672), .B2(n17191), .C1(n18976), .C2(n17191), .A(
        n17162), .ZN(n17163) );
  INV_X1 U20434 ( .A(n17163), .ZN(n17170) );
  NOR2_X1 U20435 ( .A1(n17210), .A2(n17164), .ZN(n17168) );
  NAND2_X1 U20436 ( .A1(n17165), .A2(n17164), .ZN(n17182) );
  NAND2_X1 U20437 ( .A1(n17221), .A2(n17182), .ZN(n17184) );
  AOI211_X1 U20438 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n17185), .A(n17166), .B(
        n17216), .ZN(n17167) );
  AOI221_X1 U20439 ( .B1(n17168), .B2(n19072), .C1(n17184), .C2(
        P3_REIP_REG_4__SCAN_IN), .A(n17167), .ZN(n17169) );
  OAI211_X1 U20440 ( .C1(n17172), .C2(n17171), .A(n17170), .B(n17169), .ZN(
        P3_U2667) );
  INV_X1 U20441 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n19067) );
  INV_X1 U20442 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n19068) );
  NOR2_X1 U20443 ( .A1(n19067), .A2(n19068), .ZN(n17190) );
  INV_X1 U20444 ( .A(n17190), .ZN(n17181) );
  INV_X1 U20445 ( .A(n17191), .ZN(n17217) );
  NAND2_X1 U20446 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18984), .ZN(
        n18986) );
  AOI21_X1 U20447 ( .B1(n10936), .B2(n18986), .A(n9670), .ZN(n19139) );
  AOI22_X1 U20448 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n17192), .B1(
        n17217), .B2(n19139), .ZN(n17180) );
  INV_X1 U20449 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n18163) );
  NOR2_X1 U20450 ( .A1(n18169), .A2(n18163), .ZN(n17174) );
  OAI21_X1 U20451 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17174), .A(
        n17173), .ZN(n18153) );
  AOI21_X1 U20452 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17199), .A(
        n17175), .ZN(n17198) );
  INV_X1 U20453 ( .A(n17198), .ZN(n17178) );
  AOI21_X1 U20454 ( .B1(n18153), .B2(n17178), .A(n17176), .ZN(n17177) );
  OAI21_X1 U20455 ( .B1(n18153), .B2(n17178), .A(n17177), .ZN(n17179) );
  OAI211_X1 U20456 ( .C1(n17182), .C2(n17181), .A(n17180), .B(n17179), .ZN(
        n17183) );
  AOI21_X1 U20457 ( .B1(P3_REIP_REG_3__SCAN_IN), .B2(n17184), .A(n17183), .ZN(
        n17187) );
  OAI211_X1 U20458 ( .C1(n17188), .C2(n17527), .A(n17219), .B(n17185), .ZN(
        n17186) );
  OAI211_X1 U20459 ( .C1(n17527), .C2(n17209), .A(n17187), .B(n17186), .ZN(
        P3_U2668) );
  AOI22_X1 U20460 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18163), .B1(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18169), .ZN(n18159) );
  INV_X1 U20461 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17558) );
  INV_X1 U20462 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17553) );
  NAND2_X1 U20463 ( .A1(n17558), .A2(n17553), .ZN(n17189) );
  AOI211_X1 U20464 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n17189), .A(n17188), .B(
        n17216), .ZN(n17197) );
  AOI211_X1 U20465 ( .C1(n19067), .C2(n19068), .A(n17190), .B(n17210), .ZN(
        n17196) );
  INV_X1 U20466 ( .A(n18984), .ZN(n18990) );
  NAND2_X1 U20467 ( .A1(n18989), .A2(n10935), .ZN(n18983) );
  OAI21_X1 U20468 ( .B1(n18990), .B2(n9715), .A(n18983), .ZN(n19148) );
  OAI22_X1 U20469 ( .A1(n19068), .A2(n17221), .B1(n19148), .B2(n17191), .ZN(
        n17195) );
  AOI22_X1 U20470 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n17192), .B1(
        n17220), .B2(P3_EBX_REG_2__SCAN_IN), .ZN(n17193) );
  INV_X1 U20471 ( .A(n17193), .ZN(n17194) );
  NOR4_X1 U20472 ( .A1(n17197), .A2(n17196), .A3(n17195), .A4(n17194), .ZN(
        n17201) );
  OAI211_X1 U20473 ( .C1(n17199), .C2(n18159), .A(n19045), .B(n17198), .ZN(
        n17200) );
  OAI211_X1 U20474 ( .C1(n17202), .C2(n18159), .A(n17201), .B(n17200), .ZN(
        P3_U2669) );
  NOR2_X1 U20475 ( .A1(n17558), .A2(n17553), .ZN(n17547) );
  AOI21_X1 U20476 ( .B1(n17558), .B2(n17553), .A(n17547), .ZN(n17203) );
  INV_X1 U20477 ( .A(n17203), .ZN(n17554) );
  NAND2_X1 U20478 ( .A1(n18989), .A2(n10931), .ZN(n19006) );
  INV_X1 U20479 ( .A(n19006), .ZN(n19157) );
  AOI22_X1 U20480 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17204), .B1(n19157), 
        .B2(n17217), .ZN(n17215) );
  NAND2_X1 U20481 ( .A1(n17205), .A2(n19045), .ZN(n17207) );
  OAI21_X1 U20482 ( .B1(n17208), .B2(n17207), .A(n17206), .ZN(n17213) );
  OAI22_X1 U20483 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n17210), .B1(n17209), 
        .B2(n17553), .ZN(n17211) );
  AOI221_X1 U20484 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17213), .C1(
        n18169), .C2(n17212), .A(n17211), .ZN(n17214) );
  OAI211_X1 U20485 ( .C1(n17216), .C2(n17554), .A(n17215), .B(n17214), .ZN(
        P3_U2670) );
  AOI22_X1 U20486 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n17218), .B1(n17217), 
        .B2(n9998), .ZN(n17224) );
  OAI21_X1 U20487 ( .B1(n17220), .B2(n17219), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n17223) );
  NAND3_X1 U20488 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n19150), .A3(
        n17221), .ZN(n17222) );
  NAND3_X1 U20489 ( .A1(n17224), .A2(n17223), .A3(n17222), .ZN(P3_U2671) );
  NOR2_X1 U20490 ( .A1(n17226), .A2(n17225), .ZN(n17309) );
  NAND4_X1 U20491 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n17269), .A4(n17309), .ZN(n17227) );
  NOR3_X1 U20492 ( .A1(n17280), .A2(n17228), .A3(n17227), .ZN(n17229) );
  NAND4_X1 U20493 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(n17229), .ZN(n17232) );
  NAND2_X1 U20494 ( .A1(n17551), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17231) );
  NAND2_X1 U20495 ( .A1(n17262), .A2(n18548), .ZN(n17230) );
  OAI22_X1 U20496 ( .A1(n17262), .A2(n17231), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17230), .ZN(P3_U2672) );
  NAND2_X1 U20497 ( .A1(n17233), .A2(n17232), .ZN(n17234) );
  NAND2_X1 U20498 ( .A1(n17234), .A2(n17551), .ZN(n17261) );
  AOI22_X1 U20499 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9670), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17235) );
  OAI21_X1 U20500 ( .B1(n11006), .B2(n17418), .A(n17235), .ZN(n17244) );
  AOI22_X1 U20501 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17242) );
  INV_X1 U20502 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17304) );
  OAI22_X1 U20503 ( .A1(n17472), .A2(n18764), .B1(n10978), .B2(n17304), .ZN(
        n17240) );
  AOI22_X1 U20504 ( .A1(n17476), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17238) );
  AOI22_X1 U20505 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17237) );
  AOI22_X1 U20506 ( .A1(n17512), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17236) );
  NAND3_X1 U20507 ( .A1(n17238), .A2(n17237), .A3(n17236), .ZN(n17239) );
  AOI211_X1 U20508 ( .C1(n17520), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n17240), .B(n17239), .ZN(n17241) );
  OAI211_X1 U20509 ( .C1(n17256), .C2(n17419), .A(n17242), .B(n17241), .ZN(
        n17243) );
  AOI211_X1 U20510 ( .C1(n16175), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n17244), .B(n17243), .ZN(n17245) );
  INV_X1 U20511 ( .A(n17245), .ZN(n17265) );
  NAND3_X1 U20512 ( .A1(n17264), .A2(n17263), .A3(n17265), .ZN(n17260) );
  AOI22_X1 U20513 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n17490), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n17476), .ZN(n17246) );
  OAI21_X1 U20514 ( .B1(n10109), .B2(n17247), .A(n17246), .ZN(n17258) );
  AOI22_X1 U20515 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17520), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17255) );
  OAI22_X1 U20516 ( .A1(n17248), .A2(n10978), .B1(n17472), .B2(n18770), .ZN(
        n17253) );
  AOI22_X1 U20517 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17456), .ZN(n17251) );
  AOI22_X1 U20518 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9671), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17250) );
  AOI22_X1 U20519 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n11129), .B1(
        n17512), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17249) );
  NAND3_X1 U20520 ( .A1(n17251), .A2(n17250), .A3(n17249), .ZN(n17252) );
  AOI211_X1 U20521 ( .C1(n17421), .C2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A(
        n17253), .B(n17252), .ZN(n17254) );
  OAI211_X1 U20522 ( .C1(n17256), .C2(n17412), .A(n17255), .B(n17254), .ZN(
        n17257) );
  AOI211_X1 U20523 ( .C1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .C2(n17494), .A(
        n17258), .B(n17257), .ZN(n17259) );
  XNOR2_X1 U20524 ( .A(n17260), .B(n17259), .ZN(n17568) );
  OAI22_X1 U20525 ( .A1(n17262), .A2(n17261), .B1(n17568), .B2(n17551), .ZN(
        P3_U2673) );
  NAND2_X1 U20526 ( .A1(n17264), .A2(n17263), .ZN(n17266) );
  XOR2_X1 U20527 ( .A(n17266), .B(n17265), .Z(n17576) );
  OAI21_X1 U20528 ( .B1(n17551), .B2(n17576), .A(n17271), .ZN(P3_U2674) );
  OAI21_X1 U20529 ( .B1(n17276), .B2(n17273), .A(n17272), .ZN(n17586) );
  NAND3_X1 U20530 ( .A1(n17275), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17551), 
        .ZN(n17274) );
  OAI221_X1 U20531 ( .B1(n17275), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17551), 
        .C2(n17586), .A(n17274), .ZN(P3_U2676) );
  AOI21_X1 U20532 ( .B1(n17277), .B2(n17282), .A(n17276), .ZN(n17587) );
  NAND2_X1 U20533 ( .A1(n17555), .A2(n17587), .ZN(n17278) );
  OAI221_X1 U20534 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17281), .C1(n17280), 
        .C2(n17279), .A(n17278), .ZN(P3_U2677) );
  AOI21_X1 U20535 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17551), .A(n17289), .ZN(
        n17285) );
  OAI21_X1 U20536 ( .B1(n17284), .B2(n17283), .A(n17282), .ZN(n17596) );
  OAI22_X1 U20537 ( .A1(n17286), .A2(n17285), .B1(n17551), .B2(n17596), .ZN(
        P3_U2678) );
  AOI21_X1 U20538 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17551), .A(n17295), .ZN(
        n17288) );
  XNOR2_X1 U20539 ( .A(n17287), .B(n17291), .ZN(n17602) );
  OAI22_X1 U20540 ( .A1(n17289), .A2(n17288), .B1(n17551), .B2(n17602), .ZN(
        P3_U2679) );
  AOI22_X1 U20541 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(n17551), .B1(
        P3_EBX_REG_22__SCAN_IN), .B2(n17290), .ZN(n17294) );
  OAI21_X1 U20542 ( .B1(n17293), .B2(n17292), .A(n17291), .ZN(n17608) );
  OAI22_X1 U20543 ( .A1(n17295), .A2(n17294), .B1(n17551), .B2(n17608), .ZN(
        P3_U2680) );
  AOI22_X1 U20544 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17296) );
  OAI21_X1 U20545 ( .B1(n10970), .B2(n17418), .A(n17296), .ZN(n17306) );
  AOI22_X1 U20546 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17303) );
  AOI22_X1 U20547 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17297) );
  OAI21_X1 U20548 ( .B1(n10109), .B2(n18764), .A(n17297), .ZN(n17301) );
  AOI22_X1 U20549 ( .A1(n17494), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10961), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17299) );
  AOI22_X1 U20550 ( .A1(n17508), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9671), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17298) );
  OAI211_X1 U20551 ( .C1(n10978), .C2(n17419), .A(n17299), .B(n17298), .ZN(
        n17300) );
  AOI211_X1 U20552 ( .C1(n17512), .C2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n17301), .B(n17300), .ZN(n17302) );
  OAI211_X1 U20553 ( .C1(n17511), .C2(n17304), .A(n17303), .B(n17302), .ZN(
        n17305) );
  AOI211_X1 U20554 ( .C1(n17421), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n17306), .B(n17305), .ZN(n17610) );
  NAND3_X1 U20555 ( .A1(n17308), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17551), 
        .ZN(n17307) );
  OAI221_X1 U20556 ( .B1(n17308), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17551), 
        .C2(n17610), .A(n17307), .ZN(P3_U2681) );
  NOR2_X1 U20557 ( .A1(n17555), .A2(n17309), .ZN(n17335) );
  AOI22_X1 U20558 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17495), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17321) );
  AOI22_X1 U20559 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17320) );
  OAI22_X1 U20560 ( .A1(n11006), .A2(n17310), .B1(n10948), .B2(n17537), .ZN(
        n17318) );
  AOI22_X1 U20561 ( .A1(n10981), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17512), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17316) );
  AOI22_X1 U20562 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17312) );
  AOI22_X1 U20563 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10961), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17311) );
  OAI211_X1 U20564 ( .C1(n10978), .C2(n17313), .A(n17312), .B(n17311), .ZN(
        n17314) );
  AOI21_X1 U20565 ( .B1(n11129), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n17314), .ZN(n17315) );
  OAI211_X1 U20566 ( .C1(n9672), .C2(n18589), .A(n17316), .B(n17315), .ZN(
        n17317) );
  NAND3_X1 U20567 ( .A1(n17321), .A2(n17320), .A3(n17319), .ZN(n17616) );
  AOI22_X1 U20568 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17335), .B1(n17555), 
        .B2(n17616), .ZN(n17322) );
  OAI21_X1 U20569 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17323), .A(n17322), .ZN(
        P3_U2682) );
  AOI22_X1 U20570 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17324) );
  OAI21_X1 U20571 ( .B1(n10109), .B2(n18758), .A(n17324), .ZN(n17334) );
  AOI22_X1 U20572 ( .A1(n10981), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17331) );
  OAI22_X1 U20573 ( .A1(n10949), .A2(n17437), .B1(n17474), .B2(n17540), .ZN(
        n17329) );
  AOI22_X1 U20574 ( .A1(n17508), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17494), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17327) );
  AOI22_X1 U20575 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17326) );
  AOI22_X1 U20576 ( .A1(n17512), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17514), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17325) );
  NAND3_X1 U20577 ( .A1(n17327), .A2(n17326), .A3(n17325), .ZN(n17328) );
  AOI211_X1 U20578 ( .C1(n9671), .C2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n17329), .B(n17328), .ZN(n17330) );
  OAI211_X1 U20579 ( .C1(n17511), .C2(n17332), .A(n17331), .B(n17330), .ZN(
        n17333) );
  AOI211_X1 U20580 ( .C1(n17421), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n17334), .B(n17333), .ZN(n17624) );
  OAI21_X1 U20581 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17336), .A(n17335), .ZN(
        n17337) );
  OAI21_X1 U20582 ( .B1(n17624), .B2(n17551), .A(n17337), .ZN(P3_U2683) );
  NAND2_X1 U20583 ( .A1(n18548), .A2(n17338), .ZN(n17351) );
  NOR2_X1 U20584 ( .A1(n17555), .A2(n17338), .ZN(n17366) );
  AOI22_X1 U20585 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17508), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17349) );
  AOI22_X1 U20586 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17348) );
  AOI22_X1 U20587 ( .A1(n17512), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17347) );
  OAI22_X1 U20588 ( .A1(n10948), .A2(n17544), .B1(n10978), .B2(n17452), .ZN(
        n17345) );
  AOI22_X1 U20589 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17520), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17343) );
  AOI22_X1 U20590 ( .A1(n17494), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9671), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17342) );
  AOI22_X1 U20591 ( .A1(n17476), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17341) );
  NAND2_X1 U20592 ( .A1(n17339), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n17340) );
  NAND4_X1 U20593 ( .A1(n17343), .A2(n17342), .A3(n17341), .A4(n17340), .ZN(
        n17344) );
  AOI211_X1 U20594 ( .C1(n17421), .C2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A(
        n17345), .B(n17344), .ZN(n17346) );
  NAND4_X1 U20595 ( .A1(n17349), .A2(n17348), .A3(n17347), .A4(n17346), .ZN(
        n17625) );
  AOI22_X1 U20596 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17366), .B1(n17555), 
        .B2(n17625), .ZN(n17350) );
  OAI21_X1 U20597 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17351), .A(n17350), .ZN(
        P3_U2684) );
  AOI22_X1 U20598 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17494), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17352) );
  OAI21_X1 U20599 ( .B1(n17511), .B2(n17353), .A(n17352), .ZN(n17364) );
  AOI22_X1 U20600 ( .A1(n10981), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17508), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17362) );
  AOI22_X1 U20601 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10961), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17354) );
  OAI21_X1 U20602 ( .B1(n17455), .B2(n17355), .A(n17354), .ZN(n17360) );
  AOI22_X1 U20603 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17357) );
  AOI22_X1 U20604 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9671), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17356) );
  OAI211_X1 U20605 ( .C1(n10978), .C2(n17358), .A(n17357), .B(n17356), .ZN(
        n17359) );
  AOI211_X1 U20606 ( .C1(n17512), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n17360), .B(n17359), .ZN(n17361) );
  OAI211_X1 U20607 ( .C1(n10970), .C2(n17471), .A(n17362), .B(n17361), .ZN(
        n17363) );
  AOI211_X1 U20608 ( .C1(n17421), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n17364), .B(n17363), .ZN(n17633) );
  NAND2_X1 U20609 ( .A1(n17365), .A2(n17369), .ZN(n17367) );
  NAND2_X1 U20610 ( .A1(n17367), .A2(n17366), .ZN(n17368) );
  OAI21_X1 U20611 ( .B1(n17633), .B2(n17551), .A(n17368), .ZN(P3_U2685) );
  INV_X1 U20612 ( .A(n17369), .ZN(n17383) );
  AOI22_X1 U20613 ( .A1(n18548), .A2(n17370), .B1(P3_EBX_REG_17__SCAN_IN), 
        .B2(n17551), .ZN(n17382) );
  AOI22_X1 U20614 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17371) );
  OAI21_X1 U20615 ( .B1(n10109), .B2(n18749), .A(n17371), .ZN(n17381) );
  AOI22_X1 U20616 ( .A1(n17403), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17379) );
  OAI22_X1 U20617 ( .A1(n10946), .A2(n17372), .B1(n17472), .B2(n17493), .ZN(
        n17377) );
  AOI22_X1 U20618 ( .A1(n17456), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10961), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17375) );
  AOI22_X1 U20619 ( .A1(n17508), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17494), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17374) );
  AOI22_X1 U20620 ( .A1(n17512), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17514), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17373) );
  NAND3_X1 U20621 ( .A1(n17375), .A2(n17374), .A3(n17373), .ZN(n17376) );
  AOI211_X1 U20622 ( .C1(n17495), .C2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n17377), .B(n17376), .ZN(n17378) );
  OAI211_X1 U20623 ( .C1(n9672), .C2(n18579), .A(n17379), .B(n17378), .ZN(
        n17380) );
  AOI211_X1 U20624 ( .C1(n16175), .C2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A(
        n17381), .B(n17380), .ZN(n17641) );
  OAI22_X1 U20625 ( .A1(n17383), .A2(n17382), .B1(n17641), .B2(n17551), .ZN(
        P3_U2686) );
  NAND2_X1 U20626 ( .A1(n17551), .A2(n17384), .ZN(n17416) );
  AOI22_X1 U20627 ( .A1(n10981), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17494), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17394) );
  INV_X1 U20628 ( .A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17510) );
  AOI22_X1 U20629 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17420), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17386) );
  AOI22_X1 U20630 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17385) );
  OAI211_X1 U20631 ( .C1(n10978), .C2(n17510), .A(n17386), .B(n17385), .ZN(
        n17392) );
  AOI22_X1 U20632 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17508), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17390) );
  AOI22_X1 U20633 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17389) );
  AOI22_X1 U20634 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17388) );
  NAND2_X1 U20635 ( .A1(n11129), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n17387) );
  NAND4_X1 U20636 ( .A1(n17390), .A2(n17389), .A3(n17388), .A4(n17387), .ZN(
        n17391) );
  AOI211_X1 U20637 ( .C1(n17512), .C2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A(
        n17392), .B(n17391), .ZN(n17393) );
  OAI211_X1 U20638 ( .C1(n9672), .C2(n18576), .A(n17394), .B(n17393), .ZN(
        n17642) );
  NOR4_X1 U20639 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17397), .A3(n17396), .A4(
        n17395), .ZN(n17398) );
  AOI22_X1 U20640 ( .A1(n17555), .A2(n17642), .B1(n17447), .B2(n17398), .ZN(
        n17399) );
  OAI21_X1 U20641 ( .B1(n17400), .B2(n17416), .A(n17399), .ZN(P3_U2687) );
  AOI22_X1 U20642 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n17420), .B1(
        n17508), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17401) );
  OAI21_X1 U20643 ( .B1(n17402), .B2(n11006), .A(n17401), .ZN(n17414) );
  AOI22_X1 U20644 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n9667), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17490), .ZN(n17411) );
  INV_X1 U20645 ( .A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17405) );
  AOI22_X1 U20646 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17339), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17456), .ZN(n17404) );
  OAI21_X1 U20647 ( .B1(n17455), .B2(n17405), .A(n17404), .ZN(n17409) );
  AOI22_X1 U20648 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n9720), .ZN(n17407) );
  AOI22_X1 U20649 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17476), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n9670), .ZN(n17406) );
  OAI211_X1 U20650 ( .C1(n17460), .C2(n17529), .A(n17407), .B(n17406), .ZN(
        n17408) );
  AOI211_X1 U20651 ( .C1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .C2(n17514), .A(
        n17409), .B(n17408), .ZN(n17410) );
  OAI211_X1 U20652 ( .C1(n17511), .C2(n17412), .A(n17411), .B(n17410), .ZN(
        n17413) );
  AOI211_X1 U20653 ( .C1(n17421), .C2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A(
        n17414), .B(n17413), .ZN(n17652) );
  NOR2_X1 U20654 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17415), .ZN(n17417) );
  OAI22_X1 U20655 ( .A1(n17652), .A2(n17551), .B1(n17417), .B2(n17416), .ZN(
        P3_U2688) );
  OAI22_X1 U20656 ( .A1(n17555), .A2(n17447), .B1(P3_EBX_REG_13__SCAN_IN), 
        .B2(n17559), .ZN(n17432) );
  AOI22_X1 U20657 ( .A1(n11030), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17431) );
  AOI22_X1 U20658 ( .A1(n9671), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17430) );
  AOI22_X1 U20659 ( .A1(n17514), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17429) );
  OAI22_X1 U20660 ( .A1(n17511), .A2(n17419), .B1(n17472), .B2(n17418), .ZN(
        n17427) );
  AOI22_X1 U20661 ( .A1(n17494), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17425) );
  AOI22_X1 U20662 ( .A1(n17421), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17420), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17424) );
  AOI22_X1 U20663 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17403), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17423) );
  NAND2_X1 U20664 ( .A1(n17512), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n17422) );
  NAND4_X1 U20665 ( .A1(n17425), .A2(n17424), .A3(n17423), .A4(n17422), .ZN(
        n17426) );
  AOI211_X1 U20666 ( .C1(n17495), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(
        n17427), .B(n17426), .ZN(n17428) );
  NAND4_X1 U20667 ( .A1(n17431), .A2(n17430), .A3(n17429), .A4(n17428), .ZN(
        n17658) );
  AOI22_X1 U20668 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17432), .B1(n17555), 
        .B2(n17658), .ZN(n17433) );
  OAI21_X1 U20669 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17434), .A(n17433), .ZN(
        P3_U2689) );
  AOI22_X1 U20670 ( .A1(n9670), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17435) );
  OAI21_X1 U20671 ( .B1(n10949), .B2(n17436), .A(n17435), .ZN(n17446) );
  AOI22_X1 U20672 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17444) );
  OAI22_X1 U20673 ( .A1(n17460), .A2(n17540), .B1(n17474), .B2(n17437), .ZN(
        n17442) );
  AOI22_X1 U20674 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17508), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17440) );
  AOI22_X1 U20675 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17439) );
  AOI22_X1 U20676 ( .A1(n17514), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17438) );
  NAND3_X1 U20677 ( .A1(n17440), .A2(n17439), .A3(n17438), .ZN(n17441) );
  AOI211_X1 U20678 ( .C1(n17476), .C2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A(
        n17442), .B(n17441), .ZN(n17443) );
  OAI211_X1 U20679 ( .C1(n10946), .C2(n18758), .A(n17444), .B(n17443), .ZN(
        n17445) );
  AOI211_X1 U20680 ( .C1(n17494), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n17446), .B(n17445), .ZN(n17667) );
  INV_X1 U20681 ( .A(n17467), .ZN(n17449) );
  INV_X1 U20682 ( .A(n17447), .ZN(n17448) );
  OAI211_X1 U20683 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n17449), .A(n17448), .B(
        n17551), .ZN(n17450) );
  OAI21_X1 U20684 ( .B1(n17667), .B2(n17551), .A(n17450), .ZN(P3_U2691) );
  AOI22_X1 U20685 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10961), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17451) );
  OAI21_X1 U20686 ( .B1(n17511), .B2(n17452), .A(n17451), .ZN(n17466) );
  AOI22_X1 U20687 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9670), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17464) );
  INV_X1 U20688 ( .A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17454) );
  AOI22_X1 U20689 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17339), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17453) );
  OAI21_X1 U20690 ( .B1(n17455), .B2(n17454), .A(n17453), .ZN(n17462) );
  AOI22_X1 U20691 ( .A1(n17494), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17459) );
  AOI22_X1 U20692 ( .A1(n17508), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17457), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17458) );
  OAI211_X1 U20693 ( .C1(n17460), .C2(n17544), .A(n17459), .B(n17458), .ZN(
        n17461) );
  AOI211_X1 U20694 ( .C1(n17514), .C2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A(
        n17462), .B(n17461), .ZN(n17463) );
  OAI211_X1 U20695 ( .C1(n10946), .C2(n18755), .A(n17464), .B(n17463), .ZN(
        n17465) );
  AOI211_X1 U20696 ( .C1(n17495), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n17466), .B(n17465), .ZN(n17672) );
  OAI21_X1 U20697 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17468), .A(n17467), .ZN(
        n17469) );
  AOI22_X1 U20698 ( .A1(n17555), .A2(n17672), .B1(n17469), .B2(n17551), .ZN(
        P3_U2692) );
  NAND2_X1 U20699 ( .A1(n17551), .A2(n17486), .ZN(n17505) );
  AOI22_X1 U20700 ( .A1(n17470), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17508), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17485) );
  AOI22_X1 U20701 ( .A1(n17520), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17494), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17484) );
  OAI22_X1 U20702 ( .A1(n17472), .A2(n17471), .B1(n11128), .B2(n18582), .ZN(
        n17482) );
  OAI22_X1 U20703 ( .A1(n10946), .A2(n18752), .B1(n17474), .B2(n17473), .ZN(
        n17475) );
  AOI21_X1 U20704 ( .B1(n17514), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n17475), .ZN(n17480) );
  AOI22_X1 U20705 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17476), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17479) );
  AOI22_X1 U20706 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17478) );
  AOI22_X1 U20707 ( .A1(n17512), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17477) );
  NAND4_X1 U20708 ( .A1(n17480), .A2(n17479), .A3(n17478), .A4(n17477), .ZN(
        n17481) );
  AOI211_X1 U20709 ( .C1(n9670), .C2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A(
        n17482), .B(n17481), .ZN(n17483) );
  NAND3_X1 U20710 ( .A1(n17485), .A2(n17484), .A3(n17483), .ZN(n17676) );
  NOR3_X1 U20711 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17691), .A3(n17486), .ZN(
        n17487) );
  AOI21_X1 U20712 ( .B1(n17555), .B2(n17676), .A(n17487), .ZN(n17488) );
  OAI21_X1 U20713 ( .B1(n17489), .B2(n17505), .A(n17488), .ZN(P3_U2693) );
  AOI22_X1 U20714 ( .A1(n9671), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17491) );
  OAI21_X1 U20715 ( .B1(n11128), .B2(n18579), .A(n17491), .ZN(n17504) );
  AOI22_X1 U20716 ( .A1(n17403), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17514), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17502) );
  OAI22_X1 U20717 ( .A1(n10109), .A2(n17493), .B1(n10970), .B2(n17492), .ZN(
        n17500) );
  AOI22_X1 U20718 ( .A1(n11030), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17494), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17498) );
  AOI22_X1 U20719 ( .A1(n17495), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10961), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n17497) );
  AOI22_X1 U20720 ( .A1(n17512), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17496) );
  NAND3_X1 U20721 ( .A1(n17498), .A2(n17497), .A3(n17496), .ZN(n17499) );
  AOI211_X1 U20722 ( .C1(n10981), .C2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n17500), .B(n17499), .ZN(n17501) );
  OAI211_X1 U20723 ( .C1(n10946), .C2(n18749), .A(n17502), .B(n17501), .ZN(
        n17503) );
  AOI211_X1 U20724 ( .C1(n16175), .C2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A(
        n17504), .B(n17503), .ZN(n17680) );
  NOR2_X1 U20725 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n17526), .ZN(n17506) );
  OAI22_X1 U20726 ( .A1(n17680), .A2(n17551), .B1(n17506), .B2(n17505), .ZN(
        P3_U2694) );
  INV_X1 U20727 ( .A(n17507), .ZN(n17531) );
  OAI21_X1 U20728 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17531), .A(n17551), .ZN(
        n17525) );
  AOI22_X1 U20729 ( .A1(n17508), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17490), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17509) );
  OAI21_X1 U20730 ( .B1(n17511), .B2(n17510), .A(n17509), .ZN(n17524) );
  AOI22_X1 U20731 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9671), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17522) );
  AOI22_X1 U20732 ( .A1(n10981), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17512), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17513) );
  INV_X1 U20733 ( .A(n17513), .ZN(n17519) );
  AOI22_X1 U20734 ( .A1(n17494), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17456), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17517) );
  AOI22_X1 U20735 ( .A1(n17420), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10961), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17516) );
  AOI22_X1 U20736 ( .A1(n17514), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11129), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17515) );
  NAND3_X1 U20737 ( .A1(n17517), .A2(n17516), .A3(n17515), .ZN(n17518) );
  AOI211_X1 U20738 ( .C1(n17520), .C2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n17519), .B(n17518), .ZN(n17521) );
  OAI211_X1 U20739 ( .C1(n10946), .C2(n18746), .A(n17522), .B(n17521), .ZN(
        n17523) );
  AOI211_X1 U20740 ( .C1(n17495), .C2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n17524), .B(n17523), .ZN(n17686) );
  OAI22_X1 U20741 ( .A1(n17526), .A2(n17525), .B1(n17686), .B2(n17551), .ZN(
        P3_U2695) );
  NOR3_X1 U20742 ( .A1(n17527), .A2(n17543), .A3(n17559), .ZN(n17546) );
  NAND2_X1 U20743 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17546), .ZN(n17536) );
  NOR3_X1 U20744 ( .A1(n17528), .A2(n17532), .A3(n17536), .ZN(n17535) );
  AOI21_X1 U20745 ( .B1(P3_EBX_REG_7__SCAN_IN), .B2(n17551), .A(n17535), .ZN(
        n17530) );
  OAI22_X1 U20746 ( .A1(n17531), .A2(n17530), .B1(n17529), .B2(n17551), .ZN(
        P3_U2696) );
  NOR2_X1 U20747 ( .A1(n17532), .A2(n17536), .ZN(n17539) );
  AOI21_X1 U20748 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17551), .A(n17539), .ZN(
        n17534) );
  INV_X1 U20749 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17533) );
  OAI22_X1 U20750 ( .A1(n17535), .A2(n17534), .B1(n17533), .B2(n17551), .ZN(
        P3_U2697) );
  INV_X1 U20751 ( .A(n17536), .ZN(n17542) );
  AOI21_X1 U20752 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17551), .A(n17542), .ZN(
        n17538) );
  OAI22_X1 U20753 ( .A1(n17539), .A2(n17538), .B1(n17537), .B2(n17551), .ZN(
        P3_U2698) );
  AOI21_X1 U20754 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17551), .A(n17546), .ZN(
        n17541) );
  OAI22_X1 U20755 ( .A1(n17542), .A2(n17541), .B1(n17540), .B2(n17551), .ZN(
        P3_U2699) );
  NOR2_X1 U20756 ( .A1(n17543), .A2(n17559), .ZN(n17548) );
  AOI21_X1 U20757 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17551), .A(n17548), .ZN(
        n17545) );
  OAI22_X1 U20758 ( .A1(n17546), .A2(n17545), .B1(n17544), .B2(n17551), .ZN(
        P3_U2700) );
  INV_X1 U20759 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17550) );
  AOI211_X1 U20760 ( .C1(n17555), .C2(n17550), .A(n17549), .B(n17548), .ZN(
        P3_U2701) );
  INV_X1 U20761 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17552) );
  NAND2_X1 U20762 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17555), .ZN(
        n17556) );
  OAI221_X1 U20763 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17559), .C1(n17558), 
        .C2(n9732), .A(n17556), .ZN(P3_U2703) );
  NOR2_X1 U20764 ( .A1(n17722), .A2(n18542), .ZN(n17638) );
  INV_X1 U20765 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17789) );
  INV_X1 U20766 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17786) );
  INV_X1 U20767 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17784) );
  INV_X1 U20768 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17782) );
  INV_X1 U20769 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17768) );
  NAND4_X1 U20770 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .A4(P3_EAX_REG_10__SCAN_IN), .ZN(n17656)
         );
  NAND4_X1 U20771 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_2__SCAN_IN), 
        .A3(P3_EAX_REG_1__SCAN_IN), .A4(P3_EAX_REG_0__SCAN_IN), .ZN(n17561) );
  NAND4_X1 U20772 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_5__SCAN_IN), .A4(P3_EAX_REG_4__SCAN_IN), .ZN(n17560) );
  NOR2_X1 U20773 ( .A1(n17561), .A2(n17560), .ZN(n17655) );
  NAND4_X1 U20774 ( .A1(n17655), .A2(P3_EAX_REG_14__SCAN_IN), .A3(
        P3_EAX_REG_9__SCAN_IN), .A4(P3_EAX_REG_8__SCAN_IN), .ZN(n17562) );
  NOR3_X2 U20775 ( .A1(n17720), .A2(n17656), .A3(n17562), .ZN(n17659) );
  NAND2_X1 U20776 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n17659), .ZN(n17649) );
  NOR2_X2 U20777 ( .A1(n17768), .A2(n17649), .ZN(n17644) );
  INV_X1 U20778 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17778) );
  INV_X1 U20779 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17776) );
  INV_X1 U20780 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17774) );
  INV_X1 U20781 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17772) );
  NOR4_X1 U20782 ( .A1(n17778), .A2(n17776), .A3(n17774), .A4(n17772), .ZN(
        n17609) );
  NAND4_X1 U20783 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_17__SCAN_IN), 
        .A3(n17644), .A4(n17609), .ZN(n17604) );
  NAND2_X1 U20784 ( .A1(n18548), .A2(n17603), .ZN(n17597) );
  NAND2_X1 U20785 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17582), .ZN(n17578) );
  NAND2_X1 U20786 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17573), .ZN(n17572) );
  NOR2_X1 U20787 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n9712), .ZN(n17564) );
  NAND2_X1 U20788 ( .A1(n17722), .A2(n17572), .ZN(n17571) );
  OAI21_X1 U20789 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17653), .A(n17571), .ZN(
        n17563) );
  AOI22_X1 U20790 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17564), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17563), .ZN(n17565) );
  OAI21_X1 U20791 ( .B1(n17566), .B2(n17648), .A(n17565), .ZN(P3_U2704) );
  INV_X1 U20792 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17795) );
  NOR2_X2 U20793 ( .A1(n17567), .A2(n17722), .ZN(n17643) );
  INV_X1 U20794 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19558) );
  OAI22_X1 U20795 ( .A1(n17568), .A2(n17713), .B1(n19558), .B2(n17648), .ZN(
        n17569) );
  AOI21_X1 U20796 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17643), .A(n17569), .ZN(
        n17570) );
  OAI221_X1 U20797 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n9712), .C1(n17795), 
        .C2(n17571), .A(n17570), .ZN(P3_U2705) );
  AOI22_X1 U20798 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17643), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17638), .ZN(n17575) );
  OAI211_X1 U20799 ( .C1(n17573), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17722), .B(
        n9712), .ZN(n17574) );
  OAI211_X1 U20800 ( .C1(n17713), .C2(n17576), .A(n17575), .B(n17574), .ZN(
        P3_U2706) );
  INV_X1 U20801 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n17581) );
  AOI22_X1 U20802 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17643), .B1(n17577), .B2(
        n17718), .ZN(n17580) );
  OAI211_X1 U20803 ( .C1(n17582), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17722), .B(
        n17578), .ZN(n17579) );
  OAI211_X1 U20804 ( .C1(n17648), .C2(n17581), .A(n17580), .B(n17579), .ZN(
        P3_U2707) );
  AOI22_X1 U20805 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17643), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17638), .ZN(n17585) );
  AOI211_X1 U20806 ( .C1(n17789), .C2(n17588), .A(n17582), .B(n17684), .ZN(
        n17583) );
  INV_X1 U20807 ( .A(n17583), .ZN(n17584) );
  OAI211_X1 U20808 ( .C1(n17713), .C2(n17586), .A(n17585), .B(n17584), .ZN(
        P3_U2708) );
  INV_X1 U20809 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n17591) );
  AOI22_X1 U20810 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17643), .B1(n17587), .B2(
        n17718), .ZN(n17590) );
  OAI211_X1 U20811 ( .C1(n17592), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17722), .B(
        n17588), .ZN(n17589) );
  OAI211_X1 U20812 ( .C1(n17648), .C2(n17591), .A(n17590), .B(n17589), .ZN(
        P3_U2709) );
  AOI22_X1 U20813 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17643), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17638), .ZN(n17595) );
  AOI211_X1 U20814 ( .C1(n17786), .C2(n17598), .A(n17592), .B(n17684), .ZN(
        n17593) );
  INV_X1 U20815 ( .A(n17593), .ZN(n17594) );
  OAI211_X1 U20816 ( .C1(n17596), .C2(n17713), .A(n17595), .B(n17594), .ZN(
        P3_U2710) );
  AOI22_X1 U20817 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17643), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17638), .ZN(n17601) );
  OAI21_X1 U20818 ( .B1(n17784), .B2(n17684), .A(n17597), .ZN(n17599) );
  NAND2_X1 U20819 ( .A1(n17599), .A2(n17598), .ZN(n17600) );
  OAI211_X1 U20820 ( .C1(n17602), .C2(n17713), .A(n17601), .B(n17600), .ZN(
        P3_U2711) );
  AOI211_X1 U20821 ( .C1(n17782), .C2(n17604), .A(n17684), .B(n17603), .ZN(
        n17605) );
  AOI21_X1 U20822 ( .B1(n17638), .B2(BUF2_REG_23__SCAN_IN), .A(n17605), .ZN(
        n17607) );
  NAND2_X1 U20823 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17643), .ZN(n17606) );
  OAI211_X1 U20824 ( .C1(n17608), .C2(n17713), .A(n17607), .B(n17606), .ZN(
        P3_U2712) );
  INV_X1 U20825 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17770) );
  NAND2_X1 U20826 ( .A1(n18548), .A2(n17644), .ZN(n17634) );
  NAND2_X1 U20827 ( .A1(n17609), .A2(n17635), .ZN(n17617) );
  INV_X1 U20828 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n17611) );
  OAI22_X1 U20829 ( .A1(n17611), .A2(n17648), .B1(n17713), .B2(n17610), .ZN(
        n17612) );
  INV_X1 U20830 ( .A(n17612), .ZN(n17615) );
  NAND2_X1 U20831 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17635), .ZN(n17630) );
  NAND2_X1 U20832 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17626), .ZN(n17621) );
  INV_X1 U20833 ( .A(n17621), .ZN(n17618) );
  OAI22_X1 U20834 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17653), .B1(n17684), 
        .B2(n17618), .ZN(n17613) );
  AOI22_X1 U20835 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17643), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17613), .ZN(n17614) );
  OAI211_X1 U20836 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17617), .A(n17615), .B(
        n17614), .ZN(P3_U2713) );
  AOI22_X1 U20837 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17643), .B1(n17718), .B2(
        n17616), .ZN(n17620) );
  OAI211_X1 U20838 ( .C1(n17618), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17722), .B(
        n17617), .ZN(n17619) );
  OAI211_X1 U20839 ( .C1(n17648), .C2(n15681), .A(n17620), .B(n17619), .ZN(
        P3_U2714) );
  AOI22_X1 U20840 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17643), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17638), .ZN(n17623) );
  OAI211_X1 U20841 ( .C1(n17626), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17722), .B(
        n17621), .ZN(n17622) );
  OAI211_X1 U20842 ( .C1(n17624), .C2(n17713), .A(n17623), .B(n17622), .ZN(
        P3_U2715) );
  INV_X1 U20843 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n18527) );
  AOI22_X1 U20844 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17643), .B1(n17718), .B2(
        n17625), .ZN(n17629) );
  AOI211_X1 U20845 ( .C1(n17774), .C2(n17630), .A(n17626), .B(n17684), .ZN(
        n17627) );
  INV_X1 U20846 ( .A(n17627), .ZN(n17628) );
  OAI211_X1 U20847 ( .C1(n17648), .C2(n18527), .A(n17629), .B(n17628), .ZN(
        P3_U2716) );
  AOI22_X1 U20848 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17643), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17638), .ZN(n17632) );
  OAI211_X1 U20849 ( .C1(n17635), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17722), .B(
        n17630), .ZN(n17631) );
  OAI211_X1 U20850 ( .C1(n17633), .C2(n17713), .A(n17632), .B(n17631), .ZN(
        P3_U2717) );
  OAI21_X1 U20851 ( .B1(n17770), .B2(n17684), .A(n17634), .ZN(n17637) );
  INV_X1 U20852 ( .A(n17635), .ZN(n17636) );
  NAND2_X1 U20853 ( .A1(n17637), .A2(n17636), .ZN(n17640) );
  AOI22_X1 U20854 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17643), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17638), .ZN(n17639) );
  OAI211_X1 U20855 ( .C1(n17641), .C2(n17713), .A(n17640), .B(n17639), .ZN(
        P3_U2718) );
  AOI22_X1 U20856 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17643), .B1(n17718), .B2(
        n17642), .ZN(n17647) );
  AOI211_X1 U20857 ( .C1(n17768), .C2(n17649), .A(n17684), .B(n17644), .ZN(
        n17645) );
  INV_X1 U20858 ( .A(n17645), .ZN(n17646) );
  OAI211_X1 U20859 ( .C1(n17648), .C2(n14436), .A(n17647), .B(n17646), .ZN(
        P3_U2719) );
  NAND2_X1 U20860 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17719), .ZN(n17651) );
  OAI211_X1 U20861 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n17659), .A(n17722), .B(
        n17649), .ZN(n17650) );
  OAI211_X1 U20862 ( .C1(n17652), .C2(n17713), .A(n17651), .B(n17650), .ZN(
        P3_U2720) );
  INV_X1 U20863 ( .A(BUF2_REG_14__SCAN_IN), .ZN(n17662) );
  INV_X1 U20864 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17813) );
  INV_X1 U20865 ( .A(n17653), .ZN(n17654) );
  NAND2_X1 U20866 ( .A1(n17655), .A2(n17654), .ZN(n17693) );
  NOR2_X1 U20867 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17656), .ZN(n17657) );
  AOI22_X1 U20868 ( .A1(n17718), .A2(n17658), .B1(n17682), .B2(n17657), .ZN(
        n17661) );
  INV_X1 U20869 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17827) );
  OR3_X1 U20870 ( .A1(n17827), .A2(n17684), .A3(n17659), .ZN(n17660) );
  OAI211_X1 U20871 ( .C1(n17716), .C2(n17662), .A(n17661), .B(n17660), .ZN(
        P3_U2721) );
  INV_X1 U20872 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17819) );
  NAND2_X1 U20873 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17682), .ZN(n17677) );
  NOR2_X1 U20874 ( .A1(n17819), .A2(n17677), .ZN(n17674) );
  NAND2_X1 U20875 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17674), .ZN(n17666) );
  NAND2_X1 U20876 ( .A1(n17666), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n17665) );
  AOI22_X1 U20877 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17719), .B1(n17718), .B2(
        n17663), .ZN(n17664) );
  OAI221_X1 U20878 ( .B1(n17666), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n17665), 
        .C2(n17684), .A(n17664), .ZN(P3_U2722) );
  INV_X1 U20879 ( .A(n17666), .ZN(n17669) );
  AOI21_X1 U20880 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17722), .A(n17674), .ZN(
        n17668) );
  OAI222_X1 U20881 ( .A1(n17716), .A2(n17670), .B1(n17669), .B2(n17668), .C1(
        n17713), .C2(n17667), .ZN(P3_U2723) );
  INV_X1 U20882 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17675) );
  OAI21_X1 U20883 ( .B1(n17819), .B2(n17684), .A(n17677), .ZN(n17671) );
  INV_X1 U20884 ( .A(n17671), .ZN(n17673) );
  OAI222_X1 U20885 ( .A1(n17716), .A2(n17675), .B1(n17674), .B2(n17673), .C1(
        n17713), .C2(n17672), .ZN(P3_U2724) );
  AOI22_X1 U20886 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17719), .B1(n17718), .B2(
        n17676), .ZN(n17679) );
  OAI211_X1 U20887 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17682), .A(n17722), .B(
        n17677), .ZN(n17678) );
  NAND2_X1 U20888 ( .A1(n17679), .A2(n17678), .ZN(P3_U2725) );
  INV_X1 U20889 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17683) );
  AOI21_X1 U20890 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17722), .A(n17688), .ZN(
        n17681) );
  OAI222_X1 U20891 ( .A1(n17716), .A2(n17683), .B1(n17682), .B2(n17681), .C1(
        n17713), .C2(n17680), .ZN(P3_U2726) );
  INV_X1 U20892 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17689) );
  OAI21_X1 U20893 ( .B1(n17813), .B2(n17684), .A(n17693), .ZN(n17685) );
  INV_X1 U20894 ( .A(n17685), .ZN(n17687) );
  OAI222_X1 U20895 ( .A1(n17716), .A2(n17689), .B1(n17688), .B2(n17687), .C1(
        n17713), .C2(n17686), .ZN(P3_U2727) );
  INV_X1 U20896 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17807) );
  INV_X1 U20897 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17803) );
  NAND3_X1 U20898 ( .A1(n17690), .A2(P3_EAX_REG_1__SCAN_IN), .A3(
        P3_EAX_REG_0__SCAN_IN), .ZN(n17721) );
  NOR2_X1 U20899 ( .A1(n17691), .A2(n17721), .ZN(n17711) );
  NAND2_X1 U20900 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17711), .ZN(n17707) );
  NAND2_X1 U20901 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17710), .ZN(n17700) );
  NOR2_X1 U20902 ( .A1(n17807), .A2(n17700), .ZN(n17703) );
  NAND2_X1 U20903 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17703), .ZN(n17696) );
  AOI22_X1 U20904 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17719), .B1(n17718), .B2(
        n17692), .ZN(n17695) );
  NAND3_X1 U20905 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17722), .A3(n17693), .ZN(
        n17694) );
  OAI211_X1 U20906 ( .C1(P3_EAX_REG_7__SCAN_IN), .C2(n17696), .A(n17695), .B(
        n17694), .ZN(P3_U2728) );
  INV_X1 U20907 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18541) );
  INV_X1 U20908 ( .A(n17696), .ZN(n17699) );
  AOI21_X1 U20909 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17722), .A(n17703), .ZN(
        n17698) );
  OAI222_X1 U20910 ( .A1(n18541), .A2(n17716), .B1(n17699), .B2(n17698), .C1(
        n17713), .C2(n17697), .ZN(P3_U2729) );
  INV_X1 U20911 ( .A(n17700), .ZN(n17706) );
  AOI21_X1 U20912 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17722), .A(n17706), .ZN(
        n17702) );
  OAI222_X1 U20913 ( .A1(n18537), .A2(n17716), .B1(n17703), .B2(n17702), .C1(
        n17713), .C2(n17701), .ZN(P3_U2730) );
  INV_X1 U20914 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18532) );
  AOI21_X1 U20915 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17722), .A(n17710), .ZN(
        n17705) );
  OAI222_X1 U20916 ( .A1(n18532), .A2(n17716), .B1(n17706), .B2(n17705), .C1(
        n17713), .C2(n17704), .ZN(P3_U2731) );
  INV_X1 U20917 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18528) );
  INV_X1 U20918 ( .A(n17707), .ZN(n17715) );
  AOI21_X1 U20919 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17722), .A(n17715), .ZN(
        n17709) );
  OAI222_X1 U20920 ( .A1(n18528), .A2(n17716), .B1(n17710), .B2(n17709), .C1(
        n17713), .C2(n17708), .ZN(P3_U2732) );
  INV_X1 U20921 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18523) );
  AOI21_X1 U20922 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17722), .A(n17711), .ZN(
        n17714) );
  OAI222_X1 U20923 ( .A1(n18523), .A2(n17716), .B1(n17715), .B2(n17714), .C1(
        n17713), .C2(n17712), .ZN(P3_U2733) );
  AOI22_X1 U20924 ( .A1(n17719), .A2(BUF2_REG_1__SCAN_IN), .B1(n17718), .B2(
        n17717), .ZN(n17725) );
  NOR2_X1 U20925 ( .A1(n17720), .A2(n17797), .ZN(n17723) );
  OAI211_X1 U20926 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(n17723), .A(n17722), .B(
        n17721), .ZN(n17724) );
  NAND2_X1 U20927 ( .A1(n17725), .A2(n17724), .ZN(P3_U2734) );
  NAND2_X1 U20928 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n18019), .ZN(n19181) );
  INV_X2 U20929 ( .A(n19181), .ZN(n17761) );
  NOR2_X4 U20930 ( .A1(n17761), .A2(n17745), .ZN(n17741) );
  AND2_X1 U20931 ( .A1(n17741), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20932 ( .A1(n17745), .A2(n17727), .ZN(n17744) );
  AOI22_X1 U20933 ( .A1(n17761), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17741), .ZN(n17728) );
  OAI21_X1 U20934 ( .B1(n17795), .B2(n17744), .A(n17728), .ZN(P3_U2737) );
  INV_X1 U20935 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17793) );
  AOI22_X1 U20936 ( .A1(n17761), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17729) );
  OAI21_X1 U20937 ( .B1(n17793), .B2(n17744), .A(n17729), .ZN(P3_U2738) );
  INV_X1 U20938 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17791) );
  AOI22_X1 U20939 ( .A1(n17761), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17730) );
  OAI21_X1 U20940 ( .B1(n17791), .B2(n17744), .A(n17730), .ZN(P3_U2739) );
  AOI22_X1 U20941 ( .A1(n17761), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17731) );
  OAI21_X1 U20942 ( .B1(n17789), .B2(n17744), .A(n17731), .ZN(P3_U2740) );
  AOI22_X1 U20943 ( .A1(n17761), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17732) );
  OAI21_X1 U20944 ( .B1(n9711), .B2(n17744), .A(n17732), .ZN(P3_U2741) );
  AOI22_X1 U20945 ( .A1(n17761), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17733) );
  OAI21_X1 U20946 ( .B1(n17786), .B2(n17744), .A(n17733), .ZN(P3_U2742) );
  AOI22_X1 U20947 ( .A1(n17761), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17734) );
  OAI21_X1 U20948 ( .B1(n17784), .B2(n17744), .A(n17734), .ZN(P3_U2743) );
  AOI22_X1 U20949 ( .A1(n17761), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17735) );
  OAI21_X1 U20950 ( .B1(n17782), .B2(n17744), .A(n17735), .ZN(P3_U2744) );
  INV_X1 U20951 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17780) );
  AOI22_X1 U20952 ( .A1(n17761), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17736) );
  OAI21_X1 U20953 ( .B1(n17780), .B2(n17744), .A(n17736), .ZN(P3_U2745) );
  AOI22_X1 U20954 ( .A1(n17761), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17737) );
  OAI21_X1 U20955 ( .B1(n17778), .B2(n17744), .A(n17737), .ZN(P3_U2746) );
  AOI22_X1 U20956 ( .A1(n17761), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17738) );
  OAI21_X1 U20957 ( .B1(n17776), .B2(n17744), .A(n17738), .ZN(P3_U2747) );
  AOI22_X1 U20958 ( .A1(n17761), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17739) );
  OAI21_X1 U20959 ( .B1(n17774), .B2(n17744), .A(n17739), .ZN(P3_U2748) );
  AOI22_X1 U20960 ( .A1(n17761), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17740) );
  OAI21_X1 U20961 ( .B1(n17772), .B2(n17744), .A(n17740), .ZN(P3_U2749) );
  AOI22_X1 U20962 ( .A1(n17761), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17742) );
  OAI21_X1 U20963 ( .B1(n17770), .B2(n17744), .A(n17742), .ZN(P3_U2750) );
  AOI22_X1 U20964 ( .A1(n17761), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17743) );
  OAI21_X1 U20965 ( .B1(n17768), .B2(n17744), .A(n17743), .ZN(P3_U2751) );
  INV_X1 U20966 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17832) );
  AOI22_X1 U20967 ( .A1(n17761), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17746) );
  OAI21_X1 U20968 ( .B1(n17832), .B2(n17763), .A(n17746), .ZN(P3_U2752) );
  AOI22_X1 U20969 ( .A1(n17761), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17747) );
  OAI21_X1 U20970 ( .B1(n17827), .B2(n17763), .A(n17747), .ZN(P3_U2753) );
  INV_X1 U20971 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17825) );
  AOI22_X1 U20972 ( .A1(n17761), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17748) );
  OAI21_X1 U20973 ( .B1(n17825), .B2(n17763), .A(n17748), .ZN(P3_U2754) );
  INV_X1 U20974 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17823) );
  AOI22_X1 U20975 ( .A1(n17761), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17749) );
  OAI21_X1 U20976 ( .B1(n17823), .B2(n17763), .A(n17749), .ZN(P3_U2755) );
  AOI22_X1 U20977 ( .A1(n17761), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17750) );
  OAI21_X1 U20978 ( .B1(n17819), .B2(n17763), .A(n17750), .ZN(P3_U2756) );
  INV_X1 U20979 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17817) );
  AOI22_X1 U20980 ( .A1(n17761), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17751) );
  OAI21_X1 U20981 ( .B1(n17817), .B2(n17763), .A(n17751), .ZN(P3_U2757) );
  INV_X1 U20982 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17815) );
  AOI22_X1 U20983 ( .A1(n17761), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17752) );
  OAI21_X1 U20984 ( .B1(n17815), .B2(n17763), .A(n17752), .ZN(P3_U2758) );
  AOI22_X1 U20985 ( .A1(n17761), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17753) );
  OAI21_X1 U20986 ( .B1(n17813), .B2(n17763), .A(n17753), .ZN(P3_U2759) );
  INV_X1 U20987 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17811) );
  AOI22_X1 U20988 ( .A1(n17761), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17754) );
  OAI21_X1 U20989 ( .B1(n17811), .B2(n17763), .A(n17754), .ZN(P3_U2760) );
  INV_X1 U20990 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17809) );
  AOI22_X1 U20991 ( .A1(n17761), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17755) );
  OAI21_X1 U20992 ( .B1(n17809), .B2(n17763), .A(n17755), .ZN(P3_U2761) );
  AOI22_X1 U20993 ( .A1(n17761), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17756) );
  OAI21_X1 U20994 ( .B1(n17807), .B2(n17763), .A(n17756), .ZN(P3_U2762) );
  INV_X1 U20995 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17805) );
  AOI22_X1 U20996 ( .A1(n17761), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17757) );
  OAI21_X1 U20997 ( .B1(n17805), .B2(n17763), .A(n17757), .ZN(P3_U2763) );
  AOI22_X1 U20998 ( .A1(n17761), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17758) );
  OAI21_X1 U20999 ( .B1(n17803), .B2(n17763), .A(n17758), .ZN(P3_U2764) );
  INV_X1 U21000 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17801) );
  AOI22_X1 U21001 ( .A1(n17761), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17759) );
  OAI21_X1 U21002 ( .B1(n17801), .B2(n17763), .A(n17759), .ZN(P3_U2765) );
  INV_X1 U21003 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17799) );
  AOI22_X1 U21004 ( .A1(n17761), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17760) );
  OAI21_X1 U21005 ( .B1(n17799), .B2(n17763), .A(n17760), .ZN(P3_U2766) );
  AOI22_X1 U21006 ( .A1(n17761), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17741), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17762) );
  OAI21_X1 U21007 ( .B1(n17797), .B2(n17763), .A(n17762), .ZN(P3_U2767) );
  NOR2_X1 U21008 ( .A1(n17765), .A2(n17764), .ZN(n17766) );
  AOI22_X1 U21009 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17829), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17820), .ZN(n17767) );
  OAI21_X1 U21010 ( .B1(n17768), .B2(n17831), .A(n17767), .ZN(P3_U2768) );
  AOI22_X1 U21011 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17829), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17820), .ZN(n17769) );
  OAI21_X1 U21012 ( .B1(n17770), .B2(n17831), .A(n17769), .ZN(P3_U2769) );
  AOI22_X1 U21013 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17829), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17820), .ZN(n17771) );
  OAI21_X1 U21014 ( .B1(n17772), .B2(n17831), .A(n17771), .ZN(P3_U2770) );
  AOI22_X1 U21015 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17821), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17820), .ZN(n17773) );
  OAI21_X1 U21016 ( .B1(n17774), .B2(n17831), .A(n17773), .ZN(P3_U2771) );
  AOI22_X1 U21017 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17821), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17820), .ZN(n17775) );
  OAI21_X1 U21018 ( .B1(n17776), .B2(n17831), .A(n17775), .ZN(P3_U2772) );
  AOI22_X1 U21019 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17821), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17820), .ZN(n17777) );
  OAI21_X1 U21020 ( .B1(n17778), .B2(n17831), .A(n17777), .ZN(P3_U2773) );
  AOI22_X1 U21021 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17821), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17820), .ZN(n17779) );
  OAI21_X1 U21022 ( .B1(n17780), .B2(n17831), .A(n17779), .ZN(P3_U2774) );
  AOI22_X1 U21023 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17821), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17820), .ZN(n17781) );
  OAI21_X1 U21024 ( .B1(n17782), .B2(n17831), .A(n17781), .ZN(P3_U2775) );
  AOI22_X1 U21025 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17821), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17820), .ZN(n17783) );
  OAI21_X1 U21026 ( .B1(n17784), .B2(n17831), .A(n17783), .ZN(P3_U2776) );
  AOI22_X1 U21027 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17821), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17820), .ZN(n17785) );
  OAI21_X1 U21028 ( .B1(n17786), .B2(n17831), .A(n17785), .ZN(P3_U2777) );
  AOI22_X1 U21029 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17821), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17820), .ZN(n17787) );
  OAI21_X1 U21030 ( .B1(n9711), .B2(n17831), .A(n17787), .ZN(P3_U2778) );
  AOI22_X1 U21031 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17821), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17820), .ZN(n17788) );
  OAI21_X1 U21032 ( .B1(n17789), .B2(n17831), .A(n17788), .ZN(P3_U2779) );
  AOI22_X1 U21033 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17829), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17820), .ZN(n17790) );
  OAI21_X1 U21034 ( .B1(n17791), .B2(n17831), .A(n17790), .ZN(P3_U2780) );
  AOI22_X1 U21035 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17829), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17820), .ZN(n17792) );
  OAI21_X1 U21036 ( .B1(n17793), .B2(n17831), .A(n17792), .ZN(P3_U2781) );
  AOI22_X1 U21037 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17829), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17820), .ZN(n17794) );
  OAI21_X1 U21038 ( .B1(n17795), .B2(n17831), .A(n17794), .ZN(P3_U2782) );
  AOI22_X1 U21039 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17829), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17820), .ZN(n17796) );
  OAI21_X1 U21040 ( .B1(n17797), .B2(n17831), .A(n17796), .ZN(P3_U2783) );
  AOI22_X1 U21041 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17829), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17820), .ZN(n17798) );
  OAI21_X1 U21042 ( .B1(n17799), .B2(n17831), .A(n17798), .ZN(P3_U2784) );
  AOI22_X1 U21043 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17829), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17820), .ZN(n17800) );
  OAI21_X1 U21044 ( .B1(n17801), .B2(n17831), .A(n17800), .ZN(P3_U2785) );
  AOI22_X1 U21045 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17829), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17820), .ZN(n17802) );
  OAI21_X1 U21046 ( .B1(n17803), .B2(n17831), .A(n17802), .ZN(P3_U2786) );
  AOI22_X1 U21047 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17829), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17828), .ZN(n17804) );
  OAI21_X1 U21048 ( .B1(n17805), .B2(n17831), .A(n17804), .ZN(P3_U2787) );
  AOI22_X1 U21049 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17829), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17828), .ZN(n17806) );
  OAI21_X1 U21050 ( .B1(n17807), .B2(n17831), .A(n17806), .ZN(P3_U2788) );
  AOI22_X1 U21051 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17829), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17828), .ZN(n17808) );
  OAI21_X1 U21052 ( .B1(n17809), .B2(n17831), .A(n17808), .ZN(P3_U2789) );
  AOI22_X1 U21053 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17829), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17828), .ZN(n17810) );
  OAI21_X1 U21054 ( .B1(n17811), .B2(n17831), .A(n17810), .ZN(P3_U2790) );
  AOI22_X1 U21055 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17829), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17828), .ZN(n17812) );
  OAI21_X1 U21056 ( .B1(n17813), .B2(n17831), .A(n17812), .ZN(P3_U2791) );
  AOI22_X1 U21057 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17829), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17828), .ZN(n17814) );
  OAI21_X1 U21058 ( .B1(n17815), .B2(n17831), .A(n17814), .ZN(P3_U2792) );
  AOI22_X1 U21059 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17821), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17820), .ZN(n17816) );
  OAI21_X1 U21060 ( .B1(n17817), .B2(n17831), .A(n17816), .ZN(P3_U2793) );
  AOI22_X1 U21061 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17829), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17828), .ZN(n17818) );
  OAI21_X1 U21062 ( .B1(n17819), .B2(n17831), .A(n17818), .ZN(P3_U2794) );
  AOI22_X1 U21063 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17821), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17820), .ZN(n17822) );
  OAI21_X1 U21064 ( .B1(n17823), .B2(n17831), .A(n17822), .ZN(P3_U2795) );
  AOI22_X1 U21065 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17829), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17828), .ZN(n17824) );
  OAI21_X1 U21066 ( .B1(n17825), .B2(n17831), .A(n17824), .ZN(P3_U2796) );
  AOI22_X1 U21067 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17829), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17828), .ZN(n17826) );
  OAI21_X1 U21068 ( .B1(n17827), .B2(n17831), .A(n17826), .ZN(P3_U2797) );
  AOI22_X1 U21069 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17829), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17828), .ZN(n17830) );
  OAI21_X1 U21070 ( .B1(n17832), .B2(n17831), .A(n17830), .ZN(P3_U2798) );
  AOI22_X1 U21071 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17834), .B1(
        n18036), .B2(n17833), .ZN(n17844) );
  NOR2_X1 U21072 ( .A1(n17836), .A2(n17835), .ZN(n17837) );
  XOR2_X1 U21073 ( .A(n18080), .B(n17837), .Z(n18193) );
  AOI22_X1 U21074 ( .A1(n18075), .A2(n18193), .B1(n17839), .B2(n17838), .ZN(
        n17843) );
  OAI21_X1 U21075 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17841), .A(
        n17840), .ZN(n17842) );
  NAND2_X1 U21076 ( .A1(n18499), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n18194) );
  NAND4_X1 U21077 ( .A1(n17844), .A2(n17843), .A3(n17842), .A4(n18194), .ZN(
        P3_U2803) );
  AOI21_X1 U21078 ( .B1(n17845), .B2(n18545), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17853) );
  AOI22_X1 U21079 ( .A1(n18499), .A2(P3_REIP_REG_26__SCAN_IN), .B1(n17846), 
        .B2(n18170), .ZN(n17852) );
  OAI21_X1 U21080 ( .B1(n17848), .B2(n18186), .A(n17847), .ZN(n18198) );
  NAND2_X1 U21081 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17855) );
  NOR2_X1 U21082 ( .A1(n17855), .A2(n17878), .ZN(n18184) );
  NAND2_X1 U21083 ( .A1(n18184), .A2(n18186), .ZN(n18202) );
  OAI22_X1 U21084 ( .A1(n17849), .A2(n18186), .B1(n17989), .B2(n18202), .ZN(
        n17850) );
  AOI21_X1 U21085 ( .B1(n18075), .B2(n18198), .A(n17850), .ZN(n17851) );
  OAI211_X1 U21086 ( .C1(n17854), .C2(n17853), .A(n17852), .B(n17851), .ZN(
        P3_U2804) );
  NOR2_X1 U21087 ( .A1(n18313), .A2(n17878), .ZN(n18222) );
  INV_X1 U21088 ( .A(n18222), .ZN(n17869) );
  NOR2_X1 U21089 ( .A1(n17881), .A2(n17869), .ZN(n17856) );
  OAI22_X1 U21090 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17856), .B1(
        n17855), .B2(n17869), .ZN(n18215) );
  AND2_X1 U21091 ( .A1(n11668), .A2(n18545), .ZN(n17886) );
  AOI211_X1 U21092 ( .C1(n18019), .C2(n17891), .A(n17886), .B(n18118), .ZN(
        n17894) );
  OAI21_X1 U21093 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17929), .A(
        n17894), .ZN(n17873) );
  NOR2_X1 U21094 ( .A1(n17941), .A2(n11668), .ZN(n17875) );
  OAI211_X1 U21095 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17875), .B(n17857), .ZN(n17859) );
  NOR2_X1 U21096 ( .A1(n18482), .A2(n19114), .ZN(n18210) );
  INV_X1 U21097 ( .A(n18210), .ZN(n17858) );
  OAI211_X1 U21098 ( .C1(n18024), .C2(n17860), .A(n17859), .B(n17858), .ZN(
        n17861) );
  AOI21_X1 U21099 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n17873), .A(
        n17861), .ZN(n17867) );
  NOR3_X1 U21100 ( .A1(n17878), .A2(n18312), .A3(n17881), .ZN(n17862) );
  XOR2_X1 U21101 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17862), .Z(
        n18212) );
  AOI21_X1 U21102 ( .B1(n18066), .B2(n17864), .A(n17863), .ZN(n17865) );
  XOR2_X1 U21103 ( .A(n17865), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n18211) );
  AOI22_X1 U21104 ( .A1(n18150), .A2(n18212), .B1(n18075), .B2(n18211), .ZN(
        n17866) );
  OAI211_X1 U21105 ( .C1(n18027), .C2(n18215), .A(n17867), .B(n17866), .ZN(
        P3_U2805) );
  NAND2_X1 U21106 ( .A1(n18241), .A2(n17868), .ZN(n18220) );
  AOI22_X1 U21107 ( .A1(n18090), .A2(n17869), .B1(n18150), .B2(n18220), .ZN(
        n17898) );
  AOI22_X1 U21108 ( .A1(n18349), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n18036), 
        .B2(n17870), .ZN(n17871) );
  INV_X1 U21109 ( .A(n17871), .ZN(n17872) );
  AOI221_X1 U21110 ( .B1(n17875), .B2(n17874), .C1(n17873), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17872), .ZN(n17880) );
  OAI21_X1 U21111 ( .B1(n17877), .B2(n17881), .A(n17876), .ZN(n18217) );
  NOR2_X1 U21112 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17878), .ZN(
        n18216) );
  AOI22_X1 U21113 ( .A1(n18075), .A2(n18217), .B1(n17914), .B2(n18216), .ZN(
        n17879) );
  OAI211_X1 U21114 ( .C1(n17898), .C2(n17881), .A(n17880), .B(n17879), .ZN(
        P3_U2806) );
  NAND2_X1 U21115 ( .A1(n18218), .A2(n17914), .ZN(n17899) );
  OAI22_X1 U21116 ( .A1(n17900), .A2(n17882), .B1(n18066), .B2(n18239), .ZN(
        n17883) );
  NOR2_X1 U21117 ( .A1(n17883), .A2(n17935), .ZN(n17884) );
  XOR2_X1 U21118 ( .A(n17884), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n18229) );
  INV_X1 U21119 ( .A(n17885), .ZN(n17889) );
  AOI22_X1 U21120 ( .A1(n18349), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n17887), 
        .B2(n17886), .ZN(n17888) );
  OAI21_X1 U21121 ( .B1(n18024), .B2(n17889), .A(n17888), .ZN(n17896) );
  NAND2_X1 U21122 ( .A1(n17890), .A2(n17893), .ZN(n17892) );
  OAI22_X1 U21123 ( .A1(n17894), .A2(n17893), .B1(n17892), .B2(n17891), .ZN(
        n17895) );
  AOI211_X1 U21124 ( .C1(n18075), .C2(n18229), .A(n17896), .B(n17895), .ZN(
        n17897) );
  OAI221_X1 U21125 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17899), 
        .C1(n18223), .C2(n17898), .A(n17897), .ZN(P3_U2807) );
  INV_X1 U21126 ( .A(n17900), .ZN(n17901) );
  INV_X1 U21127 ( .A(n18247), .ZN(n18238) );
  XOR2_X1 U21128 ( .A(n18239), .B(n17902), .Z(n18254) );
  AOI22_X1 U21129 ( .A1(n18090), .A2(n18313), .B1(n18150), .B2(n18312), .ZN(
        n17988) );
  OAI21_X1 U21130 ( .B1(n18247), .B2(n17934), .A(n17988), .ZN(n17925) );
  AOI21_X1 U21131 ( .B1(n17907), .B2(n17976), .A(n18118), .ZN(n17903) );
  INV_X1 U21132 ( .A(n17903), .ZN(n17904) );
  AOI21_X1 U21133 ( .B1(n18019), .B2(n17905), .A(n17904), .ZN(n17931) );
  OAI21_X1 U21134 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17929), .A(
        n17931), .ZN(n17917) );
  AOI22_X1 U21135 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17917), .B1(
        n18036), .B2(n17906), .ZN(n17910) );
  NOR2_X1 U21136 ( .A1(n17941), .A2(n17907), .ZN(n17919) );
  OAI211_X1 U21137 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17919), .B(n17908), .ZN(n17909) );
  OAI211_X1 U21138 ( .C1(n19108), .C2(n18482), .A(n17910), .B(n17909), .ZN(
        n17911) );
  AOI21_X1 U21139 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17925), .A(
        n17911), .ZN(n17913) );
  NAND3_X1 U21140 ( .A1(n18247), .A2(n17914), .A3(n18239), .ZN(n17912) );
  OAI211_X1 U21141 ( .C1(n18093), .C2(n18254), .A(n17913), .B(n17912), .ZN(
        P3_U2808) );
  OR2_X1 U21142 ( .A1(n17923), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n18263) );
  NAND2_X1 U21143 ( .A1(n18286), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n18243) );
  INV_X1 U21144 ( .A(n18243), .ZN(n18257) );
  NAND2_X1 U21145 ( .A1(n17914), .A2(n18257), .ZN(n17951) );
  OAI22_X1 U21146 ( .A1(n18482), .A2(n19107), .B1(n18024), .B2(n17915), .ZN(
        n17916) );
  AOI221_X1 U21147 ( .B1(n17919), .B2(n17918), .C1(n17917), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17916), .ZN(n17927) );
  NAND3_X1 U21148 ( .A1(n18066), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17920), .ZN(n17946) );
  INV_X1 U21149 ( .A(n17921), .ZN(n17959) );
  OAI22_X1 U21150 ( .A1(n17923), .A2(n17946), .B1(n17922), .B2(n17959), .ZN(
        n17924) );
  XOR2_X1 U21151 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n17924), .Z(
        n18256) );
  AOI22_X1 U21152 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17925), .B1(
        n18075), .B2(n18256), .ZN(n17926) );
  OAI211_X1 U21153 ( .C1(n18263), .C2(n17951), .A(n17927), .B(n17926), .ZN(
        P3_U2809) );
  NAND2_X1 U21154 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17928), .ZN(
        n18272) );
  AOI21_X1 U21155 ( .B1(n13359), .B2(n18545), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17930) );
  OAI22_X1 U21156 ( .A1(n17931), .A2(n17930), .B1(n18482), .B2(n19104), .ZN(
        n17932) );
  AOI221_X1 U21157 ( .B1(n18036), .B2(n17933), .C1(n17890), .C2(n17933), .A(
        n17932), .ZN(n17939) );
  INV_X1 U21158 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17936) );
  NOR2_X1 U21159 ( .A1(n17936), .A2(n18243), .ZN(n18268) );
  OAI21_X1 U21160 ( .B1(n17934), .B2(n18268), .A(n17988), .ZN(n17948) );
  XOR2_X1 U21161 ( .A(n17937), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(
        n18264) );
  AOI22_X1 U21162 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17948), .B1(
        n18075), .B2(n18264), .ZN(n17938) );
  OAI211_X1 U21163 ( .C1(n17951), .C2(n18272), .A(n17939), .B(n17938), .ZN(
        P3_U2810) );
  INV_X1 U21164 ( .A(n18138), .ZN(n18171) );
  OAI21_X1 U21165 ( .B1(n18118), .B2(n13361), .A(n18171), .ZN(n17971) );
  OAI21_X1 U21166 ( .B1(n17940), .B2(n17977), .A(n17971), .ZN(n17954) );
  NOR2_X1 U21167 ( .A1(n17941), .A2(n13361), .ZN(n17956) );
  OAI211_X1 U21168 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17956), .B(n17942), .ZN(n17943) );
  NAND2_X1 U21169 ( .A1(n18349), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n18275) );
  OAI211_X1 U21170 ( .C1(n18024), .C2(n17944), .A(n17943), .B(n18275), .ZN(
        n17945) );
  AOI21_X1 U21171 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17954), .A(
        n17945), .ZN(n17950) );
  OAI21_X1 U21172 ( .B1(n17957), .B2(n17959), .A(n17946), .ZN(n17947) );
  XOR2_X1 U21173 ( .A(n17947), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n18273) );
  AOI22_X1 U21174 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17948), .B1(
        n18075), .B2(n18273), .ZN(n17949) );
  OAI211_X1 U21175 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17951), .A(
        n17950), .B(n17949), .ZN(P3_U2811) );
  NAND2_X1 U21176 ( .A1(n18286), .A2(n17958), .ZN(n18290) );
  OAI22_X1 U21177 ( .A1(n18482), .A2(n19100), .B1(n18024), .B2(n17952), .ZN(
        n17953) );
  AOI221_X1 U21178 ( .B1(n17956), .B2(n17955), .C1(n17954), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17953), .ZN(n17962) );
  OAI21_X1 U21179 ( .B1(n18286), .B2(n17989), .A(n17988), .ZN(n17969) );
  OAI21_X1 U21180 ( .B1(n18080), .B2(n17958), .A(n17957), .ZN(n17960) );
  XOR2_X1 U21181 ( .A(n17960), .B(n17959), .Z(n18281) );
  AOI22_X1 U21182 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17969), .B1(
        n18075), .B2(n18281), .ZN(n17961) );
  OAI211_X1 U21183 ( .C1(n17989), .C2(n18290), .A(n17962), .B(n17961), .ZN(
        P3_U2812) );
  AOI21_X1 U21184 ( .B1(n17963), .B2(n18545), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17972) );
  INV_X1 U21185 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n18295) );
  OAI21_X1 U21186 ( .B1(n18310), .B2(n17989), .A(n18295), .ZN(n17968) );
  AOI21_X1 U21187 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17965), .A(
        n17964), .ZN(n18298) );
  OAI22_X1 U21188 ( .A1(n18160), .A2(n17966), .B1(n18298), .B2(n18093), .ZN(
        n17967) );
  AOI21_X1 U21189 ( .B1(n17969), .B2(n17968), .A(n17967), .ZN(n17970) );
  NAND2_X1 U21190 ( .A1(n18499), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n18296) );
  OAI211_X1 U21191 ( .C1(n17972), .C2(n17971), .A(n17970), .B(n18296), .ZN(
        P3_U2813) );
  NAND2_X1 U21192 ( .A1(n18066), .A2(n18029), .ZN(n18056) );
  AOI22_X1 U21193 ( .A1(n18068), .A2(n18280), .B1(n9675), .B2(n18080), .ZN(
        n17974) );
  XOR2_X1 U21194 ( .A(n18310), .B(n17974), .Z(n18307) );
  AOI21_X1 U21195 ( .B1(n17976), .B2(n17975), .A(n18118), .ZN(n18007) );
  OAI21_X1 U21196 ( .B1(n17978), .B2(n17977), .A(n18007), .ZN(n17997) );
  AOI22_X1 U21197 ( .A1(n18349), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17997), .ZN(n17984) );
  NAND2_X1 U21198 ( .A1(n17979), .A2(n17980), .ZN(n18039) );
  NOR2_X1 U21199 ( .A1(n17981), .A2(n18039), .ZN(n17996) );
  OAI211_X1 U21200 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17996), .B(n17982), .ZN(n17983) );
  OAI211_X1 U21201 ( .C1(n18024), .C2(n17985), .A(n17984), .B(n17983), .ZN(
        n17986) );
  AOI21_X1 U21202 ( .B1(n18075), .B2(n18307), .A(n17986), .ZN(n17987) );
  OAI221_X1 U21203 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17989), 
        .C1(n18310), .C2(n17988), .A(n17987), .ZN(P3_U2814) );
  AOI21_X1 U21204 ( .B1(n18314), .B2(n18004), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18319) );
  NAND2_X1 U21205 ( .A1(n18090), .A2(n18313), .ZN(n18003) );
  INV_X1 U21206 ( .A(n18335), .ZN(n18329) );
  NOR3_X1 U21207 ( .A1(n18372), .A2(n18329), .A3(n18328), .ZN(n18012) );
  NOR2_X1 U21208 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18012), .ZN(
        n18321) );
  NAND2_X1 U21209 ( .A1(n18150), .A2(n18312), .ZN(n17994) );
  NOR3_X1 U21210 ( .A1(n17990), .A2(n18328), .A3(n18363), .ZN(n17991) );
  AOI21_X1 U21211 ( .B1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n17991), .A(
        n18014), .ZN(n17992) );
  AOI221_X1 U21212 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18362), 
        .C1(n18080), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17992), .ZN(
        n17993) );
  XNOR2_X1 U21213 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17993), .ZN(
        n18326) );
  OAI22_X1 U21214 ( .A1(n18321), .A2(n17994), .B1(n18093), .B2(n18326), .ZN(
        n18001) );
  AOI22_X1 U21215 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17997), .B1(
        n17996), .B2(n17995), .ZN(n17998) );
  NAND2_X1 U21216 ( .A1(n18499), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n18324) );
  OAI211_X1 U21217 ( .C1(n18024), .C2(n17999), .A(n17998), .B(n18324), .ZN(
        n18000) );
  NOR2_X1 U21218 ( .A1(n18001), .A2(n18000), .ZN(n18002) );
  OAI21_X1 U21219 ( .B1(n18319), .B2(n18003), .A(n18002), .ZN(P3_U2815) );
  NOR2_X1 U21220 ( .A1(n18370), .A2(n18352), .ZN(n18355) );
  NAND2_X1 U21221 ( .A1(n18004), .A2(n18314), .ZN(n18005) );
  OAI221_X1 U21222 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18355), .A(n18005), .ZN(
        n18344) );
  NOR2_X1 U21223 ( .A1(n18006), .A2(n18741), .ZN(n18044) );
  NAND2_X1 U21224 ( .A1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18044), .ZN(
        n18049) );
  AOI221_X1 U21225 ( .B1(n18021), .B2(n18008), .C1(n18049), .C2(n18008), .A(
        n18007), .ZN(n18009) );
  NOR2_X1 U21226 ( .A1(n18482), .A2(n19093), .ZN(n18337) );
  AOI211_X1 U21227 ( .C1(n18010), .C2(n18170), .A(n18009), .B(n18337), .ZN(
        n18017) );
  NAND2_X1 U21228 ( .A1(n18335), .A2(n18011), .ZN(n18013) );
  AOI21_X1 U21229 ( .B1(n18328), .B2(n18013), .A(n18012), .ZN(n18341) );
  AOI22_X1 U21230 ( .A1(n18068), .A2(n18335), .B1(n18014), .B2(n18362), .ZN(
        n18015) );
  XOR2_X1 U21231 ( .A(n18328), .B(n18015), .Z(n18340) );
  AOI22_X1 U21232 ( .A1(n18150), .A2(n18341), .B1(n18075), .B2(n18340), .ZN(
        n18016) );
  OAI211_X1 U21233 ( .C1(n18027), .C2(n18344), .A(n18017), .B(n18016), .ZN(
        P3_U2816) );
  INV_X1 U21234 ( .A(n18352), .ZN(n18331) );
  NAND2_X1 U21235 ( .A1(n18331), .A2(n18333), .ZN(n18361) );
  AOI21_X1 U21236 ( .B1(n18019), .B2(n18018), .A(n18118), .ZN(n18020) );
  OAI21_X1 U21237 ( .B1(n17979), .B2(n18081), .A(n18020), .ZN(n18037) );
  NOR2_X1 U21238 ( .A1(n18482), .A2(n19090), .ZN(n18026) );
  OAI21_X1 U21239 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n18021), .ZN(n18022) );
  OAI22_X1 U21240 ( .A1(n18024), .A2(n18023), .B1(n18039), .B2(n18022), .ZN(
        n18025) );
  AOI211_X1 U21241 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18037), .A(
        n18026), .B(n18025), .ZN(n18033) );
  NOR2_X1 U21242 ( .A1(n18352), .A2(n18372), .ZN(n18350) );
  OAI22_X1 U21243 ( .A1(n18355), .A2(n18027), .B1(n18350), .B2(n18180), .ZN(
        n18041) );
  AOI22_X1 U21244 ( .A1(n18331), .A2(n18029), .B1(n18080), .B2(n18362), .ZN(
        n18030) );
  AOI21_X1 U21245 ( .B1(n18028), .B2(n18080), .A(n18030), .ZN(n18031) );
  XOR2_X1 U21246 ( .A(n18031), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n18348) );
  AOI22_X1 U21247 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18041), .B1(
        n18075), .B2(n18348), .ZN(n18032) );
  OAI211_X1 U21248 ( .C1(n9664), .C2(n18361), .A(n18033), .B(n18032), .ZN(
        P3_U2817) );
  OAI21_X1 U21249 ( .B1(n18363), .B2(n18056), .A(n18028), .ZN(n18034) );
  XOR2_X1 U21250 ( .A(n18034), .B(n18362), .Z(n18369) );
  NOR2_X1 U21251 ( .A1(n9664), .A2(n18363), .ZN(n18042) );
  AOI22_X1 U21252 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18037), .B1(
        n18036), .B2(n18035), .ZN(n18038) );
  NAND2_X1 U21253 ( .A1(n18349), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18367) );
  OAI211_X1 U21254 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n18039), .A(
        n18038), .B(n18367), .ZN(n18040) );
  AOI221_X1 U21255 ( .B1(n18042), .B2(n18362), .C1(n18041), .C2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n18040), .ZN(n18043) );
  OAI21_X1 U21256 ( .B1(n18369), .B2(n18093), .A(n18043), .ZN(P3_U2818) );
  NAND2_X1 U21257 ( .A1(n18376), .A2(n18052), .ZN(n18384) );
  INV_X1 U21258 ( .A(n18044), .ZN(n18060) );
  OAI21_X1 U21259 ( .B1(n18138), .B2(n18045), .A(n18060), .ZN(n18048) );
  NAND2_X1 U21260 ( .A1(n18499), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n18382) );
  OAI21_X1 U21261 ( .B1(n18160), .B2(n18046), .A(n18382), .ZN(n18047) );
  AOI21_X1 U21262 ( .B1(n18049), .B2(n18048), .A(n18047), .ZN(n18054) );
  AOI22_X1 U21263 ( .A1(n18090), .A2(n18370), .B1(n18150), .B2(n18372), .ZN(
        n18077) );
  OAI21_X1 U21264 ( .B1(n18376), .B2(n9664), .A(n18077), .ZN(n18062) );
  AOI21_X1 U21265 ( .B1(n18376), .B2(n18068), .A(n18050), .ZN(n18051) );
  XOR2_X1 U21266 ( .A(n18052), .B(n18051), .Z(n18380) );
  AOI22_X1 U21267 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18062), .B1(
        n18075), .B2(n18380), .ZN(n18053) );
  OAI211_X1 U21268 ( .C1(n9664), .C2(n18384), .A(n18054), .B(n18053), .ZN(
        P3_U2819) );
  OAI21_X1 U21269 ( .B1(n18392), .B2(n18056), .A(n18055), .ZN(n18057) );
  XOR2_X1 U21270 ( .A(n18057), .B(n18378), .Z(n18391) );
  NOR3_X1 U21271 ( .A1(n18097), .A2(n18083), .A3(n18741), .ZN(n18071) );
  NAND2_X1 U21272 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n18071), .ZN(
        n18070) );
  OAI21_X1 U21273 ( .B1(n18138), .B2(n18058), .A(n18070), .ZN(n18059) );
  AOI22_X1 U21274 ( .A1(n18349), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18060), 
        .B2(n18059), .ZN(n18065) );
  OAI21_X1 U21275 ( .B1(n9664), .B2(n18392), .A(n18378), .ZN(n18061) );
  AOI22_X1 U21276 ( .A1(n18063), .A2(n18170), .B1(n18062), .B2(n18061), .ZN(
        n18064) );
  OAI211_X1 U21277 ( .C1(n18391), .C2(n18093), .A(n18065), .B(n18064), .ZN(
        P3_U2820) );
  NOR2_X1 U21278 ( .A1(n18066), .A2(n11255), .ZN(n18067) );
  NOR2_X1 U21279 ( .A1(n18068), .A2(n18067), .ZN(n18069) );
  XOR2_X1 U21280 ( .A(n18069), .B(n18392), .Z(n18398) );
  OAI211_X1 U21281 ( .C1(n18071), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n18171), .B(n18070), .ZN(n18072) );
  NAND2_X1 U21282 ( .A1(n18349), .A2(P3_REIP_REG_9__SCAN_IN), .ZN(n18400) );
  OAI211_X1 U21283 ( .C1(n18160), .C2(n18073), .A(n18072), .B(n18400), .ZN(
        n18074) );
  AOI21_X1 U21284 ( .B1(n18075), .B2(n18398), .A(n18074), .ZN(n18076) );
  OAI221_X1 U21285 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n9664), .C1(
        n18392), .C2(n18077), .A(n18076), .ZN(P3_U2821) );
  OAI21_X1 U21286 ( .B1(n18414), .B2(n18080), .A(n18079), .ZN(n18417) );
  OAI21_X1 U21287 ( .B1(n18082), .B2(n18081), .A(n18176), .ZN(n18100) );
  NOR2_X1 U21288 ( .A1(n18097), .A2(n18098), .ZN(n18084) );
  OAI211_X1 U21289 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18084), .A(
        n18545), .B(n18083), .ZN(n18085) );
  NAND2_X1 U21290 ( .A1(n18499), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n18408) );
  OAI211_X1 U21291 ( .C1(n18160), .C2(n18086), .A(n18085), .B(n18408), .ZN(
        n18087) );
  AOI21_X1 U21292 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18100), .A(
        n18087), .ZN(n18092) );
  AOI21_X1 U21293 ( .B1(n18089), .B2(n18278), .A(n18088), .ZN(n18412) );
  AOI22_X1 U21294 ( .A1(n18090), .A2(n18414), .B1(n18150), .B2(n18412), .ZN(
        n18091) );
  OAI211_X1 U21295 ( .C1(n18093), .C2(n18417), .A(n18092), .B(n18091), .ZN(
        P3_U2822) );
  NAND2_X1 U21296 ( .A1(n18095), .A2(n18094), .ZN(n18096) );
  XOR2_X1 U21297 ( .A(n18096), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18428) );
  NOR2_X1 U21298 ( .A1(n18097), .A2(n18741), .ZN(n18099) );
  NOR2_X1 U21299 ( .A1(n18482), .A2(n19078), .ZN(n18419) );
  AOI221_X1 U21300 ( .B1(n18100), .B2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C1(
        n18099), .C2(n18098), .A(n18419), .ZN(n18105) );
  INV_X1 U21301 ( .A(n11058), .ZN(n18101) );
  AOI21_X1 U21302 ( .B1(n18423), .B2(n18102), .A(n18101), .ZN(n18424) );
  AOI22_X1 U21303 ( .A1(n9729), .A2(n18424), .B1(n18103), .B2(n18170), .ZN(
        n18104) );
  OAI211_X1 U21304 ( .C1(n18180), .C2(n18428), .A(n18105), .B(n18104), .ZN(
        P3_U2823) );
  AOI21_X1 U21305 ( .B1(n18433), .B2(n18107), .A(n18106), .ZN(n18436) );
  NOR2_X1 U21306 ( .A1(n18112), .A2(n18741), .ZN(n18108) );
  AOI22_X1 U21307 ( .A1(n18150), .A2(n18436), .B1(n18108), .B2(n18113), .ZN(
        n18117) );
  AOI21_X1 U21308 ( .B1(n18111), .B2(n18110), .A(n18109), .ZN(n18435) );
  OAI21_X1 U21309 ( .B1(n18741), .B2(n18112), .A(n18171), .ZN(n18128) );
  OAI22_X1 U21310 ( .A1(n18160), .A2(n18114), .B1(n18113), .B2(n18128), .ZN(
        n18115) );
  AOI21_X1 U21311 ( .B1(n9729), .B2(n18435), .A(n18115), .ZN(n18116) );
  OAI211_X1 U21312 ( .C1(n18482), .C2(n19076), .A(n18117), .B(n18116), .ZN(
        P3_U2824) );
  NOR2_X1 U21313 ( .A1(n18118), .A2(n18132), .ZN(n18137) );
  AOI21_X1 U21314 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18137), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n18129) );
  AOI21_X1 U21315 ( .B1(n18121), .B2(n18120), .A(n18119), .ZN(n18440) );
  AOI22_X1 U21316 ( .A1(n18150), .A2(n18440), .B1(n18499), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n18127) );
  OAI21_X1 U21317 ( .B1(n18123), .B2(n9790), .A(n18122), .ZN(n18124) );
  XOR2_X1 U21318 ( .A(n18124), .B(n18439), .Z(n18441) );
  AOI22_X1 U21319 ( .A1(n9729), .A2(n18441), .B1(n18125), .B2(n18170), .ZN(
        n18126) );
  OAI211_X1 U21320 ( .C1(n18129), .C2(n18128), .A(n18127), .B(n18126), .ZN(
        P3_U2825) );
  AOI21_X1 U21321 ( .B1(n18450), .B2(n18131), .A(n18130), .ZN(n18454) );
  NOR3_X1 U21322 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18132), .A3(
        n18741), .ZN(n18133) );
  NOR2_X1 U21323 ( .A1(n18482), .A2(n19072), .ZN(n18453) );
  AOI211_X1 U21324 ( .C1(n9729), .C2(n18454), .A(n18133), .B(n18453), .ZN(
        n18140) );
  AOI21_X1 U21325 ( .B1(n18136), .B2(n18135), .A(n18134), .ZN(n18455) );
  NOR2_X1 U21326 ( .A1(n18138), .A2(n18137), .ZN(n18149) );
  AOI22_X1 U21327 ( .A1(n18150), .A2(n18455), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18149), .ZN(n18139) );
  OAI211_X1 U21328 ( .C1(n18160), .C2(n18141), .A(n18140), .B(n18139), .ZN(
        P3_U2826) );
  AOI21_X1 U21329 ( .B1(n18465), .B2(n18143), .A(n18142), .ZN(n18459) );
  AOI22_X1 U21330 ( .A1(n9729), .A2(n18459), .B1(n18499), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n18152) );
  AOI21_X1 U21331 ( .B1(n18146), .B2(n18145), .A(n18144), .ZN(n18462) );
  AOI21_X1 U21332 ( .B1(n18176), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18147) );
  INV_X1 U21333 ( .A(n18147), .ZN(n18148) );
  AOI22_X1 U21334 ( .A1(n18150), .A2(n18462), .B1(n18149), .B2(n18148), .ZN(
        n18151) );
  OAI211_X1 U21335 ( .C1(n18160), .C2(n18153), .A(n18152), .B(n18151), .ZN(
        P3_U2827) );
  AOI21_X1 U21336 ( .B1(n18156), .B2(n18155), .A(n18154), .ZN(n18478) );
  NOR2_X1 U21337 ( .A1(n18482), .A2(n19068), .ZN(n18477) );
  XNOR2_X1 U21338 ( .A(n18158), .B(n18157), .ZN(n18475) );
  OAI22_X1 U21339 ( .A1(n18160), .A2(n18159), .B1(n18180), .B2(n18475), .ZN(
        n18161) );
  AOI211_X1 U21340 ( .C1(n9729), .C2(n18478), .A(n18477), .B(n18161), .ZN(
        n18162) );
  OAI221_X1 U21341 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18741), .C1(
        n18163), .C2(n18176), .A(n18162), .ZN(P3_U2828) );
  NAND2_X1 U21342 ( .A1(n19163), .A2(n18164), .ZN(n18165) );
  XNOR2_X1 U21343 ( .A(n18165), .B(n18167), .ZN(n18493) );
  AOI21_X1 U21344 ( .B1(n18174), .B2(n18167), .A(n18166), .ZN(n18486) );
  AOI22_X1 U21345 ( .A1(n9729), .A2(n18486), .B1(n18499), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18173) );
  AOI22_X1 U21346 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18171), .B1(
        n18170), .B2(n18169), .ZN(n18172) );
  OAI211_X1 U21347 ( .C1(n18493), .C2(n18180), .A(n18173), .B(n18172), .ZN(
        P3_U2829) );
  OAI21_X1 U21348 ( .B1(n18175), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18174), .ZN(n18502) );
  INV_X1 U21349 ( .A(n18502), .ZN(n18181) );
  OAI21_X1 U21350 ( .B1(n19033), .B2(n19189), .A(n18176), .ZN(n18177) );
  AOI22_X1 U21351 ( .A1(n18349), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18177), .ZN(n18178) );
  OAI221_X1 U21352 ( .B1(n18181), .B2(n18180), .C1(n18502), .C2(n18179), .A(
        n18178), .ZN(P3_U2830) );
  OAI21_X1 U21353 ( .B1(n18494), .B2(n18196), .A(n18182), .ZN(n18192) );
  NOR2_X1 U21354 ( .A1(n18992), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18472) );
  NOR2_X1 U21355 ( .A1(n18472), .A2(n18183), .ZN(n18282) );
  INV_X1 U21356 ( .A(n18447), .ZN(n18470) );
  AOI21_X1 U21357 ( .B1(n18282), .B2(n18184), .A(n18470), .ZN(n18204) );
  OAI21_X1 U21358 ( .B1(n18188), .B2(n18354), .A(n18187), .ZN(n18189) );
  AOI21_X1 U21359 ( .B1(n18966), .B2(n18190), .A(n18189), .ZN(n18197) );
  OAI211_X1 U21360 ( .C1(n19004), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n18197), .ZN(n18191) );
  AOI22_X1 U21361 ( .A1(n18399), .A2(n18193), .B1(n18192), .B2(n18191), .ZN(
        n18195) );
  OAI211_X1 U21362 ( .C1(n18495), .C2(n18196), .A(n18195), .B(n18194), .ZN(
        P3_U2835) );
  INV_X1 U21363 ( .A(n18255), .ZN(n18237) );
  OAI21_X1 U21364 ( .B1(n18197), .B2(n18494), .A(n18495), .ZN(n18199) );
  AOI22_X1 U21365 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18199), .B1(
        n18399), .B2(n18198), .ZN(n18201) );
  NAND2_X1 U21366 ( .A1(n18499), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n18200) );
  OAI211_X1 U21367 ( .C1(n18202), .C2(n18237), .A(n18201), .B(n18200), .ZN(
        P3_U2836) );
  NAND3_X1 U21368 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n18203), .ZN(n18205) );
  AOI21_X1 U21369 ( .B1(n19000), .B2(n18205), .A(n18204), .ZN(n18208) );
  NAND4_X1 U21370 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n18218), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A4(n18206), .ZN(n18207) );
  AOI221_X1 U21371 ( .B1(n18208), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n18207), .C2(n11067), .A(n18494), .ZN(n18209) );
  AOI211_X1 U21372 ( .C1(n18489), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n18210), .B(n18209), .ZN(n18214) );
  AOI22_X1 U21373 ( .A1(n18498), .A2(n18212), .B1(n18399), .B2(n18211), .ZN(
        n18213) );
  OAI211_X1 U21374 ( .C1(n18345), .C2(n18215), .A(n18214), .B(n18213), .ZN(
        P3_U2837) );
  AOI22_X1 U21375 ( .A1(n18399), .A2(n18217), .B1(n18255), .B2(n18216), .ZN(
        n18228) );
  AOI21_X1 U21376 ( .B1(n18218), .B2(n18282), .A(n18470), .ZN(n18219) );
  OAI21_X1 U21377 ( .B1(n18222), .B2(n18354), .A(n18221), .ZN(n18226) );
  AOI211_X1 U21378 ( .C1(n19000), .C2(n18224), .A(n18223), .B(n18226), .ZN(
        n18225) );
  NOR2_X1 U21379 ( .A1(n18499), .A2(n18225), .ZN(n18232) );
  OAI211_X1 U21380 ( .C1(n18407), .C2(n18226), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n18232), .ZN(n18227) );
  OAI211_X1 U21381 ( .C1(n19112), .C2(n18482), .A(n18228), .B(n18227), .ZN(
        P3_U2838) );
  INV_X1 U21382 ( .A(n18229), .ZN(n18236) );
  NAND2_X1 U21383 ( .A1(n18499), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n18235) );
  NOR3_X1 U21384 ( .A1(n18489), .A2(n18231), .A3(n18230), .ZN(n18233) );
  OAI21_X1 U21385 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n18233), .A(
        n18232), .ZN(n18234) );
  OAI211_X1 U21386 ( .C1(n18236), .C2(n18418), .A(n18235), .B(n18234), .ZN(
        P3_U2839) );
  OAI22_X1 U21387 ( .A1(n18239), .A2(n18494), .B1(n18238), .B2(n18237), .ZN(
        n18251) );
  OAI22_X1 U21388 ( .A1(n18242), .A2(n18354), .B1(n18241), .B2(n18240), .ZN(
        n18306) );
  AOI221_X1 U21389 ( .B1(n18244), .B2(n19000), .C1(n18243), .C2(n19000), .A(
        n18306), .ZN(n18245) );
  OAI221_X1 U21390 ( .B1(n19004), .B2(n18246), .C1(n19004), .C2(n18268), .A(
        n18245), .ZN(n18265) );
  NOR2_X1 U21391 ( .A1(n18966), .A2(n18371), .ZN(n18375) );
  OAI22_X1 U21392 ( .A1(n19004), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n18247), .B2(n18375), .ZN(n18248) );
  AOI22_X1 U21393 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18489), .B1(
        n18251), .B2(n18250), .ZN(n18253) );
  NAND2_X1 U21394 ( .A1(n18499), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n18252) );
  OAI211_X1 U21395 ( .C1(n18254), .C2(n18418), .A(n18253), .B(n18252), .ZN(
        P3_U2840) );
  NAND2_X1 U21396 ( .A1(n18255), .A2(n18257), .ZN(n18277) );
  AOI22_X1 U21397 ( .A1(n18349), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18399), 
        .B2(n18256), .ZN(n18262) );
  OAI221_X1 U21398 ( .B1(n18992), .B2(n18299), .C1(n18992), .C2(n18257), .A(
        n18429), .ZN(n18266) );
  NAND2_X1 U21399 ( .A1(n18469), .A2(n18992), .ZN(n18332) );
  INV_X1 U21400 ( .A(n18332), .ZN(n18488) );
  OAI21_X1 U21401 ( .B1(n18259), .B2(n18488), .A(n18258), .ZN(n18260) );
  OAI211_X1 U21402 ( .C1(n18266), .C2(n18260), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18482), .ZN(n18261) );
  OAI211_X1 U21403 ( .C1(n18263), .C2(n18277), .A(n18262), .B(n18261), .ZN(
        P3_U2841) );
  AOI22_X1 U21404 ( .A1(n18349), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n18399), 
        .B2(n18264), .ZN(n18271) );
  NOR2_X1 U21405 ( .A1(n18266), .A2(n18265), .ZN(n18267) );
  AOI221_X1 U21406 ( .B1(n18268), .B2(n18267), .C1(n18375), .C2(n18267), .A(
        n18349), .ZN(n18274) );
  NOR3_X1 U21407 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18488), .A3(
        n19029), .ZN(n18269) );
  OAI21_X1 U21408 ( .B1(n18274), .B2(n18269), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n18270) );
  OAI211_X1 U21409 ( .C1(n18277), .C2(n18272), .A(n18271), .B(n18270), .ZN(
        P3_U2842) );
  AOI22_X1 U21410 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18274), .B1(
        n18399), .B2(n18273), .ZN(n18276) );
  OAI211_X1 U21411 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n18277), .A(
        n18276), .B(n18275), .ZN(P3_U2843) );
  OAI22_X1 U21412 ( .A1(n18448), .A2(n18469), .B1(n18446), .B2(n18467), .ZN(
        n18460) );
  NAND3_X1 U21413 ( .A1(n18429), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18460), .ZN(n18458) );
  NOR3_X1 U21414 ( .A1(n18450), .A2(n18439), .A3(n18458), .ZN(n18434) );
  NAND3_X1 U21415 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n18434), .ZN(n18409) );
  AOI22_X1 U21416 ( .A1(n18280), .A2(n18347), .B1(n18429), .B2(n18279), .ZN(
        n18311) );
  AOI22_X1 U21417 ( .A1(n18349), .A2(P3_REIP_REG_18__SCAN_IN), .B1(n18399), 
        .B2(n18281), .ZN(n18289) );
  AOI21_X1 U21418 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18282), .A(
        n18470), .ZN(n18283) );
  AOI211_X1 U21419 ( .C1(n19000), .C2(n18284), .A(n18283), .B(n18306), .ZN(
        n18285) );
  OAI21_X1 U21420 ( .B1(n18286), .B2(n18375), .A(n18285), .ZN(n18291) );
  OAI21_X1 U21421 ( .B1(n18470), .B2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n18429), .ZN(n18287) );
  OAI211_X1 U21422 ( .C1(n18291), .C2(n18287), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B(n18482), .ZN(n18288) );
  OAI211_X1 U21423 ( .C1(n18311), .C2(n18290), .A(n18289), .B(n18288), .ZN(
        P3_U2844) );
  AOI21_X1 U21424 ( .B1(n18291), .B2(n18429), .A(n18489), .ZN(n18292) );
  INV_X1 U21425 ( .A(n18292), .ZN(n18294) );
  OAI21_X1 U21426 ( .B1(n18310), .B2(n18311), .A(n18295), .ZN(n18293) );
  OAI21_X1 U21427 ( .B1(n18295), .B2(n18294), .A(n18293), .ZN(n18297) );
  OAI211_X1 U21428 ( .C1(n18298), .C2(n18418), .A(n18297), .B(n18296), .ZN(
        P3_U2845) );
  AOI21_X1 U21429 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18992), .A(
        n18299), .ZN(n18302) );
  AOI22_X1 U21430 ( .A1(n18977), .A2(n18301), .B1(n18300), .B2(n19000), .ZN(
        n18395) );
  INV_X1 U21431 ( .A(n18395), .ZN(n18327) );
  AOI211_X1 U21432 ( .C1(n18304), .C2(n18303), .A(n18302), .B(n18327), .ZN(
        n18317) );
  OAI21_X1 U21433 ( .B1(n18451), .B2(n18317), .A(n18495), .ZN(n18305) );
  OAI21_X1 U21434 ( .B1(n18306), .B2(n18305), .A(n18482), .ZN(n18309) );
  AOI22_X1 U21435 ( .A1(n18499), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18399), 
        .B2(n18307), .ZN(n18308) );
  OAI221_X1 U21436 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18311), 
        .C1(n18310), .C2(n18309), .A(n18308), .ZN(P3_U2846) );
  NAND2_X1 U21437 ( .A1(n18966), .A2(n18312), .ZN(n18322) );
  NAND2_X1 U21438 ( .A1(n18371), .A2(n18313), .ZN(n18320) );
  AND3_X1 U21439 ( .A1(n18460), .A2(n18420), .A3(n18314), .ZN(n18315) );
  AOI21_X1 U21440 ( .B1(n18316), .B2(n18315), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18318) );
  OAI222_X1 U21441 ( .A1(n18322), .A2(n18321), .B1(n18320), .B2(n18319), .C1(
        n18318), .C2(n18317), .ZN(n18323) );
  AOI22_X1 U21442 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18489), .B1(
        n18429), .B2(n18323), .ZN(n18325) );
  OAI211_X1 U21443 ( .C1(n18418), .C2(n18326), .A(n18325), .B(n18324), .ZN(
        P3_U2847) );
  AOI211_X1 U21444 ( .C1(n18977), .C2(n18329), .A(n18328), .B(n18327), .ZN(
        n18330) );
  NAND2_X1 U21445 ( .A1(n19002), .A2(n18373), .ZN(n18393) );
  OAI211_X1 U21446 ( .C1(n18331), .C2(n18488), .A(n18330), .B(n18393), .ZN(
        n18336) );
  AOI21_X1 U21447 ( .B1(n18333), .B2(n18332), .A(n18336), .ZN(n18334) );
  OAI21_X1 U21448 ( .B1(n18334), .B2(n18494), .A(n18495), .ZN(n18339) );
  AND3_X1 U21449 ( .A1(n18336), .A2(n18347), .A3(n18335), .ZN(n18338) );
  AOI211_X1 U21450 ( .C1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18339), .A(
        n18338), .B(n18337), .ZN(n18343) );
  AOI22_X1 U21451 ( .A1(n18498), .A2(n18341), .B1(n18399), .B2(n18340), .ZN(
        n18342) );
  OAI211_X1 U21452 ( .C1(n18345), .C2(n18344), .A(n18343), .B(n18342), .ZN(
        P3_U2848) );
  OAI22_X1 U21453 ( .A1(n18372), .A2(n18492), .B1(n18370), .B2(n18345), .ZN(
        n18346) );
  AOI22_X1 U21454 ( .A1(n18349), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18399), 
        .B2(n18348), .ZN(n18360) );
  INV_X1 U21455 ( .A(n18350), .ZN(n18357) );
  AOI21_X1 U21456 ( .B1(n18351), .B2(n18395), .A(n18386), .ZN(n18377) );
  OAI21_X1 U21457 ( .B1(n18352), .B2(n18373), .A(n19002), .ZN(n18353) );
  OAI21_X1 U21458 ( .B1(n18355), .B2(n18354), .A(n18353), .ZN(n18356) );
  OAI211_X1 U21459 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18386), .A(
        n18429), .B(n18364), .ZN(n18358) );
  NAND3_X1 U21460 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18482), .A3(
        n18358), .ZN(n18359) );
  OAI211_X1 U21461 ( .C1(n18402), .C2(n18361), .A(n18360), .B(n18359), .ZN(
        P3_U2849) );
  OAI22_X1 U21462 ( .A1(n18402), .A2(n18363), .B1(n18362), .B2(n18494), .ZN(
        n18366) );
  NAND2_X1 U21463 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18364), .ZN(
        n18365) );
  AOI22_X1 U21464 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18489), .B1(
        n18366), .B2(n18365), .ZN(n18368) );
  OAI211_X1 U21465 ( .C1(n18369), .C2(n18418), .A(n18368), .B(n18367), .ZN(
        P3_U2850) );
  AOI22_X1 U21466 ( .A1(n18966), .A2(n18372), .B1(n18371), .B2(n18370), .ZN(
        n18394) );
  OAI21_X1 U21467 ( .B1(n18392), .B2(n18373), .A(n19002), .ZN(n18374) );
  OAI211_X1 U21468 ( .C1(n18376), .C2(n18375), .A(n18394), .B(n18374), .ZN(
        n18388) );
  OAI21_X1 U21469 ( .B1(n18379), .B2(n18494), .A(n18495), .ZN(n18381) );
  AOI22_X1 U21470 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18381), .B1(
        n18399), .B2(n18380), .ZN(n18383) );
  OAI211_X1 U21471 ( .C1(n18402), .C2(n18384), .A(n18383), .B(n18382), .ZN(
        P3_U2851) );
  NOR3_X1 U21472 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18402), .A3(
        n18392), .ZN(n18385) );
  AOI21_X1 U21473 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n18499), .A(n18385), 
        .ZN(n18390) );
  OAI211_X1 U21474 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18386), .A(
        n18429), .B(n18395), .ZN(n18387) );
  OAI211_X1 U21475 ( .C1(n18388), .C2(n18387), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18482), .ZN(n18389) );
  OAI211_X1 U21476 ( .C1(n18391), .C2(n18418), .A(n18390), .B(n18389), .ZN(
        P3_U2852) );
  NOR2_X1 U21477 ( .A1(n18499), .A2(n18392), .ZN(n18397) );
  NAND4_X1 U21478 ( .A1(n18395), .A2(n18429), .A3(n18394), .A4(n18393), .ZN(
        n18396) );
  AOI22_X1 U21479 ( .A1(n18399), .A2(n18398), .B1(n18397), .B2(n18396), .ZN(
        n18401) );
  OAI211_X1 U21480 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18402), .A(
        n18401), .B(n18400), .ZN(P3_U2853) );
  INV_X1 U21481 ( .A(n18403), .ZN(n18404) );
  OAI21_X1 U21482 ( .B1(n18472), .B2(n18404), .A(n18447), .ZN(n18405) );
  OAI21_X1 U21483 ( .B1(n18406), .B2(n18469), .A(n18405), .ZN(n18430) );
  AOI211_X1 U21484 ( .C1(n18407), .C2(n18433), .A(n18423), .B(n18430), .ZN(
        n18421) );
  OAI21_X1 U21485 ( .B1(n18421), .B2(n18483), .A(n18495), .ZN(n18411) );
  OAI21_X1 U21486 ( .B1(n18409), .B2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n18408), .ZN(n18410) );
  AOI21_X1 U21487 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n18411), .A(
        n18410), .ZN(n18416) );
  AOI22_X1 U21488 ( .A1(n18414), .A2(n18413), .B1(n18498), .B2(n18412), .ZN(
        n18415) );
  OAI211_X1 U21489 ( .C1(n18418), .C2(n18417), .A(n18416), .B(n18415), .ZN(
        P3_U2854) );
  AOI21_X1 U21490 ( .B1(n18489), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18419), .ZN(n18427) );
  NAND2_X1 U21491 ( .A1(n18420), .A2(n18460), .ZN(n18422) );
  AOI221_X1 U21492 ( .B1(n18433), .B2(n18423), .C1(n18422), .C2(n18423), .A(
        n18421), .ZN(n18425) );
  AOI22_X1 U21493 ( .A1(n18429), .A2(n18425), .B1(n18487), .B2(n18424), .ZN(
        n18426) );
  OAI211_X1 U21494 ( .C1(n18492), .C2(n18428), .A(n18427), .B(n18426), .ZN(
        P3_U2855) );
  AOI21_X1 U21495 ( .B1(n18430), .B2(n18429), .A(n18489), .ZN(n18431) );
  INV_X1 U21496 ( .A(n18431), .ZN(n18442) );
  NOR2_X1 U21497 ( .A1(n18482), .A2(n19076), .ZN(n18432) );
  AOI221_X1 U21498 ( .B1(n18434), .B2(n18433), .C1(n18442), .C2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n18432), .ZN(n18438) );
  AOI22_X1 U21499 ( .A1(n18498), .A2(n18436), .B1(n18487), .B2(n18435), .ZN(
        n18437) );
  NAND2_X1 U21500 ( .A1(n18438), .A2(n18437), .ZN(P3_U2856) );
  NAND2_X1 U21501 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18439), .ZN(
        n18445) );
  AOI22_X1 U21502 ( .A1(n18499), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18498), 
        .B2(n18440), .ZN(n18444) );
  AOI22_X1 U21503 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18442), .B1(
        n18487), .B2(n18441), .ZN(n18443) );
  OAI211_X1 U21504 ( .C1(n18458), .C2(n18445), .A(n18444), .B(n18443), .ZN(
        P3_U2857) );
  AOI211_X1 U21505 ( .C1(n18447), .C2(n18446), .A(n18472), .B(n18465), .ZN(
        n18449) );
  NAND2_X1 U21506 ( .A1(n19000), .A2(n18448), .ZN(n18480) );
  AOI21_X1 U21507 ( .B1(n18449), .B2(n18480), .A(n18494), .ZN(n18461) );
  NOR2_X1 U21508 ( .A1(n18489), .A2(n18461), .ZN(n18466) );
  AOI211_X1 U21509 ( .C1(n18451), .C2(n18495), .A(n18466), .B(n18450), .ZN(
        n18452) );
  AOI211_X1 U21510 ( .C1(n18487), .C2(n18454), .A(n18453), .B(n18452), .ZN(
        n18457) );
  NAND2_X1 U21511 ( .A1(n18498), .A2(n18455), .ZN(n18456) );
  OAI211_X1 U21512 ( .C1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n18458), .A(
        n18457), .B(n18456), .ZN(P3_U2858) );
  AOI22_X1 U21513 ( .A1(n18499), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18487), 
        .B2(n18459), .ZN(n18464) );
  AOI22_X1 U21514 ( .A1(n18498), .A2(n18462), .B1(n18461), .B2(n18460), .ZN(
        n18463) );
  OAI211_X1 U21515 ( .C1(n18466), .C2(n18465), .A(n18464), .B(n18463), .ZN(
        P3_U2859) );
  OR2_X1 U21516 ( .A1(n19145), .A2(n18467), .ZN(n18474) );
  NAND2_X1 U21517 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18468) );
  OAI22_X1 U21518 ( .A1(n18470), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n18469), .B2(n18468), .ZN(n18471) );
  NOR2_X1 U21519 ( .A1(n18472), .A2(n18471), .ZN(n18473) );
  MUX2_X1 U21520 ( .A(n18474), .B(n18473), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n18481) );
  OAI22_X1 U21521 ( .A1(n11027), .A2(n18495), .B1(n18492), .B2(n18475), .ZN(
        n18476) );
  AOI211_X1 U21522 ( .C1(n18487), .C2(n18478), .A(n18477), .B(n18476), .ZN(
        n18479) );
  OAI221_X1 U21523 ( .B1(n18494), .B2(n18481), .C1(n18494), .C2(n18480), .A(
        n18479), .ZN(P3_U2860) );
  NOR2_X1 U21524 ( .A1(n18482), .A2(n19067), .ZN(n18485) );
  AOI211_X1 U21525 ( .C1(n19004), .C2(n19163), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18483), .ZN(n18484) );
  AOI211_X1 U21526 ( .C1(n18487), .C2(n18486), .A(n18485), .B(n18484), .ZN(
        n18491) );
  NOR3_X1 U21527 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18488), .A3(
        n18494), .ZN(n18497) );
  OAI21_X1 U21528 ( .B1(n18489), .B2(n18497), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18490) );
  OAI211_X1 U21529 ( .C1(n18493), .C2(n18492), .A(n18491), .B(n18490), .ZN(
        P3_U2861) );
  AOI221_X1 U21530 ( .B1(n19004), .B2(n18495), .C1(n18494), .C2(n18495), .A(
        n19163), .ZN(n18496) );
  AOI211_X1 U21531 ( .C1(n18498), .C2(n18502), .A(n18497), .B(n18496), .ZN(
        n18501) );
  NAND2_X1 U21532 ( .A1(n18499), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18500) );
  OAI211_X1 U21533 ( .C1(n18503), .C2(n18502), .A(n18501), .B(n18500), .ZN(
        P3_U2862) );
  AOI21_X1 U21534 ( .B1(n18506), .B2(n18505), .A(n18504), .ZN(n19030) );
  OAI21_X1 U21535 ( .B1(n19030), .B2(n18552), .A(n18511), .ZN(n18507) );
  OAI221_X1 U21536 ( .B1(n19008), .B2(n19179), .C1(n19008), .C2(n18511), .A(
        n18507), .ZN(P3_U2863) );
  NAND2_X1 U21537 ( .A1(n19015), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18819) );
  INV_X1 U21538 ( .A(n18819), .ZN(n18796) );
  NAND2_X1 U21539 ( .A1(n19018), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18645) );
  INV_X1 U21540 ( .A(n18645), .ZN(n18694) );
  NOR2_X1 U21541 ( .A1(n18796), .A2(n18694), .ZN(n18509) );
  OAI22_X1 U21542 ( .A1(n18510), .A2(n19018), .B1(n18509), .B2(n18508), .ZN(
        P3_U2866) );
  NOR2_X1 U21543 ( .A1(n19019), .A2(n18511), .ZN(P3_U2867) );
  NOR2_X2 U21544 ( .A1(n18741), .A2(n14436), .ZN(n18909) );
  INV_X1 U21545 ( .A(n18909), .ZN(n18853) );
  NAND2_X1 U21546 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18513) );
  NAND2_X1 U21547 ( .A1(n19008), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18771) );
  NOR2_X2 U21548 ( .A1(n18513), .A2(n18771), .ZN(n18901) );
  INV_X1 U21549 ( .A(n18901), .ZN(n18571) );
  INV_X1 U21550 ( .A(n18667), .ZN(n18879) );
  NOR2_X1 U21551 ( .A1(n19018), .A2(n18512), .ZN(n18911) );
  NAND2_X1 U21552 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18911), .ZN(
        n18593) );
  NOR2_X1 U21553 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18715) );
  NOR2_X1 U21554 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18599) );
  NAND2_X1 U21555 ( .A1(n18715), .A2(n18599), .ZN(n18619) );
  NAND2_X1 U21556 ( .A1(n18593), .A2(n18619), .ZN(n18514) );
  INV_X1 U21557 ( .A(n18514), .ZN(n18572) );
  NOR2_X1 U21558 ( .A1(n19042), .A2(n18572), .ZN(n18546) );
  NOR2_X1 U21559 ( .A1(n18513), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18912) );
  NAND2_X1 U21560 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18912), .ZN(
        n18965) );
  INV_X1 U21561 ( .A(n18965), .ZN(n18943) );
  NAND2_X1 U21562 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18545), .ZN(n18916) );
  INV_X1 U21563 ( .A(n18916), .ZN(n18849) );
  AOI22_X1 U21564 ( .A1(n18908), .A2(n18546), .B1(n18943), .B2(n18849), .ZN(
        n18519) );
  NAND2_X1 U21565 ( .A1(n19010), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18743) );
  AND2_X1 U21566 ( .A1(n18771), .A2(n18743), .ZN(n18820) );
  NOR2_X1 U21567 ( .A1(n18820), .A2(n18513), .ZN(n18874) );
  AOI21_X1 U21568 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18667), .ZN(n18821) );
  AOI22_X1 U21569 ( .A1(n18545), .A2(n18874), .B1(n18821), .B2(n18514), .ZN(
        n18549) );
  INV_X1 U21570 ( .A(n18619), .ZN(n18612) );
  NAND2_X1 U21571 ( .A1(n18516), .A2(n18515), .ZN(n18547) );
  NOR2_X2 U21572 ( .A1(n18517), .A2(n18547), .ZN(n18913) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18549), .B1(
        n18612), .B2(n18913), .ZN(n18518) );
  OAI211_X1 U21574 ( .C1(n18853), .C2(n18571), .A(n18519), .B(n18518), .ZN(
        P3_U2868) );
  NAND2_X1 U21575 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18545), .ZN(n18922) );
  NAND2_X1 U21576 ( .A1(n18545), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18857) );
  INV_X1 U21577 ( .A(n18857), .ZN(n18918) );
  INV_X1 U21578 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18520) );
  NOR2_X2 U21579 ( .A1(n18667), .A2(n18520), .ZN(n18917) );
  AOI22_X1 U21580 ( .A1(n18901), .A2(n18918), .B1(n18546), .B2(n18917), .ZN(
        n18522) );
  NOR2_X2 U21581 ( .A1(n19186), .A2(n18547), .ZN(n18919) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18549), .B1(
        n18612), .B2(n18919), .ZN(n18521) );
  OAI211_X1 U21583 ( .C1(n18965), .C2(n18922), .A(n18522), .B(n18521), .ZN(
        P3_U2869) );
  NAND2_X1 U21584 ( .A1(n18545), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18887) );
  NOR2_X2 U21585 ( .A1(n18667), .A2(n18523), .ZN(n18923) );
  NAND2_X1 U21586 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18545), .ZN(n18928) );
  INV_X1 U21587 ( .A(n18928), .ZN(n18884) );
  AOI22_X1 U21588 ( .A1(n18546), .A2(n18923), .B1(n18943), .B2(n18884), .ZN(
        n18526) );
  NOR2_X2 U21589 ( .A1(n18524), .A2(n18547), .ZN(n18925) );
  AOI22_X1 U21590 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18549), .B1(
        n18612), .B2(n18925), .ZN(n18525) );
  OAI211_X1 U21591 ( .C1(n18571), .C2(n18887), .A(n18526), .B(n18525), .ZN(
        P3_U2870) );
  NOR2_X1 U21592 ( .A1(n18741), .A2(n18527), .ZN(n18930) );
  INV_X1 U21593 ( .A(n18930), .ZN(n18833) );
  NOR2_X2 U21594 ( .A1(n18667), .A2(n18528), .ZN(n18929) );
  NAND2_X1 U21595 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18545), .ZN(n18934) );
  INV_X1 U21596 ( .A(n18934), .ZN(n18830) );
  AOI22_X1 U21597 ( .A1(n18546), .A2(n18929), .B1(n18943), .B2(n18830), .ZN(
        n18531) );
  NOR2_X2 U21598 ( .A1(n18529), .A2(n18547), .ZN(n18931) );
  AOI22_X1 U21599 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18549), .B1(
        n18612), .B2(n18931), .ZN(n18530) );
  OAI211_X1 U21600 ( .C1(n18571), .C2(n18833), .A(n18531), .B(n18530), .ZN(
        P3_U2871) );
  NAND2_X1 U21601 ( .A1(n18545), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18940) );
  NOR2_X2 U21602 ( .A1(n18667), .A2(n18532), .ZN(n18935) );
  NAND2_X1 U21603 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18545), .ZN(n18808) );
  INV_X1 U21604 ( .A(n18808), .ZN(n18936) );
  AOI22_X1 U21605 ( .A1(n18546), .A2(n18935), .B1(n18943), .B2(n18936), .ZN(
        n18535) );
  NOR2_X2 U21606 ( .A1(n18533), .A2(n18547), .ZN(n18937) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18549), .B1(
        n18612), .B2(n18937), .ZN(n18534) );
  OAI211_X1 U21608 ( .C1(n18571), .C2(n18940), .A(n18535), .B(n18534), .ZN(
        P3_U2872) );
  INV_X1 U21609 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18536) );
  NOR2_X1 U21610 ( .A1(n18536), .A2(n18741), .ZN(n18836) );
  INV_X1 U21611 ( .A(n18836), .ZN(n18948) );
  NAND2_X1 U21612 ( .A1(n18545), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18839) );
  INV_X1 U21613 ( .A(n18839), .ZN(n18942) );
  NOR2_X2 U21614 ( .A1(n18667), .A2(n18537), .ZN(n18941) );
  AOI22_X1 U21615 ( .A1(n18901), .A2(n18942), .B1(n18546), .B2(n18941), .ZN(
        n18540) );
  NOR2_X2 U21616 ( .A1(n18538), .A2(n18547), .ZN(n18944) );
  AOI22_X1 U21617 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18549), .B1(
        n18612), .B2(n18944), .ZN(n18539) );
  OAI211_X1 U21618 ( .C1(n18965), .C2(n18948), .A(n18540), .B(n18539), .ZN(
        P3_U2873) );
  NOR2_X1 U21619 ( .A1(n19558), .A2(n18741), .ZN(n18950) );
  INV_X1 U21620 ( .A(n18950), .ZN(n18898) );
  NAND2_X1 U21621 ( .A1(n18545), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18954) );
  INV_X1 U21622 ( .A(n18954), .ZN(n18895) );
  NOR2_X2 U21623 ( .A1(n18667), .A2(n18541), .ZN(n18949) );
  AOI22_X1 U21624 ( .A1(n18901), .A2(n18895), .B1(n18546), .B2(n18949), .ZN(
        n18544) );
  NOR2_X2 U21625 ( .A1(n18542), .A2(n18547), .ZN(n18951) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18549), .B1(
        n18612), .B2(n18951), .ZN(n18543) );
  OAI211_X1 U21627 ( .C1(n18965), .C2(n18898), .A(n18544), .B(n18543), .ZN(
        P3_U2874) );
  NAND2_X1 U21628 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18545), .ZN(n18964) );
  AND2_X1 U21629 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18879), .ZN(n18956) );
  NAND2_X1 U21630 ( .A1(n18545), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18906) );
  INV_X1 U21631 ( .A(n18906), .ZN(n18958) );
  AOI22_X1 U21632 ( .A1(n18546), .A2(n18956), .B1(n18943), .B2(n18958), .ZN(
        n18551) );
  NOR2_X2 U21633 ( .A1(n18548), .A2(n18547), .ZN(n18959) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18549), .B1(
        n18612), .B2(n18959), .ZN(n18550) );
  OAI211_X1 U21635 ( .C1(n18571), .C2(n18964), .A(n18551), .B(n18550), .ZN(
        P3_U2875) );
  INV_X1 U21636 ( .A(n18599), .ZN(n18598) );
  NAND2_X1 U21637 ( .A1(n19010), .A2(n18795), .ZN(n18742) );
  NOR2_X1 U21638 ( .A1(n18598), .A2(n18742), .ZN(n18567) );
  AOI22_X1 U21639 ( .A1(n18909), .A2(n18960), .B1(n18908), .B2(n18567), .ZN(
        n18554) );
  NOR2_X1 U21640 ( .A1(n18667), .A2(n18552), .ZN(n18910) );
  INV_X1 U21641 ( .A(n18910), .ZN(n18739) );
  NOR2_X1 U21642 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18739), .ZN(
        n18643) );
  AOI22_X1 U21643 ( .A1(n18545), .A2(n18911), .B1(n18599), .B2(n18643), .ZN(
        n18568) );
  NOR2_X1 U21644 ( .A1(n18598), .A2(n18743), .ZN(n18635) );
  AOI22_X1 U21645 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18568), .B1(
        n18913), .B2(n18635), .ZN(n18553) );
  OAI211_X1 U21646 ( .C1(n18571), .C2(n18916), .A(n18554), .B(n18553), .ZN(
        P3_U2876) );
  AOI22_X1 U21647 ( .A1(n18960), .A2(n18918), .B1(n18917), .B2(n18567), .ZN(
        n18556) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18568), .B1(
        n18919), .B2(n18635), .ZN(n18555) );
  OAI211_X1 U21649 ( .C1(n18571), .C2(n18922), .A(n18556), .B(n18555), .ZN(
        P3_U2877) );
  AOI22_X1 U21650 ( .A1(n18901), .A2(n18884), .B1(n18923), .B2(n18567), .ZN(
        n18558) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18568), .B1(
        n18925), .B2(n18639), .ZN(n18557) );
  OAI211_X1 U21652 ( .C1(n18593), .C2(n18887), .A(n18558), .B(n18557), .ZN(
        P3_U2878) );
  AOI22_X1 U21653 ( .A1(n18960), .A2(n18930), .B1(n18929), .B2(n18567), .ZN(
        n18560) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18568), .B1(
        n18931), .B2(n18639), .ZN(n18559) );
  OAI211_X1 U21655 ( .C1(n18571), .C2(n18934), .A(n18560), .B(n18559), .ZN(
        P3_U2879) );
  INV_X1 U21656 ( .A(n18940), .ZN(n18805) );
  AOI22_X1 U21657 ( .A1(n18960), .A2(n18805), .B1(n18935), .B2(n18567), .ZN(
        n18562) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18568), .B1(
        n18937), .B2(n18635), .ZN(n18561) );
  OAI211_X1 U21659 ( .C1(n18571), .C2(n18808), .A(n18562), .B(n18561), .ZN(
        P3_U2880) );
  AOI22_X1 U21660 ( .A1(n18901), .A2(n18836), .B1(n18941), .B2(n18567), .ZN(
        n18564) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18568), .B1(
        n18944), .B2(n18635), .ZN(n18563) );
  OAI211_X1 U21662 ( .C1(n18593), .C2(n18839), .A(n18564), .B(n18563), .ZN(
        P3_U2881) );
  AOI22_X1 U21663 ( .A1(n18960), .A2(n18895), .B1(n18949), .B2(n18567), .ZN(
        n18566) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18568), .B1(
        n18951), .B2(n18639), .ZN(n18565) );
  OAI211_X1 U21665 ( .C1(n18571), .C2(n18898), .A(n18566), .B(n18565), .ZN(
        P3_U2882) );
  INV_X1 U21666 ( .A(n18964), .ZN(n18900) );
  AOI22_X1 U21667 ( .A1(n18960), .A2(n18900), .B1(n18956), .B2(n18567), .ZN(
        n18570) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18568), .B1(
        n18959), .B2(n18639), .ZN(n18569) );
  OAI211_X1 U21669 ( .C1(n18571), .C2(n18906), .A(n18570), .B(n18569), .ZN(
        P3_U2883) );
  NOR2_X2 U21670 ( .A1(n18771), .A2(n18598), .ZN(n18654) );
  NOR2_X1 U21671 ( .A1(n18639), .A2(n18654), .ZN(n18620) );
  OAI21_X1 U21672 ( .B1(n18876), .B2(n18572), .A(n18620), .ZN(n18573) );
  OAI211_X1 U21673 ( .C1(n19138), .C2(n18654), .A(n18573), .B(n18879), .ZN(
        n18595) );
  INV_X1 U21674 ( .A(n18595), .ZN(n18590) );
  NOR2_X1 U21675 ( .A1(n19042), .A2(n18620), .ZN(n18594) );
  AOI22_X1 U21676 ( .A1(n18960), .A2(n18849), .B1(n18908), .B2(n18594), .ZN(
        n18575) );
  AOI22_X1 U21677 ( .A1(n18909), .A2(n18612), .B1(n18913), .B2(n18654), .ZN(
        n18574) );
  OAI211_X1 U21678 ( .C1(n18590), .C2(n18576), .A(n18575), .B(n18574), .ZN(
        P3_U2884) );
  INV_X1 U21679 ( .A(n18922), .ZN(n18854) );
  AOI22_X1 U21680 ( .A1(n18960), .A2(n18854), .B1(n18917), .B2(n18594), .ZN(
        n18578) );
  AOI22_X1 U21681 ( .A1(n18612), .A2(n18918), .B1(n18919), .B2(n18654), .ZN(
        n18577) );
  OAI211_X1 U21682 ( .C1(n18590), .C2(n18579), .A(n18578), .B(n18577), .ZN(
        P3_U2885) );
  INV_X1 U21683 ( .A(n18887), .ZN(n18924) );
  AOI22_X1 U21684 ( .A1(n18612), .A2(n18924), .B1(n18923), .B2(n18594), .ZN(
        n18581) );
  AOI22_X1 U21685 ( .A1(n18960), .A2(n18884), .B1(n18925), .B2(n18654), .ZN(
        n18580) );
  OAI211_X1 U21686 ( .C1(n18590), .C2(n18582), .A(n18581), .B(n18580), .ZN(
        P3_U2886) );
  AOI22_X1 U21687 ( .A1(n18612), .A2(n18930), .B1(n18929), .B2(n18594), .ZN(
        n18584) );
  AOI22_X1 U21688 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18595), .B1(
        n18931), .B2(n18654), .ZN(n18583) );
  OAI211_X1 U21689 ( .C1(n18593), .C2(n18934), .A(n18584), .B(n18583), .ZN(
        P3_U2887) );
  AOI22_X1 U21690 ( .A1(n18612), .A2(n18805), .B1(n18935), .B2(n18594), .ZN(
        n18586) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18595), .B1(
        n18937), .B2(n18654), .ZN(n18585) );
  OAI211_X1 U21692 ( .C1(n18593), .C2(n18808), .A(n18586), .B(n18585), .ZN(
        P3_U2888) );
  AOI22_X1 U21693 ( .A1(n18612), .A2(n18942), .B1(n18941), .B2(n18594), .ZN(
        n18588) );
  AOI22_X1 U21694 ( .A1(n18960), .A2(n18836), .B1(n18944), .B2(n18654), .ZN(
        n18587) );
  OAI211_X1 U21695 ( .C1(n18590), .C2(n18589), .A(n18588), .B(n18587), .ZN(
        P3_U2889) );
  AOI22_X1 U21696 ( .A1(n18612), .A2(n18895), .B1(n18949), .B2(n18594), .ZN(
        n18592) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18595), .B1(
        n18951), .B2(n18654), .ZN(n18591) );
  OAI211_X1 U21698 ( .C1(n18593), .C2(n18898), .A(n18592), .B(n18591), .ZN(
        P3_U2890) );
  AOI22_X1 U21699 ( .A1(n18960), .A2(n18958), .B1(n18956), .B2(n18594), .ZN(
        n18597) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18595), .B1(
        n18959), .B2(n18654), .ZN(n18596) );
  OAI211_X1 U21701 ( .C1(n18619), .C2(n18964), .A(n18597), .B(n18596), .ZN(
        P3_U2891) );
  NOR2_X1 U21702 ( .A1(n19010), .A2(n18598), .ZN(n18644) );
  AND2_X1 U21703 ( .A1(n18795), .A2(n18644), .ZN(n18615) );
  AOI22_X1 U21704 ( .A1(n18909), .A2(n18639), .B1(n18908), .B2(n18615), .ZN(
        n18601) );
  NAND2_X1 U21705 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18644), .ZN(
        n18690) );
  INV_X1 U21706 ( .A(n18690), .ZN(n18681) );
  AOI21_X1 U21707 ( .B1(n19010), .B2(n18876), .A(n18667), .ZN(n18693) );
  OAI211_X1 U21708 ( .C1(n18681), .C2(n19138), .A(n18599), .B(n18693), .ZN(
        n18616) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18616), .B1(
        n18913), .B2(n18681), .ZN(n18600) );
  OAI211_X1 U21710 ( .C1(n18619), .C2(n18916), .A(n18601), .B(n18600), .ZN(
        P3_U2892) );
  AOI22_X1 U21711 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18616), .B1(
        n18917), .B2(n18615), .ZN(n18603) );
  AOI22_X1 U21712 ( .A1(n18919), .A2(n18681), .B1(n18918), .B2(n18635), .ZN(
        n18602) );
  OAI211_X1 U21713 ( .C1(n18619), .C2(n18922), .A(n18603), .B(n18602), .ZN(
        P3_U2893) );
  AOI22_X1 U21714 ( .A1(n18924), .A2(n18639), .B1(n18923), .B2(n18615), .ZN(
        n18605) );
  AOI22_X1 U21715 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18616), .B1(
        n18925), .B2(n18681), .ZN(n18604) );
  OAI211_X1 U21716 ( .C1(n18619), .C2(n18928), .A(n18605), .B(n18604), .ZN(
        P3_U2894) );
  INV_X1 U21717 ( .A(n18635), .ZN(n18626) );
  AOI22_X1 U21718 ( .A1(n18612), .A2(n18830), .B1(n18929), .B2(n18615), .ZN(
        n18607) );
  AOI22_X1 U21719 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18616), .B1(
        n18931), .B2(n18681), .ZN(n18606) );
  OAI211_X1 U21720 ( .C1(n18833), .C2(n18626), .A(n18607), .B(n18606), .ZN(
        P3_U2895) );
  AOI22_X1 U21721 ( .A1(n18805), .A2(n18635), .B1(n18935), .B2(n18615), .ZN(
        n18609) );
  AOI22_X1 U21722 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18616), .B1(
        n18937), .B2(n18681), .ZN(n18608) );
  OAI211_X1 U21723 ( .C1(n18619), .C2(n18808), .A(n18609), .B(n18608), .ZN(
        P3_U2896) );
  AOI22_X1 U21724 ( .A1(n18612), .A2(n18836), .B1(n18941), .B2(n18615), .ZN(
        n18611) );
  AOI22_X1 U21725 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18616), .B1(
        n18944), .B2(n18681), .ZN(n18610) );
  OAI211_X1 U21726 ( .C1(n18839), .C2(n18626), .A(n18611), .B(n18610), .ZN(
        P3_U2897) );
  AOI22_X1 U21727 ( .A1(n18612), .A2(n18950), .B1(n18949), .B2(n18615), .ZN(
        n18614) );
  AOI22_X1 U21728 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18616), .B1(
        n18951), .B2(n18681), .ZN(n18613) );
  OAI211_X1 U21729 ( .C1(n18954), .C2(n18626), .A(n18614), .B(n18613), .ZN(
        P3_U2898) );
  AOI22_X1 U21730 ( .A1(n18900), .A2(n18635), .B1(n18956), .B2(n18615), .ZN(
        n18618) );
  AOI22_X1 U21731 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18616), .B1(
        n18959), .B2(n18681), .ZN(n18617) );
  OAI211_X1 U21732 ( .C1(n18619), .C2(n18906), .A(n18618), .B(n18617), .ZN(
        P3_U2899) );
  INV_X1 U21733 ( .A(n18654), .ZN(n18665) );
  NAND2_X1 U21734 ( .A1(n18715), .A2(n18694), .ZN(n18714) );
  NOR2_X1 U21735 ( .A1(n18681), .A2(n18701), .ZN(n18669) );
  NOR2_X1 U21736 ( .A1(n19042), .A2(n18669), .ZN(n18638) );
  AOI22_X1 U21737 ( .A1(n18908), .A2(n18638), .B1(n18849), .B2(n18639), .ZN(
        n18623) );
  OAI22_X1 U21738 ( .A1(n18620), .A2(n18741), .B1(n18669), .B2(n18667), .ZN(
        n18621) );
  OAI21_X1 U21739 ( .B1(n18701), .B2(n19138), .A(n18621), .ZN(n18640) );
  AOI22_X1 U21740 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18640), .B1(
        n18913), .B2(n18701), .ZN(n18622) );
  OAI211_X1 U21741 ( .C1(n18853), .C2(n18665), .A(n18623), .B(n18622), .ZN(
        P3_U2900) );
  AOI22_X1 U21742 ( .A1(n18918), .A2(n18654), .B1(n18917), .B2(n18638), .ZN(
        n18625) );
  AOI22_X1 U21743 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18640), .B1(
        n18919), .B2(n18701), .ZN(n18624) );
  OAI211_X1 U21744 ( .C1(n18922), .C2(n18626), .A(n18625), .B(n18624), .ZN(
        P3_U2901) );
  AOI22_X1 U21745 ( .A1(n18884), .A2(n18639), .B1(n18923), .B2(n18638), .ZN(
        n18628) );
  AOI22_X1 U21746 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18640), .B1(
        n18925), .B2(n18701), .ZN(n18627) );
  OAI211_X1 U21747 ( .C1(n18887), .C2(n18665), .A(n18628), .B(n18627), .ZN(
        P3_U2902) );
  AOI22_X1 U21748 ( .A1(n18929), .A2(n18638), .B1(n18830), .B2(n18639), .ZN(
        n18630) );
  AOI22_X1 U21749 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18640), .B1(
        n18931), .B2(n18701), .ZN(n18629) );
  OAI211_X1 U21750 ( .C1(n18833), .C2(n18665), .A(n18630), .B(n18629), .ZN(
        P3_U2903) );
  AOI22_X1 U21751 ( .A1(n18936), .A2(n18639), .B1(n18935), .B2(n18638), .ZN(
        n18632) );
  AOI22_X1 U21752 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18640), .B1(
        n18937), .B2(n18701), .ZN(n18631) );
  OAI211_X1 U21753 ( .C1(n18940), .C2(n18665), .A(n18632), .B(n18631), .ZN(
        P3_U2904) );
  AOI22_X1 U21754 ( .A1(n18836), .A2(n18635), .B1(n18941), .B2(n18638), .ZN(
        n18634) );
  AOI22_X1 U21755 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18640), .B1(
        n18944), .B2(n18701), .ZN(n18633) );
  OAI211_X1 U21756 ( .C1(n18839), .C2(n18665), .A(n18634), .B(n18633), .ZN(
        P3_U2905) );
  AOI22_X1 U21757 ( .A1(n18950), .A2(n18635), .B1(n18949), .B2(n18638), .ZN(
        n18637) );
  AOI22_X1 U21758 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18640), .B1(
        n18951), .B2(n18701), .ZN(n18636) );
  OAI211_X1 U21759 ( .C1(n18954), .C2(n18665), .A(n18637), .B(n18636), .ZN(
        P3_U2906) );
  AOI22_X1 U21760 ( .A1(n18958), .A2(n18639), .B1(n18956), .B2(n18638), .ZN(
        n18642) );
  AOI22_X1 U21761 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18640), .B1(
        n18959), .B2(n18701), .ZN(n18641) );
  OAI211_X1 U21762 ( .C1(n18964), .C2(n18665), .A(n18642), .B(n18641), .ZN(
        P3_U2907) );
  NOR2_X1 U21763 ( .A1(n18645), .A2(n18742), .ZN(n18661) );
  AOI22_X1 U21764 ( .A1(n18909), .A2(n18681), .B1(n18908), .B2(n18661), .ZN(
        n18647) );
  AOI22_X1 U21765 ( .A1(n18545), .A2(n18644), .B1(n18694), .B2(n18643), .ZN(
        n18662) );
  NOR2_X2 U21766 ( .A1(n18645), .A2(n18743), .ZN(n18734) );
  AOI22_X1 U21767 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18662), .B1(
        n18913), .B2(n18734), .ZN(n18646) );
  OAI211_X1 U21768 ( .C1(n18916), .C2(n18665), .A(n18647), .B(n18646), .ZN(
        P3_U2908) );
  AOI22_X1 U21769 ( .A1(n18854), .A2(n18654), .B1(n18917), .B2(n18661), .ZN(
        n18649) );
  AOI22_X1 U21770 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18662), .B1(
        n18919), .B2(n18734), .ZN(n18648) );
  OAI211_X1 U21771 ( .C1(n18857), .C2(n18690), .A(n18649), .B(n18648), .ZN(
        P3_U2909) );
  AOI22_X1 U21772 ( .A1(n18924), .A2(n18681), .B1(n18923), .B2(n18661), .ZN(
        n18651) );
  AOI22_X1 U21773 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18662), .B1(
        n18925), .B2(n18734), .ZN(n18650) );
  OAI211_X1 U21774 ( .C1(n18928), .C2(n18665), .A(n18651), .B(n18650), .ZN(
        P3_U2910) );
  AOI22_X1 U21775 ( .A1(n18929), .A2(n18661), .B1(n18830), .B2(n18654), .ZN(
        n18653) );
  AOI22_X1 U21776 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18662), .B1(
        n18931), .B2(n18734), .ZN(n18652) );
  OAI211_X1 U21777 ( .C1(n18833), .C2(n18690), .A(n18653), .B(n18652), .ZN(
        P3_U2911) );
  AOI22_X1 U21778 ( .A1(n18936), .A2(n18654), .B1(n18935), .B2(n18661), .ZN(
        n18656) );
  AOI22_X1 U21779 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18662), .B1(
        n18937), .B2(n18734), .ZN(n18655) );
  OAI211_X1 U21780 ( .C1(n18940), .C2(n18690), .A(n18656), .B(n18655), .ZN(
        P3_U2912) );
  AOI22_X1 U21781 ( .A1(n18942), .A2(n18681), .B1(n18941), .B2(n18661), .ZN(
        n18658) );
  AOI22_X1 U21782 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18662), .B1(
        n18944), .B2(n18734), .ZN(n18657) );
  OAI211_X1 U21783 ( .C1(n18948), .C2(n18665), .A(n18658), .B(n18657), .ZN(
        P3_U2913) );
  AOI22_X1 U21784 ( .A1(n18949), .A2(n18661), .B1(n18895), .B2(n18681), .ZN(
        n18660) );
  AOI22_X1 U21785 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18662), .B1(
        n18951), .B2(n18734), .ZN(n18659) );
  OAI211_X1 U21786 ( .C1(n18898), .C2(n18665), .A(n18660), .B(n18659), .ZN(
        P3_U2914) );
  AOI22_X1 U21787 ( .A1(n18900), .A2(n18681), .B1(n18956), .B2(n18661), .ZN(
        n18664) );
  AOI22_X1 U21788 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18662), .B1(
        n18959), .B2(n18734), .ZN(n18663) );
  OAI211_X1 U21789 ( .C1(n18906), .C2(n18665), .A(n18664), .B(n18663), .ZN(
        P3_U2915) );
  INV_X1 U21790 ( .A(n18734), .ZN(n18729) );
  INV_X1 U21791 ( .A(n18771), .ZN(n18666) );
  NAND2_X1 U21792 ( .A1(n18694), .A2(n18666), .ZN(n18737) );
  NAND2_X1 U21793 ( .A1(n18729), .A2(n18737), .ZN(n18716) );
  INV_X1 U21794 ( .A(n18716), .ZN(n18668) );
  NOR2_X1 U21795 ( .A1(n19042), .A2(n18668), .ZN(n18686) );
  AOI22_X1 U21796 ( .A1(n18909), .A2(n18701), .B1(n18908), .B2(n18686), .ZN(
        n18672) );
  OAI22_X1 U21797 ( .A1(n18669), .A2(n18741), .B1(n18668), .B2(n18667), .ZN(
        n18670) );
  OAI21_X1 U21798 ( .B1(n18766), .B2(n19138), .A(n18670), .ZN(n18687) );
  AOI22_X1 U21799 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18687), .B1(
        n18913), .B2(n18766), .ZN(n18671) );
  OAI211_X1 U21800 ( .C1(n18916), .C2(n18690), .A(n18672), .B(n18671), .ZN(
        P3_U2916) );
  AOI22_X1 U21801 ( .A1(n18918), .A2(n18701), .B1(n18917), .B2(n18686), .ZN(
        n18674) );
  AOI22_X1 U21802 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18687), .B1(
        n18919), .B2(n18766), .ZN(n18673) );
  OAI211_X1 U21803 ( .C1(n18922), .C2(n18690), .A(n18674), .B(n18673), .ZN(
        P3_U2917) );
  AOI22_X1 U21804 ( .A1(n18924), .A2(n18701), .B1(n18923), .B2(n18686), .ZN(
        n18676) );
  AOI22_X1 U21805 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18687), .B1(
        n18925), .B2(n18766), .ZN(n18675) );
  OAI211_X1 U21806 ( .C1(n18928), .C2(n18690), .A(n18676), .B(n18675), .ZN(
        P3_U2918) );
  AOI22_X1 U21807 ( .A1(n18929), .A2(n18686), .B1(n18830), .B2(n18681), .ZN(
        n18678) );
  AOI22_X1 U21808 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18687), .B1(
        n18931), .B2(n18766), .ZN(n18677) );
  OAI211_X1 U21809 ( .C1(n18833), .C2(n18714), .A(n18678), .B(n18677), .ZN(
        P3_U2919) );
  AOI22_X1 U21810 ( .A1(n18936), .A2(n18681), .B1(n18935), .B2(n18686), .ZN(
        n18680) );
  AOI22_X1 U21811 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18687), .B1(
        n18937), .B2(n18766), .ZN(n18679) );
  OAI211_X1 U21812 ( .C1(n18940), .C2(n18714), .A(n18680), .B(n18679), .ZN(
        P3_U2920) );
  AOI22_X1 U21813 ( .A1(n18836), .A2(n18681), .B1(n18941), .B2(n18686), .ZN(
        n18683) );
  AOI22_X1 U21814 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18687), .B1(
        n18944), .B2(n18766), .ZN(n18682) );
  OAI211_X1 U21815 ( .C1(n18839), .C2(n18714), .A(n18683), .B(n18682), .ZN(
        P3_U2921) );
  AOI22_X1 U21816 ( .A1(n18949), .A2(n18686), .B1(n18895), .B2(n18701), .ZN(
        n18685) );
  AOI22_X1 U21817 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18687), .B1(
        n18951), .B2(n18766), .ZN(n18684) );
  OAI211_X1 U21818 ( .C1(n18898), .C2(n18690), .A(n18685), .B(n18684), .ZN(
        P3_U2922) );
  AOI22_X1 U21819 ( .A1(n18900), .A2(n18701), .B1(n18956), .B2(n18686), .ZN(
        n18689) );
  AOI22_X1 U21820 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18687), .B1(
        n18959), .B2(n18766), .ZN(n18688) );
  OAI211_X1 U21821 ( .C1(n18906), .C2(n18690), .A(n18689), .B(n18688), .ZN(
        P3_U2923) );
  NAND2_X1 U21822 ( .A1(n18691), .A2(n19018), .ZN(n18740) );
  NOR2_X1 U21823 ( .A1(n19042), .A2(n18740), .ZN(n18710) );
  AOI22_X1 U21824 ( .A1(n18909), .A2(n18734), .B1(n18908), .B2(n18710), .ZN(
        n18696) );
  NAND3_X1 U21825 ( .A1(n18694), .A2(n18693), .A3(n18692), .ZN(n18711) );
  NOR2_X2 U21826 ( .A1(n19008), .A2(n18740), .ZN(n18787) );
  AOI22_X1 U21827 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18711), .B1(
        n18913), .B2(n18787), .ZN(n18695) );
  OAI211_X1 U21828 ( .C1(n18916), .C2(n18714), .A(n18696), .B(n18695), .ZN(
        P3_U2924) );
  AOI22_X1 U21829 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18711), .B1(
        n18917), .B2(n18710), .ZN(n18698) );
  AOI22_X1 U21830 ( .A1(n18919), .A2(n18787), .B1(n18918), .B2(n18734), .ZN(
        n18697) );
  OAI211_X1 U21831 ( .C1(n18922), .C2(n18714), .A(n18698), .B(n18697), .ZN(
        P3_U2925) );
  AOI22_X1 U21832 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18711), .B1(
        n18923), .B2(n18710), .ZN(n18700) );
  AOI22_X1 U21833 ( .A1(n18924), .A2(n18734), .B1(n18925), .B2(n18787), .ZN(
        n18699) );
  OAI211_X1 U21834 ( .C1(n18928), .C2(n18714), .A(n18700), .B(n18699), .ZN(
        P3_U2926) );
  AOI22_X1 U21835 ( .A1(n18929), .A2(n18710), .B1(n18830), .B2(n18701), .ZN(
        n18703) );
  AOI22_X1 U21836 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18711), .B1(
        n18931), .B2(n18787), .ZN(n18702) );
  OAI211_X1 U21837 ( .C1(n18833), .C2(n18729), .A(n18703), .B(n18702), .ZN(
        P3_U2927) );
  AOI22_X1 U21838 ( .A1(n18805), .A2(n18734), .B1(n18935), .B2(n18710), .ZN(
        n18705) );
  AOI22_X1 U21839 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18711), .B1(
        n18937), .B2(n18787), .ZN(n18704) );
  OAI211_X1 U21840 ( .C1(n18808), .C2(n18714), .A(n18705), .B(n18704), .ZN(
        P3_U2928) );
  AOI22_X1 U21841 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18711), .B1(
        n18941), .B2(n18710), .ZN(n18707) );
  AOI22_X1 U21842 ( .A1(n18944), .A2(n18787), .B1(n18942), .B2(n18734), .ZN(
        n18706) );
  OAI211_X1 U21843 ( .C1(n18948), .C2(n18714), .A(n18707), .B(n18706), .ZN(
        P3_U2929) );
  AOI22_X1 U21844 ( .A1(n18949), .A2(n18710), .B1(n18895), .B2(n18734), .ZN(
        n18709) );
  AOI22_X1 U21845 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18711), .B1(
        n18951), .B2(n18787), .ZN(n18708) );
  OAI211_X1 U21846 ( .C1(n18898), .C2(n18714), .A(n18709), .B(n18708), .ZN(
        P3_U2930) );
  AOI22_X1 U21847 ( .A1(n18900), .A2(n18734), .B1(n18956), .B2(n18710), .ZN(
        n18713) );
  AOI22_X1 U21848 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18711), .B1(
        n18959), .B2(n18787), .ZN(n18712) );
  OAI211_X1 U21849 ( .C1(n18906), .C2(n18714), .A(n18713), .B(n18712), .ZN(
        P3_U2931) );
  INV_X1 U21850 ( .A(n18787), .ZN(n18794) );
  INV_X1 U21851 ( .A(n18715), .ZN(n19011) );
  NOR2_X2 U21852 ( .A1(n19011), .A2(n18819), .ZN(n18815) );
  INV_X1 U21853 ( .A(n18815), .ZN(n18811) );
  NAND2_X1 U21854 ( .A1(n18794), .A2(n18811), .ZN(n18772) );
  OAI221_X1 U21855 ( .B1(n18772), .B2(n18773), .C1(n18772), .C2(n18716), .A(
        n18821), .ZN(n18733) );
  AND2_X1 U21856 ( .A1(n18795), .A2(n18772), .ZN(n18732) );
  AOI22_X1 U21857 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18733), .B1(
        n18908), .B2(n18732), .ZN(n18718) );
  AOI22_X1 U21858 ( .A1(n18909), .A2(n18766), .B1(n18913), .B2(n18815), .ZN(
        n18717) );
  OAI211_X1 U21859 ( .C1(n18916), .C2(n18729), .A(n18718), .B(n18717), .ZN(
        P3_U2932) );
  AOI22_X1 U21860 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18733), .B1(
        n18917), .B2(n18732), .ZN(n18720) );
  AOI22_X1 U21861 ( .A1(n18919), .A2(n18815), .B1(n18918), .B2(n18766), .ZN(
        n18719) );
  OAI211_X1 U21862 ( .C1(n18922), .C2(n18729), .A(n18720), .B(n18719), .ZN(
        P3_U2933) );
  AOI22_X1 U21863 ( .A1(n18924), .A2(n18766), .B1(n18923), .B2(n18732), .ZN(
        n18722) );
  AOI22_X1 U21864 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18733), .B1(
        n18925), .B2(n18815), .ZN(n18721) );
  OAI211_X1 U21865 ( .C1(n18928), .C2(n18729), .A(n18722), .B(n18721), .ZN(
        P3_U2934) );
  AOI22_X1 U21866 ( .A1(n18930), .A2(n18766), .B1(n18929), .B2(n18732), .ZN(
        n18724) );
  AOI22_X1 U21867 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18733), .B1(
        n18931), .B2(n18815), .ZN(n18723) );
  OAI211_X1 U21868 ( .C1(n18934), .C2(n18729), .A(n18724), .B(n18723), .ZN(
        P3_U2935) );
  AOI22_X1 U21869 ( .A1(n18805), .A2(n18766), .B1(n18935), .B2(n18732), .ZN(
        n18726) );
  AOI22_X1 U21870 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18733), .B1(
        n18937), .B2(n18815), .ZN(n18725) );
  OAI211_X1 U21871 ( .C1(n18808), .C2(n18729), .A(n18726), .B(n18725), .ZN(
        P3_U2936) );
  AOI22_X1 U21872 ( .A1(n18942), .A2(n18766), .B1(n18941), .B2(n18732), .ZN(
        n18728) );
  AOI22_X1 U21873 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18733), .B1(
        n18944), .B2(n18815), .ZN(n18727) );
  OAI211_X1 U21874 ( .C1(n18948), .C2(n18729), .A(n18728), .B(n18727), .ZN(
        P3_U2937) );
  AOI22_X1 U21875 ( .A1(n18950), .A2(n18734), .B1(n18949), .B2(n18732), .ZN(
        n18731) );
  AOI22_X1 U21876 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18733), .B1(
        n18951), .B2(n18815), .ZN(n18730) );
  OAI211_X1 U21877 ( .C1(n18954), .C2(n18737), .A(n18731), .B(n18730), .ZN(
        P3_U2938) );
  AOI22_X1 U21878 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18733), .B1(
        n18956), .B2(n18732), .ZN(n18736) );
  AOI22_X1 U21879 ( .A1(n18959), .A2(n18815), .B1(n18958), .B2(n18734), .ZN(
        n18735) );
  OAI211_X1 U21880 ( .C1(n18964), .C2(n18737), .A(n18736), .B(n18735), .ZN(
        P3_U2939) );
  NAND2_X1 U21881 ( .A1(n18796), .A2(n19010), .ZN(n18738) );
  OAI22_X1 U21882 ( .A1(n18741), .A2(n18740), .B1(n18739), .B2(n18738), .ZN(
        n18769) );
  NOR2_X1 U21883 ( .A1(n18819), .A2(n18742), .ZN(n18765) );
  AOI22_X1 U21884 ( .A1(n18909), .A2(n18787), .B1(n18908), .B2(n18765), .ZN(
        n18745) );
  NOR2_X2 U21885 ( .A1(n18819), .A2(n18743), .ZN(n18845) );
  AOI22_X1 U21886 ( .A1(n18913), .A2(n18845), .B1(n18849), .B2(n18766), .ZN(
        n18744) );
  OAI211_X1 U21887 ( .C1(n18746), .C2(n18769), .A(n18745), .B(n18744), .ZN(
        P3_U2940) );
  AOI22_X1 U21888 ( .A1(n18854), .A2(n18766), .B1(n18917), .B2(n18765), .ZN(
        n18748) );
  AOI22_X1 U21889 ( .A1(n18919), .A2(n18845), .B1(n18918), .B2(n18787), .ZN(
        n18747) );
  OAI211_X1 U21890 ( .C1(n18749), .C2(n18769), .A(n18748), .B(n18747), .ZN(
        P3_U2941) );
  AOI22_X1 U21891 ( .A1(n18884), .A2(n18766), .B1(n18923), .B2(n18765), .ZN(
        n18751) );
  AOI22_X1 U21892 ( .A1(n18924), .A2(n18787), .B1(n18925), .B2(n18845), .ZN(
        n18750) );
  OAI211_X1 U21893 ( .C1(n18752), .C2(n18769), .A(n18751), .B(n18750), .ZN(
        P3_U2942) );
  AOI22_X1 U21894 ( .A1(n18930), .A2(n18787), .B1(n18929), .B2(n18765), .ZN(
        n18754) );
  AOI22_X1 U21895 ( .A1(n18931), .A2(n18845), .B1(n18830), .B2(n18766), .ZN(
        n18753) );
  OAI211_X1 U21896 ( .C1(n18755), .C2(n18769), .A(n18754), .B(n18753), .ZN(
        P3_U2943) );
  AOI22_X1 U21897 ( .A1(n18936), .A2(n18766), .B1(n18935), .B2(n18765), .ZN(
        n18757) );
  AOI22_X1 U21898 ( .A1(n18805), .A2(n18787), .B1(n18937), .B2(n18845), .ZN(
        n18756) );
  OAI211_X1 U21899 ( .C1(n18758), .C2(n18769), .A(n18757), .B(n18756), .ZN(
        P3_U2944) );
  AOI22_X1 U21900 ( .A1(n18942), .A2(n18787), .B1(n18941), .B2(n18765), .ZN(
        n18760) );
  AOI22_X1 U21901 ( .A1(n18836), .A2(n18766), .B1(n18944), .B2(n18845), .ZN(
        n18759) );
  OAI211_X1 U21902 ( .C1(n18761), .C2(n18769), .A(n18760), .B(n18759), .ZN(
        P3_U2945) );
  AOI22_X1 U21903 ( .A1(n18950), .A2(n18766), .B1(n18949), .B2(n18765), .ZN(
        n18763) );
  AOI22_X1 U21904 ( .A1(n18951), .A2(n18845), .B1(n18895), .B2(n18787), .ZN(
        n18762) );
  OAI211_X1 U21905 ( .C1(n18764), .C2(n18769), .A(n18763), .B(n18762), .ZN(
        P3_U2946) );
  AOI22_X1 U21906 ( .A1(n18958), .A2(n18766), .B1(n18956), .B2(n18765), .ZN(
        n18768) );
  AOI22_X1 U21907 ( .A1(n18900), .A2(n18787), .B1(n18959), .B2(n18845), .ZN(
        n18767) );
  OAI211_X1 U21908 ( .C1(n18770), .C2(n18769), .A(n18768), .B(n18767), .ZN(
        P3_U2947) );
  INV_X1 U21909 ( .A(n18845), .ZN(n18842) );
  NOR2_X2 U21910 ( .A1(n18819), .A2(n18771), .ZN(n18870) );
  INV_X1 U21911 ( .A(n18870), .ZN(n18868) );
  AOI21_X1 U21912 ( .B1(n18842), .B2(n18868), .A(n19042), .ZN(n18790) );
  AOI22_X1 U21913 ( .A1(n18909), .A2(n18815), .B1(n18908), .B2(n18790), .ZN(
        n18776) );
  NAND2_X1 U21914 ( .A1(n18842), .A2(n18868), .ZN(n18774) );
  OAI221_X1 U21915 ( .B1(n18774), .B2(n18773), .C1(n18774), .C2(n18772), .A(
        n18821), .ZN(n18791) );
  AOI22_X1 U21916 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18791), .B1(
        n18913), .B2(n18870), .ZN(n18775) );
  OAI211_X1 U21917 ( .C1(n18916), .C2(n18794), .A(n18776), .B(n18775), .ZN(
        P3_U2948) );
  AOI22_X1 U21918 ( .A1(n18918), .A2(n18815), .B1(n18917), .B2(n18790), .ZN(
        n18778) );
  AOI22_X1 U21919 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18791), .B1(
        n18919), .B2(n18870), .ZN(n18777) );
  OAI211_X1 U21920 ( .C1(n18922), .C2(n18794), .A(n18778), .B(n18777), .ZN(
        P3_U2949) );
  AOI22_X1 U21921 ( .A1(n18924), .A2(n18815), .B1(n18923), .B2(n18790), .ZN(
        n18780) );
  AOI22_X1 U21922 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18791), .B1(
        n18925), .B2(n18870), .ZN(n18779) );
  OAI211_X1 U21923 ( .C1(n18928), .C2(n18794), .A(n18780), .B(n18779), .ZN(
        P3_U2950) );
  AOI22_X1 U21924 ( .A1(n18930), .A2(n18815), .B1(n18929), .B2(n18790), .ZN(
        n18782) );
  AOI22_X1 U21925 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18791), .B1(
        n18931), .B2(n18870), .ZN(n18781) );
  OAI211_X1 U21926 ( .C1(n18934), .C2(n18794), .A(n18782), .B(n18781), .ZN(
        P3_U2951) );
  AOI22_X1 U21927 ( .A1(n18936), .A2(n18787), .B1(n18935), .B2(n18790), .ZN(
        n18784) );
  AOI22_X1 U21928 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18791), .B1(
        n18937), .B2(n18870), .ZN(n18783) );
  OAI211_X1 U21929 ( .C1(n18940), .C2(n18811), .A(n18784), .B(n18783), .ZN(
        P3_U2952) );
  AOI22_X1 U21930 ( .A1(n18836), .A2(n18787), .B1(n18941), .B2(n18790), .ZN(
        n18786) );
  AOI22_X1 U21931 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18791), .B1(
        n18944), .B2(n18870), .ZN(n18785) );
  OAI211_X1 U21932 ( .C1(n18839), .C2(n18811), .A(n18786), .B(n18785), .ZN(
        P3_U2953) );
  AOI22_X1 U21933 ( .A1(n18950), .A2(n18787), .B1(n18949), .B2(n18790), .ZN(
        n18789) );
  AOI22_X1 U21934 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18791), .B1(
        n18951), .B2(n18870), .ZN(n18788) );
  OAI211_X1 U21935 ( .C1(n18954), .C2(n18811), .A(n18789), .B(n18788), .ZN(
        P3_U2954) );
  AOI22_X1 U21936 ( .A1(n18900), .A2(n18815), .B1(n18956), .B2(n18790), .ZN(
        n18793) );
  AOI22_X1 U21937 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18791), .B1(
        n18959), .B2(n18870), .ZN(n18792) );
  OAI211_X1 U21938 ( .C1(n18906), .C2(n18794), .A(n18793), .B(n18792), .ZN(
        P3_U2955) );
  NOR2_X1 U21939 ( .A1(n19010), .A2(n18819), .ZN(n18850) );
  AND2_X1 U21940 ( .A1(n18795), .A2(n18850), .ZN(n18814) );
  AOI22_X1 U21941 ( .A1(n18909), .A2(n18845), .B1(n18908), .B2(n18814), .ZN(
        n18798) );
  OAI211_X1 U21942 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18545), .A(
        n18910), .B(n18796), .ZN(n18816) );
  NAND2_X1 U21943 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18850), .ZN(
        n18905) );
  AOI22_X1 U21944 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18816), .B1(
        n18913), .B2(n18890), .ZN(n18797) );
  OAI211_X1 U21945 ( .C1(n18916), .C2(n18811), .A(n18798), .B(n18797), .ZN(
        P3_U2956) );
  AOI22_X1 U21946 ( .A1(n18918), .A2(n18845), .B1(n18917), .B2(n18814), .ZN(
        n18800) );
  AOI22_X1 U21947 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18816), .B1(
        n18919), .B2(n18890), .ZN(n18799) );
  OAI211_X1 U21948 ( .C1(n18922), .C2(n18811), .A(n18800), .B(n18799), .ZN(
        P3_U2957) );
  AOI22_X1 U21949 ( .A1(n18884), .A2(n18815), .B1(n18923), .B2(n18814), .ZN(
        n18802) );
  AOI22_X1 U21950 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18816), .B1(
        n18925), .B2(n18890), .ZN(n18801) );
  OAI211_X1 U21951 ( .C1(n18887), .C2(n18842), .A(n18802), .B(n18801), .ZN(
        P3_U2958) );
  AOI22_X1 U21952 ( .A1(n18929), .A2(n18814), .B1(n18830), .B2(n18815), .ZN(
        n18804) );
  AOI22_X1 U21953 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18816), .B1(
        n18931), .B2(n18890), .ZN(n18803) );
  OAI211_X1 U21954 ( .C1(n18833), .C2(n18842), .A(n18804), .B(n18803), .ZN(
        P3_U2959) );
  AOI22_X1 U21955 ( .A1(n18805), .A2(n18845), .B1(n18935), .B2(n18814), .ZN(
        n18807) );
  AOI22_X1 U21956 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18816), .B1(
        n18937), .B2(n18890), .ZN(n18806) );
  OAI211_X1 U21957 ( .C1(n18808), .C2(n18811), .A(n18807), .B(n18806), .ZN(
        P3_U2960) );
  AOI22_X1 U21958 ( .A1(n18942), .A2(n18845), .B1(n18941), .B2(n18814), .ZN(
        n18810) );
  AOI22_X1 U21959 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18816), .B1(
        n18944), .B2(n18890), .ZN(n18809) );
  OAI211_X1 U21960 ( .C1(n18948), .C2(n18811), .A(n18810), .B(n18809), .ZN(
        P3_U2961) );
  AOI22_X1 U21961 ( .A1(n18950), .A2(n18815), .B1(n18949), .B2(n18814), .ZN(
        n18813) );
  AOI22_X1 U21962 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18816), .B1(
        n18951), .B2(n18890), .ZN(n18812) );
  OAI211_X1 U21963 ( .C1(n18954), .C2(n18842), .A(n18813), .B(n18812), .ZN(
        P3_U2962) );
  AOI22_X1 U21964 ( .A1(n18958), .A2(n18815), .B1(n18956), .B2(n18814), .ZN(
        n18818) );
  AOI22_X1 U21965 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18816), .B1(
        n18959), .B2(n18890), .ZN(n18817) );
  OAI211_X1 U21966 ( .C1(n18964), .C2(n18842), .A(n18818), .B(n18817), .ZN(
        P3_U2963) );
  NOR3_X1 U21967 ( .A1(n18820), .A2(n18819), .A3(n18876), .ZN(n18823) );
  INV_X1 U21968 ( .A(n18912), .ZN(n18848) );
  NOR2_X2 U21969 ( .A1(n18848), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18957) );
  NOR2_X1 U21970 ( .A1(n18890), .A2(n18957), .ZN(n18877) );
  INV_X1 U21971 ( .A(n18877), .ZN(n18822) );
  OAI21_X1 U21972 ( .B1(n18823), .B2(n18822), .A(n18821), .ZN(n18844) );
  NOR2_X1 U21973 ( .A1(n19042), .A2(n18877), .ZN(n18843) );
  AOI22_X1 U21974 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18844), .B1(
        n18908), .B2(n18843), .ZN(n18825) );
  AOI22_X1 U21975 ( .A1(n18909), .A2(n18870), .B1(n18913), .B2(n18957), .ZN(
        n18824) );
  OAI211_X1 U21976 ( .C1(n18916), .C2(n18842), .A(n18825), .B(n18824), .ZN(
        P3_U2964) );
  AOI22_X1 U21977 ( .A1(n18918), .A2(n18870), .B1(n18917), .B2(n18843), .ZN(
        n18827) );
  AOI22_X1 U21978 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18844), .B1(
        n18919), .B2(n18957), .ZN(n18826) );
  OAI211_X1 U21979 ( .C1(n18922), .C2(n18842), .A(n18827), .B(n18826), .ZN(
        P3_U2965) );
  AOI22_X1 U21980 ( .A1(n18924), .A2(n18870), .B1(n18923), .B2(n18843), .ZN(
        n18829) );
  AOI22_X1 U21981 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18844), .B1(
        n18925), .B2(n18957), .ZN(n18828) );
  OAI211_X1 U21982 ( .C1(n18928), .C2(n18842), .A(n18829), .B(n18828), .ZN(
        P3_U2966) );
  AOI22_X1 U21983 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18844), .B1(
        n18929), .B2(n18843), .ZN(n18832) );
  AOI22_X1 U21984 ( .A1(n18931), .A2(n18957), .B1(n18830), .B2(n18845), .ZN(
        n18831) );
  OAI211_X1 U21985 ( .C1(n18833), .C2(n18868), .A(n18832), .B(n18831), .ZN(
        P3_U2967) );
  AOI22_X1 U21986 ( .A1(n18936), .A2(n18845), .B1(n18935), .B2(n18843), .ZN(
        n18835) );
  AOI22_X1 U21987 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18844), .B1(
        n18937), .B2(n18957), .ZN(n18834) );
  OAI211_X1 U21988 ( .C1(n18940), .C2(n18868), .A(n18835), .B(n18834), .ZN(
        P3_U2968) );
  AOI22_X1 U21989 ( .A1(n18836), .A2(n18845), .B1(n18941), .B2(n18843), .ZN(
        n18838) );
  AOI22_X1 U21990 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18844), .B1(
        n18944), .B2(n18957), .ZN(n18837) );
  OAI211_X1 U21991 ( .C1(n18839), .C2(n18868), .A(n18838), .B(n18837), .ZN(
        P3_U2969) );
  AOI22_X1 U21992 ( .A1(n18949), .A2(n18843), .B1(n18895), .B2(n18870), .ZN(
        n18841) );
  AOI22_X1 U21993 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18844), .B1(
        n18951), .B2(n18957), .ZN(n18840) );
  OAI211_X1 U21994 ( .C1(n18898), .C2(n18842), .A(n18841), .B(n18840), .ZN(
        P3_U2970) );
  AOI22_X1 U21995 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18844), .B1(
        n18956), .B2(n18843), .ZN(n18847) );
  AOI22_X1 U21996 ( .A1(n18959), .A2(n18957), .B1(n18958), .B2(n18845), .ZN(
        n18846) );
  OAI211_X1 U21997 ( .C1(n18964), .C2(n18868), .A(n18847), .B(n18846), .ZN(
        P3_U2971) );
  NOR2_X1 U21998 ( .A1(n19042), .A2(n18848), .ZN(n18869) );
  AOI22_X1 U21999 ( .A1(n18908), .A2(n18869), .B1(n18849), .B2(n18870), .ZN(
        n18852) );
  AOI22_X1 U22000 ( .A1(n18545), .A2(n18850), .B1(n18912), .B2(n18910), .ZN(
        n18871) );
  AOI22_X1 U22001 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18871), .B1(
        n18913), .B2(n18943), .ZN(n18851) );
  OAI211_X1 U22002 ( .C1(n18853), .C2(n18905), .A(n18852), .B(n18851), .ZN(
        P3_U2972) );
  AOI22_X1 U22003 ( .A1(n18854), .A2(n18870), .B1(n18917), .B2(n18869), .ZN(
        n18856) );
  AOI22_X1 U22004 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18871), .B1(
        n18943), .B2(n18919), .ZN(n18855) );
  OAI211_X1 U22005 ( .C1(n18857), .C2(n18905), .A(n18856), .B(n18855), .ZN(
        P3_U2973) );
  AOI22_X1 U22006 ( .A1(n18884), .A2(n18870), .B1(n18923), .B2(n18869), .ZN(
        n18859) );
  AOI22_X1 U22007 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18871), .B1(
        n18943), .B2(n18925), .ZN(n18858) );
  OAI211_X1 U22008 ( .C1(n18887), .C2(n18905), .A(n18859), .B(n18858), .ZN(
        P3_U2974) );
  AOI22_X1 U22009 ( .A1(n18930), .A2(n18890), .B1(n18929), .B2(n18869), .ZN(
        n18861) );
  AOI22_X1 U22010 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18871), .B1(
        n18943), .B2(n18931), .ZN(n18860) );
  OAI211_X1 U22011 ( .C1(n18934), .C2(n18868), .A(n18861), .B(n18860), .ZN(
        P3_U2975) );
  AOI22_X1 U22012 ( .A1(n18936), .A2(n18870), .B1(n18935), .B2(n18869), .ZN(
        n18863) );
  AOI22_X1 U22013 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18871), .B1(
        n18943), .B2(n18937), .ZN(n18862) );
  OAI211_X1 U22014 ( .C1(n18940), .C2(n18905), .A(n18863), .B(n18862), .ZN(
        P3_U2976) );
  AOI22_X1 U22015 ( .A1(n18942), .A2(n18890), .B1(n18941), .B2(n18869), .ZN(
        n18865) );
  AOI22_X1 U22016 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18871), .B1(
        n18943), .B2(n18944), .ZN(n18864) );
  OAI211_X1 U22017 ( .C1(n18948), .C2(n18868), .A(n18865), .B(n18864), .ZN(
        P3_U2977) );
  AOI22_X1 U22018 ( .A1(n18949), .A2(n18869), .B1(n18895), .B2(n18890), .ZN(
        n18867) );
  AOI22_X1 U22019 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18871), .B1(
        n18943), .B2(n18951), .ZN(n18866) );
  OAI211_X1 U22020 ( .C1(n18898), .C2(n18868), .A(n18867), .B(n18866), .ZN(
        P3_U2978) );
  AOI22_X1 U22021 ( .A1(n18958), .A2(n18870), .B1(n18956), .B2(n18869), .ZN(
        n18873) );
  AOI22_X1 U22022 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18871), .B1(
        n18943), .B2(n18959), .ZN(n18872) );
  OAI211_X1 U22023 ( .C1(n18964), .C2(n18905), .A(n18873), .B(n18872), .ZN(
        P3_U2979) );
  INV_X1 U22024 ( .A(n18874), .ZN(n18875) );
  NOR2_X1 U22025 ( .A1(n19042), .A2(n18875), .ZN(n18899) );
  AOI22_X1 U22026 ( .A1(n18909), .A2(n18957), .B1(n18908), .B2(n18899), .ZN(
        n18881) );
  OAI21_X1 U22027 ( .B1(n18877), .B2(n18876), .A(n18875), .ZN(n18878) );
  OAI211_X1 U22028 ( .C1(n18901), .C2(n19138), .A(n18879), .B(n18878), .ZN(
        n18902) );
  AOI22_X1 U22029 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18902), .B1(
        n18901), .B2(n18913), .ZN(n18880) );
  OAI211_X1 U22030 ( .C1(n18916), .C2(n18905), .A(n18881), .B(n18880), .ZN(
        P3_U2980) );
  AOI22_X1 U22031 ( .A1(n18918), .A2(n18957), .B1(n18917), .B2(n18899), .ZN(
        n18883) );
  AOI22_X1 U22032 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18902), .B1(
        n18901), .B2(n18919), .ZN(n18882) );
  OAI211_X1 U22033 ( .C1(n18922), .C2(n18905), .A(n18883), .B(n18882), .ZN(
        P3_U2981) );
  INV_X1 U22034 ( .A(n18957), .ZN(n18947) );
  AOI22_X1 U22035 ( .A1(n18884), .A2(n18890), .B1(n18923), .B2(n18899), .ZN(
        n18886) );
  AOI22_X1 U22036 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18902), .B1(
        n18901), .B2(n18925), .ZN(n18885) );
  OAI211_X1 U22037 ( .C1(n18887), .C2(n18947), .A(n18886), .B(n18885), .ZN(
        P3_U2982) );
  AOI22_X1 U22038 ( .A1(n18930), .A2(n18957), .B1(n18929), .B2(n18899), .ZN(
        n18889) );
  AOI22_X1 U22039 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18902), .B1(
        n18901), .B2(n18931), .ZN(n18888) );
  OAI211_X1 U22040 ( .C1(n18934), .C2(n18905), .A(n18889), .B(n18888), .ZN(
        P3_U2983) );
  AOI22_X1 U22041 ( .A1(n18936), .A2(n18890), .B1(n18935), .B2(n18899), .ZN(
        n18892) );
  AOI22_X1 U22042 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18902), .B1(
        n18901), .B2(n18937), .ZN(n18891) );
  OAI211_X1 U22043 ( .C1(n18940), .C2(n18947), .A(n18892), .B(n18891), .ZN(
        P3_U2984) );
  AOI22_X1 U22044 ( .A1(n18942), .A2(n18957), .B1(n18941), .B2(n18899), .ZN(
        n18894) );
  AOI22_X1 U22045 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18902), .B1(
        n18901), .B2(n18944), .ZN(n18893) );
  OAI211_X1 U22046 ( .C1(n18948), .C2(n18905), .A(n18894), .B(n18893), .ZN(
        P3_U2985) );
  AOI22_X1 U22047 ( .A1(n18949), .A2(n18899), .B1(n18895), .B2(n18957), .ZN(
        n18897) );
  AOI22_X1 U22048 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18902), .B1(
        n18901), .B2(n18951), .ZN(n18896) );
  OAI211_X1 U22049 ( .C1(n18898), .C2(n18905), .A(n18897), .B(n18896), .ZN(
        P3_U2986) );
  AOI22_X1 U22050 ( .A1(n18900), .A2(n18957), .B1(n18956), .B2(n18899), .ZN(
        n18904) );
  AOI22_X1 U22051 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18902), .B1(
        n18901), .B2(n18959), .ZN(n18903) );
  OAI211_X1 U22052 ( .C1(n18906), .C2(n18905), .A(n18904), .B(n18903), .ZN(
        P3_U2987) );
  INV_X1 U22053 ( .A(n18911), .ZN(n18907) );
  NOR2_X1 U22054 ( .A1(n19042), .A2(n18907), .ZN(n18955) );
  AOI22_X1 U22055 ( .A1(n18909), .A2(n18943), .B1(n18908), .B2(n18955), .ZN(
        n18915) );
  AOI22_X1 U22056 ( .A1(n18545), .A2(n18912), .B1(n18911), .B2(n18910), .ZN(
        n18961) );
  AOI22_X1 U22057 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18961), .B1(
        n18960), .B2(n18913), .ZN(n18914) );
  OAI211_X1 U22058 ( .C1(n18916), .C2(n18947), .A(n18915), .B(n18914), .ZN(
        P3_U2988) );
  AOI22_X1 U22059 ( .A1(n18943), .A2(n18918), .B1(n18917), .B2(n18955), .ZN(
        n18921) );
  AOI22_X1 U22060 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18961), .B1(
        n18960), .B2(n18919), .ZN(n18920) );
  OAI211_X1 U22061 ( .C1(n18922), .C2(n18947), .A(n18921), .B(n18920), .ZN(
        P3_U2989) );
  AOI22_X1 U22062 ( .A1(n18943), .A2(n18924), .B1(n18923), .B2(n18955), .ZN(
        n18927) );
  AOI22_X1 U22063 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18961), .B1(
        n18960), .B2(n18925), .ZN(n18926) );
  OAI211_X1 U22064 ( .C1(n18928), .C2(n18947), .A(n18927), .B(n18926), .ZN(
        P3_U2990) );
  AOI22_X1 U22065 ( .A1(n18943), .A2(n18930), .B1(n18929), .B2(n18955), .ZN(
        n18933) );
  AOI22_X1 U22066 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18961), .B1(
        n18960), .B2(n18931), .ZN(n18932) );
  OAI211_X1 U22067 ( .C1(n18934), .C2(n18947), .A(n18933), .B(n18932), .ZN(
        P3_U2991) );
  AOI22_X1 U22068 ( .A1(n18936), .A2(n18957), .B1(n18935), .B2(n18955), .ZN(
        n18939) );
  AOI22_X1 U22069 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18961), .B1(
        n18960), .B2(n18937), .ZN(n18938) );
  OAI211_X1 U22070 ( .C1(n18965), .C2(n18940), .A(n18939), .B(n18938), .ZN(
        P3_U2992) );
  AOI22_X1 U22071 ( .A1(n18943), .A2(n18942), .B1(n18941), .B2(n18955), .ZN(
        n18946) );
  AOI22_X1 U22072 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18961), .B1(
        n18960), .B2(n18944), .ZN(n18945) );
  OAI211_X1 U22073 ( .C1(n18948), .C2(n18947), .A(n18946), .B(n18945), .ZN(
        P3_U2993) );
  AOI22_X1 U22074 ( .A1(n18950), .A2(n18957), .B1(n18949), .B2(n18955), .ZN(
        n18953) );
  AOI22_X1 U22075 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18961), .B1(
        n18960), .B2(n18951), .ZN(n18952) );
  OAI211_X1 U22076 ( .C1(n18965), .C2(n18954), .A(n18953), .B(n18952), .ZN(
        P3_U2994) );
  AOI22_X1 U22077 ( .A1(n18958), .A2(n18957), .B1(n18956), .B2(n18955), .ZN(
        n18963) );
  AOI22_X1 U22078 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18961), .B1(
        n18960), .B2(n18959), .ZN(n18962) );
  OAI211_X1 U22079 ( .C1(n18965), .C2(n18964), .A(n18963), .B(n18962), .ZN(
        P3_U2995) );
  NOR2_X1 U22080 ( .A1(n19000), .A2(n18966), .ZN(n18968) );
  OAI222_X1 U22081 ( .A1(n18972), .A2(n18971), .B1(n18970), .B2(n18969), .C1(
        n18968), .C2(n18967), .ZN(n19178) );
  OAI21_X1 U22082 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18973), .ZN(n18975) );
  OAI211_X1 U22083 ( .C1(n19001), .C2(n18976), .A(n18975), .B(n18974), .ZN(
        n19024) );
  NOR2_X1 U22084 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18977), .ZN(
        n19005) );
  INV_X1 U22085 ( .A(n19005), .ZN(n18978) );
  AOI22_X1 U22086 ( .A1(n18984), .A2(n18978), .B1(n19000), .B2(n18983), .ZN(
        n18979) );
  NOR2_X1 U22087 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18979), .ZN(
        n19140) );
  OAI21_X1 U22088 ( .B1(n18982), .B2(n18981), .A(n18980), .ZN(n18988) );
  OAI21_X1 U22089 ( .B1(n18984), .B2(n19004), .A(n18983), .ZN(n18985) );
  AOI21_X1 U22090 ( .B1(n18986), .B2(n18988), .A(n18985), .ZN(n19141) );
  AOI21_X1 U22091 ( .B1(n19141), .B2(n19001), .A(n10936), .ZN(n18987) );
  AOI21_X1 U22092 ( .B1(n19001), .B2(n19140), .A(n18987), .ZN(n19022) );
  INV_X1 U22093 ( .A(n19001), .ZN(n19013) );
  AOI21_X1 U22094 ( .B1(n9997), .B2(n18993), .A(n18988), .ZN(n18998) );
  NAND2_X1 U22095 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18989), .ZN(
        n18997) );
  OAI211_X1 U22096 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n18991), .B(n18990), .ZN(
        n18996) );
  NOR2_X1 U22097 ( .A1(n18992), .A2(n9998), .ZN(n18994) );
  OAI211_X1 U22098 ( .C1(n18994), .C2(n18993), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n10935), .ZN(n18995) );
  OAI211_X1 U22099 ( .C1(n18998), .C2(n18997), .A(n18996), .B(n18995), .ZN(
        n18999) );
  AOI21_X1 U22100 ( .B1(n19000), .B2(n19148), .A(n18999), .ZN(n19151) );
  AOI22_X1 U22101 ( .A1(n19013), .A2(n10935), .B1(n19151), .B2(n19001), .ZN(
        n19017) );
  NOR2_X1 U22102 ( .A1(n19003), .A2(n19002), .ZN(n19007) );
  AOI22_X1 U22103 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19004), .B1(
        n19007), .B2(n9716), .ZN(n19161) );
  OAI22_X1 U22104 ( .A1(n19007), .A2(n19006), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n19005), .ZN(n19158) );
  OR3_X1 U22105 ( .A1(n19161), .A2(n19010), .A3(n19008), .ZN(n19009) );
  AOI22_X1 U22106 ( .A1(n19161), .A2(n19010), .B1(n19158), .B2(n19009), .ZN(
        n19012) );
  OAI21_X1 U22107 ( .B1(n19013), .B2(n19012), .A(n19011), .ZN(n19016) );
  AND2_X1 U22108 ( .A1(n19017), .A2(n19016), .ZN(n19014) );
  OAI221_X1 U22109 ( .B1(n19017), .B2(n19016), .C1(n19015), .C2(n19014), .A(
        n19019), .ZN(n19021) );
  AOI21_X1 U22110 ( .B1(n19019), .B2(n19018), .A(n19017), .ZN(n19020) );
  AOI222_X1 U22111 ( .A1(n19022), .A2(n19021), .B1(n19022), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n19021), .C2(n19020), .ZN(
        n19023) );
  NOR4_X1 U22112 ( .A1(n19025), .A2(n19178), .A3(n19024), .A4(n19023), .ZN(
        n19037) );
  INV_X1 U22113 ( .A(n19149), .ZN(n19160) );
  AOI22_X1 U22114 ( .A1(n19160), .A2(n19189), .B1(n19182), .B2(n17761), .ZN(
        n19026) );
  INV_X1 U22115 ( .A(n19026), .ZN(n19032) );
  OAI211_X1 U22116 ( .C1(n19028), .C2(n19027), .A(n19180), .B(n19037), .ZN(
        n19137) );
  NAND2_X1 U22117 ( .A1(n19182), .A2(n19029), .ZN(n19038) );
  NAND2_X1 U22118 ( .A1(n19137), .A2(n19038), .ZN(n19040) );
  NOR2_X1 U22119 ( .A1(n19030), .A2(n19040), .ZN(n19031) );
  MUX2_X1 U22120 ( .A(n19032), .B(n19031), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n19035) );
  NAND2_X1 U22121 ( .A1(n19033), .A2(n19042), .ZN(n19034) );
  OAI211_X1 U22122 ( .C1(n19037), .C2(n19036), .A(n19035), .B(n19034), .ZN(
        P3_U2996) );
  NOR2_X1 U22123 ( .A1(n19187), .A2(n19181), .ZN(n19044) );
  NOR3_X1 U22124 ( .A1(n19147), .A2(n19039), .A3(n19038), .ZN(n19047) );
  NOR3_X1 U22125 ( .A1(n19042), .A2(n19041), .A3(n19040), .ZN(n19043) );
  OR4_X1 U22126 ( .A1(n19045), .A2(n19044), .A3(n19047), .A4(n19043), .ZN(
        P3_U2997) );
  NOR4_X1 U22127 ( .A1(n19189), .A2(n19048), .A3(n19047), .A4(n19046), .ZN(
        P3_U2998) );
  AND2_X1 U22128 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n19049), .ZN(
        P3_U2999) );
  AND2_X1 U22129 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n19049), .ZN(
        P3_U3000) );
  AND2_X1 U22130 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n19049), .ZN(
        P3_U3001) );
  AND2_X1 U22131 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n19049), .ZN(
        P3_U3002) );
  AND2_X1 U22132 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n19049), .ZN(
        P3_U3003) );
  AND2_X1 U22133 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n19049), .ZN(
        P3_U3004) );
  AND2_X1 U22134 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n19049), .ZN(
        P3_U3005) );
  AND2_X1 U22135 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n19049), .ZN(
        P3_U3006) );
  AND2_X1 U22136 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n19049), .ZN(
        P3_U3007) );
  AND2_X1 U22137 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n19049), .ZN(
        P3_U3008) );
  AND2_X1 U22138 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n19049), .ZN(
        P3_U3009) );
  AND2_X1 U22139 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n19049), .ZN(
        P3_U3010) );
  AND2_X1 U22140 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n19049), .ZN(
        P3_U3011) );
  AND2_X1 U22141 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n19049), .ZN(
        P3_U3012) );
  AND2_X1 U22142 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n19049), .ZN(
        P3_U3013) );
  AND2_X1 U22143 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n19049), .ZN(
        P3_U3014) );
  AND2_X1 U22144 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n19049), .ZN(
        P3_U3015) );
  AND2_X1 U22145 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n19049), .ZN(
        P3_U3016) );
  AND2_X1 U22146 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n19049), .ZN(
        P3_U3017) );
  AND2_X1 U22147 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n19049), .ZN(
        P3_U3018) );
  AND2_X1 U22148 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n19049), .ZN(
        P3_U3019) );
  AND2_X1 U22149 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n19049), .ZN(
        P3_U3020) );
  AND2_X1 U22150 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n19049), .ZN(P3_U3021) );
  AND2_X1 U22151 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n19049), .ZN(P3_U3022) );
  AND2_X1 U22152 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n19049), .ZN(P3_U3023) );
  AND2_X1 U22153 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n19049), .ZN(P3_U3024) );
  AND2_X1 U22154 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n19049), .ZN(P3_U3025) );
  AND2_X1 U22155 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n19049), .ZN(P3_U3026) );
  AND2_X1 U22156 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n19049), .ZN(P3_U3027) );
  AND2_X1 U22157 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n19049), .ZN(P3_U3028) );
  NAND2_X1 U22158 ( .A1(n19182), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n19059) );
  INV_X1 U22159 ( .A(n19059), .ZN(n19057) );
  OAI21_X1 U22160 ( .B1(n19050), .B2(n20946), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19051) );
  AOI22_X1 U22161 ( .A1(n19057), .A2(n19065), .B1(n19194), .B2(n19051), .ZN(
        n19053) );
  INV_X1 U22162 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n19052) );
  NAND3_X1 U22163 ( .A1(NA), .A2(n19063), .A3(n19052), .ZN(n19058) );
  OAI211_X1 U22164 ( .C1(P3_STATE_REG_0__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n19053), .B(n19058), .ZN(P3_U3029) );
  NOR2_X1 U22165 ( .A1(n19065), .A2(n20946), .ZN(n19061) );
  NOR2_X1 U22166 ( .A1(n19063), .A2(n19061), .ZN(n19054) );
  AOI21_X1 U22167 ( .B1(n19054), .B2(P3_REQUESTPENDING_REG_SCAN_IN), .A(n19057), .ZN(n19055) );
  OAI211_X1 U22168 ( .C1(n20946), .C2(n19056), .A(n19055), .B(n19184), .ZN(
        P3_U3030) );
  AOI21_X1 U22169 ( .B1(n19063), .B2(n19058), .A(n19057), .ZN(n19064) );
  OAI22_X1 U22170 ( .A1(NA), .A2(n19059), .B1(P3_STATE_REG_1__SCAN_IN), .B2(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n19060) );
  OAI22_X1 U22171 ( .A1(n19061), .A2(n19060), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n19062) );
  OAI22_X1 U22172 ( .A1(n19064), .A2(n19065), .B1(n19063), .B2(n19062), .ZN(
        P3_U3031) );
  OAI222_X1 U22173 ( .A1(n19067), .A2(n19129), .B1(n19066), .B2(n19126), .C1(
        n19068), .C2(n19124), .ZN(P3_U3032) );
  INV_X1 U22174 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n19070) );
  OAI222_X1 U22175 ( .A1(n19124), .A2(n19070), .B1(n19069), .B2(n19126), .C1(
        n19068), .C2(n19129), .ZN(P3_U3033) );
  OAI222_X1 U22176 ( .A1(n19124), .A2(n19072), .B1(n19071), .B2(n19126), .C1(
        n19070), .C2(n19129), .ZN(P3_U3034) );
  INV_X1 U22177 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n19075) );
  OAI222_X1 U22178 ( .A1(n19124), .A2(n19075), .B1(n19073), .B2(n19126), .C1(
        n19072), .C2(n19129), .ZN(P3_U3035) );
  OAI222_X1 U22179 ( .A1(n19075), .A2(n19129), .B1(n19074), .B2(n19126), .C1(
        n19076), .C2(n19124), .ZN(P3_U3036) );
  OAI222_X1 U22180 ( .A1(n19124), .A2(n19078), .B1(n19077), .B2(n19126), .C1(
        n19076), .C2(n19129), .ZN(P3_U3037) );
  OAI222_X1 U22181 ( .A1(n19124), .A2(n19080), .B1(n19079), .B2(n19126), .C1(
        n19078), .C2(n19129), .ZN(P3_U3038) );
  OAI222_X1 U22182 ( .A1(n19124), .A2(n19082), .B1(n19081), .B2(n19126), .C1(
        n19080), .C2(n19129), .ZN(P3_U3039) );
  OAI222_X1 U22183 ( .A1(n19124), .A2(n19084), .B1(n19083), .B2(n19126), .C1(
        n19082), .C2(n19129), .ZN(P3_U3040) );
  INV_X1 U22184 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n19086) );
  OAI222_X1 U22185 ( .A1(n19124), .A2(n19086), .B1(n19085), .B2(n19126), .C1(
        n19084), .C2(n19129), .ZN(P3_U3041) );
  OAI222_X1 U22186 ( .A1(n19124), .A2(n19088), .B1(n19087), .B2(n19126), .C1(
        n19086), .C2(n19129), .ZN(P3_U3042) );
  OAI222_X1 U22187 ( .A1(n19124), .A2(n19090), .B1(n19089), .B2(n19126), .C1(
        n19088), .C2(n19129), .ZN(P3_U3043) );
  OAI222_X1 U22188 ( .A1(n19124), .A2(n19093), .B1(n19091), .B2(n19126), .C1(
        n19090), .C2(n19129), .ZN(P3_U3044) );
  OAI222_X1 U22189 ( .A1(n19093), .A2(n19129), .B1(n19092), .B2(n19126), .C1(
        n19094), .C2(n19124), .ZN(P3_U3045) );
  OAI222_X1 U22190 ( .A1(n19124), .A2(n19096), .B1(n19095), .B2(n19126), .C1(
        n19094), .C2(n19129), .ZN(P3_U3046) );
  OAI222_X1 U22191 ( .A1(n19124), .A2(n19099), .B1(n19097), .B2(n19126), .C1(
        n19096), .C2(n19129), .ZN(P3_U3047) );
  OAI222_X1 U22192 ( .A1(n19099), .A2(n19129), .B1(n19098), .B2(n19126), .C1(
        n19100), .C2(n19124), .ZN(P3_U3048) );
  INV_X1 U22193 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n19102) );
  OAI222_X1 U22194 ( .A1(n19124), .A2(n19102), .B1(n19101), .B2(n19126), .C1(
        n19100), .C2(n19129), .ZN(P3_U3049) );
  OAI222_X1 U22195 ( .A1(n19124), .A2(n19104), .B1(n19103), .B2(n19126), .C1(
        n19102), .C2(n19129), .ZN(P3_U3050) );
  OAI222_X1 U22196 ( .A1(n19124), .A2(n19107), .B1(n19105), .B2(n19126), .C1(
        n19104), .C2(n19129), .ZN(P3_U3051) );
  OAI222_X1 U22197 ( .A1(n19107), .A2(n19129), .B1(n19106), .B2(n19126), .C1(
        n19108), .C2(n19124), .ZN(P3_U3052) );
  OAI222_X1 U22198 ( .A1(n19124), .A2(n19111), .B1(n19109), .B2(n19126), .C1(
        n19108), .C2(n19129), .ZN(P3_U3053) );
  OAI222_X1 U22199 ( .A1(n19111), .A2(n19129), .B1(n19110), .B2(n19126), .C1(
        n19112), .C2(n19124), .ZN(P3_U3054) );
  OAI222_X1 U22200 ( .A1(n19124), .A2(n19114), .B1(n19113), .B2(n19126), .C1(
        n19112), .C2(n19129), .ZN(P3_U3055) );
  OAI222_X1 U22201 ( .A1(n19124), .A2(n19116), .B1(n19115), .B2(n19126), .C1(
        n19114), .C2(n19129), .ZN(P3_U3056) );
  OAI222_X1 U22202 ( .A1(n19124), .A2(n19118), .B1(n19117), .B2(n19126), .C1(
        n19116), .C2(n19129), .ZN(P3_U3057) );
  INV_X1 U22203 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n19121) );
  OAI222_X1 U22204 ( .A1(n19124), .A2(n19121), .B1(n19119), .B2(n19126), .C1(
        n19118), .C2(n19129), .ZN(P3_U3058) );
  OAI222_X1 U22205 ( .A1(n19121), .A2(n19129), .B1(n19120), .B2(n19126), .C1(
        n19122), .C2(n19124), .ZN(P3_U3059) );
  OAI222_X1 U22206 ( .A1(n19124), .A2(n19128), .B1(n19123), .B2(n19126), .C1(
        n19122), .C2(n19129), .ZN(P3_U3060) );
  INV_X1 U22207 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19127) );
  OAI222_X1 U22208 ( .A1(n19129), .A2(n19128), .B1(n19127), .B2(n19126), .C1(
        n19125), .C2(n19124), .ZN(P3_U3061) );
  MUX2_X1 U22209 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .B(P3_BE_N_REG_3__SCAN_IN), .S(n19194), .Z(P3_U3274) );
  MUX2_X1 U22210 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .B(P3_BE_N_REG_2__SCAN_IN), .S(n19194), .Z(P3_U3275) );
  OAI22_X1 U22211 ( .A1(n19194), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n19126), .ZN(n19130) );
  INV_X1 U22212 ( .A(n19130), .ZN(P3_U3276) );
  OAI22_X1 U22213 ( .A1(n19194), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n19126), .ZN(n19131) );
  INV_X1 U22214 ( .A(n19131), .ZN(P3_U3277) );
  OAI21_X1 U22215 ( .B1(n19135), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n19133), 
        .ZN(n19132) );
  INV_X1 U22216 ( .A(n19132), .ZN(P3_U3280) );
  OAI21_X1 U22217 ( .B1(n19135), .B2(n19134), .A(n19133), .ZN(P3_U3281) );
  OAI221_X1 U22218 ( .B1(n19138), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n19138), 
        .C2(n19137), .A(n19136), .ZN(P3_U3282) );
  INV_X1 U22219 ( .A(n19150), .ZN(n19162) );
  AOI22_X1 U22220 ( .A1(n19162), .A2(n19140), .B1(n19160), .B2(n19139), .ZN(
        n19144) );
  INV_X1 U22221 ( .A(n19166), .ZN(n19164) );
  OAI21_X1 U22222 ( .B1(n19150), .B2(n19141), .A(n19164), .ZN(n19142) );
  INV_X1 U22223 ( .A(n19142), .ZN(n19143) );
  OAI22_X1 U22224 ( .A1(n19166), .A2(n19144), .B1(n19143), .B2(n10936), .ZN(
        P3_U3285) );
  OAI22_X1 U22225 ( .A1(n19146), .A2(n19145), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n19156) );
  INV_X1 U22226 ( .A(n19156), .ZN(n19153) );
  NOR2_X1 U22227 ( .A1(n19147), .A2(n19163), .ZN(n19155) );
  OAI22_X1 U22228 ( .A1(n19151), .A2(n19150), .B1(n19149), .B2(n19148), .ZN(
        n19152) );
  AOI21_X1 U22229 ( .B1(n19153), .B2(n19155), .A(n19152), .ZN(n19154) );
  AOI22_X1 U22230 ( .A1(n19166), .A2(n10935), .B1(n19154), .B2(n19164), .ZN(
        P3_U3288) );
  AOI222_X1 U22231 ( .A1(n19158), .A2(n19162), .B1(n19160), .B2(n19157), .C1(
        n19156), .C2(n19155), .ZN(n19159) );
  AOI22_X1 U22232 ( .A1(n19166), .A2(n9997), .B1(n19159), .B2(n19164), .ZN(
        P3_U3289) );
  AOI222_X1 U22233 ( .A1(n19163), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n19162), 
        .B2(n19161), .C1(n9716), .C2(n19160), .ZN(n19165) );
  AOI22_X1 U22234 ( .A1(n19166), .A2(n9715), .B1(n19165), .B2(n19164), .ZN(
        P3_U3290) );
  INV_X1 U22235 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n19173) );
  INV_X1 U22236 ( .A(n19167), .ZN(n19174) );
  AOI211_X1 U22237 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(n19168), 
        .ZN(n19169) );
  AOI21_X1 U22238 ( .B1(P3_BYTEENABLE_REG_2__SCAN_IN), .B2(n19174), .A(n19169), 
        .ZN(n19170) );
  OAI21_X1 U22239 ( .B1(n19173), .B2(n19171), .A(n19170), .ZN(P3_U3292) );
  INV_X1 U22240 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19175) );
  NOR2_X1 U22241 ( .A1(n19174), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n19172) );
  AOI22_X1 U22242 ( .A1(n19175), .A2(n19174), .B1(n19173), .B2(n19172), .ZN(
        P3_U3293) );
  INV_X1 U22243 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n19176) );
  AOI22_X1 U22244 ( .A1(n19126), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n19176), 
        .B2(n19194), .ZN(P3_U3294) );
  MUX2_X1 U22245 ( .A(P3_MORE_REG_SCAN_IN), .B(n19178), .S(n19177), .Z(
        P3_U3295) );
  OAI22_X1 U22246 ( .A1(n19182), .A2(n19181), .B1(n19180), .B2(n19179), .ZN(
        n19183) );
  NOR2_X1 U22247 ( .A1(n19202), .A2(n19183), .ZN(n19193) );
  AOI21_X1 U22248 ( .B1(n19186), .B2(n19185), .A(n19184), .ZN(n19188) );
  OAI211_X1 U22249 ( .C1(n19195), .C2(n19188), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n19187), .ZN(n19190) );
  AOI21_X1 U22250 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n19190), .A(n19189), 
        .ZN(n19192) );
  NAND2_X1 U22251 ( .A1(n19193), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n19191) );
  OAI21_X1 U22252 ( .B1(n19193), .B2(n19192), .A(n19191), .ZN(P3_U3296) );
  MUX2_X1 U22253 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .B(P3_M_IO_N_REG_SCAN_IN), 
        .S(n19194), .Z(P3_U3297) );
  INV_X1 U22254 ( .A(n19195), .ZN(n19197) );
  OAI21_X1 U22255 ( .B1(n19199), .B2(P3_READREQUEST_REG_SCAN_IN), .A(n19198), 
        .ZN(n19196) );
  OAI21_X1 U22256 ( .B1(n19198), .B2(n19197), .A(n19196), .ZN(P3_U3298) );
  NOR2_X1 U22257 ( .A1(n19199), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n19201)
         );
  OAI21_X1 U22258 ( .B1(n19202), .B2(n19201), .A(n19200), .ZN(P3_U3299) );
  INV_X1 U22259 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n20101) );
  NAND2_X1 U22260 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20101), .ZN(n20093) );
  NOR2_X1 U22261 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(P2_STATE_REG_1__SCAN_IN), 
        .ZN(n20090) );
  INV_X1 U22262 ( .A(n20090), .ZN(n19203) );
  OAI21_X1 U22263 ( .B1(n20086), .B2(n20093), .A(n19203), .ZN(n20158) );
  AOI21_X1 U22264 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n20158), .ZN(n19204) );
  INV_X1 U22265 ( .A(n19204), .ZN(P2_U2815) );
  INV_X1 U22266 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n19207) );
  OAI22_X1 U22267 ( .A1(n19208), .A2(n19207), .B1(n19206), .B2(n19205), .ZN(
        P2_U2816) );
  AOI22_X1 U22268 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(n20234), .B1(n20094), .B2(
        n20086), .ZN(n19209) );
  OAI21_X1 U22269 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n20234), .A(n19209), 
        .ZN(P2_U2817) );
  OAI21_X1 U22270 ( .B1(n20094), .B2(BS16), .A(n20158), .ZN(n20156) );
  OAI21_X1 U22271 ( .B1(n20158), .B2(n20226), .A(n20156), .ZN(P2_U2818) );
  NOR2_X1 U22272 ( .A1(n19211), .A2(n19210), .ZN(n20211) );
  OAI21_X1 U22273 ( .B1(n20211), .B2(n19213), .A(n19212), .ZN(P2_U2819) );
  NOR4_X1 U22274 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19217) );
  NOR4_X1 U22275 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19216) );
  NOR4_X1 U22276 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19215) );
  NOR4_X1 U22277 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19214) );
  NAND4_X1 U22278 ( .A1(n19217), .A2(n19216), .A3(n19215), .A4(n19214), .ZN(
        n19223) );
  NOR4_X1 U22279 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19221) );
  AOI211_X1 U22280 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19220) );
  NOR4_X1 U22281 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19219) );
  NOR4_X1 U22282 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19218) );
  NAND4_X1 U22283 ( .A1(n19221), .A2(n19220), .A3(n19219), .A4(n19218), .ZN(
        n19222) );
  NOR2_X1 U22284 ( .A1(n19223), .A2(n19222), .ZN(n19234) );
  INV_X1 U22285 ( .A(n19234), .ZN(n19232) );
  NOR2_X1 U22286 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n19232), .ZN(n19226) );
  INV_X1 U22287 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19224) );
  AOI22_X1 U22288 ( .A1(n19226), .A2(n19227), .B1(n19232), .B2(n19224), .ZN(
        P2_U2820) );
  OR3_X1 U22289 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n19231) );
  INV_X1 U22290 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19225) );
  AOI22_X1 U22291 ( .A1(n19226), .A2(n19231), .B1(n19232), .B2(n19225), .ZN(
        P2_U2821) );
  INV_X1 U22292 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20157) );
  NAND2_X1 U22293 ( .A1(n19226), .A2(n20157), .ZN(n19230) );
  OAI21_X1 U22294 ( .B1(n20102), .B2(n19227), .A(n19234), .ZN(n19228) );
  OAI21_X1 U22295 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n19234), .A(n19228), 
        .ZN(n19229) );
  OAI221_X1 U22296 ( .B1(n19230), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n19230), .C2(P2_REIP_REG_0__SCAN_IN), .A(n19229), .ZN(P2_U2822) );
  INV_X1 U22297 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19233) );
  OAI221_X1 U22298 ( .B1(n19234), .B2(n19233), .C1(n19232), .C2(n19231), .A(
        n19230), .ZN(P2_U2823) );
  NAND2_X1 U22299 ( .A1(n19235), .A2(n19237), .ZN(n19254) );
  INV_X1 U22300 ( .A(n19245), .ZN(n19236) );
  AOI211_X1 U22301 ( .C1(n19384), .C2(n19237), .A(n19236), .B(n19411), .ZN(
        n19239) );
  OAI22_X1 U22302 ( .A1(n19413), .A2(n10011), .B1(n20131), .B2(n19417), .ZN(
        n19238) );
  AOI211_X1 U22303 ( .C1(n19431), .C2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n19239), .B(n19238), .ZN(n19244) );
  AOI222_X1 U22304 ( .A1(n19242), .A2(n19361), .B1(n19241), .B2(n19403), .C1(
        n19240), .C2(n19441), .ZN(n19243) );
  OAI211_X1 U22305 ( .C1(n19245), .C2(n19254), .A(n19244), .B(n19243), .ZN(
        P2_U2834) );
  INV_X1 U22306 ( .A(n19246), .ZN(n19252) );
  AOI22_X1 U22307 ( .A1(n19437), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19431), .ZN(n19247) );
  OAI21_X1 U22308 ( .B1(n19248), .B2(n19400), .A(n19247), .ZN(n19249) );
  AOI21_X1 U22309 ( .B1(n19250), .B2(n19441), .A(n19249), .ZN(n19251) );
  OAI21_X1 U22310 ( .B1(n19252), .B2(n19434), .A(n19251), .ZN(n19253) );
  AOI21_X1 U22311 ( .B1(n9778), .B2(n19361), .A(n19253), .ZN(n19258) );
  INV_X1 U22312 ( .A(n19254), .ZN(n19255) );
  OAI21_X1 U22313 ( .B1(n19256), .B2(n19260), .A(n19255), .ZN(n19257) );
  OAI211_X1 U22314 ( .C1(n19260), .C2(n19259), .A(n19258), .B(n19257), .ZN(
        P2_U2835) );
  NAND2_X1 U22315 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n19431), .ZN(
        n19261) );
  OAI211_X1 U22316 ( .C1(n19417), .C2(n20127), .A(n19341), .B(n19261), .ZN(
        n19262) );
  AOI21_X1 U22317 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n19432), .A(n19262), .ZN(
        n19263) );
  OAI21_X1 U22318 ( .B1(n19264), .B2(n19434), .A(n19263), .ZN(n19265) );
  INV_X1 U22319 ( .A(n19265), .ZN(n19272) );
  NAND2_X1 U22320 ( .A1(n19384), .A2(n19266), .ZN(n19268) );
  XNOR2_X1 U22321 ( .A(n19268), .B(n19267), .ZN(n19270) );
  AOI22_X1 U22322 ( .A1(n19270), .A2(n19443), .B1(n19269), .B2(n19441), .ZN(
        n19271) );
  OAI211_X1 U22323 ( .C1(n19273), .C2(n19447), .A(n19272), .B(n19271), .ZN(
        P2_U2836) );
  NOR2_X1 U22324 ( .A1(n19419), .A2(n19274), .ZN(n19276) );
  XOR2_X1 U22325 ( .A(n19276), .B(n19275), .Z(n19287) );
  OAI22_X1 U22326 ( .A1(n19400), .A2(n19277), .B1(n19397), .B2(n9810), .ZN(
        n19278) );
  INV_X1 U22327 ( .A(n19278), .ZN(n19279) );
  OAI21_X1 U22328 ( .B1(n19280), .B2(n19434), .A(n19279), .ZN(n19281) );
  AOI211_X1 U22329 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n19437), .A(n19500), 
        .B(n19281), .ZN(n19286) );
  INV_X1 U22330 ( .A(n19282), .ZN(n19283) );
  AOI22_X1 U22331 ( .A1(n19284), .A2(n19361), .B1(n19283), .B2(n19441), .ZN(
        n19285) );
  OAI211_X1 U22332 ( .C1(n19411), .C2(n19287), .A(n19286), .B(n19285), .ZN(
        P2_U2837) );
  NAND2_X1 U22333 ( .A1(n19384), .A2(n19288), .ZN(n19289) );
  XOR2_X1 U22334 ( .A(n19290), .B(n19289), .Z(n19300) );
  NOR2_X1 U22335 ( .A1(n19417), .A2(n20123), .ZN(n19291) );
  AOI211_X1 U22336 ( .C1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n19431), .A(
        n19500), .B(n19291), .ZN(n19292) );
  OAI21_X1 U22337 ( .B1(n19293), .B2(n19400), .A(n19292), .ZN(n19294) );
  AOI21_X1 U22338 ( .B1(n19295), .B2(n19403), .A(n19294), .ZN(n19299) );
  AOI22_X1 U22339 ( .A1(n19297), .A2(n19361), .B1(n19296), .B2(n19441), .ZN(
        n19298) );
  OAI211_X1 U22340 ( .C1(n19411), .C2(n19300), .A(n19299), .B(n19298), .ZN(
        P2_U2838) );
  NOR2_X1 U22341 ( .A1(n19419), .A2(n19301), .ZN(n19303) );
  XOR2_X1 U22342 ( .A(n19303), .B(n19302), .Z(n19313) );
  OR2_X1 U22343 ( .A1(n19304), .A2(n19434), .ZN(n19308) );
  NAND2_X1 U22344 ( .A1(n19431), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n19305) );
  OAI211_X1 U22345 ( .C1(n19417), .C2(n15977), .A(n19341), .B(n19305), .ZN(
        n19306) );
  AOI21_X1 U22346 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n19432), .A(n19306), .ZN(
        n19307) );
  AND2_X1 U22347 ( .A1(n19308), .A2(n19307), .ZN(n19312) );
  AOI22_X1 U22348 ( .A1(n19310), .A2(n19361), .B1(n19309), .B2(n19441), .ZN(
        n19311) );
  OAI211_X1 U22349 ( .C1(n19411), .C2(n19313), .A(n19312), .B(n19311), .ZN(
        P2_U2839) );
  NOR2_X1 U22350 ( .A1(n19417), .A2(n20120), .ZN(n19314) );
  AOI211_X1 U22351 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n19431), .A(
        n19500), .B(n19314), .ZN(n19315) );
  OAI21_X1 U22352 ( .B1(n19316), .B2(n19400), .A(n19315), .ZN(n19317) );
  AOI21_X1 U22353 ( .B1(n19318), .B2(n19403), .A(n19317), .ZN(n19325) );
  NAND2_X1 U22354 ( .A1(n19384), .A2(n19319), .ZN(n19320) );
  XNOR2_X1 U22355 ( .A(n19321), .B(n19320), .ZN(n19323) );
  AOI22_X1 U22356 ( .A1(n19323), .A2(n19443), .B1(n19322), .B2(n19441), .ZN(
        n19324) );
  OAI211_X1 U22357 ( .C1(n19326), .C2(n19447), .A(n19325), .B(n19324), .ZN(
        P2_U2840) );
  NOR2_X1 U22358 ( .A1(n19419), .A2(n19337), .ZN(n19328) );
  XOR2_X1 U22359 ( .A(n19328), .B(n19327), .Z(n19335) );
  OAI21_X1 U22360 ( .B1(n11567), .B2(n19417), .A(n19395), .ZN(n19331) );
  OAI22_X1 U22361 ( .A1(n19329), .A2(n19434), .B1(n10768), .B2(n19400), .ZN(
        n19330) );
  AOI211_X1 U22362 ( .C1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n19431), .A(
        n19331), .B(n19330), .ZN(n19334) );
  AOI22_X1 U22363 ( .A1(n19332), .A2(n19441), .B1(n19454), .B2(n19361), .ZN(
        n19333) );
  OAI211_X1 U22364 ( .C1(n19411), .C2(n19335), .A(n19334), .B(n19333), .ZN(
        P2_U2841) );
  AOI211_X1 U22365 ( .C1(n19348), .C2(n19338), .A(n19337), .B(n19336), .ZN(
        n19346) );
  NAND2_X1 U22366 ( .A1(n19339), .A2(n19403), .ZN(n19344) );
  NAND2_X1 U22367 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19431), .ZN(
        n19340) );
  OAI211_X1 U22368 ( .C1(n19417), .C2(n11564), .A(n19341), .B(n19340), .ZN(
        n19342) );
  AOI21_X1 U22369 ( .B1(P2_EBX_REG_13__SCAN_IN), .B2(n19432), .A(n19342), .ZN(
        n19343) );
  NAND2_X1 U22370 ( .A1(n19344), .A2(n19343), .ZN(n19345) );
  NOR2_X1 U22371 ( .A1(n19346), .A2(n19345), .ZN(n19351) );
  AOI22_X1 U22372 ( .A1(n19349), .A2(n19348), .B1(n19347), .B2(n19441), .ZN(
        n19350) );
  OAI211_X1 U22373 ( .C1(n19352), .C2(n19447), .A(n19351), .B(n19350), .ZN(
        P2_U2842) );
  NOR2_X1 U22374 ( .A1(n19419), .A2(n19353), .ZN(n19355) );
  XOR2_X1 U22375 ( .A(n19355), .B(n19354), .Z(n19364) );
  NAND2_X1 U22376 ( .A1(n19356), .A2(n19403), .ZN(n19358) );
  NAND2_X1 U22377 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19431), .ZN(
        n19357) );
  OAI211_X1 U22378 ( .C1(n19413), .C2(n19359), .A(n19358), .B(n19357), .ZN(
        n19360) );
  AOI211_X1 U22379 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19437), .A(n19500), 
        .B(n19360), .ZN(n19363) );
  AOI22_X1 U22380 ( .A1(n10090), .A2(n19441), .B1(n19458), .B2(n19361), .ZN(
        n19362) );
  OAI211_X1 U22381 ( .C1(n19411), .C2(n19364), .A(n19363), .B(n19362), .ZN(
        P2_U2843) );
  AOI21_X1 U22382 ( .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n19431), .A(
        n19500), .ZN(n19365) );
  OAI21_X1 U22383 ( .B1(n19417), .B2(n11523), .A(n19365), .ZN(n19370) );
  INV_X1 U22384 ( .A(n19366), .ZN(n19368) );
  AOI211_X1 U22385 ( .C1(P2_EBX_REG_11__SCAN_IN), .C2(n19368), .A(n19434), .B(
        n19367), .ZN(n19369) );
  AOI211_X1 U22386 ( .C1(n19432), .C2(P2_EBX_REG_11__SCAN_IN), .A(n19370), .B(
        n19369), .ZN(n19377) );
  NAND2_X1 U22387 ( .A1(n19384), .A2(n19371), .ZN(n19372) );
  XNOR2_X1 U22388 ( .A(n19373), .B(n19372), .ZN(n19375) );
  AOI22_X1 U22389 ( .A1(n19375), .A2(n19443), .B1(n19374), .B2(n19441), .ZN(
        n19376) );
  OAI211_X1 U22390 ( .C1(n19378), .C2(n19447), .A(n19377), .B(n19376), .ZN(
        P2_U2844) );
  AOI22_X1 U22391 ( .A1(n19379), .A2(n19403), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n19432), .ZN(n19380) );
  OAI21_X1 U22392 ( .B1(n19381), .B2(n19397), .A(n19380), .ZN(n19382) );
  AOI211_X1 U22393 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n19437), .A(n19500), .B(
        n19382), .ZN(n19390) );
  NAND2_X1 U22394 ( .A1(n19384), .A2(n19383), .ZN(n19385) );
  XNOR2_X1 U22395 ( .A(n19386), .B(n19385), .ZN(n19388) );
  AOI22_X1 U22396 ( .A1(n19388), .A2(n19443), .B1(n19387), .B2(n19441), .ZN(
        n19389) );
  OAI211_X1 U22397 ( .C1(n19391), .C2(n19447), .A(n19390), .B(n19389), .ZN(
        P2_U2846) );
  NAND2_X1 U22398 ( .A1(n19384), .A2(n19392), .ZN(n19393) );
  XOR2_X1 U22399 ( .A(n19394), .B(n19393), .Z(n19410) );
  OAI21_X1 U22400 ( .B1(n19397), .B2(n19396), .A(n19395), .ZN(n19398) );
  AOI21_X1 U22401 ( .B1(n19437), .B2(P2_REIP_REG_7__SCAN_IN), .A(n19398), .ZN(
        n19399) );
  OAI21_X1 U22402 ( .B1(n19401), .B2(n19400), .A(n19399), .ZN(n19402) );
  AOI21_X1 U22403 ( .B1(n19404), .B2(n19403), .A(n19402), .ZN(n19409) );
  OAI22_X1 U22404 ( .A1(n19406), .A2(n19447), .B1(n19405), .B2(n19422), .ZN(
        n19407) );
  INV_X1 U22405 ( .A(n19407), .ZN(n19408) );
  OAI211_X1 U22406 ( .C1(n19411), .C2(n19410), .A(n19409), .B(n19408), .ZN(
        P2_U2848) );
  OAI22_X1 U22407 ( .A1(n19414), .A2(n19434), .B1(n19413), .B2(n19412), .ZN(
        n19415) );
  INV_X1 U22408 ( .A(n19415), .ZN(n19416) );
  OAI211_X1 U22409 ( .C1(n20109), .C2(n19417), .A(n19395), .B(n19416), .ZN(
        n19429) );
  NOR2_X1 U22410 ( .A1(n19419), .A2(n19418), .ZN(n19420) );
  XNOR2_X1 U22411 ( .A(n19421), .B(n19420), .ZN(n19426) );
  OAI22_X1 U22412 ( .A1(n19424), .A2(n19447), .B1(n19423), .B2(n19422), .ZN(
        n19425) );
  AOI21_X1 U22413 ( .B1(n19426), .B2(n19443), .A(n19425), .ZN(n19427) );
  INV_X1 U22414 ( .A(n19427), .ZN(n19428) );
  AOI211_X1 U22415 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19431), .A(
        n19429), .B(n19428), .ZN(n19430) );
  INV_X1 U22416 ( .A(n19430), .ZN(P2_U2849) );
  AOI22_X1 U22417 ( .A1(n19432), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19431), .ZN(n19433) );
  OAI21_X1 U22418 ( .B1(n19435), .B2(n19434), .A(n19433), .ZN(n19436) );
  AOI211_X1 U22419 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19437), .A(n19500), .B(
        n19436), .ZN(n19446) );
  NAND2_X1 U22420 ( .A1(n19384), .A2(n19438), .ZN(n19439) );
  XNOR2_X1 U22421 ( .A(n19440), .B(n19439), .ZN(n19444) );
  AOI22_X1 U22422 ( .A1(n19444), .A2(n19443), .B1(n19442), .B2(n19441), .ZN(
        n19445) );
  OAI211_X1 U22423 ( .C1(n19447), .C2(n19470), .A(n19446), .B(n19445), .ZN(
        P2_U2850) );
  AOI22_X1 U22424 ( .A1(n19450), .A2(BUF2_REG_31__SCAN_IN), .B1(n19449), .B2(
        n19448), .ZN(n19453) );
  AOI22_X1 U22425 ( .A1(n19451), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19462), .ZN(n19452) );
  NAND2_X1 U22426 ( .A1(n19453), .A2(n19452), .ZN(P2_U2888) );
  INV_X1 U22427 ( .A(n19454), .ZN(n19457) );
  AOI22_X1 U22428 ( .A1(n19464), .A2(n19455), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19462), .ZN(n19456) );
  OAI21_X1 U22429 ( .B1(n19471), .B2(n19457), .A(n19456), .ZN(P2_U2905) );
  INV_X1 U22430 ( .A(n19458), .ZN(n19461) );
  AOI22_X1 U22431 ( .A1(n19464), .A2(n19459), .B1(P2_EAX_REG_12__SCAN_IN), 
        .B2(n19462), .ZN(n19460) );
  OAI21_X1 U22432 ( .B1(n19471), .B2(n19461), .A(n19460), .ZN(P2_U2907) );
  AOI22_X1 U22433 ( .A1(n19464), .A2(n19463), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19462), .ZN(n19469) );
  OR3_X1 U22434 ( .A1(n19467), .A2(n19466), .A3(n19465), .ZN(n19468) );
  OAI211_X1 U22435 ( .C1(n19471), .C2(n19470), .A(n19469), .B(n19468), .ZN(
        P2_U2914) );
  AND2_X1 U22436 ( .A1(n19484), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22437 ( .A1(n19497), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19473) );
  OAI21_X1 U22438 ( .B1(n13453), .B2(n19499), .A(n19473), .ZN(P2_U2936) );
  AOI22_X1 U22439 ( .A1(n19497), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19474) );
  OAI21_X1 U22440 ( .B1(n11584), .B2(n19499), .A(n19474), .ZN(P2_U2937) );
  AOI22_X1 U22441 ( .A1(n19497), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19475) );
  OAI21_X1 U22442 ( .B1(n13426), .B2(n19499), .A(n19475), .ZN(P2_U2938) );
  AOI22_X1 U22443 ( .A1(n19497), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19476) );
  OAI21_X1 U22444 ( .B1(n11541), .B2(n19499), .A(n19476), .ZN(P2_U2939) );
  AOI22_X1 U22445 ( .A1(n19497), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19477) );
  OAI21_X1 U22446 ( .B1(n13514), .B2(n19499), .A(n19477), .ZN(P2_U2940) );
  AOI22_X1 U22447 ( .A1(n19497), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19478) );
  OAI21_X1 U22448 ( .B1(n13520), .B2(n19499), .A(n19478), .ZN(P2_U2941) );
  AOI22_X1 U22449 ( .A1(n19497), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19479) );
  OAI21_X1 U22450 ( .B1(n19480), .B2(n19499), .A(n19479), .ZN(P2_U2942) );
  AOI22_X1 U22451 ( .A1(n19497), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19481) );
  OAI21_X1 U22452 ( .B1(n13423), .B2(n19499), .A(n19481), .ZN(P2_U2943) );
  AOI22_X1 U22453 ( .A1(n19497), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19482) );
  OAI21_X1 U22454 ( .B1(n19483), .B2(n19499), .A(n19482), .ZN(P2_U2944) );
  AOI22_X1 U22455 ( .A1(n19497), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19484), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19485) );
  OAI21_X1 U22456 ( .B1(n19486), .B2(n19499), .A(n19485), .ZN(P2_U2945) );
  INV_X1 U22457 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19488) );
  AOI22_X1 U22458 ( .A1(n19497), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19487) );
  OAI21_X1 U22459 ( .B1(n19488), .B2(n19499), .A(n19487), .ZN(P2_U2946) );
  AOI22_X1 U22460 ( .A1(n19497), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19489) );
  OAI21_X1 U22461 ( .B1(n14276), .B2(n19499), .A(n19489), .ZN(P2_U2947) );
  INV_X1 U22462 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19491) );
  AOI22_X1 U22463 ( .A1(n19497), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19490) );
  OAI21_X1 U22464 ( .B1(n19491), .B2(n19499), .A(n19490), .ZN(P2_U2948) );
  AOI22_X1 U22465 ( .A1(n19497), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19492) );
  OAI21_X1 U22466 ( .B1(n19493), .B2(n19499), .A(n19492), .ZN(P2_U2949) );
  AOI22_X1 U22467 ( .A1(n19497), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19494) );
  OAI21_X1 U22468 ( .B1(n19495), .B2(n19499), .A(n19494), .ZN(P2_U2950) );
  AOI22_X1 U22469 ( .A1(n19497), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19496), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19498) );
  OAI21_X1 U22470 ( .B1(n13487), .B2(n19499), .A(n19498), .ZN(P2_U2951) );
  AOI22_X1 U22471 ( .A1(n19501), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19500), .ZN(n19508) );
  AOI222_X1 U22472 ( .A1(n19506), .A2(n19505), .B1(n19504), .B2(n19503), .C1(
        n10923), .C2(n19502), .ZN(n19507) );
  OAI211_X1 U22473 ( .C1(n19510), .C2(n19509), .A(n19508), .B(n19507), .ZN(
        P2_U3010) );
  NAND2_X1 U22474 ( .A1(n20175), .A2(n20182), .ZN(n19629) );
  INV_X1 U22475 ( .A(n19629), .ZN(n19632) );
  NAND2_X1 U22476 ( .A1(n19632), .A2(n20193), .ZN(n19577) );
  NOR2_X1 U22477 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19577), .ZN(
        n19566) );
  INV_X1 U22478 ( .A(n19566), .ZN(n19511) );
  AND2_X1 U22479 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19511), .ZN(n19512) );
  NAND2_X1 U22480 ( .A1(n19525), .A2(n19512), .ZN(n19518) );
  OAI21_X1 U22481 ( .B1(n20071), .B2(n19596), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19514) );
  NAND2_X1 U22482 ( .A1(n19514), .A2(n20170), .ZN(n19529) );
  AOI221_X1 U22483 ( .B1(n20067), .B2(n20195), .C1(n19529), .C2(n20195), .A(
        n19566), .ZN(n19515) );
  INV_X1 U22484 ( .A(n19515), .ZN(n19516) );
  AND2_X1 U22485 ( .A1(n20022), .A2(n19516), .ZN(n19517) );
  NOR2_X1 U22486 ( .A1(n20016), .A2(n20226), .ZN(n20183) );
  AOI22_X1 U22487 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19563), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19562), .ZN(n19917) );
  INV_X1 U22488 ( .A(n19917), .ZN(n20025) );
  NOR2_X2 U22489 ( .A1(n19522), .A2(n19564), .ZN(n20017) );
  AOI22_X1 U22490 ( .A1(n20025), .A2(n20071), .B1(n20017), .B2(n19566), .ZN(
        n19531) );
  NOR2_X1 U22491 ( .A1(n20067), .A2(n19566), .ZN(n19528) );
  INV_X1 U22492 ( .A(n19525), .ZN(n19526) );
  OAI21_X1 U22493 ( .B1(n19526), .B2(n19566), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19527) );
  AOI22_X1 U22494 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19563), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19562), .ZN(n20028) );
  AOI22_X1 U22495 ( .A1(n19524), .A2(n19568), .B1(n19596), .B2(n19914), .ZN(
        n19530) );
  OAI211_X1 U22496 ( .C1(n19539), .C2(n19532), .A(n19531), .B(n19530), .ZN(
        P2_U3048) );
  AOI22_X1 U22497 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19562), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19563), .ZN(n19994) );
  NOR2_X2 U22498 ( .A1(n9730), .A2(n19564), .ZN(n20029) );
  AOI22_X1 U22499 ( .A1(n20030), .A2(n20071), .B1(n20029), .B2(n19566), .ZN(
        n19536) );
  AOI22_X1 U22500 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19563), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19562), .ZN(n20033) );
  INV_X1 U22501 ( .A(n20033), .ZN(n19991) );
  AOI22_X1 U22502 ( .A1(n19534), .A2(n19568), .B1(n19596), .B2(n19991), .ZN(
        n19535) );
  OAI211_X1 U22503 ( .C1(n19539), .C2(n19537), .A(n19536), .B(n19535), .ZN(
        P2_U3049) );
  AOI22_X1 U22504 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19563), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19562), .ZN(n20039) );
  AOI22_X1 U22505 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19563), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19562), .ZN(n19923) );
  NOR2_X2 U22506 ( .A1(n19538), .A2(n19564), .ZN(n20034) );
  AOI22_X1 U22507 ( .A1(n20036), .A2(n20071), .B1(n20034), .B2(n19566), .ZN(
        n19542) );
  NOR2_X2 U22508 ( .A1(n19540), .A2(n19947), .ZN(n20035) );
  AOI22_X1 U22509 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19569), .B1(
        n20035), .B2(n19568), .ZN(n19541) );
  OAI211_X1 U22510 ( .C1(n20039), .C2(n19572), .A(n19542), .B(n19541), .ZN(
        P2_U3050) );
  AOI22_X1 U22511 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19563), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19562), .ZN(n19962) );
  AOI22_X1 U22512 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19562), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19563), .ZN(n20045) );
  INV_X1 U22513 ( .A(n20045), .ZN(n19959) );
  NOR2_X2 U22514 ( .A1(n19543), .A2(n19564), .ZN(n20040) );
  AOI22_X1 U22515 ( .A1(n19959), .A2(n20071), .B1(n20040), .B2(n19566), .ZN(
        n19546) );
  NOR2_X2 U22516 ( .A1(n19544), .A2(n19947), .ZN(n20041) );
  AOI22_X1 U22517 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19569), .B1(
        n20041), .B2(n19568), .ZN(n19545) );
  OAI211_X1 U22518 ( .C1(n19962), .C2(n19572), .A(n19546), .B(n19545), .ZN(
        P2_U3051) );
  AOI22_X1 U22519 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19562), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19563), .ZN(n20002) );
  AOI22_X1 U22520 ( .A1(n20071), .A2(n20048), .B1(n9656), .B2(n19566), .ZN(
        n19549) );
  NOR2_X2 U22521 ( .A1(n19547), .A2(n19947), .ZN(n20047) );
  AOI22_X1 U22522 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19569), .B1(
        n20047), .B2(n19568), .ZN(n19548) );
  OAI211_X1 U22523 ( .C1(n20051), .C2(n19572), .A(n19549), .B(n19548), .ZN(
        P2_U3052) );
  INV_X1 U22524 ( .A(n19563), .ZN(n19555) );
  INV_X1 U22525 ( .A(n19562), .ZN(n19557) );
  AOI22_X1 U22526 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19562), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19563), .ZN(n20057) );
  NOR2_X2 U22527 ( .A1(n19551), .A2(n19564), .ZN(n20052) );
  AOI22_X1 U22528 ( .A1(n19965), .A2(n20071), .B1(n20052), .B2(n19566), .ZN(
        n19554) );
  NOR2_X2 U22529 ( .A1(n19552), .A2(n19947), .ZN(n20053) );
  AOI22_X1 U22530 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19569), .B1(
        n20053), .B2(n19568), .ZN(n19553) );
  OAI211_X1 U22531 ( .C1(n19968), .C2(n19572), .A(n19554), .B(n19553), .ZN(
        P2_U3053) );
  AOI22_X1 U22532 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19563), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19562), .ZN(n20065) );
  NOR2_X2 U22533 ( .A1(n10203), .A2(n19564), .ZN(n20058) );
  AOI22_X1 U22534 ( .A1(n20060), .A2(n20071), .B1(n20058), .B2(n19566), .ZN(
        n19561) );
  NOR2_X2 U22535 ( .A1(n19559), .A2(n19947), .ZN(n20059) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19569), .B1(
        n20059), .B2(n19568), .ZN(n19560) );
  OAI211_X1 U22537 ( .C1(n20065), .C2(n19572), .A(n19561), .B(n19560), .ZN(
        P2_U3054) );
  AOI22_X1 U22538 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19562), .B1(
        BUF1_REG_23__SCAN_IN), .B2(n19563), .ZN(n19977) );
  AOI22_X1 U22539 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19563), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19562), .ZN(n20076) );
  INV_X1 U22540 ( .A(n20076), .ZN(n19972) );
  NOR2_X2 U22541 ( .A1(n19565), .A2(n19564), .ZN(n20066) );
  AOI22_X1 U22542 ( .A1(n19972), .A2(n20071), .B1(n20066), .B2(n19566), .ZN(
        n19571) );
  NOR2_X2 U22543 ( .A1(n19567), .A2(n19947), .ZN(n20068) );
  AOI22_X1 U22544 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19569), .B1(
        n20068), .B2(n19568), .ZN(n19570) );
  OAI211_X1 U22545 ( .C1(n19977), .C2(n19572), .A(n19571), .B(n19570), .ZN(
        P2_U3055) );
  INV_X1 U22546 ( .A(n19576), .ZN(n19574) );
  NAND2_X1 U22547 ( .A1(n20193), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19810) );
  NOR2_X1 U22548 ( .A1(n19810), .A2(n19629), .ZN(n19594) );
  OAI21_X1 U22549 ( .B1(n19574), .B2(n19594), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19575) );
  OAI21_X1 U22550 ( .B1(n19577), .B2(n20016), .A(n19575), .ZN(n19595) );
  AOI22_X1 U22551 ( .A1(n19595), .A2(n19524), .B1(n20017), .B2(n19594), .ZN(
        n19581) );
  AOI21_X1 U22552 ( .B1(n19576), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19579) );
  NAND2_X1 U22553 ( .A1(n20167), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19752) );
  OAI21_X1 U22554 ( .B1(n19752), .B2(n19811), .A(n19577), .ZN(n19578) );
  OAI211_X1 U22555 ( .C1(n19594), .C2(n19579), .A(n19578), .B(n20022), .ZN(
        n19597) );
  AOI22_X1 U22556 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19597), .B1(
        n19596), .B2(n20025), .ZN(n19580) );
  OAI211_X1 U22557 ( .C1(n20028), .C2(n19628), .A(n19581), .B(n19580), .ZN(
        P2_U3056) );
  AOI22_X1 U22558 ( .A1(n19595), .A2(n19534), .B1(n20029), .B2(n19594), .ZN(
        n19583) );
  AOI22_X1 U22559 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19597), .B1(
        n19596), .B2(n20030), .ZN(n19582) );
  OAI211_X1 U22560 ( .C1(n20033), .C2(n19628), .A(n19583), .B(n19582), .ZN(
        P2_U3057) );
  AOI22_X1 U22561 ( .A1(n19595), .A2(n20035), .B1(n20034), .B2(n19594), .ZN(
        n19585) );
  AOI22_X1 U22562 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19597), .B1(
        n19596), .B2(n20036), .ZN(n19584) );
  OAI211_X1 U22563 ( .C1(n20039), .C2(n19628), .A(n19585), .B(n19584), .ZN(
        P2_U3058) );
  AOI22_X1 U22564 ( .A1(n19595), .A2(n20041), .B1(n20040), .B2(n19594), .ZN(
        n19587) );
  AOI22_X1 U22565 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19597), .B1(
        n19596), .B2(n19959), .ZN(n19586) );
  OAI211_X1 U22566 ( .C1(n19962), .C2(n19628), .A(n19587), .B(n19586), .ZN(
        P2_U3059) );
  AOI22_X1 U22567 ( .A1(n19595), .A2(n20047), .B1(n9656), .B2(n19594), .ZN(
        n19589) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19597), .B1(
        n19596), .B2(n20048), .ZN(n19588) );
  OAI211_X1 U22569 ( .C1(n20051), .C2(n19628), .A(n19589), .B(n19588), .ZN(
        P2_U3060) );
  AOI22_X1 U22570 ( .A1(n19595), .A2(n20053), .B1(n20052), .B2(n19594), .ZN(
        n19591) );
  AOI22_X1 U22571 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19597), .B1(
        n19596), .B2(n19965), .ZN(n19590) );
  OAI211_X1 U22572 ( .C1(n19968), .C2(n19628), .A(n19591), .B(n19590), .ZN(
        P2_U3061) );
  AOI22_X1 U22573 ( .A1(n19595), .A2(n20059), .B1(n20058), .B2(n19594), .ZN(
        n19593) );
  AOI22_X1 U22574 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19597), .B1(
        n19596), .B2(n20060), .ZN(n19592) );
  OAI211_X1 U22575 ( .C1(n20065), .C2(n19628), .A(n19593), .B(n19592), .ZN(
        P2_U3062) );
  AOI22_X1 U22576 ( .A1(n19595), .A2(n20068), .B1(n20066), .B2(n19594), .ZN(
        n19599) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19597), .B1(
        n19596), .B2(n19972), .ZN(n19598) );
  OAI211_X1 U22578 ( .C1(n19977), .C2(n19628), .A(n19599), .B(n19598), .ZN(
        P2_U3063) );
  INV_X1 U22579 ( .A(n10492), .ZN(n19600) );
  NOR2_X1 U22580 ( .A1(n20193), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19839) );
  AND2_X1 U22581 ( .A1(n19839), .A2(n19632), .ZN(n19623) );
  OAI21_X1 U22582 ( .B1(n19600), .B2(n19623), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19601) );
  OR2_X1 U22583 ( .A1(n19841), .A2(n19629), .ZN(n19604) );
  NAND2_X1 U22584 ( .A1(n19601), .A2(n19604), .ZN(n19624) );
  AOI22_X1 U22585 ( .A1(n19624), .A2(n19524), .B1(n20017), .B2(n19623), .ZN(
        n19610) );
  INV_X1 U22586 ( .A(n19623), .ZN(n19602) );
  OAI21_X1 U22587 ( .B1(n10492), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19602), 
        .ZN(n19607) );
  INV_X1 U22588 ( .A(n19628), .ZN(n19603) );
  OAI21_X1 U22589 ( .B1(n19652), .B2(n19603), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19605) );
  NAND2_X1 U22590 ( .A1(n19605), .A2(n19604), .ZN(n19606) );
  MUX2_X1 U22591 ( .A(n19607), .B(n19606), .S(n20170), .Z(n19608) );
  NAND2_X1 U22592 ( .A1(n19608), .A2(n20022), .ZN(n19625) );
  AOI22_X1 U22593 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19625), .B1(
        n19652), .B2(n19914), .ZN(n19609) );
  OAI211_X1 U22594 ( .C1(n19917), .C2(n19628), .A(n19610), .B(n19609), .ZN(
        P2_U3064) );
  AOI22_X1 U22595 ( .A1(n19624), .A2(n19534), .B1(n20029), .B2(n19623), .ZN(
        n19612) );
  AOI22_X1 U22596 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19625), .B1(
        n19652), .B2(n19991), .ZN(n19611) );
  OAI211_X1 U22597 ( .C1(n19994), .C2(n19628), .A(n19612), .B(n19611), .ZN(
        P2_U3065) );
  AOI22_X1 U22598 ( .A1(n19624), .A2(n20035), .B1(n20034), .B2(n19623), .ZN(
        n19614) );
  INV_X1 U22599 ( .A(n20039), .ZN(n19920) );
  AOI22_X1 U22600 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19625), .B1(
        n19652), .B2(n19920), .ZN(n19613) );
  OAI211_X1 U22601 ( .C1(n19923), .C2(n19628), .A(n19614), .B(n19613), .ZN(
        P2_U3066) );
  AOI22_X1 U22602 ( .A1(n19624), .A2(n20041), .B1(n20040), .B2(n19623), .ZN(
        n19616) );
  INV_X1 U22603 ( .A(n19962), .ZN(n20042) );
  AOI22_X1 U22604 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19625), .B1(
        n19652), .B2(n20042), .ZN(n19615) );
  OAI211_X1 U22605 ( .C1(n20045), .C2(n19628), .A(n19616), .B(n19615), .ZN(
        P2_U3067) );
  AOI22_X1 U22606 ( .A1(n19624), .A2(n20047), .B1(n9656), .B2(n19623), .ZN(
        n19618) );
  INV_X1 U22607 ( .A(n20051), .ZN(n19999) );
  AOI22_X1 U22608 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19625), .B1(
        n19652), .B2(n19999), .ZN(n19617) );
  OAI211_X1 U22609 ( .C1(n20002), .C2(n19628), .A(n19618), .B(n19617), .ZN(
        P2_U3068) );
  AOI22_X1 U22610 ( .A1(n19624), .A2(n20053), .B1(n20052), .B2(n19623), .ZN(
        n19620) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19625), .B1(
        n19652), .B2(n20054), .ZN(n19619) );
  OAI211_X1 U22612 ( .C1(n20057), .C2(n19628), .A(n19620), .B(n19619), .ZN(
        P2_U3069) );
  AOI22_X1 U22613 ( .A1(n19624), .A2(n20059), .B1(n20058), .B2(n19623), .ZN(
        n19622) );
  INV_X1 U22614 ( .A(n20065), .ZN(n19930) );
  AOI22_X1 U22615 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19625), .B1(
        n19652), .B2(n19930), .ZN(n19621) );
  OAI211_X1 U22616 ( .C1(n19933), .C2(n19628), .A(n19622), .B(n19621), .ZN(
        P2_U3070) );
  AOI22_X1 U22617 ( .A1(n19624), .A2(n20068), .B1(n20066), .B2(n19623), .ZN(
        n19627) );
  INV_X1 U22618 ( .A(n19977), .ZN(n20070) );
  AOI22_X1 U22619 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19625), .B1(
        n19652), .B2(n20070), .ZN(n19626) );
  OAI211_X1 U22620 ( .C1(n20076), .C2(n19628), .A(n19627), .B(n19626), .ZN(
        P2_U3071) );
  NOR2_X1 U22621 ( .A1(n19872), .A2(n19629), .ZN(n19656) );
  AOI22_X1 U22622 ( .A1(n19914), .A2(n19687), .B1(n19656), .B2(n20017), .ZN(
        n19641) );
  AOI21_X1 U22623 ( .B1(n19630), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19634) );
  INV_X1 U22624 ( .A(n19752), .ZN(n19631) );
  AOI21_X1 U22625 ( .B1(n19631), .B2(n20164), .A(n20016), .ZN(n19635) );
  NAND2_X1 U22626 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19632), .ZN(
        n19638) );
  NAND2_X1 U22627 ( .A1(n19635), .A2(n19638), .ZN(n19633) );
  OAI211_X1 U22628 ( .C1(n19656), .C2(n19634), .A(n19633), .B(n20022), .ZN(
        n19658) );
  INV_X1 U22629 ( .A(n19635), .ZN(n19639) );
  OAI21_X1 U22630 ( .B1(n19636), .B2(n19656), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19637) );
  AOI22_X1 U22631 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19658), .B1(
        n19524), .B2(n19657), .ZN(n19640) );
  OAI211_X1 U22632 ( .C1(n19917), .C2(n19661), .A(n19641), .B(n19640), .ZN(
        P2_U3072) );
  AOI22_X1 U22633 ( .A1(n20030), .A2(n19652), .B1(n19656), .B2(n20029), .ZN(
        n19643) );
  AOI22_X1 U22634 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19658), .B1(
        n19534), .B2(n19657), .ZN(n19642) );
  OAI211_X1 U22635 ( .C1(n20033), .C2(n19655), .A(n19643), .B(n19642), .ZN(
        P2_U3073) );
  AOI22_X1 U22636 ( .A1(n20036), .A2(n19652), .B1(n19656), .B2(n20034), .ZN(
        n19645) );
  AOI22_X1 U22637 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19658), .B1(
        n20035), .B2(n19657), .ZN(n19644) );
  OAI211_X1 U22638 ( .C1(n20039), .C2(n19655), .A(n19645), .B(n19644), .ZN(
        P2_U3074) );
  AOI22_X1 U22639 ( .A1(n19959), .A2(n19652), .B1(n19656), .B2(n20040), .ZN(
        n19647) );
  AOI22_X1 U22640 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19658), .B1(
        n20041), .B2(n19657), .ZN(n19646) );
  OAI211_X1 U22641 ( .C1(n19962), .C2(n19655), .A(n19647), .B(n19646), .ZN(
        P2_U3075) );
  AOI22_X1 U22642 ( .A1(n19652), .A2(n20048), .B1(n19656), .B2(n9656), .ZN(
        n19649) );
  AOI22_X1 U22643 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19658), .B1(
        n20047), .B2(n19657), .ZN(n19648) );
  OAI211_X1 U22644 ( .C1(n20051), .C2(n19655), .A(n19649), .B(n19648), .ZN(
        P2_U3076) );
  AOI22_X1 U22645 ( .A1(n19965), .A2(n19652), .B1(n19656), .B2(n20052), .ZN(
        n19651) );
  AOI22_X1 U22646 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19658), .B1(
        n20053), .B2(n19657), .ZN(n19650) );
  OAI211_X1 U22647 ( .C1(n19968), .C2(n19655), .A(n19651), .B(n19650), .ZN(
        P2_U3077) );
  AOI22_X1 U22648 ( .A1(n20060), .A2(n19652), .B1(n19656), .B2(n20058), .ZN(
        n19654) );
  AOI22_X1 U22649 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19658), .B1(
        n20059), .B2(n19657), .ZN(n19653) );
  OAI211_X1 U22650 ( .C1(n20065), .C2(n19655), .A(n19654), .B(n19653), .ZN(
        P2_U3078) );
  AOI22_X1 U22651 ( .A1(n20070), .A2(n19687), .B1(n19656), .B2(n20066), .ZN(
        n19660) );
  AOI22_X1 U22652 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19658), .B1(
        n20068), .B2(n19657), .ZN(n19659) );
  OAI211_X1 U22653 ( .C1(n20076), .C2(n19661), .A(n19660), .B(n19659), .ZN(
        P2_U3079) );
  NOR2_X1 U22654 ( .A1(n19663), .A2(n19662), .ZN(n19906) );
  NAND2_X1 U22655 ( .A1(n19906), .A2(n20175), .ZN(n19669) );
  INV_X1 U22656 ( .A(n19664), .ZN(n19666) );
  NAND3_X1 U22657 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n20175), .A3(
        n20193), .ZN(n19697) );
  NOR2_X1 U22658 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19697), .ZN(
        n19685) );
  OAI21_X1 U22659 ( .B1(n19666), .B2(n19685), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19665) );
  OAI21_X1 U22660 ( .B1(n19669), .B2(n20016), .A(n19665), .ZN(n19686) );
  AOI22_X1 U22661 ( .A1(n19686), .A2(n19524), .B1(n20017), .B2(n19685), .ZN(
        n19672) );
  OAI21_X1 U22662 ( .B1(n19687), .B2(n19711), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19668) );
  AOI211_X1 U22663 ( .C1(n19666), .C2(n20195), .A(n19685), .B(n20170), .ZN(
        n19667) );
  AOI211_X1 U22664 ( .C1(n19669), .C2(n19668), .A(n19947), .B(n19667), .ZN(
        n19670) );
  AOI22_X1 U22665 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19688), .B1(
        n19687), .B2(n20025), .ZN(n19671) );
  OAI211_X1 U22666 ( .C1(n20028), .C2(n19718), .A(n19672), .B(n19671), .ZN(
        P2_U3080) );
  AOI22_X1 U22667 ( .A1(n19686), .A2(n19534), .B1(n20029), .B2(n19685), .ZN(
        n19674) );
  AOI22_X1 U22668 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19688), .B1(
        n19687), .B2(n20030), .ZN(n19673) );
  OAI211_X1 U22669 ( .C1(n20033), .C2(n19718), .A(n19674), .B(n19673), .ZN(
        P2_U3081) );
  AOI22_X1 U22670 ( .A1(n19686), .A2(n20035), .B1(n20034), .B2(n19685), .ZN(
        n19676) );
  AOI22_X1 U22671 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19688), .B1(
        n19687), .B2(n20036), .ZN(n19675) );
  OAI211_X1 U22672 ( .C1(n20039), .C2(n19718), .A(n19676), .B(n19675), .ZN(
        P2_U3082) );
  AOI22_X1 U22673 ( .A1(n19686), .A2(n20041), .B1(n20040), .B2(n19685), .ZN(
        n19678) );
  AOI22_X1 U22674 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19688), .B1(
        n19687), .B2(n19959), .ZN(n19677) );
  OAI211_X1 U22675 ( .C1(n19962), .C2(n19718), .A(n19678), .B(n19677), .ZN(
        P2_U3083) );
  AOI22_X1 U22676 ( .A1(n19686), .A2(n20047), .B1(n9656), .B2(n19685), .ZN(
        n19680) );
  AOI22_X1 U22677 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19688), .B1(
        n19687), .B2(n20048), .ZN(n19679) );
  OAI211_X1 U22678 ( .C1(n20051), .C2(n19718), .A(n19680), .B(n19679), .ZN(
        P2_U3084) );
  AOI22_X1 U22679 ( .A1(n19686), .A2(n20053), .B1(n20052), .B2(n19685), .ZN(
        n19682) );
  AOI22_X1 U22680 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19688), .B1(
        n19687), .B2(n19965), .ZN(n19681) );
  OAI211_X1 U22681 ( .C1(n19968), .C2(n19718), .A(n19682), .B(n19681), .ZN(
        P2_U3085) );
  AOI22_X1 U22682 ( .A1(n19686), .A2(n20059), .B1(n20058), .B2(n19685), .ZN(
        n19684) );
  AOI22_X1 U22683 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19688), .B1(
        n19687), .B2(n20060), .ZN(n19683) );
  OAI211_X1 U22684 ( .C1(n20065), .C2(n19718), .A(n19684), .B(n19683), .ZN(
        P2_U3086) );
  AOI22_X1 U22685 ( .A1(n19686), .A2(n20068), .B1(n20066), .B2(n19685), .ZN(
        n19690) );
  AOI22_X1 U22686 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19688), .B1(
        n19687), .B2(n19972), .ZN(n19689) );
  OAI211_X1 U22687 ( .C1(n19977), .C2(n19718), .A(n19690), .B(n19689), .ZN(
        P2_U3087) );
  INV_X1 U22688 ( .A(n19940), .ZN(n19951) );
  NOR2_X1 U22689 ( .A1(n20202), .A2(n19697), .ZN(n19725) );
  AOI22_X1 U22690 ( .A1(n19914), .A2(n19745), .B1(n19725), .B2(n20017), .ZN(
        n19700) );
  OAI21_X1 U22691 ( .B1(n19752), .B2(n19940), .A(n20170), .ZN(n19698) );
  INV_X1 U22692 ( .A(n19697), .ZN(n19694) );
  INV_X1 U22693 ( .A(n19725), .ZN(n19691) );
  OAI211_X1 U22694 ( .C1(n19692), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19691), 
        .B(n20016), .ZN(n19693) );
  OAI211_X1 U22695 ( .C1(n19698), .C2(n19694), .A(n20022), .B(n19693), .ZN(
        n19715) );
  OAI21_X1 U22696 ( .B1(n19695), .B2(n19725), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19696) );
  OAI21_X1 U22697 ( .B1(n19698), .B2(n19697), .A(n19696), .ZN(n19714) );
  AOI22_X1 U22698 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19715), .B1(
        n19524), .B2(n19714), .ZN(n19699) );
  OAI211_X1 U22699 ( .C1(n19917), .C2(n19718), .A(n19700), .B(n19699), .ZN(
        P2_U3088) );
  AOI22_X1 U22700 ( .A1(n20030), .A2(n19711), .B1(n20029), .B2(n19725), .ZN(
        n19702) );
  AOI22_X1 U22701 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19715), .B1(
        n19534), .B2(n19714), .ZN(n19701) );
  OAI211_X1 U22702 ( .C1(n20033), .C2(n19742), .A(n19702), .B(n19701), .ZN(
        P2_U3089) );
  AOI22_X1 U22703 ( .A1(n19920), .A2(n19745), .B1(n19725), .B2(n20034), .ZN(
        n19704) );
  AOI22_X1 U22704 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19715), .B1(
        n20035), .B2(n19714), .ZN(n19703) );
  OAI211_X1 U22705 ( .C1(n19923), .C2(n19718), .A(n19704), .B(n19703), .ZN(
        P2_U3090) );
  AOI22_X1 U22706 ( .A1(n19959), .A2(n19711), .B1(n19725), .B2(n20040), .ZN(
        n19706) );
  AOI22_X1 U22707 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19715), .B1(
        n20041), .B2(n19714), .ZN(n19705) );
  OAI211_X1 U22708 ( .C1(n19962), .C2(n19742), .A(n19706), .B(n19705), .ZN(
        P2_U3091) );
  AOI22_X1 U22709 ( .A1(n19999), .A2(n19745), .B1(n19725), .B2(n9656), .ZN(
        n19708) );
  AOI22_X1 U22710 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19715), .B1(
        n20047), .B2(n19714), .ZN(n19707) );
  OAI211_X1 U22711 ( .C1(n20002), .C2(n19718), .A(n19708), .B(n19707), .ZN(
        P2_U3092) );
  AOI22_X1 U22712 ( .A1(n20054), .A2(n19745), .B1(n19725), .B2(n20052), .ZN(
        n19710) );
  AOI22_X1 U22713 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19715), .B1(
        n20053), .B2(n19714), .ZN(n19709) );
  OAI211_X1 U22714 ( .C1(n20057), .C2(n19718), .A(n19710), .B(n19709), .ZN(
        P2_U3093) );
  AOI22_X1 U22715 ( .A1(n20060), .A2(n19711), .B1(n19725), .B2(n20058), .ZN(
        n19713) );
  AOI22_X1 U22716 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19715), .B1(
        n20059), .B2(n19714), .ZN(n19712) );
  OAI211_X1 U22717 ( .C1(n20065), .C2(n19742), .A(n19713), .B(n19712), .ZN(
        P2_U3094) );
  AOI22_X1 U22718 ( .A1(n20070), .A2(n19745), .B1(n19725), .B2(n20066), .ZN(
        n19717) );
  AOI22_X1 U22719 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19715), .B1(
        n20068), .B2(n19714), .ZN(n19716) );
  OAI211_X1 U22720 ( .C1(n20076), .C2(n19718), .A(n19717), .B(n19716), .ZN(
        P2_U3095) );
  NAND2_X1 U22721 ( .A1(n20175), .A2(n19979), .ZN(n19751) );
  NOR2_X1 U22722 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19751), .ZN(
        n19743) );
  NOR2_X1 U22723 ( .A1(n19725), .A2(n19743), .ZN(n19720) );
  OR2_X1 U22724 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19720), .ZN(n19723) );
  INV_X1 U22725 ( .A(n19721), .ZN(n19722) );
  NOR3_X1 U22726 ( .A1(n19722), .A2(n19743), .A3(n19942), .ZN(n19726) );
  AOI21_X1 U22727 ( .B1(n19942), .B2(n19723), .A(n19726), .ZN(n19744) );
  AOI22_X1 U22728 ( .A1(n19744), .A2(n19524), .B1(n20017), .B2(n19743), .ZN(
        n19729) );
  AOI21_X1 U22729 ( .B1(n19742), .B2(n19778), .A(n20226), .ZN(n19724) );
  AOI221_X1 U22730 ( .B1(n20195), .B2(n19725), .C1(n20195), .C2(n19724), .A(
        n19743), .ZN(n19727) );
  AOI22_X1 U22731 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n20025), .ZN(n19728) );
  OAI211_X1 U22732 ( .C1(n20028), .C2(n19778), .A(n19729), .B(n19728), .ZN(
        P2_U3096) );
  AOI22_X1 U22733 ( .A1(n19744), .A2(n19534), .B1(n20029), .B2(n19743), .ZN(
        n19731) );
  AOI22_X1 U22734 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n20030), .ZN(n19730) );
  OAI211_X1 U22735 ( .C1(n20033), .C2(n19778), .A(n19731), .B(n19730), .ZN(
        P2_U3097) );
  AOI22_X1 U22736 ( .A1(n19744), .A2(n20035), .B1(n20034), .B2(n19743), .ZN(
        n19733) );
  AOI22_X1 U22737 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19746), .B1(
        n19767), .B2(n19920), .ZN(n19732) );
  OAI211_X1 U22738 ( .C1(n19923), .C2(n19742), .A(n19733), .B(n19732), .ZN(
        P2_U3098) );
  AOI22_X1 U22739 ( .A1(n19744), .A2(n20041), .B1(n20040), .B2(n19743), .ZN(
        n19735) );
  AOI22_X1 U22740 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19746), .B1(
        n19767), .B2(n20042), .ZN(n19734) );
  OAI211_X1 U22741 ( .C1(n20045), .C2(n19742), .A(n19735), .B(n19734), .ZN(
        P2_U3099) );
  AOI22_X1 U22742 ( .A1(n19744), .A2(n20047), .B1(n9656), .B2(n19743), .ZN(
        n19737) );
  AOI22_X1 U22743 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n20048), .ZN(n19736) );
  OAI211_X1 U22744 ( .C1(n20051), .C2(n19778), .A(n19737), .B(n19736), .ZN(
        P2_U3100) );
  AOI22_X1 U22745 ( .A1(n19744), .A2(n20053), .B1(n20052), .B2(n19743), .ZN(
        n19739) );
  AOI22_X1 U22746 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19746), .B1(
        n19767), .B2(n20054), .ZN(n19738) );
  OAI211_X1 U22747 ( .C1(n20057), .C2(n19742), .A(n19739), .B(n19738), .ZN(
        P2_U3101) );
  AOI22_X1 U22748 ( .A1(n19744), .A2(n20059), .B1(n20058), .B2(n19743), .ZN(
        n19741) );
  AOI22_X1 U22749 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19746), .B1(
        n19767), .B2(n19930), .ZN(n19740) );
  OAI211_X1 U22750 ( .C1(n19933), .C2(n19742), .A(n19741), .B(n19740), .ZN(
        P2_U3102) );
  AOI22_X1 U22751 ( .A1(n19744), .A2(n20068), .B1(n20066), .B2(n19743), .ZN(
        n19748) );
  AOI22_X1 U22752 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19746), .B1(
        n19745), .B2(n19972), .ZN(n19747) );
  OAI211_X1 U22753 ( .C1(n19977), .C2(n19778), .A(n19748), .B(n19747), .ZN(
        P2_U3103) );
  NOR2_X1 U22754 ( .A1(n20202), .A2(n19751), .ZN(n19785) );
  OR3_X1 U22755 ( .A1(n19749), .A2(n19785), .A3(n19942), .ZN(n19753) );
  INV_X1 U22756 ( .A(n19753), .ZN(n19750) );
  AOI211_X2 U22757 ( .C1(n19751), .C2(n19942), .A(n20079), .B(n19750), .ZN(
        n19774) );
  AOI22_X1 U22758 ( .A1(n19774), .A2(n19524), .B1(n20017), .B2(n19785), .ZN(
        n19760) );
  INV_X1 U22759 ( .A(n19751), .ZN(n19756) );
  NOR2_X1 U22760 ( .A1(n19752), .A2(n20020), .ZN(n20169) );
  OAI211_X1 U22761 ( .C1(n20195), .C2(n19785), .A(n19753), .B(n20022), .ZN(
        n19754) );
  INV_X1 U22762 ( .A(n19754), .ZN(n19755) );
  OAI21_X1 U22763 ( .B1(n19756), .B2(n20169), .A(n19755), .ZN(n19775) );
  INV_X1 U22764 ( .A(n20020), .ZN(n19757) );
  AOI22_X1 U22765 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19775), .B1(
        n19805), .B2(n19914), .ZN(n19759) );
  OAI211_X1 U22766 ( .C1(n19917), .C2(n19778), .A(n19760), .B(n19759), .ZN(
        P2_U3104) );
  AOI22_X1 U22767 ( .A1(n19774), .A2(n19534), .B1(n20029), .B2(n19785), .ZN(
        n19762) );
  AOI22_X1 U22768 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19775), .B1(
        n19805), .B2(n19991), .ZN(n19761) );
  OAI211_X1 U22769 ( .C1(n19994), .C2(n19778), .A(n19762), .B(n19761), .ZN(
        P2_U3105) );
  AOI22_X1 U22770 ( .A1(n19774), .A2(n20035), .B1(n20034), .B2(n19785), .ZN(
        n19764) );
  AOI22_X1 U22771 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19775), .B1(
        n19805), .B2(n19920), .ZN(n19763) );
  OAI211_X1 U22772 ( .C1(n19923), .C2(n19778), .A(n19764), .B(n19763), .ZN(
        P2_U3106) );
  AOI22_X1 U22773 ( .A1(n19774), .A2(n20041), .B1(n20040), .B2(n19785), .ZN(
        n19766) );
  AOI22_X1 U22774 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19775), .B1(
        n19767), .B2(n19959), .ZN(n19765) );
  OAI211_X1 U22775 ( .C1(n19962), .C2(n19803), .A(n19766), .B(n19765), .ZN(
        P2_U3107) );
  AOI22_X1 U22776 ( .A1(n19774), .A2(n20047), .B1(n9656), .B2(n19785), .ZN(
        n19769) );
  AOI22_X1 U22777 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19775), .B1(
        n19767), .B2(n20048), .ZN(n19768) );
  OAI211_X1 U22778 ( .C1(n20051), .C2(n19803), .A(n19769), .B(n19768), .ZN(
        P2_U3108) );
  AOI22_X1 U22779 ( .A1(n19774), .A2(n20053), .B1(n20052), .B2(n19785), .ZN(
        n19771) );
  AOI22_X1 U22780 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19775), .B1(
        n19805), .B2(n20054), .ZN(n19770) );
  OAI211_X1 U22781 ( .C1(n20057), .C2(n19778), .A(n19771), .B(n19770), .ZN(
        P2_U3109) );
  AOI22_X1 U22782 ( .A1(n19774), .A2(n20059), .B1(n20058), .B2(n19785), .ZN(
        n19773) );
  AOI22_X1 U22783 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19775), .B1(
        n19805), .B2(n19930), .ZN(n19772) );
  OAI211_X1 U22784 ( .C1(n19933), .C2(n19778), .A(n19773), .B(n19772), .ZN(
        P2_U3110) );
  AOI22_X1 U22785 ( .A1(n19774), .A2(n20068), .B1(n20066), .B2(n19785), .ZN(
        n19777) );
  AOI22_X1 U22786 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19775), .B1(
        n19805), .B2(n20070), .ZN(n19776) );
  OAI211_X1 U22787 ( .C1(n20076), .C2(n19778), .A(n19777), .B(n19776), .ZN(
        P2_U3111) );
  NAND2_X1 U22788 ( .A1(n20182), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19877) );
  INV_X1 U22789 ( .A(n19877), .ZN(n19873) );
  NAND2_X1 U22790 ( .A1(n19873), .A2(n20193), .ZN(n19817) );
  NOR2_X1 U22791 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19817), .ZN(
        n19804) );
  AOI22_X1 U22792 ( .A1(n19914), .A2(n19829), .B1(n20017), .B2(n19804), .ZN(
        n19790) );
  AOI21_X1 U22793 ( .B1(n19803), .B2(n19838), .A(n20226), .ZN(n19780) );
  NOR2_X1 U22794 ( .A1(n19780), .A2(n20016), .ZN(n19784) );
  INV_X1 U22795 ( .A(n19785), .ZN(n19782) );
  INV_X1 U22796 ( .A(n10487), .ZN(n19786) );
  AOI21_X1 U22797 ( .B1(n19786), .B2(n20195), .A(n20170), .ZN(n19781) );
  AOI21_X1 U22798 ( .B1(n19784), .B2(n19782), .A(n19781), .ZN(n19783) );
  OAI21_X1 U22799 ( .B1(n19804), .B2(n19783), .A(n20022), .ZN(n19807) );
  OAI21_X1 U22800 ( .B1(n19804), .B2(n19785), .A(n19784), .ZN(n19788) );
  OAI21_X1 U22801 ( .B1(n19786), .B2(n19804), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19787) );
  AOI22_X1 U22802 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19807), .B1(
        n19524), .B2(n19806), .ZN(n19789) );
  OAI211_X1 U22803 ( .C1(n19917), .C2(n19803), .A(n19790), .B(n19789), .ZN(
        P2_U3112) );
  AOI22_X1 U22804 ( .A1(n19991), .A2(n19829), .B1(n20029), .B2(n19804), .ZN(
        n19792) );
  AOI22_X1 U22805 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19807), .B1(
        n19534), .B2(n19806), .ZN(n19791) );
  OAI211_X1 U22806 ( .C1(n19994), .C2(n19803), .A(n19792), .B(n19791), .ZN(
        P2_U3113) );
  AOI22_X1 U22807 ( .A1(n20036), .A2(n19805), .B1(n20034), .B2(n19804), .ZN(
        n19794) );
  AOI22_X1 U22808 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19807), .B1(
        n20035), .B2(n19806), .ZN(n19793) );
  OAI211_X1 U22809 ( .C1(n20039), .C2(n19838), .A(n19794), .B(n19793), .ZN(
        P2_U3114) );
  AOI22_X1 U22810 ( .A1(n20042), .A2(n19829), .B1(n20040), .B2(n19804), .ZN(
        n19796) );
  AOI22_X1 U22811 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19807), .B1(
        n20041), .B2(n19806), .ZN(n19795) );
  OAI211_X1 U22812 ( .C1(n20045), .C2(n19803), .A(n19796), .B(n19795), .ZN(
        P2_U3115) );
  AOI22_X1 U22813 ( .A1(n19805), .A2(n20048), .B1(n9656), .B2(n19804), .ZN(
        n19798) );
  AOI22_X1 U22814 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19807), .B1(
        n20047), .B2(n19806), .ZN(n19797) );
  OAI211_X1 U22815 ( .C1(n20051), .C2(n19838), .A(n19798), .B(n19797), .ZN(
        P2_U3116) );
  AOI22_X1 U22816 ( .A1(n19965), .A2(n19805), .B1(n20052), .B2(n19804), .ZN(
        n19800) );
  AOI22_X1 U22817 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19807), .B1(
        n20053), .B2(n19806), .ZN(n19799) );
  OAI211_X1 U22818 ( .C1(n19968), .C2(n19838), .A(n19800), .B(n19799), .ZN(
        P2_U3117) );
  AOI22_X1 U22819 ( .A1(n19930), .A2(n19829), .B1(n20058), .B2(n19804), .ZN(
        n19802) );
  AOI22_X1 U22820 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19807), .B1(
        n20059), .B2(n19806), .ZN(n19801) );
  OAI211_X1 U22821 ( .C1(n19933), .C2(n19803), .A(n19802), .B(n19801), .ZN(
        P2_U3118) );
  AOI22_X1 U22822 ( .A1(n19972), .A2(n19805), .B1(n20066), .B2(n19804), .ZN(
        n19809) );
  AOI22_X1 U22823 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19807), .B1(
        n20068), .B2(n19806), .ZN(n19808) );
  OAI211_X1 U22824 ( .C1(n19977), .C2(n19838), .A(n19809), .B(n19808), .ZN(
        P2_U3119) );
  NOR2_X1 U22825 ( .A1(n19810), .A2(n19877), .ZN(n19842) );
  AOI22_X1 U22826 ( .A1(n19914), .A2(n19867), .B1(n20017), .B2(n19842), .ZN(
        n19820) );
  OR2_X1 U22827 ( .A1(n20167), .A2(n20226), .ZN(n20021) );
  OAI21_X1 U22828 ( .B1(n20021), .B2(n19811), .A(n20170), .ZN(n19818) );
  INV_X1 U22829 ( .A(n19817), .ZN(n19812) );
  NOR2_X1 U22830 ( .A1(n19818), .A2(n19812), .ZN(n19813) );
  AOI211_X1 U22831 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n10480), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19813), .ZN(n19814) );
  OAI21_X1 U22832 ( .B1(n19842), .B2(n19814), .A(n20022), .ZN(n19835) );
  INV_X1 U22833 ( .A(n10480), .ZN(n19815) );
  OAI21_X1 U22834 ( .B1(n19815), .B2(n19842), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19816) );
  AOI22_X1 U22835 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19835), .B1(
        n19524), .B2(n19834), .ZN(n19819) );
  OAI211_X1 U22836 ( .C1(n19917), .C2(n19838), .A(n19820), .B(n19819), .ZN(
        P2_U3120) );
  AOI22_X1 U22837 ( .A1(n19991), .A2(n19867), .B1(n20029), .B2(n19842), .ZN(
        n19822) );
  AOI22_X1 U22838 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19835), .B1(
        n19534), .B2(n19834), .ZN(n19821) );
  OAI211_X1 U22839 ( .C1(n19994), .C2(n19838), .A(n19822), .B(n19821), .ZN(
        P2_U3121) );
  AOI22_X1 U22840 ( .A1(n19920), .A2(n19867), .B1(n20034), .B2(n19842), .ZN(
        n19824) );
  AOI22_X1 U22841 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19835), .B1(
        n20035), .B2(n19834), .ZN(n19823) );
  OAI211_X1 U22842 ( .C1(n19923), .C2(n19838), .A(n19824), .B(n19823), .ZN(
        P2_U3122) );
  AOI22_X1 U22843 ( .A1(n19959), .A2(n19829), .B1(n20040), .B2(n19842), .ZN(
        n19826) );
  AOI22_X1 U22844 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19835), .B1(
        n20041), .B2(n19834), .ZN(n19825) );
  OAI211_X1 U22845 ( .C1(n19962), .C2(n19864), .A(n19826), .B(n19825), .ZN(
        P2_U3123) );
  AOI22_X1 U22846 ( .A1(n19829), .A2(n20048), .B1(n9656), .B2(n19842), .ZN(
        n19828) );
  AOI22_X1 U22847 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19835), .B1(
        n20047), .B2(n19834), .ZN(n19827) );
  OAI211_X1 U22848 ( .C1(n20051), .C2(n19864), .A(n19828), .B(n19827), .ZN(
        P2_U3124) );
  AOI22_X1 U22849 ( .A1(n19965), .A2(n19829), .B1(n20052), .B2(n19842), .ZN(
        n19831) );
  AOI22_X1 U22850 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19835), .B1(
        n20053), .B2(n19834), .ZN(n19830) );
  OAI211_X1 U22851 ( .C1(n19968), .C2(n19864), .A(n19831), .B(n19830), .ZN(
        P2_U3125) );
  AOI22_X1 U22852 ( .A1(n19930), .A2(n19867), .B1(n20058), .B2(n19842), .ZN(
        n19833) );
  AOI22_X1 U22853 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19835), .B1(
        n20059), .B2(n19834), .ZN(n19832) );
  OAI211_X1 U22854 ( .C1(n19933), .C2(n19838), .A(n19833), .B(n19832), .ZN(
        P2_U3126) );
  AOI22_X1 U22855 ( .A1(n20070), .A2(n19867), .B1(n20066), .B2(n19842), .ZN(
        n19837) );
  AOI22_X1 U22856 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19835), .B1(
        n20068), .B2(n19834), .ZN(n19836) );
  OAI211_X1 U22857 ( .C1(n20076), .C2(n19838), .A(n19837), .B(n19836), .ZN(
        P2_U3127) );
  INV_X1 U22858 ( .A(n9750), .ZN(n19845) );
  NAND2_X1 U22859 ( .A1(n19839), .A2(n19873), .ZN(n19846) );
  INV_X1 U22860 ( .A(n19846), .ZN(n19865) );
  OAI21_X1 U22861 ( .B1(n19845), .B2(n19865), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19840) );
  OAI21_X1 U22862 ( .B1(n19877), .B2(n19841), .A(n19840), .ZN(n19866) );
  AOI22_X1 U22863 ( .A1(n19866), .A2(n19524), .B1(n20017), .B2(n19865), .ZN(
        n19851) );
  OAI21_X1 U22864 ( .B1(n19867), .B2(n19902), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19844) );
  INV_X1 U22865 ( .A(n19842), .ZN(n19843) );
  AOI21_X1 U22866 ( .B1(n19844), .B2(n19843), .A(n20016), .ZN(n19849) );
  NAND3_X1 U22867 ( .A1(n19845), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n20195), 
        .ZN(n19847) );
  NAND2_X1 U22868 ( .A1(n19847), .A2(n19846), .ZN(n19848) );
  OAI21_X1 U22869 ( .B1(n19849), .B2(n19848), .A(n20022), .ZN(n19868) );
  AOI22_X1 U22870 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19868), .B1(
        n19902), .B2(n19914), .ZN(n19850) );
  OAI211_X1 U22871 ( .C1(n19917), .C2(n19864), .A(n19851), .B(n19850), .ZN(
        P2_U3128) );
  AOI22_X1 U22872 ( .A1(n19866), .A2(n19534), .B1(n20029), .B2(n19865), .ZN(
        n19853) );
  AOI22_X1 U22873 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19868), .B1(
        n19902), .B2(n19991), .ZN(n19852) );
  OAI211_X1 U22874 ( .C1(n19994), .C2(n19864), .A(n19853), .B(n19852), .ZN(
        P2_U3129) );
  AOI22_X1 U22875 ( .A1(n19866), .A2(n20035), .B1(n20034), .B2(n19865), .ZN(
        n19855) );
  AOI22_X1 U22876 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19868), .B1(
        n19867), .B2(n20036), .ZN(n19854) );
  OAI211_X1 U22877 ( .C1(n20039), .C2(n19895), .A(n19855), .B(n19854), .ZN(
        P2_U3130) );
  AOI22_X1 U22878 ( .A1(n19866), .A2(n20041), .B1(n20040), .B2(n19865), .ZN(
        n19857) );
  AOI22_X1 U22879 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19868), .B1(
        n19867), .B2(n19959), .ZN(n19856) );
  OAI211_X1 U22880 ( .C1(n19962), .C2(n19895), .A(n19857), .B(n19856), .ZN(
        P2_U3131) );
  AOI22_X1 U22881 ( .A1(n19866), .A2(n20047), .B1(n9656), .B2(n19865), .ZN(
        n19859) );
  AOI22_X1 U22882 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19868), .B1(
        n19867), .B2(n20048), .ZN(n19858) );
  OAI211_X1 U22883 ( .C1(n20051), .C2(n19895), .A(n19859), .B(n19858), .ZN(
        P2_U3132) );
  AOI22_X1 U22884 ( .A1(n19866), .A2(n20053), .B1(n20052), .B2(n19865), .ZN(
        n19861) );
  AOI22_X1 U22885 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19868), .B1(
        n19867), .B2(n19965), .ZN(n19860) );
  OAI211_X1 U22886 ( .C1(n19968), .C2(n19895), .A(n19861), .B(n19860), .ZN(
        P2_U3133) );
  AOI22_X1 U22887 ( .A1(n19866), .A2(n20059), .B1(n20058), .B2(n19865), .ZN(
        n19863) );
  AOI22_X1 U22888 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19868), .B1(
        n19902), .B2(n19930), .ZN(n19862) );
  OAI211_X1 U22889 ( .C1(n19933), .C2(n19864), .A(n19863), .B(n19862), .ZN(
        P2_U3134) );
  AOI22_X1 U22890 ( .A1(n19866), .A2(n20068), .B1(n20066), .B2(n19865), .ZN(
        n19870) );
  AOI22_X1 U22891 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19868), .B1(
        n19867), .B2(n19972), .ZN(n19869) );
  OAI211_X1 U22892 ( .C1(n19977), .C2(n19895), .A(n19870), .B(n19869), .ZN(
        P2_U3135) );
  INV_X1 U22893 ( .A(n19872), .ZN(n19874) );
  NAND2_X1 U22894 ( .A1(n19874), .A2(n19873), .ZN(n19880) );
  AND2_X1 U22895 ( .A1(n19880), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19875) );
  NAND2_X1 U22896 ( .A1(n19876), .A2(n19875), .ZN(n19881) );
  NOR2_X1 U22897 ( .A1(n20193), .A2(n19877), .ZN(n19884) );
  INV_X1 U22898 ( .A(n19884), .ZN(n19878) );
  OAI21_X1 U22899 ( .B1(n19878), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19942), 
        .ZN(n19879) );
  AND2_X1 U22900 ( .A1(n19881), .A2(n19879), .ZN(n19901) );
  INV_X1 U22901 ( .A(n19880), .ZN(n19900) );
  AOI22_X1 U22902 ( .A1(n19901), .A2(n19524), .B1(n20017), .B2(n19900), .ZN(
        n19886) );
  INV_X1 U22903 ( .A(n20021), .ZN(n19950) );
  OAI211_X1 U22904 ( .C1(n19900), .C2(n20195), .A(n19881), .B(n20022), .ZN(
        n19882) );
  INV_X1 U22905 ( .A(n19882), .ZN(n19883) );
  OAI221_X1 U22906 ( .B1(n19884), .B2(n20164), .C1(n19884), .C2(n19950), .A(
        n19883), .ZN(n19903) );
  AOI22_X1 U22907 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19903), .B1(
        n19902), .B2(n20025), .ZN(n19885) );
  OAI211_X1 U22908 ( .C1(n20028), .C2(n19939), .A(n19886), .B(n19885), .ZN(
        P2_U3136) );
  AOI22_X1 U22909 ( .A1(n19901), .A2(n19534), .B1(n20029), .B2(n19900), .ZN(
        n19888) );
  AOI22_X1 U22910 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19903), .B1(
        n19902), .B2(n20030), .ZN(n19887) );
  OAI211_X1 U22911 ( .C1(n20033), .C2(n19939), .A(n19888), .B(n19887), .ZN(
        P2_U3137) );
  AOI22_X1 U22912 ( .A1(n19901), .A2(n20035), .B1(n20034), .B2(n19900), .ZN(
        n19890) );
  AOI22_X1 U22913 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19903), .B1(
        n19909), .B2(n19920), .ZN(n19889) );
  OAI211_X1 U22914 ( .C1(n19923), .C2(n19895), .A(n19890), .B(n19889), .ZN(
        P2_U3138) );
  AOI22_X1 U22915 ( .A1(n19901), .A2(n20041), .B1(n20040), .B2(n19900), .ZN(
        n19892) );
  AOI22_X1 U22916 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19903), .B1(
        n19909), .B2(n20042), .ZN(n19891) );
  OAI211_X1 U22917 ( .C1(n20045), .C2(n19895), .A(n19892), .B(n19891), .ZN(
        P2_U3139) );
  AOI22_X1 U22918 ( .A1(n19901), .A2(n20047), .B1(n9656), .B2(n19900), .ZN(
        n19894) );
  AOI22_X1 U22919 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19903), .B1(
        n19909), .B2(n19999), .ZN(n19893) );
  OAI211_X1 U22920 ( .C1(n20002), .C2(n19895), .A(n19894), .B(n19893), .ZN(
        P2_U3140) );
  AOI22_X1 U22921 ( .A1(n19901), .A2(n20053), .B1(n20052), .B2(n19900), .ZN(
        n19897) );
  AOI22_X1 U22922 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19903), .B1(
        n19902), .B2(n19965), .ZN(n19896) );
  OAI211_X1 U22923 ( .C1(n19968), .C2(n19939), .A(n19897), .B(n19896), .ZN(
        P2_U3141) );
  AOI22_X1 U22924 ( .A1(n19901), .A2(n20059), .B1(n20058), .B2(n19900), .ZN(
        n19899) );
  AOI22_X1 U22925 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19903), .B1(
        n19902), .B2(n20060), .ZN(n19898) );
  OAI211_X1 U22926 ( .C1(n20065), .C2(n19939), .A(n19899), .B(n19898), .ZN(
        P2_U3142) );
  AOI22_X1 U22927 ( .A1(n19901), .A2(n20068), .B1(n20066), .B2(n19900), .ZN(
        n19905) );
  AOI22_X1 U22928 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19903), .B1(
        n19902), .B2(n19972), .ZN(n19904) );
  OAI211_X1 U22929 ( .C1(n19977), .C2(n19939), .A(n19905), .B(n19904), .ZN(
        P2_U3143) );
  NAND2_X1 U22930 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19906), .ZN(
        n19911) );
  OR2_X1 U22931 ( .A1(n19911), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19908) );
  INV_X1 U22932 ( .A(n10486), .ZN(n19907) );
  NAND3_X1 U22933 ( .A1(n20193), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19944) );
  NOR2_X1 U22934 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19944), .ZN(
        n19934) );
  NOR3_X1 U22935 ( .A1(n19907), .A2(n19934), .A3(n19942), .ZN(n19910) );
  AOI21_X1 U22936 ( .B1(n19942), .B2(n19908), .A(n19910), .ZN(n19935) );
  AOI22_X1 U22937 ( .A1(n19935), .A2(n19524), .B1(n20017), .B2(n19934), .ZN(
        n19916) );
  OAI21_X1 U22938 ( .B1(n19909), .B2(n19973), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19912) );
  AOI211_X1 U22939 ( .C1(n19912), .C2(n19911), .A(n19947), .B(n19910), .ZN(
        n19913) );
  AOI22_X1 U22940 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19936), .B1(
        n19973), .B2(n19914), .ZN(n19915) );
  OAI211_X1 U22941 ( .C1(n19917), .C2(n19939), .A(n19916), .B(n19915), .ZN(
        P2_U3144) );
  AOI22_X1 U22942 ( .A1(n19935), .A2(n19534), .B1(n20029), .B2(n19934), .ZN(
        n19919) );
  AOI22_X1 U22943 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19936), .B1(
        n19973), .B2(n19991), .ZN(n19918) );
  OAI211_X1 U22944 ( .C1(n19994), .C2(n19939), .A(n19919), .B(n19918), .ZN(
        P2_U3145) );
  AOI22_X1 U22945 ( .A1(n19935), .A2(n20035), .B1(n20034), .B2(n19934), .ZN(
        n19922) );
  AOI22_X1 U22946 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19936), .B1(
        n19973), .B2(n19920), .ZN(n19921) );
  OAI211_X1 U22947 ( .C1(n19923), .C2(n19939), .A(n19922), .B(n19921), .ZN(
        P2_U3146) );
  AOI22_X1 U22948 ( .A1(n19935), .A2(n20041), .B1(n20040), .B2(n19934), .ZN(
        n19925) );
  AOI22_X1 U22949 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19936), .B1(
        n19973), .B2(n20042), .ZN(n19924) );
  OAI211_X1 U22950 ( .C1(n20045), .C2(n19939), .A(n19925), .B(n19924), .ZN(
        P2_U3147) );
  AOI22_X1 U22951 ( .A1(n19935), .A2(n20047), .B1(n9656), .B2(n19934), .ZN(
        n19927) );
  AOI22_X1 U22952 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19936), .B1(
        n19973), .B2(n19999), .ZN(n19926) );
  OAI211_X1 U22953 ( .C1(n20002), .C2(n19939), .A(n19927), .B(n19926), .ZN(
        P2_U3148) );
  AOI22_X1 U22954 ( .A1(n19935), .A2(n20053), .B1(n20052), .B2(n19934), .ZN(
        n19929) );
  AOI22_X1 U22955 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19936), .B1(
        n19973), .B2(n20054), .ZN(n19928) );
  OAI211_X1 U22956 ( .C1(n20057), .C2(n19939), .A(n19929), .B(n19928), .ZN(
        P2_U3149) );
  AOI22_X1 U22957 ( .A1(n19935), .A2(n20059), .B1(n20058), .B2(n19934), .ZN(
        n19932) );
  AOI22_X1 U22958 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19936), .B1(
        n19973), .B2(n19930), .ZN(n19931) );
  OAI211_X1 U22959 ( .C1(n19933), .C2(n19939), .A(n19932), .B(n19931), .ZN(
        P2_U3150) );
  AOI22_X1 U22960 ( .A1(n19935), .A2(n20068), .B1(n20066), .B2(n19934), .ZN(
        n19938) );
  AOI22_X1 U22961 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19936), .B1(
        n19973), .B2(n20070), .ZN(n19937) );
  OAI211_X1 U22962 ( .C1(n20076), .C2(n19939), .A(n19938), .B(n19937), .ZN(
        P2_U3151) );
  INV_X1 U22963 ( .A(n10479), .ZN(n19943) );
  NOR2_X1 U22964 ( .A1(n20202), .A2(n19944), .ZN(n19981) );
  NOR3_X1 U22965 ( .A1(n19943), .A2(n19981), .A3(n19942), .ZN(n19946) );
  INV_X1 U22966 ( .A(n19944), .ZN(n19952) );
  AOI21_X1 U22967 ( .B1(n20195), .B2(n19952), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19945) );
  AOI22_X1 U22968 ( .A1(n19971), .A2(n19524), .B1(n20017), .B2(n19981), .ZN(
        n19954) );
  INV_X1 U22969 ( .A(n19981), .ZN(n19948) );
  AOI211_X1 U22970 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19948), .A(n19947), 
        .B(n19946), .ZN(n19949) );
  OAI221_X1 U22971 ( .B1(n19952), .B2(n19951), .C1(n19952), .C2(n19950), .A(
        n19949), .ZN(n19974) );
  AOI22_X1 U22972 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19974), .B1(
        n19973), .B2(n20025), .ZN(n19953) );
  OAI211_X1 U22973 ( .C1(n20028), .C2(n20013), .A(n19954), .B(n19953), .ZN(
        P2_U3152) );
  AOI22_X1 U22974 ( .A1(n19971), .A2(n19534), .B1(n20029), .B2(n19981), .ZN(
        n19956) );
  AOI22_X1 U22975 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19974), .B1(
        n19973), .B2(n20030), .ZN(n19955) );
  OAI211_X1 U22976 ( .C1(n20033), .C2(n20013), .A(n19956), .B(n19955), .ZN(
        P2_U3153) );
  AOI22_X1 U22977 ( .A1(n19971), .A2(n20035), .B1(n20034), .B2(n19981), .ZN(
        n19958) );
  AOI22_X1 U22978 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19974), .B1(
        n19973), .B2(n20036), .ZN(n19957) );
  OAI211_X1 U22979 ( .C1(n20039), .C2(n20013), .A(n19958), .B(n19957), .ZN(
        P2_U3154) );
  AOI22_X1 U22980 ( .A1(n19971), .A2(n20041), .B1(n20040), .B2(n19981), .ZN(
        n19961) );
  AOI22_X1 U22981 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19974), .B1(
        n19973), .B2(n19959), .ZN(n19960) );
  OAI211_X1 U22982 ( .C1(n19962), .C2(n20013), .A(n19961), .B(n19960), .ZN(
        P2_U3155) );
  AOI22_X1 U22983 ( .A1(n19971), .A2(n20047), .B1(n9656), .B2(n19981), .ZN(
        n19964) );
  AOI22_X1 U22984 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19974), .B1(
        n19973), .B2(n20048), .ZN(n19963) );
  OAI211_X1 U22985 ( .C1(n20051), .C2(n20013), .A(n19964), .B(n19963), .ZN(
        P2_U3156) );
  AOI22_X1 U22986 ( .A1(n19971), .A2(n20053), .B1(n20052), .B2(n19981), .ZN(
        n19967) );
  AOI22_X1 U22987 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19974), .B1(
        n19973), .B2(n19965), .ZN(n19966) );
  OAI211_X1 U22988 ( .C1(n19968), .C2(n20013), .A(n19967), .B(n19966), .ZN(
        P2_U3157) );
  AOI22_X1 U22989 ( .A1(n19971), .A2(n20059), .B1(n20058), .B2(n19981), .ZN(
        n19970) );
  AOI22_X1 U22990 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19974), .B1(
        n19973), .B2(n20060), .ZN(n19969) );
  OAI211_X1 U22991 ( .C1(n20065), .C2(n20013), .A(n19970), .B(n19969), .ZN(
        P2_U3158) );
  AOI22_X1 U22992 ( .A1(n19971), .A2(n20068), .B1(n20066), .B2(n19981), .ZN(
        n19976) );
  AOI22_X1 U22993 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19974), .B1(
        n19973), .B2(n19972), .ZN(n19975) );
  OAI211_X1 U22994 ( .C1(n19977), .C2(n20013), .A(n19976), .B(n19975), .ZN(
        P2_U3159) );
  INV_X1 U22995 ( .A(n20013), .ZN(n20005) );
  NAND2_X1 U22996 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19979), .ZN(
        n20019) );
  NOR2_X1 U22997 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20019), .ZN(
        n20008) );
  AOI22_X1 U22998 ( .A1(n20025), .A2(n20005), .B1(n20017), .B2(n20008), .ZN(
        n19990) );
  AOI21_X1 U22999 ( .B1(n10483), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19983) );
  AOI21_X1 U23000 ( .B1(n20075), .B2(n20013), .A(n20226), .ZN(n19980) );
  NOR2_X1 U23001 ( .A1(n19980), .A2(n20016), .ZN(n19984) );
  NOR2_X1 U23002 ( .A1(n20008), .A2(n19981), .ZN(n19987) );
  NAND2_X1 U23003 ( .A1(n19984), .A2(n19987), .ZN(n19982) );
  OAI211_X1 U23004 ( .C1(n20008), .C2(n19983), .A(n19982), .B(n20022), .ZN(
        n20010) );
  INV_X1 U23005 ( .A(n19984), .ZN(n19988) );
  INV_X1 U23006 ( .A(n10483), .ZN(n19985) );
  OAI21_X1 U23007 ( .B1(n19985), .B2(n20008), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19986) );
  AOI22_X1 U23008 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20010), .B1(
        n19524), .B2(n20009), .ZN(n19989) );
  OAI211_X1 U23009 ( .C1(n20028), .C2(n20075), .A(n19990), .B(n19989), .ZN(
        P2_U3160) );
  AOI22_X1 U23010 ( .A1(n19991), .A2(n20061), .B1(n20029), .B2(n20008), .ZN(
        n19993) );
  AOI22_X1 U23011 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20010), .B1(
        n19534), .B2(n20009), .ZN(n19992) );
  OAI211_X1 U23012 ( .C1(n19994), .C2(n20013), .A(n19993), .B(n19992), .ZN(
        P2_U3161) );
  AOI22_X1 U23013 ( .A1(n20036), .A2(n20005), .B1(n20034), .B2(n20008), .ZN(
        n19996) );
  AOI22_X1 U23014 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20010), .B1(
        n20035), .B2(n20009), .ZN(n19995) );
  OAI211_X1 U23015 ( .C1(n20039), .C2(n20075), .A(n19996), .B(n19995), .ZN(
        P2_U3162) );
  AOI22_X1 U23016 ( .A1(n20042), .A2(n20061), .B1(n20040), .B2(n20008), .ZN(
        n19998) );
  AOI22_X1 U23017 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20010), .B1(
        n20041), .B2(n20009), .ZN(n19997) );
  OAI211_X1 U23018 ( .C1(n20045), .C2(n20013), .A(n19998), .B(n19997), .ZN(
        P2_U3163) );
  AOI22_X1 U23019 ( .A1(n19999), .A2(n20061), .B1(n9656), .B2(n20008), .ZN(
        n20001) );
  AOI22_X1 U23020 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20010), .B1(
        n20047), .B2(n20009), .ZN(n20000) );
  OAI211_X1 U23021 ( .C1(n20002), .C2(n20013), .A(n20001), .B(n20000), .ZN(
        P2_U3164) );
  AOI22_X1 U23022 ( .A1(n20054), .A2(n20061), .B1(n20052), .B2(n20008), .ZN(
        n20004) );
  AOI22_X1 U23023 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20010), .B1(
        n20053), .B2(n20009), .ZN(n20003) );
  OAI211_X1 U23024 ( .C1(n20057), .C2(n20013), .A(n20004), .B(n20003), .ZN(
        P2_U3165) );
  AOI22_X1 U23025 ( .A1(n20060), .A2(n20005), .B1(n20058), .B2(n20008), .ZN(
        n20007) );
  AOI22_X1 U23026 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20010), .B1(
        n20059), .B2(n20009), .ZN(n20006) );
  OAI211_X1 U23027 ( .C1(n20065), .C2(n20075), .A(n20007), .B(n20006), .ZN(
        P2_U3166) );
  AOI22_X1 U23028 ( .A1(n20070), .A2(n20061), .B1(n20066), .B2(n20008), .ZN(
        n20012) );
  AOI22_X1 U23029 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20010), .B1(
        n20068), .B2(n20009), .ZN(n20011) );
  OAI211_X1 U23030 ( .C1(n20076), .C2(n20013), .A(n20012), .B(n20011), .ZN(
        P2_U3167) );
  INV_X1 U23031 ( .A(n20018), .ZN(n20014) );
  OAI21_X1 U23032 ( .B1(n20014), .B2(n20067), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n20015) );
  OAI21_X1 U23033 ( .B1(n20019), .B2(n20016), .A(n20015), .ZN(n20069) );
  AOI22_X1 U23034 ( .A1(n20069), .A2(n19524), .B1(n20067), .B2(n20017), .ZN(
        n20027) );
  AOI21_X1 U23035 ( .B1(n9653), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n20024) );
  OAI21_X1 U23036 ( .B1(n20021), .B2(n20020), .A(n20019), .ZN(n20023) );
  OAI211_X1 U23037 ( .C1(n20067), .C2(n20024), .A(n20023), .B(n20022), .ZN(
        n20072) );
  AOI22_X1 U23038 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20072), .B1(
        n20061), .B2(n20025), .ZN(n20026) );
  OAI211_X1 U23039 ( .C1(n20028), .C2(n20064), .A(n20027), .B(n20026), .ZN(
        P2_U3168) );
  AOI22_X1 U23040 ( .A1(n20069), .A2(n19534), .B1(n20067), .B2(n20029), .ZN(
        n20032) );
  AOI22_X1 U23041 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20072), .B1(
        n20061), .B2(n20030), .ZN(n20031) );
  OAI211_X1 U23042 ( .C1(n20033), .C2(n20064), .A(n20032), .B(n20031), .ZN(
        P2_U3169) );
  AOI22_X1 U23043 ( .A1(n20069), .A2(n20035), .B1(n20067), .B2(n20034), .ZN(
        n20038) );
  AOI22_X1 U23044 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20072), .B1(
        n20061), .B2(n20036), .ZN(n20037) );
  OAI211_X1 U23045 ( .C1(n20039), .C2(n20064), .A(n20038), .B(n20037), .ZN(
        P2_U3170) );
  AOI22_X1 U23046 ( .A1(n20069), .A2(n20041), .B1(n20067), .B2(n20040), .ZN(
        n20044) );
  AOI22_X1 U23047 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20072), .B1(
        n20071), .B2(n20042), .ZN(n20043) );
  OAI211_X1 U23048 ( .C1(n20045), .C2(n20075), .A(n20044), .B(n20043), .ZN(
        P2_U3171) );
  AOI22_X1 U23049 ( .A1(n20069), .A2(n20047), .B1(n20067), .B2(n9656), .ZN(
        n20050) );
  AOI22_X1 U23050 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20072), .B1(
        n20061), .B2(n20048), .ZN(n20049) );
  OAI211_X1 U23051 ( .C1(n20051), .C2(n20064), .A(n20050), .B(n20049), .ZN(
        P2_U3172) );
  AOI22_X1 U23052 ( .A1(n20069), .A2(n20053), .B1(n20067), .B2(n20052), .ZN(
        n20056) );
  AOI22_X1 U23053 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20072), .B1(
        n20071), .B2(n20054), .ZN(n20055) );
  OAI211_X1 U23054 ( .C1(n20057), .C2(n20075), .A(n20056), .B(n20055), .ZN(
        P2_U3173) );
  AOI22_X1 U23055 ( .A1(n20069), .A2(n20059), .B1(n20067), .B2(n20058), .ZN(
        n20063) );
  AOI22_X1 U23056 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20072), .B1(
        n20061), .B2(n20060), .ZN(n20062) );
  OAI211_X1 U23057 ( .C1(n20065), .C2(n20064), .A(n20063), .B(n20062), .ZN(
        P2_U3174) );
  AOI22_X1 U23058 ( .A1(n20069), .A2(n20068), .B1(n20067), .B2(n20066), .ZN(
        n20074) );
  AOI22_X1 U23059 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20072), .B1(
        n20071), .B2(n20070), .ZN(n20073) );
  OAI211_X1 U23060 ( .C1(n20076), .C2(n20075), .A(n20074), .B(n20073), .ZN(
        P2_U3175) );
  INV_X1 U23061 ( .A(n20077), .ZN(n20081) );
  INV_X1 U23062 ( .A(n20078), .ZN(n20080) );
  OR4_X1 U23063 ( .A1(n20081), .A2(P2_STATE2_REG_1__SCAN_IN), .A3(n20080), 
        .A4(n20079), .ZN(n20082) );
  OAI221_X1 U23064 ( .B1(n14795), .B2(n20084), .C1(n14795), .C2(n20083), .A(
        n20082), .ZN(P2_U3177) );
  AND2_X1 U23065 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n20085), .ZN(
        P2_U3179) );
  AND2_X1 U23066 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n20085), .ZN(
        P2_U3180) );
  AND2_X1 U23067 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n20085), .ZN(
        P2_U3181) );
  AND2_X1 U23068 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n20085), .ZN(
        P2_U3182) );
  AND2_X1 U23069 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n20085), .ZN(
        P2_U3183) );
  AND2_X1 U23070 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n20085), .ZN(
        P2_U3184) );
  AND2_X1 U23071 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n20085), .ZN(
        P2_U3185) );
  AND2_X1 U23072 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n20085), .ZN(
        P2_U3186) );
  AND2_X1 U23073 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n20085), .ZN(
        P2_U3187) );
  AND2_X1 U23074 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n20085), .ZN(
        P2_U3188) );
  AND2_X1 U23075 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n20085), .ZN(
        P2_U3189) );
  AND2_X1 U23076 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n20085), .ZN(
        P2_U3190) );
  AND2_X1 U23077 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n20085), .ZN(
        P2_U3191) );
  AND2_X1 U23078 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n20085), .ZN(
        P2_U3192) );
  AND2_X1 U23079 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n20085), .ZN(
        P2_U3193) );
  AND2_X1 U23080 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n20085), .ZN(
        P2_U3194) );
  AND2_X1 U23081 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n20085), .ZN(
        P2_U3195) );
  AND2_X1 U23082 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n20085), .ZN(
        P2_U3196) );
  AND2_X1 U23083 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n20085), .ZN(
        P2_U3197) );
  AND2_X1 U23084 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n20085), .ZN(
        P2_U3198) );
  AND2_X1 U23085 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n20085), .ZN(
        P2_U3199) );
  AND2_X1 U23086 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n20085), .ZN(
        P2_U3200) );
  AND2_X1 U23087 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n20085), .ZN(P2_U3201) );
  AND2_X1 U23088 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n20085), .ZN(P2_U3202) );
  AND2_X1 U23089 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n20085), .ZN(P2_U3203) );
  AND2_X1 U23090 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n20085), .ZN(P2_U3204) );
  AND2_X1 U23091 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n20085), .ZN(P2_U3205) );
  AND2_X1 U23092 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n20085), .ZN(P2_U3206) );
  AND2_X1 U23093 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n20085), .ZN(P2_U3207) );
  AND2_X1 U23094 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n20085), .ZN(P2_U3208) );
  AND2_X1 U23095 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n20215), .ZN(n20097) );
  INV_X1 U23096 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n20232) );
  NOR3_X1 U23097 ( .A1(n20097), .A2(n20232), .A3(n20086), .ZN(n20089) );
  OAI211_X1 U23098 ( .C1(HOLD), .C2(n20232), .A(n20234), .B(n20087), .ZN(
        n20088) );
  NAND2_X1 U23099 ( .A1(NA), .A2(n20090), .ZN(n20095) );
  OAI211_X1 U23100 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n20089), .A(n20088), 
        .B(n20095), .ZN(P2_U3209) );
  NAND2_X1 U23101 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n20946), .ZN(n20096) );
  AOI211_X1 U23102 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(n20096), .A(n20090), 
        .B(n20232), .ZN(n20091) );
  NOR3_X1 U23103 ( .A1(n20219), .A2(n20097), .A3(n20091), .ZN(n20092) );
  OAI21_X1 U23104 ( .B1(n20946), .B2(n20093), .A(n20092), .ZN(P2_U3210) );
  INV_X1 U23105 ( .A(NA), .ZN(n21055) );
  AOI22_X1 U23106 ( .A1(n20094), .A2(n20232), .B1(n20097), .B2(n21055), .ZN(
        n20100) );
  OAI21_X1 U23107 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n20099) );
  OAI211_X1 U23108 ( .C1(n20097), .C2(n20096), .A(P2_STATE_REG_2__SCAN_IN), 
        .B(n20095), .ZN(n20098) );
  OAI21_X1 U23109 ( .B1(n20100), .B2(n20099), .A(n20098), .ZN(P2_U3211) );
  OAI222_X1 U23110 ( .A1(n20151), .A2(n20104), .B1(n20103), .B2(n20233), .C1(
        n20102), .C2(n20147), .ZN(P2_U3212) );
  OAI222_X1 U23111 ( .A1(n20151), .A2(n11419), .B1(n20105), .B2(n20233), .C1(
        n20104), .C2(n20147), .ZN(P2_U3213) );
  OAI222_X1 U23112 ( .A1(n20151), .A2(n14221), .B1(n20106), .B2(n20233), .C1(
        n11419), .C2(n20147), .ZN(P2_U3214) );
  OAI222_X1 U23113 ( .A1(n20151), .A2(n14463), .B1(n20107), .B2(n20233), .C1(
        n14221), .C2(n20147), .ZN(P2_U3215) );
  OAI222_X1 U23114 ( .A1(n20151), .A2(n20109), .B1(n20108), .B2(n20233), .C1(
        n14463), .C2(n20147), .ZN(P2_U3216) );
  OAI222_X1 U23115 ( .A1(n20151), .A2(n20111), .B1(n20110), .B2(n20233), .C1(
        n20109), .C2(n20147), .ZN(P2_U3217) );
  OAI222_X1 U23116 ( .A1(n20151), .A2(n11438), .B1(n20112), .B2(n20233), .C1(
        n20111), .C2(n20147), .ZN(P2_U3218) );
  OAI222_X1 U23117 ( .A1(n20151), .A2(n16056), .B1(n20113), .B2(n20233), .C1(
        n11438), .C2(n20147), .ZN(P2_U3219) );
  OAI222_X1 U23118 ( .A1(n20151), .A2(n11478), .B1(n20114), .B2(n20233), .C1(
        n16056), .C2(n20147), .ZN(P2_U3220) );
  OAI222_X1 U23119 ( .A1(n20151), .A2(n11523), .B1(n20115), .B2(n20233), .C1(
        n11478), .C2(n20147), .ZN(P2_U3221) );
  OAI222_X1 U23120 ( .A1(n20151), .A2(n11526), .B1(n20116), .B2(n20233), .C1(
        n11523), .C2(n20147), .ZN(P2_U3222) );
  OAI222_X1 U23121 ( .A1(n20151), .A2(n11564), .B1(n20117), .B2(n20233), .C1(
        n11526), .C2(n20147), .ZN(P2_U3223) );
  OAI222_X1 U23122 ( .A1(n20151), .A2(n11567), .B1(n20118), .B2(n20233), .C1(
        n11564), .C2(n20147), .ZN(P2_U3224) );
  OAI222_X1 U23123 ( .A1(n20151), .A2(n20120), .B1(n20119), .B2(n20233), .C1(
        n11567), .C2(n20147), .ZN(P2_U3225) );
  OAI222_X1 U23124 ( .A1(n20151), .A2(n15977), .B1(n20121), .B2(n20233), .C1(
        n20120), .C2(n20147), .ZN(P2_U3226) );
  OAI222_X1 U23125 ( .A1(n20151), .A2(n20123), .B1(n20122), .B2(n20233), .C1(
        n15977), .C2(n20147), .ZN(P2_U3227) );
  OAI222_X1 U23126 ( .A1(n20151), .A2(n20125), .B1(n20124), .B2(n20233), .C1(
        n20123), .C2(n20147), .ZN(P2_U3228) );
  OAI222_X1 U23127 ( .A1(n20151), .A2(n20127), .B1(n20126), .B2(n20233), .C1(
        n20125), .C2(n20147), .ZN(P2_U3229) );
  OAI222_X1 U23128 ( .A1(n20151), .A2(n20129), .B1(n20128), .B2(n20233), .C1(
        n20127), .C2(n20147), .ZN(P2_U3230) );
  OAI222_X1 U23129 ( .A1(n20151), .A2(n20131), .B1(n20130), .B2(n20233), .C1(
        n20129), .C2(n20147), .ZN(P2_U3231) );
  OAI222_X1 U23130 ( .A1(n20151), .A2(n11619), .B1(n20132), .B2(n20233), .C1(
        n20131), .C2(n20147), .ZN(P2_U3232) );
  OAI222_X1 U23131 ( .A1(n20151), .A2(n20134), .B1(n20133), .B2(n20233), .C1(
        n11619), .C2(n20147), .ZN(P2_U3233) );
  OAI222_X1 U23132 ( .A1(n20151), .A2(n20136), .B1(n20135), .B2(n20233), .C1(
        n20134), .C2(n20147), .ZN(P2_U3234) );
  OAI222_X1 U23133 ( .A1(n20151), .A2(n20138), .B1(n20137), .B2(n20233), .C1(
        n20136), .C2(n20147), .ZN(P2_U3235) );
  OAI222_X1 U23134 ( .A1(n20151), .A2(n20140), .B1(n20139), .B2(n20233), .C1(
        n20138), .C2(n20147), .ZN(P2_U3236) );
  OAI222_X1 U23135 ( .A1(n20151), .A2(n20143), .B1(n20141), .B2(n20233), .C1(
        n20140), .C2(n20147), .ZN(P2_U3237) );
  OAI222_X1 U23136 ( .A1(n20147), .A2(n20143), .B1(n20142), .B2(n20233), .C1(
        n15720), .C2(n20151), .ZN(P2_U3238) );
  OAI222_X1 U23137 ( .A1(n20151), .A2(n20145), .B1(n20144), .B2(n20233), .C1(
        n15720), .C2(n20147), .ZN(P2_U3239) );
  OAI222_X1 U23138 ( .A1(n20151), .A2(n20148), .B1(n20146), .B2(n20233), .C1(
        n20145), .C2(n20147), .ZN(P2_U3240) );
  INV_X1 U23139 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n20149) );
  OAI222_X1 U23140 ( .A1(n20151), .A2(n20150), .B1(n20149), .B2(n20233), .C1(
        n20148), .C2(n20147), .ZN(P2_U3241) );
  OAI22_X1 U23141 ( .A1(n20234), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n20233), .ZN(n20152) );
  INV_X1 U23142 ( .A(n20152), .ZN(P2_U3585) );
  MUX2_X1 U23143 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n20234), .Z(P2_U3586) );
  OAI22_X1 U23144 ( .A1(n20234), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n20233), .ZN(n20153) );
  INV_X1 U23145 ( .A(n20153), .ZN(P2_U3587) );
  OAI22_X1 U23146 ( .A1(n20234), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n20233), .ZN(n20154) );
  INV_X1 U23147 ( .A(n20154), .ZN(P2_U3588) );
  OAI21_X1 U23148 ( .B1(n20158), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n20156), 
        .ZN(n20155) );
  INV_X1 U23149 ( .A(n20155), .ZN(P2_U3591) );
  OAI21_X1 U23150 ( .B1(n20158), .B2(n20157), .A(n20156), .ZN(P2_U3592) );
  INV_X1 U23151 ( .A(n20159), .ZN(n20160) );
  OAI22_X1 U23152 ( .A1(n20167), .A2(n20161), .B1(n20165), .B2(n20160), .ZN(
        n20163) );
  MUX2_X1 U23153 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20163), .S(
        n20162), .Z(P2_U3596) );
  NAND2_X1 U23154 ( .A1(n20164), .A2(n20183), .ZN(n20176) );
  NAND3_X1 U23155 ( .A1(n20190), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n20165), 
        .ZN(n20166) );
  NAND2_X1 U23156 ( .A1(n20166), .A2(n20194), .ZN(n20177) );
  NAND2_X1 U23157 ( .A1(n20176), .A2(n20177), .ZN(n20173) );
  INV_X1 U23158 ( .A(n20167), .ZN(n20172) );
  INV_X1 U23159 ( .A(n20168), .ZN(n20171) );
  AOI222_X1 U23160 ( .A1(n20173), .A2(n20172), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n20171), .C1(n20170), .C2(n20169), .ZN(n20174) );
  AOI22_X1 U23161 ( .A1(n20203), .A2(n20175), .B1(n20174), .B2(n20200), .ZN(
        P2_U3602) );
  OAI21_X1 U23162 ( .B1(n20178), .B2(n20177), .A(n20176), .ZN(n20179) );
  AOI21_X1 U23163 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n20180), .A(n20179), 
        .ZN(n20181) );
  AOI22_X1 U23164 ( .A1(n20203), .A2(n20182), .B1(n20181), .B2(n20200), .ZN(
        P2_U3603) );
  INV_X1 U23165 ( .A(n20183), .ZN(n20189) );
  INV_X1 U23166 ( .A(n20184), .ZN(n20185) );
  NAND3_X1 U23167 ( .A1(n20190), .A2(n20194), .A3(n20185), .ZN(n20188) );
  NAND2_X1 U23168 ( .A1(n20186), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n20187) );
  OAI211_X1 U23169 ( .C1(n20190), .C2(n20189), .A(n20188), .B(n20187), .ZN(
        n20191) );
  INV_X1 U23170 ( .A(n20191), .ZN(n20192) );
  AOI22_X1 U23171 ( .A1(n20203), .A2(n20193), .B1(n20192), .B2(n20200), .ZN(
        P2_U3604) );
  INV_X1 U23172 ( .A(n20194), .ZN(n20196) );
  OAI22_X1 U23173 ( .A1(n20197), .A2(n20196), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20195), .ZN(n20198) );
  AOI21_X1 U23174 ( .B1(n20199), .B2(P2_STATE2_REG_2__SCAN_IN), .A(n20198), 
        .ZN(n20201) );
  AOI22_X1 U23175 ( .A1(n20203), .A2(n20202), .B1(n20201), .B2(n20200), .ZN(
        P2_U3605) );
  INV_X1 U23176 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n20204) );
  AOI22_X1 U23177 ( .A1(n20233), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n20204), 
        .B2(n20234), .ZN(P2_U3608) );
  AOI22_X1 U23178 ( .A1(n20208), .A2(n20207), .B1(n20206), .B2(n20205), .ZN(
        n20209) );
  NAND2_X1 U23179 ( .A1(n20210), .A2(n20209), .ZN(n20212) );
  MUX2_X1 U23180 ( .A(P2_MORE_REG_SCAN_IN), .B(n20212), .S(n20211), .Z(
        P2_U3609) );
  OAI21_X1 U23181 ( .B1(n20215), .B2(n20214), .A(n20213), .ZN(n20216) );
  AOI21_X1 U23182 ( .B1(n20195), .B2(n20217), .A(n20216), .ZN(n20231) );
  NOR4_X1 U23183 ( .A1(n10221), .A2(n9730), .A3(n20219), .A4(n20218), .ZN(
        n20223) );
  AOI21_X1 U23184 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n20221), .A(n20220), 
        .ZN(n20222) );
  NOR2_X1 U23185 ( .A1(n20223), .A2(n20222), .ZN(n20230) );
  INV_X1 U23186 ( .A(n20231), .ZN(n20228) );
  OAI211_X1 U23187 ( .C1(n20226), .C2(n20225), .A(n20224), .B(n9730), .ZN(
        n20227) );
  AND2_X1 U23188 ( .A1(n20228), .A2(n20227), .ZN(n20229) );
  AOI22_X1 U23189 ( .A1(n20232), .A2(n20231), .B1(n20230), .B2(n20229), .ZN(
        P2_U3610) );
  OAI22_X1 U23190 ( .A1(n20234), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n20233), .ZN(n20235) );
  INV_X1 U23191 ( .A(n20235), .ZN(P2_U3611) );
  AND2_X1 U23192 ( .A1(n20955), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n20236) );
  INV_X1 U23193 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n21173) );
  AOI21_X1 U23194 ( .B1(n20236), .B2(n21173), .A(n21031), .ZN(P1_U2802) );
  INV_X2 U23195 ( .A(n21031), .ZN(n21032) );
  NOR2_X1 U23196 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n20959) );
  OAI21_X1 U23197 ( .B1(n20959), .B2(P1_D_C_N_REG_SCAN_IN), .A(n21032), .ZN(
        n20237) );
  OAI21_X1 U23198 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n21032), .A(n20237), 
        .ZN(P1_U2804) );
  AOI21_X1 U23199 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20955), .A(n21031), 
        .ZN(n20945) );
  OAI21_X1 U23200 ( .B1(BS16), .B2(n20959), .A(n20945), .ZN(n21006) );
  OAI21_X1 U23201 ( .B1(n20945), .B2(n21170), .A(n21006), .ZN(P1_U2805) );
  OAI21_X1 U23202 ( .B1(n20239), .B2(n21212), .A(n20238), .ZN(P1_U2806) );
  NOR4_X1 U23203 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n20243) );
  NOR4_X1 U23204 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n20242) );
  NOR4_X1 U23205 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n20241) );
  NOR4_X1 U23206 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n20240) );
  NAND4_X1 U23207 ( .A1(n20243), .A2(n20242), .A3(n20241), .A4(n20240), .ZN(
        n20249) );
  NOR4_X1 U23208 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20247) );
  AOI211_X1 U23209 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_2__SCAN_IN), .B(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n20246) );
  NOR4_X1 U23210 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n20245) );
  NOR4_X1 U23211 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n20244) );
  NAND4_X1 U23212 ( .A1(n20247), .A2(n20246), .A3(n20245), .A4(n20244), .ZN(
        n20248) );
  NOR2_X1 U23213 ( .A1(n20249), .A2(n20248), .ZN(n21017) );
  INV_X1 U23214 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n20251) );
  NOR3_X1 U23215 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n20252) );
  OAI21_X1 U23216 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n20252), .A(n21017), .ZN(
        n20250) );
  OAI21_X1 U23217 ( .B1(n21017), .B2(n20251), .A(n20250), .ZN(P1_U2807) );
  INV_X1 U23218 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20254) );
  NOR2_X1 U23219 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21012) );
  OAI21_X1 U23220 ( .B1(n20252), .B2(n21012), .A(n21017), .ZN(n20253) );
  OAI21_X1 U23221 ( .B1(n21017), .B2(n20254), .A(n20253), .ZN(P1_U2808) );
  OR2_X1 U23222 ( .A1(n20256), .A2(n20255), .ZN(n20267) );
  AOI22_X1 U23223 ( .A1(n20258), .A2(n20338), .B1(n20320), .B2(n20257), .ZN(
        n20259) );
  OAI211_X1 U23224 ( .C1(n20335), .C2(n20260), .A(n20259), .B(n20289), .ZN(
        n20261) );
  AOI21_X1 U23225 ( .B1(n20321), .B2(P1_EBX_REG_9__SCAN_IN), .A(n20261), .ZN(
        n20266) );
  INV_X1 U23226 ( .A(n20262), .ZN(n20264) );
  AOI22_X1 U23227 ( .A1(n20264), .A2(n20287), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n20263), .ZN(n20265) );
  OAI211_X1 U23228 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n20267), .A(n20266), .B(
        n20265), .ZN(P1_U2831) );
  OAI22_X1 U23229 ( .A1(n20269), .A2(n20306), .B1(n20351), .B2(n20268), .ZN(
        n20274) );
  NAND4_X1 U23230 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(n20301), .A4(n20270), .ZN(n20271) );
  OAI211_X1 U23231 ( .C1(n20272), .C2(n20340), .A(n20271), .B(n20289), .ZN(
        n20273) );
  AOI211_X1 U23232 ( .C1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n20323), .A(
        n20274), .B(n20273), .ZN(n20280) );
  AND2_X1 U23233 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n20277) );
  NOR2_X1 U23234 ( .A1(n20276), .A2(n20275), .ZN(n20311) );
  AOI21_X1 U23235 ( .B1(n20277), .B2(n20311), .A(n20312), .ZN(n20286) );
  AOI22_X1 U23236 ( .A1(n20278), .A2(n20287), .B1(n20286), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n20279) );
  NAND2_X1 U23237 ( .A1(n20280), .A2(n20279), .ZN(P1_U2833) );
  INV_X1 U23238 ( .A(n20281), .ZN(n20283) );
  AOI22_X1 U23239 ( .A1(n20283), .A2(n20338), .B1(n20320), .B2(n20282), .ZN(
        n20292) );
  AOI22_X1 U23240 ( .A1(n20321), .A2(P1_EBX_REG_6__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20323), .ZN(n20291) );
  INV_X1 U23241 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20284) );
  OAI21_X1 U23242 ( .B1(n20312), .B2(n20311), .A(P1_REIP_REG_5__SCAN_IN), .ZN(
        n20300) );
  NAND2_X1 U23243 ( .A1(n20284), .A2(n20300), .ZN(n20285) );
  AOI22_X1 U23244 ( .A1(n20288), .A2(n20287), .B1(n20286), .B2(n20285), .ZN(
        n20290) );
  NAND4_X1 U23245 ( .A1(n20292), .A2(n20291), .A3(n20290), .A4(n20289), .ZN(
        P1_U2834) );
  INV_X1 U23246 ( .A(n20293), .ZN(n20295) );
  AOI22_X1 U23247 ( .A1(n20295), .A2(n20338), .B1(n20320), .B2(n20294), .ZN(
        n20304) );
  AOI21_X1 U23248 ( .B1(n20323), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n20310), .ZN(n20296) );
  OAI21_X1 U23249 ( .B1(n20340), .B2(n20297), .A(n20296), .ZN(n20298) );
  AOI21_X1 U23250 ( .B1(n20299), .B2(n20315), .A(n20298), .ZN(n20303) );
  OAI21_X1 U23251 ( .B1(P1_REIP_REG_5__SCAN_IN), .B2(n20301), .A(n20300), .ZN(
        n20302) );
  NAND3_X1 U23252 ( .A1(n20304), .A2(n20303), .A3(n20302), .ZN(P1_U2835) );
  INV_X1 U23253 ( .A(n20433), .ZN(n20305) );
  AOI22_X1 U23254 ( .A1(n20321), .A2(P1_EBX_REG_4__SCAN_IN), .B1(n20320), .B2(
        n20305), .ZN(n20318) );
  INV_X1 U23255 ( .A(n20346), .ZN(n20307) );
  OAI22_X1 U23256 ( .A1(n20308), .A2(n20307), .B1(n20426), .B2(n20306), .ZN(
        n20309) );
  AOI211_X1 U23257 ( .C1(n20323), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20310), .B(n20309), .ZN(n20317) );
  NAND2_X1 U23258 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n20319) );
  INV_X1 U23259 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20963) );
  OAI21_X1 U23260 ( .B1(n20319), .B2(n20333), .A(n20963), .ZN(n20314) );
  NOR2_X1 U23261 ( .A1(n20312), .A2(n20311), .ZN(n20313) );
  AOI22_X1 U23262 ( .A1(n20421), .A2(n20315), .B1(n20314), .B2(n20313), .ZN(
        n20316) );
  NAND3_X1 U23263 ( .A1(n20318), .A2(n20317), .A3(n20316), .ZN(P1_U2836) );
  OAI21_X1 U23264 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(P1_REIP_REG_2__SCAN_IN), 
        .A(n20319), .ZN(n20332) );
  AOI22_X1 U23265 ( .A1(n20321), .A2(P1_EBX_REG_3__SCAN_IN), .B1(n20320), .B2(
        n20441), .ZN(n20331) );
  INV_X1 U23266 ( .A(n20322), .ZN(n20324) );
  AOI22_X1 U23267 ( .A1(n20338), .A2(n20324), .B1(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n20323), .ZN(n20325) );
  OAI21_X1 U23268 ( .B1(n20326), .B2(n13964), .A(n20325), .ZN(n20329) );
  NOR2_X1 U23269 ( .A1(n20327), .A2(n20342), .ZN(n20328) );
  AOI211_X1 U23270 ( .C1(n20346), .C2(n13856), .A(n20329), .B(n20328), .ZN(
        n20330) );
  OAI211_X1 U23271 ( .C1(n20333), .C2(n20332), .A(n20331), .B(n20330), .ZN(
        P1_U2837) );
  OAI22_X1 U23272 ( .A1(n20335), .A2(n20337), .B1(n13702), .B2(n20334), .ZN(
        n20336) );
  AOI21_X1 U23273 ( .B1(n20338), .B2(n20337), .A(n20336), .ZN(n20339) );
  OAI21_X1 U23274 ( .B1(n20341), .B2(n20340), .A(n20339), .ZN(n20345) );
  NOR2_X1 U23275 ( .A1(n20343), .A2(n20342), .ZN(n20344) );
  AOI211_X1 U23276 ( .C1(n20346), .C2(n20841), .A(n20345), .B(n20344), .ZN(
        n20349) );
  NAND2_X1 U23277 ( .A1(n20347), .A2(n13702), .ZN(n20348) );
  OAI211_X1 U23278 ( .C1(n20351), .C2(n20350), .A(n20349), .B(n20348), .ZN(
        P1_U2839) );
  AOI22_X1 U23279 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20353) );
  OAI21_X1 U23280 ( .B1(n13665), .B2(n20375), .A(n20353), .ZN(P1_U2921) );
  AOI22_X1 U23281 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20354) );
  OAI21_X1 U23282 ( .B1(n14575), .B2(n20375), .A(n20354), .ZN(P1_U2922) );
  AOI22_X1 U23283 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20355) );
  OAI21_X1 U23284 ( .B1(n14530), .B2(n20375), .A(n20355), .ZN(P1_U2923) );
  AOI22_X1 U23285 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20356) );
  OAI21_X1 U23286 ( .B1(n14491), .B2(n20375), .A(n20356), .ZN(P1_U2924) );
  AOI22_X1 U23287 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20357) );
  OAI21_X1 U23288 ( .B1(n14553), .B2(n20375), .A(n20357), .ZN(P1_U2925) );
  AOI22_X1 U23289 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20358) );
  OAI21_X1 U23290 ( .B1(n14581), .B2(n20375), .A(n20358), .ZN(P1_U2926) );
  AOI22_X1 U23291 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20359) );
  OAI21_X1 U23292 ( .B1(n14441), .B2(n20375), .A(n20359), .ZN(P1_U2927) );
  AOI22_X1 U23293 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n21028), .B1(n16268), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20360) );
  OAI21_X1 U23294 ( .B1(n14418), .B2(n20375), .A(n20360), .ZN(P1_U2928) );
  AOI22_X1 U23295 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20373), .B1(n16268), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20361) );
  OAI21_X1 U23296 ( .B1(n12137), .B2(n20375), .A(n20361), .ZN(P1_U2929) );
  AOI22_X1 U23297 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20373), .B1(n16268), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20362) );
  OAI21_X1 U23298 ( .B1(n20363), .B2(n20375), .A(n20362), .ZN(P1_U2930) );
  AOI22_X1 U23299 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20373), .B1(n16268), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20364) );
  OAI21_X1 U23300 ( .B1(n14095), .B2(n20375), .A(n20364), .ZN(P1_U2931) );
  AOI22_X1 U23301 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20373), .B1(n16268), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20365) );
  OAI21_X1 U23302 ( .B1(n20366), .B2(n20375), .A(n20365), .ZN(P1_U2932) );
  AOI22_X1 U23303 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20373), .B1(n16268), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20367) );
  OAI21_X1 U23304 ( .B1(n20368), .B2(n20375), .A(n20367), .ZN(P1_U2933) );
  AOI22_X1 U23305 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20373), .B1(n16268), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20369) );
  OAI21_X1 U23306 ( .B1(n20370), .B2(n20375), .A(n20369), .ZN(P1_U2934) );
  AOI22_X1 U23307 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20373), .B1(n16268), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20371) );
  OAI21_X1 U23308 ( .B1(n20372), .B2(n20375), .A(n20371), .ZN(P1_U2935) );
  AOI22_X1 U23309 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20373), .B1(n16268), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20374) );
  OAI21_X1 U23310 ( .B1(n20376), .B2(n20375), .A(n20374), .ZN(P1_U2936) );
  AOI22_X1 U23311 ( .A1(n20413), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20383), .ZN(n20379) );
  INV_X1 U23312 ( .A(n20377), .ZN(n20378) );
  NAND2_X1 U23313 ( .A1(n20398), .A2(n20378), .ZN(n20400) );
  NAND2_X1 U23314 ( .A1(n20379), .A2(n20400), .ZN(P1_U2945) );
  AOI22_X1 U23315 ( .A1(n20413), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20383), .ZN(n20382) );
  INV_X1 U23316 ( .A(n20380), .ZN(n20381) );
  NAND2_X1 U23317 ( .A1(n20398), .A2(n20381), .ZN(n20402) );
  NAND2_X1 U23318 ( .A1(n20382), .A2(n20402), .ZN(P1_U2946) );
  AOI22_X1 U23319 ( .A1(n20413), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20383), .ZN(n20386) );
  INV_X1 U23320 ( .A(n20384), .ZN(n20385) );
  NAND2_X1 U23321 ( .A1(n20398), .A2(n20385), .ZN(n20404) );
  NAND2_X1 U23322 ( .A1(n20386), .A2(n20404), .ZN(P1_U2947) );
  AOI22_X1 U23323 ( .A1(n20413), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20412), .ZN(n20389) );
  INV_X1 U23324 ( .A(n20387), .ZN(n20388) );
  NAND2_X1 U23325 ( .A1(n20398), .A2(n20388), .ZN(n20406) );
  NAND2_X1 U23326 ( .A1(n20389), .A2(n20406), .ZN(P1_U2948) );
  AOI22_X1 U23327 ( .A1(n20413), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20412), .ZN(n20392) );
  INV_X1 U23328 ( .A(n20390), .ZN(n20391) );
  NAND2_X1 U23329 ( .A1(n20398), .A2(n20391), .ZN(n20408) );
  NAND2_X1 U23330 ( .A1(n20392), .A2(n20408), .ZN(P1_U2949) );
  AOI22_X1 U23331 ( .A1(n20413), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20412), .ZN(n20395) );
  INV_X1 U23332 ( .A(n20393), .ZN(n20394) );
  NAND2_X1 U23333 ( .A1(n20398), .A2(n20394), .ZN(n20410) );
  NAND2_X1 U23334 ( .A1(n20395), .A2(n20410), .ZN(P1_U2950) );
  AOI22_X1 U23335 ( .A1(n20413), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20383), .ZN(n20399) );
  INV_X1 U23336 ( .A(n20396), .ZN(n20397) );
  NAND2_X1 U23337 ( .A1(n20398), .A2(n20397), .ZN(n20414) );
  NAND2_X1 U23338 ( .A1(n20399), .A2(n20414), .ZN(P1_U2951) );
  AOI22_X1 U23339 ( .A1(n20413), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20412), .ZN(n20401) );
  NAND2_X1 U23340 ( .A1(n20401), .A2(n20400), .ZN(P1_U2960) );
  AOI22_X1 U23341 ( .A1(n20413), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20383), .ZN(n20403) );
  NAND2_X1 U23342 ( .A1(n20403), .A2(n20402), .ZN(P1_U2961) );
  AOI22_X1 U23343 ( .A1(n20413), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20412), .ZN(n20405) );
  NAND2_X1 U23344 ( .A1(n20405), .A2(n20404), .ZN(P1_U2962) );
  AOI22_X1 U23345 ( .A1(n20413), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20383), .ZN(n20407) );
  NAND2_X1 U23346 ( .A1(n20407), .A2(n20406), .ZN(P1_U2963) );
  AOI22_X1 U23347 ( .A1(n20413), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20412), .ZN(n20409) );
  NAND2_X1 U23348 ( .A1(n20409), .A2(n20408), .ZN(P1_U2964) );
  AOI22_X1 U23349 ( .A1(n20413), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20412), .ZN(n20411) );
  NAND2_X1 U23350 ( .A1(n20411), .A2(n20410), .ZN(P1_U2965) );
  AOI22_X1 U23351 ( .A1(n20413), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20412), .ZN(n20415) );
  NAND2_X1 U23352 ( .A1(n20415), .A2(n20414), .ZN(P1_U2966) );
  AOI22_X1 U23353 ( .A1(n20416), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20473), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20425) );
  OR2_X1 U23354 ( .A1(n20418), .A2(n20417), .ZN(n20419) );
  NAND2_X1 U23355 ( .A1(n20420), .A2(n20419), .ZN(n20431) );
  INV_X1 U23356 ( .A(n20431), .ZN(n20423) );
  AOI22_X1 U23357 ( .A1(n20423), .A2(n20422), .B1(n16364), .B2(n20421), .ZN(
        n20424) );
  OAI211_X1 U23358 ( .C1(n20427), .C2(n20426), .A(n20425), .B(n20424), .ZN(
        P1_U2995) );
  NOR2_X1 U23359 ( .A1(n20428), .A2(n20454), .ZN(n20429) );
  AOI211_X1 U23360 ( .C1(n20450), .C2(n20456), .A(n20429), .B(n20449), .ZN(
        n20448) );
  AOI211_X1 U23361 ( .C1(n20438), .C2(n20447), .A(n20430), .B(n20442), .ZN(
        n20436) );
  NOR2_X1 U23362 ( .A1(n20431), .A2(n20470), .ZN(n20435) );
  OAI22_X1 U23363 ( .A1(n20433), .A2(n20469), .B1(n20963), .B2(n20432), .ZN(
        n20434) );
  NOR3_X1 U23364 ( .A1(n20436), .A2(n20435), .A3(n20434), .ZN(n20437) );
  OAI21_X1 U23365 ( .B1(n20448), .B2(n20438), .A(n20437), .ZN(P1_U3027) );
  AOI21_X1 U23366 ( .B1(n20441), .B2(n20440), .A(n20439), .ZN(n20446) );
  INV_X1 U23367 ( .A(n20442), .ZN(n20443) );
  AOI22_X1 U23368 ( .A1(n20444), .A2(n20452), .B1(n20447), .B2(n20443), .ZN(
        n20445) );
  OAI211_X1 U23369 ( .C1(n20448), .C2(n20447), .A(n20446), .B(n20445), .ZN(
        P1_U3028) );
  AOI21_X1 U23370 ( .B1(n20451), .B2(n20450), .A(n20449), .ZN(n20463) );
  NAND3_X1 U23371 ( .A1(n20453), .A2(n13898), .A3(n20452), .ZN(n20459) );
  OAI21_X1 U23372 ( .B1(n20456), .B2(n20455), .A(n20454), .ZN(n20457) );
  AOI22_X1 U23373 ( .A1(n20467), .A2(n20457), .B1(n20473), .B2(
        P1_REIP_REG_2__SCAN_IN), .ZN(n20458) );
  OAI211_X1 U23374 ( .C1(n20469), .C2(n20460), .A(n20459), .B(n20458), .ZN(
        n20461) );
  INV_X1 U23375 ( .A(n20461), .ZN(n20462) );
  OAI221_X1 U23376 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20465), .C1(
        n20464), .C2(n20463), .A(n20462), .ZN(P1_U3029) );
  NOR3_X1 U23377 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n20467), .A3(
        n20466), .ZN(n20477) );
  OAI22_X1 U23378 ( .A1(n20471), .A2(n20470), .B1(n20469), .B2(n20468), .ZN(
        n20472) );
  AOI21_X1 U23379 ( .B1(n20473), .B2(P1_REIP_REG_0__SCAN_IN), .A(n20472), .ZN(
        n20474) );
  OAI221_X1 U23380 ( .B1(n20477), .B2(n20476), .C1(n20477), .C2(n20475), .A(
        n20474), .ZN(P1_U3031) );
  NOR2_X1 U23381 ( .A1(n12578), .A2(n20478), .ZN(P1_U3032) );
  AOI22_X1 U23382 ( .A1(n20926), .A2(n20849), .B1(n20497), .B2(n20883), .ZN(
        n20480) );
  AOI22_X1 U23383 ( .A1(n20882), .A2(n20499), .B1(n20526), .B2(n20889), .ZN(
        n20479) );
  OAI211_X1 U23384 ( .C1(n20498), .C2(n20481), .A(n20480), .B(n20479), .ZN(
        P1_U3033) );
  AOI22_X1 U23385 ( .A1(n20926), .A2(n20895), .B1(n20497), .B2(n20894), .ZN(
        n20483) );
  AOI22_X1 U23386 ( .A1(n20893), .A2(n20499), .B1(n20526), .B2(n20781), .ZN(
        n20482) );
  OAI211_X1 U23387 ( .C1(n20498), .C2(n20484), .A(n20483), .B(n20482), .ZN(
        P1_U3034) );
  AOI22_X1 U23388 ( .A1(n20926), .A2(n20901), .B1(n20497), .B2(n20900), .ZN(
        n20486) );
  AOI22_X1 U23389 ( .A1(n20899), .A2(n20499), .B1(n20526), .B2(n20784), .ZN(
        n20485) );
  OAI211_X1 U23390 ( .C1(n20498), .C2(n20487), .A(n20486), .B(n20485), .ZN(
        P1_U3035) );
  INV_X1 U23391 ( .A(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n20490) );
  AOI22_X1 U23392 ( .A1(n20926), .A2(n20907), .B1(n20497), .B2(n20906), .ZN(
        n20489) );
  AOI22_X1 U23393 ( .A1(n20905), .A2(n20499), .B1(n20526), .B2(n20787), .ZN(
        n20488) );
  OAI211_X1 U23394 ( .C1(n20498), .C2(n20490), .A(n20489), .B(n20488), .ZN(
        P1_U3036) );
  AOI22_X1 U23395 ( .A1(n20926), .A2(n20919), .B1(n20497), .B2(n20918), .ZN(
        n20492) );
  AOI22_X1 U23396 ( .A1(n20917), .A2(n20499), .B1(n20526), .B2(n20792), .ZN(
        n20491) );
  OAI211_X1 U23397 ( .C1(n20498), .C2(n20493), .A(n20492), .B(n20491), .ZN(
        P1_U3038) );
  INV_X1 U23398 ( .A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n20496) );
  AOI22_X1 U23399 ( .A1(n20926), .A2(n20865), .B1(n20497), .B2(n20924), .ZN(
        n20495) );
  AOI22_X1 U23400 ( .A1(n20923), .A2(n20499), .B1(n20526), .B2(n20925), .ZN(
        n20494) );
  OAI211_X1 U23401 ( .C1(n20498), .C2(n20496), .A(n20495), .B(n20494), .ZN(
        P1_U3039) );
  AOI22_X1 U23402 ( .A1(n20926), .A2(n20935), .B1(n20497), .B2(n20934), .ZN(
        n20502) );
  INV_X1 U23403 ( .A(n20498), .ZN(n20500) );
  AOI22_X1 U23404 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20500), .B1(
        n20932), .B2(n20499), .ZN(n20501) );
  OAI211_X1 U23405 ( .C1(n20941), .C2(n20511), .A(n20502), .B(n20501), .ZN(
        P1_U3040) );
  NOR2_X1 U23406 ( .A1(n20733), .A2(n20505), .ZN(n20525) );
  INV_X1 U23407 ( .A(n20568), .ZN(n20504) );
  INV_X1 U23408 ( .A(n20503), .ZN(n20734) );
  AOI21_X1 U23409 ( .B1(n20504), .B2(n20734), .A(n20525), .ZN(n20506) );
  OAI22_X1 U23410 ( .A1(n20506), .A2(n20880), .B1(n20505), .B2(n12006), .ZN(
        n20524) );
  AOI22_X1 U23411 ( .A1(n20883), .A2(n20525), .B1(n20524), .B2(n20882), .ZN(
        n20510) );
  OAI211_X1 U23412 ( .C1(n20580), .C2(n21170), .A(n20811), .B(n20506), .ZN(
        n20507) );
  OAI211_X1 U23413 ( .C1(n20811), .C2(n20508), .A(n20886), .B(n20507), .ZN(
        n20527) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20527), .B1(
        n20553), .B2(n20889), .ZN(n20509) );
  OAI211_X1 U23415 ( .C1(n20892), .C2(n20511), .A(n20510), .B(n20509), .ZN(
        P1_U3041) );
  AOI22_X1 U23416 ( .A1(n20894), .A2(n20525), .B1(n20524), .B2(n20893), .ZN(
        n20513) );
  AOI22_X1 U23417 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20527), .B1(
        n20526), .B2(n20895), .ZN(n20512) );
  OAI211_X1 U23418 ( .C1(n20898), .C2(n20560), .A(n20513), .B(n20512), .ZN(
        P1_U3042) );
  AOI22_X1 U23419 ( .A1(n20900), .A2(n20525), .B1(n20524), .B2(n20899), .ZN(
        n20515) );
  AOI22_X1 U23420 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20527), .B1(
        n20526), .B2(n20901), .ZN(n20514) );
  OAI211_X1 U23421 ( .C1(n20904), .C2(n20560), .A(n20515), .B(n20514), .ZN(
        P1_U3043) );
  AOI22_X1 U23422 ( .A1(n20906), .A2(n20525), .B1(n20524), .B2(n20905), .ZN(
        n20517) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20527), .B1(
        n20526), .B2(n20907), .ZN(n20516) );
  OAI211_X1 U23424 ( .C1(n20910), .C2(n20560), .A(n20517), .B(n20516), .ZN(
        P1_U3044) );
  AOI22_X1 U23425 ( .A1(n20912), .A2(n20525), .B1(n20524), .B2(n20911), .ZN(
        n20519) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20527), .B1(
        n20526), .B2(n20859), .ZN(n20518) );
  OAI211_X1 U23427 ( .C1(n20862), .C2(n20560), .A(n20519), .B(n20518), .ZN(
        P1_U3045) );
  AOI22_X1 U23428 ( .A1(n20918), .A2(n20525), .B1(n20524), .B2(n20917), .ZN(
        n20521) );
  AOI22_X1 U23429 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20527), .B1(
        n20526), .B2(n20919), .ZN(n20520) );
  OAI211_X1 U23430 ( .C1(n20922), .C2(n20560), .A(n20521), .B(n20520), .ZN(
        P1_U3046) );
  AOI22_X1 U23431 ( .A1(n20924), .A2(n20525), .B1(n20524), .B2(n20923), .ZN(
        n20523) );
  AOI22_X1 U23432 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20527), .B1(
        n20865), .B2(n20526), .ZN(n20522) );
  OAI211_X1 U23433 ( .C1(n20868), .C2(n20560), .A(n20523), .B(n20522), .ZN(
        P1_U3047) );
  AOI22_X1 U23434 ( .A1(n20934), .A2(n20525), .B1(n20524), .B2(n20932), .ZN(
        n20529) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20527), .B1(
        n20526), .B2(n20935), .ZN(n20528) );
  OAI211_X1 U23436 ( .C1(n20941), .C2(n20560), .A(n20529), .B(n20528), .ZN(
        P1_U3048) );
  NOR3_X1 U23437 ( .A1(n20611), .A2(n20553), .A3(n20880), .ZN(n20530) );
  INV_X1 U23438 ( .A(n20766), .ZN(n20671) );
  NOR2_X1 U23439 ( .A1(n20530), .A2(n20671), .ZN(n20537) );
  INV_X1 U23440 ( .A(n20537), .ZN(n20531) );
  NOR2_X1 U23441 ( .A1(n20568), .A2(n14392), .ZN(n20536) );
  INV_X1 U23442 ( .A(n20883), .ZN(n20572) );
  NOR3_X1 U23443 ( .A1(n20532), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20574) );
  NAND2_X1 U23444 ( .A1(n20733), .A2(n20574), .ZN(n20559) );
  OAI22_X1 U23445 ( .A1(n20588), .A2(n20852), .B1(n20572), .B2(n20559), .ZN(
        n20533) );
  INV_X1 U23446 ( .A(n20533), .ZN(n20539) );
  NOR2_X1 U23447 ( .A1(n10112), .A2(n12006), .ZN(n20677) );
  INV_X1 U23448 ( .A(n20773), .ZN(n20534) );
  AOI211_X1 U23449 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n20559), .A(n20677), 
        .B(n20534), .ZN(n20535) );
  AOI22_X1 U23450 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20562), .B1(
        n20553), .B2(n20849), .ZN(n20538) );
  OAI211_X1 U23451 ( .C1(n20565), .C2(n9680), .A(n20539), .B(n20538), .ZN(
        P1_U3049) );
  INV_X1 U23452 ( .A(n20894), .ZN(n20583) );
  OAI22_X1 U23453 ( .A1(n20588), .A2(n20898), .B1(n20583), .B2(n20559), .ZN(
        n20540) );
  INV_X1 U23454 ( .A(n20540), .ZN(n20542) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20562), .B1(
        n20553), .B2(n20895), .ZN(n20541) );
  OAI211_X1 U23456 ( .C1(n20565), .C2(n9678), .A(n20542), .B(n20541), .ZN(
        P1_U3050) );
  INV_X1 U23457 ( .A(n20900), .ZN(n20587) );
  OAI22_X1 U23458 ( .A1(n20560), .A2(n20747), .B1(n20587), .B2(n20559), .ZN(
        n20543) );
  INV_X1 U23459 ( .A(n20543), .ZN(n20545) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20562), .B1(
        n20611), .B2(n20784), .ZN(n20544) );
  OAI211_X1 U23461 ( .C1(n20565), .C2(n9679), .A(n20545), .B(n20544), .ZN(
        P1_U3051) );
  INV_X1 U23462 ( .A(n20906), .ZN(n20592) );
  OAI22_X1 U23463 ( .A1(n20588), .A2(n20910), .B1(n20592), .B2(n20559), .ZN(
        n20546) );
  INV_X1 U23464 ( .A(n20546), .ZN(n20548) );
  AOI22_X1 U23465 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20562), .B1(
        n20553), .B2(n20907), .ZN(n20547) );
  OAI211_X1 U23466 ( .C1(n20565), .C2(n9676), .A(n20548), .B(n20547), .ZN(
        P1_U3052) );
  INV_X1 U23467 ( .A(n20912), .ZN(n20596) );
  OAI22_X1 U23468 ( .A1(n20588), .A2(n20862), .B1(n20596), .B2(n20559), .ZN(
        n20549) );
  INV_X1 U23469 ( .A(n20549), .ZN(n20551) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20562), .B1(
        n20553), .B2(n20859), .ZN(n20550) );
  OAI211_X1 U23471 ( .C1(n20565), .C2(n9677), .A(n20551), .B(n20550), .ZN(
        P1_U3053) );
  INV_X1 U23472 ( .A(n20918), .ZN(n20600) );
  OAI22_X1 U23473 ( .A1(n20588), .A2(n20922), .B1(n20600), .B2(n20559), .ZN(
        n20552) );
  INV_X1 U23474 ( .A(n20552), .ZN(n20555) );
  AOI22_X1 U23475 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20562), .B1(
        n20553), .B2(n20919), .ZN(n20554) );
  OAI211_X1 U23476 ( .C1(n20565), .C2(n9682), .A(n20555), .B(n20554), .ZN(
        P1_U3054) );
  INV_X1 U23477 ( .A(n20924), .ZN(n20604) );
  OAI22_X1 U23478 ( .A1(n20560), .A2(n20930), .B1(n20604), .B2(n20559), .ZN(
        n20556) );
  INV_X1 U23479 ( .A(n20556), .ZN(n20558) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20562), .B1(
        n20611), .B2(n20925), .ZN(n20557) );
  OAI211_X1 U23481 ( .C1(n20565), .C2(n20797), .A(n20558), .B(n20557), .ZN(
        P1_U3055) );
  INV_X1 U23482 ( .A(n20934), .ZN(n20609) );
  OAI22_X1 U23483 ( .A1(n20560), .A2(n20764), .B1(n20609), .B2(n20559), .ZN(
        n20561) );
  INV_X1 U23484 ( .A(n20561), .ZN(n20564) );
  AOI22_X1 U23485 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20562), .B1(
        n20611), .B2(n20799), .ZN(n20563) );
  OAI211_X1 U23486 ( .C1(n20565), .C2(n9681), .A(n20564), .B(n20563), .ZN(
        P1_U3056) );
  INV_X1 U23487 ( .A(n20580), .ZN(n20567) );
  OAI21_X1 U23488 ( .B1(n20567), .B2(n20880), .A(n20566), .ZN(n20576) );
  OR2_X1 U23489 ( .A1(n20568), .A2(n20876), .ZN(n20570) );
  INV_X1 U23490 ( .A(n20569), .ZN(n20806) );
  NAND2_X1 U23491 ( .A1(n20806), .A2(n20768), .ZN(n20608) );
  AND2_X1 U23492 ( .A1(n20570), .A2(n20608), .ZN(n20577) );
  INV_X1 U23493 ( .A(n20577), .ZN(n20571) );
  OAI22_X1 U23494 ( .A1(n20588), .A2(n20892), .B1(n20572), .B2(n20608), .ZN(
        n20573) );
  INV_X1 U23495 ( .A(n20573), .ZN(n20582) );
  INV_X1 U23496 ( .A(n20574), .ZN(n20575) );
  AOI22_X1 U23497 ( .A1(n20577), .A2(n20576), .B1(n20880), .B2(n20575), .ZN(
        n20578) );
  NAND2_X1 U23498 ( .A1(n20886), .A2(n20578), .ZN(n20612) );
  AOI22_X1 U23499 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20612), .B1(
        n20640), .B2(n20889), .ZN(n20581) );
  OAI211_X1 U23500 ( .C1(n20615), .C2(n9680), .A(n20582), .B(n20581), .ZN(
        P1_U3057) );
  OAI22_X1 U23501 ( .A1(n20620), .A2(n20898), .B1(n20583), .B2(n20608), .ZN(
        n20584) );
  INV_X1 U23502 ( .A(n20584), .ZN(n20586) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20612), .B1(
        n20611), .B2(n20895), .ZN(n20585) );
  OAI211_X1 U23504 ( .C1(n20615), .C2(n9678), .A(n20586), .B(n20585), .ZN(
        P1_U3058) );
  OAI22_X1 U23505 ( .A1(n20588), .A2(n20747), .B1(n20587), .B2(n20608), .ZN(
        n20589) );
  INV_X1 U23506 ( .A(n20589), .ZN(n20591) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20612), .B1(
        n20640), .B2(n20784), .ZN(n20590) );
  OAI211_X1 U23508 ( .C1(n20615), .C2(n9679), .A(n20591), .B(n20590), .ZN(
        P1_U3059) );
  OAI22_X1 U23509 ( .A1(n20620), .A2(n20910), .B1(n20592), .B2(n20608), .ZN(
        n20593) );
  INV_X1 U23510 ( .A(n20593), .ZN(n20595) );
  AOI22_X1 U23511 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20612), .B1(
        n20611), .B2(n20907), .ZN(n20594) );
  OAI211_X1 U23512 ( .C1(n20615), .C2(n9676), .A(n20595), .B(n20594), .ZN(
        P1_U3060) );
  OAI22_X1 U23513 ( .A1(n20620), .A2(n20862), .B1(n20596), .B2(n20608), .ZN(
        n20597) );
  INV_X1 U23514 ( .A(n20597), .ZN(n20599) );
  AOI22_X1 U23515 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20612), .B1(
        n20611), .B2(n20859), .ZN(n20598) );
  OAI211_X1 U23516 ( .C1(n20615), .C2(n9677), .A(n20599), .B(n20598), .ZN(
        P1_U3061) );
  OAI22_X1 U23517 ( .A1(n20620), .A2(n20922), .B1(n20600), .B2(n20608), .ZN(
        n20601) );
  INV_X1 U23518 ( .A(n20601), .ZN(n20603) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20612), .B1(
        n20611), .B2(n20919), .ZN(n20602) );
  OAI211_X1 U23520 ( .C1(n20615), .C2(n9682), .A(n20603), .B(n20602), .ZN(
        P1_U3062) );
  OAI22_X1 U23521 ( .A1(n20620), .A2(n20868), .B1(n20604), .B2(n20608), .ZN(
        n20605) );
  INV_X1 U23522 ( .A(n20605), .ZN(n20607) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20612), .B1(
        n20611), .B2(n20865), .ZN(n20606) );
  OAI211_X1 U23524 ( .C1(n20615), .C2(n20797), .A(n20607), .B(n20606), .ZN(
        P1_U3063) );
  OAI22_X1 U23525 ( .A1(n20620), .A2(n20941), .B1(n20609), .B2(n20608), .ZN(
        n20610) );
  INV_X1 U23526 ( .A(n20610), .ZN(n20614) );
  AOI22_X1 U23527 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20612), .B1(
        n20611), .B2(n20935), .ZN(n20613) );
  OAI211_X1 U23528 ( .C1(n20615), .C2(n9681), .A(n20614), .B(n20613), .ZN(
        P1_U3064) );
  INV_X1 U23529 ( .A(n20649), .ZN(n20617) );
  NOR3_X1 U23530 ( .A1(n16225), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20648) );
  INV_X1 U23531 ( .A(n20648), .ZN(n20645) );
  NOR2_X1 U23532 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20645), .ZN(
        n20639) );
  INV_X1 U23533 ( .A(n20674), .ZN(n20843) );
  INV_X1 U23534 ( .A(n20673), .ZN(n20644) );
  NAND3_X1 U23535 ( .A1(n20644), .A2(n20811), .A3(n14392), .ZN(n20618) );
  OAI21_X1 U23536 ( .B1(n20843), .B2(n20619), .A(n20618), .ZN(n20638) );
  AOI22_X1 U23537 ( .A1(n20883), .A2(n20639), .B1(n20882), .B2(n20638), .ZN(
        n20625) );
  AOI21_X1 U23538 ( .B1(n20620), .B2(n20669), .A(n21170), .ZN(n20621) );
  AOI21_X1 U23539 ( .B1(n20644), .B2(n14392), .A(n20621), .ZN(n20622) );
  NOR2_X1 U23540 ( .A1(n20622), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20623) );
  AOI22_X1 U23541 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20849), .ZN(n20624) );
  OAI211_X1 U23542 ( .C1(n20852), .C2(n20669), .A(n20625), .B(n20624), .ZN(
        P1_U3065) );
  AOI22_X1 U23543 ( .A1(n20894), .A2(n20639), .B1(n20893), .B2(n20638), .ZN(
        n20627) );
  AOI22_X1 U23544 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20895), .ZN(n20626) );
  OAI211_X1 U23545 ( .C1(n20898), .C2(n20669), .A(n20627), .B(n20626), .ZN(
        P1_U3066) );
  AOI22_X1 U23546 ( .A1(n20900), .A2(n20639), .B1(n20899), .B2(n20638), .ZN(
        n20629) );
  AOI22_X1 U23547 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20641), .B1(
        n20901), .B2(n20640), .ZN(n20628) );
  OAI211_X1 U23548 ( .C1(n20904), .C2(n20669), .A(n20629), .B(n20628), .ZN(
        P1_U3067) );
  AOI22_X1 U23549 ( .A1(n20906), .A2(n20639), .B1(n20905), .B2(n20638), .ZN(
        n20631) );
  AOI22_X1 U23550 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20907), .ZN(n20630) );
  OAI211_X1 U23551 ( .C1(n20910), .C2(n20669), .A(n20631), .B(n20630), .ZN(
        P1_U3068) );
  AOI22_X1 U23552 ( .A1(n20912), .A2(n20639), .B1(n20911), .B2(n20638), .ZN(
        n20633) );
  AOI22_X1 U23553 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20859), .ZN(n20632) );
  OAI211_X1 U23554 ( .C1(n20862), .C2(n20669), .A(n20633), .B(n20632), .ZN(
        P1_U3069) );
  AOI22_X1 U23555 ( .A1(n20918), .A2(n20639), .B1(n20917), .B2(n20638), .ZN(
        n20635) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20919), .ZN(n20634) );
  OAI211_X1 U23557 ( .C1(n20922), .C2(n20669), .A(n20635), .B(n20634), .ZN(
        P1_U3070) );
  AOI22_X1 U23558 ( .A1(n20924), .A2(n20639), .B1(n20923), .B2(n20638), .ZN(
        n20637) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20865), .ZN(n20636) );
  OAI211_X1 U23560 ( .C1(n20868), .C2(n20669), .A(n20637), .B(n20636), .ZN(
        P1_U3071) );
  AOI22_X1 U23561 ( .A1(n20934), .A2(n20639), .B1(n20932), .B2(n20638), .ZN(
        n20643) );
  AOI22_X1 U23562 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20935), .ZN(n20642) );
  OAI211_X1 U23563 ( .C1(n20941), .C2(n20669), .A(n20643), .B(n20642), .ZN(
        P1_U3072) );
  NOR2_X1 U23564 ( .A1(n20733), .A2(n20645), .ZN(n20665) );
  AOI21_X1 U23565 ( .B1(n20644), .B2(n20734), .A(n20665), .ZN(n20646) );
  OAI22_X1 U23566 ( .A1(n20646), .A2(n20880), .B1(n20645), .B2(n12006), .ZN(
        n20664) );
  AOI22_X1 U23567 ( .A1(n20883), .A2(n20665), .B1(n20882), .B2(n20664), .ZN(
        n20651) );
  OAI211_X1 U23568 ( .C1(n20649), .C2(n21170), .A(n20811), .B(n20646), .ZN(
        n20647) );
  OAI211_X1 U23569 ( .C1(n20811), .C2(n20648), .A(n20886), .B(n20647), .ZN(
        n20666) );
  AOI22_X1 U23570 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20666), .B1(
        n20698), .B2(n20889), .ZN(n20650) );
  OAI211_X1 U23571 ( .C1(n20892), .C2(n20669), .A(n20651), .B(n20650), .ZN(
        P1_U3073) );
  AOI22_X1 U23572 ( .A1(n20894), .A2(n20665), .B1(n20893), .B2(n20664), .ZN(
        n20653) );
  AOI22_X1 U23573 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20666), .B1(
        n20698), .B2(n20781), .ZN(n20652) );
  OAI211_X1 U23574 ( .C1(n20744), .C2(n20669), .A(n20653), .B(n20652), .ZN(
        P1_U3074) );
  AOI22_X1 U23575 ( .A1(n20900), .A2(n20665), .B1(n20899), .B2(n20664), .ZN(
        n20655) );
  AOI22_X1 U23576 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20666), .B1(
        n20698), .B2(n20784), .ZN(n20654) );
  OAI211_X1 U23577 ( .C1(n20747), .C2(n20669), .A(n20655), .B(n20654), .ZN(
        P1_U3075) );
  AOI22_X1 U23578 ( .A1(n20906), .A2(n20665), .B1(n20905), .B2(n20664), .ZN(
        n20657) );
  AOI22_X1 U23579 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20666), .B1(
        n20698), .B2(n20787), .ZN(n20656) );
  OAI211_X1 U23580 ( .C1(n20750), .C2(n20669), .A(n20657), .B(n20656), .ZN(
        P1_U3076) );
  AOI22_X1 U23581 ( .A1(n20912), .A2(n20665), .B1(n20911), .B2(n20664), .ZN(
        n20659) );
  AOI22_X1 U23582 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20666), .B1(
        n20698), .B2(n20913), .ZN(n20658) );
  OAI211_X1 U23583 ( .C1(n20916), .C2(n20669), .A(n20659), .B(n20658), .ZN(
        P1_U3077) );
  AOI22_X1 U23584 ( .A1(n20918), .A2(n20665), .B1(n20917), .B2(n20664), .ZN(
        n20661) );
  AOI22_X1 U23585 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20666), .B1(
        n20698), .B2(n20792), .ZN(n20660) );
  OAI211_X1 U23586 ( .C1(n20755), .C2(n20669), .A(n20661), .B(n20660), .ZN(
        P1_U3078) );
  AOI22_X1 U23587 ( .A1(n20924), .A2(n20665), .B1(n20923), .B2(n20664), .ZN(
        n20663) );
  AOI22_X1 U23588 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20666), .B1(
        n20698), .B2(n20925), .ZN(n20662) );
  OAI211_X1 U23589 ( .C1(n20930), .C2(n20669), .A(n20663), .B(n20662), .ZN(
        P1_U3079) );
  AOI22_X1 U23590 ( .A1(n20934), .A2(n20665), .B1(n20932), .B2(n20664), .ZN(
        n20668) );
  AOI22_X1 U23591 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20666), .B1(
        n20698), .B2(n20799), .ZN(n20667) );
  OAI211_X1 U23592 ( .C1(n20764), .C2(n20669), .A(n20668), .B(n20667), .ZN(
        P1_U3080) );
  NOR3_X1 U23593 ( .A1(n20698), .A2(n20699), .A3(n20880), .ZN(n20672) );
  NOR2_X1 U23594 ( .A1(n20672), .A2(n20671), .ZN(n20682) );
  INV_X1 U23595 ( .A(n20682), .ZN(n20675) );
  NOR2_X1 U23596 ( .A1(n20673), .A2(n14392), .ZN(n20681) );
  NOR2_X1 U23597 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20676), .ZN(
        n20697) );
  AOI22_X1 U23598 ( .A1(n20698), .A2(n20849), .B1(n20883), .B2(n20697), .ZN(
        n20684) );
  INV_X1 U23599 ( .A(n20677), .ZN(n20678) );
  OAI211_X1 U23600 ( .C1(n20774), .C2(n20697), .A(n20678), .B(n20847), .ZN(
        n20679) );
  INV_X1 U23601 ( .A(n20679), .ZN(n20680) );
  AOI22_X1 U23602 ( .A1(n20700), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n20889), .B2(n20699), .ZN(n20683) );
  OAI211_X1 U23603 ( .C1(n20703), .C2(n9680), .A(n20684), .B(n20683), .ZN(
        P1_U3081) );
  AOI22_X1 U23604 ( .A1(n20698), .A2(n20895), .B1(n20894), .B2(n20697), .ZN(
        n20686) );
  AOI22_X1 U23605 ( .A1(n20700), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n20781), .B2(n20699), .ZN(n20685) );
  OAI211_X1 U23606 ( .C1(n20703), .C2(n9678), .A(n20686), .B(n20685), .ZN(
        P1_U3082) );
  AOI22_X1 U23607 ( .A1(n20698), .A2(n20901), .B1(n20900), .B2(n20697), .ZN(
        n20688) );
  AOI22_X1 U23608 ( .A1(n20700), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n20784), .B2(n20699), .ZN(n20687) );
  OAI211_X1 U23609 ( .C1(n20703), .C2(n9679), .A(n20688), .B(n20687), .ZN(
        P1_U3083) );
  AOI22_X1 U23610 ( .A1(n20698), .A2(n20907), .B1(n20906), .B2(n20697), .ZN(
        n20690) );
  AOI22_X1 U23611 ( .A1(n20700), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n20787), .B2(n20699), .ZN(n20689) );
  OAI211_X1 U23612 ( .C1(n20703), .C2(n9676), .A(n20690), .B(n20689), .ZN(
        P1_U3084) );
  AOI22_X1 U23613 ( .A1(n20698), .A2(n20859), .B1(n20912), .B2(n20697), .ZN(
        n20692) );
  AOI22_X1 U23614 ( .A1(n20700), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n20913), .B2(n20699), .ZN(n20691) );
  OAI211_X1 U23615 ( .C1(n20703), .C2(n9677), .A(n20692), .B(n20691), .ZN(
        P1_U3085) );
  AOI22_X1 U23616 ( .A1(n20698), .A2(n20919), .B1(n20918), .B2(n20697), .ZN(
        n20694) );
  AOI22_X1 U23617 ( .A1(n20700), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n20792), .B2(n20699), .ZN(n20693) );
  OAI211_X1 U23618 ( .C1(n20703), .C2(n9682), .A(n20694), .B(n20693), .ZN(
        P1_U3086) );
  AOI22_X1 U23619 ( .A1(n20698), .A2(n20865), .B1(n20924), .B2(n20697), .ZN(
        n20696) );
  AOI22_X1 U23620 ( .A1(n20700), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n20925), .B2(n20699), .ZN(n20695) );
  OAI211_X1 U23621 ( .C1(n20703), .C2(n20797), .A(n20696), .B(n20695), .ZN(
        P1_U3087) );
  AOI22_X1 U23622 ( .A1(n20698), .A2(n20935), .B1(n20934), .B2(n20697), .ZN(
        n20702) );
  AOI22_X1 U23623 ( .A1(n20700), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n20799), .B2(n20699), .ZN(n20701) );
  OAI211_X1 U23624 ( .C1(n20703), .C2(n9681), .A(n20702), .B(n20701), .ZN(
        P1_U3088) );
  NOR3_X1 U23625 ( .A1(n20768), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20738) );
  INV_X1 U23626 ( .A(n20738), .ZN(n20735) );
  NOR2_X1 U23627 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20735), .ZN(
        n20728) );
  AND2_X1 U23628 ( .A1(n13856), .A2(n13542), .ZN(n20805) );
  AOI21_X1 U23629 ( .B1(n20805), .B2(n14392), .A(n20728), .ZN(n20710) );
  INV_X1 U23630 ( .A(n20706), .ZN(n20707) );
  OAI22_X1 U23631 ( .A1(n20710), .A2(n20880), .B1(n20708), .B2(n20707), .ZN(
        n20727) );
  AOI22_X1 U23632 ( .A1(n20883), .A2(n20728), .B1(n20882), .B2(n20727), .ZN(
        n20714) );
  INV_X1 U23633 ( .A(n20763), .ZN(n20709) );
  OAI21_X1 U23634 ( .B1(n20709), .B2(n20729), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20711) );
  NAND2_X1 U23635 ( .A1(n20711), .A2(n20710), .ZN(n20712) );
  AOI22_X1 U23636 ( .A1(n20730), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n20849), .B2(n20729), .ZN(n20713) );
  OAI211_X1 U23637 ( .C1(n20852), .C2(n20763), .A(n20714), .B(n20713), .ZN(
        P1_U3097) );
  AOI22_X1 U23638 ( .A1(n20894), .A2(n20728), .B1(n20893), .B2(n20727), .ZN(
        n20716) );
  AOI22_X1 U23639 ( .A1(n20730), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n20895), .B2(n20729), .ZN(n20715) );
  OAI211_X1 U23640 ( .C1(n20898), .C2(n20763), .A(n20716), .B(n20715), .ZN(
        P1_U3098) );
  AOI22_X1 U23641 ( .A1(n20900), .A2(n20728), .B1(n20899), .B2(n20727), .ZN(
        n20718) );
  AOI22_X1 U23642 ( .A1(n20730), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n20901), .B2(n20729), .ZN(n20717) );
  OAI211_X1 U23643 ( .C1(n20904), .C2(n20763), .A(n20718), .B(n20717), .ZN(
        P1_U3099) );
  AOI22_X1 U23644 ( .A1(n20906), .A2(n20728), .B1(n20905), .B2(n20727), .ZN(
        n20720) );
  AOI22_X1 U23645 ( .A1(n20730), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n20907), .B2(n20729), .ZN(n20719) );
  OAI211_X1 U23646 ( .C1(n20910), .C2(n20763), .A(n20720), .B(n20719), .ZN(
        P1_U3100) );
  AOI22_X1 U23647 ( .A1(n20912), .A2(n20728), .B1(n20911), .B2(n20727), .ZN(
        n20722) );
  AOI22_X1 U23648 ( .A1(n20730), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n20859), .B2(n20729), .ZN(n20721) );
  OAI211_X1 U23649 ( .C1(n20862), .C2(n20763), .A(n20722), .B(n20721), .ZN(
        P1_U3101) );
  AOI22_X1 U23650 ( .A1(n20918), .A2(n20728), .B1(n20917), .B2(n20727), .ZN(
        n20724) );
  AOI22_X1 U23651 ( .A1(n20730), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n20919), .B2(n20729), .ZN(n20723) );
  OAI211_X1 U23652 ( .C1(n20922), .C2(n20763), .A(n20724), .B(n20723), .ZN(
        P1_U3102) );
  AOI22_X1 U23653 ( .A1(n20924), .A2(n20728), .B1(n20923), .B2(n20727), .ZN(
        n20726) );
  AOI22_X1 U23654 ( .A1(n20730), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n20865), .B2(n20729), .ZN(n20725) );
  OAI211_X1 U23655 ( .C1(n20868), .C2(n20763), .A(n20726), .B(n20725), .ZN(
        P1_U3103) );
  AOI22_X1 U23656 ( .A1(n20934), .A2(n20728), .B1(n20932), .B2(n20727), .ZN(
        n20732) );
  AOI22_X1 U23657 ( .A1(n20730), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n20935), .B2(n20729), .ZN(n20731) );
  OAI211_X1 U23658 ( .C1(n20941), .C2(n20763), .A(n20732), .B(n20731), .ZN(
        P1_U3104) );
  NOR2_X1 U23659 ( .A1(n20733), .A2(n20735), .ZN(n20759) );
  AOI21_X1 U23660 ( .B1(n20805), .B2(n20734), .A(n20759), .ZN(n20736) );
  OAI22_X1 U23661 ( .A1(n20736), .A2(n20880), .B1(n20735), .B2(n12006), .ZN(
        n20758) );
  AOI22_X1 U23662 ( .A1(n20883), .A2(n20759), .B1(n20882), .B2(n20758), .ZN(
        n20741) );
  OAI211_X1 U23663 ( .C1(n20812), .C2(n21170), .A(n20811), .B(n20736), .ZN(
        n20737) );
  OAI211_X1 U23664 ( .C1(n20811), .C2(n20738), .A(n20886), .B(n20737), .ZN(
        n20760) );
  AOI22_X1 U23665 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20760), .B1(
        n20800), .B2(n20889), .ZN(n20740) );
  OAI211_X1 U23666 ( .C1(n20892), .C2(n20763), .A(n20741), .B(n20740), .ZN(
        P1_U3105) );
  AOI22_X1 U23667 ( .A1(n20894), .A2(n20759), .B1(n20893), .B2(n20758), .ZN(
        n20743) );
  AOI22_X1 U23668 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20760), .B1(
        n20800), .B2(n20781), .ZN(n20742) );
  OAI211_X1 U23669 ( .C1(n20744), .C2(n20763), .A(n20743), .B(n20742), .ZN(
        P1_U3106) );
  AOI22_X1 U23670 ( .A1(n20900), .A2(n20759), .B1(n20899), .B2(n20758), .ZN(
        n20746) );
  AOI22_X1 U23671 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20760), .B1(
        n20800), .B2(n20784), .ZN(n20745) );
  OAI211_X1 U23672 ( .C1(n20747), .C2(n20763), .A(n20746), .B(n20745), .ZN(
        P1_U3107) );
  AOI22_X1 U23673 ( .A1(n20906), .A2(n20759), .B1(n20905), .B2(n20758), .ZN(
        n20749) );
  AOI22_X1 U23674 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20760), .B1(
        n20800), .B2(n20787), .ZN(n20748) );
  OAI211_X1 U23675 ( .C1(n20750), .C2(n20763), .A(n20749), .B(n20748), .ZN(
        P1_U3108) );
  AOI22_X1 U23676 ( .A1(n20912), .A2(n20759), .B1(n20911), .B2(n20758), .ZN(
        n20752) );
  AOI22_X1 U23677 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20760), .B1(
        n20800), .B2(n20913), .ZN(n20751) );
  OAI211_X1 U23678 ( .C1(n20916), .C2(n20763), .A(n20752), .B(n20751), .ZN(
        P1_U3109) );
  AOI22_X1 U23679 ( .A1(n20918), .A2(n20759), .B1(n20917), .B2(n20758), .ZN(
        n20754) );
  AOI22_X1 U23680 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20760), .B1(
        n20800), .B2(n20792), .ZN(n20753) );
  OAI211_X1 U23681 ( .C1(n20755), .C2(n20763), .A(n20754), .B(n20753), .ZN(
        P1_U3110) );
  AOI22_X1 U23682 ( .A1(n20924), .A2(n20759), .B1(n20923), .B2(n20758), .ZN(
        n20757) );
  AOI22_X1 U23683 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20760), .B1(
        n20800), .B2(n20925), .ZN(n20756) );
  OAI211_X1 U23684 ( .C1(n20930), .C2(n20763), .A(n20757), .B(n20756), .ZN(
        P1_U3111) );
  AOI22_X1 U23685 ( .A1(n20934), .A2(n20759), .B1(n20932), .B2(n20758), .ZN(
        n20762) );
  AOI22_X1 U23686 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20760), .B1(
        n20800), .B2(n20799), .ZN(n20761) );
  OAI211_X1 U23687 ( .C1(n20764), .C2(n20763), .A(n20762), .B(n20761), .ZN(
        P1_U3112) );
  INV_X1 U23688 ( .A(n20800), .ZN(n20765) );
  NAND2_X1 U23689 ( .A1(n20765), .A2(n20811), .ZN(n20767) );
  OAI21_X1 U23690 ( .B1(n20767), .B2(n20834), .A(n20766), .ZN(n20777) );
  AND2_X1 U23691 ( .A1(n20805), .A2(n20841), .ZN(n20772) );
  OR2_X1 U23692 ( .A1(n20769), .A2(n20768), .ZN(n20842) );
  INV_X1 U23693 ( .A(n20842), .ZN(n20770) );
  NAND3_X1 U23694 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n16225), .ZN(n20814) );
  NOR2_X1 U23695 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20814), .ZN(
        n20798) );
  AOI22_X1 U23696 ( .A1(n20834), .A2(n20889), .B1(n20883), .B2(n20798), .ZN(
        n20780) );
  INV_X1 U23697 ( .A(n20772), .ZN(n20776) );
  NAND2_X1 U23698 ( .A1(n20842), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20846) );
  OAI211_X1 U23699 ( .C1(n20774), .C2(n20798), .A(n20846), .B(n20773), .ZN(
        n20775) );
  AOI21_X1 U23700 ( .B1(n20777), .B2(n20776), .A(n20775), .ZN(n20778) );
  AOI22_X1 U23701 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20801), .B1(
        n20800), .B2(n20849), .ZN(n20779) );
  OAI211_X1 U23702 ( .C1(n20804), .C2(n9680), .A(n20780), .B(n20779), .ZN(
        P1_U3113) );
  AOI22_X1 U23703 ( .A1(n20800), .A2(n20895), .B1(n20894), .B2(n20798), .ZN(
        n20783) );
  AOI22_X1 U23704 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20801), .B1(
        n20834), .B2(n20781), .ZN(n20782) );
  OAI211_X1 U23705 ( .C1(n20804), .C2(n9678), .A(n20783), .B(n20782), .ZN(
        P1_U3114) );
  AOI22_X1 U23706 ( .A1(n20800), .A2(n20901), .B1(n20900), .B2(n20798), .ZN(
        n20786) );
  AOI22_X1 U23707 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20801), .B1(
        n20834), .B2(n20784), .ZN(n20785) );
  OAI211_X1 U23708 ( .C1(n20804), .C2(n9679), .A(n20786), .B(n20785), .ZN(
        P1_U3115) );
  AOI22_X1 U23709 ( .A1(n20834), .A2(n20787), .B1(n20906), .B2(n20798), .ZN(
        n20789) );
  AOI22_X1 U23710 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20801), .B1(
        n20800), .B2(n20907), .ZN(n20788) );
  OAI211_X1 U23711 ( .C1(n20804), .C2(n9676), .A(n20789), .B(n20788), .ZN(
        P1_U3116) );
  AOI22_X1 U23712 ( .A1(n20800), .A2(n20859), .B1(n20912), .B2(n20798), .ZN(
        n20791) );
  AOI22_X1 U23713 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20801), .B1(
        n20834), .B2(n20913), .ZN(n20790) );
  OAI211_X1 U23714 ( .C1(n20804), .C2(n9677), .A(n20791), .B(n20790), .ZN(
        P1_U3117) );
  AOI22_X1 U23715 ( .A1(n20834), .A2(n20792), .B1(n20918), .B2(n20798), .ZN(
        n20794) );
  AOI22_X1 U23716 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20801), .B1(
        n20800), .B2(n20919), .ZN(n20793) );
  OAI211_X1 U23717 ( .C1(n20804), .C2(n9682), .A(n20794), .B(n20793), .ZN(
        P1_U3118) );
  AOI22_X1 U23718 ( .A1(n20800), .A2(n20865), .B1(n20924), .B2(n20798), .ZN(
        n20796) );
  AOI22_X1 U23719 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20801), .B1(
        n20834), .B2(n20925), .ZN(n20795) );
  OAI211_X1 U23720 ( .C1(n20804), .C2(n20797), .A(n20796), .B(n20795), .ZN(
        P1_U3119) );
  AOI22_X1 U23721 ( .A1(n20834), .A2(n20799), .B1(n20934), .B2(n20798), .ZN(
        n20803) );
  AOI22_X1 U23722 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20801), .B1(
        n20800), .B2(n20935), .ZN(n20802) );
  OAI211_X1 U23723 ( .C1(n20804), .C2(n9681), .A(n20803), .B(n20802), .ZN(
        P1_U3120) );
  INV_X1 U23724 ( .A(n20805), .ZN(n20807) );
  NAND2_X1 U23725 ( .A1(n20806), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20809) );
  OAI21_X1 U23726 ( .B1(n20807), .B2(n20876), .A(n20809), .ZN(n20816) );
  INV_X1 U23727 ( .A(n20816), .ZN(n20808) );
  OAI22_X1 U23728 ( .A1(n20808), .A2(n20880), .B1(n20814), .B2(n12006), .ZN(
        n20833) );
  INV_X1 U23729 ( .A(n20809), .ZN(n20832) );
  AOI22_X1 U23730 ( .A1(n20833), .A2(n20882), .B1(n20883), .B2(n20832), .ZN(
        n20819) );
  AOI21_X1 U23731 ( .B1(n20812), .B2(n20811), .A(n20810), .ZN(n20817) );
  AOI21_X1 U23732 ( .B1(n20880), .B2(n20814), .A(n20813), .ZN(n20815) );
  AOI22_X1 U23733 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20835), .B1(
        n20834), .B2(n20849), .ZN(n20818) );
  OAI211_X1 U23734 ( .C1(n20852), .C2(n20838), .A(n20819), .B(n20818), .ZN(
        P1_U3121) );
  AOI22_X1 U23735 ( .A1(n20833), .A2(n20893), .B1(n20894), .B2(n20832), .ZN(
        n20821) );
  AOI22_X1 U23736 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20835), .B1(
        n20834), .B2(n20895), .ZN(n20820) );
  OAI211_X1 U23737 ( .C1(n20898), .C2(n20838), .A(n20821), .B(n20820), .ZN(
        P1_U3122) );
  AOI22_X1 U23738 ( .A1(n20833), .A2(n20899), .B1(n20900), .B2(n20832), .ZN(
        n20823) );
  AOI22_X1 U23739 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20835), .B1(
        n20834), .B2(n20901), .ZN(n20822) );
  OAI211_X1 U23740 ( .C1(n20904), .C2(n20838), .A(n20823), .B(n20822), .ZN(
        P1_U3123) );
  AOI22_X1 U23741 ( .A1(n20833), .A2(n20905), .B1(n20906), .B2(n20832), .ZN(
        n20825) );
  AOI22_X1 U23742 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20835), .B1(
        n20834), .B2(n20907), .ZN(n20824) );
  OAI211_X1 U23743 ( .C1(n20910), .C2(n20838), .A(n20825), .B(n20824), .ZN(
        P1_U3124) );
  AOI22_X1 U23744 ( .A1(n20833), .A2(n20911), .B1(n20912), .B2(n20832), .ZN(
        n20827) );
  AOI22_X1 U23745 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20835), .B1(
        n20834), .B2(n20859), .ZN(n20826) );
  OAI211_X1 U23746 ( .C1(n20862), .C2(n20838), .A(n20827), .B(n20826), .ZN(
        P1_U3125) );
  AOI22_X1 U23747 ( .A1(n20833), .A2(n20917), .B1(n20918), .B2(n20832), .ZN(
        n20829) );
  AOI22_X1 U23748 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20835), .B1(
        n20834), .B2(n20919), .ZN(n20828) );
  OAI211_X1 U23749 ( .C1(n20922), .C2(n20838), .A(n20829), .B(n20828), .ZN(
        P1_U3126) );
  AOI22_X1 U23750 ( .A1(n20833), .A2(n20923), .B1(n20924), .B2(n20832), .ZN(
        n20831) );
  AOI22_X1 U23751 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20835), .B1(
        n20834), .B2(n20865), .ZN(n20830) );
  OAI211_X1 U23752 ( .C1(n20868), .C2(n20838), .A(n20831), .B(n20830), .ZN(
        P1_U3127) );
  AOI22_X1 U23753 ( .A1(n20833), .A2(n20932), .B1(n20934), .B2(n20832), .ZN(
        n20837) );
  AOI22_X1 U23754 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20835), .B1(
        n20834), .B2(n20935), .ZN(n20836) );
  OAI211_X1 U23755 ( .C1(n20941), .C2(n20838), .A(n20837), .B(n20836), .ZN(
        P1_U3128) );
  INV_X1 U23756 ( .A(n20887), .ZN(n20879) );
  NOR2_X1 U23757 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20879), .ZN(
        n20870) );
  INV_X1 U23758 ( .A(n20840), .ZN(n20878) );
  NAND2_X1 U23759 ( .A1(n20878), .A2(n20841), .ZN(n20844) );
  OAI22_X1 U23760 ( .A1(n20844), .A2(n20880), .B1(n20843), .B2(n20842), .ZN(
        n20869) );
  AOI22_X1 U23761 ( .A1(n20883), .A2(n20870), .B1(n20882), .B2(n20869), .ZN(
        n20851) );
  OAI21_X1 U23762 ( .B1(n20936), .B2(n20871), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20845) );
  AOI21_X1 U23763 ( .B1(n20845), .B2(n20844), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20848) );
  AOI22_X1 U23764 ( .A1(n20872), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n20849), .B2(n20871), .ZN(n20850) );
  OAI211_X1 U23765 ( .C1(n20852), .C2(n20929), .A(n20851), .B(n20850), .ZN(
        P1_U3145) );
  AOI22_X1 U23766 ( .A1(n20894), .A2(n20870), .B1(n20893), .B2(n20869), .ZN(
        n20854) );
  AOI22_X1 U23767 ( .A1(n20872), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n20871), .B2(n20895), .ZN(n20853) );
  OAI211_X1 U23768 ( .C1(n20898), .C2(n20929), .A(n20854), .B(n20853), .ZN(
        P1_U3146) );
  AOI22_X1 U23769 ( .A1(n20900), .A2(n20870), .B1(n20899), .B2(n20869), .ZN(
        n20856) );
  AOI22_X1 U23770 ( .A1(n20872), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n20871), .B2(n20901), .ZN(n20855) );
  OAI211_X1 U23771 ( .C1(n20904), .C2(n20929), .A(n20856), .B(n20855), .ZN(
        P1_U3147) );
  AOI22_X1 U23772 ( .A1(n20906), .A2(n20870), .B1(n20905), .B2(n20869), .ZN(
        n20858) );
  AOI22_X1 U23773 ( .A1(n20872), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n20871), .B2(n20907), .ZN(n20857) );
  OAI211_X1 U23774 ( .C1(n20910), .C2(n20929), .A(n20858), .B(n20857), .ZN(
        P1_U3148) );
  AOI22_X1 U23775 ( .A1(n20912), .A2(n20870), .B1(n20911), .B2(n20869), .ZN(
        n20861) );
  AOI22_X1 U23776 ( .A1(n20872), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n20859), .B2(n20871), .ZN(n20860) );
  OAI211_X1 U23777 ( .C1(n20862), .C2(n20929), .A(n20861), .B(n20860), .ZN(
        P1_U3149) );
  AOI22_X1 U23778 ( .A1(n20918), .A2(n20870), .B1(n20917), .B2(n20869), .ZN(
        n20864) );
  AOI22_X1 U23779 ( .A1(n20872), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n20871), .B2(n20919), .ZN(n20863) );
  OAI211_X1 U23780 ( .C1(n20922), .C2(n20929), .A(n20864), .B(n20863), .ZN(
        P1_U3150) );
  AOI22_X1 U23781 ( .A1(n20924), .A2(n20870), .B1(n20923), .B2(n20869), .ZN(
        n20867) );
  AOI22_X1 U23782 ( .A1(n20872), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n20871), .B2(n20865), .ZN(n20866) );
  OAI211_X1 U23783 ( .C1(n20868), .C2(n20929), .A(n20867), .B(n20866), .ZN(
        P1_U3151) );
  AOI22_X1 U23784 ( .A1(n20934), .A2(n20870), .B1(n20932), .B2(n20869), .ZN(
        n20874) );
  AOI22_X1 U23785 ( .A1(n20872), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n20871), .B2(n20935), .ZN(n20873) );
  OAI211_X1 U23786 ( .C1(n20941), .C2(n20929), .A(n20874), .B(n20873), .ZN(
        P1_U3152) );
  INV_X1 U23787 ( .A(n20875), .ZN(n20933) );
  INV_X1 U23788 ( .A(n20876), .ZN(n20877) );
  AOI21_X1 U23789 ( .B1(n20878), .B2(n20877), .A(n20933), .ZN(n20881) );
  OAI22_X1 U23790 ( .A1(n20881), .A2(n20880), .B1(n12006), .B2(n20879), .ZN(
        n20931) );
  AOI22_X1 U23791 ( .A1(n20883), .A2(n20933), .B1(n20882), .B2(n20931), .ZN(
        n20891) );
  NOR2_X1 U23792 ( .A1(n20885), .A2(n20884), .ZN(n20888) );
  OAI21_X1 U23793 ( .B1(n20888), .B2(n20887), .A(n20886), .ZN(n20937) );
  AOI22_X1 U23794 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20937), .B1(
        n20926), .B2(n20889), .ZN(n20890) );
  OAI211_X1 U23795 ( .C1(n20892), .C2(n20929), .A(n20891), .B(n20890), .ZN(
        P1_U3153) );
  AOI22_X1 U23796 ( .A1(n20894), .A2(n20933), .B1(n20893), .B2(n20931), .ZN(
        n20897) );
  AOI22_X1 U23797 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20937), .B1(
        n20936), .B2(n20895), .ZN(n20896) );
  OAI211_X1 U23798 ( .C1(n20898), .C2(n20940), .A(n20897), .B(n20896), .ZN(
        P1_U3154) );
  AOI22_X1 U23799 ( .A1(n20900), .A2(n20933), .B1(n20899), .B2(n20931), .ZN(
        n20903) );
  AOI22_X1 U23800 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20937), .B1(
        n20936), .B2(n20901), .ZN(n20902) );
  OAI211_X1 U23801 ( .C1(n20904), .C2(n20940), .A(n20903), .B(n20902), .ZN(
        P1_U3155) );
  AOI22_X1 U23802 ( .A1(n20906), .A2(n20933), .B1(n20905), .B2(n20931), .ZN(
        n20909) );
  AOI22_X1 U23803 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20937), .B1(
        n20936), .B2(n20907), .ZN(n20908) );
  OAI211_X1 U23804 ( .C1(n20910), .C2(n20940), .A(n20909), .B(n20908), .ZN(
        P1_U3156) );
  AOI22_X1 U23805 ( .A1(n20912), .A2(n20933), .B1(n20911), .B2(n20931), .ZN(
        n20915) );
  AOI22_X1 U23806 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20937), .B1(
        n20926), .B2(n20913), .ZN(n20914) );
  OAI211_X1 U23807 ( .C1(n20916), .C2(n20929), .A(n20915), .B(n20914), .ZN(
        P1_U3157) );
  AOI22_X1 U23808 ( .A1(n20918), .A2(n20933), .B1(n20917), .B2(n20931), .ZN(
        n20921) );
  AOI22_X1 U23809 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20937), .B1(
        n20936), .B2(n20919), .ZN(n20920) );
  OAI211_X1 U23810 ( .C1(n20922), .C2(n20940), .A(n20921), .B(n20920), .ZN(
        P1_U3158) );
  AOI22_X1 U23811 ( .A1(n20924), .A2(n20933), .B1(n20923), .B2(n20931), .ZN(
        n20928) );
  AOI22_X1 U23812 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20937), .B1(
        n20926), .B2(n20925), .ZN(n20927) );
  OAI211_X1 U23813 ( .C1(n20930), .C2(n20929), .A(n20928), .B(n20927), .ZN(
        P1_U3159) );
  AOI22_X1 U23814 ( .A1(n20934), .A2(n20933), .B1(n20932), .B2(n20931), .ZN(
        n20939) );
  AOI22_X1 U23815 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20937), .B1(
        n20936), .B2(n20935), .ZN(n20938) );
  OAI211_X1 U23816 ( .C1(n20941), .C2(n20940), .A(n20939), .B(n20938), .ZN(
        P1_U3160) );
  NOR2_X1 U23817 ( .A1(n21023), .A2(n20942), .ZN(n20944) );
  OAI21_X1 U23818 ( .B1(n20944), .B2(n12006), .A(n20943), .ZN(P1_U3163) );
  AND2_X1 U23819 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n21008), .ZN(
        P1_U3164) );
  AND2_X1 U23820 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n21008), .ZN(
        P1_U3165) );
  AND2_X1 U23821 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n21008), .ZN(
        P1_U3166) );
  AND2_X1 U23822 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n21008), .ZN(
        P1_U3167) );
  AND2_X1 U23823 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n21008), .ZN(
        P1_U3168) );
  AND2_X1 U23824 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n21008), .ZN(
        P1_U3169) );
  AND2_X1 U23825 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n21008), .ZN(
        P1_U3170) );
  AND2_X1 U23826 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n21008), .ZN(
        P1_U3171) );
  AND2_X1 U23827 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n21008), .ZN(
        P1_U3172) );
  AND2_X1 U23828 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n21008), .ZN(
        P1_U3173) );
  AND2_X1 U23829 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n21008), .ZN(
        P1_U3174) );
  AND2_X1 U23830 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n21008), .ZN(
        P1_U3175) );
  AND2_X1 U23831 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n21008), .ZN(
        P1_U3176) );
  AND2_X1 U23832 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n21008), .ZN(
        P1_U3177) );
  AND2_X1 U23833 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n21008), .ZN(
        P1_U3178) );
  AND2_X1 U23834 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n21008), .ZN(
        P1_U3179) );
  AND2_X1 U23835 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n21008), .ZN(
        P1_U3180) );
  AND2_X1 U23836 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n21008), .ZN(
        P1_U3181) );
  AND2_X1 U23837 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n21008), .ZN(
        P1_U3182) );
  AND2_X1 U23838 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n21008), .ZN(
        P1_U3183) );
  AND2_X1 U23839 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n21008), .ZN(
        P1_U3184) );
  AND2_X1 U23840 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n21008), .ZN(
        P1_U3185) );
  AND2_X1 U23841 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n21008), .ZN(P1_U3186) );
  AND2_X1 U23842 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n21008), .ZN(P1_U3187) );
  AND2_X1 U23843 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n21008), .ZN(P1_U3188) );
  AND2_X1 U23844 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n21008), .ZN(P1_U3189) );
  AND2_X1 U23845 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n21008), .ZN(P1_U3190) );
  AND2_X1 U23846 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n21008), .ZN(P1_U3191) );
  AND2_X1 U23847 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n21008), .ZN(P1_U3192) );
  AND2_X1 U23848 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n21008), .ZN(P1_U3193) );
  NOR2_X1 U23849 ( .A1(n21176), .A2(NA), .ZN(n20951) );
  NOR2_X1 U23850 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20947) );
  OAI22_X1 U23851 ( .A1(n20951), .A2(n20948), .B1(n20947), .B2(n20946), .ZN(
        n20949) );
  AOI21_X1 U23852 ( .B1(n21032), .B2(n20949), .A(n20959), .ZN(n20950) );
  OAI21_X1 U23853 ( .B1(n21027), .B2(n20955), .A(n20950), .ZN(P1_U3194) );
  OAI211_X1 U23854 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20951), .A(
        P1_STATE_REG_1__SCAN_IN), .B(n21018), .ZN(n20952) );
  INV_X1 U23855 ( .A(n20952), .ZN(n20953) );
  AOI221_X1 U23856 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20954), .C1(n21055), 
        .C2(n20954), .A(n20953), .ZN(n20958) );
  AOI21_X1 U23857 ( .B1(n21018), .B2(n21055), .A(n20955), .ZN(n20957) );
  OAI211_X1 U23858 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21176), .A(
        P1_STATE_REG_0__SCAN_IN), .B(HOLD), .ZN(n20956) );
  OAI22_X1 U23859 ( .A1(n20959), .A2(n20958), .B1(n20957), .B2(n20956), .ZN(
        P1_U3196) );
  OR2_X1 U23860 ( .A1(n21032), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20987) );
  NOR2_X1 U23861 ( .A1(n20960), .A2(n21032), .ZN(n20997) );
  INV_X1 U23862 ( .A(n20997), .ZN(n20984) );
  INV_X1 U23863 ( .A(n20984), .ZN(n21000) );
  AOI222_X1 U23864 ( .A1(n20999), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n21000), .ZN(n20961) );
  INV_X1 U23865 ( .A(n20961), .ZN(P1_U3197) );
  AOI222_X1 U23866 ( .A1(n21000), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20999), .ZN(n20962) );
  INV_X1 U23867 ( .A(n20962), .ZN(P1_U3198) );
  OAI222_X1 U23868 ( .A1(n20984), .A2(n13964), .B1(n20964), .B2(n21031), .C1(
        n20963), .C2(n20987), .ZN(P1_U3199) );
  AOI222_X1 U23869 ( .A1(n20999), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n21000), .ZN(n20965) );
  INV_X1 U23870 ( .A(n20965), .ZN(P1_U3200) );
  AOI222_X1 U23871 ( .A1(n21000), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20999), .ZN(n20966) );
  INV_X1 U23872 ( .A(n20966), .ZN(P1_U3201) );
  AOI222_X1 U23873 ( .A1(n21000), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20999), .ZN(n20967) );
  INV_X1 U23874 ( .A(n20967), .ZN(P1_U3202) );
  AOI222_X1 U23875 ( .A1(n21000), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20999), .ZN(n20968) );
  INV_X1 U23876 ( .A(n20968), .ZN(P1_U3203) );
  AOI222_X1 U23877 ( .A1(n21000), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n20999), .ZN(n20969) );
  INV_X1 U23878 ( .A(n20969), .ZN(P1_U3204) );
  AOI222_X1 U23879 ( .A1(n21000), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20999), .ZN(n20970) );
  INV_X1 U23880 ( .A(n20970), .ZN(P1_U3205) );
  AOI22_X1 U23881 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n21032), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n20999), .ZN(n20971) );
  OAI21_X1 U23882 ( .B1(n20972), .B2(n20984), .A(n20971), .ZN(P1_U3206) );
  AOI22_X1 U23883 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n21032), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20999), .ZN(n20973) );
  OAI21_X1 U23884 ( .B1(n20974), .B2(n20984), .A(n20973), .ZN(P1_U3207) );
  AOI22_X1 U23885 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(n21032), .B1(
        P1_REIP_REG_12__SCAN_IN), .B2(n20997), .ZN(n20975) );
  OAI21_X1 U23886 ( .B1(n20977), .B2(n20987), .A(n20975), .ZN(P1_U3208) );
  AOI22_X1 U23887 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n21032), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20999), .ZN(n20976) );
  OAI21_X1 U23888 ( .B1(n20977), .B2(n20984), .A(n20976), .ZN(P1_U3209) );
  AOI22_X1 U23889 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n21032), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n21000), .ZN(n20978) );
  OAI21_X1 U23890 ( .B1(n15253), .B2(n20987), .A(n20978), .ZN(P1_U3210) );
  AOI222_X1 U23891 ( .A1(n21000), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20999), .ZN(n20979) );
  INV_X1 U23892 ( .A(n20979), .ZN(P1_U3211) );
  AOI22_X1 U23893 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n21032), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20999), .ZN(n20980) );
  OAI21_X1 U23894 ( .B1(n20981), .B2(n20984), .A(n20980), .ZN(P1_U3212) );
  INV_X1 U23895 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20985) );
  AOI22_X1 U23896 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n21032), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n21000), .ZN(n20982) );
  OAI21_X1 U23897 ( .B1(n20985), .B2(n20987), .A(n20982), .ZN(P1_U3213) );
  AOI22_X1 U23898 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n21032), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20999), .ZN(n20983) );
  OAI21_X1 U23899 ( .B1(n20985), .B2(n20984), .A(n20983), .ZN(P1_U3214) );
  AOI22_X1 U23900 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n21032), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20997), .ZN(n20986) );
  OAI21_X1 U23901 ( .B1(n15207), .B2(n20987), .A(n20986), .ZN(P1_U3215) );
  AOI222_X1 U23902 ( .A1(n21000), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20999), .ZN(n20988) );
  INV_X1 U23903 ( .A(n20988), .ZN(P1_U3216) );
  AOI222_X1 U23904 ( .A1(n20997), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20999), .ZN(n20989) );
  INV_X1 U23905 ( .A(n20989), .ZN(P1_U3217) );
  AOI222_X1 U23906 ( .A1(n21000), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20999), .ZN(n20990) );
  INV_X1 U23907 ( .A(n20990), .ZN(P1_U3218) );
  AOI222_X1 U23908 ( .A1(n20997), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20999), .ZN(n20991) );
  INV_X1 U23909 ( .A(n20991), .ZN(P1_U3219) );
  AOI222_X1 U23910 ( .A1(n20997), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20999), .ZN(n20992) );
  INV_X1 U23911 ( .A(n20992), .ZN(P1_U3220) );
  AOI222_X1 U23912 ( .A1(n20997), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20999), .ZN(n20993) );
  INV_X1 U23913 ( .A(n20993), .ZN(P1_U3221) );
  AOI222_X1 U23914 ( .A1(n21000), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20999), .ZN(n20994) );
  INV_X1 U23915 ( .A(n20994), .ZN(P1_U3222) );
  AOI222_X1 U23916 ( .A1(n20997), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20999), .ZN(n20995) );
  INV_X1 U23917 ( .A(n20995), .ZN(P1_U3223) );
  AOI222_X1 U23918 ( .A1(n21000), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20999), .ZN(n20996) );
  INV_X1 U23919 ( .A(n20996), .ZN(P1_U3224) );
  AOI222_X1 U23920 ( .A1(n20997), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20999), .ZN(n20998) );
  INV_X1 U23921 ( .A(n20998), .ZN(P1_U3225) );
  AOI222_X1 U23922 ( .A1(n21000), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n21032), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20999), .ZN(n21001) );
  INV_X1 U23923 ( .A(n21001), .ZN(P1_U3226) );
  OAI22_X1 U23924 ( .A1(n21032), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n21031), .ZN(n21002) );
  INV_X1 U23925 ( .A(n21002), .ZN(P1_U3458) );
  OAI22_X1 U23926 ( .A1(n21032), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n21031), .ZN(n21003) );
  INV_X1 U23927 ( .A(n21003), .ZN(P1_U3459) );
  OAI22_X1 U23928 ( .A1(n21032), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n21031), .ZN(n21004) );
  INV_X1 U23929 ( .A(n21004), .ZN(P1_U3460) );
  OAI22_X1 U23930 ( .A1(n21032), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n21031), .ZN(n21005) );
  INV_X1 U23931 ( .A(n21005), .ZN(P1_U3461) );
  INV_X1 U23932 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n21011) );
  INV_X1 U23933 ( .A(n21006), .ZN(n21007) );
  AOI21_X1 U23934 ( .B1(n21011), .B2(n21008), .A(n21007), .ZN(P1_U3464) );
  AOI21_X1 U23935 ( .B1(n21008), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n21007), 
        .ZN(n21009) );
  INV_X1 U23936 ( .A(n21009), .ZN(P1_U3465) );
  NOR3_X1 U23937 ( .A1(n21011), .A2(P1_REIP_REG_0__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .ZN(n21010) );
  AOI221_X1 U23938 ( .B1(n21012), .B2(n21011), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n21010), .ZN(n21014) );
  INV_X1 U23939 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21013) );
  INV_X1 U23940 ( .A(n21017), .ZN(n21015) );
  AOI22_X1 U23941 ( .A1(n21017), .A2(n21014), .B1(n21013), .B2(n21015), .ZN(
        P1_U3481) );
  NOR2_X1 U23942 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n21016) );
  INV_X1 U23943 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n21054) );
  AOI22_X1 U23944 ( .A1(n21017), .A2(n21016), .B1(n21054), .B2(n21015), .ZN(
        P1_U3482) );
  AOI22_X1 U23945 ( .A1(n21031), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n21092), 
        .B2(n21032), .ZN(P1_U3483) );
  AOI211_X1 U23946 ( .C1(n21019), .C2(n21170), .A(n12006), .B(n21018), .ZN(
        n21021) );
  AND2_X1 U23947 ( .A1(n21021), .A2(n21020), .ZN(n21024) );
  OAI21_X1 U23948 ( .B1(n21024), .B2(n21023), .A(n21022), .ZN(n21030) );
  AOI211_X1 U23949 ( .C1(n21028), .C2(n21027), .A(n21026), .B(n21025), .ZN(
        n21029) );
  MUX2_X1 U23950 ( .A(n21030), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n21029), 
        .Z(P1_U3485) );
  OAI22_X1 U23951 ( .A1(n21032), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n21031), .ZN(n21033) );
  INV_X1 U23952 ( .A(n21033), .ZN(P1_U3486) );
  INV_X1 U23953 ( .A(keyinput_f21), .ZN(n21128) );
  AOI22_X1 U23954 ( .A1(n21036), .A2(keyinput_f15), .B1(n21035), .B2(
        keyinput_f10), .ZN(n21034) );
  OAI221_X1 U23955 ( .B1(n21036), .B2(keyinput_f15), .C1(n21035), .C2(
        keyinput_f10), .A(n21034), .ZN(n21126) );
  INV_X1 U23956 ( .A(READY2), .ZN(n21039) );
  AOI22_X1 U23957 ( .A1(n21039), .A2(keyinput_f37), .B1(n21038), .B2(
        keyinput_f55), .ZN(n21037) );
  OAI221_X1 U23958 ( .B1(n21039), .B2(keyinput_f37), .C1(n21038), .C2(
        keyinput_f55), .A(n21037), .ZN(n21125) );
  INV_X1 U23959 ( .A(keyinput_f35), .ZN(n21041) );
  OAI22_X1 U23960 ( .A1(n21042), .A2(keyinput_f13), .B1(n21041), .B2(BS16), 
        .ZN(n21040) );
  AOI221_X1 U23961 ( .B1(n21042), .B2(keyinput_f13), .C1(BS16), .C2(n21041), 
        .A(n21040), .ZN(n21059) );
  INV_X1 U23962 ( .A(keyinput_f50), .ZN(n21044) );
  AOI22_X1 U23963 ( .A1(n21171), .A2(keyinput_f12), .B1(
        P1_BYTEENABLE_REG_2__SCAN_IN), .B2(n21044), .ZN(n21043) );
  OAI221_X1 U23964 ( .B1(n21171), .B2(keyinput_f12), .C1(n21044), .C2(
        P1_BYTEENABLE_REG_2__SCAN_IN), .A(n21043), .ZN(n21053) );
  INV_X1 U23965 ( .A(DATAI_1_), .ZN(n21046) );
  AOI22_X1 U23966 ( .A1(n21047), .A2(keyinput_f59), .B1(keyinput_f31), .B2(
        n21046), .ZN(n21045) );
  OAI221_X1 U23967 ( .B1(n21047), .B2(keyinput_f59), .C1(n21046), .C2(
        keyinput_f31), .A(n21045), .ZN(n21052) );
  AOI22_X1 U23968 ( .A1(n21193), .A2(keyinput_f11), .B1(n21138), .B2(
        keyinput_f4), .ZN(n21048) );
  OAI221_X1 U23969 ( .B1(n21193), .B2(keyinput_f11), .C1(n21138), .C2(
        keyinput_f4), .A(n21048), .ZN(n21051) );
  AOI22_X1 U23970 ( .A1(n21173), .A2(keyinput_f39), .B1(n21209), .B2(
        keyinput_f5), .ZN(n21049) );
  OAI221_X1 U23971 ( .B1(n21173), .B2(keyinput_f39), .C1(n21209), .C2(
        keyinput_f5), .A(n21049), .ZN(n21050) );
  NOR4_X1 U23972 ( .A1(n21053), .A2(n21052), .A3(n21051), .A4(n21050), .ZN(
        n21058) );
  XOR2_X1 U23973 ( .A(keyinput_f48), .B(n21054), .Z(n21057) );
  XOR2_X1 U23974 ( .A(keyinput_f34), .B(n21055), .Z(n21056) );
  NAND4_X1 U23975 ( .A1(n21059), .A2(n21058), .A3(n21057), .A4(n21056), .ZN(
        n21124) );
  OAI22_X1 U23976 ( .A1(DATAI_26_), .A2(keyinput_f6), .B1(HOLD), .B2(
        keyinput_f33), .ZN(n21060) );
  AOI221_X1 U23977 ( .B1(DATAI_26_), .B2(keyinput_f6), .C1(keyinput_f33), .C2(
        HOLD), .A(n21060), .ZN(n21122) );
  OAI22_X1 U23978 ( .A1(DATAI_24_), .A2(keyinput_f8), .B1(DATAI_8_), .B2(
        keyinput_f24), .ZN(n21061) );
  AOI221_X1 U23979 ( .B1(DATAI_24_), .B2(keyinput_f8), .C1(keyinput_f24), .C2(
        DATAI_8_), .A(n21061), .ZN(n21121) );
  AOI22_X1 U23980 ( .A1(DATAI_9_), .A2(keyinput_f23), .B1(DATAI_25_), .B2(
        keyinput_f7), .ZN(n21062) );
  OAI221_X1 U23981 ( .B1(DATAI_9_), .B2(keyinput_f23), .C1(DATAI_25_), .C2(
        keyinput_f7), .A(n21062), .ZN(n21069) );
  AOI22_X1 U23982 ( .A1(keyinput_f42), .A2(P1_D_C_N_REG_SCAN_IN), .B1(
        DATAI_31_), .B2(keyinput_f1), .ZN(n21063) );
  OAI221_X1 U23983 ( .B1(keyinput_f42), .B2(P1_D_C_N_REG_SCAN_IN), .C1(
        DATAI_31_), .C2(keyinput_f1), .A(n21063), .ZN(n21068) );
  AOI22_X1 U23984 ( .A1(P1_READREQUEST_REG_SCAN_IN), .A2(keyinput_f38), .B1(
        READY1), .B2(keyinput_f36), .ZN(n21064) );
  OAI221_X1 U23985 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_f38), .C1(
        READY1), .C2(keyinput_f36), .A(n21064), .ZN(n21067) );
  AOI22_X1 U23986 ( .A1(DATAI_15_), .A2(keyinput_f17), .B1(DATAI_16_), .B2(
        keyinput_f16), .ZN(n21065) );
  OAI221_X1 U23987 ( .B1(DATAI_15_), .B2(keyinput_f17), .C1(DATAI_16_), .C2(
        keyinput_f16), .A(n21065), .ZN(n21066) );
  NOR4_X1 U23988 ( .A1(n21069), .A2(n21068), .A3(n21067), .A4(n21066), .ZN(
        n21073) );
  OAI22_X1 U23989 ( .A1(n21071), .A2(keyinput_f20), .B1(keyinput_f27), .B2(
        DATAI_5_), .ZN(n21070) );
  AOI221_X1 U23990 ( .B1(n21071), .B2(keyinput_f20), .C1(DATAI_5_), .C2(
        keyinput_f27), .A(n21070), .ZN(n21072) );
  OAI211_X1 U23991 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(keyinput_f44), .A(
        n21073), .B(n21072), .ZN(n21074) );
  AOI21_X1 U23992 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_f44), .A(
        n21074), .ZN(n21120) );
  OAI22_X1 U23993 ( .A1(DATAI_30_), .A2(keyinput_f2), .B1(DATAI_4_), .B2(
        keyinput_f28), .ZN(n21075) );
  AOI221_X1 U23994 ( .B1(DATAI_30_), .B2(keyinput_f2), .C1(keyinput_f28), .C2(
        DATAI_4_), .A(n21075), .ZN(n21082) );
  OAI22_X1 U23995 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(keyinput_f63), .B1(
        DATAI_10_), .B2(keyinput_f22), .ZN(n21076) );
  AOI221_X1 U23996 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(keyinput_f63), .C1(
        keyinput_f22), .C2(DATAI_10_), .A(n21076), .ZN(n21081) );
  INV_X1 U23997 ( .A(DATAI_2_), .ZN(n21211) );
  OAI22_X1 U23998 ( .A1(n21211), .A2(keyinput_f30), .B1(keyinput_f9), .B2(
        DATAI_23_), .ZN(n21077) );
  AOI221_X1 U23999 ( .B1(n21211), .B2(keyinput_f30), .C1(DATAI_23_), .C2(
        keyinput_f9), .A(n21077), .ZN(n21080) );
  OAI22_X1 U24000 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(keyinput_f62), .B1(
        keyinput_f0), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n21078) );
  AOI221_X1 U24001 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_f62), .C1(
        P1_MEMORYFETCH_REG_SCAN_IN), .C2(keyinput_f0), .A(n21078), .ZN(n21079)
         );
  NAND4_X1 U24002 ( .A1(n21082), .A2(n21081), .A3(n21080), .A4(n21079), .ZN(
        n21118) );
  OAI22_X1 U24003 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(keyinput_f56), .B1(
        keyinput_f40), .B2(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21083) );
  AOI221_X1 U24004 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(keyinput_f56), .C1(
        P1_CODEFETCH_REG_SCAN_IN), .C2(keyinput_f40), .A(n21083), .ZN(n21090)
         );
  OAI22_X1 U24005 ( .A1(DATAI_13_), .A2(keyinput_f19), .B1(keyinput_f51), .B2(
        P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n21084) );
  AOI221_X1 U24006 ( .B1(DATAI_13_), .B2(keyinput_f19), .C1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .C2(keyinput_f51), .A(n21084), .ZN(
        n21089) );
  OAI22_X1 U24007 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(keyinput_f61), .B1(
        P1_FLUSH_REG_SCAN_IN), .B2(keyinput_f46), .ZN(n21085) );
  AOI221_X1 U24008 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput_f61), .C1(
        keyinput_f46), .C2(P1_FLUSH_REG_SCAN_IN), .A(n21085), .ZN(n21088) );
  OAI22_X1 U24009 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_f57), .B1(
        DATAI_14_), .B2(keyinput_f18), .ZN(n21086) );
  AOI221_X1 U24010 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_f57), .C1(
        keyinput_f18), .C2(DATAI_14_), .A(n21086), .ZN(n21087) );
  NAND4_X1 U24011 ( .A1(n21090), .A2(n21089), .A3(n21088), .A4(n21087), .ZN(
        n21117) );
  OAI22_X1 U24012 ( .A1(n21093), .A2(keyinput_f60), .B1(n21092), .B2(
        keyinput_f47), .ZN(n21091) );
  AOI221_X1 U24013 ( .B1(n21093), .B2(keyinput_f60), .C1(keyinput_f47), .C2(
        n21092), .A(n21091), .ZN(n21102) );
  INV_X1 U24014 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n21174) );
  OAI22_X1 U24015 ( .A1(n21174), .A2(keyinput_f58), .B1(n21176), .B2(
        keyinput_f43), .ZN(n21094) );
  AOI221_X1 U24016 ( .B1(n21174), .B2(keyinput_f58), .C1(keyinput_f43), .C2(
        n21176), .A(n21094), .ZN(n21101) );
  INV_X1 U24017 ( .A(DATAI_0_), .ZN(n21208) );
  OAI22_X1 U24018 ( .A1(n21096), .A2(keyinput_f54), .B1(n21208), .B2(
        keyinput_f32), .ZN(n21095) );
  AOI221_X1 U24019 ( .B1(n21096), .B2(keyinput_f54), .C1(keyinput_f32), .C2(
        n21208), .A(n21095), .ZN(n21100) );
  INV_X1 U24020 ( .A(DATAI_3_), .ZN(n21098) );
  OAI22_X1 U24021 ( .A1(n13779), .A2(keyinput_f26), .B1(n21098), .B2(
        keyinput_f29), .ZN(n21097) );
  AOI221_X1 U24022 ( .B1(n13779), .B2(keyinput_f26), .C1(keyinput_f29), .C2(
        n21098), .A(n21097), .ZN(n21099) );
  NAND4_X1 U24023 ( .A1(n21102), .A2(n21101), .A3(n21100), .A4(n21099), .ZN(
        n21116) );
  OAI22_X1 U24024 ( .A1(n21201), .A2(keyinput_f3), .B1(n13792), .B2(
        keyinput_f25), .ZN(n21103) );
  AOI221_X1 U24025 ( .B1(n21201), .B2(keyinput_f3), .C1(keyinput_f25), .C2(
        n13792), .A(n21103), .ZN(n21114) );
  INV_X1 U24026 ( .A(keyinput_f41), .ZN(n21105) );
  OAI22_X1 U24027 ( .A1(n21106), .A2(keyinput_f45), .B1(n21105), .B2(
        P1_M_IO_N_REG_SCAN_IN), .ZN(n21104) );
  AOI221_X1 U24028 ( .B1(n21106), .B2(keyinput_f45), .C1(P1_M_IO_N_REG_SCAN_IN), .C2(n21105), .A(n21104), .ZN(n21113) );
  OAI22_X1 U24029 ( .A1(n21185), .A2(keyinput_f52), .B1(n21108), .B2(
        keyinput_f53), .ZN(n21107) );
  AOI221_X1 U24030 ( .B1(n21185), .B2(keyinput_f52), .C1(keyinput_f53), .C2(
        n21108), .A(n21107), .ZN(n21112) );
  INV_X1 U24031 ( .A(keyinput_f49), .ZN(n21110) );
  OAI22_X1 U24032 ( .A1(n21198), .A2(keyinput_f14), .B1(n21110), .B2(
        P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n21109) );
  AOI221_X1 U24033 ( .B1(n21198), .B2(keyinput_f14), .C1(
        P1_BYTEENABLE_REG_1__SCAN_IN), .C2(n21110), .A(n21109), .ZN(n21111) );
  NAND4_X1 U24034 ( .A1(n21114), .A2(n21113), .A3(n21112), .A4(n21111), .ZN(
        n21115) );
  NOR4_X1 U24035 ( .A1(n21118), .A2(n21117), .A3(n21116), .A4(n21115), .ZN(
        n21119) );
  NAND4_X1 U24036 ( .A1(n21122), .A2(n21121), .A3(n21120), .A4(n21119), .ZN(
        n21123) );
  NOR4_X1 U24037 ( .A1(n21126), .A2(n21125), .A3(n21124), .A4(n21123), .ZN(
        n21127) );
  AOI221_X1 U24038 ( .B1(DATAI_11_), .B2(keyinput_f21), .C1(n21129), .C2(
        n21128), .A(n21127), .ZN(n21230) );
  AOI22_X1 U24039 ( .A1(P1_BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput_g51), .B1(
        DATAI_25_), .B2(keyinput_g7), .ZN(n21130) );
  OAI221_X1 U24040 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_g51), 
        .C1(DATAI_25_), .C2(keyinput_g7), .A(n21130), .ZN(n21137) );
  AOI22_X1 U24041 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(keyinput_g61), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(keyinput_g59), .ZN(n21131) );
  OAI221_X1 U24042 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(keyinput_g61), .C1(
        P1_REIP_REG_24__SCAN_IN), .C2(keyinput_g59), .A(n21131), .ZN(n21136)
         );
  AOI22_X1 U24043 ( .A1(P1_BYTEENABLE_REG_0__SCAN_IN), .A2(keyinput_g48), .B1(
        HOLD), .B2(keyinput_g33), .ZN(n21132) );
  OAI221_X1 U24044 ( .B1(P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_g48), 
        .C1(HOLD), .C2(keyinput_g33), .A(n21132), .ZN(n21135) );
  AOI22_X1 U24045 ( .A1(DATAI_19_), .A2(keyinput_g13), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(keyinput_g60), .ZN(n21133) );
  OAI221_X1 U24046 ( .B1(DATAI_19_), .B2(keyinput_g13), .C1(
        P1_REIP_REG_23__SCAN_IN), .C2(keyinput_g60), .A(n21133), .ZN(n21134)
         );
  NOR4_X1 U24047 ( .A1(n21137), .A2(n21136), .A3(n21135), .A4(n21134), .ZN(
        n21166) );
  XOR2_X1 U24048 ( .A(n21138), .B(keyinput_g4), .Z(n21146) );
  AOI22_X1 U24049 ( .A1(DATAI_30_), .A2(keyinput_g2), .B1(n21140), .B2(
        keyinput_g1), .ZN(n21139) );
  OAI221_X1 U24050 ( .B1(DATAI_30_), .B2(keyinput_g2), .C1(n21140), .C2(
        keyinput_g1), .A(n21139), .ZN(n21145) );
  AOI22_X1 U24051 ( .A1(P1_W_R_N_REG_SCAN_IN), .A2(keyinput_g47), .B1(DATAI_1_), .B2(keyinput_g31), .ZN(n21141) );
  OAI221_X1 U24052 ( .B1(P1_W_R_N_REG_SCAN_IN), .B2(keyinput_g47), .C1(
        DATAI_1_), .C2(keyinput_g31), .A(n21141), .ZN(n21144) );
  AOI22_X1 U24053 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_g57), .B1(
        P1_REIP_REG_28__SCAN_IN), .B2(keyinput_g55), .ZN(n21142) );
  OAI221_X1 U24054 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_g57), .C1(
        P1_REIP_REG_28__SCAN_IN), .C2(keyinput_g55), .A(n21142), .ZN(n21143)
         );
  NOR4_X1 U24055 ( .A1(n21146), .A2(n21145), .A3(n21144), .A4(n21143), .ZN(
        n21165) );
  AOI22_X1 U24056 ( .A1(READY2), .A2(keyinput_g37), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(keyinput_g62), .ZN(n21147) );
  OAI221_X1 U24057 ( .B1(READY2), .B2(keyinput_g37), .C1(
        P1_REIP_REG_21__SCAN_IN), .C2(keyinput_g62), .A(n21147), .ZN(n21154)
         );
  AOI22_X1 U24058 ( .A1(P1_BYTEENABLE_REG_1__SCAN_IN), .A2(keyinput_g49), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(keyinput_g41), .ZN(n21148) );
  OAI221_X1 U24059 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(keyinput_g49), 
        .C1(P1_M_IO_N_REG_SCAN_IN), .C2(keyinput_g41), .A(n21148), .ZN(n21153)
         );
  AOI22_X1 U24060 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput_g42), .B1(
        P1_READREQUEST_REG_SCAN_IN), .B2(keyinput_g38), .ZN(n21149) );
  OAI221_X1 U24061 ( .B1(P1_D_C_N_REG_SCAN_IN), .B2(keyinput_g42), .C1(
        P1_READREQUEST_REG_SCAN_IN), .C2(keyinput_g38), .A(n21149), .ZN(n21152) );
  AOI22_X1 U24062 ( .A1(P1_BYTEENABLE_REG_2__SCAN_IN), .A2(keyinput_g50), .B1(
        P1_REIP_REG_29__SCAN_IN), .B2(keyinput_g54), .ZN(n21150) );
  OAI221_X1 U24063 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_g50), 
        .C1(P1_REIP_REG_29__SCAN_IN), .C2(keyinput_g54), .A(n21150), .ZN(
        n21151) );
  NOR4_X1 U24064 ( .A1(n21154), .A2(n21153), .A3(n21152), .A4(n21151), .ZN(
        n21164) );
  AOI22_X1 U24065 ( .A1(DATAI_7_), .A2(keyinput_g25), .B1(DATAI_13_), .B2(
        keyinput_g19), .ZN(n21155) );
  OAI221_X1 U24066 ( .B1(DATAI_7_), .B2(keyinput_g25), .C1(DATAI_13_), .C2(
        keyinput_g19), .A(n21155), .ZN(n21162) );
  AOI22_X1 U24067 ( .A1(DATAI_3_), .A2(keyinput_g29), .B1(DATAI_23_), .B2(
        keyinput_g9), .ZN(n21156) );
  OAI221_X1 U24068 ( .B1(DATAI_3_), .B2(keyinput_g29), .C1(DATAI_23_), .C2(
        keyinput_g9), .A(n21156), .ZN(n21161) );
  AOI22_X1 U24069 ( .A1(P1_MORE_REG_SCAN_IN), .A2(keyinput_g45), .B1(DATAI_24_), .B2(keyinput_g8), .ZN(n21157) );
  OAI221_X1 U24070 ( .B1(P1_MORE_REG_SCAN_IN), .B2(keyinput_g45), .C1(
        DATAI_24_), .C2(keyinput_g8), .A(n21157), .ZN(n21160) );
  AOI22_X1 U24071 ( .A1(DATAI_17_), .A2(keyinput_g15), .B1(DATAI_10_), .B2(
        keyinput_g22), .ZN(n21158) );
  OAI221_X1 U24072 ( .B1(DATAI_17_), .B2(keyinput_g15), .C1(DATAI_10_), .C2(
        keyinput_g22), .A(n21158), .ZN(n21159) );
  NOR4_X1 U24073 ( .A1(n21162), .A2(n21161), .A3(n21160), .A4(n21159), .ZN(
        n21163) );
  NAND4_X1 U24074 ( .A1(n21166), .A2(n21165), .A3(n21164), .A4(n21163), .ZN(
        n21228) );
  AOI22_X1 U24075 ( .A1(n21168), .A2(keyinput_g23), .B1(keyinput_g0), .B2(
        n13458), .ZN(n21167) );
  OAI221_X1 U24076 ( .B1(n21168), .B2(keyinput_g23), .C1(n13458), .C2(
        keyinput_g0), .A(n21167), .ZN(n21181) );
  AOI22_X1 U24077 ( .A1(n21171), .A2(keyinput_g12), .B1(n21170), .B2(
        keyinput_g44), .ZN(n21169) );
  OAI221_X1 U24078 ( .B1(n21171), .B2(keyinput_g12), .C1(n21170), .C2(
        keyinput_g44), .A(n21169), .ZN(n21180) );
  AOI22_X1 U24079 ( .A1(n21174), .A2(keyinput_g58), .B1(keyinput_g39), .B2(
        n21173), .ZN(n21172) );
  OAI221_X1 U24080 ( .B1(n21174), .B2(keyinput_g58), .C1(n21173), .C2(
        keyinput_g39), .A(n21172), .ZN(n21179) );
  AOI22_X1 U24081 ( .A1(n21177), .A2(keyinput_g6), .B1(keyinput_g43), .B2(
        n21176), .ZN(n21175) );
  OAI221_X1 U24082 ( .B1(n21177), .B2(keyinput_g6), .C1(n21176), .C2(
        keyinput_g43), .A(n21175), .ZN(n21178) );
  NOR4_X1 U24083 ( .A1(n21181), .A2(n21180), .A3(n21179), .A4(n21178), .ZN(
        n21226) );
  AOI22_X1 U24084 ( .A1(NA), .A2(keyinput_g34), .B1(P1_REIP_REG_30__SCAN_IN), 
        .B2(keyinput_g53), .ZN(n21182) );
  OAI221_X1 U24085 ( .B1(NA), .B2(keyinput_g34), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(keyinput_g53), .A(n21182), .ZN(n21191) );
  AOI22_X1 U24086 ( .A1(DATAI_6_), .A2(keyinput_g26), .B1(DATAI_12_), .B2(
        keyinput_g20), .ZN(n21183) );
  OAI221_X1 U24087 ( .B1(DATAI_6_), .B2(keyinput_g26), .C1(DATAI_12_), .C2(
        keyinput_g20), .A(n21183), .ZN(n21190) );
  AOI22_X1 U24088 ( .A1(n21185), .A2(keyinput_g52), .B1(keyinput_g63), .B2(
        n15207), .ZN(n21184) );
  OAI221_X1 U24089 ( .B1(n21185), .B2(keyinput_g52), .C1(n15207), .C2(
        keyinput_g63), .A(n21184), .ZN(n21189) );
  AOI22_X1 U24090 ( .A1(DATAI_22_), .A2(keyinput_g10), .B1(n21187), .B2(
        keyinput_g16), .ZN(n21186) );
  OAI221_X1 U24091 ( .B1(DATAI_22_), .B2(keyinput_g10), .C1(n21187), .C2(
        keyinput_g16), .A(n21186), .ZN(n21188) );
  NOR4_X1 U24092 ( .A1(n21191), .A2(n21190), .A3(n21189), .A4(n21188), .ZN(
        n21225) );
  AOI22_X1 U24093 ( .A1(n21194), .A2(keyinput_g40), .B1(n21193), .B2(
        keyinput_g11), .ZN(n21192) );
  OAI221_X1 U24094 ( .B1(n21194), .B2(keyinput_g40), .C1(n21193), .C2(
        keyinput_g11), .A(n21192), .ZN(n21206) );
  INV_X1 U24095 ( .A(DATAI_4_), .ZN(n21196) );
  AOI22_X1 U24096 ( .A1(n21196), .A2(keyinput_g28), .B1(keyinput_g17), .B2(
        n13661), .ZN(n21195) );
  OAI221_X1 U24097 ( .B1(n21196), .B2(keyinput_g28), .C1(n13661), .C2(
        keyinput_g17), .A(n21195), .ZN(n21205) );
  AOI22_X1 U24098 ( .A1(n21199), .A2(keyinput_g56), .B1(keyinput_g14), .B2(
        n21198), .ZN(n21197) );
  OAI221_X1 U24099 ( .B1(n21199), .B2(keyinput_g56), .C1(n21198), .C2(
        keyinput_g14), .A(n21197), .ZN(n21204) );
  AOI22_X1 U24100 ( .A1(n21202), .A2(keyinput_g24), .B1(n21201), .B2(
        keyinput_g3), .ZN(n21200) );
  OAI221_X1 U24101 ( .B1(n21202), .B2(keyinput_g24), .C1(n21201), .C2(
        keyinput_g3), .A(n21200), .ZN(n21203) );
  NOR4_X1 U24102 ( .A1(n21206), .A2(n21205), .A3(n21204), .A4(n21203), .ZN(
        n21224) );
  AOI22_X1 U24103 ( .A1(n21209), .A2(keyinput_g5), .B1(keyinput_g32), .B2(
        n21208), .ZN(n21207) );
  OAI221_X1 U24104 ( .B1(n21209), .B2(keyinput_g5), .C1(n21208), .C2(
        keyinput_g32), .A(n21207), .ZN(n21222) );
  AOI22_X1 U24105 ( .A1(n21212), .A2(keyinput_g46), .B1(n21211), .B2(
        keyinput_g30), .ZN(n21210) );
  OAI221_X1 U24106 ( .B1(n21212), .B2(keyinput_g46), .C1(n21211), .C2(
        keyinput_g30), .A(n21210), .ZN(n21221) );
  INV_X1 U24107 ( .A(READY1), .ZN(n21215) );
  INV_X1 U24108 ( .A(DATAI_5_), .ZN(n21214) );
  AOI22_X1 U24109 ( .A1(n21215), .A2(keyinput_g36), .B1(keyinput_g27), .B2(
        n21214), .ZN(n21213) );
  OAI221_X1 U24110 ( .B1(n21215), .B2(keyinput_g36), .C1(n21214), .C2(
        keyinput_g27), .A(n21213), .ZN(n21220) );
  INV_X1 U24111 ( .A(BS16), .ZN(n21218) );
  AOI22_X1 U24112 ( .A1(n21218), .A2(keyinput_g35), .B1(n21217), .B2(
        keyinput_g18), .ZN(n21216) );
  OAI221_X1 U24113 ( .B1(n21218), .B2(keyinput_g35), .C1(n21217), .C2(
        keyinput_g18), .A(n21216), .ZN(n21219) );
  NOR4_X1 U24114 ( .A1(n21222), .A2(n21221), .A3(n21220), .A4(n21219), .ZN(
        n21223) );
  NAND4_X1 U24115 ( .A1(n21226), .A2(n21225), .A3(n21224), .A4(n21223), .ZN(
        n21227) );
  OAI22_X1 U24116 ( .A1(DATAI_11_), .A2(keyinput_g21), .B1(n21228), .B2(n21227), .ZN(n21229) );
  AOI211_X1 U24117 ( .C1(DATAI_11_), .C2(keyinput_g21), .A(n21230), .B(n21229), 
        .ZN(n21232) );
  AOI22_X1 U24118 ( .A1(n16846), .A2(P3_ADDRESS_REG_29__SCAN_IN), .B1(
        P2_ADDRESS_REG_29__SCAN_IN), .B2(n16848), .ZN(n21231) );
  XNOR2_X1 U24119 ( .A(n21232), .B(n21231), .ZN(U355) );
  NOR2_X1 U11245 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10369) );
  INV_X1 U11517 ( .A(n10099), .ZN(n12929) );
  NAND2_X1 U15299 ( .A1(n12015), .A2(n11975), .ZN(n12033) );
  AND2_X1 U11106 ( .A1(n13298), .A2(n13297), .ZN(n9738) );
  NAND2_X2 U11284 ( .A1(n19004), .A2(n18992), .ZN(n18447) );
  NOR2_X2 U14987 ( .A1(n9725), .A2(n16856), .ZN(n18150) );
  AND2_X1 U12786 ( .A1(n14953), .A2(n9785), .ZN(n14904) );
  INV_X1 U11232 ( .A(n18176), .ZN(n18118) );
  CLKBUF_X1 U11147 ( .A(n12450), .Z(n12548) );
  NAND3_X2 U11153 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13115) );
  XNOR2_X1 U11170 ( .A(n11972), .B(n11973), .ZN(n12011) );
  CLKBUF_X1 U11172 ( .A(n10284), .Z(n10661) );
  CLKBUF_X1 U11186 ( .A(n10977), .Z(n9720) );
  NAND2_X1 U11225 ( .A1(n12011), .A2(n13237), .ZN(n12015) );
  CLKBUF_X1 U11237 ( .A(n10661), .Z(n10662) );
  CLKBUF_X1 U11238 ( .A(n11397), .Z(n11638) );
  CLKBUF_X1 U11272 ( .A(n13230), .Z(n15783) );
  CLKBUF_X1 U11300 ( .A(n10318), .Z(n10321) );
  INV_X1 U11313 ( .A(n17470), .ZN(n17511) );
  CLKBUF_X1 U11481 ( .A(n14893), .Z(n14894) );
  CLKBUF_X2 U11565 ( .A(n11390), .Z(n13338) );
  CLKBUF_X2 U11703 ( .A(n9684), .Z(n9730) );
  CLKBUF_X1 U12460 ( .A(n18168), .Z(n9729) );
  INV_X1 U12802 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14807) );
  CLKBUF_X1 U12832 ( .A(n18078), .Z(n9664) );
  OR2_X1 U13381 ( .A1(n11315), .A2(n19564), .ZN(n21233) );
  CLKBUF_X1 U15273 ( .A(n11866), .Z(n12383) );
  CLKBUF_X1 U15284 ( .A(n17821), .Z(n17829) );
endmodule

