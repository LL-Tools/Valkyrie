

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput0, keyinput1, keyinput2, 
        keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, 
        keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, 
        keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, 
        keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, 
        keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, 
        keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, 
        keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, 
        keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, 
        keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, 
        keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, 
        keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862;

  NAND2_X1 U3408 ( .A1(n5684), .A2(n4335), .ZN(n5649) );
  OAI21_X1 U3409 ( .B1(n6357), .B2(n3113), .A(n3010), .ZN(n3009) );
  XNOR2_X1 U3410 ( .A(n3055), .B(n3389), .ZN(n3514) );
  OAI21_X1 U3411 ( .B1(n3490), .B2(n3489), .A(n3488), .ZN(n3057) );
  INV_X2 U3412 ( .A(n3674), .ZN(n3977) );
  AND2_X2 U3413 ( .A1(n3322), .A2(n3986), .ZN(n4297) );
  CLKBUF_X2 U3414 ( .A(n3287), .Z(n3965) );
  CLKBUF_X2 U3415 ( .A(n3263), .Z(n3964) );
  OR2_X1 U3416 ( .A1(n3328), .A2(n3322), .ZN(n5491) );
  AND4_X1 U3417 ( .A1(n3186), .A2(n3185), .A3(n3184), .A4(n3183), .ZN(n3202)
         );
  BUF_X2 U3418 ( .A(n3242), .Z(n3863) );
  AND2_X2 U3419 ( .A1(n4506), .A2(n5179), .ZN(n3926) );
  NAND2_X1 U3420 ( .A1(n3369), .A2(n3370), .ZN(n2960) );
  AND2_X1 U3421 ( .A1(n5684), .A2(n4335), .ZN(n2961) );
  NAND2_X1 U3422 ( .A1(n3369), .A2(n3370), .ZN(n3441) );
  INV_X1 U3423 ( .A(n3788), .ZN(n3900) );
  CLKBUF_X2 U3424 ( .A(n3381), .Z(n3864) );
  NAND2_X1 U3425 ( .A1(n3496), .A2(n3436), .ZN(n3489) );
  AND2_X1 U3426 ( .A1(n3018), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3176)
         );
  AND2_X1 U3427 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4719) );
  INV_X1 U3428 ( .A(n3328), .ZN(n3285) );
  AND2_X2 U3429 ( .A1(n5254), .A2(n4192), .ZN(n5232) );
  INV_X1 U3430 ( .A(n6266), .ZN(n6280) );
  INV_X1 U3431 ( .A(n3546), .ZN(n3674) );
  NAND2_X1 U3432 ( .A1(n4183), .A2(n4182), .ZN(n5848) );
  OR2_X1 U3433 ( .A1(n5888), .A2(n3004), .ZN(n5872) );
  NOR2_X2 U3434 ( .A1(n6029), .A2(n4126), .ZN(n6032) );
  OR2_X1 U3435 ( .A1(n5275), .A2(n5257), .ZN(n5259) );
  OR2_X1 U3436 ( .A1(n4488), .A2(n4415), .ZN(n4489) );
  NAND2_X1 U3437 ( .A1(n4596), .A2(n4598), .ZN(n4597) );
  INV_X1 U3438 ( .A(n5641), .ZN(n5645) );
  AND2_X2 U3439 ( .A1(n4506), .A2(n3176), .ZN(n2962) );
  AND2_X2 U3440 ( .A1(n5179), .A2(n3155), .ZN(n2963) );
  NAND2_X1 U3441 ( .A1(n3058), .A2(n4323), .ZN(n5779) );
  AOI21_X1 U3442 ( .B1(n5660), .B2(n5667), .A(n3082), .ZN(n5661) );
  OAI22_X1 U3443 ( .A1(n5861), .A2(n5667), .B1(n5678), .B2(n5650), .ZN(n5651)
         );
  NAND2_X1 U3444 ( .A1(n2961), .A2(n3134), .ZN(n5667) );
  AND2_X4 U34450 ( .A1(n3176), .A2(n3155), .ZN(n3243) );
  NOR2_X4 U34460 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3178) );
  OR2_X1 U34470 ( .A1(n5852), .A2(n6345), .ZN(n4339) );
  NAND2_X1 U34480 ( .A1(n3009), .A2(n4308), .ZN(n5152) );
  AOI21_X1 U3449 ( .B1(n3085), .B2(n3087), .A(n2987), .ZN(n3083) );
  AOI21_X1 U3450 ( .B1(n3090), .B2(n3089), .A(n2978), .ZN(n3088) );
  AND2_X1 U34510 ( .A1(n3112), .A2(n4296), .ZN(n3010) );
  AND2_X1 U34520 ( .A1(n3013), .A2(n3011), .ZN(n4970) );
  NAND2_X1 U34530 ( .A1(n5200), .A2(n5199), .ZN(n5234) );
  OR2_X1 U3454 ( .A1(n5941), .A2(n5834), .ZN(n5921) );
  NOR2_X1 U34550 ( .A1(n3120), .A2(n3116), .ZN(n3115) );
  NAND2_X1 U34560 ( .A1(n3015), .A2(n3080), .ZN(n6367) );
  NAND2_X2 U3457 ( .A1(n5645), .A2(n4628), .ZN(n4987) );
  INV_X2 U3458 ( .A(n4329), .ZN(n2964) );
  AOI21_X1 U34590 ( .B1(n4256), .B2(n4297), .A(n4255), .ZN(n6366) );
  NOR2_X1 U34600 ( .A1(n6016), .A2(n6436), .ZN(n6041) );
  CLKBUF_X1 U34610 ( .A(n4251), .Z(n6670) );
  NAND2_X1 U34620 ( .A1(n4460), .A2(n4697), .ZN(n6016) );
  NAND2_X2 U34630 ( .A1(n4460), .A2(n4449), .ZN(n6381) );
  INV_X2 U34640 ( .A(n4905), .ZN(n4592) );
  NOR2_X2 U34650 ( .A1(n6690), .A2(n4205), .ZN(n5547) );
  NAND2_X1 U3466 ( .A1(n4260), .A2(n4259), .ZN(n4428) );
  NAND2_X1 U3467 ( .A1(n3057), .A2(n3056), .ZN(n3513) );
  NAND2_X1 U34680 ( .A1(n3459), .A2(n3458), .ZN(n4733) );
  INV_X2 U34690 ( .A(n4729), .ZN(n4642) );
  CLKBUF_X1 U34700 ( .A(n4635), .Z(n6144) );
  NAND2_X1 U34710 ( .A1(n3490), .A2(n3489), .ZN(n3056) );
  CLKBUF_X1 U34720 ( .A(n4729), .Z(n6461) );
  NAND2_X1 U34730 ( .A1(n3039), .A2(n4046), .ZN(n4488) );
  NAND2_X1 U34740 ( .A1(n2990), .A2(n3016), .ZN(n3496) );
  OAI21_X1 U3475 ( .B1(n4042), .B2(n2983), .A(n3037), .ZN(n3039) );
  OR2_X1 U3476 ( .A1(n4027), .A2(n4026), .ZN(n4042) );
  AND3_X1 U3477 ( .A1(n3356), .A2(n3358), .A3(n3357), .ZN(n3354) );
  NAND2_X1 U3478 ( .A1(n4092), .A2(n4091), .ZN(n3154) );
  NAND2_X1 U3479 ( .A1(n3316), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3317) );
  NAND3_X1 U3480 ( .A1(n3314), .A2(n3313), .A3(n3312), .ZN(n3348) );
  MUX2_X1 U3481 ( .A(n3437), .B(n4311), .S(n3432), .Z(n3499) );
  AND2_X1 U3482 ( .A1(n3310), .A2(n3324), .ZN(n3314) );
  NOR2_X1 U3483 ( .A1(n3433), .A2(n6747), .ZN(n4311) );
  AND2_X2 U3484 ( .A1(n3346), .A2(n3334), .ZN(n4039) );
  CLKBUF_X1 U3485 ( .A(n3325), .Z(n3326) );
  INV_X2 U3486 ( .A(n4527), .ZN(n5204) );
  OR2_X1 U3487 ( .A1(n3431), .A2(n3430), .ZN(n4266) );
  NAND2_X2 U3488 ( .A1(n3285), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3315) );
  AND2_X2 U3489 ( .A1(n3328), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3346) );
  INV_X1 U3490 ( .A(n3308), .ZN(n3325) );
  NAND2_X1 U3491 ( .A1(n2969), .A2(n2980), .ZN(n3135) );
  NAND2_X1 U3492 ( .A1(n2970), .A2(n2981), .ZN(n3341) );
  NAND4_X2 U3493 ( .A1(n3234), .A2(n3233), .A3(n3232), .A4(n3231), .ZN(n3282)
         );
  AND4_X1 U3494 ( .A1(n3212), .A2(n3211), .A3(n3210), .A4(n3209), .ZN(n3213)
         );
  AND4_X1 U3495 ( .A1(n3207), .A2(n3206), .A3(n3205), .A4(n3204), .ZN(n3214)
         );
  AND4_X1 U3496 ( .A1(n3230), .A2(n3229), .A3(n3228), .A4(n3227), .ZN(n3231)
         );
  AND4_X1 U3497 ( .A1(n3222), .A2(n3221), .A3(n3220), .A4(n3219), .ZN(n3233)
         );
  AND4_X1 U3498 ( .A1(n3247), .A2(n3246), .A3(n3245), .A4(n3244), .ZN(n3248)
         );
  AND4_X1 U3499 ( .A1(n3218), .A2(n3217), .A3(n3216), .A4(n3215), .ZN(n3234)
         );
  AND4_X1 U3500 ( .A1(n3241), .A2(n3240), .A3(n3239), .A4(n3238), .ZN(n3249)
         );
  BUF_X2 U3501 ( .A(n3295), .Z(n3920) );
  BUF_X2 U3502 ( .A(n3863), .Z(n3958) );
  NOR2_X1 U3503 ( .A1(n6358), .A2(n4667), .ZN(n6631) );
  BUF_X2 U3504 ( .A(n3243), .Z(n3963) );
  BUF_X2 U3505 ( .A(n3375), .Z(n3825) );
  OR2_X2 U3506 ( .A1(n6666), .A2(n6672), .ZN(n6358) );
  BUF_X2 U3507 ( .A(n3926), .Z(n3944) );
  BUF_X2 U3508 ( .A(n3273), .Z(n3882) );
  BUF_X2 U3509 ( .A(n3288), .Z(n2965) );
  INV_X2 U3510 ( .A(n4373), .ZN(n2966) );
  OAI211_X1 U3511 ( .C1(n3355), .C2(n3339), .A(n3354), .B(n3359), .ZN(n3077)
         );
  AND2_X4 U3513 ( .A1(n3008), .A2(n3007), .ZN(n4506) );
  OR2_X1 U3514 ( .A1(n3545), .A2(n3544), .ZN(n4300) );
  NAND2_X1 U3515 ( .A1(n2971), .A2(n3020), .ZN(n3645) );
  NOR2_X1 U3516 ( .A1(n4544), .A2(n2999), .ZN(n3020) );
  OR2_X1 U3517 ( .A1(n3421), .A2(n3420), .ZN(n4315) );
  INV_X1 U3518 ( .A(n3342), .ZN(n4065) );
  NAND2_X1 U3519 ( .A1(n3022), .A2(n2998), .ZN(n5243) );
  INV_X1 U3520 ( .A(n5296), .ZN(n3022) );
  INV_X1 U3521 ( .A(n3108), .ZN(n3107) );
  NOR2_X1 U3522 ( .A1(n3799), .A2(n5716), .ZN(n3075) );
  NAND2_X1 U3523 ( .A1(n3646), .A2(n3658), .ZN(n3024) );
  NAND2_X1 U3524 ( .A1(n6367), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3012)
         );
  INV_X1 U3525 ( .A(n3516), .ZN(n3685) );
  INV_X1 U3526 ( .A(n3086), .ZN(n3085) );
  OAI21_X1 U3527 ( .B1(n2968), .B2(n3087), .A(n4328), .ZN(n3086) );
  AND2_X1 U3528 ( .A1(n4733), .A2(n3096), .ZN(n3095) );
  NOR2_X1 U3529 ( .A1(n3097), .A2(n3554), .ZN(n3096) );
  INV_X1 U3530 ( .A(n3168), .ZN(n3097) );
  NAND2_X1 U3531 ( .A1(n6026), .A2(n6795), .ZN(n3054) );
  AND2_X1 U3532 ( .A1(n2979), .A2(n3151), .ZN(n3150) );
  INV_X1 U3533 ( .A(n5397), .ZN(n3151) );
  INV_X1 U3534 ( .A(n3115), .ZN(n3089) );
  NAND2_X2 U3535 ( .A1(n5350), .A2(n4527), .ZN(n5196) );
  NAND2_X1 U3536 ( .A1(n4428), .A2(n4262), .ZN(n3080) );
  NAND2_X1 U3537 ( .A1(n3701), .A2(n3169), .ZN(n3312) );
  AND4_X1 U3538 ( .A1(n3267), .A2(n3266), .A3(n3265), .A4(n3264), .ZN(n3280)
         );
  NAND2_X1 U3539 ( .A1(n3287), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3265) );
  AND2_X1 U3540 ( .A1(n5538), .A2(EBX_REG_12__SCAN_IN), .ZN(n3067) );
  NAND2_X1 U3541 ( .A1(n3876), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3895)
         );
  INV_X1 U3542 ( .A(n3877), .ZN(n3876) );
  NAND2_X1 U3543 ( .A1(n3128), .A2(n2977), .ZN(n3127) );
  INV_X1 U3544 ( .A(n5779), .ZN(n3128) );
  NAND2_X1 U3545 ( .A1(n5994), .A2(n5999), .ZN(n6045) );
  INV_X1 U3546 ( .A(n4263), .ZN(n6146) );
  OR2_X1 U3547 ( .A1(n6647), .A2(n4638), .ZN(n4639) );
  INV_X1 U3548 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6657) );
  INV_X1 U3549 ( .A(n5865), .ZN(n4197) );
  AND2_X2 U3550 ( .A1(n3339), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3177)
         );
  NAND2_X1 U3551 ( .A1(n3026), .A2(n3025), .ZN(n4004) );
  NAND2_X1 U3552 ( .A1(n3986), .A2(n3350), .ZN(n3025) );
  NAND2_X1 U3553 ( .A1(n3447), .A2(n3027), .ZN(n3026) );
  AND2_X1 U3554 ( .A1(n3986), .A2(n3315), .ZN(n3027) );
  NAND2_X1 U3555 ( .A1(n3997), .A2(n3308), .ZN(n3092) );
  INV_X1 U3556 ( .A(n3315), .ZN(n3388) );
  AND2_X1 U3557 ( .A1(n3353), .A2(n3352), .ZN(n3359) );
  AOI21_X1 U3558 ( .B1(n3863), .B2(INSTQUEUE_REG_2__4__SCAN_IN), .A(n3203), 
        .ZN(n3206) );
  AOI22_X1 U3559 ( .A1(n3286), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        INSTQUEUE_REG_4__4__SCAN_IN), .B2(n2962), .ZN(n3210) );
  AOI21_X1 U3560 ( .B1(n3243), .B2(INSTQUEUE_REG_6__4__SCAN_IN), .A(n3208), 
        .ZN(n3212) );
  AND2_X1 U3561 ( .A1(n3295), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3208) );
  OR2_X1 U3562 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n6681), .ZN(n4028)
         );
  NAND2_X1 U3563 ( .A1(n4032), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4035) );
  OR2_X1 U3564 ( .A1(n4034), .A2(n4035), .ZN(n4057) );
  INV_X1 U3565 ( .A(n4151), .ZN(n3146) );
  NAND2_X1 U3566 ( .A1(n3741), .A2(n3021), .ZN(n5296) );
  AND2_X1 U3567 ( .A1(n3000), .A2(n3740), .ZN(n3021) );
  INV_X1 U3568 ( .A(n3157), .ZN(n3156) );
  NAND2_X1 U3569 ( .A1(n5335), .A2(n3159), .ZN(n3158) );
  INV_X1 U3570 ( .A(n5348), .ZN(n3159) );
  NOR2_X1 U3571 ( .A1(n3163), .A2(n3162), .ZN(n3161) );
  INV_X1 U3572 ( .A(n5391), .ZN(n3162) );
  NAND2_X1 U3573 ( .A1(n3690), .A2(n5419), .ZN(n3163) );
  AND2_X1 U3574 ( .A1(n3643), .A2(n3642), .ZN(n3644) );
  INV_X1 U3575 ( .A(n5161), .ZN(n3164) );
  AND2_X1 U3576 ( .A1(n3618), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3619)
         );
  NOR2_X1 U3577 ( .A1(n5498), .A2(n3063), .ZN(n3062) );
  INV_X1 U3578 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3063) );
  NAND2_X1 U3579 ( .A1(n4281), .A2(n4297), .ZN(n3102) );
  INV_X1 U3580 ( .A(n5188), .ZN(n3855) );
  AND2_X1 U3581 ( .A1(n4073), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3518) );
  NAND2_X1 U3582 ( .A1(n3135), .A2(n3322), .ZN(n4074) );
  INV_X1 U3583 ( .A(n4327), .ZN(n3087) );
  NAND2_X1 U3584 ( .A1(n4158), .A2(n3148), .ZN(n3147) );
  INV_X1 U3585 ( .A(n5324), .ZN(n3148) );
  NAND2_X1 U3586 ( .A1(n3044), .A2(n2986), .ZN(n5693) );
  INV_X1 U3587 ( .A(n5723), .ZN(n3043) );
  AND2_X1 U3588 ( .A1(n3122), .A2(n2984), .ZN(n2968) );
  INV_X1 U3589 ( .A(n5412), .ZN(n3152) );
  AND2_X1 U3590 ( .A1(n3117), .A2(n2975), .ZN(n3090) );
  INV_X1 U3591 ( .A(n5812), .ZN(n3120) );
  INV_X1 U3592 ( .A(n5138), .ZN(n3116) );
  AND2_X1 U3593 ( .A1(n3118), .A2(n5813), .ZN(n3117) );
  NAND2_X1 U3594 ( .A1(n5812), .A2(n3119), .ZN(n3118) );
  INV_X1 U3595 ( .A(n4320), .ZN(n3119) );
  NAND2_X1 U3596 ( .A1(n4305), .A2(n4304), .ZN(n4309) );
  NAND2_X1 U3597 ( .A1(n4527), .A2(n4177), .ZN(n4170) );
  AND2_X1 U3598 ( .A1(n4662), .A2(n3308), .ZN(n4073) );
  INV_X1 U3599 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4748) );
  AND4_X1 U3600 ( .A1(n3299), .A2(n3298), .A3(n3297), .A4(n3296), .ZN(n3300)
         );
  AOI22_X1 U3601 ( .A1(n3287), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3286), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U3602 ( .A1(n4036), .A2(n4035), .ZN(n4056) );
  OR2_X1 U3603 ( .A1(n4034), .A2(n4033), .ZN(n4036) );
  AND2_X1 U3604 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6446), .ZN(n4033)
         );
  OR2_X1 U3605 ( .A1(n5530), .A2(n5463), .ZN(n5472) );
  AND3_X1 U3606 ( .A1(n4065), .A2(n4064), .A3(n4063), .ZN(n4086) );
  AND2_X1 U3607 ( .A1(n5591), .A2(n3017), .ZN(n4063) );
  AND2_X1 U3608 ( .A1(n4253), .A2(n3003), .ZN(n3017) );
  AND2_X1 U3609 ( .A1(n4569), .A2(n4061), .ZN(n4629) );
  INV_X1 U3610 ( .A(n4464), .ZN(n4465) );
  CLKBUF_X1 U3611 ( .A(n4070), .Z(n4071) );
  OR2_X1 U3612 ( .A1(n4903), .A2(n4420), .ZN(n4464) );
  AND2_X1 U3613 ( .A1(n3985), .A2(n3166), .ZN(n3106) );
  CLKBUF_X1 U3614 ( .A(n5243), .Z(n5244) );
  NAND2_X1 U3615 ( .A1(n3075), .A2(n3852), .ZN(n3877) );
  OR2_X1 U3616 ( .A1(n5323), .A2(n3158), .ZN(n3157) );
  CLKBUF_X1 U3617 ( .A(n5296), .Z(n5297) );
  AND2_X1 U3618 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3691) );
  OR2_X1 U3619 ( .A1(n3656), .A2(n3655), .ZN(n3657) );
  INV_X1 U3620 ( .A(n3024), .ZN(n3023) );
  NOR2_X1 U3621 ( .A1(n4968), .A2(n4631), .ZN(n3078) );
  INV_X1 U3622 ( .A(n4544), .ZN(n3019) );
  NAND2_X1 U3623 ( .A1(n3061), .A2(n3062), .ZN(n3572) );
  NOR2_X1 U3624 ( .A1(n3519), .A2(n3060), .ZN(n3529) );
  NAND2_X1 U3625 ( .A1(n4520), .A2(n4521), .ZN(n3015) );
  NAND2_X1 U3626 ( .A1(n4488), .A2(n6654), .ZN(n4903) );
  NAND2_X1 U3627 ( .A1(n4093), .A2(n4177), .ZN(n5205) );
  NAND2_X1 U3628 ( .A1(n3134), .A2(n3005), .ZN(n3130) );
  OR2_X1 U3629 ( .A1(n5823), .A2(n3033), .ZN(n3031) );
  NAND2_X1 U3630 ( .A1(n6016), .A2(n3002), .ZN(n3033) );
  AND2_X1 U3631 ( .A1(n3035), .A2(n3002), .ZN(n3032) );
  NOR2_X1 U3632 ( .A1(n5926), .A2(n5825), .ZN(n3035) );
  NAND2_X1 U3633 ( .A1(n6056), .A2(n6016), .ZN(n3034) );
  NAND2_X1 U3634 ( .A1(n3046), .A2(n3054), .ZN(n3045) );
  INV_X1 U3635 ( .A(n3049), .ZN(n3046) );
  AOI21_X1 U3636 ( .B1(n3051), .B2(n3053), .A(n3050), .ZN(n3049) );
  INV_X1 U3637 ( .A(n5731), .ZN(n3050) );
  OR2_X1 U3638 ( .A1(n5703), .A2(n3047), .ZN(n3044) );
  NAND2_X1 U3639 ( .A1(n3051), .A2(n3054), .ZN(n3047) );
  INV_X1 U3640 ( .A(n5693), .ZN(n5722) );
  NAND2_X1 U3641 ( .A1(n3121), .A2(n2968), .ZN(n5703) );
  NOR2_X1 U3642 ( .A1(n6026), .A2(n5988), .ZN(n3126) );
  NAND2_X1 U3643 ( .A1(n5786), .A2(n5787), .ZN(n3058) );
  NAND2_X1 U3644 ( .A1(n5152), .A2(n4310), .ZN(n5139) );
  NAND2_X1 U3645 ( .A1(n5139), .A2(n5138), .ZN(n5137) );
  NAND2_X1 U3646 ( .A1(n3496), .A2(n3500), .ZN(n4729) );
  XNOR2_X1 U3647 ( .A(n4748), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6464)
         );
  AND4_X1 U3648 ( .A1(n3272), .A2(n3271), .A3(n3270), .A4(n3269), .ZN(n3279)
         );
  AND4_X1 U3649 ( .A1(n3262), .A2(n3261), .A3(n3260), .A4(n3259), .ZN(n3281)
         );
  CLKBUF_X2 U3650 ( .A(n3341), .Z(n4662) );
  OR2_X1 U3651 ( .A1(n6670), .A2(n4752), .ZN(n4756) );
  INV_X1 U3652 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n5093) );
  INV_X1 U3653 ( .A(n4738), .ZN(n4737) );
  OAI21_X1 U3654 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .A(
        n4347), .ZN(n4208) );
  NAND2_X1 U3655 ( .A1(n6266), .A2(n5801), .ZN(n5450) );
  NOR2_X1 U3656 ( .A1(n6282), .A2(n5454), .ZN(n3069) );
  OAI21_X1 U3657 ( .B1(n5570), .B2(n5453), .A(n3066), .ZN(n3065) );
  AND2_X1 U3658 ( .A1(n3068), .A2(n2991), .ZN(n3066) );
  AND2_X1 U3659 ( .A1(n5191), .A2(n3076), .ZN(n6266) );
  NOR2_X1 U3660 ( .A1(n5547), .A2(n4722), .ZN(n3076) );
  NOR2_X1 U3661 ( .A1(n4206), .A2(n5547), .ZN(n6267) );
  OR2_X1 U3662 ( .A1(n5191), .A2(n4722), .ZN(n4206) );
  INV_X1 U3663 ( .A(n6279), .ZN(n5570) );
  AND2_X1 U3664 ( .A1(n4188), .A2(n4191), .ZN(n5665) );
  NAND2_X1 U3665 ( .A1(n4189), .A2(n4190), .ZN(n4191) );
  NAND2_X1 U3666 ( .A1(n5857), .A2(n5856), .ZN(n3137) );
  NOR2_X1 U3667 ( .A1(n5874), .A2(n3040), .ZN(n5853) );
  AND2_X1 U3668 ( .A1(n5972), .A2(n5861), .ZN(n3040) );
  OR2_X1 U3669 ( .A1(n5232), .A2(n4193), .ZN(n5865) );
  NAND2_X1 U3670 ( .A1(n2976), .A2(n3041), .ZN(n5874) );
  NAND2_X1 U3671 ( .A1(n5972), .A2(n3004), .ZN(n3041) );
  NAND2_X1 U3672 ( .A1(n3042), .A2(n2985), .ZN(n5906) );
  INV_X1 U3673 ( .A(n5923), .ZN(n3042) );
  INV_X1 U3674 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6681) );
  INV_X1 U3675 ( .A(n6671), .ZN(n6677) );
  INV_X1 U3676 ( .A(n6144), .ZN(n6675) );
  AND3_X1 U3677 ( .A1(n6152), .A2(n6151), .A3(n6150), .ZN(n6185) );
  INV_X1 U3678 ( .A(n6147), .ZN(n6192) );
  INV_X1 U3679 ( .A(n6623), .ZN(n6492) );
  AND2_X1 U3680 ( .A1(n4004), .A2(n3998), .ZN(n3028) );
  AND2_X1 U3681 ( .A1(n6463), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3994)
         );
  AND2_X1 U3682 ( .A1(n4016), .A2(n4011), .ZN(n4014) );
  AND2_X1 U3683 ( .A1(n3111), .A2(n5261), .ZN(n3110) );
  INV_X1 U3684 ( .A(n5271), .ZN(n3111) );
  OR2_X1 U3685 ( .A1(n3483), .A2(n3482), .ZN(n4289) );
  NAND2_X1 U3686 ( .A1(n3098), .A2(n3460), .ZN(n3553) );
  AND2_X1 U3687 ( .A1(n4733), .A2(n3168), .ZN(n3098) );
  OR2_X1 U3688 ( .A1(n3470), .A2(n3469), .ZN(n4290) );
  OR2_X1 U3689 ( .A1(n3402), .A2(n3401), .ZN(n4265) );
  CLKBUF_X1 U3690 ( .A(n2963), .Z(n3728) );
  AOI21_X1 U3691 ( .B1(n3499), .B2(n3497), .A(n4311), .ZN(n3436) );
  NAND2_X1 U3693 ( .A1(n3329), .A2(n4051), .ZN(n4080) );
  AND2_X1 U3694 ( .A1(n3282), .A2(n3308), .ZN(n3169) );
  NAND4_X1 U3695 ( .A1(n3351), .A2(n3236), .A3(n3350), .A4(n3388), .ZN(n3357)
         );
  NAND2_X1 U3696 ( .A1(n4472), .A2(n3167), .ZN(n3356) );
  AND2_X1 U3697 ( .A1(n4073), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3167) );
  INV_X1 U3698 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4010) );
  AOI21_X1 U3699 ( .B1(n3295), .B2(INSTQUEUE_REG_14__2__SCAN_IN), .A(n3294), 
        .ZN(n3296) );
  AND2_X1 U3700 ( .A1(n2962), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3294) );
  AOI22_X1 U3701 ( .A1(n3375), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3258) );
  OR2_X1 U3702 ( .A1(n3457), .A2(n3456), .ZN(n4274) );
  NAND2_X1 U3703 ( .A1(n3447), .A2(n3315), .ZN(n4013) );
  INV_X1 U3704 ( .A(n4013), .ZN(n4037) );
  AOI21_X1 U3705 ( .B1(n4037), .B2(n4297), .A(n4057), .ZN(n4041) );
  NAND2_X1 U3706 ( .A1(n4039), .A2(n4297), .ZN(n4043) );
  OR2_X1 U3707 ( .A1(n3892), .A2(n3891), .ZN(n3898) );
  NOR2_X1 U3708 ( .A1(n4190), .A2(n5246), .ZN(n3166) );
  NAND2_X1 U3709 ( .A1(n3109), .A2(n5287), .ZN(n3108) );
  INV_X1 U3710 ( .A(n5298), .ZN(n3109) );
  NOR2_X1 U3711 ( .A1(n4510), .A2(n6747), .ZN(n3953) );
  NAND2_X1 U3712 ( .A1(n3535), .A2(n3534), .ZN(n3484) );
  AOI21_X1 U3713 ( .B1(n3125), .B2(n3123), .A(n2988), .ZN(n3122) );
  INV_X1 U3714 ( .A(n2977), .ZN(n3123) );
  NAND2_X1 U3715 ( .A1(n4107), .A2(n3143), .ZN(n3142) );
  INV_X1 U3716 ( .A(n4633), .ZN(n3143) );
  INV_X1 U3717 ( .A(n4549), .ZN(n4107) );
  NAND2_X1 U3718 ( .A1(n5204), .A2(n4089), .ZN(n4128) );
  AOI22_X1 U3719 ( .A1(n4039), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3388), 
        .B2(n4252), .ZN(n3389) );
  NAND2_X1 U3720 ( .A1(n3100), .A2(n3099), .ZN(n3055) );
  NAND2_X1 U3721 ( .A1(n4252), .A2(n4064), .ZN(n3099) );
  OR2_X1 U3722 ( .A1(n6670), .A2(n4733), .ZN(n6510) );
  NAND2_X1 U3723 ( .A1(n3295), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3192)
         );
  AND4_X1 U3724 ( .A1(n3292), .A2(n3291), .A3(n3290), .A4(n3289), .ZN(n3301)
         );
  AOI22_X1 U3725 ( .A1(n2963), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3263), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3179) );
  AOI22_X1 U3726 ( .A1(n3295), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3243), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3174) );
  AOI22_X1 U3727 ( .A1(n2962), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3286), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3173) );
  NAND2_X1 U3728 ( .A1(n3214), .A2(n3213), .ZN(n3333) );
  AOI22_X1 U3729 ( .A1(n2962), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n2963), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3247) );
  CLKBUF_X1 U3730 ( .A(n3349), .Z(n3992) );
  AND2_X1 U3731 ( .A1(n4025), .A2(n4024), .ZN(n4026) );
  INV_X1 U3732 ( .A(n3038), .ZN(n3037) );
  OAI22_X1 U3733 ( .A1(n4041), .A2(n4040), .B1(n4056), .B2(n4037), .ZN(n3038)
         );
  NAND2_X1 U3734 ( .A1(n5177), .A2(n6747), .ZN(n4237) );
  AND2_X1 U3735 ( .A1(n4058), .A2(n4057), .ZN(n4419) );
  OR2_X1 U3736 ( .A1(n4047), .A2(n3285), .ZN(n4420) );
  OR2_X1 U3737 ( .A1(n5328), .A2(n4215), .ZN(n4218) );
  INV_X1 U3738 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5327) );
  AND2_X1 U3739 ( .A1(n4145), .A2(n5349), .ZN(n5352) );
  NAND2_X1 U3740 ( .A1(n6247), .A2(REIP_REG_12__SCAN_IN), .ZN(n3068) );
  XNOR2_X1 U3741 ( .A(n2960), .B(n4857), .ZN(n4635) );
  NAND2_X1 U3742 ( .A1(n3077), .A2(n3390), .ZN(n3391) );
  AND2_X1 U3743 ( .A1(n4169), .A2(n4168), .ZN(n5257) );
  OR2_X1 U3744 ( .A1(n5336), .A2(n3144), .ZN(n5275) );
  INV_X1 U3745 ( .A(n3147), .ZN(n3145) );
  AND2_X1 U3746 ( .A1(n4113), .A2(n4112), .ZN(n4964) );
  XNOR2_X1 U3747 ( .A(n3154), .B(n4456), .ZN(n4528) );
  NAND2_X1 U3748 ( .A1(n4528), .A2(n4527), .ZN(n4526) );
  NOR2_X1 U3749 ( .A1(n4476), .A2(n4085), .ZN(n4458) );
  INV_X1 U3750 ( .A(n4073), .ZN(n4439) );
  AND3_X1 U3751 ( .A1(n3622), .A2(n3621), .A3(n3620), .ZN(n5161) );
  NAND2_X1 U3752 ( .A1(n3981), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4201)
         );
  NOR2_X1 U3753 ( .A1(n3895), .A2(n3072), .ZN(n3981) );
  NAND2_X1 U3754 ( .A1(n3073), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n3072)
         );
  NOR2_X1 U3755 ( .A1(n5671), .A2(n3074), .ZN(n3073) );
  OR2_X1 U3756 ( .A1(n3798), .A2(n5327), .ZN(n3799) );
  INV_X1 U3757 ( .A(n3075), .ZN(n3853) );
  AND2_X1 U3758 ( .A1(n3771), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3772)
         );
  NAND2_X1 U3759 ( .A1(n3772), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3798)
         );
  NOR2_X1 U3760 ( .A1(n3738), .A2(n5750), .ZN(n3771) );
  NOR2_X1 U3761 ( .A1(n5378), .A2(n3105), .ZN(n3104) );
  INV_X1 U3762 ( .A(n3161), .ZN(n3105) );
  INV_X1 U3763 ( .A(n5418), .ZN(n3160) );
  AND2_X1 U3764 ( .A1(n3637), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3638)
         );
  NAND2_X1 U3765 ( .A1(n6357), .A2(n4280), .ZN(n5001) );
  AOI21_X1 U3766 ( .B1(n4273), .B2(n3685), .A(n3531), .ZN(n4601) );
  NAND2_X1 U3767 ( .A1(n3014), .A2(n6440), .ZN(n3013) );
  NAND2_X1 U3768 ( .A1(n3012), .A2(n6366), .ZN(n3011) );
  INV_X1 U3769 ( .A(n6367), .ZN(n3014) );
  NAND2_X1 U3770 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3519) );
  AND2_X1 U3771 ( .A1(n3512), .A2(n3511), .ZN(n4609) );
  NOR2_X1 U3772 ( .A1(n3130), .A2(n5845), .ZN(n3129) );
  NAND2_X1 U3773 ( .A1(n3084), .A2(n3083), .ZN(n5686) );
  NOR3_X1 U3774 ( .A1(n5336), .A2(n4151), .A3(n3147), .ZN(n5301) );
  NOR3_X1 U3775 ( .A1(n5336), .A2(n4151), .A3(n5324), .ZN(n5326) );
  AND2_X1 U3776 ( .A1(n5441), .A2(n2982), .ZN(n5379) );
  INV_X1 U3777 ( .A(n5380), .ZN(n3149) );
  NAND2_X1 U3778 ( .A1(n5441), .A2(n3150), .ZN(n5399) );
  NAND2_X1 U3779 ( .A1(n3121), .A2(n3122), .ZN(n5765) );
  NAND2_X1 U3780 ( .A1(n5441), .A2(n2979), .ZN(n5414) );
  NAND2_X1 U3781 ( .A1(n3088), .A2(n3059), .ZN(n5786) );
  NAND2_X1 U3782 ( .A1(n5822), .A2(n5821), .ZN(n6000) );
  NAND2_X1 U3783 ( .A1(n5139), .A2(n3115), .ZN(n3101) );
  NOR2_X1 U3784 ( .A1(n4604), .A2(n3139), .ZN(n4984) );
  OR2_X1 U3785 ( .A1(n3142), .A2(n3140), .ZN(n3139) );
  INV_X1 U3786 ( .A(n4964), .ZN(n3140) );
  NAND2_X1 U3787 ( .A1(n6041), .A2(n5824), .ZN(n6042) );
  OR2_X1 U3788 ( .A1(n5823), .A2(n6434), .ZN(n6043) );
  NOR2_X1 U3789 ( .A1(n4604), .A2(n3142), .ZN(n4965) );
  NAND2_X1 U3790 ( .A1(n3141), .A2(n4107), .ZN(n4632) );
  INV_X1 U3791 ( .A(n4604), .ZN(n3141) );
  NAND2_X1 U3792 ( .A1(n6355), .A2(n6354), .ZN(n6357) );
  NAND2_X1 U3793 ( .A1(n4456), .A2(n4527), .ZN(n3153) );
  AND2_X1 U3794 ( .A1(n3081), .A2(n3080), .ZN(n4520) );
  NAND2_X1 U3795 ( .A1(n4261), .A2(n6800), .ZN(n3081) );
  NOR2_X1 U3796 ( .A1(n3348), .A2(n4051), .ZN(n4451) );
  OR2_X1 U3797 ( .A1(n4822), .A2(n6144), .ZN(n4933) );
  NOR2_X1 U3798 ( .A1(n4825), .A2(n6461), .ZN(n6075) );
  OR2_X1 U3799 ( .A1(n6117), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6115)
         );
  NOR2_X1 U3800 ( .A1(n6510), .A2(n6068), .ZN(n4788) );
  AND2_X1 U3801 ( .A1(n5092), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4789)
         );
  AND2_X1 U3802 ( .A1(n4786), .A2(n6681), .ZN(n5092) );
  AND3_X1 U3803 ( .A1(n6681), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6516) );
  NOR2_X1 U3804 ( .A1(n6510), .A2(n6146), .ZN(n6462) );
  AND2_X1 U3805 ( .A1(n4823), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6143)
         );
  OR2_X1 U3806 ( .A1(n5049), .A2(n4642), .ZN(n6074) );
  NOR2_X1 U3808 ( .A1(n5049), .A2(n6461), .ZN(n5089) );
  AND2_X1 U3809 ( .A1(n5056), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4754)
         );
  NOR2_X1 U3810 ( .A1(n5055), .A2(n5093), .ZN(n4689) );
  AND2_X1 U3811 ( .A1(n4786), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5056)
         );
  NOR2_X1 U3812 ( .A1(n6070), .A2(n4636), .ZN(n6472) );
  OR2_X1 U3813 ( .A1(n4863), .A2(n6657), .ZN(n6139) );
  NOR2_X1 U3814 ( .A1(n5055), .A2(n4650), .ZN(n6513) );
  INV_X1 U3815 ( .A(n4859), .ZN(n4740) );
  OR2_X1 U3816 ( .A1(n6670), .A2(n4734), .ZN(n4738) );
  OR2_X1 U3817 ( .A1(n4429), .A2(n3992), .ZN(n6209) );
  AND2_X1 U3818 ( .A1(n4722), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4062) );
  AND2_X1 U3819 ( .A1(n6747), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6723) );
  INV_X1 U3820 ( .A(STATE_REG_2__SCAN_IN), .ZN(n4367) );
  INV_X1 U3821 ( .A(n6654), .ZN(n6223) );
  INV_X1 U3822 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6469) );
  INV_X1 U3823 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5213) );
  OR2_X1 U3824 ( .A1(n5278), .A2(n4216), .ZN(n5263) );
  NOR2_X1 U3825 ( .A1(n5511), .A2(n4227), .ZN(n5538) );
  AND2_X1 U3826 ( .A1(n5386), .A2(n4211), .ZN(n5343) );
  INV_X1 U3827 ( .A(n6251), .ZN(n6273) );
  INV_X1 U3828 ( .A(n6249), .ZN(n6272) );
  NOR2_X1 U3829 ( .A1(n5472), .A2(n5464), .ZN(n6271) );
  INV_X1 U3830 ( .A(n5538), .ZN(n6276) );
  NOR2_X1 U3831 ( .A1(n5511), .A2(n4207), .ZN(n5553) );
  CLKBUF_X1 U3832 ( .A(n4504), .Z(n4505) );
  AND2_X2 U3833 ( .A1(n4629), .A2(n4066), .ZN(n5641) );
  NOR2_X1 U3834 ( .A1(n4629), .A2(n4628), .ZN(n5642) );
  INV_X1 U3835 ( .A(n5642), .ZN(n5647) );
  AND2_X1 U3836 ( .A1(n4908), .A2(n4907), .ZN(n6321) );
  NOR2_X2 U3837 ( .A1(n6321), .A2(n6331), .ZN(n6330) );
  INV_X1 U3838 ( .A(n6330), .ZN(n6337) );
  INV_X1 U3839 ( .A(n6321), .ZN(n6336) );
  INV_X2 U3840 ( .A(n4551), .ZN(n4593) );
  NAND2_X1 U3841 ( .A1(n4465), .A2(n4048), .ZN(n4569) );
  AOI21_X1 U3842 ( .B1(READY_N), .B2(n4071), .A(n4464), .ZN(n4551) );
  XNOR2_X1 U3843 ( .A(n4202), .B(n5213), .ZN(n5191) );
  OR2_X1 U3844 ( .A1(n4201), .A2(n4228), .ZN(n4202) );
  XNOR2_X1 U3845 ( .A(n5189), .B(n5592), .ZN(n5209) );
  INV_X1 U3846 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5671) );
  AOI21_X1 U3847 ( .B1(n5246), .B2(n5244), .A(n5245), .ZN(n5673) );
  AND2_X1 U3848 ( .A1(n3895), .A2(n3878), .ZN(n5688) );
  INV_X1 U3849 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5716) );
  NOR2_X1 U3850 ( .A1(n5347), .A2(n3157), .ZN(n5309) );
  INV_X1 U3851 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U3852 ( .A1(n3692), .A2(n2974), .ZN(n3737) );
  NAND2_X1 U3853 ( .A1(n3692), .A2(n3691), .ZN(n3721) );
  NAND2_X1 U3854 ( .A1(n3023), .A2(n3659), .ZN(n5431) );
  AND2_X1 U3855 ( .A1(n3061), .A2(n2972), .ZN(n3577) );
  OR2_X1 U3856 ( .A1(n4978), .A2(n4980), .ZN(n6283) );
  NOR2_X1 U3857 ( .A1(n3547), .A2(n5498), .ZN(n3548) );
  NAND2_X1 U3858 ( .A1(n5816), .A2(n4620), .ZN(n6375) );
  INV_X1 U3859 ( .A(n5816), .ZN(n6365) );
  INV_X1 U3860 ( .A(n6375), .ZN(n5818) );
  OR2_X2 U3861 ( .A1(n4903), .A2(n6209), .ZN(n6345) );
  INV_X1 U3862 ( .A(n6358), .ZN(n6370) );
  XNOR2_X1 U3863 ( .A(n5208), .B(n5207), .ZN(n5842) );
  INV_X1 U3864 ( .A(n5203), .ZN(n5208) );
  XNOR2_X1 U3865 ( .A(n3131), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5844)
         );
  NAND2_X1 U3866 ( .A1(n3133), .A2(n3132), .ZN(n3131) );
  NAND2_X1 U3867 ( .A1(n5658), .A2(n5187), .ZN(n3132) );
  NAND2_X1 U3868 ( .A1(n5678), .A2(n3129), .ZN(n3133) );
  OAI21_X1 U3869 ( .B1(n5649), .B2(n3130), .A(n3103), .ZN(n4338) );
  NAND2_X1 U3870 ( .A1(n5649), .A2(n4337), .ZN(n3103) );
  NAND2_X1 U3871 ( .A1(n3036), .A2(n3029), .ZN(n5827) );
  AND2_X1 U3872 ( .A1(n3031), .A2(n3030), .ZN(n3029) );
  NAND2_X1 U3873 ( .A1(n3044), .A2(n3045), .ZN(n5724) );
  NAND2_X1 U3874 ( .A1(n3048), .A2(n3051), .ZN(n5730) );
  NAND2_X1 U3875 ( .A1(n5703), .A2(n3052), .ZN(n3048) );
  NAND2_X1 U3876 ( .A1(n5703), .A2(n4327), .ZN(n5739) );
  INV_X1 U3877 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U3878 ( .A1(n3127), .A2(n3124), .ZN(n5772) );
  INV_X1 U3879 ( .A(n3126), .ZN(n3124) );
  NAND2_X1 U3880 ( .A1(n5137), .A2(n4320), .ZN(n5815) );
  INV_X1 U3881 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6400) );
  NOR2_X1 U3882 ( .A1(n6041), .A2(n6059), .ZN(n6425) );
  AND2_X1 U3883 ( .A1(n6045), .A2(n5828), .ZN(n6441) );
  INV_X1 U3884 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6463) );
  INV_X1 U3885 ( .A(n6146), .ZN(n6068) );
  INV_X1 U3886 ( .A(n4505), .ZN(n6070) );
  INV_X1 U3887 ( .A(n6672), .ZN(n6515) );
  NAND2_X1 U3888 ( .A1(n2960), .A2(n3374), .ZN(n4636) );
  OR2_X1 U3889 ( .A1(n6672), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6676) );
  INV_X1 U3890 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6446) );
  OAI21_X1 U3891 ( .B1(n4726), .B2(n6665), .A(n5055), .ZN(n6682) );
  AND2_X1 U3892 ( .A1(n4451), .A2(n3322), .ZN(n6196) );
  INV_X1 U3893 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3008) );
  INV_X1 U3894 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5174) );
  AOI21_X1 U3895 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6747), .A(n4497), .ZN(
        n5180) );
  INV_X1 U3896 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3006) );
  AND2_X1 U3897 ( .A1(n4451), .A2(n3350), .ZN(n4723) );
  NOR2_X1 U3898 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n5177) );
  INV_X1 U3899 ( .A(n5180), .ZN(n5176) );
  OR2_X1 U3900 ( .A1(n4928), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4958)
         );
  AND2_X1 U3901 ( .A1(n6081), .A2(n6080), .ZN(n6106) );
  NAND2_X1 U3902 ( .A1(n5089), .A2(n6677), .ZN(n6460) );
  NAND2_X1 U3903 ( .A1(n4788), .A2(n6461), .ZN(n5132) );
  NAND2_X1 U3904 ( .A1(n6516), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6700) );
  NAND2_X1 U3905 ( .A1(n4644), .A2(n4642), .ZN(n5015) );
  NOR2_X2 U3906 ( .A1(n4643), .A2(n4642), .ZN(n6147) );
  INV_X1 U3907 ( .A(n6585), .ZN(n5042) );
  INV_X1 U3908 ( .A(n5015), .ZN(n5044) );
  AND2_X1 U3909 ( .A1(n6556), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6584)
         );
  NOR2_X1 U3910 ( .A1(n6677), .A2(n6074), .ZN(n6585) );
  NOR2_X1 U3911 ( .A1(n6358), .A2(n4688), .ZN(n6563) );
  INV_X1 U3912 ( .A(n6586), .ZN(n5088) );
  INV_X1 U3913 ( .A(n6468), .ZN(n6566) );
  INV_X1 U3914 ( .A(n6601), .ZN(n6571) );
  INV_X1 U3915 ( .A(n6608), .ZN(n6574) );
  INV_X1 U3916 ( .A(n6615), .ZN(n6577) );
  INV_X1 U3917 ( .A(n6622), .ZN(n6580) );
  NAND2_X1 U3918 ( .A1(n4689), .A2(n3308), .ZN(n6539) );
  NAND2_X1 U3919 ( .A1(n4753), .A2(n4642), .ZN(n4862) );
  NOR2_X2 U3920 ( .A1(n4756), .A2(n4642), .ZN(n5085) );
  INV_X1 U3921 ( .A(n6637), .ZN(n6590) );
  AOI21_X1 U3922 ( .B1(n5056), .B2(STATE2_REG_2__SCAN_IN), .A(n4750), .ZN(
        n4785) );
  INV_X1 U3923 ( .A(n6563), .ZN(n6481) );
  NOR2_X1 U3924 ( .A1(n4988), .A2(n5055), .ZN(n6468) );
  NOR2_X1 U3925 ( .A1(n6358), .A2(n4687), .ZN(n6558) );
  NAND2_X1 U3926 ( .A1(n6370), .A2(DATAI_18_), .ZN(n6520) );
  INV_X1 U3927 ( .A(n6616), .ZN(n6530) );
  NAND2_X1 U3928 ( .A1(n6370), .A2(DATAI_22_), .ZN(n6540) );
  NAND2_X1 U3929 ( .A1(n4737), .A2(n6461), .ZN(n6594) );
  NOR2_X1 U3930 ( .A1(n4671), .A2(n5055), .ZN(n6593) );
  NOR2_X1 U3931 ( .A1(n6358), .A2(n4672), .ZN(n6596) );
  NOR2_X1 U3932 ( .A1(n4677), .A2(n5055), .ZN(n6601) );
  NOR2_X1 U3933 ( .A1(n4682), .A2(n5055), .ZN(n6608) );
  NOR2_X1 U3934 ( .A1(n4654), .A2(n5055), .ZN(n6615) );
  INV_X1 U3935 ( .A(n6534), .ZN(n6621) );
  NOR2_X1 U3936 ( .A1(n4640), .A2(n5055), .ZN(n6622) );
  NOR2_X1 U3937 ( .A1(n6358), .A2(n4645), .ZN(n6623) );
  NOR2_X1 U3938 ( .A1(n6358), .A2(n4641), .ZN(n6624) );
  NOR2_X1 U3939 ( .A1(n4666), .A2(n5055), .ZN(n6629) );
  AND2_X1 U3940 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4740), .ZN(n6636)
         );
  NOR2_X1 U3941 ( .A1(n4660), .A2(n5055), .ZN(n6637) );
  NOR2_X2 U3942 ( .A1(n4738), .A2(n6461), .ZN(n6640) );
  INV_X1 U3943 ( .A(n6594), .ZN(n6642) );
  NOR2_X1 U3944 ( .A1(n6358), .A2(n6784), .ZN(n6641) );
  AND2_X1 U3945 ( .A1(n4488), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6647) );
  AND2_X1 U3946 ( .A1(n4062), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6654) );
  NOR2_X1 U3947 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6694) );
  NOR2_X1 U3948 ( .A1(n4373), .A2(n4353), .ZN(n4363) );
  AOI21_X1 U3949 ( .B1(n4367), .B2(STATE_REG_1__SCAN_IN), .A(n4352), .ZN(n4353) );
  OR2_X1 U3950 ( .A1(n4208), .A2(STATE_REG_0__SCAN_IN), .ZN(n4906) );
  OR2_X1 U3951 ( .A1(n2966), .A2(STATE_REG_2__SCAN_IN), .ZN(n4372) );
  AND2_X1 U3952 ( .A1(n4234), .A2(n4233), .ZN(n4235) );
  NAND2_X1 U3953 ( .A1(n3070), .A2(n3064), .ZN(U2815) );
  INV_X1 U3954 ( .A(n5452), .ZN(n3070) );
  NOR2_X1 U3955 ( .A1(n3069), .A2(n3065), .ZN(n3064) );
  AND2_X1 U3956 ( .A1(n4186), .A2(n4185), .ZN(n4187) );
  OR2_X1 U3957 ( .A1(n5848), .A2(n6295), .ZN(n4186) );
  AOI21_X1 U3958 ( .B1(n4197), .B2(n4196), .A(n4195), .ZN(n4198) );
  NOR2_X1 U3959 ( .A1(n6302), .A2(n4194), .ZN(n4195) );
  AOI211_X1 U3960 ( .C1(n3138), .C2(n6433), .A(n5855), .B(n3136), .ZN(n5858)
         );
  NAND2_X1 U3961 ( .A1(n3137), .A2(n5854), .ZN(n3136) );
  INV_X2 U3962 ( .A(n3322), .ZN(n3350) );
  INV_X1 U3963 ( .A(n3165), .ZN(n4997) );
  INV_X1 U3964 ( .A(n3282), .ZN(n3997) );
  INV_X1 U3965 ( .A(n5491), .ZN(n3340) );
  OR2_X1 U3966 ( .A1(n5347), .A2(n3158), .ZN(n5322) );
  NAND2_X1 U3967 ( .A1(n3741), .A2(n3740), .ZN(n5347) );
  AND2_X1 U3968 ( .A1(n4978), .A2(n2994), .ZN(n2967) );
  NOR2_X1 U3969 ( .A1(n3163), .A2(n3160), .ZN(n5390) );
  AND4_X1 U3970 ( .A1(n3175), .A2(n3174), .A3(n3173), .A4(n3172), .ZN(n2969)
         );
  NAND2_X1 U3971 ( .A1(n4978), .A2(n2993), .ZN(n5158) );
  INV_X1 U3972 ( .A(n5675), .ZN(n3134) );
  AND4_X1 U3973 ( .A1(n3252), .A2(n3251), .A3(n3256), .A4(n3250), .ZN(n2970)
         );
  AND2_X1 U3974 ( .A1(n3078), .A2(n4979), .ZN(n2971) );
  INV_X1 U3975 ( .A(n3311), .ZN(n3701) );
  AND2_X1 U3976 ( .A1(n3062), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n2972)
         );
  AND3_X1 U3977 ( .A1(n3092), .A2(n3135), .A3(n3341), .ZN(n2973) );
  OR2_X1 U3978 ( .A1(n3334), .A2(n6747), .ZN(n3447) );
  NAND2_X1 U3979 ( .A1(n4978), .A2(n4998), .ZN(n3165) );
  NAND2_X1 U3980 ( .A1(n2964), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3094) );
  INV_X1 U3981 ( .A(n5972), .ZN(n6380) );
  OR2_X1 U3982 ( .A1(n6045), .A2(n6434), .ZN(n5972) );
  OR2_X1 U3983 ( .A1(n5738), .A2(n3093), .ZN(n3051) );
  AND2_X1 U3984 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n3691), .ZN(n2974)
         );
  OR2_X1 U3985 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3797) );
  INV_X2 U3986 ( .A(n3797), .ZN(n3982) );
  INV_X4 U3987 ( .A(n2964), .ZN(n6026) );
  INV_X1 U3988 ( .A(n3396), .ZN(n3966) );
  NAND2_X1 U3989 ( .A1(n3917), .A2(n3916), .ZN(n4189) );
  NAND2_X1 U3990 ( .A1(n3301), .A2(n3300), .ZN(n3311) );
  NAND2_X1 U3991 ( .A1(n5418), .A2(n3161), .ZN(n5377) );
  XNOR2_X1 U3992 ( .A(n3517), .B(n4733), .ZN(n4245) );
  NOR2_X1 U3993 ( .A1(n5270), .A2(n5271), .ZN(n5260) );
  NOR2_X1 U3994 ( .A1(n5296), .A2(n5298), .ZN(n5286) );
  OR2_X1 U3995 ( .A1(n4329), .A2(n4321), .ZN(n2975) );
  NOR2_X1 U3996 ( .A1(n5234), .A2(n5233), .ZN(n3138) );
  NOR2_X1 U3997 ( .A1(n5906), .A2(n5830), .ZN(n2976) );
  NAND2_X1 U3998 ( .A1(n4329), .A2(n5988), .ZN(n2977) );
  NAND2_X2 U3999 ( .A1(n4253), .A2(n3328), .ZN(n4093) );
  INV_X1 U4000 ( .A(n3295), .ZN(n3415) );
  NAND2_X1 U4001 ( .A1(n5792), .A2(n4322), .ZN(n2978) );
  NAND2_X1 U4002 ( .A1(n3016), .A2(n3410), .ZN(n3501) );
  AND2_X1 U4003 ( .A1(n5425), .A2(n3152), .ZN(n2979) );
  NAND2_X1 U4004 ( .A1(n3101), .A2(n3117), .ZN(n5793) );
  AND4_X1 U4005 ( .A1(n3182), .A2(n3181), .A3(n3180), .A4(n3179), .ZN(n2980)
         );
  NOR2_X1 U4006 ( .A1(n4188), .A2(n5221), .ZN(n5590) );
  AND3_X1 U4007 ( .A1(n3253), .A2(n3258), .A3(n3257), .ZN(n2981) );
  AND2_X1 U4008 ( .A1(n3092), .A2(n3341), .ZN(n4076) );
  AND2_X1 U4009 ( .A1(n3150), .A2(n3149), .ZN(n2982) );
  NAND2_X1 U4010 ( .A1(n3659), .A2(n3024), .ZN(n5418) );
  INV_X1 U4011 ( .A(n4631), .ZN(n3552) );
  AND2_X1 U4012 ( .A1(n4041), .A2(n4040), .ZN(n2983) );
  NOR2_X1 U4013 ( .A1(n4324), .A2(n3126), .ZN(n3125) );
  NAND2_X1 U4014 ( .A1(n4329), .A2(n4325), .ZN(n2984) );
  NAND2_X1 U4015 ( .A1(n5972), .A2(n5835), .ZN(n2985) );
  INV_X1 U4016 ( .A(n3053), .ZN(n3052) );
  NAND2_X1 U4017 ( .A1(n4327), .A2(n3094), .ZN(n3053) );
  AND2_X1 U4018 ( .A1(n3045), .A2(n3043), .ZN(n2986) );
  AND2_X1 U4019 ( .A1(n2964), .A2(n4331), .ZN(n2987) );
  AND2_X1 U4020 ( .A1(n4329), .A2(n5984), .ZN(n2988) );
  OR2_X1 U4021 ( .A1(n5336), .A2(n4151), .ZN(n2989) );
  AND2_X1 U4022 ( .A1(n3410), .A2(n6747), .ZN(n2990) );
  OR2_X1 U4023 ( .A1(n3387), .A2(n3386), .ZN(n4252) );
  NOR2_X1 U4024 ( .A1(n5451), .A2(n3067), .ZN(n2991) );
  NOR2_X1 U4025 ( .A1(n5347), .A2(n5348), .ZN(n2992) );
  INV_X1 U4026 ( .A(n3094), .ZN(n3093) );
  INV_X2 U4027 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6747) );
  NOR2_X1 U4028 ( .A1(n4662), .A2(n6657), .ZN(n3546) );
  INV_X1 U4029 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3339) );
  INV_X1 U4030 ( .A(n3135), .ZN(n4253) );
  INV_X1 U4031 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3007) );
  AND2_X1 U4032 ( .A1(n2971), .A2(n3019), .ZN(n4978) );
  NAND2_X1 U4033 ( .A1(n5441), .A2(n5425), .ZN(n5411) );
  AND2_X1 U4034 ( .A1(n3607), .A2(n4998), .ZN(n2993) );
  AND2_X1 U4035 ( .A1(n2993), .A2(n3164), .ZN(n2994) );
  INV_X1 U4036 ( .A(n6433), .ZN(n6034) );
  AND2_X1 U4037 ( .A1(n4460), .A2(n4455), .ZN(n6433) );
  NAND2_X1 U4038 ( .A1(n3019), .A2(n3552), .ZN(n4967) );
  AND2_X1 U4039 ( .A1(n3019), .A2(n3078), .ZN(n2995) );
  OR2_X1 U4040 ( .A1(n3895), .A2(n5262), .ZN(n2996) );
  OR3_X1 U4041 ( .A1(n3895), .A2(n5262), .A3(n5671), .ZN(n2997) );
  AND3_X1 U4042 ( .A1(n4065), .A2(n3340), .A3(n4253), .ZN(n4472) );
  AND2_X1 U4043 ( .A1(n3110), .A2(n3107), .ZN(n2998) );
  INV_X1 U4044 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5758) );
  NAND2_X1 U4045 ( .A1(n2994), .A2(n5164), .ZN(n2999) );
  AND2_X1 U4046 ( .A1(n5310), .A2(n3156), .ZN(n3000) );
  AND2_X1 U4047 ( .A1(n2974), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3001)
         );
  INV_X1 U4048 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3060) );
  AND2_X1 U4049 ( .A1(n4472), .A2(n4073), .ZN(n4445) );
  INV_X1 U4050 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3018) );
  AND2_X1 U4051 ( .A1(n5831), .A2(n5931), .ZN(n3002) );
  INV_X1 U4052 ( .A(n3547), .ZN(n3061) );
  AND2_X1 U4053 ( .A1(n3308), .A2(n4062), .ZN(n3003) );
  INV_X1 U4054 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n3074) );
  NAND2_X1 U4055 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3004) );
  INV_X1 U4056 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n4722) );
  INV_X1 U4057 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3071) );
  AND2_X1 U4058 ( .A1(n5648), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3005)
         );
  AND2_X2 U4059 ( .A1(n3006), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5179)
         );
  NAND3_X1 U4060 ( .A1(n5152), .A2(n3090), .A3(n4310), .ZN(n3059) );
  INV_X1 U4061 ( .A(n3405), .ZN(n3016) );
  OAI21_X1 U4062 ( .B1(n3333), .B2(n3308), .A(n3341), .ZN(n3309) );
  INV_X2 U4063 ( .A(n5243), .ZN(n3917) );
  NAND2_X1 U4064 ( .A1(n3659), .A2(n3646), .ZN(n5432) );
  AND2_X4 U4065 ( .A1(n4506), .A2(n3178), .ZN(n3381) );
  NAND2_X1 U4066 ( .A1(n4043), .A2(n3028), .ZN(n4002) );
  NAND2_X2 U4067 ( .A1(n4444), .A2(n4443), .ZN(n4460) );
  NAND2_X1 U4068 ( .A1(n5822), .A2(n3032), .ZN(n3030) );
  OR2_X1 U4069 ( .A1(n5823), .A2(n3034), .ZN(n3036) );
  INV_X1 U4070 ( .A(n6043), .ZN(n5928) );
  NAND2_X1 U4071 ( .A1(n4076), .A2(n3235), .ZN(n3323) );
  INV_X2 U4072 ( .A(n3517), .ZN(n3460) );
  NAND2_X2 U4073 ( .A1(n3513), .A2(n3514), .ZN(n3517) );
  NAND3_X1 U4074 ( .A1(n3061), .A2(n2972), .A3(PHYADDRPOINTER_REG_8__SCAN_IN), 
        .ZN(n3592) );
  NAND2_X1 U4075 ( .A1(n3692), .A2(n3001), .ZN(n3738) );
  NAND2_X1 U4076 ( .A1(n3405), .A2(n3077), .ZN(n3373) );
  AND2_X2 U4077 ( .A1(n4733), .A2(n3460), .ZN(n3535) );
  NAND2_X1 U4078 ( .A1(n3079), .A2(n4270), .ZN(n4521) );
  NAND2_X1 U4079 ( .A1(n4263), .A2(n4297), .ZN(n3079) );
  AND2_X1 U4080 ( .A1(n5659), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3082)
         );
  NAND2_X2 U4081 ( .A1(n4333), .A2(n4332), .ZN(n5684) );
  NAND2_X1 U4082 ( .A1(n3121), .A2(n3085), .ZN(n3084) );
  INV_X1 U4083 ( .A(n3332), .ZN(n3091) );
  NAND2_X2 U4084 ( .A1(n3325), .A2(n3282), .ZN(n3332) );
  AND2_X2 U4085 ( .A1(n2973), .A2(n4077), .ZN(n3343) );
  NAND2_X1 U4086 ( .A1(n3091), .A2(n3235), .ZN(n4077) );
  NAND2_X1 U4088 ( .A1(n3460), .A2(n3095), .ZN(n4287) );
  XNOR2_X1 U4089 ( .A(n3535), .B(n3473), .ZN(n4273) );
  NAND3_X1 U4090 ( .A1(n3441), .A2(n6747), .A3(n3374), .ZN(n3100) );
  XNOR2_X2 U4091 ( .A(n4286), .B(n6060), .ZN(n5000) );
  NAND2_X2 U4092 ( .A1(n3102), .A2(n4285), .ZN(n4286) );
  AND2_X1 U4093 ( .A1(n4474), .A2(n3327), .ZN(n3330) );
  OAI211_X1 U4094 ( .C1(n4474), .C2(n6747), .A(n3306), .B(n3305), .ZN(n3307)
         );
  NAND2_X1 U4095 ( .A1(n3236), .A2(n3237), .ZN(n4474) );
  NAND2_X1 U4096 ( .A1(n5418), .A2(n3104), .ZN(n5364) );
  NAND2_X1 U4097 ( .A1(n3917), .A2(n3166), .ZN(n4188) );
  NAND2_X1 U4098 ( .A1(n3917), .A2(n3106), .ZN(n5189) );
  OR2_X1 U4099 ( .A1(n5296), .A2(n3108), .ZN(n5270) );
  NAND2_X1 U4100 ( .A1(n5000), .A2(n3114), .ZN(n3112) );
  INV_X1 U4101 ( .A(n5000), .ZN(n3113) );
  INV_X1 U4102 ( .A(n4280), .ZN(n3114) );
  NAND2_X1 U4103 ( .A1(n5001), .A2(n5000), .ZN(n5147) );
  NAND2_X1 U4104 ( .A1(n3135), .A2(n3332), .ZN(n3324) );
  NAND3_X1 U4105 ( .A1(n3146), .A2(n3145), .A3(n4165), .ZN(n3144) );
  NAND2_X1 U4106 ( .A1(n3154), .A2(n3153), .ZN(n4616) );
  NAND2_X1 U4107 ( .A1(n4545), .A2(n4546), .ZN(n4544) );
  AND2_X2 U4108 ( .A1(n3155), .A2(n4719), .ZN(n3295) );
  AND2_X2 U4109 ( .A1(n3155), .A2(n3178), .ZN(n3242) );
  AND2_X2 U4110 ( .A1(n3171), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3155)
         );
  NAND3_X1 U4111 ( .A1(n3301), .A2(n3300), .A3(n3997), .ZN(n3342) );
  NAND2_X1 U4112 ( .A1(n5418), .A2(n5419), .ZN(n5403) );
  NAND3_X1 U4113 ( .A1(n3358), .A2(n3357), .A3(n3356), .ZN(n3362) );
  OR2_X2 U4114 ( .A1(n5201), .A2(n4181), .ZN(n4183) );
  AOI21_X1 U4115 ( .B1(n5209), .B2(n6370), .A(n5192), .ZN(n5193) );
  INV_X1 U4116 ( .A(n5842), .ZN(n5572) );
  INV_X1 U4117 ( .A(n5665), .ZN(n5606) );
  AOI22_X1 U4118 ( .A1(n3293), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3209) );
  AND2_X1 U4119 ( .A1(n4618), .A2(n4617), .ZN(n6432) );
  NAND2_X1 U4120 ( .A1(n4099), .A2(n4098), .ZN(n4618) );
  INV_X1 U4121 ( .A(n4616), .ZN(n4099) );
  INV_X1 U4122 ( .A(n3349), .ZN(n3236) );
  NAND2_X1 U4123 ( .A1(n3235), .A2(n3282), .ZN(n3349) );
  AND3_X1 U4124 ( .A1(n3331), .A2(n3330), .A3(n4080), .ZN(n3338) );
  INV_X2 U4125 ( .A(n4177), .ZN(n5350) );
  INV_X1 U4126 ( .A(n4200), .ZN(n4244) );
  OAI21_X1 U4127 ( .B1(n5590), .B2(n5593), .A(n5189), .ZN(n4200) );
  INV_X1 U4128 ( .A(READY_N), .ZN(n6692) );
  NAND2_X1 U4129 ( .A1(n6302), .A2(n5591), .ZN(n6295) );
  INV_X1 U4130 ( .A(n6295), .ZN(n4196) );
  INV_X1 U4131 ( .A(n5588), .ZN(n6299) );
  INV_X1 U4132 ( .A(n6345), .ZN(n6369) );
  AND2_X1 U4133 ( .A1(n3534), .A2(n3533), .ZN(n3168) );
  AND2_X1 U4134 ( .A1(n3345), .A2(n3346), .ZN(n3170) );
  INV_X1 U4135 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6844) );
  NAND2_X1 U4136 ( .A1(n6657), .A2(n5093), .ZN(n6672) );
  INV_X1 U4137 ( .A(DATAI_31_), .ZN(n6784) );
  INV_X1 U4138 ( .A(DATAI_7_), .ZN(n4660) );
  INV_X1 U4139 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4032) );
  AOI21_X1 U4140 ( .B1(n4245), .B2(n3685), .A(n3524), .ZN(n4533) );
  INV_X1 U4141 ( .A(n3268), .ZN(n3396) );
  AOI22_X1 U4142 ( .A1(n3375), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3289) );
  INV_X1 U4143 ( .A(n4252), .ZN(n4246) );
  AOI22_X1 U4144 ( .A1(n3293), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3172) );
  AND4_X1 U4145 ( .A1(n3226), .A2(n3225), .A3(n3224), .A4(n3223), .ZN(n3232)
         );
  NAND2_X1 U4146 ( .A1(n3268), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3272)
         );
  CLKBUF_X2 U4147 ( .A(n3293), .Z(n3921) );
  NAND2_X1 U4148 ( .A1(n2963), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3190)
         );
  INV_X1 U4149 ( .A(n5246), .ZN(n3916) );
  INV_X1 U4150 ( .A(n5433), .ZN(n3658) );
  INV_X1 U4151 ( .A(n4297), .ZN(n4312) );
  AND4_X1 U4152 ( .A1(n3277), .A2(n3276), .A3(n3275), .A4(n3274), .ZN(n3278)
         );
  AND2_X1 U4153 ( .A1(n3990), .A2(n4009), .ZN(n4054) );
  AND2_X1 U4154 ( .A1(n3255), .A2(n3254), .ZN(n3256) );
  INV_X1 U4155 ( .A(n5366), .ZN(n3740) );
  AND2_X1 U4156 ( .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3852) );
  INV_X1 U4157 ( .A(n5157), .ZN(n3607) );
  OR2_X1 U4158 ( .A1(n3702), .A2(n3332), .ZN(n4510) );
  AND2_X1 U4159 ( .A1(n5277), .A2(n4220), .ZN(n5247) );
  INV_X1 U4160 ( .A(n5511), .ZN(n5211) );
  INV_X1 U4161 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4228) );
  AND2_X1 U4162 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5648) );
  INV_X1 U4163 ( .A(n5687), .ZN(n4332) );
  AND2_X1 U4164 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5931) );
  INV_X1 U4165 ( .A(n4615), .ZN(n4098) );
  NAND2_X1 U4166 ( .A1(n4045), .A2(n4044), .ZN(n4046) );
  AND2_X1 U4167 ( .A1(n6143), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4646)
         );
  INV_X1 U4168 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5262) );
  AND2_X1 U4169 ( .A1(n5343), .A2(n4212), .ZN(n5305) );
  INV_X1 U4170 ( .A(n5530), .ZN(n5532) );
  OR2_X1 U4171 ( .A1(n5547), .A2(n5093), .ZN(n6251) );
  AND2_X1 U4172 ( .A1(n5311), .A2(n5299), .ZN(n4158) );
  AND2_X1 U4173 ( .A1(n4140), .A2(n4139), .ZN(n5397) );
  INV_X1 U4174 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n6754) );
  INV_X1 U4175 ( .A(n5206), .ZN(n5207) );
  OR2_X1 U4176 ( .A1(n6026), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5676)
         );
  AND2_X1 U4177 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5910) );
  INV_X1 U4178 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5973) );
  INV_X1 U4179 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5988) );
  INV_X1 U4180 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6046) );
  INV_X1 U4181 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6062) );
  OR2_X1 U4182 ( .A1(n4237), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6412) );
  AND2_X1 U4183 ( .A1(n4493), .A2(n4492), .ZN(n6198) );
  OR2_X1 U4184 ( .A1(n6671), .A2(n4820), .ZN(n4825) );
  AND2_X1 U4185 ( .A1(n5092), .A2(n6463), .ZN(n5130) );
  NAND2_X1 U4186 ( .A1(n6462), .A2(n4642), .ZN(n6703) );
  NOR2_X1 U4187 ( .A1(n6677), .A2(n4820), .ZN(n4644) );
  INV_X1 U4188 ( .A(DATAI_16_), .ZN(n4688) );
  AND2_X1 U4189 ( .A1(n4748), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4786)
         );
  NAND2_X1 U4190 ( .A1(n3446), .A2(n3445), .ZN(n4857) );
  INV_X1 U4191 ( .A(DATAI_29_), .ZN(n4641) );
  AND2_X1 U4192 ( .A1(n6144), .A2(n6552), .ZN(n4749) );
  OR2_X1 U4193 ( .A1(n4421), .A2(n6223), .ZN(n6221) );
  NAND2_X1 U4194 ( .A1(n4464), .A2(n6221), .ZN(n6690) );
  OR2_X1 U4195 ( .A1(n5848), .A2(n5570), .ZN(n4234) );
  INV_X1 U4196 ( .A(n6276), .ZN(n6260) );
  AND2_X1 U4197 ( .A1(n5553), .A2(n4527), .ZN(n6279) );
  OR2_X1 U4198 ( .A1(n6302), .A2(n4184), .ZN(n4185) );
  INV_X1 U4199 ( .A(n6302), .ZN(n5584) );
  NOR2_X2 U4200 ( .A1(n5641), .A2(n4439), .ZN(n5636) );
  AND2_X1 U4201 ( .A1(n6321), .A2(n3328), .ZN(n6306) );
  AND2_X1 U4202 ( .A1(n4909), .A2(n6747), .ZN(n6331) );
  INV_X1 U4203 ( .A(DATAI_6_), .ZN(n4666) );
  INV_X1 U4204 ( .A(n4569), .ZN(n4572) );
  AND2_X1 U4205 ( .A1(n5431), .A2(n5434), .ZN(n6291) );
  NAND2_X1 U4206 ( .A1(n6345), .A2(n4238), .ZN(n5816) );
  INV_X1 U4207 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5956) );
  INV_X1 U4208 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6036) );
  AND2_X1 U4209 ( .A1(n5153), .A2(n5152), .ZN(n6396) );
  AND2_X1 U4210 ( .A1(n6435), .A2(n6441), .ZN(n6059) );
  INV_X1 U4211 ( .A(n6016), .ZN(n6434) );
  NAND2_X1 U4212 ( .A1(n4639), .A2(n6747), .ZN(n5055) );
  NAND2_X1 U4213 ( .A1(n4932), .A2(n4931), .ZN(n4957) );
  OAI211_X1 U4214 ( .C1(n4830), .C2(n4829), .A(n6513), .B(n4828), .ZN(n4853)
         );
  NOR2_X1 U4215 ( .A1(n4825), .A2(n4642), .ZN(n4926) );
  OAI21_X1 U4216 ( .B1(n6079), .B2(n6082), .A(n6476), .ZN(n6104) );
  INV_X1 U4217 ( .A(n6460), .ZN(n5134) );
  OAI211_X1 U4218 ( .C1(n6515), .C2(n5092), .A(n4793), .B(n6513), .ZN(n4816)
         );
  INV_X1 U4219 ( .A(n6470), .ZN(n6497) );
  OAI211_X1 U4220 ( .C1(n6515), .C2(n6143), .A(n4651), .B(n6513), .ZN(n4692)
         );
  OAI211_X1 U4221 ( .C1(n5020), .C2(n6553), .A(n5019), .B(n5018), .ZN(n5045)
         );
  OAI21_X1 U4222 ( .B1(n6562), .B2(n6561), .A(n6560), .ZN(n6587) );
  AND2_X1 U4223 ( .A1(n5089), .A2(n6671), .ZN(n6586) );
  OAI211_X1 U4224 ( .C1(n6515), .C2(n5056), .A(n4759), .B(n6513), .ZN(n4782)
         );
  INV_X1 U4225 ( .A(n4862), .ZN(n4898) );
  NOR2_X1 U4226 ( .A1(n6358), .A2(n4673), .ZN(n6595) );
  NOR2_X1 U4227 ( .A1(n6358), .A2(n4656), .ZN(n6616) );
  NOR2_X1 U4228 ( .A1(n6358), .A2(n4661), .ZN(n6639) );
  AND2_X1 U4229 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n4909) );
  INV_X1 U4230 ( .A(STATE_REG_0__SCAN_IN), .ZN(n4352) );
  INV_X1 U4231 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6228) );
  INV_X1 U4232 ( .A(n6267), .ZN(n6282) );
  INV_X1 U4233 ( .A(n5544), .ZN(n5561) );
  NAND2_X1 U4234 ( .A1(n5665), .A2(n6299), .ZN(n4199) );
  INV_X1 U4235 ( .A(n5728), .ZN(n5625) );
  INV_X1 U4236 ( .A(n6291), .ZN(n5644) );
  INV_X1 U4237 ( .A(DATAI_3_), .ZN(n4682) );
  INV_X1 U4238 ( .A(n6306), .ZN(n5008) );
  INV_X1 U4239 ( .A(n6331), .ZN(n6335) );
  INV_X1 U4240 ( .A(UWORD_REG_9__SCAN_IN), .ZN(n6816) );
  INV_X1 U4241 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6826) );
  INV_X1 U4242 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6738) );
  INV_X1 U4243 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6420) );
  INV_X1 U4244 ( .A(n4926), .ZN(n4963) );
  AOI22_X1 U4245 ( .A1(n4827), .A2(n4829), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4824), .ZN(n4856) );
  INV_X1 U4246 ( .A(n6075), .ZN(n6110) );
  INV_X1 U4247 ( .A(n6456), .ZN(n6137) );
  AOI22_X1 U4248 ( .A1(n4792), .A2(n4787), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5092), .ZN(n4819) );
  NAND2_X1 U4249 ( .A1(n6462), .A2(n6461), .ZN(n6702) );
  AOI21_X1 U4250 ( .B1(n6516), .B2(STATE2_REG_2__SCAN_IN), .A(n6505), .ZN(
        n6706) );
  NAND2_X1 U4251 ( .A1(n6370), .A2(DATAI_19_), .ZN(n6525) );
  AOI22_X1 U4252 ( .A1(n4649), .A2(n4637), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6143), .ZN(n4695) );
  AOI22_X1 U4253 ( .A1(n5017), .A2(n6553), .B1(n6464), .B2(n5014), .ZN(n5048)
         );
  AOI22_X1 U4254 ( .A1(n6559), .A2(n6561), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6556), .ZN(n6591) );
  INV_X1 U4255 ( .A(n6624), .ZN(n6535) );
  INV_X1 U4256 ( .A(n6593), .ZN(n6705) );
  INV_X1 U4257 ( .A(n6629), .ZN(n6583) );
  NOR2_X1 U4258 ( .A1(n4861), .A2(n4860), .ZN(n4901) );
  AOI21_X1 U4259 ( .B1(n4736), .B2(n4739), .A(n4735), .ZN(n6646) );
  INV_X1 U4260 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6244) );
  INV_X1 U4261 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6815) );
  INV_X1 U4262 ( .A(REIP_REG_24__SCAN_IN), .ZN(n5293) );
  AND2_X1 U4263 ( .A1(n4352), .A2(STATE_REG_1__SCAN_IN), .ZN(n4373) );
  NAND2_X1 U4264 ( .A1(n4199), .A2(n4198), .ZN(U2831) );
  AND2_X2 U4265 ( .A1(n3177), .A2(n3176), .ZN(n3375) );
  AND2_X2 U4266 ( .A1(n3177), .A2(n4719), .ZN(n3288) );
  AOI22_X1 U4267 ( .A1(n3375), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3175) );
  INV_X1 U4268 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3171) );
  AND2_X4 U4269 ( .A1(n3177), .A2(n3178), .ZN(n3286) );
  AND2_X4 U4270 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4507) );
  AND2_X2 U4271 ( .A1(n3178), .A2(n4507), .ZN(n3293) );
  AND2_X4 U4272 ( .A1(n4719), .A2(n4507), .ZN(n3273) );
  AND2_X2 U4273 ( .A1(n3176), .A2(n4507), .ZN(n3380) );
  AND2_X2 U4274 ( .A1(n5179), .A2(n3177), .ZN(n3287) );
  AOI22_X1 U4275 ( .A1(n3380), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3182) );
  AND2_X4 U4276 ( .A1(n5179), .A2(n4507), .ZN(n3268) );
  AOI22_X1 U4277 ( .A1(n3242), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4278 ( .A1(n3926), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3381), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3180) );
  NAND2_X1 U4279 ( .A1(n3380), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3186) );
  NAND2_X1 U4280 ( .A1(n2962), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3185) );
  NAND2_X1 U4281 ( .A1(n3242), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3184) );
  NAND2_X1 U4282 ( .A1(n3926), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3183) );
  NAND2_X1 U4283 ( .A1(n3243), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3189) );
  NAND2_X1 U4284 ( .A1(n3288), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3188)
         );
  NAND2_X1 U4285 ( .A1(n3293), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3187) );
  NAND2_X1 U4287 ( .A1(n3286), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3194) );
  NAND2_X1 U4288 ( .A1(n3375), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3193) );
  NAND2_X1 U4289 ( .A1(n3273), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3191)
         );
  NAND2_X1 U4291 ( .A1(n3268), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3198)
         );
  NAND2_X1 U4292 ( .A1(n3287), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3197) );
  NAND2_X1 U4293 ( .A1(n3381), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3196) );
  NAND2_X1 U4294 ( .A1(n3263), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3195)
         );
  AND4_X2 U4295 ( .A1(n3198), .A2(n3197), .A3(n3196), .A4(n3195), .ZN(n3199)
         );
  NAND4_X4 U4296 ( .A1(n3202), .A2(n3201), .A3(n3200), .A4(n3199), .ZN(n3322)
         );
  INV_X1 U4297 ( .A(n4074), .ZN(n3237) );
  AOI22_X1 U4298 ( .A1(n3380), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3207) );
  AND2_X1 U4299 ( .A1(n3268), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3203) );
  AOI22_X1 U4300 ( .A1(n3926), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3381), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3205) );
  AOI22_X1 U4301 ( .A1(n3263), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        INSTQUEUE_REG_10__4__SCAN_IN), .B2(n2963), .ZN(n3204) );
  AOI22_X1 U4302 ( .A1(n3375), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3211) );
  INV_X1 U4303 ( .A(n3333), .ZN(n3235) );
  NAND2_X1 U4304 ( .A1(n3242), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3218) );
  NAND2_X1 U4305 ( .A1(n3380), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U4306 ( .A1(n3287), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3216) );
  NAND2_X1 U4307 ( .A1(n3268), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3215)
         );
  NAND2_X1 U4308 ( .A1(n3286), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3222) );
  NAND2_X1 U4309 ( .A1(n2962), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U4310 ( .A1(n3273), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3220)
         );
  NAND2_X1 U4311 ( .A1(n3375), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3219) );
  NAND2_X1 U4312 ( .A1(n3288), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3226)
         );
  NAND2_X1 U4313 ( .A1(n3243), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3225) );
  NAND2_X1 U4314 ( .A1(n3295), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3224)
         );
  NAND2_X1 U4315 ( .A1(n3293), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3223) );
  NAND2_X1 U4316 ( .A1(n3926), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3230) );
  NAND2_X1 U4317 ( .A1(n2963), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3229)
         );
  NAND2_X1 U4318 ( .A1(n3381), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3228) );
  NAND2_X1 U4319 ( .A1(n3263), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3227)
         );
  AOI22_X1 U4320 ( .A1(n3375), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3241) );
  AOI22_X1 U4321 ( .A1(n3926), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3239) );
  AOI22_X1 U4322 ( .A1(n3295), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3238) );
  AOI22_X1 U4323 ( .A1(n3242), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3381), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3246) );
  AOI22_X1 U4324 ( .A1(n3380), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3263), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3245) );
  AOI22_X1 U4325 ( .A1(n3243), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3244) );
  NAND2_X2 U4326 ( .A1(n3249), .A2(n3248), .ZN(n3308) );
  BUF_X8 U4327 ( .A(n3286), .Z(n3956) );
  AOI22_X1 U4328 ( .A1(n3956), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        INSTQUEUE_REG_4__7__SCAN_IN), .B2(n2962), .ZN(n3253) );
  AOI22_X1 U4329 ( .A1(n3243), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3295), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3252) );
  AOI22_X1 U4330 ( .A1(n3863), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3381), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3251) );
  AOI22_X1 U4331 ( .A1(n2963), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3250) );
  AOI22_X1 U4332 ( .A1(n3293), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3257) );
  AOI22_X1 U4333 ( .A1(n3287), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3263), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3255) );
  AOI22_X1 U4334 ( .A1(n3380), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3254) );
  NAND2_X1 U4335 ( .A1(n3243), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3262) );
  NAND2_X1 U4336 ( .A1(n3286), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3261) );
  NAND2_X1 U4337 ( .A1(n3295), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3260)
         );
  NAND2_X1 U4338 ( .A1(n2962), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3259) );
  NAND2_X1 U4339 ( .A1(n2963), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3267)
         );
  NAND2_X1 U4340 ( .A1(n3380), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3266) );
  NAND2_X1 U4341 ( .A1(n3263), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3264)
         );
  NAND2_X1 U4342 ( .A1(n3242), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3271) );
  NAND2_X1 U4343 ( .A1(n3926), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3270) );
  NAND2_X1 U4344 ( .A1(n3381), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3269) );
  NAND2_X1 U4345 ( .A1(n3288), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3277)
         );
  NAND2_X1 U4346 ( .A1(n3375), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3276) );
  NAND2_X1 U4347 ( .A1(n3293), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3275) );
  NAND2_X1 U4348 ( .A1(n3273), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3274)
         );
  NAND4_X4 U4349 ( .A1(n3281), .A2(n3280), .A3(n3279), .A4(n3278), .ZN(n3328)
         );
  NAND2_X1 U4350 ( .A1(n3350), .A2(n3328), .ZN(n4070) );
  NAND2_X1 U4351 ( .A1(n3346), .A2(n3332), .ZN(n3283) );
  OAI21_X1 U4352 ( .B1(n6747), .B2(n4070), .A(n3283), .ZN(n3284) );
  NAND2_X1 U4353 ( .A1(n3323), .A2(n3284), .ZN(n3306) );
  NAND2_X1 U4354 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n4347) );
  NAND2_X1 U4355 ( .A1(n3350), .A2(n4208), .ZN(n3345) );
  NAND3_X1 U4356 ( .A1(n3997), .A2(n3345), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3303) );
  AOI22_X1 U4357 ( .A1(n3286), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4358 ( .A1(n3287), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3263), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4359 ( .A1(n3380), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3381), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3290) );
  AOI22_X1 U4360 ( .A1(n3243), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4361 ( .A1(n3863), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4362 ( .A1(n2963), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3926), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3297) );
  NAND2_X1 U4363 ( .A1(n3311), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3302) );
  OAI211_X1 U4364 ( .C1(n3315), .C2(n3350), .A(n3303), .B(n3302), .ZN(n3304)
         );
  INV_X1 U4365 ( .A(n3304), .ZN(n3305) );
  INV_X1 U4366 ( .A(n3307), .ZN(n3319) );
  INV_X1 U4367 ( .A(n3309), .ZN(n3310) );
  NAND2_X1 U4368 ( .A1(n3311), .A2(n3349), .ZN(n3313) );
  NAND2_X1 U4369 ( .A1(n3348), .A2(n3388), .ZN(n3318) );
  INV_X1 U4370 ( .A(n3343), .ZN(n3316) );
  NAND3_X2 U4371 ( .A1(n3319), .A2(n3318), .A3(n3317), .ZN(n3363) );
  NAND2_X1 U4372 ( .A1(n3363), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3321) );
  MUX2_X1 U4373 ( .A(n4062), .B(n4237), .S(n6463), .Z(n3320) );
  NAND2_X1 U4374 ( .A1(n3321), .A2(n3320), .ZN(n3406) );
  NAND2_X1 U4375 ( .A1(n3348), .A2(n3340), .ZN(n4083) );
  INV_X1 U4376 ( .A(n4070), .ZN(n4302) );
  OAI21_X1 U4377 ( .B1(n3323), .B2(n3324), .A(n4302), .ZN(n3331) );
  NAND2_X1 U4378 ( .A1(n5177), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6653) );
  AOI21_X1 U4379 ( .B1(n3326), .B2(n4253), .A(n6653), .ZN(n3327) );
  NAND2_X1 U4380 ( .A1(n3701), .A2(n3328), .ZN(n4049) );
  AND2_X1 U4381 ( .A1(n4049), .A2(n5491), .ZN(n3329) );
  OR2_X1 U4382 ( .A1(n3349), .A2(n3328), .ZN(n4051) );
  BUF_X1 U4383 ( .A(n3333), .Z(n3334) );
  NAND2_X1 U4384 ( .A1(n3332), .A2(n3334), .ZN(n3335) );
  NAND2_X1 U4385 ( .A1(n3343), .A2(n3335), .ZN(n3336) );
  NAND2_X1 U4386 ( .A1(n3336), .A2(n3322), .ZN(n3337) );
  NAND3_X1 U4387 ( .A1(n4083), .A2(n3338), .A3(n3337), .ZN(n3407) );
  AND2_X2 U4388 ( .A1(n3406), .A2(n3407), .ZN(n3405) );
  INV_X1 U4389 ( .A(n3363), .ZN(n3355) );
  NOR2_X1 U4390 ( .A1(n3342), .A2(n3334), .ZN(n3344) );
  NAND2_X1 U4391 ( .A1(n3344), .A2(n3343), .ZN(n4047) );
  INV_X1 U4392 ( .A(n4047), .ZN(n3347) );
  NAND2_X1 U4393 ( .A1(n3347), .A2(n3170), .ZN(n3358) );
  INV_X1 U4394 ( .A(n3348), .ZN(n3351) );
  INV_X1 U4395 ( .A(n4237), .ZN(n3444) );
  NAND2_X1 U4396 ( .A1(n3444), .A2(n6464), .ZN(n3353) );
  INV_X1 U4397 ( .A(n4062), .ZN(n3366) );
  NAND2_X1 U4398 ( .A1(n3366), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3352) );
  INV_X1 U4399 ( .A(n3359), .ZN(n3360) );
  OR2_X1 U4400 ( .A1(n3360), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3361)
         );
  NAND2_X1 U4401 ( .A1(n3362), .A2(n3361), .ZN(n3390) );
  NAND2_X1 U4402 ( .A1(n3373), .A2(n3390), .ZN(n3369) );
  BUF_X2 U4403 ( .A(n3363), .Z(n3442) );
  NAND2_X1 U4404 ( .A1(n3442), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3368) );
  NAND2_X1 U4405 ( .A1(n4010), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U4406 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3364) );
  NAND2_X1 U4407 ( .A1(n3364), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3365) );
  OAI21_X1 U4408 ( .B1(n6117), .B2(n6463), .A(n3365), .ZN(n4863) );
  AOI22_X1 U4409 ( .A1(n4863), .A2(n3444), .B1(n3366), .B2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3367) );
  NAND2_X1 U4410 ( .A1(n3368), .A2(n3367), .ZN(n3370) );
  INV_X1 U4411 ( .A(n3370), .ZN(n3371) );
  AND2_X1 U4412 ( .A1(n3371), .A2(n3390), .ZN(n3372) );
  NAND2_X1 U4413 ( .A1(n3373), .A2(n3372), .ZN(n3374) );
  AOI22_X1 U4414 ( .A1(n3825), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4415 ( .A1(n3963), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3378) );
  INV_X1 U4416 ( .A(n2962), .ZN(n3785) );
  INV_X2 U4417 ( .A(n3785), .ZN(n3939) );
  AOI22_X1 U4418 ( .A1(n3939), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4419 ( .A1(n3921), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3376) );
  NAND4_X1 U4420 ( .A1(n3379), .A2(n3378), .A3(n3377), .A4(n3376), .ZN(n3387)
         );
  INV_X1 U4421 ( .A(n3380), .ZN(n5181) );
  AOI22_X1 U4422 ( .A1(n3957), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3385) );
  AOI22_X1 U4423 ( .A1(n3958), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4424 ( .A1(n3944), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4425 ( .A1(n3728), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3382) );
  NAND4_X1 U4426 ( .A1(n3385), .A2(n3384), .A3(n3383), .A4(n3382), .ZN(n3386)
         );
  XNOR2_X1 U4427 ( .A(n3405), .B(n3391), .ZN(n4504) );
  NAND2_X1 U4428 ( .A1(n4504), .A2(n6747), .ZN(n3404) );
  INV_X1 U4429 ( .A(n3447), .ZN(n4064) );
  AOI22_X1 U4430 ( .A1(n3939), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3728), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4431 ( .A1(n3944), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3958), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4432 ( .A1(n2965), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3393) );
  AOI22_X1 U4433 ( .A1(n3965), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3392) );
  NAND4_X1 U4434 ( .A1(n3395), .A2(n3394), .A3(n3393), .A4(n3392), .ZN(n3402)
         );
  AOI22_X1 U4435 ( .A1(n3963), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4436 ( .A1(n3957), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3399) );
  AOI22_X1 U4437 ( .A1(n3966), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3381), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3398) );
  AOI22_X1 U4438 ( .A1(n3825), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3397) );
  NAND4_X1 U4439 ( .A1(n3400), .A2(n3399), .A3(n3398), .A4(n3397), .ZN(n3401)
         );
  NAND2_X1 U4440 ( .A1(n4064), .A2(n4265), .ZN(n3403) );
  INV_X1 U4442 ( .A(n3406), .ZN(n3409) );
  INV_X1 U4443 ( .A(n3407), .ZN(n3408) );
  NAND2_X1 U4444 ( .A1(n3409), .A2(n3408), .ZN(n3410) );
  AOI22_X1 U4445 ( .A1(n3825), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3414) );
  AOI22_X1 U4446 ( .A1(n3965), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3863), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3413) );
  AOI22_X1 U4447 ( .A1(n3939), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3412) );
  INV_X1 U4448 ( .A(n3728), .ZN(n3788) );
  AOI22_X1 U4449 ( .A1(n3728), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3411) );
  NAND4_X1 U4450 ( .A1(n3414), .A2(n3413), .A3(n3412), .A4(n3411), .ZN(n3421)
         );
  AOI22_X1 U4451 ( .A1(n3295), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3419) );
  AOI22_X1 U4452 ( .A1(n3957), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3418) );
  AOI22_X1 U4453 ( .A1(n3268), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3381), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3417) );
  AOI22_X1 U4454 ( .A1(n3963), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3416) );
  NAND4_X1 U4455 ( .A1(n3419), .A2(n3418), .A3(n3417), .A4(n3416), .ZN(n3420)
         );
  NOR2_X1 U4456 ( .A1(n3447), .A2(n4315), .ZN(n3437) );
  NAND2_X1 U4457 ( .A1(n3235), .A2(n4315), .ZN(n3433) );
  AOI22_X1 U4458 ( .A1(n3963), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4459 ( .A1(n3939), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3424) );
  AOI22_X1 U4460 ( .A1(n3957), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4461 ( .A1(n3958), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3422) );
  NAND4_X1 U4462 ( .A1(n3425), .A2(n3424), .A3(n3423), .A4(n3422), .ZN(n3431)
         );
  AOI22_X1 U4463 ( .A1(n3965), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4464 ( .A1(n3295), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4465 ( .A1(n3728), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4466 ( .A1(n3825), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3426) );
  NAND4_X1 U4467 ( .A1(n3429), .A2(n3428), .A3(n3427), .A4(n3426), .ZN(n3430)
         );
  INV_X1 U4468 ( .A(n4266), .ZN(n3432) );
  NOR2_X1 U4469 ( .A1(n4266), .A2(n6747), .ZN(n3435) );
  NAND2_X1 U4470 ( .A1(n4039), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3434) );
  OAI211_X1 U4471 ( .C1(n3346), .C2(n3435), .A(n3434), .B(n3433), .ZN(n3497)
         );
  INV_X1 U4472 ( .A(n4265), .ZN(n3440) );
  NAND2_X1 U4473 ( .A1(n4039), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3439) );
  INV_X1 U4474 ( .A(n3437), .ZN(n3438) );
  OAI211_X1 U4475 ( .C1(n3440), .C2(n3315), .A(n3439), .B(n3438), .ZN(n3488)
         );
  NAND2_X1 U4476 ( .A1(n3442), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3446) );
  NAND3_X1 U4477 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4859) );
  AOI21_X1 U4478 ( .B1(n6700), .B2(n6681), .A(n6636), .ZN(n5098) );
  NOR2_X1 U4479 ( .A1(n4062), .A2(n6681), .ZN(n3443) );
  AOI21_X1 U4480 ( .B1(n5098), .B2(n3444), .A(n3443), .ZN(n3445) );
  NAND2_X1 U4481 ( .A1(n4635), .A2(n6747), .ZN(n3459) );
  AOI22_X1 U4482 ( .A1(n3825), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4483 ( .A1(n3963), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4484 ( .A1(n3939), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4485 ( .A1(n3921), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3448) );
  NAND4_X1 U4486 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), .ZN(n3457)
         );
  INV_X2 U4487 ( .A(n5181), .ZN(n3957) );
  AOI22_X1 U4488 ( .A1(n3957), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4489 ( .A1(n3958), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4490 ( .A1(n3944), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4491 ( .A1(n3900), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3452) );
  NAND4_X1 U4492 ( .A1(n3455), .A2(n3454), .A3(n3453), .A4(n3452), .ZN(n3456)
         );
  AOI22_X1 U4493 ( .A1(n4039), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4013), 
        .B2(n4274), .ZN(n3458) );
  NAND2_X1 U4494 ( .A1(n4039), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3472) );
  AOI22_X1 U4495 ( .A1(n3825), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4496 ( .A1(n3963), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3463) );
  AOI22_X1 U4497 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3939), .B1(n3956), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3462) );
  AOI22_X1 U4498 ( .A1(n3921), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3461) );
  NAND4_X1 U4499 ( .A1(n3464), .A2(n3463), .A3(n3462), .A4(n3461), .ZN(n3470)
         );
  AOI22_X1 U4500 ( .A1(n3957), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4501 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n3863), .B1(n3966), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4502 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n3944), .B1(n3864), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4503 ( .A1(n3900), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3465) );
  NAND4_X1 U4504 ( .A1(n3468), .A2(n3467), .A3(n3466), .A4(n3465), .ZN(n3469)
         );
  NAND2_X1 U4505 ( .A1(n4013), .A2(n4290), .ZN(n3471) );
  NAND2_X1 U4506 ( .A1(n3472), .A2(n3471), .ZN(n3534) );
  INV_X1 U4507 ( .A(n3534), .ZN(n3473) );
  AOI22_X1 U4508 ( .A1(n3825), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3477) );
  AOI22_X1 U4509 ( .A1(n3963), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3476) );
  AOI22_X1 U4510 ( .A1(n3939), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3475) );
  AOI22_X1 U4511 ( .A1(n3921), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3474) );
  NAND4_X1 U4512 ( .A1(n3477), .A2(n3476), .A3(n3475), .A4(n3474), .ZN(n3483)
         );
  AOI22_X1 U4513 ( .A1(n3957), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3481) );
  AOI22_X1 U4514 ( .A1(n3958), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3480) );
  INV_X1 U4515 ( .A(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n6840) );
  AOI22_X1 U4516 ( .A1(n3944), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3479) );
  AOI22_X1 U4517 ( .A1(n3900), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3478) );
  NAND4_X1 U4518 ( .A1(n3481), .A2(n3480), .A3(n3479), .A4(n3478), .ZN(n3482)
         );
  AOI22_X1 U4519 ( .A1(n4039), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4013), 
        .B2(n4289), .ZN(n3532) );
  XNOR2_X2 U4520 ( .A(n3484), .B(n3533), .ZN(n4281) );
  NAND2_X1 U4521 ( .A1(n3326), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3516) );
  NAND2_X1 U4522 ( .A1(n4281), .A2(n3685), .ZN(n3487) );
  NAND2_X1 U4523 ( .A1(n3529), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3547)
         );
  XNOR2_X1 U4524 ( .A(n3547), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U4525 ( .A1(n6657), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5188) );
  OAI22_X1 U4526 ( .A1(n5495), .A2(n3797), .B1(n5188), .B2(n5498), .ZN(n3485)
         );
  AOI21_X1 U4527 ( .B1(n3546), .B2(EAX_REG_5__SCAN_IN), .A(n3485), .ZN(n3486)
         );
  NAND2_X1 U4528 ( .A1(n3487), .A2(n3486), .ZN(n4545) );
  XNOR2_X1 U4529 ( .A(n3489), .B(n3488), .ZN(n3491) );
  XNOR2_X1 U4530 ( .A(n3491), .B(n3490), .ZN(n4263) );
  NAND2_X1 U4531 ( .A1(n4263), .A2(n3685), .ZN(n3495) );
  AOI22_X1 U4532 ( .A1(n3977), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6657), .ZN(n3493) );
  NAND2_X1 U4533 ( .A1(n3518), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3492) );
  AND2_X1 U4534 ( .A1(n3493), .A2(n3492), .ZN(n3494) );
  NAND2_X1 U4535 ( .A1(n3495), .A2(n3494), .ZN(n4596) );
  INV_X1 U4536 ( .A(n3497), .ZN(n3498) );
  XNOR2_X1 U4537 ( .A(n3499), .B(n3498), .ZN(n3500) );
  NAND2_X1 U4538 ( .A1(n4729), .A2(n3326), .ZN(n4499) );
  OR2_X1 U4539 ( .A1(n3501), .A2(n3516), .ZN(n3505) );
  AOI22_X1 U4540 ( .A1(n3977), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6657), .ZN(n3503) );
  NAND2_X1 U4541 ( .A1(n3518), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3502) );
  AND2_X1 U4542 ( .A1(n3503), .A2(n3502), .ZN(n3504) );
  NAND2_X1 U4543 ( .A1(n3505), .A2(n3504), .ZN(n3507) );
  AND2_X1 U4544 ( .A1(n3507), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3506) );
  NAND2_X1 U4545 ( .A1(n4499), .A2(n3506), .ZN(n4502) );
  INV_X1 U4546 ( .A(n3507), .ZN(n4500) );
  NAND2_X1 U4547 ( .A1(n4500), .A2(n3982), .ZN(n3508) );
  NAND2_X1 U4548 ( .A1(n4502), .A2(n3508), .ZN(n4598) );
  NAND2_X1 U4549 ( .A1(n3518), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3512) );
  INV_X1 U4550 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5535) );
  OAI21_X1 U4551 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3519), .ZN(n6374) );
  NAND2_X1 U4552 ( .A1(n3982), .A2(n6374), .ZN(n3509) );
  OAI21_X1 U4553 ( .B1(n5535), .B2(n5188), .A(n3509), .ZN(n3510) );
  AOI21_X1 U4554 ( .B1(n3546), .B2(EAX_REG_2__SCAN_IN), .A(n3510), .ZN(n3511)
         );
  NOR2_X2 U4555 ( .A1(n4597), .A2(n4609), .ZN(n4534) );
  OR2_X1 U4556 ( .A1(n3514), .A2(n3513), .ZN(n3515) );
  NAND2_X1 U4557 ( .A1(n3517), .A2(n3515), .ZN(n4251) );
  OAI21_X1 U4558 ( .B1(n4251), .B2(n3516), .A(n5188), .ZN(n4611) );
  NAND2_X1 U4559 ( .A1(n4597), .A2(n4609), .ZN(n4535) );
  INV_X1 U4560 ( .A(n3518), .ZN(n3528) );
  INV_X1 U4561 ( .A(n3529), .ZN(n3521) );
  NAND2_X1 U4562 ( .A1(n3060), .A2(n3519), .ZN(n3520) );
  NAND2_X1 U4563 ( .A1(n3521), .A2(n3520), .ZN(n5522) );
  AOI22_X1 U4564 ( .A1(n5522), .A2(n3982), .B1(n3855), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3523) );
  NAND2_X1 U4565 ( .A1(n3546), .A2(EAX_REG_3__SCAN_IN), .ZN(n3522) );
  OAI211_X1 U4566 ( .C1(n3528), .C2(n3018), .A(n3523), .B(n3522), .ZN(n3524)
         );
  INV_X1 U4567 ( .A(n4533), .ZN(n3525) );
  OAI211_X1 U4568 ( .C1(n4534), .C2(n4611), .A(n4535), .B(n3525), .ZN(n4537)
         );
  NAND2_X1 U4569 ( .A1(n6657), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3527)
         );
  NAND2_X1 U4570 ( .A1(n3546), .A2(EAX_REG_4__SCAN_IN), .ZN(n3526) );
  OAI211_X1 U4571 ( .C1(n3528), .C2(n4032), .A(n3527), .B(n3526), .ZN(n3530)
         );
  OAI21_X1 U4572 ( .B1(n3529), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3547), 
        .ZN(n6363) );
  MUX2_X1 U4573 ( .A(n3530), .B(n6363), .S(n3982), .Z(n3531) );
  NOR2_X2 U4574 ( .A1(n4537), .A2(n4601), .ZN(n4546) );
  INV_X1 U4575 ( .A(n3532), .ZN(n3533) );
  AOI22_X1 U4576 ( .A1(n3825), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4577 ( .A1(n3963), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4578 ( .A1(n3939), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4579 ( .A1(n3921), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3536) );
  NAND4_X1 U4580 ( .A1(n3539), .A2(n3538), .A3(n3537), .A4(n3536), .ZN(n3545)
         );
  AOI22_X1 U4581 ( .A1(n3957), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4582 ( .A1(n3958), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4583 ( .A1(n3944), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4584 ( .A1(n3900), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3540) );
  NAND4_X1 U4585 ( .A1(n3543), .A2(n3542), .A3(n3541), .A4(n3540), .ZN(n3544)
         );
  AOI22_X1 U4586 ( .A1(n4039), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4013), 
        .B2(n4300), .ZN(n3554) );
  NAND2_X1 U4587 ( .A1(n3553), .A2(n3554), .ZN(n4288) );
  INV_X1 U4588 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4994) );
  INV_X1 U4589 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5498) );
  OR2_X1 U4590 ( .A1(n3548), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3549) );
  NAND2_X1 U4591 ( .A1(n3572), .A2(n3549), .ZN(n6353) );
  AOI22_X1 U4592 ( .A1(n6353), .A2(n3982), .B1(n3855), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3550) );
  OAI21_X1 U4593 ( .B1(n3674), .B2(n4994), .A(n3550), .ZN(n3551) );
  AOI21_X1 U4594 ( .B1(n4288), .B2(n3685), .A(n3551), .ZN(n4631) );
  NAND2_X1 U4595 ( .A1(n4039), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3556) );
  NAND2_X1 U4596 ( .A1(n4013), .A2(n4315), .ZN(n3555) );
  NAND2_X1 U4597 ( .A1(n3556), .A2(n3555), .ZN(n3557) );
  XNOR2_X1 U4598 ( .A(n4287), .B(n3557), .ZN(n4298) );
  INV_X1 U4599 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4995) );
  INV_X1 U4600 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3558) );
  XNOR2_X1 U4601 ( .A(n3572), .B(n3558), .ZN(n5473) );
  NAND2_X1 U4602 ( .A1(n5473), .A2(n3982), .ZN(n3560) );
  NAND2_X1 U4603 ( .A1(n3855), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3559)
         );
  OAI211_X1 U4604 ( .C1(n3674), .C2(n4995), .A(n3560), .B(n3559), .ZN(n3561)
         );
  AOI21_X1 U4605 ( .B1(n4298), .B2(n3685), .A(n3561), .ZN(n4968) );
  AOI22_X1 U4606 ( .A1(n3939), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4607 ( .A1(n3957), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4608 ( .A1(n3958), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3563) );
  AOI22_X1 U4609 ( .A1(n3920), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3562) );
  NAND4_X1 U4610 ( .A1(n3565), .A2(n3564), .A3(n3563), .A4(n3562), .ZN(n3571)
         );
  AOI22_X1 U4611 ( .A1(n3825), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3569) );
  AOI22_X1 U4612 ( .A1(n3965), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3568) );
  AOI22_X1 U4613 ( .A1(n3900), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3567) );
  AOI22_X1 U4614 ( .A1(n3963), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3566) );
  NAND4_X1 U4615 ( .A1(n3569), .A2(n3568), .A3(n3567), .A4(n3566), .ZN(n3570)
         );
  OAI21_X1 U4616 ( .B1(n3571), .B2(n3570), .A(n3685), .ZN(n3576) );
  NAND2_X1 U4617 ( .A1(n3546), .A2(EAX_REG_8__SCAN_IN), .ZN(n3575) );
  XNOR2_X1 U4618 ( .A(n3577), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6281) );
  NAND2_X1 U4619 ( .A1(n6281), .A2(n3982), .ZN(n3574) );
  NAND2_X1 U4620 ( .A1(n3855), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3573)
         );
  NAND4_X1 U4621 ( .A1(n3576), .A2(n3575), .A3(n3574), .A4(n3573), .ZN(n4979)
         );
  XNOR2_X1 U4622 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .B(n3592), .ZN(n6265) );
  AOI22_X1 U4623 ( .A1(n3825), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3581) );
  AOI22_X1 U4624 ( .A1(n3939), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4625 ( .A1(n3957), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3958), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4626 ( .A1(n3920), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3578) );
  NAND4_X1 U4627 ( .A1(n3581), .A2(n3580), .A3(n3579), .A4(n3578), .ZN(n3587)
         );
  AOI22_X1 U4628 ( .A1(n3900), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3585) );
  AOI22_X1 U4629 ( .A1(n3963), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3584) );
  AOI22_X1 U4630 ( .A1(n3966), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3583) );
  AOI22_X1 U4631 ( .A1(n3944), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3582) );
  NAND4_X1 U4632 ( .A1(n3585), .A2(n3584), .A3(n3583), .A4(n3582), .ZN(n3586)
         );
  OR2_X1 U4633 ( .A1(n3587), .A2(n3586), .ZN(n3588) );
  AOI22_X1 U4634 ( .A1(n3685), .A2(n3588), .B1(n3855), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3590) );
  NAND2_X1 U4635 ( .A1(n3546), .A2(EAX_REG_9__SCAN_IN), .ZN(n3589) );
  OAI211_X1 U4636 ( .C1(n6265), .C2(n3797), .A(n3590), .B(n3589), .ZN(n4998)
         );
  INV_X1 U4637 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3591) );
  NOR2_X1 U4638 ( .A1(n3592), .A2(n3591), .ZN(n3618) );
  XNOR2_X1 U4639 ( .A(n3618), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5807)
         );
  AOI22_X1 U4640 ( .A1(n3825), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3243), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3596) );
  AOI22_X1 U4641 ( .A1(n3958), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4642 ( .A1(n3957), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4643 ( .A1(n3900), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3593) );
  NAND4_X1 U4644 ( .A1(n3596), .A2(n3595), .A3(n3594), .A4(n3593), .ZN(n3602)
         );
  AOI22_X1 U4645 ( .A1(n3939), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3600) );
  AOI22_X1 U4646 ( .A1(n3965), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4647 ( .A1(n2965), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4648 ( .A1(n3920), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3597) );
  NAND4_X1 U4649 ( .A1(n3600), .A2(n3599), .A3(n3598), .A4(n3597), .ZN(n3601)
         );
  OAI21_X1 U4650 ( .B1(n3602), .B2(n3601), .A(n3685), .ZN(n3605) );
  NAND2_X1 U4651 ( .A1(n3977), .A2(EAX_REG_10__SCAN_IN), .ZN(n3604) );
  NAND2_X1 U4652 ( .A1(n3855), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3603)
         );
  NAND3_X1 U4653 ( .A1(n3605), .A2(n3604), .A3(n3603), .ZN(n3606) );
  AOI21_X1 U4654 ( .B1(n5807), .B2(n3982), .A(n3606), .ZN(n5157) );
  AOI22_X1 U4655 ( .A1(n3825), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3611) );
  AOI22_X1 U4656 ( .A1(n3966), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3610) );
  AOI22_X1 U4657 ( .A1(n3944), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3609) );
  AOI22_X1 U4658 ( .A1(n3900), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3608) );
  NAND4_X1 U4659 ( .A1(n3611), .A2(n3610), .A3(n3609), .A4(n3608), .ZN(n3617)
         );
  AOI22_X1 U4660 ( .A1(n3920), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4661 ( .A1(n3939), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3614) );
  AOI22_X1 U4662 ( .A1(n3957), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3958), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3613) );
  AOI22_X1 U4663 ( .A1(n3963), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3612) );
  NAND4_X1 U4664 ( .A1(n3615), .A2(n3614), .A3(n3613), .A4(n3612), .ZN(n3616)
         );
  OAI21_X1 U4665 ( .B1(n3617), .B2(n3616), .A(n3685), .ZN(n3622) );
  NAND2_X1 U4666 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n3619), .ZN(n3636)
         );
  OAI21_X1 U4667 ( .B1(PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n3619), .A(n3636), 
        .ZN(n6340) );
  AOI22_X1 U4668 ( .A1(n3982), .A2(n6340), .B1(n3855), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3621) );
  NAND2_X1 U4669 ( .A1(n3546), .A2(EAX_REG_11__SCAN_IN), .ZN(n3620) );
  XNOR2_X1 U4670 ( .A(n3636), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5801)
         );
  AOI22_X1 U4671 ( .A1(n3977), .A2(EAX_REG_12__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6657), .ZN(n3623) );
  MUX2_X1 U4672 ( .A(n5801), .B(n3623), .S(n3797), .Z(n3635) );
  AOI22_X1 U4673 ( .A1(n3965), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3627) );
  AOI22_X1 U4674 ( .A1(n3957), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4675 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3966), .B1(n3864), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4676 ( .A1(n3963), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3624) );
  NAND4_X1 U4677 ( .A1(n3627), .A2(n3626), .A3(n3625), .A4(n3624), .ZN(n3633)
         );
  AOI22_X1 U4678 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n3939), .B1(n3728), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4679 ( .A1(n3825), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4680 ( .A1(n3956), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4681 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n3863), .B1(n3964), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3628) );
  NAND4_X1 U4682 ( .A1(n3631), .A2(n3630), .A3(n3629), .A4(n3628), .ZN(n3632)
         );
  OAI21_X1 U4683 ( .B1(n3633), .B2(n3632), .A(n3685), .ZN(n3634) );
  NAND2_X1 U4684 ( .A1(n3635), .A2(n3634), .ZN(n5164) );
  NAND2_X1 U4685 ( .A1(n3546), .A2(EAX_REG_13__SCAN_IN), .ZN(n3643) );
  INV_X1 U4686 ( .A(n3636), .ZN(n3637) );
  NAND2_X1 U4687 ( .A1(n3638), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3675)
         );
  INV_X1 U4688 ( .A(n3638), .ZN(n3640) );
  INV_X1 U4689 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3639) );
  NAND2_X1 U4690 ( .A1(n3640), .A2(n3639), .ZN(n3641) );
  NAND2_X1 U4691 ( .A1(n3675), .A2(n3641), .ZN(n5789) );
  AOI22_X1 U4692 ( .A1(n5789), .A2(n3982), .B1(PHYADDRPOINTER_REG_13__SCAN_IN), 
        .B2(n3855), .ZN(n3642) );
  OR2_X2 U4693 ( .A1(n3645), .A2(n3644), .ZN(n3659) );
  NAND2_X1 U4694 ( .A1(n3645), .A2(n3644), .ZN(n3646) );
  AOI22_X1 U4695 ( .A1(n3825), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4696 ( .A1(n3958), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4697 ( .A1(n3965), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4698 ( .A1(n3956), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3647) );
  NAND4_X1 U4699 ( .A1(n3650), .A2(n3649), .A3(n3648), .A4(n3647), .ZN(n3656)
         );
  AOI22_X1 U4700 ( .A1(n3939), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3654) );
  AOI22_X1 U4701 ( .A1(n3957), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4702 ( .A1(n3963), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4703 ( .A1(n3900), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3651) );
  NAND4_X1 U4704 ( .A1(n3654), .A2(n3653), .A3(n3652), .A4(n3651), .ZN(n3655)
         );
  NAND2_X1 U4705 ( .A1(n3685), .A2(n3657), .ZN(n5433) );
  INV_X1 U4706 ( .A(EAX_REG_14__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4707 ( .A1(n3825), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3663) );
  AOI22_X1 U4708 ( .A1(n3965), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3662) );
  AOI22_X1 U4709 ( .A1(n3957), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3661) );
  AOI22_X1 U4710 ( .A1(n3920), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3660) );
  NAND4_X1 U4711 ( .A1(n3663), .A2(n3662), .A3(n3661), .A4(n3660), .ZN(n3669)
         );
  AOI22_X1 U4712 ( .A1(n3939), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3728), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4713 ( .A1(n3958), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3666) );
  AOI22_X1 U4714 ( .A1(n3963), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3665) );
  AOI22_X1 U4715 ( .A1(n3864), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3664) );
  NAND4_X1 U4716 ( .A1(n3667), .A2(n3666), .A3(n3665), .A4(n3664), .ZN(n3668)
         );
  OAI21_X1 U4717 ( .B1(n3669), .B2(n3668), .A(n3685), .ZN(n3672) );
  INV_X1 U4718 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3670) );
  XNOR2_X1 U4719 ( .A(n3675), .B(n3670), .ZN(n5782) );
  AOI22_X1 U4720 ( .A1(n5782), .A2(n3982), .B1(PHYADDRPOINTER_REG_14__SCAN_IN), 
        .B2(n3855), .ZN(n3671) );
  OAI211_X1 U4721 ( .C1(n3674), .C2(n3673), .A(n3672), .B(n3671), .ZN(n5419)
         );
  INV_X1 U4722 ( .A(n3675), .ZN(n3692) );
  NAND2_X1 U4723 ( .A1(n3692), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3676)
         );
  XNOR2_X1 U4724 ( .A(n3676), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5405)
         );
  AOI22_X1 U4725 ( .A1(n3546), .A2(EAX_REG_15__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n3855), .ZN(n3689) );
  AOI22_X1 U4726 ( .A1(n3957), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4727 ( .A1(n3958), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3679) );
  AOI22_X1 U4728 ( .A1(n2965), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3678) );
  AOI22_X1 U4729 ( .A1(n3900), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3677) );
  NAND4_X1 U4730 ( .A1(n3680), .A2(n3679), .A3(n3678), .A4(n3677), .ZN(n3687)
         );
  AOI22_X1 U4731 ( .A1(n3963), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3684) );
  AOI22_X1 U4732 ( .A1(n3939), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3683) );
  AOI22_X1 U4733 ( .A1(n3944), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4734 ( .A1(n3825), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3681) );
  NAND4_X1 U4735 ( .A1(n3684), .A2(n3683), .A3(n3682), .A4(n3681), .ZN(n3686)
         );
  OAI21_X1 U4736 ( .B1(n3687), .B2(n3686), .A(n3685), .ZN(n3688) );
  OAI211_X1 U4737 ( .C1(n5405), .C2(n3797), .A(n3689), .B(n3688), .ZN(n3690)
         );
  INV_X1 U4738 ( .A(n3690), .ZN(n5404) );
  XNOR2_X1 U4739 ( .A(n3721), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5769)
         );
  AOI22_X1 U4740 ( .A1(n3900), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3696) );
  AOI22_X1 U4741 ( .A1(n3966), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3695) );
  AOI22_X1 U4742 ( .A1(n3957), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3694) );
  AOI22_X1 U4743 ( .A1(n3921), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3693) );
  NAND4_X1 U4744 ( .A1(n3696), .A2(n3695), .A3(n3694), .A4(n3693), .ZN(n3704)
         );
  AOI22_X1 U4745 ( .A1(n3825), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4746 ( .A1(n3963), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4747 ( .A1(n3939), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3698) );
  AOI22_X1 U4748 ( .A1(n3944), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3958), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3697) );
  NAND4_X1 U4749 ( .A1(n3700), .A2(n3699), .A3(n3698), .A4(n3697), .ZN(n3703)
         );
  NAND3_X1 U4750 ( .A1(n3701), .A2(n3334), .A3(n4662), .ZN(n3702) );
  OAI21_X1 U4751 ( .B1(n3704), .B2(n3703), .A(n3953), .ZN(n3706) );
  AOI22_X1 U4752 ( .A1(n3977), .A2(EAX_REG_16__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n3855), .ZN(n3705) );
  OAI211_X1 U4753 ( .C1(n5769), .C2(n3797), .A(n3706), .B(n3705), .ZN(n5391)
         );
  AOI22_X1 U4754 ( .A1(n3825), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3710) );
  AOI22_X1 U4755 ( .A1(n3957), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4756 ( .A1(n3900), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3708) );
  AOI22_X1 U4757 ( .A1(n3864), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3707) );
  NAND4_X1 U4758 ( .A1(n3710), .A2(n3709), .A3(n3708), .A4(n3707), .ZN(n3718)
         );
  AOI22_X1 U4759 ( .A1(n3939), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4760 ( .A1(n3963), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3715) );
  NAND2_X1 U4761 ( .A1(n3958), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3712) );
  NAND2_X1 U4762 ( .A1(n3921), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3711) );
  AND3_X1 U4763 ( .A1(n3712), .A2(n3797), .A3(n3711), .ZN(n3714) );
  AOI22_X1 U4764 ( .A1(n3944), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3713) );
  NAND4_X1 U4765 ( .A1(n3716), .A2(n3715), .A3(n3714), .A4(n3713), .ZN(n3717)
         );
  INV_X1 U4766 ( .A(n3953), .ZN(n3979) );
  NAND2_X1 U4767 ( .A1(n3979), .A2(n3797), .ZN(n3776) );
  OAI21_X1 U4768 ( .B1(n3718), .B2(n3717), .A(n3776), .ZN(n3720) );
  AOI22_X1 U4769 ( .A1(n3977), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6657), .ZN(n3719) );
  NAND2_X1 U4770 ( .A1(n3720), .A2(n3719), .ZN(n3723) );
  XNOR2_X1 U4771 ( .A(n3737), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5762)
         );
  NAND2_X1 U4772 ( .A1(n5762), .A2(n3982), .ZN(n3722) );
  NAND2_X1 U4773 ( .A1(n3723), .A2(n3722), .ZN(n5378) );
  INV_X1 U4774 ( .A(n5364), .ZN(n3741) );
  AOI22_X1 U4775 ( .A1(n3825), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3727) );
  AOI22_X1 U4776 ( .A1(n3863), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3726) );
  AOI22_X1 U4777 ( .A1(n3920), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3725) );
  AOI22_X1 U4778 ( .A1(n3956), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3724) );
  NAND4_X1 U4779 ( .A1(n3727), .A2(n3726), .A3(n3725), .A4(n3724), .ZN(n3734)
         );
  AOI22_X1 U4780 ( .A1(n3939), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3728), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3732) );
  AOI22_X1 U4781 ( .A1(n3957), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4782 ( .A1(n3963), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3730) );
  AOI22_X1 U4783 ( .A1(n3944), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3729) );
  NAND4_X1 U4784 ( .A1(n3732), .A2(n3731), .A3(n3730), .A4(n3729), .ZN(n3733)
         );
  OAI21_X1 U4785 ( .B1(n3734), .B2(n3733), .A(n3953), .ZN(n3736) );
  AOI22_X1 U4786 ( .A1(n3977), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6657), .ZN(n3735) );
  AND2_X1 U4787 ( .A1(n3736), .A2(n3735), .ZN(n3739) );
  AOI21_X1 U4788 ( .B1(n5750), .B2(n3738), .A(n3771), .ZN(n5748) );
  MUX2_X1 U4789 ( .A(n3739), .B(n5748), .S(n3982), .Z(n5366) );
  AOI22_X1 U4790 ( .A1(n3963), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3745) );
  AOI22_X1 U4791 ( .A1(n2965), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3744) );
  AOI22_X1 U4792 ( .A1(n3863), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4793 ( .A1(n3944), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3742) );
  NAND4_X1 U4794 ( .A1(n3745), .A2(n3744), .A3(n3743), .A4(n3742), .ZN(n3753)
         );
  AOI22_X1 U4795 ( .A1(n3825), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3939), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4796 ( .A1(n3957), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3750) );
  NAND2_X1 U4797 ( .A1(n3268), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3747)
         );
  NAND2_X1 U4798 ( .A1(n3921), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3746) );
  AND3_X1 U4799 ( .A1(n3747), .A2(n3797), .A3(n3746), .ZN(n3749) );
  AOI22_X1 U4800 ( .A1(n3900), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3748) );
  NAND4_X1 U4801 ( .A1(n3751), .A2(n3750), .A3(n3749), .A4(n3748), .ZN(n3752)
         );
  OAI21_X1 U4802 ( .B1(n3753), .B2(n3752), .A(n3776), .ZN(n3755) );
  AOI22_X1 U4803 ( .A1(n3977), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6657), .ZN(n3754) );
  NAND2_X1 U4804 ( .A1(n3755), .A2(n3754), .ZN(n3758) );
  INV_X1 U4805 ( .A(n3771), .ZN(n3756) );
  XNOR2_X1 U4806 ( .A(n3756), .B(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5744)
         );
  NAND2_X1 U4807 ( .A1(n5744), .A2(n3982), .ZN(n3757) );
  NAND2_X1 U4808 ( .A1(n3758), .A2(n3757), .ZN(n5348) );
  AOI22_X1 U4809 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3958), .B1(n3268), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4810 ( .A1(n3963), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4811 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3900), .B1(n3964), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3760) );
  AOI22_X1 U4812 ( .A1(n3825), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3759) );
  NAND4_X1 U4813 ( .A1(n3762), .A2(n3761), .A3(n3760), .A4(n3759), .ZN(n3768)
         );
  AOI22_X1 U4814 ( .A1(n2965), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4815 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n3957), .B1(n3965), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4816 ( .A1(n3939), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3764) );
  AOI22_X1 U4817 ( .A1(n3944), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3763) );
  NAND4_X1 U4818 ( .A1(n3766), .A2(n3765), .A3(n3764), .A4(n3763), .ZN(n3767)
         );
  OAI21_X1 U4819 ( .B1(n3768), .B2(n3767), .A(n3953), .ZN(n3770) );
  AOI22_X1 U4820 ( .A1(n3977), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6657), .ZN(n3769) );
  NAND2_X1 U4821 ( .A1(n3770), .A2(n3769), .ZN(n3775) );
  INV_X1 U4822 ( .A(n3772), .ZN(n3773) );
  INV_X1 U4823 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5340) );
  NAND2_X1 U4824 ( .A1(n3773), .A2(n5340), .ZN(n3774) );
  NAND2_X1 U4825 ( .A1(n3798), .A2(n3774), .ZN(n5734) );
  MUX2_X1 U4826 ( .A(n3775), .B(n5734), .S(n3982), .Z(n5335) );
  XOR2_X1 U4827 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n3798), .Z(n5726) );
  INV_X1 U4828 ( .A(n3776), .ZN(n3795) );
  AOI22_X1 U4829 ( .A1(n3963), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3958), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4830 ( .A1(n3956), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4831 ( .A1(n3825), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4832 ( .A1(n3964), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3777) );
  NAND4_X1 U4833 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3777), .ZN(n3792)
         );
  INV_X1 U4834 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4877) );
  AOI22_X1 U4835 ( .A1(n3965), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3782) );
  AOI21_X1 U4836 ( .B1(n2965), .B2(INSTQUEUE_REG_0__5__SCAN_IN), .A(n3982), 
        .ZN(n3781) );
  OAI211_X1 U4837 ( .C1(n3396), .C2(n4877), .A(n3782), .B(n3781), .ZN(n3791)
         );
  INV_X1 U4838 ( .A(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3784) );
  INV_X1 U4839 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3783) );
  OAI22_X1 U4840 ( .A1(n3785), .A2(n3784), .B1(n5181), .B2(n3783), .ZN(n3790)
         );
  INV_X1 U4841 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3787) );
  INV_X1 U4842 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3786) );
  OAI22_X1 U4843 ( .A1(n3788), .A2(n3787), .B1(n3415), .B2(n3786), .ZN(n3789)
         );
  NOR4_X1 U4844 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(n3794)
         );
  AOI22_X1 U4845 ( .A1(n3977), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6657), .ZN(n3793) );
  OAI21_X1 U4846 ( .B1(n3795), .B2(n3794), .A(n3793), .ZN(n3796) );
  OAI21_X1 U4847 ( .B1(n5726), .B2(n3797), .A(n3796), .ZN(n5323) );
  NAND2_X1 U4848 ( .A1(n3799), .A2(n5716), .ZN(n3800) );
  AND2_X1 U4849 ( .A1(n3853), .A2(n3800), .ZN(n5720) );
  OAI21_X1 U4850 ( .B1(PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6469), .A(n6657), 
        .ZN(n3801) );
  INV_X1 U4851 ( .A(n3801), .ZN(n3802) );
  AOI21_X1 U4852 ( .B1(n3546), .B2(EAX_REG_22__SCAN_IN), .A(n3802), .ZN(n3814)
         );
  AOI22_X1 U4853 ( .A1(n3825), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3806) );
  AOI22_X1 U4854 ( .A1(n3939), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3805) );
  AOI22_X1 U4855 ( .A1(n3920), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3804) );
  AOI22_X1 U4856 ( .A1(n3963), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3803) );
  NAND4_X1 U4857 ( .A1(n3806), .A2(n3805), .A3(n3804), .A4(n3803), .ZN(n3812)
         );
  AOI22_X1 U4858 ( .A1(n3958), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3810) );
  AOI22_X1 U4859 ( .A1(n3900), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4860 ( .A1(n3944), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4861 ( .A1(n3957), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3807) );
  NAND4_X1 U4862 ( .A1(n3810), .A2(n3809), .A3(n3808), .A4(n3807), .ZN(n3811)
         );
  OAI21_X1 U4863 ( .B1(n3812), .B2(n3811), .A(n3953), .ZN(n3813) );
  AOI22_X1 U4864 ( .A1(n5720), .A2(n3982), .B1(n3814), .B2(n3813), .ZN(n5310)
         );
  AOI22_X1 U4865 ( .A1(n3939), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3957), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4866 ( .A1(n3963), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4867 ( .A1(n3863), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4868 ( .A1(n3825), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3815) );
  NAND4_X1 U4869 ( .A1(n3818), .A2(n3817), .A3(n3816), .A4(n3815), .ZN(n3824)
         );
  AOI22_X1 U4870 ( .A1(n3900), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4871 ( .A1(n3944), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4872 ( .A1(n2965), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4873 ( .A1(n3965), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3819) );
  NAND4_X1 U4874 ( .A1(n3822), .A2(n3821), .A3(n3820), .A4(n3819), .ZN(n3823)
         );
  NOR2_X1 U4875 ( .A1(n3824), .A2(n3823), .ZN(n3840) );
  AOI22_X1 U4876 ( .A1(n3939), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4877 ( .A1(n3963), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4878 ( .A1(n3944), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4879 ( .A1(n3825), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3826) );
  NAND4_X1 U4880 ( .A1(n3829), .A2(n3828), .A3(n3827), .A4(n3826), .ZN(n3835)
         );
  AOI22_X1 U4881 ( .A1(n3900), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4882 ( .A1(n3958), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4883 ( .A1(n2965), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4884 ( .A1(n3957), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3830) );
  NAND4_X1 U4885 ( .A1(n3833), .A2(n3832), .A3(n3831), .A4(n3830), .ZN(n3834)
         );
  NOR2_X1 U4886 ( .A1(n3835), .A2(n3834), .ZN(n3841) );
  XOR2_X1 U4887 ( .A(n3840), .B(n3841), .Z(n3838) );
  INV_X1 U4888 ( .A(EAX_REG_23__SCAN_IN), .ZN(n3836) );
  INV_X1 U4889 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5708) );
  OAI22_X1 U4890 ( .A1(n3674), .A2(n3836), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5708), .ZN(n3837) );
  AOI21_X1 U4891 ( .B1(n3953), .B2(n3838), .A(n3837), .ZN(n3839) );
  XNOR2_X1 U4892 ( .A(n3853), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5710)
         );
  MUX2_X1 U4893 ( .A(n3839), .B(n5710), .S(n3982), .Z(n5298) );
  OR2_X1 U4894 ( .A1(n3841), .A2(n3840), .ZN(n3872) );
  AOI22_X1 U4895 ( .A1(n3957), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4896 ( .A1(n3965), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3958), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4897 ( .A1(n2965), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3843) );
  INV_X1 U4898 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n6752) );
  AOI22_X1 U4899 ( .A1(n3926), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3842) );
  NAND4_X1 U4900 ( .A1(n3845), .A2(n3844), .A3(n3843), .A4(n3842), .ZN(n3851)
         );
  AOI22_X1 U4901 ( .A1(n3825), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3243), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4902 ( .A1(n3920), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4903 ( .A1(n3939), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4904 ( .A1(n3900), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3846) );
  NAND4_X1 U4905 ( .A1(n3849), .A2(n3848), .A3(n3847), .A4(n3846), .ZN(n3850)
         );
  NOR2_X1 U4906 ( .A1(n3851), .A2(n3850), .ZN(n3871) );
  XNOR2_X1 U4907 ( .A(n3872), .B(n3871), .ZN(n3858) );
  INV_X1 U4908 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5289) );
  OAI21_X1 U4909 ( .B1(n3853), .B2(n5708), .A(n5289), .ZN(n3854) );
  NAND2_X1 U4910 ( .A1(n3877), .A2(n3854), .ZN(n5698) );
  NAND2_X1 U4911 ( .A1(n5698), .A2(n3982), .ZN(n3857) );
  AOI22_X1 U4912 ( .A1(n3977), .A2(EAX_REG_24__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n3855), .ZN(n3856) );
  OAI211_X1 U4913 ( .C1(n3858), .C2(n3979), .A(n3857), .B(n3856), .ZN(n5287)
         );
  AOI22_X1 U4914 ( .A1(n3825), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4915 ( .A1(n3963), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4916 ( .A1(n3939), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4917 ( .A1(n3921), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3859) );
  NAND4_X1 U4918 ( .A1(n3862), .A2(n3861), .A3(n3860), .A4(n3859), .ZN(n3870)
         );
  AOI22_X1 U4919 ( .A1(n3957), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4920 ( .A1(n3863), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4921 ( .A1(n3944), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4922 ( .A1(n3900), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3865) );
  NAND4_X1 U4923 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(n3869)
         );
  NOR2_X1 U4924 ( .A1(n3870), .A2(n3869), .ZN(n3881) );
  OR2_X1 U4925 ( .A1(n3872), .A2(n3871), .ZN(n3880) );
  XOR2_X1 U4926 ( .A(n3881), .B(n3880), .Z(n3875) );
  INV_X1 U4927 ( .A(EAX_REG_25__SCAN_IN), .ZN(n3873) );
  OAI22_X1 U4928 ( .A1(n3674), .A2(n3873), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6754), .ZN(n3874) );
  AOI21_X1 U4929 ( .B1(n3875), .B2(n3953), .A(n3874), .ZN(n3879) );
  NAND2_X1 U4930 ( .A1(n3877), .A2(n6754), .ZN(n3878) );
  MUX2_X1 U4931 ( .A(n3879), .B(n5688), .S(n3982), .Z(n5271) );
  NOR2_X1 U4932 ( .A1(n3881), .A2(n3880), .ZN(n3899) );
  AOI22_X1 U4933 ( .A1(n3825), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4934 ( .A1(n3963), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4935 ( .A1(n3939), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4936 ( .A1(n3921), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3882), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3883) );
  NAND4_X1 U4937 ( .A1(n3886), .A2(n3885), .A3(n3884), .A4(n3883), .ZN(n3892)
         );
  AOI22_X1 U4938 ( .A1(n3957), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4939 ( .A1(n3958), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3268), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4940 ( .A1(n3926), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3864), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4941 ( .A1(n3900), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3887) );
  NAND4_X1 U4942 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n3891)
         );
  XNOR2_X1 U4943 ( .A(n3899), .B(n3898), .ZN(n3894) );
  AOI22_X1 U4944 ( .A1(n3977), .A2(EAX_REG_26__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n6657), .ZN(n3893) );
  OAI21_X1 U4945 ( .B1(n3894), .B2(n3979), .A(n3893), .ZN(n3897) );
  NAND2_X1 U4946 ( .A1(n3895), .A2(n5262), .ZN(n3896) );
  NAND2_X1 U4947 ( .A1(n2996), .A2(n3896), .ZN(n5680) );
  MUX2_X1 U4948 ( .A(n3897), .B(n5680), .S(n3982), .Z(n5261) );
  NAND2_X1 U4949 ( .A1(n3899), .A2(n3898), .ZN(n3918) );
  AOI22_X1 U4950 ( .A1(n3243), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3939), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4951 ( .A1(n3825), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n2965), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4952 ( .A1(n3921), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4953 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n3900), .B1(n3964), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3901) );
  NAND4_X1 U4954 ( .A1(n3904), .A2(n3903), .A3(n3902), .A4(n3901), .ZN(n3910)
         );
  AOI22_X1 U4955 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3956), .B1(n3920), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4956 ( .A1(n3957), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4957 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3966), .B1(n3958), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4958 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3944), .B1(n3381), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3905) );
  NAND4_X1 U4959 ( .A1(n3908), .A2(n3907), .A3(n3906), .A4(n3905), .ZN(n3909)
         );
  NOR2_X1 U4960 ( .A1(n3910), .A2(n3909), .ZN(n3919) );
  XOR2_X1 U4961 ( .A(n3918), .B(n3919), .Z(n3913) );
  INV_X1 U4962 ( .A(EAX_REG_27__SCAN_IN), .ZN(n3911) );
  OAI22_X1 U4963 ( .A1(n3674), .A2(n3911), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5671), .ZN(n3912) );
  AOI21_X1 U4964 ( .B1(n3913), .B2(n3953), .A(n3912), .ZN(n3915) );
  INV_X1 U4965 ( .A(n2996), .ZN(n3914) );
  XOR2_X1 U4966 ( .A(n3914), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .Z(n5669) );
  MUX2_X1 U4967 ( .A(n3915), .B(n5669), .S(n3982), .Z(n5246) );
  NOR2_X1 U4968 ( .A1(n3919), .A2(n3918), .ZN(n3938) );
  AOI22_X1 U4969 ( .A1(n3825), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4970 ( .A1(n3243), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3920), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4971 ( .A1(n3939), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4972 ( .A1(n3921), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3922) );
  NAND4_X1 U4973 ( .A1(n3925), .A2(n3924), .A3(n3923), .A4(n3922), .ZN(n3932)
         );
  AOI22_X1 U4974 ( .A1(n3957), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3965), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3930) );
  AOI22_X1 U4975 ( .A1(n3958), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3966), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4976 ( .A1(n3926), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3381), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4977 ( .A1(n3900), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3927) );
  NAND4_X1 U4978 ( .A1(n3930), .A2(n3929), .A3(n3928), .A4(n3927), .ZN(n3931)
         );
  OR2_X1 U4979 ( .A1(n3932), .A2(n3931), .ZN(n3937) );
  XOR2_X1 U4980 ( .A(n3938), .B(n3937), .Z(n3935) );
  INV_X1 U4981 ( .A(EAX_REG_28__SCAN_IN), .ZN(n3933) );
  OAI22_X1 U4982 ( .A1(n3674), .A2(n3933), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3074), .ZN(n3934) );
  AOI21_X1 U4983 ( .B1(n3935), .B2(n3953), .A(n3934), .ZN(n3936) );
  AOI21_X1 U4984 ( .B1(n3074), .B2(n2997), .A(n3981), .ZN(n5662) );
  MUX2_X1 U4985 ( .A(n3936), .B(n5662), .S(n3982), .Z(n4190) );
  NAND2_X1 U4986 ( .A1(n3938), .A2(n3937), .ZN(n3973) );
  AOI22_X1 U4987 ( .A1(n3825), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3288), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4988 ( .A1(n3939), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4989 ( .A1(n3957), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3958), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4990 ( .A1(n3920), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3940) );
  NAND4_X1 U4991 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(n3950)
         );
  AOI22_X1 U4992 ( .A1(n3965), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3944), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4993 ( .A1(n3243), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3921), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4994 ( .A1(n3966), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3381), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4995 ( .A1(n3900), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3945) );
  NAND4_X1 U4996 ( .A1(n3948), .A2(n3947), .A3(n3946), .A4(n3945), .ZN(n3949)
         );
  NOR2_X1 U4997 ( .A1(n3950), .A2(n3949), .ZN(n3974) );
  XOR2_X1 U4998 ( .A(n3973), .B(n3974), .Z(n3954) );
  INV_X1 U4999 ( .A(EAX_REG_29__SCAN_IN), .ZN(n3951) );
  INV_X1 U5000 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5654) );
  OAI22_X1 U5001 ( .A1(n3674), .A2(n3951), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5654), .ZN(n3952) );
  AOI21_X1 U5002 ( .B1(n3954), .B2(n3953), .A(n3952), .ZN(n3955) );
  XOR2_X1 U5003 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .B(n3981), .Z(n5652) );
  MUX2_X1 U5004 ( .A(n3955), .B(n5652), .S(n3982), .Z(n5221) );
  AOI22_X1 U5005 ( .A1(n3920), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3956), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U5006 ( .A1(n3957), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3728), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U5007 ( .A1(n3944), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3958), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U5008 ( .A1(n3825), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3293), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3959) );
  NAND4_X1 U5009 ( .A1(n3962), .A2(n3961), .A3(n3960), .A4(n3959), .ZN(n3972)
         );
  AOI22_X1 U5010 ( .A1(n3963), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3939), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3970) );
  AOI22_X1 U5011 ( .A1(n3965), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3964), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3969) );
  AOI22_X1 U5012 ( .A1(n3966), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3381), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U5013 ( .A1(n2965), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3967) );
  NAND4_X1 U5014 ( .A1(n3970), .A2(n3969), .A3(n3968), .A4(n3967), .ZN(n3971)
         );
  NOR2_X1 U5015 ( .A1(n3972), .A2(n3971), .ZN(n3976) );
  NOR2_X1 U5016 ( .A1(n3974), .A2(n3973), .ZN(n3975) );
  XOR2_X1 U5017 ( .A(n3976), .B(n3975), .Z(n3980) );
  AOI22_X1 U5018 ( .A1(n3977), .A2(EAX_REG_30__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6657), .ZN(n3978) );
  OAI21_X1 U5019 ( .B1(n3980), .B2(n3979), .A(n3978), .ZN(n3983) );
  XNOR2_X1 U5020 ( .A(n4201), .B(n4228), .ZN(n4242) );
  MUX2_X1 U5021 ( .A(n3983), .B(n4242), .S(n3982), .Z(n5593) );
  INV_X1 U5022 ( .A(n5593), .ZN(n3984) );
  NOR2_X1 U5023 ( .A1(n3984), .A2(n5221), .ZN(n3985) );
  INV_X1 U5025 ( .A(n3994), .ZN(n3988) );
  XNOR2_X1 U5026 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3989) );
  INV_X1 U5027 ( .A(n3989), .ZN(n3987) );
  NAND2_X1 U5028 ( .A1(n3988), .A2(n3987), .ZN(n3990) );
  NAND2_X1 U5029 ( .A1(n3994), .A2(n3989), .ZN(n4009) );
  NAND2_X1 U5030 ( .A1(n3350), .A2(n3986), .ZN(n3991) );
  AND2_X1 U5031 ( .A1(n3991), .A2(n5491), .ZN(n4020) );
  AND2_X1 U5032 ( .A1(n3171), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3993)
         );
  NOR2_X1 U5033 ( .A1(n3994), .A2(n3993), .ZN(n3999) );
  NAND2_X1 U5034 ( .A1(n3992), .A2(n3999), .ZN(n3995) );
  NAND2_X1 U5035 ( .A1(n3995), .A2(n3346), .ZN(n3996) );
  OAI211_X1 U5036 ( .C1(n4043), .C2(n4054), .A(n4020), .B(n3996), .ZN(n4003)
         );
  INV_X1 U5037 ( .A(n4054), .ZN(n3998) );
  INV_X1 U5038 ( .A(n3999), .ZN(n4000) );
  OAI21_X1 U5039 ( .B1(n4037), .B2(n4000), .A(n4043), .ZN(n4001) );
  NAND3_X1 U5040 ( .A1(n4003), .A2(n4002), .A3(n4001), .ZN(n4007) );
  INV_X1 U5041 ( .A(n4004), .ZN(n4005) );
  NAND3_X1 U5042 ( .A1(n4005), .A2(STATE2_REG_0__SCAN_IN), .A3(n4054), .ZN(
        n4006) );
  NAND2_X1 U5043 ( .A1(n4007), .A2(n4006), .ZN(n4023) );
  NAND2_X1 U5044 ( .A1(n4748), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4008) );
  NAND2_X1 U5045 ( .A1(n4009), .A2(n4008), .ZN(n4015) );
  NAND2_X1 U5046 ( .A1(n4010), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4016) );
  NAND2_X1 U5047 ( .A1(n5174), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4011) );
  INV_X1 U5048 ( .A(n4014), .ZN(n4012) );
  XNOR2_X1 U5049 ( .A(n4015), .B(n4012), .ZN(n4053) );
  INV_X1 U5050 ( .A(n4039), .ZN(n4025) );
  NAND2_X1 U5051 ( .A1(n4013), .A2(n4053), .ZN(n4019) );
  OAI211_X1 U5052 ( .C1(n4053), .C2(n4025), .A(n4020), .B(n4019), .ZN(n4022)
         );
  NAND2_X1 U5053 ( .A1(n4015), .A2(n4014), .ZN(n4017) );
  NAND2_X1 U5054 ( .A1(n4017), .A2(n4016), .ZN(n4029) );
  XNOR2_X1 U5055 ( .A(n6681), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4018)
         );
  XNOR2_X1 U5056 ( .A(n4029), .B(n4018), .ZN(n4052) );
  OAI22_X1 U5057 ( .A1(n4020), .A2(n4019), .B1(n4052), .B2(n4312), .ZN(n4021)
         );
  AOI21_X1 U5058 ( .B1(n4023), .B2(n4022), .A(n4021), .ZN(n4027) );
  INV_X1 U5059 ( .A(n4052), .ZN(n4024) );
  NAND2_X1 U5060 ( .A1(n4029), .A2(n4028), .ZN(n4031) );
  NAND2_X1 U5061 ( .A1(n6681), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4030) );
  NAND2_X1 U5062 ( .A1(n4031), .A2(n4030), .ZN(n4034) );
  INV_X1 U5063 ( .A(n4057), .ZN(n4038) );
  AOI22_X1 U5064 ( .A1(n4039), .A2(n4038), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6747), .ZN(n4040) );
  INV_X1 U5065 ( .A(n4043), .ZN(n4045) );
  INV_X1 U5066 ( .A(n4056), .ZN(n4044) );
  AND2_X1 U5067 ( .A1(n3322), .A2(n6692), .ZN(n4048) );
  NAND2_X1 U5068 ( .A1(n4510), .A2(n4049), .ZN(n4050) );
  NAND2_X1 U5069 ( .A1(n3343), .A2(n4050), .ZN(n4429) );
  NOR2_X1 U5070 ( .A1(n4429), .A2(n5491), .ZN(n4696) );
  NAND2_X1 U5071 ( .A1(n4488), .A2(n4696), .ZN(n4060) );
  NAND3_X1 U5072 ( .A1(n4054), .A2(n4053), .A3(n4052), .ZN(n4055) );
  NAND2_X1 U5073 ( .A1(n4056), .A2(n4055), .ZN(n4058) );
  NOR2_X1 U5074 ( .A1(n4419), .A2(READY_N), .ZN(n4434) );
  NAND2_X1 U5075 ( .A1(n4723), .A2(n4434), .ZN(n4059) );
  NAND2_X1 U5076 ( .A1(n4060), .A2(n4059), .ZN(n4491) );
  NAND2_X1 U5077 ( .A1(n4491), .A2(n6654), .ZN(n4061) );
  INV_X1 U5078 ( .A(n4662), .ZN(n5591) );
  NAND2_X1 U5079 ( .A1(n4086), .A2(n3340), .ZN(n4066) );
  NAND2_X1 U5080 ( .A1(n3332), .A2(n4662), .ZN(n4628) );
  NAND2_X1 U5081 ( .A1(n5636), .A2(DATAI_30_), .ZN(n4068) );
  NOR2_X2 U5082 ( .A1(n4629), .A2(n3986), .ZN(n5635) );
  AOI22_X1 U5083 ( .A1(n5635), .A2(DATAI_14_), .B1(n5641), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n4067) );
  AND2_X1 U5084 ( .A1(n4068), .A2(n4067), .ZN(n4069) );
  OAI21_X1 U5085 ( .B1(n4200), .B2(n4987), .A(n4069), .ZN(U2861) );
  NAND2_X1 U5086 ( .A1(n4297), .A2(n3326), .ZN(n4415) );
  NAND2_X1 U5087 ( .A1(n3323), .A2(n3328), .ZN(n4072) );
  MUX2_X1 U5088 ( .A(n4071), .B(n4072), .S(n3332), .Z(n4430) );
  NAND2_X1 U5089 ( .A1(n3285), .A2(n3322), .ZN(n5510) );
  OR2_X1 U5090 ( .A1(n5510), .A2(n3311), .ZN(n4484) );
  NAND2_X1 U5091 ( .A1(n4484), .A2(n4073), .ZN(n4075) );
  BUF_X4 U5092 ( .A(n4074), .Z(n4177) );
  OAI21_X1 U5093 ( .B1(n4075), .B2(n5205), .A(n4253), .ZN(n4082) );
  NAND2_X1 U5094 ( .A1(n4076), .A2(n4077), .ZN(n4079) );
  NAND2_X1 U5095 ( .A1(n4079), .A2(n5350), .ZN(n4081) );
  AND3_X1 U5096 ( .A1(n4082), .A2(n4081), .A3(n4080), .ZN(n4084) );
  NAND3_X1 U5097 ( .A1(n4430), .A2(n4084), .A3(n4083), .ZN(n4476) );
  NOR2_X1 U5098 ( .A1(n4474), .A2(n3328), .ZN(n4085) );
  NAND2_X1 U5099 ( .A1(n4458), .A2(n6654), .ZN(n4088) );
  NAND2_X1 U5101 ( .A1(n4086), .A2(n4527), .ZN(n4087) );
  OAI21_X4 U5102 ( .B1(n4489), .B2(n4088), .A(n4087), .ZN(n6302) );
  NAND2_X2 U5103 ( .A1(n4662), .A2(n6302), .ZN(n5588) );
  MUX2_X1 U5104 ( .A(n5196), .B(n4093), .S(EBX_REG_1__SCAN_IN), .Z(n4092) );
  INV_X1 U5105 ( .A(n4093), .ZN(n4089) );
  NAND2_X1 U5106 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4090)
         );
  AND2_X1 U5107 ( .A1(n4128), .A2(n4090), .ZN(n4091) );
  NAND2_X1 U5108 ( .A1(n4093), .A2(EBX_REG_0__SCAN_IN), .ZN(n4095) );
  INV_X1 U5109 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U5110 ( .A1(n4177), .A2(n5562), .ZN(n4094) );
  NAND2_X1 U5111 ( .A1(n4095), .A2(n4094), .ZN(n4456) );
  MUX2_X1 U5112 ( .A(n5196), .B(n4093), .S(EBX_REG_2__SCAN_IN), .Z(n4097) );
  NAND2_X1 U5113 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4096)
         );
  AND3_X1 U5114 ( .A1(n4097), .A2(n4128), .A3(n4096), .ZN(n4615) );
  NAND2_X1 U5115 ( .A1(n4177), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4100)
         );
  OAI211_X1 U5116 ( .C1(n5204), .C2(EBX_REG_3__SCAN_IN), .A(n4093), .B(n4100), 
        .ZN(n4101) );
  OAI21_X1 U5117 ( .B1(n4170), .B2(EBX_REG_3__SCAN_IN), .A(n4101), .ZN(n4539)
         );
  NOR2_X2 U5118 ( .A1(n4618), .A2(n4539), .ZN(n4603) );
  OR2_X1 U5119 ( .A1(n5196), .A2(EBX_REG_4__SCAN_IN), .ZN(n4105) );
  NAND2_X1 U5120 ( .A1(n4093), .A2(n6420), .ZN(n4103) );
  INV_X1 U5121 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4606) );
  NAND2_X1 U5122 ( .A1(n4527), .A2(n4606), .ZN(n4102) );
  NAND3_X1 U5123 ( .A1(n4103), .A2(n4177), .A3(n4102), .ZN(n4104) );
  NAND2_X1 U5124 ( .A1(n4105), .A2(n4104), .ZN(n4602) );
  NAND2_X1 U5125 ( .A1(n4603), .A2(n4602), .ZN(n4604) );
  MUX2_X1 U5126 ( .A(n4170), .B(n4177), .S(EBX_REG_5__SCAN_IN), .Z(n4106) );
  OAI21_X1 U5127 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n5205), .A(n4106), 
        .ZN(n4549) );
  OR2_X1 U5128 ( .A1(n5196), .A2(EBX_REG_6__SCAN_IN), .ZN(n4111) );
  NAND2_X1 U5129 ( .A1(n4093), .A2(n6062), .ZN(n4109) );
  INV_X1 U5130 ( .A(EBX_REG_6__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U5131 ( .A1(n4527), .A2(n5485), .ZN(n4108) );
  NAND3_X1 U5132 ( .A1(n4109), .A2(n4177), .A3(n4108), .ZN(n4110) );
  AND2_X1 U5133 ( .A1(n4111), .A2(n4110), .ZN(n4633) );
  MUX2_X1 U5134 ( .A(n4170), .B(n4177), .S(EBX_REG_7__SCAN_IN), .Z(n4113) );
  INV_X1 U5135 ( .A(n5205), .ZN(n4176) );
  NAND2_X1 U5136 ( .A1(n6400), .A2(n4176), .ZN(n4112) );
  OR2_X1 U5137 ( .A1(n5196), .A2(EBX_REG_8__SCAN_IN), .ZN(n4117) );
  NAND2_X1 U5138 ( .A1(n4093), .A2(n6046), .ZN(n4115) );
  INV_X1 U5139 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6275) );
  NAND2_X1 U5140 ( .A1(n4527), .A2(n6275), .ZN(n4114) );
  NAND3_X1 U5141 ( .A1(n4115), .A2(n4177), .A3(n4114), .ZN(n4116) );
  NAND2_X1 U5142 ( .A1(n4117), .A2(n4116), .ZN(n4983) );
  NAND2_X1 U5143 ( .A1(n4984), .A2(n4983), .ZN(n4982) );
  NAND2_X1 U5144 ( .A1(n4177), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4118)
         );
  OAI211_X1 U5145 ( .C1(n5204), .C2(EBX_REG_9__SCAN_IN), .A(n4093), .B(n4118), 
        .ZN(n4119) );
  OAI21_X1 U5146 ( .B1(n4170), .B2(EBX_REG_9__SCAN_IN), .A(n4119), .ZN(n6259)
         );
  OR2_X2 U5147 ( .A1(n4982), .A2(n6259), .ZN(n6029) );
  MUX2_X1 U5148 ( .A(n5196), .B(n4093), .S(EBX_REG_10__SCAN_IN), .Z(n4122) );
  NAND2_X1 U5149 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n5204), .ZN(n4120) );
  AND2_X1 U5150 ( .A1(n4128), .A2(n4120), .ZN(n4121) );
  NAND2_X1 U5151 ( .A1(n4122), .A2(n4121), .ZN(n6031) );
  INV_X1 U5152 ( .A(n4170), .ZN(n4161) );
  INV_X1 U5153 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6298) );
  NAND2_X1 U5154 ( .A1(n4161), .A2(n6298), .ZN(n4125) );
  NAND2_X1 U5155 ( .A1(n4177), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4123) );
  OAI211_X1 U5156 ( .C1(n5204), .C2(EBX_REG_11__SCAN_IN), .A(n4093), .B(n4123), 
        .ZN(n4124) );
  AND2_X1 U5157 ( .A1(n4125), .A2(n4124), .ZN(n6030) );
  NAND2_X1 U5158 ( .A1(n6031), .A2(n6030), .ZN(n4126) );
  MUX2_X1 U5159 ( .A(n5196), .B(n4093), .S(EBX_REG_12__SCAN_IN), .Z(n4130) );
  NAND2_X1 U5160 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4127) );
  AND2_X1 U5161 ( .A1(n4128), .A2(n4127), .ZN(n4129) );
  NAND2_X1 U5162 ( .A1(n4130), .A2(n4129), .ZN(n5439) );
  INV_X1 U5163 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U5164 ( .A1(n4161), .A2(n6293), .ZN(n4133) );
  NAND2_X1 U5165 ( .A1(n4177), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4131) );
  OAI211_X1 U5166 ( .C1(n5204), .C2(EBX_REG_13__SCAN_IN), .A(n4093), .B(n4131), 
        .ZN(n4132) );
  AND2_X1 U5167 ( .A1(n4133), .A2(n4132), .ZN(n5438) );
  AND2_X1 U5168 ( .A1(n5439), .A2(n5438), .ZN(n4134) );
  AND2_X2 U5169 ( .A1(n6032), .A2(n4134), .ZN(n5441) );
  MUX2_X1 U5170 ( .A(n5196), .B(n4093), .S(EBX_REG_14__SCAN_IN), .Z(n4136) );
  NAND2_X1 U5171 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4135) );
  NAND2_X1 U5172 ( .A1(n4136), .A2(n4135), .ZN(n5425) );
  NAND2_X1 U5173 ( .A1(n4177), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4137) );
  OAI211_X1 U5174 ( .C1(EBX_REG_15__SCAN_IN), .C2(n5204), .A(n4093), .B(n4137), 
        .ZN(n4138) );
  OAI21_X1 U5175 ( .B1(n4170), .B2(EBX_REG_15__SCAN_IN), .A(n4138), .ZN(n5412)
         );
  MUX2_X1 U5176 ( .A(n5196), .B(n4093), .S(EBX_REG_16__SCAN_IN), .Z(n4140) );
  NAND2_X1 U5177 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4139) );
  NAND2_X1 U5178 ( .A1(n4177), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4141) );
  OAI211_X1 U5179 ( .C1(EBX_REG_17__SCAN_IN), .C2(n5204), .A(n4093), .B(n4141), 
        .ZN(n4142) );
  OAI21_X1 U5180 ( .B1(n4170), .B2(EBX_REG_17__SCAN_IN), .A(n4142), .ZN(n5380)
         );
  MUX2_X1 U5181 ( .A(n5196), .B(n4093), .S(EBX_REG_19__SCAN_IN), .Z(n4144) );
  NAND2_X1 U5182 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n4143) );
  NAND2_X1 U5183 ( .A1(n4144), .A2(n4143), .ZN(n5353) );
  NAND2_X1 U5184 ( .A1(n5379), .A2(n5353), .ZN(n5336) );
  INV_X1 U5185 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6818) );
  OR2_X1 U5186 ( .A1(n5205), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4145)
         );
  INV_X1 U5187 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5583) );
  NAND2_X1 U5188 ( .A1(n4527), .A2(n5583), .ZN(n5349) );
  OR2_X1 U5189 ( .A1(n5205), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4147)
         );
  NAND2_X1 U5190 ( .A1(n4527), .A2(n6818), .ZN(n4146) );
  NAND2_X1 U5191 ( .A1(n4147), .A2(n4146), .ZN(n5337) );
  NAND2_X1 U5192 ( .A1(n5352), .A2(n5337), .ZN(n4150) );
  INV_X1 U5193 ( .A(n5352), .ZN(n4148) );
  NAND2_X1 U5194 ( .A1(n4148), .A2(n4177), .ZN(n4149) );
  OAI211_X1 U5195 ( .C1(n4177), .C2(n6818), .A(n4150), .B(n4149), .ZN(n4151)
         );
  MUX2_X1 U5196 ( .A(n4170), .B(n4177), .S(EBX_REG_21__SCAN_IN), .Z(n4152) );
  OAI21_X1 U5197 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5205), .A(n4152), 
        .ZN(n5324) );
  MUX2_X1 U5198 ( .A(n5196), .B(n4093), .S(EBX_REG_22__SCAN_IN), .Z(n4154) );
  NAND2_X1 U5199 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4153) );
  NAND2_X1 U5200 ( .A1(n4154), .A2(n4153), .ZN(n5311) );
  INV_X1 U5201 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5578) );
  NAND2_X1 U5202 ( .A1(n4161), .A2(n5578), .ZN(n4157) );
  NAND2_X1 U5203 ( .A1(n4177), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4155) );
  OAI211_X1 U5204 ( .C1(EBX_REG_23__SCAN_IN), .C2(n5204), .A(n4093), .B(n4155), 
        .ZN(n4156) );
  AND2_X1 U5205 ( .A1(n4157), .A2(n4156), .ZN(n5299) );
  MUX2_X1 U5206 ( .A(n5196), .B(n4093), .S(EBX_REG_24__SCAN_IN), .Z(n4160) );
  NAND2_X1 U5207 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4159) );
  NAND2_X1 U5208 ( .A1(n4160), .A2(n4159), .ZN(n5288) );
  INV_X1 U5209 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5575) );
  NAND2_X1 U5210 ( .A1(n4161), .A2(n5575), .ZN(n4164) );
  NAND2_X1 U5211 ( .A1(n4177), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4162) );
  OAI211_X1 U5212 ( .C1(EBX_REG_25__SCAN_IN), .C2(n5204), .A(n4093), .B(n4162), 
        .ZN(n4163) );
  AND2_X1 U5213 ( .A1(n4164), .A2(n4163), .ZN(n5272) );
  AND2_X1 U5214 ( .A1(n5288), .A2(n5272), .ZN(n4165) );
  OR2_X1 U5215 ( .A1(n5196), .A2(EBX_REG_26__SCAN_IN), .ZN(n4169) );
  INV_X1 U5216 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n4166) );
  NAND2_X1 U5217 ( .A1(n4093), .A2(n4166), .ZN(n4167) );
  OAI211_X1 U5218 ( .C1(EBX_REG_26__SCAN_IN), .C2(n5204), .A(n4167), .B(n4177), 
        .ZN(n4168) );
  MUX2_X1 U5219 ( .A(n4170), .B(n4177), .S(EBX_REG_27__SCAN_IN), .Z(n4171) );
  OAI21_X1 U5220 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5205), .A(n4171), 
        .ZN(n5252) );
  NOR2_X4 U5221 ( .A1(n5259), .A2(n5252), .ZN(n5254) );
  OR2_X1 U5222 ( .A1(n5196), .A2(EBX_REG_28__SCAN_IN), .ZN(n4174) );
  INV_X1 U5223 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4336) );
  NAND2_X1 U5224 ( .A1(n4093), .A2(n4336), .ZN(n4172) );
  OAI211_X1 U5225 ( .C1(EBX_REG_28__SCAN_IN), .C2(n5204), .A(n4172), .B(n4177), 
        .ZN(n4173) );
  NAND2_X1 U5226 ( .A1(n4174), .A2(n4173), .ZN(n4192) );
  INV_X1 U5227 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5856) );
  NOR2_X1 U5228 ( .A1(n5204), .A2(EBX_REG_29__SCAN_IN), .ZN(n4175) );
  AOI21_X1 U5229 ( .B1(n4176), .B2(n5856), .A(n4175), .ZN(n5227) );
  NAND2_X1 U5230 ( .A1(n5232), .A2(n5227), .ZN(n5195) );
  AND2_X1 U5231 ( .A1(n5195), .A2(n4177), .ZN(n5201) );
  NAND2_X1 U5232 ( .A1(n5195), .A2(n5232), .ZN(n4180) );
  AND2_X1 U5233 ( .A1(n5204), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4178)
         );
  AOI21_X1 U5234 ( .B1(n5205), .B2(EBX_REG_30__SCAN_IN), .A(n4178), .ZN(n5202)
         );
  INV_X1 U5235 ( .A(n5202), .ZN(n4179) );
  NAND2_X1 U5236 ( .A1(n4180), .A2(n4179), .ZN(n4181) );
  OAI211_X1 U5237 ( .C1(n5232), .C2(n4177), .A(n5195), .B(n5202), .ZN(n4182)
         );
  INV_X1 U5238 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4184) );
  OAI21_X1 U5239 ( .B1(n4200), .B2(n5588), .A(n4187), .ZN(U2829) );
  NOR2_X1 U5240 ( .A1(n5254), .A2(n4192), .ZN(n4193) );
  INV_X1 U5241 ( .A(EBX_REG_28__SCAN_IN), .ZN(n4194) );
  INV_X1 U5242 ( .A(n4419), .ZN(n4203) );
  NAND2_X1 U5243 ( .A1(n4451), .A2(n4203), .ZN(n4421) );
  AND3_X1 U5244 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .A3(
        n6694), .ZN(n6649) );
  INV_X1 U5245 ( .A(n6649), .ZN(n4204) );
  NAND2_X1 U5246 ( .A1(n6723), .A2(n3982), .ZN(n6659) );
  NAND3_X1 U5247 ( .A1(n6412), .A2(n4204), .A3(n6659), .ZN(n4205) );
  NAND2_X1 U5248 ( .A1(n4244), .A2(n6267), .ZN(n4236) );
  OR2_X1 U5249 ( .A1(n5547), .A2(n6657), .ZN(n5511) );
  NAND2_X1 U5250 ( .A1(n6692), .A2(n6469), .ZN(n4223) );
  NAND2_X1 U5251 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4223), .ZN(n4207) );
  NAND2_X1 U5252 ( .A1(n3350), .A2(n4906), .ZN(n4438) );
  INV_X1 U5253 ( .A(n4223), .ZN(n4224) );
  AND3_X1 U5254 ( .A1(n4438), .A2(n3328), .A3(n4224), .ZN(n4209) );
  NAND2_X2 U5255 ( .A1(n5211), .A2(n4209), .ZN(n5530) );
  INV_X1 U5256 ( .A(n5547), .ZN(n5504) );
  NAND2_X1 U5257 ( .A1(n5530), .A2(n5504), .ZN(n5564) );
  INV_X1 U5258 ( .A(REIP_REG_14__SCAN_IN), .ZN(n4368) );
  INV_X1 U5259 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6411) );
  NAND3_X1 U5260 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n5512) );
  NOR2_X1 U5261 ( .A1(n6411), .A2(n5512), .ZN(n5462) );
  NAND2_X1 U5262 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5462), .ZN(n5435) );
  NAND2_X1 U5263 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .ZN(
        n5466) );
  NOR2_X1 U5264 ( .A1(n6844), .A2(n5466), .ZN(n5455) );
  NAND4_X1 U5265 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5455), .A3(
        REIP_REG_10__SCAN_IN), .A4(REIP_REG_9__SCAN_IN), .ZN(n5436) );
  NOR2_X1 U5266 ( .A1(n5435), .A2(n5436), .ZN(n5444) );
  NAND3_X1 U5267 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .A3(
        n5444), .ZN(n5420) );
  NOR2_X1 U5268 ( .A1(n4368), .A2(n5420), .ZN(n5421) );
  NAND4_X1 U5269 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5421), .A3(
        REIP_REG_16__SCAN_IN), .A4(REIP_REG_15__SCAN_IN), .ZN(n5355) );
  OR2_X1 U5270 ( .A1(n5547), .A2(n5355), .ZN(n4210) );
  NAND2_X1 U5271 ( .A1(n5564), .A2(n4210), .ZN(n5386) );
  NAND3_X1 U5272 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        REIP_REG_20__SCAN_IN), .ZN(n4213) );
  NAND2_X1 U5273 ( .A1(n5564), .A2(n4213), .ZN(n4211) );
  AND2_X1 U5274 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5314) );
  NAND2_X1 U5275 ( .A1(n5314), .A2(REIP_REG_23__SCAN_IN), .ZN(n4215) );
  NAND2_X1 U5276 ( .A1(n5564), .A2(n4215), .ZN(n4212) );
  NOR2_X1 U5277 ( .A1(n4213), .A2(n5355), .ZN(n4214) );
  NAND2_X1 U5278 ( .A1(n5532), .A2(n4214), .ZN(n5328) );
  OR2_X1 U5279 ( .A1(n4218), .A2(REIP_REG_24__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U5280 ( .A1(n5305), .A2(n5291), .ZN(n5278) );
  NAND2_X1 U5281 ( .A1(REIP_REG_25__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .ZN(
        n4219) );
  AND2_X1 U5282 ( .A1(n5532), .A2(n4219), .ZN(n4216) );
  NAND2_X1 U5283 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n4221) );
  AND2_X1 U5284 ( .A1(n5532), .A2(n4221), .ZN(n4217) );
  NOR2_X1 U5285 ( .A1(n5263), .A2(n4217), .ZN(n5240) );
  INV_X1 U5286 ( .A(n5240), .ZN(n5226) );
  NOR2_X1 U5287 ( .A1(n4218), .A2(n5293), .ZN(n5277) );
  INV_X1 U5288 ( .A(n4219), .ZN(n4220) );
  INV_X1 U5289 ( .A(n4221), .ZN(n4222) );
  NAND2_X1 U5290 ( .A1(n5247), .A2(n4222), .ZN(n5224) );
  XNOR2_X1 U5291 ( .A(REIP_REG_30__SCAN_IN), .B(REIP_REG_29__SCAN_IN), .ZN(
        n4231) );
  NOR2_X1 U5292 ( .A1(n4906), .A2(n4223), .ZN(n6218) );
  NOR2_X1 U5293 ( .A1(n4071), .A2(n6218), .ZN(n5210) );
  NOR2_X1 U5294 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4224), .ZN(n4225) );
  AND2_X1 U5295 ( .A1(n3328), .A2(n4225), .ZN(n4226) );
  NOR2_X1 U5296 ( .A1(n5210), .A2(n4226), .ZN(n4227) );
  OAI22_X1 U5297 ( .A1(n6280), .A2(n4242), .B1(n6251), .B2(n4228), .ZN(n4229)
         );
  AOI21_X1 U5298 ( .B1(EBX_REG_30__SCAN_IN), .B2(n6260), .A(n4229), .ZN(n4230)
         );
  OAI21_X1 U5299 ( .B1(n5224), .B2(n4231), .A(n4230), .ZN(n4232) );
  AOI21_X1 U5300 ( .B1(n5226), .B2(REIP_REG_30__SCAN_IN), .A(n4232), .ZN(n4233) );
  NAND2_X1 U5301 ( .A1(n4236), .A2(n4235), .ZN(U2797) );
  NAND2_X1 U5302 ( .A1(n6723), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6666) );
  NAND2_X1 U5303 ( .A1(n4237), .A2(n6672), .ZN(n6691) );
  NAND2_X1 U5304 ( .A1(n6691), .A2(n6747), .ZN(n4238) );
  NAND2_X1 U5305 ( .A1(n6747), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4240) );
  NAND2_X1 U5306 ( .A1(n6469), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4239) );
  NAND2_X1 U5307 ( .A1(n4240), .A2(n4239), .ZN(n4620) );
  INV_X2 U5308 ( .A(n6412), .ZN(n6364) );
  NAND2_X1 U5309 ( .A1(n6364), .A2(REIP_REG_30__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U5310 ( .A1(n6365), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4241)
         );
  OAI211_X1 U5311 ( .C1(n6375), .C2(n4242), .A(n5847), .B(n4241), .ZN(n4243)
         );
  AOI21_X1 U5312 ( .B1(n4244), .B2(n6370), .A(n4243), .ZN(n4340) );
  NAND2_X1 U5313 ( .A1(n4245), .A2(n4297), .ZN(n4250) );
  NAND2_X1 U5314 ( .A1(n4266), .A2(n4265), .ZN(n4264) );
  NAND2_X1 U5315 ( .A1(n4264), .A2(n4246), .ZN(n4275) );
  INV_X1 U5316 ( .A(n4274), .ZN(n4247) );
  XNOR2_X1 U5317 ( .A(n4275), .B(n4247), .ZN(n4248) );
  NAND2_X1 U5318 ( .A1(n4248), .A2(n4302), .ZN(n4249) );
  NAND2_X1 U5319 ( .A1(n4250), .A2(n4249), .ZN(n4271) );
  INV_X1 U5320 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6429) );
  XNOR2_X1 U5321 ( .A(n4271), .B(n6429), .ZN(n4971) );
  INV_X1 U5322 ( .A(n4251), .ZN(n4256) );
  XNOR2_X1 U5323 ( .A(n4264), .B(n4252), .ZN(n4254) );
  NAND2_X1 U5324 ( .A1(n3285), .A2(n3135), .ZN(n4257) );
  OAI21_X1 U5325 ( .B1(n4254), .B2(n4071), .A(n4257), .ZN(n4255) );
  NAND2_X1 U5326 ( .A1(n4642), .A2(n4297), .ZN(n4260) );
  OAI21_X1 U5327 ( .B1(n4071), .B2(n4266), .A(n4257), .ZN(n4258) );
  INV_X1 U5328 ( .A(n4258), .ZN(n4259) );
  NAND2_X1 U5329 ( .A1(n4428), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4261)
         );
  INV_X1 U5330 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6800) );
  AND2_X1 U5331 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4262) );
  OAI21_X1 U5332 ( .B1(n4266), .B2(n4265), .A(n4264), .ZN(n4267) );
  INV_X1 U5333 ( .A(n4267), .ZN(n4269) );
  NAND3_X1 U5334 ( .A1(n3701), .A2(n3986), .A3(n3135), .ZN(n4268) );
  AOI21_X1 U5335 ( .B1(n4269), .B2(n4302), .A(n4268), .ZN(n4270) );
  INV_X1 U5336 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6440) );
  NAND2_X1 U5337 ( .A1(n4971), .A2(n4970), .ZN(n4973) );
  NAND2_X1 U5338 ( .A1(n4271), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4272)
         );
  NAND2_X1 U5339 ( .A1(n4973), .A2(n4272), .ZN(n6355) );
  NAND2_X1 U5340 ( .A1(n4273), .A2(n4297), .ZN(n4278) );
  NAND2_X1 U5341 ( .A1(n4275), .A2(n4274), .ZN(n4292) );
  XNOR2_X1 U5342 ( .A(n4292), .B(n4290), .ZN(n4276) );
  NAND2_X1 U5343 ( .A1(n4276), .A2(n4302), .ZN(n4277) );
  NAND2_X1 U5344 ( .A1(n4278), .A2(n4277), .ZN(n4279) );
  XNOR2_X1 U5345 ( .A(n4279), .B(n6420), .ZN(n6354) );
  NAND2_X1 U5346 ( .A1(n4279), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4280)
         );
  INV_X1 U5347 ( .A(n4290), .ZN(n4282) );
  OR2_X1 U5348 ( .A1(n4292), .A2(n4282), .ZN(n4283) );
  XNOR2_X1 U5349 ( .A(n4283), .B(n4289), .ZN(n4284) );
  NAND2_X1 U5350 ( .A1(n4284), .A2(n4302), .ZN(n4285) );
  INV_X1 U5351 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U5352 ( .A1(n4286), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n5146)
         );
  NAND3_X1 U5353 ( .A1(n4287), .A2(n4297), .A3(n4288), .ZN(n4295) );
  NAND2_X1 U5354 ( .A1(n4290), .A2(n4289), .ZN(n4291) );
  OR2_X1 U5355 ( .A1(n4292), .A2(n4291), .ZN(n4299) );
  XNOR2_X1 U5356 ( .A(n4299), .B(n4300), .ZN(n4293) );
  NAND2_X1 U5357 ( .A1(n4293), .A2(n4302), .ZN(n4294) );
  NAND2_X1 U5358 ( .A1(n4295), .A2(n4294), .ZN(n5148) );
  NAND2_X1 U5359 ( .A1(n5148), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n5150)
         );
  AND2_X1 U5360 ( .A1(n5146), .A2(n5150), .ZN(n4296) );
  NAND2_X1 U5361 ( .A1(n4298), .A2(n4297), .ZN(n4305) );
  INV_X1 U5362 ( .A(n4299), .ZN(n4301) );
  NAND2_X1 U5363 ( .A1(n4301), .A2(n4300), .ZN(n4317) );
  XNOR2_X1 U5364 ( .A(n4317), .B(n4315), .ZN(n4303) );
  NAND2_X1 U5365 ( .A1(n4303), .A2(n4302), .ZN(n4304) );
  XNOR2_X1 U5366 ( .A(n4309), .B(n6400), .ZN(n5149) );
  INV_X1 U5367 ( .A(n5148), .ZN(n4306) );
  NAND2_X1 U5368 ( .A1(n4306), .A2(n6062), .ZN(n4307) );
  AND2_X1 U5369 ( .A1(n5149), .A2(n4307), .ZN(n4308) );
  NAND2_X1 U5370 ( .A1(n4309), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4310)
         );
  INV_X1 U5371 ( .A(n4311), .ZN(n4313) );
  NOR2_X1 U5372 ( .A1(n4313), .A2(n4312), .ZN(n4314) );
  NAND2_X2 U5373 ( .A1(n4287), .A2(n4314), .ZN(n4329) );
  INV_X1 U5374 ( .A(n4315), .ZN(n4316) );
  OR3_X1 U5375 ( .A1(n4317), .A2(n4316), .A3(n4071), .ZN(n4318) );
  NAND2_X1 U5376 ( .A1(n4329), .A2(n4318), .ZN(n4319) );
  XNOR2_X1 U5377 ( .A(n4319), .B(n6046), .ZN(n5138) );
  NAND2_X1 U5378 ( .A1(n4319), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4320)
         );
  INV_X1 U5379 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6376) );
  NAND2_X1 U5380 ( .A1(n4329), .A2(n6376), .ZN(n5812) );
  OR2_X1 U5381 ( .A1(n4329), .A2(n6376), .ZN(n5813) );
  INV_X1 U5382 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5805) );
  INV_X1 U5383 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6018) );
  AND3_X1 U5384 ( .A1(n5805), .A2(n6036), .A3(n6018), .ZN(n4321) );
  NAND2_X1 U5385 ( .A1(n6026), .A2(n6018), .ZN(n5792) );
  NAND2_X1 U5386 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U5387 ( .A1(n6026), .A2(n5795), .ZN(n4322) );
  XNOR2_X1 U5388 ( .A(n6026), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5787)
         );
  INV_X1 U5389 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U5390 ( .A1(n6026), .A2(n5998), .ZN(n4323) );
  NOR2_X1 U5391 ( .A1(n4329), .A2(n5984), .ZN(n4324) );
  AND2_X1 U5392 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5831) );
  NAND2_X1 U5393 ( .A1(n5831), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4325) );
  INV_X1 U5394 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5947) );
  AND3_X1 U5395 ( .A1(n5973), .A2(n5956), .A3(n5947), .ZN(n4326) );
  OR2_X1 U5396 ( .A1(n6026), .A2(n4326), .ZN(n4327) );
  NAND2_X1 U5397 ( .A1(n5931), .A2(n5910), .ZN(n5702) );
  NAND2_X1 U5398 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5836) );
  OAI21_X1 U5399 ( .B1(n5702), .B2(n5836), .A(n6026), .ZN(n4328) );
  NOR2_X1 U5400 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5930) );
  NOR2_X1 U5401 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5909) );
  INV_X1 U5402 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5900) );
  INV_X1 U5403 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4330) );
  NAND4_X1 U5404 ( .A1(n5930), .A2(n5909), .A3(n5900), .A4(n4330), .ZN(n4331)
         );
  INV_X1 U5405 ( .A(n5686), .ZN(n4333) );
  INV_X1 U5406 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4334) );
  XNOR2_X1 U5407 ( .A(n6026), .B(n4334), .ZN(n5687) );
  NAND2_X1 U5408 ( .A1(n6026), .A2(n4334), .ZN(n4335) );
  NAND2_X1 U5409 ( .A1(n6026), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5675) );
  INV_X1 U5410 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5659) );
  NAND2_X1 U5411 ( .A1(n5659), .A2(n4336), .ZN(n5860) );
  OR2_X1 U5412 ( .A1(n5676), .A2(n5860), .ZN(n5650) );
  NOR2_X1 U5413 ( .A1(n5650), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4337)
         );
  XNOR2_X1 U5414 ( .A(n4338), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5852)
         );
  NAND2_X1 U5415 ( .A1(n4340), .A2(n4339), .ZN(U2956) );
  INV_X1 U5416 ( .A(STATE_REG_1__SCAN_IN), .ZN(n4343) );
  INV_X1 U5417 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4354) );
  NOR2_X1 U5418 ( .A1(n4352), .A2(n4354), .ZN(n4348) );
  AND2_X1 U5419 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n4355) );
  NAND2_X1 U5420 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n4341) );
  OAI21_X1 U5421 ( .B1(n4348), .B2(n4355), .A(n4341), .ZN(n4342) );
  OAI211_X1 U5422 ( .C1(n6692), .C2(n4343), .A(n4342), .B(n4906), .ZN(U3182)
         );
  AOI221_X1 U5423 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6692), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n4344) );
  AOI221_X1 U5424 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n4344), .C2(HOLD), .A(n4352), .ZN(n4351) );
  AND2_X1 U5425 ( .A1(n4347), .A2(n4352), .ZN(n4346) );
  INV_X1 U5426 ( .A(NA_N), .ZN(n4349) );
  NAND2_X1 U5427 ( .A1(n4349), .A2(STATE_REG_2__SCAN_IN), .ZN(n4345) );
  AND2_X1 U5428 ( .A1(n4346), .A2(n4345), .ZN(n4356) );
  AOI22_X1 U5429 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n4360) );
  INV_X1 U5430 ( .A(n4347), .ZN(n4359) );
  AOI21_X1 U5431 ( .B1(n4349), .B2(n4348), .A(n4359), .ZN(n4350) );
  OAI22_X1 U5432 ( .A1(n4351), .A2(n4356), .B1(n4360), .B2(n4350), .ZN(U3183)
         );
  INV_X1 U5433 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6812) );
  NOR2_X1 U5434 ( .A1(n4363), .A2(n6812), .ZN(U3159) );
  INV_X1 U5435 ( .A(DATAWIDTH_REG_29__SCAN_IN), .ZN(n6783) );
  NOR2_X1 U5436 ( .A1(n4363), .A2(n6783), .ZN(U3153) );
  INV_X1 U5437 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6813) );
  NOR2_X1 U5438 ( .A1(n4363), .A2(n6813), .ZN(U3155) );
  INV_X1 U5439 ( .A(DATAWIDTH_REG_11__SCAN_IN), .ZN(n6843) );
  NOR2_X1 U5440 ( .A1(n4363), .A2(n6843), .ZN(U3171) );
  OAI21_X1 U5441 ( .B1(n4355), .B2(n4354), .A(n2966), .ZN(n4358) );
  INV_X1 U5442 ( .A(n4356), .ZN(n4357) );
  OAI211_X1 U5443 ( .C1(n4360), .C2(n4359), .A(n4358), .B(n4357), .ZN(U3181)
         );
  NOR2_X1 U5444 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n4361) );
  OAI21_X1 U5445 ( .B1(BS16_N), .B2(n4361), .A(n4363), .ZN(n4364) );
  OAI21_X1 U5446 ( .B1(n4363), .B2(n6244), .A(n4364), .ZN(U3452) );
  OAI21_X1 U5447 ( .B1(n4363), .B2(n6469), .A(n4364), .ZN(U2792) );
  OAI21_X1 U5448 ( .B1(n4361), .B2(D_C_N_REG_SCAN_IN), .A(n2966), .ZN(n4362)
         );
  OAI21_X1 U5449 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n2966), .A(n4362), .ZN(
        U2791) );
  INV_X1 U5450 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6828) );
  INV_X1 U5451 ( .A(n4363), .ZN(n4366) );
  OAI21_X1 U5452 ( .B1(n4373), .B2(n6828), .A(n4366), .ZN(U2789) );
  INV_X1 U5453 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6231) );
  INV_X1 U5454 ( .A(n4364), .ZN(n4365) );
  AOI21_X1 U5455 ( .B1(n6231), .B2(n4366), .A(n4365), .ZN(U3451) );
  AND2_X1 U5456 ( .A1(n4366), .A2(DATAWIDTH_REG_26__SCAN_IN), .ZN(U3156) );
  AND2_X1 U5457 ( .A1(n4366), .A2(DATAWIDTH_REG_4__SCAN_IN), .ZN(U3178) );
  AND2_X1 U5458 ( .A1(n4366), .A2(DATAWIDTH_REG_22__SCAN_IN), .ZN(U3160) );
  AND2_X1 U5459 ( .A1(n4366), .A2(DATAWIDTH_REG_28__SCAN_IN), .ZN(U3154) );
  AND2_X1 U5460 ( .A1(n4366), .A2(DATAWIDTH_REG_24__SCAN_IN), .ZN(U3158) );
  AND2_X1 U5461 ( .A1(n4366), .A2(DATAWIDTH_REG_31__SCAN_IN), .ZN(U3151) );
  AND2_X1 U5462 ( .A1(n4366), .A2(DATAWIDTH_REG_21__SCAN_IN), .ZN(U3161) );
  AND2_X1 U5463 ( .A1(n4366), .A2(DATAWIDTH_REG_25__SCAN_IN), .ZN(U3157) );
  AND2_X1 U5464 ( .A1(n4366), .A2(DATAWIDTH_REG_30__SCAN_IN), .ZN(U3152) );
  AND2_X1 U5465 ( .A1(n4366), .A2(DATAWIDTH_REG_15__SCAN_IN), .ZN(U3167) );
  AND2_X1 U5466 ( .A1(n4366), .A2(DATAWIDTH_REG_14__SCAN_IN), .ZN(U3168) );
  AND2_X1 U5467 ( .A1(n4366), .A2(DATAWIDTH_REG_13__SCAN_IN), .ZN(U3169) );
  AND2_X1 U5468 ( .A1(n4366), .A2(DATAWIDTH_REG_12__SCAN_IN), .ZN(U3170) );
  AND2_X1 U5469 ( .A1(n4366), .A2(DATAWIDTH_REG_20__SCAN_IN), .ZN(U3162) );
  AND2_X1 U5470 ( .A1(n4366), .A2(DATAWIDTH_REG_10__SCAN_IN), .ZN(U3172) );
  AND2_X1 U5471 ( .A1(n4366), .A2(DATAWIDTH_REG_9__SCAN_IN), .ZN(U3173) );
  AND2_X1 U5472 ( .A1(n4366), .A2(DATAWIDTH_REG_5__SCAN_IN), .ZN(U3177) );
  AND2_X1 U5473 ( .A1(n4366), .A2(DATAWIDTH_REG_8__SCAN_IN), .ZN(U3174) );
  AND2_X1 U5474 ( .A1(n4366), .A2(DATAWIDTH_REG_7__SCAN_IN), .ZN(U3175) );
  AND2_X1 U5475 ( .A1(n4366), .A2(DATAWIDTH_REG_6__SCAN_IN), .ZN(U3176) );
  AND2_X1 U5476 ( .A1(n4366), .A2(DATAWIDTH_REG_17__SCAN_IN), .ZN(U3165) );
  AND2_X1 U5477 ( .A1(n4366), .A2(DATAWIDTH_REG_16__SCAN_IN), .ZN(U3166) );
  AND2_X1 U5478 ( .A1(n4366), .A2(DATAWIDTH_REG_3__SCAN_IN), .ZN(U3179) );
  AND2_X1 U5479 ( .A1(n4366), .A2(DATAWIDTH_REG_2__SCAN_IN), .ZN(U3180) );
  AND2_X1 U5480 ( .A1(n4366), .A2(DATAWIDTH_REG_19__SCAN_IN), .ZN(U3163) );
  AND2_X1 U5481 ( .A1(n4366), .A2(DATAWIDTH_REG_18__SCAN_IN), .ZN(U3164) );
  OR2_X2 U5482 ( .A1(n2966), .A2(n4367), .ZN(n4387) );
  INV_X1 U5483 ( .A(REIP_REG_13__SCAN_IN), .ZN(n4370) );
  INV_X1 U5484 ( .A(ADDRESS_REG_12__SCAN_IN), .ZN(n4369) );
  OAI222_X1 U5485 ( .A1(n4387), .A2(n4370), .B1(n4369), .B2(n4373), .C1(n4372), 
        .C2(n4368), .ZN(U3196) );
  INV_X1 U5486 ( .A(REIP_REG_29__SCAN_IN), .ZN(n4371) );
  INV_X1 U5487 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6737) );
  INV_X1 U5488 ( .A(REIP_REG_30__SCAN_IN), .ZN(n4410) );
  OAI222_X1 U5489 ( .A1(n4387), .A2(n4371), .B1(n4373), .B2(n6737), .C1(n4372), 
        .C2(n4410), .ZN(U3212) );
  INV_X1 U5490 ( .A(REIP_REG_5__SCAN_IN), .ZN(n4403) );
  INV_X1 U5491 ( .A(ADDRESS_REG_3__SCAN_IN), .ZN(n6749) );
  OAI222_X1 U5492 ( .A1(n4387), .A2(n6411), .B1(n4372), .B2(n4403), .C1(n4373), 
        .C2(n6749), .ZN(U3187) );
  INV_X1 U5493 ( .A(REIP_REG_27__SCAN_IN), .ZN(n4400) );
  INV_X1 U5494 ( .A(ADDRESS_REG_25__SCAN_IN), .ZN(n6819) );
  INV_X1 U5495 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6766) );
  OAI222_X1 U5496 ( .A1(n4372), .A2(n4400), .B1(n4373), .B2(n6819), .C1(n4387), 
        .C2(n6766), .ZN(U3209) );
  INV_X2 U5497 ( .A(n4372), .ZN(n4411) );
  AOI22_X1 U5498 ( .A1(n4411), .A2(REIP_REG_15__SCAN_IN), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n2966), .ZN(n4374) );
  OAI21_X1 U5499 ( .B1(n4368), .B2(n4387), .A(n4374), .ZN(U3197) );
  INV_X1 U5500 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6798) );
  AOI22_X1 U5501 ( .A1(n4411), .A2(REIP_REG_13__SCAN_IN), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n2966), .ZN(n4375) );
  OAI21_X1 U5502 ( .B1(n6798), .B2(n4387), .A(n4375), .ZN(U3195) );
  INV_X1 U5503 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5470) );
  AOI22_X1 U5504 ( .A1(n4411), .A2(REIP_REG_11__SCAN_IN), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n2966), .ZN(n4376) );
  OAI21_X1 U5505 ( .B1(n5470), .B2(n4387), .A(n4376), .ZN(U3193) );
  INV_X1 U5506 ( .A(REIP_REG_11__SCAN_IN), .ZN(n4378) );
  AOI22_X1 U5507 ( .A1(n4411), .A2(REIP_REG_12__SCAN_IN), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n2966), .ZN(n4377) );
  OAI21_X1 U5508 ( .B1(n4378), .B2(n4387), .A(n4377), .ZN(U3194) );
  INV_X1 U5509 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6262) );
  AOI22_X1 U5510 ( .A1(n4411), .A2(REIP_REG_10__SCAN_IN), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n2966), .ZN(n4379) );
  OAI21_X1 U5511 ( .B1(n6262), .B2(n4387), .A(n4379), .ZN(U3192) );
  AOI22_X1 U5512 ( .A1(n4411), .A2(REIP_REG_7__SCAN_IN), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n2966), .ZN(n4380) );
  OAI21_X1 U5513 ( .B1(n6844), .B2(n4387), .A(n4380), .ZN(U3189) );
  INV_X1 U5514 ( .A(REIP_REG_7__SCAN_IN), .ZN(n4382) );
  AOI22_X1 U5515 ( .A1(n4411), .A2(REIP_REG_8__SCAN_IN), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n2966), .ZN(n4381) );
  OAI21_X1 U5516 ( .B1(n4382), .B2(n4387), .A(n4381), .ZN(U3190) );
  INV_X1 U5517 ( .A(REIP_REG_8__SCAN_IN), .ZN(n5140) );
  AOI22_X1 U5518 ( .A1(n4411), .A2(REIP_REG_9__SCAN_IN), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n2966), .ZN(n4383) );
  OAI21_X1 U5519 ( .B1(n5140), .B2(n4387), .A(n4383), .ZN(U3191) );
  INV_X1 U5520 ( .A(REIP_REG_2__SCAN_IN), .ZN(n5531) );
  AOI22_X1 U5521 ( .A1(n4411), .A2(REIP_REG_3__SCAN_IN), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n2966), .ZN(n4384) );
  OAI21_X1 U5522 ( .B1(n5531), .B2(n4387), .A(n4384), .ZN(U3185) );
  INV_X1 U5523 ( .A(REIP_REG_3__SCAN_IN), .ZN(n4386) );
  AOI22_X1 U5524 ( .A1(n4411), .A2(REIP_REG_4__SCAN_IN), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n2966), .ZN(n4385) );
  OAI21_X1 U5525 ( .B1(n4386), .B2(n4387), .A(n4385), .ZN(U3186) );
  AOI22_X1 U5526 ( .A1(n4411), .A2(REIP_REG_2__SCAN_IN), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n2966), .ZN(n4388) );
  OAI21_X1 U5527 ( .B1(n6815), .B2(n4387), .A(n4388), .ZN(U3184) );
  INV_X1 U5528 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5332) );
  AOI22_X1 U5529 ( .A1(n4411), .A2(REIP_REG_22__SCAN_IN), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n2966), .ZN(n4389) );
  OAI21_X1 U5530 ( .B1(n5332), .B2(n4387), .A(n4389), .ZN(U3204) );
  INV_X1 U5531 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5407) );
  AOI22_X1 U5532 ( .A1(n4411), .A2(REIP_REG_16__SCAN_IN), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n2966), .ZN(n4390) );
  OAI21_X1 U5533 ( .B1(n5407), .B2(n4387), .A(n4390), .ZN(U3198) );
  INV_X1 U5534 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5382) );
  AOI22_X1 U5535 ( .A1(n4411), .A2(REIP_REG_17__SCAN_IN), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n2966), .ZN(n4391) );
  OAI21_X1 U5536 ( .B1(n5382), .B2(n4387), .A(n4391), .ZN(U3199) );
  INV_X1 U5537 ( .A(REIP_REG_17__SCAN_IN), .ZN(n4393) );
  AOI22_X1 U5538 ( .A1(n4411), .A2(REIP_REG_18__SCAN_IN), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n2966), .ZN(n4392) );
  OAI21_X1 U5539 ( .B1(n4393), .B2(n4387), .A(n4392), .ZN(U3200) );
  INV_X1 U5540 ( .A(REIP_REG_18__SCAN_IN), .ZN(n5339) );
  AOI22_X1 U5541 ( .A1(n4411), .A2(REIP_REG_19__SCAN_IN), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n2966), .ZN(n4394) );
  OAI21_X1 U5542 ( .B1(n5339), .B2(n4387), .A(n4394), .ZN(U3201) );
  INV_X1 U5543 ( .A(REIP_REG_19__SCAN_IN), .ZN(n4396) );
  AOI22_X1 U5544 ( .A1(n4411), .A2(REIP_REG_20__SCAN_IN), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n2966), .ZN(n4395) );
  OAI21_X1 U5545 ( .B1(n4396), .B2(n4387), .A(n4395), .ZN(U3202) );
  INV_X1 U5546 ( .A(REIP_REG_20__SCAN_IN), .ZN(n4398) );
  AOI22_X1 U5547 ( .A1(n4411), .A2(REIP_REG_21__SCAN_IN), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n2966), .ZN(n4397) );
  OAI21_X1 U5548 ( .B1(n4398), .B2(n4387), .A(n4397), .ZN(U3203) );
  AOI22_X1 U5549 ( .A1(n4411), .A2(REIP_REG_28__SCAN_IN), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n2966), .ZN(n4399) );
  OAI21_X1 U5550 ( .B1(n4400), .B2(n4387), .A(n4399), .ZN(U3210) );
  INV_X1 U5551 ( .A(REIP_REG_22__SCAN_IN), .ZN(n5319) );
  AOI22_X1 U5552 ( .A1(n4411), .A2(REIP_REG_23__SCAN_IN), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n2966), .ZN(n4401) );
  OAI21_X1 U5553 ( .B1(n5319), .B2(n4387), .A(n4401), .ZN(U3205) );
  AOI22_X1 U5554 ( .A1(n4411), .A2(REIP_REG_6__SCAN_IN), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n2966), .ZN(n4402) );
  OAI21_X1 U5555 ( .B1(n4403), .B2(n4387), .A(n4402), .ZN(U3188) );
  INV_X1 U5556 ( .A(REIP_REG_25__SCAN_IN), .ZN(n4405) );
  AOI22_X1 U5557 ( .A1(n4411), .A2(REIP_REG_26__SCAN_IN), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n2966), .ZN(n4404) );
  OAI21_X1 U5558 ( .B1(n4405), .B2(n4387), .A(n4404), .ZN(U3208) );
  INV_X1 U5559 ( .A(REIP_REG_23__SCAN_IN), .ZN(n4407) );
  AOI22_X1 U5560 ( .A1(n4411), .A2(REIP_REG_24__SCAN_IN), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n2966), .ZN(n4406) );
  OAI21_X1 U5561 ( .B1(n4407), .B2(n4387), .A(n4406), .ZN(U3206) );
  AOI22_X1 U5562 ( .A1(n4411), .A2(REIP_REG_25__SCAN_IN), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n2966), .ZN(n4408) );
  OAI21_X1 U5563 ( .B1(n5293), .B2(n4387), .A(n4408), .ZN(U3207) );
  AOI22_X1 U5564 ( .A1(n4411), .A2(REIP_REG_31__SCAN_IN), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n2966), .ZN(n4409) );
  OAI21_X1 U5565 ( .B1(n4410), .B2(n4387), .A(n4409), .ZN(U3213) );
  INV_X1 U5566 ( .A(REIP_REG_28__SCAN_IN), .ZN(n4413) );
  AOI22_X1 U5567 ( .A1(n4411), .A2(REIP_REG_29__SCAN_IN), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n2966), .ZN(n4412) );
  OAI21_X1 U5568 ( .B1(n4413), .B2(n4387), .A(n4412), .ZN(U3211) );
  INV_X1 U5569 ( .A(n6209), .ZN(n4414) );
  NOR2_X1 U5570 ( .A1(n4414), .A2(n4696), .ZN(n4448) );
  NAND2_X1 U5571 ( .A1(n4448), .A2(n4420), .ZN(n4417) );
  INV_X1 U5572 ( .A(n4415), .ZN(n4416) );
  AND2_X1 U5573 ( .A1(n4458), .A2(n4416), .ZN(n4697) );
  MUX2_X1 U5574 ( .A(n4417), .B(n4697), .S(n4488), .Z(n4418) );
  AOI21_X1 U5575 ( .B1(n4419), .B2(n4451), .A(n4418), .ZN(n6210) );
  NAND2_X1 U5576 ( .A1(n4421), .A2(n4420), .ZN(n4422) );
  OAI21_X1 U5577 ( .B1(n4488), .B2(n3340), .A(n4422), .ZN(n6224) );
  NAND3_X1 U5578 ( .A1(n5204), .A2(n5491), .A3(n4906), .ZN(n4423) );
  AND2_X1 U5579 ( .A1(n4423), .A2(n6692), .ZN(n6693) );
  NOR2_X1 U5580 ( .A1(n6224), .A2(n6693), .ZN(n6207) );
  OR2_X1 U5581 ( .A1(n6207), .A2(n6223), .ZN(n6227) );
  NAND2_X1 U5582 ( .A1(n6227), .A2(MORE_REG_SCAN_IN), .ZN(n4424) );
  OAI21_X1 U5583 ( .B1(n6210), .B2(n6227), .A(n4424), .ZN(U3471) );
  OR2_X1 U5584 ( .A1(n6672), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5356) );
  NAND2_X1 U5585 ( .A1(n4464), .A2(n5356), .ZN(n6220) );
  INV_X1 U5586 ( .A(READREQUEST_REG_SCAN_IN), .ZN(n5194) );
  NAND2_X1 U5587 ( .A1(n6221), .A2(n5194), .ZN(n4426) );
  NAND3_X1 U5588 ( .A1(n6690), .A2(n5491), .A3(n5204), .ZN(n4425) );
  OAI21_X1 U5589 ( .B1(n6220), .B2(n4426), .A(n4425), .ZN(n4427) );
  INV_X1 U5590 ( .A(n4427), .ZN(U3474) );
  XNOR2_X1 U5591 ( .A(n4428), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4627)
         );
  INV_X1 U5592 ( .A(n4429), .ZN(n4431) );
  NAND2_X1 U5593 ( .A1(n4431), .A2(n4430), .ZN(n4433) );
  INV_X1 U5594 ( .A(n4451), .ZN(n4432) );
  NAND2_X1 U5595 ( .A1(n4433), .A2(n4432), .ZN(n4485) );
  NAND2_X1 U5596 ( .A1(n3322), .A2(n4906), .ZN(n4435) );
  NAND3_X1 U5597 ( .A1(n4435), .A2(n4434), .A3(n3311), .ZN(n4436) );
  NAND3_X1 U5598 ( .A1(n4489), .A2(n4485), .A3(n4436), .ZN(n4437) );
  NAND2_X1 U5599 ( .A1(n4437), .A2(n6654), .ZN(n4444) );
  OR2_X1 U5600 ( .A1(n4047), .A2(READY_N), .ZN(n4482) );
  INV_X1 U5601 ( .A(n4438), .ZN(n4440) );
  OAI211_X1 U5602 ( .C1(n4482), .C2(n4440), .A(n3328), .B(n4439), .ZN(n4441)
         );
  NAND2_X1 U5603 ( .A1(n4441), .A2(n3701), .ZN(n4442) );
  OR2_X1 U5604 ( .A1(n4903), .A2(n4442), .ZN(n4443) );
  INV_X1 U5605 ( .A(n4723), .ZN(n4447) );
  OR2_X1 U5606 ( .A1(n4047), .A2(n5204), .ZN(n4481) );
  NAND2_X1 U5607 ( .A1(n4445), .A2(n3334), .ZN(n4446) );
  NAND4_X1 U5608 ( .A1(n4448), .A2(n4447), .A3(n4481), .A4(n4446), .ZN(n4449)
         );
  INV_X1 U5609 ( .A(n4460), .ZN(n4450) );
  NAND2_X1 U5610 ( .A1(n4450), .A2(n6412), .ZN(n4525) );
  INV_X1 U5611 ( .A(n4525), .ZN(n4453) );
  NAND2_X1 U5612 ( .A1(n4460), .A2(n6196), .ZN(n5994) );
  INV_X1 U5613 ( .A(n5994), .ZN(n4452) );
  OAI21_X1 U5614 ( .B1(n4453), .B2(n4452), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4463) );
  OR2_X1 U5615 ( .A1(n4047), .A2(n4071), .ZN(n6193) );
  NAND2_X1 U5616 ( .A1(n4445), .A2(n3235), .ZN(n4454) );
  NAND2_X1 U5617 ( .A1(n6193), .A2(n4454), .ZN(n4455) );
  OR2_X1 U5618 ( .A1(n5205), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4457)
         );
  NAND2_X1 U5619 ( .A1(n4457), .A2(n4456), .ZN(n5569) );
  INV_X1 U5620 ( .A(n5569), .ZN(n4461) );
  INV_X1 U5621 ( .A(n4458), .ZN(n4459) );
  NAND2_X1 U5622 ( .A1(n4460), .A2(n4459), .ZN(n5999) );
  AND2_X1 U5623 ( .A1(n6016), .A2(n5999), .ZN(n5996) );
  NOR2_X1 U5624 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5996), .ZN(n4523)
         );
  INV_X1 U5625 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6797) );
  NOR2_X1 U5626 ( .A1(n6412), .A2(n6797), .ZN(n4624) );
  AOI211_X1 U5627 ( .C1(n6433), .C2(n4461), .A(n4523), .B(n4624), .ZN(n4462)
         );
  OAI211_X1 U5628 ( .C1(n4627), .C2(n6381), .A(n4463), .B(n4462), .ZN(U3018)
         );
  INV_X1 U5629 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n4923) );
  NAND2_X1 U5630 ( .A1(n4572), .A2(DATAI_0_), .ZN(n4582) );
  NAND2_X1 U5631 ( .A1(n3350), .A2(n4465), .ZN(n4905) );
  NAND2_X1 U5632 ( .A1(n4592), .A2(EAX_REG_16__SCAN_IN), .ZN(n4466) );
  OAI211_X1 U5633 ( .C1(n4551), .C2(n4923), .A(n4582), .B(n4466), .ZN(U2924)
         );
  INV_X1 U5634 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n4910) );
  NAND2_X1 U5635 ( .A1(n4572), .A2(DATAI_1_), .ZN(n4580) );
  NAND2_X1 U5636 ( .A1(n4592), .A2(EAX_REG_17__SCAN_IN), .ZN(n4467) );
  OAI211_X1 U5637 ( .C1(n4551), .C2(n4910), .A(n4580), .B(n4467), .ZN(U2925)
         );
  INV_X1 U5638 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n4913) );
  NAND2_X1 U5639 ( .A1(n4572), .A2(DATAI_2_), .ZN(n4586) );
  NAND2_X1 U5640 ( .A1(n4592), .A2(EAX_REG_18__SCAN_IN), .ZN(n4468) );
  OAI211_X1 U5641 ( .C1(n4551), .C2(n4913), .A(n4586), .B(n4468), .ZN(U2926)
         );
  INV_X1 U5642 ( .A(UWORD_REG_10__SCAN_IN), .ZN(n6781) );
  NAND2_X1 U5643 ( .A1(n4572), .A2(DATAI_10_), .ZN(n4555) );
  NAND2_X1 U5644 ( .A1(n4592), .A2(EAX_REG_26__SCAN_IN), .ZN(n4469) );
  OAI211_X1 U5645 ( .C1(n4551), .C2(n6781), .A(n4555), .B(n4469), .ZN(U2934)
         );
  NAND2_X1 U5646 ( .A1(n4572), .A2(DATAI_9_), .ZN(n4552) );
  NAND2_X1 U5647 ( .A1(n4592), .A2(EAX_REG_25__SCAN_IN), .ZN(n4470) );
  OAI211_X1 U5648 ( .C1(n4551), .C2(n6816), .A(n4552), .B(n4470), .ZN(U2933)
         );
  INV_X1 U5649 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6309) );
  INV_X1 U5650 ( .A(DATAI_15_), .ZN(n6848) );
  INV_X1 U5651 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4471) );
  OAI222_X1 U5652 ( .A1(n4905), .A2(n6309), .B1(n4569), .B2(n6848), .C1(n4471), 
        .C2(n4551), .ZN(U2954) );
  INV_X1 U5653 ( .A(n4472), .ZN(n4473) );
  NAND3_X1 U5654 ( .A1(n4047), .A2(n4474), .A3(n4473), .ZN(n4475) );
  NOR2_X1 U5655 ( .A1(n4723), .A2(n4475), .ZN(n4478) );
  INV_X1 U5656 ( .A(n4476), .ZN(n4477) );
  AND2_X1 U5657 ( .A1(n4478), .A2(n4477), .ZN(n4701) );
  OAI22_X1 U5658 ( .A1(n3501), .A2(n4701), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4510), .ZN(n6195) );
  INV_X1 U5659 ( .A(n6195), .ZN(n4479) );
  INV_X1 U5660 ( .A(n5177), .ZN(n4513) );
  OAI22_X1 U5661 ( .A1(n4479), .A2(n4513), .B1(n4722), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4480) );
  AOI21_X1 U5662 ( .B1(n6647), .B2(n3171), .A(n4480), .ZN(n4495) );
  NAND2_X1 U5663 ( .A1(n6196), .A2(n6692), .ZN(n4483) );
  AOI22_X1 U5664 ( .A1(n4483), .A2(n4482), .B1(n4906), .B2(n4481), .ZN(n4487)
         );
  NAND2_X1 U5665 ( .A1(n4485), .A2(n4484), .ZN(n4486) );
  AOI21_X1 U5666 ( .B1(n4488), .B2(n4487), .A(n4486), .ZN(n4490) );
  AND2_X1 U5667 ( .A1(n4490), .A2(n4489), .ZN(n4493) );
  INV_X1 U5668 ( .A(n4491), .ZN(n4492) );
  NAND2_X1 U5669 ( .A1(n4909), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6665) );
  OAI22_X1 U5670 ( .A1(n6198), .A2(n6223), .B1(n6228), .B2(n6665), .ZN(n4497)
         );
  AOI21_X1 U5671 ( .B1(n6196), .B2(n5177), .A(n5180), .ZN(n4494) );
  OAI22_X1 U5672 ( .A1(n4495), .A2(n5180), .B1(n4494), .B2(n3007), .ZN(U3461)
         );
  INV_X1 U5673 ( .A(n4857), .ZN(n6471) );
  OR2_X1 U5674 ( .A1(n2960), .A2(n6471), .ZN(n4496) );
  XNOR2_X1 U5675 ( .A(n4496), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5514)
         );
  NAND4_X1 U5676 ( .A1(n4497), .A2(n4723), .A3(n5177), .A4(n5514), .ZN(n4498)
         );
  OAI21_X1 U5677 ( .B1(n4032), .B2(n5176), .A(n4498), .ZN(U3455) );
  NAND2_X1 U5678 ( .A1(n4499), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4501) );
  NAND2_X1 U5679 ( .A1(n4501), .A2(n4500), .ZN(n4503) );
  NAND2_X1 U5680 ( .A1(n4503), .A2(n4502), .ZN(n5560) );
  OAI222_X1 U5681 ( .A1(n5560), .A2(n5588), .B1(n6302), .B2(n5562), .C1(n5569), 
        .C2(n6295), .ZN(U2859) );
  INV_X1 U5682 ( .A(n4701), .ZN(n4713) );
  AND2_X1 U5683 ( .A1(n6196), .A2(n3339), .ZN(n4707) );
  INV_X1 U5684 ( .A(n4506), .ZN(n4508) );
  INV_X1 U5685 ( .A(n4507), .ZN(n4514) );
  NAND2_X1 U5686 ( .A1(n4508), .A2(n4514), .ZN(n4509) );
  NOR2_X1 U5687 ( .A1(n4510), .A2(n4509), .ZN(n4511) );
  OR2_X1 U5688 ( .A1(n4707), .A2(n4511), .ZN(n4512) );
  AOI21_X1 U5689 ( .B1(n4505), .B2(n4713), .A(n4512), .ZN(n6197) );
  NOR2_X1 U5690 ( .A1(n6197), .A2(n4513), .ZN(n4518) );
  NAND2_X1 U5691 ( .A1(n6647), .A2(n4514), .ZN(n5173) );
  NAND2_X1 U5692 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n5169) );
  INV_X1 U5693 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4515) );
  AOI22_X1 U5694 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4515), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6800), .ZN(n5170) );
  INV_X1 U5695 ( .A(n5170), .ZN(n4516) );
  OAI22_X1 U5696 ( .A1(n5173), .A2(n4506), .B1(n5169), .B2(n4516), .ZN(n4517)
         );
  OAI21_X1 U5697 ( .B1(n4518), .B2(n4517), .A(n5176), .ZN(n4519) );
  OAI21_X1 U5698 ( .B1(n5176), .B2(n3339), .A(n4519), .ZN(U3460) );
  XNOR2_X1 U5699 ( .A(n4521), .B(n4520), .ZN(n4993) );
  NOR2_X1 U5700 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6380), .ZN(n4531)
         );
  INV_X1 U5701 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4522) );
  NAND2_X1 U5702 ( .A1(n5994), .A2(n4522), .ZN(n5828) );
  INV_X1 U5703 ( .A(n4523), .ZN(n4524) );
  NAND2_X1 U5704 ( .A1(n4525), .A2(n4524), .ZN(n5823) );
  INV_X1 U5705 ( .A(n5823), .ZN(n6057) );
  NAND2_X1 U5706 ( .A1(n6364), .A2(REIP_REG_1__SCAN_IN), .ZN(n4989) );
  OAI21_X1 U5707 ( .B1(n4528), .B2(n4527), .A(n4526), .ZN(n4599) );
  NAND2_X1 U5708 ( .A1(n6433), .A2(n4599), .ZN(n4529) );
  OAI211_X1 U5709 ( .C1(n6057), .C2(n6800), .A(n4989), .B(n4529), .ZN(n4530)
         );
  AOI21_X1 U5710 ( .B1(n4531), .B2(n5828), .A(n4530), .ZN(n4532) );
  OAI21_X1 U5711 ( .B1(n4993), .B2(n6381), .A(n4532), .ZN(U3017) );
  OR2_X1 U5712 ( .A1(n4611), .A2(n4534), .ZN(n4536) );
  NAND2_X1 U5713 ( .A1(n4536), .A2(n4535), .ZN(n4612) );
  INV_X1 U5714 ( .A(n4537), .ZN(n4538) );
  AOI21_X1 U5715 ( .B1(n4533), .B2(n4612), .A(n4538), .ZN(n4976) );
  AND2_X1 U5716 ( .A1(n4618), .A2(n4539), .ZN(n4540) );
  NOR2_X1 U5717 ( .A1(n4603), .A2(n4540), .ZN(n6423) );
  INV_X1 U5718 ( .A(n6423), .ZN(n4541) );
  INV_X1 U5719 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6780) );
  OAI22_X1 U5720 ( .A1(n6295), .A2(n4541), .B1(n6780), .B2(n6302), .ZN(n4542)
         );
  AOI21_X1 U5721 ( .B1(n4976), .B2(n6299), .A(n4542), .ZN(n4543) );
  INV_X1 U5722 ( .A(n4543), .ZN(U2856) );
  OR2_X1 U5723 ( .A1(n4546), .A2(n4545), .ZN(n4547) );
  NAND2_X1 U5724 ( .A1(n4544), .A2(n4547), .ZN(n5502) );
  INV_X1 U5725 ( .A(n4632), .ZN(n4548) );
  AOI21_X1 U5726 ( .B1(n4549), .B2(n4604), .A(n4548), .ZN(n6404) );
  AOI22_X1 U5727 ( .A1(n6404), .A2(n4196), .B1(n5584), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n4550) );
  OAI21_X1 U5728 ( .B1(n5502), .B2(n5588), .A(n4550), .ZN(U2854) );
  INV_X1 U5729 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6318) );
  NAND2_X1 U5730 ( .A1(n4593), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4553) );
  OAI211_X1 U5731 ( .C1(n6318), .C2(n4905), .A(n4553), .B(n4552), .ZN(U2948)
         );
  NAND2_X1 U5732 ( .A1(n4593), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4554) );
  NAND2_X1 U5733 ( .A1(n4572), .A2(DATAI_8_), .ZN(n4584) );
  OAI211_X1 U5734 ( .C1(n6826), .C2(n4905), .A(n4554), .B(n4584), .ZN(U2947)
         );
  INV_X1 U5735 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6316) );
  NAND2_X1 U5736 ( .A1(n4593), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4556) );
  OAI211_X1 U5737 ( .C1(n6316), .C2(n4905), .A(n4556), .B(n4555), .ZN(U2949)
         );
  NAND2_X1 U5738 ( .A1(n4593), .A2(LWORD_REG_12__SCAN_IN), .ZN(n4557) );
  NAND2_X1 U5739 ( .A1(n4572), .A2(DATAI_12_), .ZN(n4563) );
  OAI211_X1 U5740 ( .C1(n6738), .C2(n4905), .A(n4557), .B(n4563), .ZN(U2951)
         );
  INV_X1 U5741 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6804) );
  NAND2_X1 U5742 ( .A1(n4593), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4558) );
  NAND2_X1 U5743 ( .A1(n4572), .A2(DATAI_13_), .ZN(n4566) );
  OAI211_X1 U5744 ( .C1(n6804), .C2(n4905), .A(n4558), .B(n4566), .ZN(U2952)
         );
  AOI22_X1 U5745 ( .A1(n4593), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n4592), .ZN(n4559) );
  NAND2_X1 U5746 ( .A1(n4572), .A2(DATAI_3_), .ZN(n4590) );
  NAND2_X1 U5747 ( .A1(n4559), .A2(n4590), .ZN(U2927) );
  AOI22_X1 U5748 ( .A1(n4593), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n4592), .ZN(n4560) );
  NAND2_X1 U5749 ( .A1(n4572), .A2(DATAI_11_), .ZN(n4561) );
  NAND2_X1 U5750 ( .A1(n4560), .A2(n4561), .ZN(U2950) );
  AOI22_X1 U5751 ( .A1(n4593), .A2(UWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_27__SCAN_IN), .B2(n4592), .ZN(n4562) );
  NAND2_X1 U5752 ( .A1(n4562), .A2(n4561), .ZN(U2935) );
  AOI22_X1 U5753 ( .A1(n4593), .A2(UWORD_REG_12__SCAN_IN), .B1(n4592), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n4564) );
  NAND2_X1 U5754 ( .A1(n4564), .A2(n4563), .ZN(U2936) );
  AOI22_X1 U5755 ( .A1(n4593), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n4592), .ZN(n4565) );
  NAND2_X1 U5756 ( .A1(n4572), .A2(DATAI_5_), .ZN(n4588) );
  NAND2_X1 U5757 ( .A1(n4565), .A2(n4588), .ZN(U2944) );
  AOI22_X1 U5758 ( .A1(n4593), .A2(UWORD_REG_13__SCAN_IN), .B1(n4592), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n4567) );
  NAND2_X1 U5759 ( .A1(n4567), .A2(n4566), .ZN(U2937) );
  AOI22_X1 U5760 ( .A1(n4593), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n4592), .ZN(n4568) );
  OR2_X1 U5761 ( .A1(n4569), .A2(n4666), .ZN(n4594) );
  NAND2_X1 U5762 ( .A1(n4568), .A2(n4594), .ZN(U2930) );
  AOI22_X1 U5763 ( .A1(n4593), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n4592), .ZN(n4570) );
  OR2_X1 U5764 ( .A1(n4569), .A2(n4660), .ZN(n4578) );
  NAND2_X1 U5765 ( .A1(n4570), .A2(n4578), .ZN(U2946) );
  AOI22_X1 U5766 ( .A1(n4593), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n4592), .ZN(n4571) );
  NAND2_X1 U5767 ( .A1(n4572), .A2(DATAI_4_), .ZN(n4574) );
  NAND2_X1 U5768 ( .A1(n4571), .A2(n4574), .ZN(U2928) );
  AOI22_X1 U5769 ( .A1(n4593), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n4592), .ZN(n4573) );
  NAND2_X1 U5770 ( .A1(n4572), .A2(DATAI_14_), .ZN(n4576) );
  NAND2_X1 U5771 ( .A1(n4573), .A2(n4576), .ZN(U2938) );
  AOI22_X1 U5772 ( .A1(n4593), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n4592), .ZN(n4575) );
  NAND2_X1 U5773 ( .A1(n4575), .A2(n4574), .ZN(U2943) );
  AOI22_X1 U5774 ( .A1(n4593), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n4592), .ZN(n4577) );
  NAND2_X1 U5775 ( .A1(n4577), .A2(n4576), .ZN(U2953) );
  AOI22_X1 U5776 ( .A1(n4593), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n4592), .ZN(n4579) );
  NAND2_X1 U5777 ( .A1(n4579), .A2(n4578), .ZN(U2931) );
  AOI22_X1 U5778 ( .A1(n4593), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n4592), .ZN(n4581) );
  NAND2_X1 U5779 ( .A1(n4581), .A2(n4580), .ZN(U2940) );
  AOI22_X1 U5780 ( .A1(n4593), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n4592), .ZN(n4583) );
  NAND2_X1 U5781 ( .A1(n4583), .A2(n4582), .ZN(U2939) );
  AOI22_X1 U5782 ( .A1(n4593), .A2(UWORD_REG_8__SCAN_IN), .B1(n4592), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n4585) );
  NAND2_X1 U5783 ( .A1(n4585), .A2(n4584), .ZN(U2932) );
  AOI22_X1 U5784 ( .A1(n4593), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n4592), .ZN(n4587) );
  NAND2_X1 U5785 ( .A1(n4587), .A2(n4586), .ZN(U2941) );
  AOI22_X1 U5786 ( .A1(n4593), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n4592), .ZN(n4589) );
  NAND2_X1 U5787 ( .A1(n4589), .A2(n4588), .ZN(U2929) );
  AOI22_X1 U5788 ( .A1(n4593), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n4592), .ZN(n4591) );
  NAND2_X1 U5789 ( .A1(n4591), .A2(n4590), .ZN(U2942) );
  AOI22_X1 U5790 ( .A1(n4593), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n4592), .ZN(n4595) );
  NAND2_X1 U5791 ( .A1(n4595), .A2(n4594), .ZN(U2945) );
  OAI21_X1 U5792 ( .B1(n4596), .B2(n4598), .A(n4597), .ZN(n5559) );
  AOI22_X1 U5793 ( .A1(n4196), .A2(n4599), .B1(n5584), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4600) );
  OAI21_X1 U5794 ( .B1(n5559), .B2(n5588), .A(n4600), .ZN(U2858) );
  XNOR2_X1 U5795 ( .A(n4601), .B(n4537), .ZN(n6359) );
  OR2_X1 U5796 ( .A1(n4603), .A2(n4602), .ZN(n4605) );
  AND2_X1 U5797 ( .A1(n4605), .A2(n4604), .ZN(n6414) );
  INV_X1 U5798 ( .A(n6414), .ZN(n5516) );
  OAI22_X1 U5799 ( .A1(n6295), .A2(n5516), .B1(n4606), .B2(n6302), .ZN(n4607)
         );
  INV_X1 U5800 ( .A(n4607), .ZN(n4608) );
  OAI21_X1 U5801 ( .B1(n6359), .B2(n5588), .A(n4608), .ZN(U2855) );
  INV_X1 U5802 ( .A(n4609), .ZN(n4610) );
  NOR2_X1 U5803 ( .A1(n4611), .A2(n4610), .ZN(n4614) );
  INV_X1 U5804 ( .A(n4612), .ZN(n4613) );
  AOI21_X1 U5805 ( .B1(n4614), .B2(n4597), .A(n4613), .ZN(n6371) );
  INV_X1 U5806 ( .A(n6371), .ZN(n4630) );
  NAND2_X1 U5807 ( .A1(n4616), .A2(n4615), .ZN(n4617) );
  AOI22_X1 U5808 ( .A1(n4196), .A2(n6432), .B1(n5584), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4619) );
  OAI21_X1 U5809 ( .B1(n4630), .B2(n5588), .A(n4619), .ZN(U2857) );
  INV_X1 U5810 ( .A(n5560), .ZN(n4625) );
  INV_X1 U5811 ( .A(n4620), .ZN(n4622) );
  INV_X1 U5812 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4621) );
  AOI21_X1 U5813 ( .B1(n5816), .B2(n4622), .A(n4621), .ZN(n4623) );
  AOI211_X1 U5814 ( .C1(n4625), .C2(n6370), .A(n4624), .B(n4623), .ZN(n4626)
         );
  OAI21_X1 U5815 ( .B1(n4627), .B2(n6345), .A(n4626), .ZN(U2986) );
  INV_X1 U5816 ( .A(DATAI_4_), .ZN(n4654) );
  INV_X1 U5817 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6325) );
  OAI222_X1 U5818 ( .A1(n4987), .A2(n6359), .B1(n5647), .B2(n4654), .C1(n5645), 
        .C2(n6325), .ZN(U2887) );
  INV_X1 U5819 ( .A(DATAI_1_), .ZN(n4671) );
  INV_X1 U5820 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6333) );
  OAI222_X1 U5821 ( .A1(n5559), .A2(n4987), .B1(n5647), .B2(n4671), .C1(n5645), 
        .C2(n6333), .ZN(U2890) );
  INV_X1 U5822 ( .A(n4976), .ZN(n5529) );
  INV_X1 U5823 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6327) );
  OAI222_X1 U5824 ( .A1(n5529), .A2(n4987), .B1(n5647), .B2(n4682), .C1(n5645), 
        .C2(n6327), .ZN(U2888) );
  INV_X1 U5825 ( .A(DATAI_2_), .ZN(n4677) );
  INV_X1 U5826 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6329) );
  OAI222_X1 U5827 ( .A1(n4630), .A2(n4987), .B1(n5647), .B2(n4677), .C1(n5645), 
        .C2(n6329), .ZN(U2889) );
  INV_X1 U5828 ( .A(DATAI_5_), .ZN(n4640) );
  INV_X1 U5829 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6324) );
  OAI222_X1 U5830 ( .A1(n5502), .A2(n4987), .B1(n5647), .B2(n4640), .C1(n5645), 
        .C2(n6324), .ZN(U2886) );
  XNOR2_X1 U5831 ( .A(n4544), .B(n3552), .ZN(n5488) );
  INV_X1 U5832 ( .A(n5488), .ZN(n6348) );
  AOI21_X1 U5833 ( .B1(n4633), .B2(n4632), .A(n4965), .ZN(n6065) );
  AOI22_X1 U5834 ( .A1(n6065), .A2(n4196), .B1(n5584), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4634) );
  OAI21_X1 U5835 ( .B1(n6348), .B2(n5588), .A(n4634), .ZN(U2853) );
  NAND2_X1 U5836 ( .A1(n6670), .A2(n6146), .ZN(n4820) );
  OAI21_X1 U5837 ( .B1(n4644), .B2(n6672), .A(n6676), .ZN(n4649) );
  INV_X1 U5838 ( .A(n3501), .ZN(n6552) );
  NAND2_X1 U5839 ( .A1(n6070), .A2(n4636), .ZN(n4822) );
  INV_X1 U5840 ( .A(n4822), .ZN(n6145) );
  NOR2_X1 U5841 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4823) );
  AOI21_X1 U5842 ( .B1(n4749), .B2(n6145), .A(n4646), .ZN(n4648) );
  INV_X1 U5843 ( .A(n4648), .ZN(n4637) );
  NOR2_X1 U5844 ( .A1(n4909), .A2(n6694), .ZN(n4638) );
  INV_X1 U5845 ( .A(n4644), .ZN(n4643) );
  INV_X1 U5846 ( .A(DATAI_21_), .ZN(n4645) );
  NAND2_X1 U5847 ( .A1(n4689), .A2(n3986), .ZN(n6534) );
  INV_X1 U5848 ( .A(n4646), .ZN(n4690) );
  OAI22_X1 U5849 ( .A1(n5015), .A2(n6492), .B1(n6534), .B2(n4690), .ZN(n4647)
         );
  AOI21_X1 U5850 ( .B1(n6624), .B2(n6147), .A(n4647), .ZN(n4653) );
  NAND2_X1 U5851 ( .A1(n4649), .A2(n4648), .ZN(n4651) );
  NOR2_X1 U5852 ( .A1(n5093), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4650)
         );
  NAND2_X1 U5853 ( .A1(n4692), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4652) );
  OAI211_X1 U5854 ( .C1(n4695), .C2(n6580), .A(n4653), .B(n4652), .ZN(U3097)
         );
  INV_X1 U5855 ( .A(DATAI_28_), .ZN(n4655) );
  NOR2_X2 U5856 ( .A1(n6358), .A2(n4655), .ZN(n6617) );
  INV_X1 U5857 ( .A(DATAI_20_), .ZN(n4656) );
  NAND2_X1 U5858 ( .A1(n4689), .A2(n3334), .ZN(n6529) );
  OAI22_X1 U5859 ( .A1(n5015), .A2(n6530), .B1(n6529), .B2(n4690), .ZN(n4657)
         );
  AOI21_X1 U5860 ( .B1(n6617), .B2(n6147), .A(n4657), .ZN(n4659) );
  NAND2_X1 U5861 ( .A1(n4692), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4658) );
  OAI211_X1 U5862 ( .C1(n4695), .C2(n6577), .A(n4659), .B(n4658), .ZN(U3096)
         );
  INV_X1 U5863 ( .A(DATAI_23_), .ZN(n4661) );
  INV_X1 U5864 ( .A(n6639), .ZN(n6501) );
  NAND2_X1 U5865 ( .A1(n4689), .A2(n4662), .ZN(n6545) );
  OAI22_X1 U5866 ( .A1(n5015), .A2(n6501), .B1(n6545), .B2(n4690), .ZN(n4663)
         );
  AOI21_X1 U5867 ( .B1(n6641), .B2(n6147), .A(n4663), .ZN(n4665) );
  NAND2_X1 U5868 ( .A1(n4692), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4664) );
  OAI211_X1 U5869 ( .C1(n4695), .C2(n6590), .A(n4665), .B(n4664), .ZN(U3099)
         );
  INV_X1 U5870 ( .A(DATAI_30_), .ZN(n4667) );
  OAI22_X1 U5871 ( .A1(n5015), .A2(n6540), .B1(n6539), .B2(n4690), .ZN(n4668)
         );
  AOI21_X1 U5872 ( .B1(n6631), .B2(n6147), .A(n4668), .ZN(n4670) );
  NAND2_X1 U5873 ( .A1(n4692), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4669) );
  OAI211_X1 U5874 ( .C1(n4695), .C2(n6583), .A(n4670), .B(n4669), .ZN(U3098)
         );
  INV_X1 U5875 ( .A(DATAI_25_), .ZN(n4672) );
  INV_X1 U5876 ( .A(DATAI_17_), .ZN(n4673) );
  INV_X1 U5877 ( .A(n6595), .ZN(n6704) );
  NAND2_X1 U5878 ( .A1(n4689), .A2(n3322), .ZN(n6699) );
  OAI22_X1 U5879 ( .A1(n5015), .A2(n6704), .B1(n6699), .B2(n4690), .ZN(n4674)
         );
  AOI21_X1 U5880 ( .B1(n6596), .B2(n6147), .A(n4674), .ZN(n4676) );
  NAND2_X1 U5881 ( .A1(n4692), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n4675) );
  OAI211_X1 U5882 ( .C1(n4695), .C2(n6705), .A(n4676), .B(n4675), .ZN(U3093)
         );
  INV_X1 U5883 ( .A(DATAI_26_), .ZN(n4678) );
  NOR2_X2 U5884 ( .A1(n6358), .A2(n4678), .ZN(n6603) );
  NAND2_X1 U5885 ( .A1(n4689), .A2(n3311), .ZN(n6519) );
  OAI22_X1 U5886 ( .A1(n5015), .A2(n6520), .B1(n6519), .B2(n4690), .ZN(n4679)
         );
  AOI21_X1 U5887 ( .B1(n6603), .B2(n6147), .A(n4679), .ZN(n4681) );
  NAND2_X1 U5888 ( .A1(n4692), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4680) );
  OAI211_X1 U5889 ( .C1(n4695), .C2(n6571), .A(n4681), .B(n4680), .ZN(U3094)
         );
  INV_X1 U5890 ( .A(DATAI_27_), .ZN(n4683) );
  NOR2_X2 U5891 ( .A1(n6358), .A2(n4683), .ZN(n6610) );
  NAND2_X1 U5892 ( .A1(n4689), .A2(n3135), .ZN(n6524) );
  OAI22_X1 U5893 ( .A1(n5015), .A2(n6525), .B1(n6524), .B2(n4690), .ZN(n4684)
         );
  AOI21_X1 U5894 ( .B1(n6610), .B2(n6147), .A(n4684), .ZN(n4686) );
  NAND2_X1 U5895 ( .A1(n4692), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4685) );
  OAI211_X1 U5896 ( .C1(n4695), .C2(n6574), .A(n4686), .B(n4685), .ZN(U3095)
         );
  INV_X1 U5897 ( .A(DATAI_0_), .ZN(n4988) );
  INV_X1 U5898 ( .A(DATAI_24_), .ZN(n4687) );
  NAND2_X1 U5899 ( .A1(n4689), .A2(n3328), .ZN(n6506) );
  OAI22_X1 U5900 ( .A1(n5015), .A2(n6481), .B1(n6506), .B2(n4690), .ZN(n4691)
         );
  AOI21_X1 U5901 ( .B1(n6558), .B2(n6147), .A(n4691), .ZN(n4694) );
  NAND2_X1 U5902 ( .A1(n4692), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4693) );
  OAI211_X1 U5903 ( .C1(n4695), .C2(n6566), .A(n4694), .B(n4693), .ZN(U3092)
         );
  OR2_X1 U5904 ( .A1(n4697), .A2(n4696), .ZN(n4704) );
  AOI21_X1 U5905 ( .B1(n4704), .B2(n4507), .A(n4707), .ZN(n4699) );
  NAND2_X1 U5906 ( .A1(n6196), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4698) );
  MUX2_X1 U5907 ( .A(n4699), .B(n4698), .S(n5174), .Z(n4700) );
  NOR2_X1 U5908 ( .A1(n4507), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4702)
         );
  NAND2_X1 U5909 ( .A1(n4704), .A2(n4702), .ZN(n4709) );
  OAI211_X1 U5910 ( .C1(n4701), .C2(n4636), .A(n4700), .B(n4709), .ZN(n5172)
         );
  MUX2_X1 U5911 ( .A(n5172), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(n6198), 
        .Z(n6194) );
  INV_X1 U5912 ( .A(n4702), .ZN(n4703) );
  NAND2_X1 U5913 ( .A1(n4704), .A2(n4703), .ZN(n4706) );
  NAND3_X1 U5914 ( .A1(n6196), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4705) );
  NAND2_X1 U5915 ( .A1(n4706), .A2(n4705), .ZN(n4711) );
  INV_X1 U5916 ( .A(n6196), .ZN(n4902) );
  INV_X1 U5917 ( .A(n4707), .ZN(n4708) );
  OAI211_X1 U5918 ( .C1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(n4902), .A(n4709), .B(n4708), .ZN(n4710) );
  MUX2_X1 U5919 ( .A(n4711), .B(n4710), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4712) );
  INV_X1 U5920 ( .A(n4712), .ZN(n4715) );
  NAND2_X1 U5921 ( .A1(n6144), .A2(n4713), .ZN(n4714) );
  NAND2_X1 U5922 ( .A1(n4715), .A2(n4714), .ZN(n5178) );
  INV_X1 U5923 ( .A(n6198), .ZN(n4716) );
  NAND2_X1 U5924 ( .A1(n5178), .A2(n4716), .ZN(n4718) );
  NAND2_X1 U5925 ( .A1(n6198), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4717) );
  NAND2_X1 U5926 ( .A1(n4718), .A2(n4717), .ZN(n6206) );
  NAND2_X1 U5927 ( .A1(n6194), .A2(n6206), .ZN(n4721) );
  NAND2_X1 U5928 ( .A1(n4719), .A2(n6228), .ZN(n4720) );
  MUX2_X1 U5929 ( .A(n4721), .B(n4720), .S(STATE2_REG_1__SCAN_IN), .Z(n6212)
         );
  MUX2_X1 U5930 ( .A(n6198), .B(n6228), .S(STATE2_REG_1__SCAN_IN), .Z(n4725)
         );
  AND2_X1 U5931 ( .A1(n4723), .A2(n4722), .ZN(n4724) );
  AOI22_X1 U5932 ( .A1(n4725), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(n5514), .B2(n4724), .ZN(n6211) );
  OAI21_X1 U5933 ( .B1(n6212), .B2(n4506), .A(n6211), .ZN(n4727) );
  NOR2_X1 U5934 ( .A1(n4727), .A2(FLUSH_REG_SCAN_IN), .ZN(n4726) );
  INV_X1 U5935 ( .A(n4727), .ZN(n4728) );
  NAND2_X1 U5936 ( .A1(n4728), .A2(n4909), .ZN(n6652) );
  INV_X1 U5937 ( .A(n6652), .ZN(n4731) );
  AND2_X1 U5938 ( .A1(n5093), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6674) );
  OAI22_X1 U5939 ( .A1(n6461), .A2(n6672), .B1(n6674), .B2(n3501), .ZN(n4730)
         );
  OAI21_X1 U5940 ( .B1(n4731), .B2(n4730), .A(n6682), .ZN(n4732) );
  OAI21_X1 U5941 ( .B1(n6682), .B2(n6463), .A(n4732), .ZN(U3465) );
  NAND2_X1 U5942 ( .A1(n6068), .A2(n4733), .ZN(n4734) );
  OAI21_X1 U5943 ( .B1(n4737), .B2(n6358), .A(n6676), .ZN(n4736) );
  AOI21_X1 U5944 ( .B1(n4749), .B2(n6472), .A(n6636), .ZN(n4739) );
  OAI21_X1 U5945 ( .B1(n6515), .B2(n4740), .A(n6513), .ZN(n4735) );
  INV_X1 U5946 ( .A(n6646), .ZN(n4746) );
  INV_X1 U5947 ( .A(n6558), .ZN(n6507) );
  NAND2_X1 U5948 ( .A1(n6640), .A2(n6563), .ZN(n4744) );
  OR2_X1 U5949 ( .A1(n4739), .A2(n6672), .ZN(n4742) );
  NAND2_X1 U5950 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n4740), .ZN(n4741) );
  NAND2_X1 U5951 ( .A1(n4742), .A2(n4741), .ZN(n6638) );
  INV_X1 U5952 ( .A(n6506), .ZN(n6557) );
  AOI22_X1 U5953 ( .A1(n6638), .A2(n6468), .B1(n6636), .B2(n6557), .ZN(n4743)
         );
  OAI211_X1 U5954 ( .C1(n6594), .C2(n6507), .A(n4744), .B(n4743), .ZN(n4745)
         );
  AOI21_X1 U5955 ( .B1(n4746), .B2(INSTQUEUE_REG_15__0__SCAN_IN), .A(n4745), 
        .ZN(n4747) );
  INV_X1 U5956 ( .A(n4747), .ZN(U3140) );
  INV_X1 U5957 ( .A(n4636), .ZN(n5537) );
  NAND2_X1 U5958 ( .A1(n5537), .A2(n6070), .ZN(n5050) );
  INV_X1 U5959 ( .A(n5050), .ZN(n5097) );
  AOI21_X1 U5960 ( .B1(n5097), .B2(n4749), .A(n4754), .ZN(n4757) );
  NOR2_X1 U5961 ( .A1(n4757), .A2(n6672), .ZN(n4750) );
  INV_X1 U5962 ( .A(n4733), .ZN(n4751) );
  OR2_X1 U5963 ( .A1(n4751), .A2(n6068), .ZN(n4752) );
  INV_X1 U5964 ( .A(n4756), .ZN(n4753) );
  INV_X1 U5965 ( .A(n4754), .ZN(n4780) );
  OAI22_X1 U5966 ( .A1(n4862), .A2(n6525), .B1(n6524), .B2(n4780), .ZN(n4755)
         );
  AOI21_X1 U5967 ( .B1(n6610), .B2(n5085), .A(n4755), .ZN(n4761) );
  NOR2_X1 U5968 ( .A1(n4756), .A2(n6469), .ZN(n6669) );
  INV_X1 U5969 ( .A(n6669), .ZN(n4758) );
  NAND3_X1 U5970 ( .A1(n4758), .A2(n6515), .A3(n4757), .ZN(n4759) );
  NAND2_X1 U5971 ( .A1(n4782), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n4760)
         );
  OAI211_X1 U5972 ( .C1(n4785), .C2(n6574), .A(n4761), .B(n4760), .ZN(U3127)
         );
  OAI22_X1 U5973 ( .A1(n4862), .A2(n6501), .B1(n6545), .B2(n4780), .ZN(n4762)
         );
  AOI21_X1 U5974 ( .B1(n6641), .B2(n5085), .A(n4762), .ZN(n4764) );
  NAND2_X1 U5975 ( .A1(n4782), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n4763)
         );
  OAI211_X1 U5976 ( .C1(n4785), .C2(n6590), .A(n4764), .B(n4763), .ZN(U3131)
         );
  OAI22_X1 U5977 ( .A1(n4862), .A2(n6704), .B1(n6699), .B2(n4780), .ZN(n4765)
         );
  AOI21_X1 U5978 ( .B1(n6596), .B2(n5085), .A(n4765), .ZN(n4767) );
  NAND2_X1 U5979 ( .A1(n4782), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4766)
         );
  OAI211_X1 U5980 ( .C1(n4785), .C2(n6705), .A(n4767), .B(n4766), .ZN(U3125)
         );
  OAI22_X1 U5981 ( .A1(n4862), .A2(n6481), .B1(n6506), .B2(n4780), .ZN(n4768)
         );
  AOI21_X1 U5982 ( .B1(n6558), .B2(n5085), .A(n4768), .ZN(n4770) );
  NAND2_X1 U5983 ( .A1(n4782), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4769)
         );
  OAI211_X1 U5984 ( .C1(n4785), .C2(n6566), .A(n4770), .B(n4769), .ZN(U3124)
         );
  OAI22_X1 U5985 ( .A1(n4862), .A2(n6530), .B1(n6529), .B2(n4780), .ZN(n4771)
         );
  AOI21_X1 U5986 ( .B1(n6617), .B2(n5085), .A(n4771), .ZN(n4773) );
  NAND2_X1 U5987 ( .A1(n4782), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4772)
         );
  OAI211_X1 U5988 ( .C1(n4785), .C2(n6577), .A(n4773), .B(n4772), .ZN(U3128)
         );
  OAI22_X1 U5989 ( .A1(n4862), .A2(n6540), .B1(n6539), .B2(n4780), .ZN(n4774)
         );
  AOI21_X1 U5990 ( .B1(n6631), .B2(n5085), .A(n4774), .ZN(n4776) );
  NAND2_X1 U5991 ( .A1(n4782), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4775)
         );
  OAI211_X1 U5992 ( .C1(n4785), .C2(n6583), .A(n4776), .B(n4775), .ZN(U3130)
         );
  OAI22_X1 U5993 ( .A1(n4862), .A2(n6520), .B1(n6519), .B2(n4780), .ZN(n4777)
         );
  AOI21_X1 U5994 ( .B1(n6603), .B2(n5085), .A(n4777), .ZN(n4779) );
  NAND2_X1 U5995 ( .A1(n4782), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4778)
         );
  OAI211_X1 U5996 ( .C1(n4785), .C2(n6571), .A(n4779), .B(n4778), .ZN(U3126)
         );
  OAI22_X1 U5997 ( .A1(n4862), .A2(n6492), .B1(n6534), .B2(n4780), .ZN(n4781)
         );
  AOI21_X1 U5998 ( .B1(n6624), .B2(n5085), .A(n4781), .ZN(n4784) );
  NAND2_X1 U5999 ( .A1(n4782), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4783)
         );
  OAI211_X1 U6000 ( .C1(n4785), .C2(n6580), .A(n4784), .B(n4783), .ZN(U3129)
         );
  OAI21_X1 U6001 ( .B1(n4788), .B2(n6672), .A(n6676), .ZN(n4792) );
  NOR2_X1 U6002 ( .A1(n5050), .A2(n4857), .ZN(n5090) );
  AOI21_X1 U6003 ( .B1(n5090), .B2(n6552), .A(n4789), .ZN(n4791) );
  INV_X1 U6004 ( .A(n4791), .ZN(n4787) );
  INV_X1 U6005 ( .A(n6520), .ZN(n6602) );
  NAND2_X1 U6006 ( .A1(n4788), .A2(n4642), .ZN(n6470) );
  INV_X1 U6007 ( .A(n6603), .ZN(n6162) );
  INV_X1 U6008 ( .A(n4789), .ZN(n4814) );
  OAI22_X1 U6009 ( .A1(n5132), .A2(n6162), .B1(n6519), .B2(n4814), .ZN(n4790)
         );
  AOI21_X1 U6010 ( .B1(n6602), .B2(n6497), .A(n4790), .ZN(n4795) );
  NAND2_X1 U6011 ( .A1(n4792), .A2(n4791), .ZN(n4793) );
  NAND2_X1 U6012 ( .A1(n4816), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4794) );
  OAI211_X1 U6013 ( .C1(n4819), .C2(n6571), .A(n4795), .B(n4794), .ZN(U3062)
         );
  INV_X1 U6014 ( .A(n6596), .ZN(n6701) );
  OAI22_X1 U6015 ( .A1(n5132), .A2(n6701), .B1(n6699), .B2(n4814), .ZN(n4796)
         );
  AOI21_X1 U6016 ( .B1(n6595), .B2(n6497), .A(n4796), .ZN(n4798) );
  NAND2_X1 U6017 ( .A1(n4816), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4797) );
  OAI211_X1 U6018 ( .C1(n4819), .C2(n6705), .A(n4798), .B(n4797), .ZN(U3061)
         );
  OAI22_X1 U6019 ( .A1(n5132), .A2(n6535), .B1(n6534), .B2(n4814), .ZN(n4799)
         );
  AOI21_X1 U6020 ( .B1(n6623), .B2(n6497), .A(n4799), .ZN(n4801) );
  NAND2_X1 U6021 ( .A1(n4816), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4800) );
  OAI211_X1 U6022 ( .C1(n4819), .C2(n6580), .A(n4801), .B(n4800), .ZN(U3065)
         );
  INV_X1 U6023 ( .A(n6525), .ZN(n6609) );
  INV_X1 U6024 ( .A(n6610), .ZN(n6167) );
  OAI22_X1 U6025 ( .A1(n5132), .A2(n6167), .B1(n6524), .B2(n4814), .ZN(n4802)
         );
  AOI21_X1 U6026 ( .B1(n6609), .B2(n6497), .A(n4802), .ZN(n4804) );
  NAND2_X1 U6027 ( .A1(n4816), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4803) );
  OAI211_X1 U6028 ( .C1(n4819), .C2(n6574), .A(n4804), .B(n4803), .ZN(U3063)
         );
  INV_X1 U6029 ( .A(n6641), .ZN(n6546) );
  OAI22_X1 U6030 ( .A1(n5132), .A2(n6546), .B1(n6545), .B2(n4814), .ZN(n4805)
         );
  AOI21_X1 U6031 ( .B1(n6639), .B2(n6497), .A(n4805), .ZN(n4807) );
  NAND2_X1 U6032 ( .A1(n4816), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4806) );
  OAI211_X1 U6033 ( .C1(n4819), .C2(n6590), .A(n4807), .B(n4806), .ZN(U3067)
         );
  INV_X1 U6034 ( .A(n6540), .ZN(n6630) );
  INV_X1 U6035 ( .A(n6631), .ZN(n6181) );
  OAI22_X1 U6036 ( .A1(n5132), .A2(n6181), .B1(n6539), .B2(n4814), .ZN(n4808)
         );
  AOI21_X1 U6037 ( .B1(n6630), .B2(n6497), .A(n4808), .ZN(n4810) );
  NAND2_X1 U6038 ( .A1(n4816), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4809) );
  OAI211_X1 U6039 ( .C1(n4819), .C2(n6583), .A(n4810), .B(n4809), .ZN(U3066)
         );
  INV_X1 U6040 ( .A(n6617), .ZN(n6172) );
  OAI22_X1 U6041 ( .A1(n5132), .A2(n6172), .B1(n6529), .B2(n4814), .ZN(n4811)
         );
  AOI21_X1 U6042 ( .B1(n6616), .B2(n6497), .A(n4811), .ZN(n4813) );
  NAND2_X1 U6043 ( .A1(n4816), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4812) );
  OAI211_X1 U6044 ( .C1(n4819), .C2(n6577), .A(n4813), .B(n4812), .ZN(U3064)
         );
  OAI22_X1 U6045 ( .A1(n5132), .A2(n6507), .B1(n6506), .B2(n4814), .ZN(n4815)
         );
  AOI21_X1 U6046 ( .B1(n6563), .B2(n6497), .A(n4815), .ZN(n4818) );
  NAND2_X1 U6047 ( .A1(n4816), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4817) );
  OAI211_X1 U6048 ( .C1(n4819), .C2(n6566), .A(n4818), .B(n4817), .ZN(U3060)
         );
  INV_X1 U6049 ( .A(n4825), .ZN(n4821) );
  AOI21_X1 U6050 ( .B1(n4821), .B2(STATEBS16_REG_SCAN_IN), .A(n6672), .ZN(
        n4827) );
  NAND2_X1 U6051 ( .A1(n4823), .A2(n6681), .ZN(n4928) );
  OR2_X1 U6052 ( .A1(n4928), .A2(n6463), .ZN(n4851) );
  OAI21_X1 U6053 ( .B1(n4933), .B2(n3501), .A(n4851), .ZN(n4829) );
  INV_X1 U6054 ( .A(n4928), .ZN(n4824) );
  OAI22_X1 U6055 ( .A1(n6110), .A2(n6704), .B1(n6699), .B2(n4851), .ZN(n4826)
         );
  AOI21_X1 U6056 ( .B1(n6596), .B2(n4926), .A(n4826), .ZN(n4832) );
  INV_X1 U6057 ( .A(n4827), .ZN(n4830) );
  NAND2_X1 U6058 ( .A1(n4928), .A2(n6672), .ZN(n4828) );
  NAND2_X1 U6059 ( .A1(n4853), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4831) );
  OAI211_X1 U6060 ( .C1(n4856), .C2(n6705), .A(n4832), .B(n4831), .ZN(U3029)
         );
  OAI22_X1 U6061 ( .A1(n6110), .A2(n6492), .B1(n6534), .B2(n4851), .ZN(n4833)
         );
  AOI21_X1 U6062 ( .B1(n6624), .B2(n4926), .A(n4833), .ZN(n4835) );
  NAND2_X1 U6063 ( .A1(n4853), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4834) );
  OAI211_X1 U6064 ( .C1(n4856), .C2(n6580), .A(n4835), .B(n4834), .ZN(U3033)
         );
  OAI22_X1 U6065 ( .A1(n6110), .A2(n6525), .B1(n6524), .B2(n4851), .ZN(n4836)
         );
  AOI21_X1 U6066 ( .B1(n6610), .B2(n4926), .A(n4836), .ZN(n4838) );
  NAND2_X1 U6067 ( .A1(n4853), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4837) );
  OAI211_X1 U6068 ( .C1(n4856), .C2(n6574), .A(n4838), .B(n4837), .ZN(U3031)
         );
  OAI22_X1 U6069 ( .A1(n6110), .A2(n6501), .B1(n6545), .B2(n4851), .ZN(n4839)
         );
  AOI21_X1 U6070 ( .B1(n6641), .B2(n4926), .A(n4839), .ZN(n4841) );
  NAND2_X1 U6071 ( .A1(n4853), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4840) );
  OAI211_X1 U6072 ( .C1(n4856), .C2(n6590), .A(n4841), .B(n4840), .ZN(U3035)
         );
  OAI22_X1 U6073 ( .A1(n6110), .A2(n6481), .B1(n6506), .B2(n4851), .ZN(n4842)
         );
  AOI21_X1 U6074 ( .B1(n6558), .B2(n4926), .A(n4842), .ZN(n4844) );
  NAND2_X1 U6075 ( .A1(n4853), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4843) );
  OAI211_X1 U6076 ( .C1(n4856), .C2(n6566), .A(n4844), .B(n4843), .ZN(U3028)
         );
  OAI22_X1 U6077 ( .A1(n6110), .A2(n6540), .B1(n6539), .B2(n4851), .ZN(n4845)
         );
  AOI21_X1 U6078 ( .B1(n6631), .B2(n4926), .A(n4845), .ZN(n4847) );
  NAND2_X1 U6079 ( .A1(n4853), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4846) );
  OAI211_X1 U6080 ( .C1(n4856), .C2(n6583), .A(n4847), .B(n4846), .ZN(U3034)
         );
  OAI22_X1 U6081 ( .A1(n6110), .A2(n6530), .B1(n6529), .B2(n4851), .ZN(n4848)
         );
  AOI21_X1 U6082 ( .B1(n6617), .B2(n4926), .A(n4848), .ZN(n4850) );
  NAND2_X1 U6083 ( .A1(n4853), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4849) );
  OAI211_X1 U6084 ( .C1(n4856), .C2(n6577), .A(n4850), .B(n4849), .ZN(U3032)
         );
  OAI22_X1 U6085 ( .A1(n6110), .A2(n6520), .B1(n6519), .B2(n4851), .ZN(n4852)
         );
  AOI21_X1 U6086 ( .B1(n6603), .B2(n4926), .A(n4852), .ZN(n4855) );
  NAND2_X1 U6087 ( .A1(n4853), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4854) );
  OAI211_X1 U6088 ( .C1(n4856), .C2(n6571), .A(n4855), .B(n4854), .ZN(U3030)
         );
  NAND3_X1 U6089 ( .A1(n4862), .A2(n6594), .A3(n6515), .ZN(n4858) );
  AOI22_X1 U6090 ( .A1(n4858), .A2(n6676), .B1(n6472), .B2(n4857), .ZN(n4861)
         );
  NOR2_X1 U6091 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4859), .ZN(n4895)
         );
  INV_X1 U6092 ( .A(n5055), .ZN(n4930) );
  OAI21_X1 U6093 ( .B1(n6464), .B2(n6657), .A(n4930), .ZN(n6078) );
  AOI21_X1 U6094 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6681), .A(n6078), .ZN(
        n5019) );
  OAI211_X1 U6095 ( .C1(n4895), .C2(n5093), .A(n5019), .B(n6139), .ZN(n4860)
         );
  INV_X1 U6096 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4869) );
  INV_X1 U6097 ( .A(n6524), .ZN(n6607) );
  AND2_X1 U6098 ( .A1(n6144), .A2(n6515), .ZN(n6138) );
  NAND2_X1 U6099 ( .A1(n6138), .A2(n6472), .ZN(n4865) );
  INV_X1 U6100 ( .A(n6464), .ZN(n5053) );
  NAND2_X1 U6101 ( .A1(n4863), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6150) );
  OR3_X1 U6102 ( .A1(n5053), .A2(n6150), .A3(n6681), .ZN(n4864) );
  NAND2_X1 U6103 ( .A1(n4865), .A2(n4864), .ZN(n4894) );
  AOI22_X1 U6104 ( .A1(n6607), .A2(n4895), .B1(n4894), .B2(n6608), .ZN(n4866)
         );
  OAI21_X1 U6105 ( .B1(n6594), .B2(n6525), .A(n4866), .ZN(n4867) );
  AOI21_X1 U6106 ( .B1(n6610), .B2(n4898), .A(n4867), .ZN(n4868) );
  OAI21_X1 U6107 ( .B1(n4901), .B2(n4869), .A(n4868), .ZN(U3135) );
  INV_X1 U6108 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4873) );
  INV_X1 U6109 ( .A(n6519), .ZN(n6600) );
  AOI22_X1 U6110 ( .A1(n6600), .A2(n4895), .B1(n4894), .B2(n6601), .ZN(n4870)
         );
  OAI21_X1 U6111 ( .B1(n6594), .B2(n6520), .A(n4870), .ZN(n4871) );
  AOI21_X1 U6112 ( .B1(n6603), .B2(n4898), .A(n4871), .ZN(n4872) );
  OAI21_X1 U6113 ( .B1(n4901), .B2(n4873), .A(n4872), .ZN(U3134) );
  AOI22_X1 U6114 ( .A1(n6621), .A2(n4895), .B1(n4894), .B2(n6622), .ZN(n4874)
         );
  OAI21_X1 U6115 ( .B1(n6594), .B2(n6492), .A(n4874), .ZN(n4875) );
  AOI21_X1 U6116 ( .B1(n6624), .B2(n4898), .A(n4875), .ZN(n4876) );
  OAI21_X1 U6117 ( .B1(n4901), .B2(n4877), .A(n4876), .ZN(U3137) );
  INV_X1 U6118 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4881) );
  AOI22_X1 U6119 ( .A1(n6557), .A2(n4895), .B1(n4894), .B2(n6468), .ZN(n4878)
         );
  OAI21_X1 U6120 ( .B1(n6594), .B2(n6481), .A(n4878), .ZN(n4879) );
  AOI21_X1 U6121 ( .B1(n6558), .B2(n4898), .A(n4879), .ZN(n4880) );
  OAI21_X1 U6122 ( .B1(n4901), .B2(n4881), .A(n4880), .ZN(U3132) );
  INV_X1 U6123 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4885) );
  INV_X1 U6124 ( .A(n6539), .ZN(n6628) );
  AOI22_X1 U6125 ( .A1(n6628), .A2(n4895), .B1(n4894), .B2(n6629), .ZN(n4882)
         );
  OAI21_X1 U6126 ( .B1(n6594), .B2(n6540), .A(n4882), .ZN(n4883) );
  AOI21_X1 U6127 ( .B1(n6631), .B2(n4898), .A(n4883), .ZN(n4884) );
  OAI21_X1 U6128 ( .B1(n4901), .B2(n4885), .A(n4884), .ZN(U3138) );
  INV_X1 U6129 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4889) );
  INV_X1 U6130 ( .A(n6529), .ZN(n6614) );
  AOI22_X1 U6131 ( .A1(n6614), .A2(n4895), .B1(n4894), .B2(n6615), .ZN(n4886)
         );
  OAI21_X1 U6132 ( .B1(n6594), .B2(n6530), .A(n4886), .ZN(n4887) );
  AOI21_X1 U6133 ( .B1(n6617), .B2(n4898), .A(n4887), .ZN(n4888) );
  OAI21_X1 U6134 ( .B1(n4901), .B2(n4889), .A(n4888), .ZN(U3136) );
  INV_X1 U6135 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4893) );
  INV_X1 U6136 ( .A(n6699), .ZN(n6592) );
  AOI22_X1 U6137 ( .A1(n6592), .A2(n4895), .B1(n4894), .B2(n6593), .ZN(n4890)
         );
  OAI21_X1 U6138 ( .B1(n6594), .B2(n6704), .A(n4890), .ZN(n4891) );
  AOI21_X1 U6139 ( .B1(n6596), .B2(n4898), .A(n4891), .ZN(n4892) );
  OAI21_X1 U6140 ( .B1(n4901), .B2(n4893), .A(n4892), .ZN(U3133) );
  INV_X1 U6141 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4900) );
  INV_X1 U6142 ( .A(n6545), .ZN(n6635) );
  AOI22_X1 U6143 ( .A1(n6635), .A2(n4895), .B1(n4894), .B2(n6637), .ZN(n4896)
         );
  OAI21_X1 U6144 ( .B1(n6594), .B2(n6501), .A(n4896), .ZN(n4897) );
  AOI21_X1 U6145 ( .B1(n6641), .B2(n4898), .A(n4897), .ZN(n4899) );
  OAI21_X1 U6146 ( .B1(n4901), .B2(n4900), .A(n4899), .ZN(U3139) );
  INV_X1 U6147 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4912) );
  OR2_X1 U6148 ( .A1(n4903), .A2(n4902), .ZN(n4904) );
  NAND2_X1 U6149 ( .A1(n4905), .A2(n4904), .ZN(n4908) );
  INV_X1 U6150 ( .A(n4906), .ZN(n4907) );
  INV_X1 U6151 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4911) );
  OAI222_X1 U6152 ( .A1(n4912), .A2(n6337), .B1(n5008), .B2(n4911), .C1(n6335), 
        .C2(n4910), .ZN(U2906) );
  INV_X1 U6153 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n4915) );
  INV_X1 U6154 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4914) );
  OAI222_X1 U6155 ( .A1(n4915), .A2(n6337), .B1(n5008), .B2(n4914), .C1(n6335), 
        .C2(n4913), .ZN(U2905) );
  INV_X1 U6156 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4917) );
  INV_X1 U6157 ( .A(UWORD_REG_7__SCAN_IN), .ZN(n4916) );
  OAI222_X1 U6158 ( .A1(n4917), .A2(n6337), .B1(n5008), .B2(n3836), .C1(n6335), 
        .C2(n4916), .ZN(U2900) );
  INV_X1 U6159 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n4920) );
  INV_X1 U6160 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4919) );
  INV_X1 U6161 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n4918) );
  OAI222_X1 U6162 ( .A1(n4920), .A2(n6337), .B1(n5008), .B2(n4919), .C1(n6335), 
        .C2(n4918), .ZN(U2903) );
  INV_X1 U6163 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n4922) );
  INV_X1 U6164 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n4921) );
  OAI222_X1 U6165 ( .A1(n4922), .A2(n6337), .B1(n5008), .B2(n3911), .C1(n6335), 
        .C2(n4921), .ZN(U2896) );
  INV_X1 U6166 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4925) );
  INV_X1 U6167 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4924) );
  OAI222_X1 U6168 ( .A1(n4925), .A2(n6337), .B1(n5008), .B2(n4924), .C1(n6335), 
        .C2(n4923), .ZN(U2907) );
  NOR3_X1 U6169 ( .A1(n4926), .A2(n6640), .A3(n6672), .ZN(n4927) );
  INV_X1 U6170 ( .A(n6676), .ZN(n5051) );
  OAI21_X1 U6171 ( .B1(n4927), .B2(n5051), .A(n4933), .ZN(n4932) );
  INV_X1 U6172 ( .A(n6150), .ZN(n6465) );
  OAI21_X1 U6173 ( .B1(n5098), .B2(n6464), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n4929) );
  NAND2_X1 U6174 ( .A1(n4930), .A2(n4929), .ZN(n5095) );
  AOI211_X1 U6175 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4958), .A(n6465), .B(
        n5095), .ZN(n4931) );
  NAND2_X1 U6176 ( .A1(n4957), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4938) );
  INV_X1 U6177 ( .A(n4933), .ZN(n4935) );
  NOR3_X1 U6178 ( .A1(n5098), .A2(n6464), .A3(n6139), .ZN(n4934) );
  AOI21_X1 U6179 ( .B1(n4935), .B2(n6515), .A(n4934), .ZN(n4959) );
  OAI22_X1 U6180 ( .A1(n4959), .A2(n6571), .B1(n6519), .B2(n4958), .ZN(n4936)
         );
  AOI21_X1 U6181 ( .B1(n6640), .B2(n6603), .A(n4936), .ZN(n4937) );
  OAI211_X1 U6182 ( .C1(n4963), .C2(n6520), .A(n4938), .B(n4937), .ZN(U3022)
         );
  NAND2_X1 U6183 ( .A1(n4957), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4941) );
  OAI22_X1 U6184 ( .A1(n4959), .A2(n6580), .B1(n6534), .B2(n4958), .ZN(n4939)
         );
  AOI21_X1 U6185 ( .B1(n6640), .B2(n6624), .A(n4939), .ZN(n4940) );
  OAI211_X1 U6186 ( .C1(n4963), .C2(n6492), .A(n4941), .B(n4940), .ZN(U3025)
         );
  NAND2_X1 U6187 ( .A1(n4957), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4944) );
  OAI22_X1 U6188 ( .A1(n4959), .A2(n6577), .B1(n6529), .B2(n4958), .ZN(n4942)
         );
  AOI21_X1 U6189 ( .B1(n6640), .B2(n6617), .A(n4942), .ZN(n4943) );
  OAI211_X1 U6190 ( .C1(n4963), .C2(n6530), .A(n4944), .B(n4943), .ZN(U3024)
         );
  NAND2_X1 U6191 ( .A1(n4957), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4947) );
  OAI22_X1 U6192 ( .A1(n4959), .A2(n6566), .B1(n6506), .B2(n4958), .ZN(n4945)
         );
  AOI21_X1 U6193 ( .B1(n6640), .B2(n6558), .A(n4945), .ZN(n4946) );
  OAI211_X1 U6194 ( .C1(n4963), .C2(n6481), .A(n4947), .B(n4946), .ZN(U3020)
         );
  NAND2_X1 U6195 ( .A1(n4957), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4950) );
  OAI22_X1 U6196 ( .A1(n4959), .A2(n6705), .B1(n6699), .B2(n4958), .ZN(n4948)
         );
  AOI21_X1 U6197 ( .B1(n6640), .B2(n6596), .A(n4948), .ZN(n4949) );
  OAI211_X1 U6198 ( .C1(n4963), .C2(n6704), .A(n4950), .B(n4949), .ZN(U3021)
         );
  NAND2_X1 U6199 ( .A1(n4957), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4953) );
  OAI22_X1 U6200 ( .A1(n4959), .A2(n6590), .B1(n6545), .B2(n4958), .ZN(n4951)
         );
  AOI21_X1 U6201 ( .B1(n6640), .B2(n6641), .A(n4951), .ZN(n4952) );
  OAI211_X1 U6202 ( .C1(n4963), .C2(n6501), .A(n4953), .B(n4952), .ZN(U3027)
         );
  NAND2_X1 U6203 ( .A1(n4957), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4956) );
  OAI22_X1 U6204 ( .A1(n4959), .A2(n6574), .B1(n6524), .B2(n4958), .ZN(n4954)
         );
  AOI21_X1 U6205 ( .B1(n6640), .B2(n6610), .A(n4954), .ZN(n4955) );
  OAI211_X1 U6206 ( .C1(n4963), .C2(n6525), .A(n4956), .B(n4955), .ZN(U3023)
         );
  NAND2_X1 U6207 ( .A1(n4957), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4962) );
  OAI22_X1 U6208 ( .A1(n4959), .A2(n6583), .B1(n6539), .B2(n4958), .ZN(n4960)
         );
  AOI21_X1 U6209 ( .B1(n6640), .B2(n6631), .A(n4960), .ZN(n4961) );
  OAI211_X1 U6210 ( .C1(n4963), .C2(n6540), .A(n4962), .B(n4961), .ZN(U3026)
         );
  NOR2_X1 U6211 ( .A1(n4965), .A2(n4964), .ZN(n4966) );
  OR2_X1 U6212 ( .A1(n4984), .A2(n4966), .ZN(n5475) );
  XNOR2_X1 U6213 ( .A(n4968), .B(n4967), .ZN(n5481) );
  INV_X1 U6214 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4969) );
  OAI222_X1 U6215 ( .A1(n5475), .A2(n6295), .B1(n5588), .B2(n5481), .C1(n4969), 
        .C2(n6302), .ZN(U2852) );
  OR2_X1 U6216 ( .A1(n4971), .A2(n4970), .ZN(n4972) );
  NAND2_X1 U6217 ( .A1(n4973), .A2(n4972), .ZN(n6424) );
  NAND2_X1 U6218 ( .A1(n6364), .A2(REIP_REG_3__SCAN_IN), .ZN(n6421) );
  NAND2_X1 U6219 ( .A1(n6365), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4974)
         );
  OAI211_X1 U6220 ( .C1(n6375), .C2(n5522), .A(n6421), .B(n4974), .ZN(n4975)
         );
  AOI21_X1 U6221 ( .B1(n4976), .B2(n6370), .A(n4975), .ZN(n4977) );
  OAI21_X1 U6222 ( .B1(n6345), .B2(n6424), .A(n4977), .ZN(U2983) );
  NOR2_X1 U6223 ( .A1(n2995), .A2(n4979), .ZN(n4980) );
  AOI22_X1 U6224 ( .A1(n5642), .A2(DATAI_8_), .B1(n5641), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4981) );
  OAI21_X1 U6225 ( .B1(n6283), .B2(n4987), .A(n4981), .ZN(U2883) );
  OAI21_X1 U6226 ( .B1(n4984), .B2(n4983), .A(n4982), .ZN(n4985) );
  INV_X1 U6227 ( .A(n4985), .ZN(n6278) );
  AOI22_X1 U6228 ( .A1(n6278), .A2(n4196), .B1(n5584), .B2(EBX_REG_8__SCAN_IN), 
        .ZN(n4986) );
  OAI21_X1 U6229 ( .B1(n6283), .B2(n5588), .A(n4986), .ZN(U2851) );
  INV_X1 U6230 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6746) );
  OAI222_X1 U6231 ( .A1(n5560), .A2(n4987), .B1(n5647), .B2(n4988), .C1(n5645), 
        .C2(n6746), .ZN(U2891) );
  INV_X1 U6232 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5549) );
  OAI21_X1 U6233 ( .B1(n5816), .B2(n5549), .A(n4989), .ZN(n4991) );
  NOR2_X1 U6234 ( .A1(n5559), .A2(n6358), .ZN(n4990) );
  AOI211_X1 U6235 ( .C1(n5818), .C2(n5549), .A(n4991), .B(n4990), .ZN(n4992)
         );
  OAI21_X1 U6236 ( .B1(n4993), .B2(n6345), .A(n4992), .ZN(U2985) );
  OAI222_X1 U6237 ( .A1(n5647), .A2(n4666), .B1(n4987), .B2(n6348), .C1(n4994), 
        .C2(n5645), .ZN(U2885) );
  OAI222_X1 U6238 ( .A1(n5647), .A2(n4660), .B1(n4987), .B2(n5481), .C1(n4995), 
        .C2(n5645), .ZN(U2884) );
  AOI222_X1 U6239 ( .A1(n6330), .A2(DATAO_REG_22__SCAN_IN), .B1(n6306), .B2(
        EAX_REG_22__SCAN_IN), .C1(n6331), .C2(UWORD_REG_6__SCAN_IN), .ZN(n4996) );
  INV_X1 U6240 ( .A(n4996), .ZN(U2901) );
  OAI21_X1 U6241 ( .B1(n4978), .B2(n4998), .A(n3165), .ZN(n6264) );
  AOI22_X1 U6242 ( .A1(n5642), .A2(DATAI_9_), .B1(n5641), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4999) );
  OAI21_X1 U6243 ( .B1(n6264), .B2(n4987), .A(n4999), .ZN(U2882) );
  OAI21_X1 U6244 ( .B1(n5001), .B2(n5000), .A(n5147), .ZN(n6403) );
  NAND2_X1 U6245 ( .A1(n6364), .A2(REIP_REG_5__SCAN_IN), .ZN(n6406) );
  OAI21_X1 U6246 ( .B1(n5816), .B2(n5498), .A(n6406), .ZN(n5003) );
  NOR2_X1 U6247 ( .A1(n5502), .A2(n6358), .ZN(n5002) );
  AOI211_X1 U6248 ( .C1(n5818), .C2(n5495), .A(n5003), .B(n5002), .ZN(n5004)
         );
  OAI21_X1 U6249 ( .B1(n6345), .B2(n6403), .A(n5004), .ZN(U2981) );
  INV_X1 U6250 ( .A(EAX_REG_30__SCAN_IN), .ZN(n5007) );
  NAND2_X1 U6251 ( .A1(n6330), .A2(DATAO_REG_30__SCAN_IN), .ZN(n5006) );
  NAND2_X1 U6252 ( .A1(n6331), .A2(UWORD_REG_14__SCAN_IN), .ZN(n5005) );
  OAI211_X1 U6253 ( .C1(n5008), .C2(n5007), .A(n5006), .B(n5005), .ZN(U2893)
         );
  AOI222_X1 U6254 ( .A1(EAX_REG_28__SCAN_IN), .A2(n6306), .B1(n6330), .B2(
        DATAO_REG_28__SCAN_IN), .C1(n6331), .C2(UWORD_REG_12__SCAN_IN), .ZN(
        n5009) );
  INV_X1 U6255 ( .A(n5009), .ZN(U2895) );
  AOI222_X1 U6256 ( .A1(EAX_REG_24__SCAN_IN), .A2(n6306), .B1(n6330), .B2(
        DATAO_REG_24__SCAN_IN), .C1(n6331), .C2(UWORD_REG_8__SCAN_IN), .ZN(
        n5010) );
  INV_X1 U6257 ( .A(n5010), .ZN(U2899) );
  AOI222_X1 U6258 ( .A1(EAX_REG_21__SCAN_IN), .A2(n6306), .B1(n6330), .B2(
        DATAO_REG_21__SCAN_IN), .C1(n6331), .C2(UWORD_REG_5__SCAN_IN), .ZN(
        n5011) );
  INV_X1 U6259 ( .A(n5011), .ZN(U2902) );
  AOI222_X1 U6260 ( .A1(EAX_REG_29__SCAN_IN), .A2(n6306), .B1(n6330), .B2(
        DATAO_REG_29__SCAN_IN), .C1(n6331), .C2(UWORD_REG_13__SCAN_IN), .ZN(
        n5012) );
  INV_X1 U6261 ( .A(n5012), .ZN(U2894) );
  NAND2_X1 U6262 ( .A1(n6670), .A2(n6068), .ZN(n5049) );
  AOI21_X1 U6263 ( .B1(n5042), .B2(n5015), .A(n6469), .ZN(n5013) );
  NOR2_X1 U6264 ( .A1(n5013), .A2(n6672), .ZN(n5017) );
  AND2_X1 U6265 ( .A1(n4505), .A2(n4636), .ZN(n6076) );
  AND2_X1 U6266 ( .A1(n6076), .A2(n6144), .ZN(n6553) );
  NOR2_X1 U6267 ( .A1(n6139), .A2(n6681), .ZN(n5014) );
  NOR2_X1 U6268 ( .A1(n6117), .A2(n6681), .ZN(n6556) );
  NAND2_X1 U6269 ( .A1(n6556), .A2(n6463), .ZN(n5041) );
  OAI22_X1 U6270 ( .A1(n5042), .A2(n6481), .B1(n5041), .B2(n6506), .ZN(n5016)
         );
  AOI21_X1 U6271 ( .B1(n5044), .B2(n6558), .A(n5016), .ZN(n5022) );
  INV_X1 U6272 ( .A(n5017), .ZN(n5020) );
  AOI21_X1 U6273 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n5041), .A(n6465), .ZN(
        n5018) );
  NAND2_X1 U6274 ( .A1(n5045), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n5021)
         );
  OAI211_X1 U6275 ( .C1(n5048), .C2(n6566), .A(n5022), .B(n5021), .ZN(U3100)
         );
  OAI22_X1 U6276 ( .A1(n5042), .A2(n6525), .B1(n5041), .B2(n6524), .ZN(n5023)
         );
  AOI21_X1 U6277 ( .B1(n5044), .B2(n6610), .A(n5023), .ZN(n5025) );
  NAND2_X1 U6278 ( .A1(n5045), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n5024)
         );
  OAI211_X1 U6279 ( .C1(n5048), .C2(n6574), .A(n5025), .B(n5024), .ZN(U3103)
         );
  OAI22_X1 U6280 ( .A1(n5042), .A2(n6520), .B1(n5041), .B2(n6519), .ZN(n5026)
         );
  AOI21_X1 U6281 ( .B1(n5044), .B2(n6603), .A(n5026), .ZN(n5028) );
  NAND2_X1 U6282 ( .A1(n5045), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n5027)
         );
  OAI211_X1 U6283 ( .C1(n5048), .C2(n6571), .A(n5028), .B(n5027), .ZN(U3102)
         );
  OAI22_X1 U6284 ( .A1(n5042), .A2(n6704), .B1(n5041), .B2(n6699), .ZN(n5029)
         );
  AOI21_X1 U6285 ( .B1(n5044), .B2(n6596), .A(n5029), .ZN(n5031) );
  NAND2_X1 U6286 ( .A1(n5045), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n5030)
         );
  OAI211_X1 U6287 ( .C1(n5048), .C2(n6705), .A(n5031), .B(n5030), .ZN(U3101)
         );
  OAI22_X1 U6288 ( .A1(n5042), .A2(n6540), .B1(n5041), .B2(n6539), .ZN(n5032)
         );
  AOI21_X1 U6289 ( .B1(n5044), .B2(n6631), .A(n5032), .ZN(n5034) );
  NAND2_X1 U6290 ( .A1(n5045), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n5033)
         );
  OAI211_X1 U6291 ( .C1(n5048), .C2(n6583), .A(n5034), .B(n5033), .ZN(U3106)
         );
  OAI22_X1 U6292 ( .A1(n5042), .A2(n6492), .B1(n5041), .B2(n6534), .ZN(n5035)
         );
  AOI21_X1 U6293 ( .B1(n5044), .B2(n6624), .A(n5035), .ZN(n5037) );
  NAND2_X1 U6294 ( .A1(n5045), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n5036)
         );
  OAI211_X1 U6295 ( .C1(n5048), .C2(n6580), .A(n5037), .B(n5036), .ZN(U3105)
         );
  OAI22_X1 U6296 ( .A1(n5042), .A2(n6501), .B1(n5041), .B2(n6545), .ZN(n5038)
         );
  AOI21_X1 U6297 ( .B1(n5044), .B2(n6641), .A(n5038), .ZN(n5040) );
  NAND2_X1 U6298 ( .A1(n5045), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n5039)
         );
  OAI211_X1 U6299 ( .C1(n5048), .C2(n6590), .A(n5040), .B(n5039), .ZN(U3107)
         );
  OAI22_X1 U6300 ( .A1(n5042), .A2(n6530), .B1(n5041), .B2(n6529), .ZN(n5043)
         );
  AOI21_X1 U6301 ( .B1(n5044), .B2(n6617), .A(n5043), .ZN(n5047) );
  NAND2_X1 U6302 ( .A1(n5045), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n5046)
         );
  OAI211_X1 U6303 ( .C1(n5048), .C2(n6577), .A(n5047), .B(n5046), .ZN(U3104)
         );
  NOR3_X1 U6304 ( .A1(n6586), .A2(n5085), .A3(n6672), .ZN(n5052) );
  OAI22_X1 U6305 ( .A1(n5052), .A2(n5051), .B1(n6471), .B2(n5050), .ZN(n5058)
         );
  NAND2_X1 U6306 ( .A1(n5098), .A2(n5053), .ZN(n6140) );
  AND2_X1 U6307 ( .A1(n6140), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5054) );
  NOR2_X1 U6308 ( .A1(n5055), .A2(n5054), .ZN(n6152) );
  NAND2_X1 U6309 ( .A1(n5056), .A2(n6463), .ZN(n5082) );
  NAND2_X1 U6310 ( .A1(n5082), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5057) );
  NAND4_X1 U6311 ( .A1(n5058), .A2(n6152), .A3(n6139), .A4(n5057), .ZN(n5081)
         );
  NAND2_X1 U6312 ( .A1(n5081), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5062)
         );
  INV_X1 U6313 ( .A(n6140), .ZN(n5059) );
  AOI22_X1 U6314 ( .A1(n6138), .A2(n5097), .B1(n6465), .B2(n5059), .ZN(n5083)
         );
  OAI22_X1 U6315 ( .A1(n5083), .A2(n6583), .B1(n6539), .B2(n5082), .ZN(n5060)
         );
  AOI21_X1 U6316 ( .B1(n5085), .B2(n6630), .A(n5060), .ZN(n5061) );
  OAI211_X1 U6317 ( .C1(n5088), .C2(n6181), .A(n5062), .B(n5061), .ZN(U3122)
         );
  NAND2_X1 U6318 ( .A1(n5081), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5065)
         );
  OAI22_X1 U6319 ( .A1(n5083), .A2(n6574), .B1(n6524), .B2(n5082), .ZN(n5063)
         );
  AOI21_X1 U6320 ( .B1(n5085), .B2(n6609), .A(n5063), .ZN(n5064) );
  OAI211_X1 U6321 ( .C1(n5088), .C2(n6167), .A(n5065), .B(n5064), .ZN(U3119)
         );
  NAND2_X1 U6322 ( .A1(n5081), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5068)
         );
  OAI22_X1 U6323 ( .A1(n5083), .A2(n6580), .B1(n6534), .B2(n5082), .ZN(n5066)
         );
  AOI21_X1 U6324 ( .B1(n5085), .B2(n6623), .A(n5066), .ZN(n5067) );
  OAI211_X1 U6325 ( .C1(n5088), .C2(n6535), .A(n5068), .B(n5067), .ZN(U3121)
         );
  NAND2_X1 U6326 ( .A1(n5081), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5071)
         );
  OAI22_X1 U6327 ( .A1(n5083), .A2(n6577), .B1(n6529), .B2(n5082), .ZN(n5069)
         );
  AOI21_X1 U6328 ( .B1(n5085), .B2(n6616), .A(n5069), .ZN(n5070) );
  OAI211_X1 U6329 ( .C1(n5088), .C2(n6172), .A(n5071), .B(n5070), .ZN(U3120)
         );
  NAND2_X1 U6330 ( .A1(n5081), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5074)
         );
  OAI22_X1 U6331 ( .A1(n5083), .A2(n6566), .B1(n6506), .B2(n5082), .ZN(n5072)
         );
  AOI21_X1 U6332 ( .B1(n5085), .B2(n6563), .A(n5072), .ZN(n5073) );
  OAI211_X1 U6333 ( .C1(n5088), .C2(n6507), .A(n5074), .B(n5073), .ZN(U3116)
         );
  NAND2_X1 U6334 ( .A1(n5081), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5077)
         );
  OAI22_X1 U6335 ( .A1(n5083), .A2(n6571), .B1(n6519), .B2(n5082), .ZN(n5075)
         );
  AOI21_X1 U6336 ( .B1(n5085), .B2(n6602), .A(n5075), .ZN(n5076) );
  OAI211_X1 U6337 ( .C1(n5088), .C2(n6162), .A(n5077), .B(n5076), .ZN(U3118)
         );
  NAND2_X1 U6338 ( .A1(n5081), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5080)
         );
  OAI22_X1 U6339 ( .A1(n5083), .A2(n6705), .B1(n6699), .B2(n5082), .ZN(n5078)
         );
  AOI21_X1 U6340 ( .B1(n5085), .B2(n6595), .A(n5078), .ZN(n5079) );
  OAI211_X1 U6341 ( .C1(n5088), .C2(n6701), .A(n5080), .B(n5079), .ZN(U3117)
         );
  NAND2_X1 U6342 ( .A1(n5081), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5087)
         );
  OAI22_X1 U6343 ( .A1(n5083), .A2(n6590), .B1(n6545), .B2(n5082), .ZN(n5084)
         );
  AOI21_X1 U6344 ( .B1(n5085), .B2(n6639), .A(n5084), .ZN(n5086) );
  OAI211_X1 U6345 ( .C1(n5088), .C2(n6546), .A(n5087), .B(n5086), .ZN(U3123)
         );
  NAND3_X1 U6346 ( .A1(n5132), .A2(n6460), .A3(n6515), .ZN(n5091) );
  AOI21_X1 U6347 ( .B1(n5091), .B2(n6676), .A(n5090), .ZN(n5096) );
  OAI21_X1 U6348 ( .B1(n5130), .B2(n5093), .A(n6139), .ZN(n5094) );
  NOR3_X2 U6349 ( .A1(n5096), .A2(n5095), .A3(n5094), .ZN(n5136) );
  INV_X1 U6350 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5104) );
  NAND3_X1 U6351 ( .A1(n5097), .A2(n6675), .A3(n6515), .ZN(n5100) );
  OR3_X1 U6352 ( .A1(n5098), .A2(n6464), .A3(n6150), .ZN(n5099) );
  NAND2_X1 U6353 ( .A1(n5100), .A2(n5099), .ZN(n5129) );
  AOI22_X1 U6354 ( .A1(n6600), .A2(n5130), .B1(n5129), .B2(n6601), .ZN(n5101)
         );
  OAI21_X1 U6355 ( .B1(n5132), .B2(n6520), .A(n5101), .ZN(n5102) );
  AOI21_X1 U6356 ( .B1(n6603), .B2(n5134), .A(n5102), .ZN(n5103) );
  OAI21_X1 U6357 ( .B1(n5136), .B2(n5104), .A(n5103), .ZN(U3054) );
  INV_X1 U6358 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5108) );
  AOI22_X1 U6359 ( .A1(n6628), .A2(n5130), .B1(n5129), .B2(n6629), .ZN(n5105)
         );
  OAI21_X1 U6360 ( .B1(n5132), .B2(n6540), .A(n5105), .ZN(n5106) );
  AOI21_X1 U6361 ( .B1(n6631), .B2(n5134), .A(n5106), .ZN(n5107) );
  OAI21_X1 U6362 ( .B1(n5136), .B2(n5108), .A(n5107), .ZN(U3058) );
  INV_X1 U6363 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5112) );
  AOI22_X1 U6364 ( .A1(n6635), .A2(n5130), .B1(n5129), .B2(n6637), .ZN(n5109)
         );
  OAI21_X1 U6365 ( .B1(n5132), .B2(n6501), .A(n5109), .ZN(n5110) );
  AOI21_X1 U6366 ( .B1(n6641), .B2(n5134), .A(n5110), .ZN(n5111) );
  OAI21_X1 U6367 ( .B1(n5136), .B2(n5112), .A(n5111), .ZN(U3059) );
  INV_X1 U6368 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5116) );
  AOI22_X1 U6369 ( .A1(n6614), .A2(n5130), .B1(n5129), .B2(n6615), .ZN(n5113)
         );
  OAI21_X1 U6370 ( .B1(n5132), .B2(n6530), .A(n5113), .ZN(n5114) );
  AOI21_X1 U6371 ( .B1(n6617), .B2(n5134), .A(n5114), .ZN(n5115) );
  OAI21_X1 U6372 ( .B1(n5136), .B2(n5116), .A(n5115), .ZN(U3056) );
  INV_X1 U6373 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5120) );
  AOI22_X1 U6374 ( .A1(n6621), .A2(n5130), .B1(n5129), .B2(n6622), .ZN(n5117)
         );
  OAI21_X1 U6375 ( .B1(n5132), .B2(n6492), .A(n5117), .ZN(n5118) );
  AOI21_X1 U6376 ( .B1(n6624), .B2(n5134), .A(n5118), .ZN(n5119) );
  OAI21_X1 U6377 ( .B1(n5136), .B2(n5120), .A(n5119), .ZN(U3057) );
  INV_X1 U6378 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5124) );
  AOI22_X1 U6379 ( .A1(n6557), .A2(n5130), .B1(n5129), .B2(n6468), .ZN(n5121)
         );
  OAI21_X1 U6380 ( .B1(n5132), .B2(n6481), .A(n5121), .ZN(n5122) );
  AOI21_X1 U6381 ( .B1(n6558), .B2(n5134), .A(n5122), .ZN(n5123) );
  OAI21_X1 U6382 ( .B1(n5136), .B2(n5124), .A(n5123), .ZN(U3052) );
  INV_X1 U6383 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5128) );
  AOI22_X1 U6384 ( .A1(n6607), .A2(n5130), .B1(n5129), .B2(n6608), .ZN(n5125)
         );
  OAI21_X1 U6385 ( .B1(n5132), .B2(n6525), .A(n5125), .ZN(n5126) );
  AOI21_X1 U6386 ( .B1(n6610), .B2(n5134), .A(n5126), .ZN(n5127) );
  OAI21_X1 U6387 ( .B1(n5136), .B2(n5128), .A(n5127), .ZN(U3055) );
  AOI22_X1 U6388 ( .A1(n6592), .A2(n5130), .B1(n5129), .B2(n6593), .ZN(n5131)
         );
  OAI21_X1 U6389 ( .B1(n5132), .B2(n6704), .A(n5131), .ZN(n5133) );
  AOI21_X1 U6390 ( .B1(n6596), .B2(n5134), .A(n5133), .ZN(n5135) );
  OAI21_X1 U6391 ( .B1(n5136), .B2(n6752), .A(n5135), .ZN(U3053) );
  OAI21_X1 U6392 ( .B1(n5139), .B2(n5138), .A(n5137), .ZN(n6051) );
  INV_X1 U6393 ( .A(n6283), .ZN(n5144) );
  NOR2_X1 U6394 ( .A1(n6412), .A2(n5140), .ZN(n6049) );
  INV_X1 U6395 ( .A(n6049), .ZN(n5142) );
  NAND2_X1 U6396 ( .A1(n6365), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5141)
         );
  OAI211_X1 U6397 ( .C1(n6375), .C2(n6281), .A(n5142), .B(n5141), .ZN(n5143)
         );
  AOI21_X1 U6398 ( .B1(n5144), .B2(n6370), .A(n5143), .ZN(n5145) );
  OAI21_X1 U6399 ( .B1(n6345), .B2(n6051), .A(n5145), .ZN(U2978) );
  NAND2_X1 U6400 ( .A1(n5147), .A2(n5146), .ZN(n6053) );
  XNOR2_X1 U6401 ( .A(n5148), .B(n6062), .ZN(n6052) );
  NAND2_X1 U6402 ( .A1(n6053), .A2(n6052), .ZN(n6055) );
  INV_X1 U6403 ( .A(n5149), .ZN(n5151) );
  NAND3_X1 U6404 ( .A1(n6055), .A2(n5151), .A3(n5150), .ZN(n5153) );
  NAND2_X1 U6405 ( .A1(n6396), .A2(n6369), .ZN(n5156) );
  NOR2_X1 U6406 ( .A1(n6412), .A2(n4382), .ZN(n6394) );
  NOR2_X1 U6407 ( .A1(n6375), .A2(n5473), .ZN(n5154) );
  AOI211_X1 U6408 ( .C1(n6365), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6394), 
        .B(n5154), .ZN(n5155) );
  OAI211_X1 U6409 ( .C1(n5481), .C2(n6358), .A(n5156), .B(n5155), .ZN(U2979)
         );
  OAI21_X1 U6410 ( .B1(n4997), .B2(n3607), .A(n5158), .ZN(n5811) );
  XNOR2_X1 U6411 ( .A(n6029), .B(n6031), .ZN(n6378) );
  AOI22_X1 U6412 ( .A1(n6378), .A2(n4196), .B1(EBX_REG_10__SCAN_IN), .B2(n5584), .ZN(n5159) );
  OAI21_X1 U6413 ( .B1(n5811), .B2(n5588), .A(n5159), .ZN(U2849) );
  AOI22_X1 U6414 ( .A1(n5642), .A2(DATAI_10_), .B1(n5641), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5160) );
  OAI21_X1 U6415 ( .B1(n5811), .B2(n4987), .A(n5160), .ZN(U2881) );
  AND2_X1 U6416 ( .A1(n5158), .A2(n5161), .ZN(n5162) );
  OR2_X1 U6417 ( .A1(n5162), .A2(n2967), .ZN(n6341) );
  AOI22_X1 U6418 ( .A1(n5642), .A2(DATAI_11_), .B1(n5641), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5163) );
  OAI21_X1 U6419 ( .B1(n6341), .B2(n4987), .A(n5163), .ZN(U2880) );
  XOR2_X1 U6420 ( .A(n2967), .B(n5164), .Z(n5802) );
  INV_X1 U6421 ( .A(n5802), .ZN(n5454) );
  INV_X1 U6422 ( .A(n5439), .ZN(n5165) );
  XNOR2_X1 U6423 ( .A(n6032), .B(n5165), .ZN(n6014) );
  AOI22_X1 U6424 ( .A1(n6014), .A2(n4196), .B1(n5584), .B2(EBX_REG_12__SCAN_IN), .ZN(n5166) );
  OAI21_X1 U6425 ( .B1(n5454), .B2(n5588), .A(n5166), .ZN(U2847) );
  AOI22_X1 U6426 ( .A1(n5642), .A2(DATAI_12_), .B1(n5641), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5167) );
  OAI21_X1 U6427 ( .B1(n5454), .B2(n4987), .A(n5167), .ZN(U2879) );
  NAND3_X1 U6428 ( .A1(n6647), .A2(n4507), .A3(n5174), .ZN(n5168) );
  OAI21_X1 U6429 ( .B1(n5170), .B2(n5169), .A(n5168), .ZN(n5171) );
  AOI21_X1 U6430 ( .B1(n5172), .B2(n5177), .A(n5171), .ZN(n5175) );
  AND2_X1 U6431 ( .A1(n5173), .A2(n5176), .ZN(n5185) );
  OAI22_X1 U6432 ( .A1(n5175), .A2(n5180), .B1(n5185), .B2(n5174), .ZN(U3459)
         );
  NAND3_X1 U6433 ( .A1(n5178), .A2(n5177), .A3(n5176), .ZN(n5184) );
  NOR2_X1 U6434 ( .A1(n5181), .A2(n5180), .ZN(n5182) );
  OAI21_X1 U6435 ( .B1(n5179), .B2(n5182), .A(n6647), .ZN(n5183) );
  OAI211_X1 U6436 ( .C1(n5185), .C2(n3018), .A(n5184), .B(n5183), .ZN(U3456)
         );
  OR2_X1 U6437 ( .A1(n4329), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5186)
         );
  NOR2_X1 U6438 ( .A1(n5684), .A2(n5186), .ZN(n5658) );
  NOR4_X1 U6439 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A3(INSTADDRPOINTER_REG_28__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5187) );
  INV_X1 U6440 ( .A(EAX_REG_31__SCAN_IN), .ZN(n5595) );
  OAI22_X1 U6441 ( .A1(n3674), .A2(n5595), .B1(n5188), .B2(n5213), .ZN(n5592)
         );
  NAND2_X1 U6442 ( .A1(n6364), .A2(REIP_REG_31__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U6443 ( .A1(n6365), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5190)
         );
  OAI211_X1 U6444 ( .C1(n5191), .C2(n6375), .A(n5839), .B(n5190), .ZN(n5192)
         );
  OAI21_X1 U6445 ( .B1(n5844), .B2(n6345), .A(n5193), .ZN(U2955) );
  MUX2_X1 U6446 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n2966), .Z(U3473) );
  MUX2_X1 U6447 ( .A(n5194), .B(W_R_N_REG_SCAN_IN), .S(n2966), .Z(U3470) );
  OR2_X1 U6448 ( .A1(n5195), .A2(n5350), .ZN(n5200) );
  INV_X1 U6449 ( .A(n5196), .ZN(n5198) );
  INV_X1 U6450 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5197) );
  AND2_X1 U6451 ( .A1(n5198), .A2(n5197), .ZN(n5228) );
  NAND2_X1 U6452 ( .A1(n5232), .A2(n5228), .ZN(n5199) );
  AOI21_X1 U6453 ( .B1(n5202), .B2(n5234), .A(n5201), .ZN(n5203) );
  OAI22_X1 U6454 ( .A1(n5205), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5204), .ZN(n5206) );
  NAND2_X1 U6455 ( .A1(n5209), .A2(n6267), .ZN(n5220) );
  AND2_X1 U6456 ( .A1(REIP_REG_30__SCAN_IN), .A2(REIP_REG_29__SCAN_IN), .ZN(
        n5214) );
  OAI21_X1 U6457 ( .B1(n5214), .B2(n5530), .A(n5240), .ZN(n5218) );
  NAND3_X1 U6458 ( .A1(n5211), .A2(EBX_REG_31__SCAN_IN), .A3(n5210), .ZN(n5212) );
  OAI21_X1 U6459 ( .B1(n6251), .B2(n5213), .A(n5212), .ZN(n5217) );
  INV_X1 U6460 ( .A(n5214), .ZN(n5215) );
  NOR3_X1 U6461 ( .A1(n5224), .A2(REIP_REG_31__SCAN_IN), .A3(n5215), .ZN(n5216) );
  AOI211_X1 U6462 ( .C1(n5218), .C2(REIP_REG_31__SCAN_IN), .A(n5217), .B(n5216), .ZN(n5219) );
  OAI211_X1 U6463 ( .C1(n5572), .C2(n5570), .A(n5220), .B(n5219), .ZN(U2796)
         );
  AOI21_X1 U6464 ( .B1(n5221), .B2(n4188), .A(n5590), .ZN(n5656) );
  INV_X1 U6465 ( .A(n5656), .ZN(n5603) );
  AOI22_X1 U6466 ( .A1(n6266), .A2(n5652), .B1(n6273), .B2(
        PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5223) );
  NAND2_X1 U6467 ( .A1(n6260), .A2(EBX_REG_29__SCAN_IN), .ZN(n5222) );
  OAI211_X1 U6468 ( .C1(n5224), .C2(REIP_REG_29__SCAN_IN), .A(n5223), .B(n5222), .ZN(n5225) );
  AOI21_X1 U6469 ( .B1(n5226), .B2(REIP_REG_29__SCAN_IN), .A(n5225), .ZN(n5236) );
  NAND2_X1 U6470 ( .A1(n5227), .A2(n4177), .ZN(n5230) );
  INV_X1 U6471 ( .A(n5228), .ZN(n5229) );
  NAND2_X1 U6472 ( .A1(n5230), .A2(n5229), .ZN(n5231) );
  NOR2_X1 U6473 ( .A1(n5232), .A2(n5231), .ZN(n5233) );
  NAND2_X1 U6474 ( .A1(n3138), .A2(n6279), .ZN(n5235) );
  OAI211_X1 U6475 ( .C1(n5603), .C2(n6282), .A(n5236), .B(n5235), .ZN(U2798)
         );
  AOI21_X1 U6476 ( .B1(n5247), .B2(REIP_REG_27__SCAN_IN), .A(
        REIP_REG_28__SCAN_IN), .ZN(n5239) );
  AOI22_X1 U6477 ( .A1(n6266), .A2(n5662), .B1(n6273), .B2(
        PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5238) );
  NAND2_X1 U6478 ( .A1(n6260), .A2(EBX_REG_28__SCAN_IN), .ZN(n5237) );
  OAI211_X1 U6479 ( .C1(n5240), .C2(n5239), .A(n5238), .B(n5237), .ZN(n5241)
         );
  AOI21_X1 U6480 ( .B1(n4197), .B2(n6279), .A(n5241), .ZN(n5242) );
  OAI21_X1 U6481 ( .B1(n5606), .B2(n6282), .A(n5242), .ZN(U2799) );
  INV_X1 U6482 ( .A(n4189), .ZN(n5245) );
  INV_X1 U6483 ( .A(n5673), .ZN(n5609) );
  INV_X1 U6484 ( .A(n5247), .ZN(n5250) );
  AOI22_X1 U6485 ( .A1(n6266), .A2(n5669), .B1(n6273), .B2(
        PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5249) );
  NAND2_X1 U6486 ( .A1(n6260), .A2(EBX_REG_27__SCAN_IN), .ZN(n5248) );
  OAI211_X1 U6487 ( .C1(n5250), .C2(REIP_REG_27__SCAN_IN), .A(n5249), .B(n5248), .ZN(n5251) );
  AOI21_X1 U6488 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5263), .A(n5251), .ZN(n5256) );
  AND2_X1 U6489 ( .A1(n5259), .A2(n5252), .ZN(n5253) );
  NOR2_X1 U6490 ( .A1(n5254), .A2(n5253), .ZN(n5869) );
  NAND2_X1 U6491 ( .A1(n5869), .A2(n6279), .ZN(n5255) );
  OAI211_X1 U6492 ( .C1(n5609), .C2(n6282), .A(n5256), .B(n5255), .ZN(U2800)
         );
  NAND2_X1 U6493 ( .A1(n5275), .A2(n5257), .ZN(n5258) );
  NAND2_X1 U6494 ( .A1(n5259), .A2(n5258), .ZN(n5878) );
  OAI21_X1 U6495 ( .B1(n5260), .B2(n5261), .A(n5244), .ZN(n5612) );
  INV_X1 U6496 ( .A(n5612), .ZN(n5682) );
  NAND2_X1 U6497 ( .A1(n5682), .A2(n6267), .ZN(n5269) );
  OAI22_X1 U6498 ( .A1(n6280), .A2(n5680), .B1(n6251), .B2(n5262), .ZN(n5267)
         );
  INV_X1 U6499 ( .A(n5263), .ZN(n5265) );
  AOI21_X1 U6500 ( .B1(n5277), .B2(REIP_REG_25__SCAN_IN), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5264) );
  NOR2_X1 U6501 ( .A1(n5265), .A2(n5264), .ZN(n5266) );
  AOI211_X1 U6502 ( .C1(n5538), .C2(EBX_REG_26__SCAN_IN), .A(n5267), .B(n5266), 
        .ZN(n5268) );
  OAI211_X1 U6503 ( .C1(n5878), .C2(n5570), .A(n5269), .B(n5268), .ZN(U2801)
         );
  AOI21_X1 U6504 ( .B1(n5271), .B2(n5270), .A(n5260), .ZN(n5691) );
  INV_X1 U6505 ( .A(n5691), .ZN(n5615) );
  NAND2_X1 U6506 ( .A1(n5301), .A2(n5288), .ZN(n5274) );
  INV_X1 U6507 ( .A(n5272), .ZN(n5273) );
  NAND2_X1 U6508 ( .A1(n5274), .A2(n5273), .ZN(n5276) );
  NAND2_X1 U6509 ( .A1(n5276), .A2(n5275), .ZN(n5576) );
  INV_X1 U6510 ( .A(n5576), .ZN(n5885) );
  INV_X1 U6511 ( .A(n5277), .ZN(n5283) );
  NAND2_X1 U6512 ( .A1(n5278), .A2(REIP_REG_25__SCAN_IN), .ZN(n5282) );
  INV_X1 U6513 ( .A(n5688), .ZN(n5279) );
  OAI22_X1 U6514 ( .A1(n6280), .A2(n5279), .B1(n6251), .B2(n6754), .ZN(n5280)
         );
  AOI21_X1 U6515 ( .B1(n5538), .B2(EBX_REG_25__SCAN_IN), .A(n5280), .ZN(n5281)
         );
  OAI211_X1 U6516 ( .C1(REIP_REG_25__SCAN_IN), .C2(n5283), .A(n5282), .B(n5281), .ZN(n5284) );
  AOI21_X1 U6517 ( .B1(n5885), .B2(n6279), .A(n5284), .ZN(n5285) );
  OAI21_X1 U6518 ( .B1(n5615), .B2(n6282), .A(n5285), .ZN(U2802) );
  OAI21_X1 U6519 ( .B1(n5286), .B2(n5287), .A(n5270), .ZN(n5696) );
  XNOR2_X1 U6520 ( .A(n5301), .B(n5288), .ZN(n5577) );
  INV_X1 U6521 ( .A(n5577), .ZN(n5897) );
  OAI22_X1 U6522 ( .A1(n6280), .A2(n5698), .B1(n6251), .B2(n5289), .ZN(n5290)
         );
  AOI21_X1 U6523 ( .B1(n5538), .B2(EBX_REG_24__SCAN_IN), .A(n5290), .ZN(n5292)
         );
  OAI211_X1 U6524 ( .C1(n5305), .C2(n5293), .A(n5292), .B(n5291), .ZN(n5294)
         );
  AOI21_X1 U6525 ( .B1(n5897), .B2(n6279), .A(n5294), .ZN(n5295) );
  OAI21_X1 U6526 ( .B1(n5696), .B2(n6282), .A(n5295), .ZN(U2803) );
  AOI21_X1 U6527 ( .B1(n5298), .B2(n5297), .A(n5286), .ZN(n5707) );
  INV_X1 U6528 ( .A(n5707), .ZN(n5620) );
  AOI21_X1 U6529 ( .B1(n5326), .B2(n5311), .A(n5299), .ZN(n5300) );
  OR2_X1 U6530 ( .A1(n5301), .A2(n5300), .ZN(n5904) );
  INV_X1 U6531 ( .A(n5904), .ZN(n5307) );
  INV_X1 U6532 ( .A(n5328), .ZN(n5316) );
  AOI21_X1 U6533 ( .B1(n5316), .B2(n5314), .A(REIP_REG_23__SCAN_IN), .ZN(n5304) );
  AOI22_X1 U6534 ( .A1(n6266), .A2(n5710), .B1(n6273), .B2(
        PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5303) );
  NAND2_X1 U6535 ( .A1(n6260), .A2(EBX_REG_23__SCAN_IN), .ZN(n5302) );
  OAI211_X1 U6536 ( .C1(n5305), .C2(n5304), .A(n5303), .B(n5302), .ZN(n5306)
         );
  AOI21_X1 U6537 ( .B1(n5307), .B2(n6279), .A(n5306), .ZN(n5308) );
  OAI21_X1 U6538 ( .B1(n5620), .B2(n6282), .A(n5308), .ZN(U2804) );
  OAI21_X1 U6539 ( .B1(n5309), .B2(n5310), .A(n5297), .ZN(n5717) );
  XOR2_X1 U6540 ( .A(n5311), .B(n5326), .Z(n5911) );
  INV_X1 U6541 ( .A(n5720), .ZN(n5312) );
  OAI22_X1 U6542 ( .A1(n6280), .A2(n5312), .B1(n6251), .B2(n5716), .ZN(n5313)
         );
  AOI21_X1 U6543 ( .B1(n5538), .B2(EBX_REG_22__SCAN_IN), .A(n5313), .ZN(n5318)
         );
  INV_X1 U6544 ( .A(n5314), .ZN(n5315) );
  OAI211_X1 U6545 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5316), .B(n5315), .ZN(n5317) );
  OAI211_X1 U6546 ( .C1(n5343), .C2(n5319), .A(n5318), .B(n5317), .ZN(n5320)
         );
  AOI21_X1 U6547 ( .B1(n5911), .B2(n6279), .A(n5320), .ZN(n5321) );
  OAI21_X1 U6548 ( .B1(n5717), .B2(n6282), .A(n5321), .ZN(U2805) );
  XOR2_X1 U6549 ( .A(n5323), .B(n5322), .Z(n5728) );
  AND2_X1 U6550 ( .A1(n2989), .A2(n5324), .ZN(n5325) );
  NOR2_X1 U6551 ( .A1(n5326), .A2(n5325), .ZN(n5918) );
  OAI22_X1 U6552 ( .A1(n6280), .A2(n5726), .B1(n6251), .B2(n5327), .ZN(n5330)
         );
  NOR2_X1 U6553 ( .A1(n5328), .A2(REIP_REG_21__SCAN_IN), .ZN(n5329) );
  AOI211_X1 U6554 ( .C1(EBX_REG_21__SCAN_IN), .C2(n6260), .A(n5330), .B(n5329), 
        .ZN(n5331) );
  OAI21_X1 U6555 ( .B1(n5343), .B2(n5332), .A(n5331), .ZN(n5333) );
  AOI21_X1 U6556 ( .B1(n5918), .B2(n6279), .A(n5333), .ZN(n5334) );
  OAI21_X1 U6557 ( .B1(n5625), .B2(n6282), .A(n5334), .ZN(U2806) );
  OAI21_X1 U6558 ( .B1(n2992), .B2(n5335), .A(n5322), .ZN(n5732) );
  MUX2_X1 U6559 ( .A(n5352), .B(n5350), .S(n5336), .Z(n5338) );
  XNOR2_X1 U6560 ( .A(n5338), .B(n5337), .ZN(n5581) );
  NOR3_X1 U6561 ( .A1(n5530), .A2(n5355), .A3(n5339), .ZN(n5354) );
  AOI21_X1 U6562 ( .B1(n5354), .B2(REIP_REG_19__SCAN_IN), .A(
        REIP_REG_20__SCAN_IN), .ZN(n5344) );
  OAI22_X1 U6563 ( .A1(n6280), .A2(n5734), .B1(n6251), .B2(n5340), .ZN(n5341)
         );
  AOI21_X1 U6564 ( .B1(EBX_REG_20__SCAN_IN), .B2(n6260), .A(n5341), .ZN(n5342)
         );
  OAI21_X1 U6565 ( .B1(n5344), .B2(n5343), .A(n5342), .ZN(n5345) );
  AOI21_X1 U6566 ( .B1(n5581), .B2(n6279), .A(n5345), .ZN(n5346) );
  OAI21_X1 U6567 ( .B1(n5732), .B2(n6282), .A(n5346), .ZN(U2807) );
  XNOR2_X1 U6568 ( .A(n5347), .B(n5348), .ZN(n5741) );
  INV_X1 U6569 ( .A(n5349), .ZN(n5351) );
  MUX2_X1 U6570 ( .A(n5352), .B(n5351), .S(n5350), .Z(n5370) );
  NAND2_X1 U6571 ( .A1(n5379), .A2(n5370), .ZN(n5372) );
  XNOR2_X1 U6572 ( .A(n5372), .B(n5353), .ZN(n5938) );
  INV_X1 U6573 ( .A(n5354), .ZN(n5361) );
  NOR3_X1 U6574 ( .A1(n5530), .A2(n5355), .A3(REIP_REG_18__SCAN_IN), .ZN(n5367) );
  INV_X1 U6575 ( .A(n5386), .ZN(n5375) );
  OAI21_X1 U6576 ( .B1(n5367), .B2(n5375), .A(REIP_REG_19__SCAN_IN), .ZN(n5360) );
  INV_X1 U6577 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5740) );
  NAND2_X1 U6578 ( .A1(n6266), .A2(n5744), .ZN(n5357) );
  OR2_X1 U6579 ( .A1(n5547), .A2(n5356), .ZN(n6249) );
  OAI211_X1 U6580 ( .C1(n6251), .C2(n5740), .A(n5357), .B(n6249), .ZN(n5358)
         );
  AOI21_X1 U6581 ( .B1(n5538), .B2(EBX_REG_19__SCAN_IN), .A(n5358), .ZN(n5359)
         );
  OAI211_X1 U6582 ( .C1(n5361), .C2(REIP_REG_19__SCAN_IN), .A(n5360), .B(n5359), .ZN(n5362) );
  AOI21_X1 U6583 ( .B1(n5938), .B2(n6279), .A(n5362), .ZN(n5363) );
  OAI21_X1 U6584 ( .B1(n5741), .B2(n6282), .A(n5363), .ZN(U2808) );
  INV_X1 U6585 ( .A(n5347), .ZN(n5365) );
  AOI21_X1 U6586 ( .B1(n5366), .B2(n5364), .A(n5365), .ZN(n5752) );
  INV_X1 U6587 ( .A(n5752), .ZN(n5632) );
  AOI21_X1 U6588 ( .B1(n6260), .B2(EBX_REG_18__SCAN_IN), .A(n5367), .ZN(n5369)
         );
  AOI21_X1 U6589 ( .B1(n6266), .B2(n5748), .A(n6272), .ZN(n5368) );
  OAI211_X1 U6590 ( .C1(n5750), .C2(n6251), .A(n5369), .B(n5368), .ZN(n5374)
         );
  OR2_X1 U6591 ( .A1(n5379), .A2(n5370), .ZN(n5371) );
  NAND2_X1 U6592 ( .A1(n5372), .A2(n5371), .ZN(n5950) );
  NOR2_X1 U6593 ( .A1(n5950), .A2(n5570), .ZN(n5373) );
  AOI211_X1 U6594 ( .C1(n5375), .C2(REIP_REG_18__SCAN_IN), .A(n5374), .B(n5373), .ZN(n5376) );
  OAI21_X1 U6595 ( .B1(n5632), .B2(n6282), .A(n5376), .ZN(U2809) );
  XNOR2_X1 U6596 ( .A(n5377), .B(n5378), .ZN(n5759) );
  AOI21_X1 U6597 ( .B1(n5380), .B2(n5399), .A(n5379), .ZN(n5955) );
  INV_X1 U6598 ( .A(n5421), .ZN(n5381) );
  NOR2_X1 U6599 ( .A1(n5530), .A2(n5381), .ZN(n5408) );
  NOR2_X1 U6600 ( .A1(n5382), .A2(n5407), .ZN(n5392) );
  AOI21_X1 U6601 ( .B1(n5408), .B2(n5392), .A(REIP_REG_17__SCAN_IN), .ZN(n5387) );
  AOI21_X1 U6602 ( .B1(n6266), .B2(n5762), .A(n6272), .ZN(n5383) );
  OAI21_X1 U6603 ( .B1(n5758), .B2(n6251), .A(n5383), .ZN(n5384) );
  AOI21_X1 U6604 ( .B1(n6260), .B2(EBX_REG_17__SCAN_IN), .A(n5384), .ZN(n5385)
         );
  OAI21_X1 U6605 ( .B1(n5387), .B2(n5386), .A(n5385), .ZN(n5388) );
  AOI21_X1 U6606 ( .B1(n5955), .B2(n6279), .A(n5388), .ZN(n5389) );
  OAI21_X1 U6607 ( .B1(n5759), .B2(n6282), .A(n5389), .ZN(U2810) );
  OAI21_X1 U6608 ( .B1(n5390), .B2(n5391), .A(n5377), .ZN(n5766) );
  OAI21_X1 U6609 ( .B1(n5530), .B2(n5421), .A(n5504), .ZN(n5429) );
  INV_X1 U6610 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5586) );
  INV_X1 U6611 ( .A(n5392), .ZN(n5393) );
  OAI211_X1 U6612 ( .C1(REIP_REG_16__SCAN_IN), .C2(REIP_REG_15__SCAN_IN), .A(
        n5408), .B(n5393), .ZN(n5396) );
  OAI21_X1 U6613 ( .B1(n6251), .B2(n3071), .A(n6249), .ZN(n5394) );
  AOI21_X1 U6614 ( .B1(n5769), .B2(n6266), .A(n5394), .ZN(n5395) );
  OAI211_X1 U6615 ( .C1(n5586), .C2(n6276), .A(n5396), .B(n5395), .ZN(n5401)
         );
  NAND2_X1 U6616 ( .A1(n5414), .A2(n5397), .ZN(n5398) );
  NAND2_X1 U6617 ( .A1(n5399), .A2(n5398), .ZN(n5966) );
  NOR2_X1 U6618 ( .A1(n5966), .A2(n5570), .ZN(n5400) );
  AOI211_X1 U6619 ( .C1(REIP_REG_16__SCAN_IN), .C2(n5429), .A(n5401), .B(n5400), .ZN(n5402) );
  OAI21_X1 U6620 ( .B1(n5766), .B2(n6282), .A(n5402), .ZN(U2811) );
  AOI21_X1 U6621 ( .B1(n5404), .B2(n5403), .A(n5390), .ZN(n5776) );
  INV_X1 U6622 ( .A(n5776), .ZN(n5640) );
  INV_X1 U6623 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5587) );
  INV_X1 U6624 ( .A(n5405), .ZN(n5774) );
  NOR2_X1 U6625 ( .A1(n6280), .A2(n5774), .ZN(n5406) );
  AOI211_X1 U6626 ( .C1(n6273), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n6272), 
        .B(n5406), .ZN(n5410) );
  NAND2_X1 U6627 ( .A1(n5408), .A2(n5407), .ZN(n5409) );
  OAI211_X1 U6628 ( .C1(n5587), .C2(n6276), .A(n5410), .B(n5409), .ZN(n5416)
         );
  NAND2_X1 U6629 ( .A1(n5411), .A2(n5412), .ZN(n5413) );
  NAND2_X1 U6630 ( .A1(n5414), .A2(n5413), .ZN(n5980) );
  NOR2_X1 U6631 ( .A1(n5980), .A2(n5570), .ZN(n5415) );
  AOI211_X1 U6632 ( .C1(REIP_REG_15__SCAN_IN), .C2(n5429), .A(n5416), .B(n5415), .ZN(n5417) );
  OAI21_X1 U6633 ( .B1(n5640), .B2(n6282), .A(n5417), .ZN(U2812) );
  OAI21_X1 U6634 ( .B1(n5418), .B2(n5419), .A(n5403), .ZN(n5780) );
  NOR3_X1 U6635 ( .A1(n5530), .A2(n5421), .A3(n5420), .ZN(n5422) );
  AOI21_X1 U6636 ( .B1(EBX_REG_14__SCAN_IN), .B2(n6260), .A(n5422), .ZN(n5424)
         );
  AOI21_X1 U6637 ( .B1(n6273), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6272), 
        .ZN(n5423) );
  OAI211_X1 U6638 ( .C1(n5782), .C2(n6280), .A(n5424), .B(n5423), .ZN(n5428)
         );
  OR2_X1 U6639 ( .A1(n5441), .A2(n5425), .ZN(n5426) );
  NAND2_X1 U6640 ( .A1(n5411), .A2(n5426), .ZN(n5991) );
  NOR2_X1 U6641 ( .A1(n5991), .A2(n5570), .ZN(n5427) );
  AOI211_X1 U6642 ( .C1(REIP_REG_14__SCAN_IN), .C2(n5429), .A(n5428), .B(n5427), .ZN(n5430) );
  OAI21_X1 U6643 ( .B1(n5780), .B2(n6282), .A(n5430), .ZN(U2813) );
  NAND2_X1 U6644 ( .A1(n5432), .A2(n5433), .ZN(n5434) );
  OR2_X1 U6645 ( .A1(n5547), .A2(n5435), .ZN(n5471) );
  OAI21_X1 U6646 ( .B1(n5436), .B2(n5471), .A(n5564), .ZN(n5437) );
  INV_X1 U6647 ( .A(n5437), .ZN(n6247) );
  AND3_X1 U6648 ( .A1(n5532), .A2(n5444), .A3(n6798), .ZN(n5451) );
  OAI21_X1 U6649 ( .B1(n6247), .B2(n5451), .A(REIP_REG_13__SCAN_IN), .ZN(n5448) );
  AOI21_X1 U6650 ( .B1(n6032), .B2(n5439), .A(n5438), .ZN(n5440) );
  OR2_X1 U6651 ( .A1(n5441), .A2(n5440), .ZN(n6289) );
  INV_X1 U6652 ( .A(n6289), .ZN(n6005) );
  AOI22_X1 U6653 ( .A1(EBX_REG_13__SCAN_IN), .A2(n5538), .B1(n6279), .B2(n6005), .ZN(n5447) );
  NOR2_X1 U6654 ( .A1(n6280), .A2(n5789), .ZN(n5442) );
  AOI211_X1 U6655 ( .C1(n6273), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6272), 
        .B(n5442), .ZN(n5446) );
  NAND2_X1 U6656 ( .A1(REIP_REG_12__SCAN_IN), .A2(n4370), .ZN(n6721) );
  INV_X1 U6657 ( .A(n6721), .ZN(n5443) );
  NAND3_X1 U6658 ( .A1(n5532), .A2(n5444), .A3(n5443), .ZN(n5445) );
  AND4_X1 U6659 ( .A1(n5448), .A2(n5447), .A3(n5446), .A4(n5445), .ZN(n5449)
         );
  OAI21_X1 U6660 ( .B1(n5644), .B2(n6282), .A(n5449), .ZN(U2814) );
  INV_X1 U6661 ( .A(n6014), .ZN(n5453) );
  INV_X1 U6662 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5799) );
  OAI211_X1 U6663 ( .C1(n6251), .C2(n5799), .A(n5450), .B(n6249), .ZN(n5452)
         );
  INV_X1 U6664 ( .A(n5455), .ZN(n5456) );
  OAI21_X1 U6665 ( .B1(n5456), .B2(n5471), .A(n5564), .ZN(n6287) );
  INV_X1 U6666 ( .A(n5811), .ZN(n5461) );
  INV_X1 U6667 ( .A(n5807), .ZN(n5457) );
  AOI22_X1 U6668 ( .A1(n6266), .A2(n5457), .B1(n6273), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5459) );
  AOI22_X1 U6669 ( .A1(EBX_REG_10__SCAN_IN), .A2(n5538), .B1(n6279), .B2(n6378), .ZN(n5458) );
  NAND3_X1 U6670 ( .A1(n5459), .A2(n5458), .A3(n6249), .ZN(n5460) );
  AOI21_X1 U6671 ( .B1(n5461), .B2(n6267), .A(n5460), .ZN(n5469) );
  INV_X1 U6672 ( .A(n5462), .ZN(n5463) );
  NAND2_X1 U6673 ( .A1(REIP_REG_6__SCAN_IN), .A2(REIP_REG_5__SCAN_IN), .ZN(
        n5464) );
  INV_X1 U6674 ( .A(n6271), .ZN(n5465) );
  NOR2_X1 U6675 ( .A1(n5466), .A2(n5465), .ZN(n6257) );
  NAND2_X1 U6676 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5467) );
  OAI211_X1 U6677 ( .C1(REIP_REG_10__SCAN_IN), .C2(REIP_REG_9__SCAN_IN), .A(
        n6257), .B(n5467), .ZN(n5468) );
  OAI211_X1 U6678 ( .C1(n6287), .C2(n5470), .A(n5469), .B(n5468), .ZN(U2817)
         );
  NAND2_X1 U6679 ( .A1(n5564), .A2(n5471), .ZN(n5490) );
  INV_X1 U6680 ( .A(n5490), .ZN(n5493) );
  INV_X1 U6681 ( .A(n5472), .ZN(n5494) );
  AND3_X1 U6682 ( .A1(n5494), .A2(REIP_REG_5__SCAN_IN), .A3(n6844), .ZN(n5487)
         );
  OAI21_X1 U6683 ( .B1(n5493), .B2(n5487), .A(REIP_REG_7__SCAN_IN), .ZN(n5480)
         );
  INV_X1 U6684 ( .A(n5473), .ZN(n5474) );
  AOI22_X1 U6685 ( .A1(n6266), .A2(n5474), .B1(n6273), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5477) );
  INV_X1 U6686 ( .A(n5475), .ZN(n6395) );
  AOI22_X1 U6687 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6260), .B1(n6279), .B2(n6395), 
        .ZN(n5476) );
  NAND3_X1 U6688 ( .A1(n5477), .A2(n5476), .A3(n6249), .ZN(n5478) );
  AOI21_X1 U6689 ( .B1(n6271), .B2(n4382), .A(n5478), .ZN(n5479) );
  OAI211_X1 U6690 ( .C1(n5481), .C2(n6282), .A(n5480), .B(n5479), .ZN(U2820)
         );
  NOR2_X1 U6691 ( .A1(n6280), .A2(n6353), .ZN(n5482) );
  AOI211_X1 U6692 ( .C1(n6273), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6272), 
        .B(n5482), .ZN(n5484) );
  NAND2_X1 U6693 ( .A1(n6279), .A2(n6065), .ZN(n5483) );
  OAI211_X1 U6694 ( .C1(n5485), .C2(n6276), .A(n5484), .B(n5483), .ZN(n5486)
         );
  AOI211_X1 U6695 ( .C1(n5488), .C2(n6267), .A(n5487), .B(n5486), .ZN(n5489)
         );
  OAI21_X1 U6696 ( .B1(n5490), .B2(n6844), .A(n5489), .ZN(U2821) );
  NOR2_X1 U6697 ( .A1(n5511), .A2(n5491), .ZN(n5492) );
  OR2_X1 U6698 ( .A1(n6267), .A2(n5492), .ZN(n5544) );
  OAI21_X1 U6699 ( .B1(n5494), .B2(REIP_REG_5__SCAN_IN), .A(n5493), .ZN(n5501)
         );
  AOI21_X1 U6700 ( .B1(n6266), .B2(n5495), .A(n6272), .ZN(n5497) );
  NAND2_X1 U6701 ( .A1(n6260), .A2(EBX_REG_5__SCAN_IN), .ZN(n5496) );
  OAI211_X1 U6702 ( .C1(n5498), .C2(n6251), .A(n5497), .B(n5496), .ZN(n5499)
         );
  AOI21_X1 U6703 ( .B1(n6279), .B2(n6404), .A(n5499), .ZN(n5500) );
  OAI211_X1 U6704 ( .C1(n5561), .C2(n5502), .A(n5501), .B(n5500), .ZN(U2822)
         );
  INV_X1 U6705 ( .A(n5512), .ZN(n5503) );
  OR2_X1 U6706 ( .A1(n5530), .A2(n5503), .ZN(n5505) );
  NAND2_X1 U6707 ( .A1(n5505), .A2(n5504), .ZN(n5520) );
  INV_X1 U6708 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5509) );
  INV_X1 U6709 ( .A(n6363), .ZN(n5506) );
  AOI21_X1 U6710 ( .B1(n6266), .B2(n5506), .A(n6272), .ZN(n5508) );
  NAND2_X1 U6711 ( .A1(n5538), .A2(EBX_REG_4__SCAN_IN), .ZN(n5507) );
  OAI211_X1 U6712 ( .C1(n5509), .C2(n6251), .A(n5508), .B(n5507), .ZN(n5518)
         );
  NOR2_X1 U6713 ( .A1(n5511), .A2(n5510), .ZN(n5566) );
  NOR3_X1 U6714 ( .A1(n5530), .A2(REIP_REG_4__SCAN_IN), .A3(n5512), .ZN(n5513)
         );
  AOI21_X1 U6715 ( .B1(n5514), .B2(n5566), .A(n5513), .ZN(n5515) );
  OAI21_X1 U6716 ( .B1(n5570), .B2(n5516), .A(n5515), .ZN(n5517) );
  AOI211_X1 U6717 ( .C1(REIP_REG_4__SCAN_IN), .C2(n5520), .A(n5518), .B(n5517), 
        .ZN(n5519) );
  OAI21_X1 U6718 ( .B1(n5561), .B2(n6359), .A(n5519), .ZN(U2823) );
  NOR3_X1 U6719 ( .A1(n5547), .A2(n5531), .A3(n6815), .ZN(n5521) );
  OAI21_X1 U6720 ( .B1(REIP_REG_3__SCAN_IN), .B2(n5521), .A(n5520), .ZN(n5527)
         );
  OAI22_X1 U6721 ( .A1(n6280), .A2(n5522), .B1(n6251), .B2(n3060), .ZN(n5523)
         );
  AOI21_X1 U6722 ( .B1(n5566), .B2(n6144), .A(n5523), .ZN(n5526) );
  NAND2_X1 U6723 ( .A1(n6279), .A2(n6423), .ZN(n5525) );
  NAND2_X1 U6724 ( .A1(n6260), .A2(EBX_REG_3__SCAN_IN), .ZN(n5524) );
  AND4_X1 U6725 ( .A1(n5527), .A2(n5526), .A3(n5525), .A4(n5524), .ZN(n5528)
         );
  OAI21_X1 U6726 ( .B1(n5529), .B2(n5561), .A(n5528), .ZN(U2824) );
  NOR2_X1 U6727 ( .A1(n5530), .A2(REIP_REG_1__SCAN_IN), .ZN(n5546) );
  NOR3_X1 U6728 ( .A1(n5546), .A2(n5547), .A3(n5531), .ZN(n5534) );
  AOI21_X1 U6729 ( .B1(n5532), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n5533) );
  NOR2_X1 U6730 ( .A1(n5534), .A2(n5533), .ZN(n5543) );
  OAI22_X1 U6731 ( .A1(n6280), .A2(n6374), .B1(n6251), .B2(n5535), .ZN(n5536)
         );
  AOI21_X1 U6732 ( .B1(n5537), .B2(n5566), .A(n5536), .ZN(n5541) );
  NAND2_X1 U6733 ( .A1(n6279), .A2(n6432), .ZN(n5540) );
  NAND2_X1 U6734 ( .A1(n5538), .A2(EBX_REG_2__SCAN_IN), .ZN(n5539) );
  NAND3_X1 U6735 ( .A1(n5541), .A2(n5540), .A3(n5539), .ZN(n5542) );
  AOI211_X1 U6736 ( .C1(n6371), .C2(n5544), .A(n5543), .B(n5542), .ZN(n5545)
         );
  INV_X1 U6737 ( .A(n5545), .ZN(U2825) );
  INV_X1 U6738 ( .A(n5546), .ZN(n5557) );
  NOR2_X1 U6739 ( .A1(n6280), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5551)
         );
  NAND2_X1 U6740 ( .A1(n5547), .A2(REIP_REG_1__SCAN_IN), .ZN(n5548) );
  OAI21_X1 U6741 ( .B1(n6251), .B2(n5549), .A(n5548), .ZN(n5550) );
  NOR2_X1 U6742 ( .A1(n5551), .A2(n5550), .ZN(n5556) );
  INV_X1 U6743 ( .A(n4526), .ZN(n5552) );
  AOI22_X1 U6744 ( .A1(n4505), .A2(n5566), .B1(n5553), .B2(n5552), .ZN(n5555)
         );
  NAND2_X1 U6745 ( .A1(n6260), .A2(EBX_REG_1__SCAN_IN), .ZN(n5554) );
  AND4_X1 U6746 ( .A1(n5557), .A2(n5556), .A3(n5555), .A4(n5554), .ZN(n5558)
         );
  OAI21_X1 U6747 ( .B1(n5561), .B2(n5559), .A(n5558), .ZN(U2826) );
  OAI22_X1 U6748 ( .A1(n5562), .A2(n6276), .B1(n5561), .B2(n5560), .ZN(n5563)
         );
  AOI21_X1 U6749 ( .B1(REIP_REG_0__SCAN_IN), .B2(n5564), .A(n5563), .ZN(n5568)
         );
  NAND2_X1 U6750 ( .A1(n6280), .A2(n6251), .ZN(n5565) );
  AOI22_X1 U6751 ( .A1(n5566), .A2(n6552), .B1(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n5565), .ZN(n5567) );
  OAI211_X1 U6752 ( .C1(n5570), .C2(n5569), .A(n5568), .B(n5567), .ZN(U2827)
         );
  INV_X1 U6753 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5571) );
  OAI22_X1 U6754 ( .A1(n5572), .A2(n6295), .B1(n5571), .B2(n6302), .ZN(U2828)
         );
  AOI22_X1 U6755 ( .A1(n3138), .A2(n4196), .B1(n5584), .B2(EBX_REG_29__SCAN_IN), .ZN(n5573) );
  OAI21_X1 U6756 ( .B1(n5603), .B2(n5588), .A(n5573), .ZN(U2830) );
  AOI22_X1 U6757 ( .A1(n5869), .A2(n4196), .B1(n5584), .B2(EBX_REG_27__SCAN_IN), .ZN(n5574) );
  OAI21_X1 U6758 ( .B1(n5609), .B2(n5588), .A(n5574), .ZN(U2832) );
  INV_X1 U6759 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6831) );
  OAI222_X1 U6760 ( .A1(n5878), .A2(n6295), .B1(n6831), .B2(n6302), .C1(n5612), 
        .C2(n5588), .ZN(U2833) );
  OAI222_X1 U6761 ( .A1(n5576), .A2(n6295), .B1(n5575), .B2(n6302), .C1(n5615), 
        .C2(n5588), .ZN(U2834) );
  INV_X1 U6762 ( .A(EBX_REG_24__SCAN_IN), .ZN(n6768) );
  OAI222_X1 U6763 ( .A1(n6768), .A2(n6302), .B1(n6295), .B2(n5577), .C1(n5588), 
        .C2(n5696), .ZN(U2835) );
  OAI222_X1 U6764 ( .A1(n5578), .A2(n6302), .B1(n6295), .B2(n5904), .C1(n5620), 
        .C2(n5588), .ZN(U2836) );
  AOI22_X1 U6765 ( .A1(n5911), .A2(n4196), .B1(EBX_REG_22__SCAN_IN), .B2(n5584), .ZN(n5579) );
  OAI21_X1 U6766 ( .B1(n5717), .B2(n5588), .A(n5579), .ZN(U2837) );
  AOI22_X1 U6767 ( .A1(n5918), .A2(n4196), .B1(n5584), .B2(EBX_REG_21__SCAN_IN), .ZN(n5580) );
  OAI21_X1 U6768 ( .B1(n5625), .B2(n5588), .A(n5580), .ZN(U2838) );
  INV_X1 U6769 ( .A(n5581), .ZN(n5934) );
  OAI222_X1 U6770 ( .A1(n5732), .A2(n5588), .B1(n6302), .B2(n6818), .C1(n5934), 
        .C2(n6295), .ZN(U2839) );
  INV_X1 U6771 ( .A(n5938), .ZN(n5582) );
  INV_X1 U6772 ( .A(EBX_REG_19__SCAN_IN), .ZN(n6778) );
  OAI222_X1 U6773 ( .A1(n5741), .A2(n5588), .B1(n6295), .B2(n5582), .C1(n6302), 
        .C2(n6778), .ZN(U2840) );
  OAI222_X1 U6774 ( .A1(n5950), .A2(n6295), .B1(n5583), .B2(n6302), .C1(n5632), 
        .C2(n5588), .ZN(U2841) );
  AOI22_X1 U6775 ( .A1(n5955), .A2(n4196), .B1(n5584), .B2(EBX_REG_17__SCAN_IN), .ZN(n5585) );
  OAI21_X1 U6776 ( .B1(n5759), .B2(n5588), .A(n5585), .ZN(U2842) );
  OAI222_X1 U6777 ( .A1(n5966), .A2(n6295), .B1(n5586), .B2(n6302), .C1(n5766), 
        .C2(n5588), .ZN(U2843) );
  OAI222_X1 U6778 ( .A1(n5980), .A2(n6295), .B1(n5587), .B2(n6302), .C1(n5640), 
        .C2(n5588), .ZN(U2844) );
  INV_X1 U6779 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5589) );
  OAI222_X1 U6780 ( .A1(n5991), .A2(n6295), .B1(n5589), .B2(n6302), .C1(n5780), 
        .C2(n5588), .ZN(U2845) );
  NOR3_X1 U6781 ( .A1(n5590), .A2(n5641), .A3(n5592), .ZN(n5600) );
  NAND4_X1 U6782 ( .A1(n5590), .A2(n5593), .A3(n5592), .A4(n5645), .ZN(n5597)
         );
  OAI211_X1 U6783 ( .C1(n5593), .C2(n5592), .A(n5645), .B(n5591), .ZN(n5594)
         );
  OAI21_X1 U6784 ( .B1(n5645), .B2(n5595), .A(n5594), .ZN(n5596) );
  NAND2_X1 U6785 ( .A1(n5597), .A2(n5596), .ZN(n5599) );
  INV_X1 U6786 ( .A(n5636), .ZN(n5598) );
  OAI22_X1 U6787 ( .A1(n5600), .A2(n5599), .B1(n5598), .B2(n6784), .ZN(U2860)
         );
  AOI22_X1 U6788 ( .A1(n5635), .A2(DATAI_13_), .B1(n5641), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U6789 ( .A1(n5636), .A2(DATAI_29_), .ZN(n5601) );
  OAI211_X1 U6790 ( .C1(n5603), .C2(n4987), .A(n5602), .B(n5601), .ZN(U2862)
         );
  AOI22_X1 U6791 ( .A1(n5635), .A2(DATAI_12_), .B1(n5641), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U6792 ( .A1(n5636), .A2(DATAI_28_), .ZN(n5604) );
  OAI211_X1 U6793 ( .C1(n5606), .C2(n4987), .A(n5605), .B(n5604), .ZN(U2863)
         );
  AOI22_X1 U6794 ( .A1(n5635), .A2(DATAI_11_), .B1(n5641), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U6795 ( .A1(n5636), .A2(DATAI_27_), .ZN(n5607) );
  OAI211_X1 U6796 ( .C1(n5609), .C2(n4987), .A(n5608), .B(n5607), .ZN(U2864)
         );
  AOI22_X1 U6797 ( .A1(n5635), .A2(DATAI_10_), .B1(n5641), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5611) );
  NAND2_X1 U6798 ( .A1(n5636), .A2(DATAI_26_), .ZN(n5610) );
  OAI211_X1 U6799 ( .C1(n5612), .C2(n4987), .A(n5611), .B(n5610), .ZN(U2865)
         );
  AOI22_X1 U6800 ( .A1(n5635), .A2(DATAI_9_), .B1(n5641), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U6801 ( .A1(n5636), .A2(DATAI_25_), .ZN(n5613) );
  OAI211_X1 U6802 ( .C1(n5615), .C2(n4987), .A(n5614), .B(n5613), .ZN(U2866)
         );
  AOI22_X1 U6803 ( .A1(n5635), .A2(DATAI_8_), .B1(n5641), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5617) );
  NAND2_X1 U6804 ( .A1(n5636), .A2(DATAI_24_), .ZN(n5616) );
  OAI211_X1 U6805 ( .C1(n5696), .C2(n4987), .A(n5617), .B(n5616), .ZN(U2867)
         );
  AOI22_X1 U6806 ( .A1(n5635), .A2(DATAI_7_), .B1(n5641), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U6807 ( .A1(n5636), .A2(DATAI_23_), .ZN(n5618) );
  OAI211_X1 U6808 ( .C1(n5620), .C2(n4987), .A(n5619), .B(n5618), .ZN(U2868)
         );
  AOI22_X1 U6809 ( .A1(n5635), .A2(DATAI_6_), .B1(n5641), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U6810 ( .A1(n5636), .A2(DATAI_22_), .ZN(n5621) );
  OAI211_X1 U6811 ( .C1(n5717), .C2(n4987), .A(n5622), .B(n5621), .ZN(U2869)
         );
  AOI22_X1 U6812 ( .A1(n5635), .A2(DATAI_5_), .B1(n5641), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5624) );
  NAND2_X1 U6813 ( .A1(n5636), .A2(DATAI_21_), .ZN(n5623) );
  OAI211_X1 U6814 ( .C1(n5625), .C2(n4987), .A(n5624), .B(n5623), .ZN(U2870)
         );
  AOI22_X1 U6815 ( .A1(n5635), .A2(DATAI_4_), .B1(n5641), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U6816 ( .A1(n5636), .A2(DATAI_20_), .ZN(n5626) );
  OAI211_X1 U6817 ( .C1(n5732), .C2(n4987), .A(n5627), .B(n5626), .ZN(U2871)
         );
  AOI22_X1 U6818 ( .A1(n5635), .A2(DATAI_3_), .B1(n5641), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U6819 ( .A1(n5636), .A2(DATAI_19_), .ZN(n5628) );
  OAI211_X1 U6820 ( .C1(n5741), .C2(n4987), .A(n5629), .B(n5628), .ZN(U2872)
         );
  AOI22_X1 U6821 ( .A1(n5635), .A2(DATAI_2_), .B1(n5641), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5631) );
  NAND2_X1 U6822 ( .A1(n5636), .A2(DATAI_18_), .ZN(n5630) );
  OAI211_X1 U6823 ( .C1(n5632), .C2(n4987), .A(n5631), .B(n5630), .ZN(U2873)
         );
  AOI22_X1 U6824 ( .A1(n5635), .A2(DATAI_1_), .B1(n5641), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U6825 ( .A1(n5636), .A2(DATAI_17_), .ZN(n5633) );
  OAI211_X1 U6826 ( .C1(n5759), .C2(n4987), .A(n5634), .B(n5633), .ZN(U2874)
         );
  AOI22_X1 U6827 ( .A1(n5635), .A2(DATAI_0_), .B1(n5641), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U6828 ( .A1(n5636), .A2(DATAI_16_), .ZN(n5637) );
  OAI211_X1 U6829 ( .C1(n5766), .C2(n4987), .A(n5638), .B(n5637), .ZN(U2875)
         );
  AOI22_X1 U6830 ( .A1(n5642), .A2(DATAI_15_), .B1(n5641), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5639) );
  OAI21_X1 U6831 ( .B1(n5640), .B2(n4987), .A(n5639), .ZN(U2876) );
  AOI22_X1 U6832 ( .A1(n5642), .A2(DATAI_14_), .B1(n5641), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5643) );
  OAI21_X1 U6833 ( .B1(n5780), .B2(n4987), .A(n5643), .ZN(U2877) );
  INV_X1 U6834 ( .A(DATAI_13_), .ZN(n5646) );
  OAI222_X1 U6835 ( .A1(n5647), .A2(n5646), .B1(n5645), .B2(n6804), .C1(n4987), 
        .C2(n5644), .ZN(U2878) );
  INV_X1 U6836 ( .A(n5648), .ZN(n5861) );
  INV_X1 U6837 ( .A(n5649), .ZN(n5678) );
  XNOR2_X1 U6838 ( .A(n5651), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5859)
         );
  NAND2_X1 U6839 ( .A1(n5818), .A2(n5652), .ZN(n5653) );
  NAND2_X1 U6840 ( .A1(n6364), .A2(REIP_REG_29__SCAN_IN), .ZN(n5854) );
  OAI211_X1 U6841 ( .C1(n5816), .C2(n5654), .A(n5653), .B(n5854), .ZN(n5655)
         );
  AOI21_X1 U6842 ( .B1(n5656), .B2(n6370), .A(n5655), .ZN(n5657) );
  OAI21_X1 U6843 ( .B1(n5859), .B2(n6345), .A(n5657), .ZN(U2957) );
  INV_X1 U6844 ( .A(n5658), .ZN(n5660) );
  XNOR2_X1 U6845 ( .A(n5661), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5868)
         );
  NAND2_X1 U6846 ( .A1(n5818), .A2(n5662), .ZN(n5663) );
  NAND2_X1 U6847 ( .A1(n6364), .A2(REIP_REG_28__SCAN_IN), .ZN(n5863) );
  OAI211_X1 U6848 ( .C1(n5816), .C2(n3074), .A(n5663), .B(n5863), .ZN(n5664)
         );
  AOI21_X1 U6849 ( .B1(n5665), .B2(n6370), .A(n5664), .ZN(n5666) );
  OAI21_X1 U6850 ( .B1(n6345), .B2(n5868), .A(n5666), .ZN(U2958) );
  OAI21_X1 U6851 ( .B1(n5684), .B2(n5676), .A(n5667), .ZN(n5668) );
  XNOR2_X1 U6852 ( .A(n5668), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5876)
         );
  NAND2_X1 U6853 ( .A1(n5818), .A2(n5669), .ZN(n5670) );
  NAND2_X1 U6854 ( .A1(n6364), .A2(REIP_REG_27__SCAN_IN), .ZN(n5870) );
  OAI211_X1 U6855 ( .C1(n5816), .C2(n5671), .A(n5670), .B(n5870), .ZN(n5672)
         );
  AOI21_X1 U6856 ( .B1(n5673), .B2(n6370), .A(n5672), .ZN(n5674) );
  OAI21_X1 U6857 ( .B1(n5876), .B2(n6345), .A(n5674), .ZN(U2959) );
  NAND2_X1 U6858 ( .A1(n5676), .A2(n5675), .ZN(n5677) );
  XNOR2_X1 U6859 ( .A(n5678), .B(n5677), .ZN(n5884) );
  NAND2_X1 U6860 ( .A1(n6364), .A2(REIP_REG_26__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U6861 ( .A1(n6365), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5679)
         );
  OAI211_X1 U6862 ( .C1(n6375), .C2(n5680), .A(n5877), .B(n5679), .ZN(n5681)
         );
  AOI21_X1 U6863 ( .B1(n5682), .B2(n6370), .A(n5681), .ZN(n5683) );
  OAI21_X1 U6864 ( .B1(n5884), .B2(n6345), .A(n5683), .ZN(U2960) );
  INV_X1 U6865 ( .A(n5684), .ZN(n5685) );
  AOI21_X1 U6866 ( .B1(n5687), .B2(n5686), .A(n5685), .ZN(n5892) );
  NAND2_X1 U6867 ( .A1(n5818), .A2(n5688), .ZN(n5689) );
  NAND2_X1 U6868 ( .A1(n6364), .A2(REIP_REG_25__SCAN_IN), .ZN(n5886) );
  OAI211_X1 U6869 ( .C1(n5816), .C2(n6754), .A(n5689), .B(n5886), .ZN(n5690)
         );
  AOI21_X1 U6870 ( .B1(n5691), .B2(n6370), .A(n5690), .ZN(n5692) );
  OAI21_X1 U6871 ( .B1(n5892), .B2(n6345), .A(n5692), .ZN(U2961) );
  XNOR2_X1 U6872 ( .A(n6026), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5738)
         );
  XNOR2_X1 U6873 ( .A(n6026), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5731)
         );
  INV_X1 U6874 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6795) );
  XNOR2_X1 U6875 ( .A(n2964), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5723)
         );
  NOR2_X1 U6876 ( .A1(n6026), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5713)
         );
  NAND2_X1 U6877 ( .A1(n5722), .A2(n5713), .ZN(n5705) );
  OAI21_X1 U6878 ( .B1(n2964), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5693), 
        .ZN(n5715) );
  NAND3_X1 U6879 ( .A1(n4329), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5694) );
  OAI22_X1 U6880 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n5705), .B1(n5715), .B2(n5694), .ZN(n5695) );
  XNOR2_X1 U6881 ( .A(n5695), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5899)
         );
  INV_X1 U6882 ( .A(n5696), .ZN(n5700) );
  NAND2_X1 U6883 ( .A1(n6364), .A2(REIP_REG_24__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U6884 ( .A1(n6365), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5697)
         );
  OAI211_X1 U6885 ( .C1(n6375), .C2(n5698), .A(n5893), .B(n5697), .ZN(n5699)
         );
  AOI21_X1 U6886 ( .B1(n5700), .B2(n6370), .A(n5699), .ZN(n5701) );
  OAI21_X1 U6887 ( .B1(n5899), .B2(n6345), .A(n5701), .ZN(U2962) );
  OR3_X1 U6888 ( .A1(n5703), .A2(n2964), .A3(n5702), .ZN(n5704) );
  NAND2_X1 U6889 ( .A1(n5705), .A2(n5704), .ZN(n5706) );
  XNOR2_X1 U6890 ( .A(n5706), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5908)
         );
  NAND2_X1 U6891 ( .A1(n5707), .A2(n6370), .ZN(n5712) );
  NAND2_X1 U6892 ( .A1(n6364), .A2(REIP_REG_23__SCAN_IN), .ZN(n5902) );
  OAI21_X1 U6893 ( .B1(n5816), .B2(n5708), .A(n5902), .ZN(n5709) );
  AOI21_X1 U6894 ( .B1(n5818), .B2(n5710), .A(n5709), .ZN(n5711) );
  OAI211_X1 U6895 ( .C1(n5908), .C2(n6345), .A(n5712), .B(n5711), .ZN(U2963)
         );
  AOI21_X1 U6896 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n4329), .A(n5713), 
        .ZN(n5714) );
  XNOR2_X1 U6897 ( .A(n5715), .B(n5714), .ZN(n5917) );
  NAND2_X1 U6898 ( .A1(n6364), .A2(REIP_REG_22__SCAN_IN), .ZN(n5912) );
  OAI21_X1 U6899 ( .B1(n5816), .B2(n5716), .A(n5912), .ZN(n5719) );
  NOR2_X1 U6900 ( .A1(n5717), .A2(n6358), .ZN(n5718) );
  AOI211_X1 U6901 ( .C1(n5818), .C2(n5720), .A(n5719), .B(n5718), .ZN(n5721)
         );
  OAI21_X1 U6902 ( .B1(n5917), .B2(n6345), .A(n5721), .ZN(U2964) );
  AOI21_X1 U6903 ( .B1(n5724), .B2(n5723), .A(n5722), .ZN(n5925) );
  NAND2_X1 U6904 ( .A1(n6364), .A2(REIP_REG_21__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U6905 ( .A1(n6365), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5725)
         );
  OAI211_X1 U6906 ( .C1(n6375), .C2(n5726), .A(n5919), .B(n5725), .ZN(n5727)
         );
  AOI21_X1 U6907 ( .B1(n5728), .B2(n6370), .A(n5727), .ZN(n5729) );
  OAI21_X1 U6908 ( .B1(n5925), .B2(n6345), .A(n5729), .ZN(U2965) );
  XOR2_X1 U6909 ( .A(n5731), .B(n5730), .Z(n5937) );
  INV_X1 U6910 ( .A(n5732), .ZN(n5736) );
  NAND2_X1 U6911 ( .A1(n6364), .A2(REIP_REG_20__SCAN_IN), .ZN(n5933) );
  NAND2_X1 U6912 ( .A1(n6365), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5733)
         );
  OAI211_X1 U6913 ( .C1(n6375), .C2(n5734), .A(n5933), .B(n5733), .ZN(n5735)
         );
  AOI21_X1 U6914 ( .B1(n5736), .B2(n6370), .A(n5735), .ZN(n5737) );
  OAI21_X1 U6915 ( .B1(n5937), .B2(n6345), .A(n5737), .ZN(U2966) );
  XNOR2_X1 U6916 ( .A(n5739), .B(n5738), .ZN(n5945) );
  NAND2_X1 U6917 ( .A1(n6364), .A2(REIP_REG_19__SCAN_IN), .ZN(n5939) );
  OAI21_X1 U6918 ( .B1(n5816), .B2(n5740), .A(n5939), .ZN(n5743) );
  NOR2_X1 U6919 ( .A1(n5741), .A2(n6358), .ZN(n5742) );
  AOI211_X1 U6920 ( .C1(n5818), .C2(n5744), .A(n5743), .B(n5742), .ZN(n5745)
         );
  OAI21_X1 U6921 ( .B1(n5945), .B2(n6345), .A(n5745), .ZN(U2967) );
  NAND3_X1 U6922 ( .A1(n5765), .A2(n2964), .A3(n5973), .ZN(n5754) );
  NOR3_X1 U6923 ( .A1(n5765), .A2(n2964), .A3(n5973), .ZN(n5756) );
  NAND2_X1 U6924 ( .A1(n5756), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5746) );
  OAI21_X1 U6925 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5754), .A(n5746), 
        .ZN(n5747) );
  XNOR2_X1 U6926 ( .A(n5747), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5954)
         );
  NAND2_X1 U6927 ( .A1(n5818), .A2(n5748), .ZN(n5749) );
  NAND2_X1 U6928 ( .A1(n6364), .A2(REIP_REG_18__SCAN_IN), .ZN(n5948) );
  OAI211_X1 U6929 ( .C1(n5816), .C2(n5750), .A(n5749), .B(n5948), .ZN(n5751)
         );
  AOI21_X1 U6930 ( .B1(n5752), .B2(n6370), .A(n5751), .ZN(n5753) );
  OAI21_X1 U6931 ( .B1(n5954), .B2(n6345), .A(n5753), .ZN(U2968) );
  INV_X1 U6932 ( .A(n5754), .ZN(n5755) );
  NOR2_X1 U6933 ( .A1(n5756), .A2(n5755), .ZN(n5757) );
  XNOR2_X1 U6934 ( .A(n5757), .B(n5956), .ZN(n5964) );
  NAND2_X1 U6935 ( .A1(n6364), .A2(REIP_REG_17__SCAN_IN), .ZN(n5958) );
  OAI21_X1 U6936 ( .B1(n5816), .B2(n5758), .A(n5958), .ZN(n5761) );
  NOR2_X1 U6937 ( .A1(n5759), .A2(n6358), .ZN(n5760) );
  AOI211_X1 U6938 ( .C1(n5818), .C2(n5762), .A(n5761), .B(n5760), .ZN(n5763)
         );
  OAI21_X1 U6939 ( .B1(n5964), .B2(n6345), .A(n5763), .ZN(U2969) );
  XNOR2_X1 U6940 ( .A(n6026), .B(n5973), .ZN(n5764) );
  XNOR2_X1 U6941 ( .A(n5765), .B(n5764), .ZN(n5978) );
  NAND2_X1 U6942 ( .A1(n6364), .A2(REIP_REG_16__SCAN_IN), .ZN(n5965) );
  OAI21_X1 U6943 ( .B1(n5816), .B2(n3071), .A(n5965), .ZN(n5768) );
  NOR2_X1 U6944 ( .A1(n5766), .A2(n6358), .ZN(n5767) );
  AOI211_X1 U6945 ( .C1(n5818), .C2(n5769), .A(n5768), .B(n5767), .ZN(n5770)
         );
  OAI21_X1 U6946 ( .B1(n6345), .B2(n5978), .A(n5770), .ZN(U2970) );
  XNOR2_X1 U6947 ( .A(n6026), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5771)
         );
  XNOR2_X1 U6948 ( .A(n5772), .B(n5771), .ZN(n5987) );
  NAND2_X1 U6949 ( .A1(n6364), .A2(REIP_REG_15__SCAN_IN), .ZN(n5979) );
  NAND2_X1 U6950 ( .A1(n6365), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5773)
         );
  OAI211_X1 U6951 ( .C1(n6375), .C2(n5774), .A(n5979), .B(n5773), .ZN(n5775)
         );
  AOI21_X1 U6952 ( .B1(n5776), .B2(n6370), .A(n5775), .ZN(n5777) );
  OAI21_X1 U6953 ( .B1(n5987), .B2(n6345), .A(n5777), .ZN(U2971) );
  XNOR2_X1 U6954 ( .A(n6026), .B(n5988), .ZN(n5778) );
  XNOR2_X1 U6955 ( .A(n5779), .B(n5778), .ZN(n6004) );
  INV_X1 U6956 ( .A(n5780), .ZN(n5784) );
  NAND2_X1 U6957 ( .A1(n6364), .A2(REIP_REG_14__SCAN_IN), .ZN(n5989) );
  NAND2_X1 U6958 ( .A1(n6365), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5781)
         );
  OAI211_X1 U6959 ( .C1(n6375), .C2(n5782), .A(n5989), .B(n5781), .ZN(n5783)
         );
  AOI21_X1 U6960 ( .B1(n5784), .B2(n6370), .A(n5783), .ZN(n5785) );
  OAI21_X1 U6961 ( .B1(n6345), .B2(n6004), .A(n5785), .ZN(U2972) );
  XOR2_X1 U6962 ( .A(n5787), .B(n5786), .Z(n6012) );
  NAND2_X1 U6963 ( .A1(n6364), .A2(REIP_REG_13__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U6964 ( .A1(n6365), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5788)
         );
  OAI211_X1 U6965 ( .C1(n6375), .C2(n5789), .A(n6006), .B(n5788), .ZN(n5790)
         );
  AOI21_X1 U6966 ( .B1(n6291), .B2(n6370), .A(n5790), .ZN(n5791) );
  OAI21_X1 U6967 ( .B1(n6345), .B2(n6012), .A(n5791), .ZN(U2973) );
  OAI21_X1 U6968 ( .B1(n6026), .B2(n6018), .A(n5792), .ZN(n5798) );
  INV_X1 U6969 ( .A(n5793), .ZN(n5796) );
  NAND2_X1 U6970 ( .A1(n5796), .A2(n5805), .ZN(n6025) );
  OAI21_X1 U6971 ( .B1(n6025), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n2964), 
        .ZN(n5794) );
  OAI21_X1 U6972 ( .B1(n5796), .B2(n5795), .A(n5794), .ZN(n5797) );
  XOR2_X1 U6973 ( .A(n5798), .B(n5797), .Z(n6024) );
  AND2_X1 U6974 ( .A1(n6364), .A2(REIP_REG_12__SCAN_IN), .ZN(n6013) );
  NOR2_X1 U6975 ( .A1(n5816), .A2(n5799), .ZN(n5800) );
  AOI211_X1 U6976 ( .C1(n5818), .C2(n5801), .A(n6013), .B(n5800), .ZN(n5804)
         );
  NAND2_X1 U6977 ( .A1(n5802), .A2(n6370), .ZN(n5803) );
  OAI211_X1 U6978 ( .C1(n6024), .C2(n6345), .A(n5804), .B(n5803), .ZN(U2974)
         );
  XNOR2_X1 U6979 ( .A(n6026), .B(n5805), .ZN(n5806) );
  XNOR2_X1 U6980 ( .A(n5793), .B(n5806), .ZN(n6382) );
  NAND2_X1 U6981 ( .A1(n6382), .A2(n6369), .ZN(n5810) );
  NOR2_X1 U6982 ( .A1(n6412), .A2(n5470), .ZN(n6377) );
  NOR2_X1 U6983 ( .A1(n6375), .A2(n5807), .ZN(n5808) );
  AOI211_X1 U6984 ( .C1(n6365), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6377), 
        .B(n5808), .ZN(n5809) );
  OAI211_X1 U6985 ( .C1(n6358), .C2(n5811), .A(n5810), .B(n5809), .ZN(U2976)
         );
  NAND2_X1 U6986 ( .A1(n5813), .A2(n5812), .ZN(n5814) );
  XNOR2_X1 U6987 ( .A(n5815), .B(n5814), .ZN(n6389) );
  NAND2_X1 U6988 ( .A1(n6389), .A2(n6369), .ZN(n5820) );
  NAND2_X1 U6989 ( .A1(n6364), .A2(REIP_REG_9__SCAN_IN), .ZN(n6386) );
  OAI21_X1 U6990 ( .B1(n5816), .B2(n3591), .A(n6386), .ZN(n5817) );
  AOI21_X1 U6991 ( .B1(n5818), .B2(n6265), .A(n5817), .ZN(n5819) );
  OAI211_X1 U6992 ( .C1(n6358), .C2(n6264), .A(n5820), .B(n5819), .ZN(U2977)
         );
  INV_X1 U6993 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5845) );
  NOR2_X1 U6994 ( .A1(n6429), .A2(n6420), .ZN(n6410) );
  NAND2_X1 U6995 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6410), .ZN(n6061)
         );
  NOR2_X1 U6996 ( .A1(n6062), .A2(n6061), .ZN(n5824) );
  AOI21_X1 U6997 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6436) );
  INV_X1 U6998 ( .A(n6042), .ZN(n5822) );
  NOR2_X1 U6999 ( .A1(n6400), .A2(n6046), .ZN(n6379) );
  NAND3_X1 U7000 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6379), .ZN(n5825) );
  INV_X1 U7001 ( .A(n5825), .ZN(n5821) );
  NAND2_X1 U7002 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5993) );
  NOR2_X1 U7003 ( .A1(n5993), .A2(n5998), .ZN(n5995) );
  NAND2_X1 U7004 ( .A1(n5995), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5971) );
  OR3_X1 U7005 ( .A1(n5971), .A2(n5973), .A3(n5984), .ZN(n5926) );
  INV_X1 U7006 ( .A(n6045), .ZN(n6056) );
  NOR2_X1 U7007 ( .A1(n6440), .A2(n6800), .ZN(n6435) );
  NAND2_X1 U7008 ( .A1(n6435), .A2(n5824), .ZN(n6044) );
  NOR2_X1 U7009 ( .A1(n6044), .A2(n5825), .ZN(n5967) );
  INV_X1 U7010 ( .A(n5926), .ZN(n5957) );
  NAND2_X1 U7011 ( .A1(n5967), .A2(n5957), .ZN(n5826) );
  NAND2_X1 U7012 ( .A1(n6045), .A2(n5826), .ZN(n5927) );
  NAND2_X1 U7013 ( .A1(n5827), .A2(n5927), .ZN(n5923) );
  INV_X1 U7014 ( .A(n5910), .ZN(n5835) );
  OAI21_X1 U7015 ( .B1(n6441), .B2(n6434), .A(n5836), .ZN(n5829) );
  INV_X1 U7016 ( .A(n5829), .ZN(n5830) );
  OAI21_X1 U7017 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n6380), .A(n5853), 
        .ZN(n5850) );
  AOI21_X1 U7018 ( .B1(n5845), .B2(n5972), .A(n5850), .ZN(n5840) );
  NAND2_X1 U7019 ( .A1(n6441), .A2(n5967), .ZN(n6017) );
  NAND2_X1 U7020 ( .A1(n6000), .A2(n6017), .ZN(n6037) );
  INV_X1 U7021 ( .A(n5831), .ZN(n5832) );
  NOR2_X1 U7022 ( .A1(n5926), .A2(n5832), .ZN(n5833) );
  NAND2_X1 U7023 ( .A1(n6037), .A2(n5833), .ZN(n5941) );
  INV_X1 U7024 ( .A(n5931), .ZN(n5834) );
  NOR2_X1 U7025 ( .A1(n5921), .A2(n5835), .ZN(n5901) );
  INV_X1 U7026 ( .A(n5836), .ZN(n5837) );
  NAND2_X1 U7027 ( .A1(n5901), .A2(n5837), .ZN(n5888) );
  NOR2_X1 U7028 ( .A1(n5872), .A2(n5861), .ZN(n5857) );
  NAND4_X1 U7029 ( .A1(n5857), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A4(n4515), .ZN(n5838) );
  OAI211_X1 U7030 ( .C1(n5840), .C2(n4515), .A(n5839), .B(n5838), .ZN(n5841)
         );
  AOI21_X1 U7031 ( .B1(n5842), .B2(n6433), .A(n5841), .ZN(n5843) );
  OAI21_X1 U7032 ( .B1(n5844), .B2(n6381), .A(n5843), .ZN(U2987) );
  NAND3_X1 U7033 ( .A1(n5857), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5845), .ZN(n5846) );
  OAI211_X1 U7034 ( .C1(n5848), .C2(n6034), .A(n5847), .B(n5846), .ZN(n5849)
         );
  AOI21_X1 U7035 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5850), .A(n5849), 
        .ZN(n5851) );
  OAI21_X1 U7036 ( .B1(n5852), .B2(n6381), .A(n5851), .ZN(U2988) );
  NOR2_X1 U7037 ( .A1(n5853), .A2(n5856), .ZN(n5855) );
  OAI21_X1 U7038 ( .B1(n5859), .B2(n6381), .A(n5858), .ZN(U2989) );
  INV_X1 U7039 ( .A(n5872), .ZN(n5862) );
  NAND3_X1 U7040 ( .A1(n5862), .A2(n5861), .A3(n5860), .ZN(n5864) );
  OAI211_X1 U7041 ( .C1(n6034), .C2(n5865), .A(n5864), .B(n5863), .ZN(n5866)
         );
  AOI21_X1 U7042 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n5874), .A(n5866), 
        .ZN(n5867) );
  OAI21_X1 U7043 ( .B1(n5868), .B2(n6381), .A(n5867), .ZN(U2990) );
  NAND2_X1 U7044 ( .A1(n5869), .A2(n6433), .ZN(n5871) );
  OAI211_X1 U7045 ( .C1(n5872), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5871), .B(n5870), .ZN(n5873) );
  AOI21_X1 U7046 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5874), .A(n5873), 
        .ZN(n5875) );
  OAI21_X1 U7047 ( .B1(n5876), .B2(n6381), .A(n5875), .ZN(U2991) );
  INV_X1 U7048 ( .A(n2976), .ZN(n5890) );
  OAI21_X1 U7049 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A(n3004), .ZN(n5881) );
  OAI21_X1 U7050 ( .B1(n5878), .B2(n6034), .A(n5877), .ZN(n5879) );
  INV_X1 U7051 ( .A(n5879), .ZN(n5880) );
  OAI21_X1 U7052 ( .B1(n5888), .B2(n5881), .A(n5880), .ZN(n5882) );
  AOI21_X1 U7053 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5890), .A(n5882), 
        .ZN(n5883) );
  OAI21_X1 U7054 ( .B1(n5884), .B2(n6381), .A(n5883), .ZN(U2992) );
  NAND2_X1 U7055 ( .A1(n5885), .A2(n6433), .ZN(n5887) );
  OAI211_X1 U7056 ( .C1(n5888), .C2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5887), .B(n5886), .ZN(n5889) );
  AOI21_X1 U7057 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5890), .A(n5889), 
        .ZN(n5891) );
  OAI21_X1 U7058 ( .B1(n5892), .B2(n6381), .A(n5891), .ZN(U2993) );
  INV_X1 U7059 ( .A(n5893), .ZN(n5896) );
  AOI21_X1 U7060 ( .B1(n5901), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5894) );
  NOR2_X1 U7061 ( .A1(n2976), .A2(n5894), .ZN(n5895) );
  AOI211_X1 U7062 ( .C1(n6433), .C2(n5897), .A(n5896), .B(n5895), .ZN(n5898)
         );
  OAI21_X1 U7063 ( .B1(n5899), .B2(n6381), .A(n5898), .ZN(U2994) );
  NAND2_X1 U7064 ( .A1(n5901), .A2(n5900), .ZN(n5903) );
  OAI211_X1 U7065 ( .C1(n6034), .C2(n5904), .A(n5903), .B(n5902), .ZN(n5905)
         );
  AOI21_X1 U7066 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5906), .A(n5905), 
        .ZN(n5907) );
  OAI21_X1 U7067 ( .B1(n5908), .B2(n6381), .A(n5907), .ZN(U2995) );
  NOR3_X1 U7068 ( .A1(n5921), .A2(n5910), .A3(n5909), .ZN(n5915) );
  INV_X1 U7069 ( .A(n5911), .ZN(n5913) );
  OAI21_X1 U7070 ( .B1(n5913), .B2(n6034), .A(n5912), .ZN(n5914) );
  AOI211_X1 U7071 ( .C1(INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n5923), .A(n5915), .B(n5914), .ZN(n5916) );
  OAI21_X1 U7072 ( .B1(n5917), .B2(n6381), .A(n5916), .ZN(U2996) );
  NAND2_X1 U7073 ( .A1(n5918), .A2(n6433), .ZN(n5920) );
  OAI211_X1 U7074 ( .C1(n5921), .C2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5920), .B(n5919), .ZN(n5922) );
  AOI21_X1 U7075 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5923), .A(n5922), 
        .ZN(n5924) );
  OAI21_X1 U7076 ( .B1(n5925), .B2(n6381), .A(n5924), .ZN(U2997) );
  NOR3_X1 U7077 ( .A1(n6000), .A2(n5956), .A3(n5926), .ZN(n5929) );
  OAI21_X1 U7078 ( .B1(n5929), .B2(n5928), .A(n5927), .ZN(n5962) );
  AOI21_X1 U7079 ( .B1(n6441), .B2(n5956), .A(n5962), .ZN(n5946) );
  OAI21_X1 U7080 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6380), .A(n5946), 
        .ZN(n5943) );
  OR3_X1 U7081 ( .A1(n5941), .A2(n5931), .A3(n5930), .ZN(n5932) );
  OAI211_X1 U7082 ( .C1(n5934), .C2(n6034), .A(n5933), .B(n5932), .ZN(n5935)
         );
  AOI21_X1 U7083 ( .B1(n5943), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5935), 
        .ZN(n5936) );
  OAI21_X1 U7084 ( .B1(n5937), .B2(n6381), .A(n5936), .ZN(U2998) );
  NAND2_X1 U7085 ( .A1(n5938), .A2(n6433), .ZN(n5940) );
  OAI211_X1 U7086 ( .C1(n5941), .C2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5940), .B(n5939), .ZN(n5942) );
  AOI21_X1 U7087 ( .B1(n5943), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5942), 
        .ZN(n5944) );
  OAI21_X1 U7088 ( .B1(n5945), .B2(n6381), .A(n5944), .ZN(U2999) );
  INV_X1 U7089 ( .A(n5946), .ZN(n5952) );
  NAND4_X1 U7090 ( .A1(n6037), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5957), .A4(n5947), .ZN(n5949) );
  OAI211_X1 U7091 ( .C1(n6034), .C2(n5950), .A(n5949), .B(n5948), .ZN(n5951)
         );
  AOI21_X1 U7092 ( .B1(n5952), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n5951), 
        .ZN(n5953) );
  OAI21_X1 U7093 ( .B1(n5954), .B2(n6381), .A(n5953), .ZN(U3000) );
  INV_X1 U7094 ( .A(n5955), .ZN(n5960) );
  NAND3_X1 U7095 ( .A1(n6037), .A2(n5957), .A3(n5956), .ZN(n5959) );
  OAI211_X1 U7096 ( .C1(n6034), .C2(n5960), .A(n5959), .B(n5958), .ZN(n5961)
         );
  AOI21_X1 U7097 ( .B1(n5962), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5961), 
        .ZN(n5963) );
  OAI21_X1 U7098 ( .B1(n5964), .B2(n6381), .A(n5963), .ZN(U3001) );
  XNOR2_X1 U7099 ( .A(n5973), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5976)
         );
  INV_X1 U7100 ( .A(n6037), .ZN(n6019) );
  NOR2_X1 U7101 ( .A1(n6019), .A2(n5971), .ZN(n5985) );
  OAI21_X1 U7102 ( .B1(n5966), .B2(n6034), .A(n5965), .ZN(n5975) );
  NAND2_X1 U7103 ( .A1(n6000), .A2(n6043), .ZN(n5970) );
  INV_X1 U7104 ( .A(n5967), .ZN(n5968) );
  NAND2_X1 U7105 ( .A1(n6045), .A2(n5968), .ZN(n5969) );
  NAND2_X1 U7106 ( .A1(n5970), .A2(n5969), .ZN(n6038) );
  AOI21_X1 U7107 ( .B1(n5972), .B2(n5971), .A(n6038), .ZN(n5981) );
  NOR2_X1 U7108 ( .A1(n5981), .A2(n5973), .ZN(n5974) );
  AOI211_X1 U7109 ( .C1(n5976), .C2(n5985), .A(n5975), .B(n5974), .ZN(n5977)
         );
  OAI21_X1 U7110 ( .B1(n5978), .B2(n6381), .A(n5977), .ZN(U3002) );
  OAI21_X1 U7111 ( .B1(n5980), .B2(n6034), .A(n5979), .ZN(n5983) );
  NOR2_X1 U7112 ( .A1(n5981), .A2(n5984), .ZN(n5982) );
  AOI211_X1 U7113 ( .C1(n5985), .C2(n5984), .A(n5983), .B(n5982), .ZN(n5986)
         );
  OAI21_X1 U7114 ( .B1(n5987), .B2(n6381), .A(n5986), .ZN(U3003) );
  NAND3_X1 U7115 ( .A1(n6037), .A2(n5995), .A3(n5988), .ZN(n5990) );
  OAI211_X1 U7116 ( .C1(n6034), .C2(n5991), .A(n5990), .B(n5989), .ZN(n5992)
         );
  INV_X1 U7117 ( .A(n5992), .ZN(n6003) );
  INV_X1 U7118 ( .A(n5993), .ZN(n6015) );
  OAI22_X1 U7119 ( .A1(n5996), .A2(n6015), .B1(n5995), .B2(n5994), .ZN(n5997)
         );
  OR2_X1 U7120 ( .A1(n6038), .A2(n5997), .ZN(n6010) );
  NAND2_X1 U7121 ( .A1(n6015), .A2(n5998), .ZN(n6008) );
  AOI21_X1 U7122 ( .B1(n6000), .B2(n5999), .A(n6008), .ZN(n6001) );
  OAI21_X1 U7123 ( .B1(n6010), .B2(n6001), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n6002) );
  OAI211_X1 U7124 ( .C1(n6004), .C2(n6381), .A(n6003), .B(n6002), .ZN(U3004)
         );
  NAND2_X1 U7125 ( .A1(n6005), .A2(n6433), .ZN(n6007) );
  OAI211_X1 U7126 ( .C1(n6019), .C2(n6008), .A(n6007), .B(n6006), .ZN(n6009)
         );
  AOI21_X1 U7127 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n6010), .A(n6009), 
        .ZN(n6011) );
  OAI21_X1 U7128 ( .B1(n6012), .B2(n6381), .A(n6011), .ZN(U3005) );
  AOI21_X1 U7129 ( .B1(n6014), .B2(n6433), .A(n6013), .ZN(n6023) );
  AOI21_X1 U7130 ( .B1(n6017), .B2(n6016), .A(n6015), .ZN(n6021) );
  OAI21_X1 U7131 ( .B1(n6019), .B2(n6036), .A(n6018), .ZN(n6020) );
  OAI21_X1 U7132 ( .B1(n6021), .B2(n6038), .A(n6020), .ZN(n6022) );
  OAI211_X1 U7133 ( .C1(n6024), .C2(n6381), .A(n6023), .B(n6022), .ZN(U3006)
         );
  AOI22_X1 U7134 ( .A1(n6025), .A2(n2964), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n5793), .ZN(n6028) );
  XNOR2_X1 U7135 ( .A(n6026), .B(n6036), .ZN(n6027) );
  XNOR2_X1 U7136 ( .A(n6028), .B(n6027), .ZN(n6346) );
  INV_X1 U7137 ( .A(n6029), .ZN(n6258) );
  AOI21_X1 U7138 ( .B1(n6258), .B2(n6031), .A(n6030), .ZN(n6033) );
  OR2_X1 U7139 ( .A1(n6033), .A2(n6032), .ZN(n6294) );
  NAND2_X1 U7140 ( .A1(n6364), .A2(REIP_REG_11__SCAN_IN), .ZN(n6338) );
  OAI21_X1 U7141 ( .B1(n6294), .B2(n6034), .A(n6338), .ZN(n6035) );
  AOI21_X1 U7142 ( .B1(n6037), .B2(n6036), .A(n6035), .ZN(n6040) );
  NAND2_X1 U7143 ( .A1(n6038), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6039) );
  OAI211_X1 U7144 ( .C1(n6346), .C2(n6381), .A(n6040), .B(n6039), .ZN(U3007)
         );
  NOR3_X1 U7145 ( .A1(n6425), .A2(n6061), .A3(n6062), .ZN(n6397) );
  OAI21_X1 U7146 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6397), .ZN(n6047) );
  AOI22_X1 U7147 ( .A1(n6045), .A2(n6044), .B1(n6043), .B2(n6042), .ZN(n6401)
         );
  OAI22_X1 U7148 ( .A1(n6379), .A2(n6047), .B1(n6401), .B2(n6046), .ZN(n6048)
         );
  AOI211_X1 U7149 ( .C1(n6433), .C2(n6278), .A(n6049), .B(n6048), .ZN(n6050)
         );
  OAI21_X1 U7150 ( .B1(n6381), .B2(n6051), .A(n6050), .ZN(U3010) );
  OR2_X1 U7151 ( .A1(n6053), .A2(n6052), .ZN(n6054) );
  NAND2_X1 U7152 ( .A1(n6055), .A2(n6054), .ZN(n6349) );
  OAI22_X1 U7154 ( .A1(n6057), .A2(n6434), .B1(n6056), .B2(n6435), .ZN(n6437)
         );
  AOI21_X1 U7155 ( .B1(n6434), .B2(n6436), .A(n6437), .ZN(n6430) );
  OAI21_X1 U7156 ( .B1(n6410), .B2(n6380), .A(n6430), .ZN(n6058) );
  AOI221_X1 U7157 ( .B1(n6434), .B2(n6060), .C1(n6059), .C2(n6060), .A(n6058), 
        .ZN(n6409) );
  OAI33_X1 U7158 ( .A1(1'b0), .A2(n6409), .A3(n6062), .B1(
        INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6425), .B3(n6061), .ZN(n6064) );
  INV_X1 U7159 ( .A(n6064), .ZN(n6067) );
  NOR2_X1 U7160 ( .A1(n6412), .A2(n6844), .ZN(n6347) );
  AOI21_X1 U7161 ( .B1(n6065), .B2(n6433), .A(n6347), .ZN(n6066) );
  OAI211_X1 U7162 ( .C1(n6381), .C2(n6349), .A(n6067), .B(n6066), .ZN(U3012)
         );
  NAND2_X1 U7163 ( .A1(n6068), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6509) );
  OAI211_X1 U7164 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6068), .A(n6509), .B(
        n6515), .ZN(n6069) );
  OAI21_X1 U7165 ( .B1(n6674), .B2(n6070), .A(n6069), .ZN(n6071) );
  MUX2_X1 U7166 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n6071), .S(n6682), 
        .Z(U3464) );
  XNOR2_X1 U7167 ( .A(n6670), .B(n6509), .ZN(n6072) );
  OAI22_X1 U7168 ( .A1(n6072), .A2(n6672), .B1(n6674), .B2(n4636), .ZN(n6073)
         );
  MUX2_X1 U7169 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n6073), .S(n6682), 
        .Z(U3463) );
  NOR2_X2 U7170 ( .A1(n6074), .A2(n6671), .ZN(n6455) );
  OAI21_X1 U7171 ( .B1(n6075), .B2(n6455), .A(n6676), .ZN(n6077) );
  NAND2_X1 U7172 ( .A1(n6675), .A2(n6076), .ZN(n6112) );
  AOI21_X1 U7173 ( .B1(n6077), .B2(n6112), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n6079) );
  NOR2_X1 U7174 ( .A1(n6115), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6082)
         );
  AOI21_X1 U7175 ( .B1(STATE2_REG_2__SCAN_IN), .B2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n6078), .ZN(n6476) );
  NAND2_X1 U7176 ( .A1(n6104), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6085) );
  OR2_X1 U7177 ( .A1(n6112), .A2(n6672), .ZN(n6081) );
  INV_X1 U7178 ( .A(n6139), .ZN(n6473) );
  NAND3_X1 U7179 ( .A1(n6473), .A2(n6464), .A3(n6681), .ZN(n6080) );
  INV_X1 U7180 ( .A(n6082), .ZN(n6105) );
  OAI22_X1 U7181 ( .A1(n6106), .A2(n6566), .B1(n6506), .B2(n6105), .ZN(n6083)
         );
  AOI21_X1 U7182 ( .B1(n6455), .B2(n6563), .A(n6083), .ZN(n6084) );
  OAI211_X1 U7183 ( .C1(n6110), .C2(n6507), .A(n6085), .B(n6084), .ZN(U3036)
         );
  NAND2_X1 U7184 ( .A1(n6104), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6088) );
  OAI22_X1 U7185 ( .A1(n6106), .A2(n6705), .B1(n6699), .B2(n6105), .ZN(n6086)
         );
  AOI21_X1 U7186 ( .B1(n6455), .B2(n6595), .A(n6086), .ZN(n6087) );
  OAI211_X1 U7187 ( .C1(n6110), .C2(n6701), .A(n6088), .B(n6087), .ZN(U3037)
         );
  NAND2_X1 U7188 ( .A1(n6104), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n6091) );
  OAI22_X1 U7189 ( .A1(n6106), .A2(n6571), .B1(n6519), .B2(n6105), .ZN(n6089)
         );
  AOI21_X1 U7190 ( .B1(n6455), .B2(n6602), .A(n6089), .ZN(n6090) );
  OAI211_X1 U7191 ( .C1(n6110), .C2(n6162), .A(n6091), .B(n6090), .ZN(U3038)
         );
  NAND2_X1 U7192 ( .A1(n6104), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n6094) );
  OAI22_X1 U7193 ( .A1(n6106), .A2(n6574), .B1(n6524), .B2(n6105), .ZN(n6092)
         );
  AOI21_X1 U7194 ( .B1(n6455), .B2(n6609), .A(n6092), .ZN(n6093) );
  OAI211_X1 U7195 ( .C1(n6110), .C2(n6167), .A(n6094), .B(n6093), .ZN(U3039)
         );
  NAND2_X1 U7196 ( .A1(n6104), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n6097) );
  OAI22_X1 U7197 ( .A1(n6106), .A2(n6577), .B1(n6529), .B2(n6105), .ZN(n6095)
         );
  AOI21_X1 U7198 ( .B1(n6455), .B2(n6616), .A(n6095), .ZN(n6096) );
  OAI211_X1 U7199 ( .C1(n6110), .C2(n6172), .A(n6097), .B(n6096), .ZN(U3040)
         );
  NAND2_X1 U7200 ( .A1(n6104), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n6100) );
  OAI22_X1 U7201 ( .A1(n6106), .A2(n6580), .B1(n6534), .B2(n6105), .ZN(n6098)
         );
  AOI21_X1 U7202 ( .B1(n6455), .B2(n6623), .A(n6098), .ZN(n6099) );
  OAI211_X1 U7203 ( .C1(n6110), .C2(n6535), .A(n6100), .B(n6099), .ZN(U3041)
         );
  NAND2_X1 U7204 ( .A1(n6104), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n6103) );
  OAI22_X1 U7205 ( .A1(n6106), .A2(n6583), .B1(n6539), .B2(n6105), .ZN(n6101)
         );
  AOI21_X1 U7206 ( .B1(n6455), .B2(n6630), .A(n6101), .ZN(n6102) );
  OAI211_X1 U7207 ( .C1(n6110), .C2(n6181), .A(n6103), .B(n6102), .ZN(U3042)
         );
  NAND2_X1 U7208 ( .A1(n6104), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6109) );
  OAI22_X1 U7209 ( .A1(n6106), .A2(n6590), .B1(n6545), .B2(n6105), .ZN(n6107)
         );
  AOI21_X1 U7210 ( .B1(n6455), .B2(n6639), .A(n6107), .ZN(n6108) );
  OAI211_X1 U7211 ( .C1(n6110), .C2(n6546), .A(n6109), .B(n6108), .ZN(U3043)
         );
  INV_X1 U7212 ( .A(n6509), .ZN(n6111) );
  AOI21_X1 U7213 ( .B1(n6111), .B2(n6670), .A(n6672), .ZN(n6551) );
  INV_X1 U7214 ( .A(n6551), .ZN(n6120) );
  OR2_X1 U7215 ( .A1(n6112), .A2(n3501), .ZN(n6114) );
  INV_X1 U7216 ( .A(n6115), .ZN(n6113) );
  NAND2_X1 U7217 ( .A1(n6113), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6453) );
  AND2_X1 U7218 ( .A1(n6114), .A2(n6453), .ZN(n6116) );
  OAI22_X1 U7219 ( .A1(n6120), .A2(n6116), .B1(n6657), .B2(n6115), .ZN(n6456)
         );
  INV_X1 U7220 ( .A(n6116), .ZN(n6119) );
  NAND2_X1 U7221 ( .A1(n6672), .A2(n6117), .ZN(n6118) );
  AND2_X1 U7222 ( .A1(n6513), .A2(n6118), .ZN(n6560) );
  OAI211_X1 U7223 ( .C1(n6120), .C2(n6119), .A(n6560), .B(n6681), .ZN(n6457)
         );
  NOR2_X1 U7224 ( .A1(n6460), .A2(n6481), .ZN(n6122) );
  INV_X1 U7225 ( .A(n6455), .ZN(n6133) );
  OAI22_X1 U7226 ( .A1(n6133), .A2(n6507), .B1(n6506), .B2(n6453), .ZN(n6121)
         );
  AOI211_X1 U7227 ( .C1(n6457), .C2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n6122), 
        .B(n6121), .ZN(n6123) );
  OAI21_X1 U7228 ( .B1(n6137), .B2(n6566), .A(n6123), .ZN(U3044) );
  NOR2_X1 U7229 ( .A1(n6460), .A2(n6704), .ZN(n6125) );
  OAI22_X1 U7230 ( .A1(n6133), .A2(n6701), .B1(n6699), .B2(n6453), .ZN(n6124)
         );
  AOI211_X1 U7231 ( .C1(n6457), .C2(INSTQUEUE_REG_3__1__SCAN_IN), .A(n6125), 
        .B(n6124), .ZN(n6126) );
  OAI21_X1 U7232 ( .B1(n6137), .B2(n6705), .A(n6126), .ZN(U3045) );
  NOR2_X1 U7233 ( .A1(n6460), .A2(n6492), .ZN(n6128) );
  OAI22_X1 U7234 ( .A1(n6133), .A2(n6535), .B1(n6534), .B2(n6453), .ZN(n6127)
         );
  AOI211_X1 U7235 ( .C1(n6457), .C2(INSTQUEUE_REG_3__5__SCAN_IN), .A(n6128), 
        .B(n6127), .ZN(n6129) );
  OAI21_X1 U7236 ( .B1(n6137), .B2(n6580), .A(n6129), .ZN(U3049) );
  NOR2_X1 U7237 ( .A1(n6460), .A2(n6540), .ZN(n6131) );
  OAI22_X1 U7238 ( .A1(n6133), .A2(n6181), .B1(n6539), .B2(n6453), .ZN(n6130)
         );
  AOI211_X1 U7239 ( .C1(n6457), .C2(INSTQUEUE_REG_3__6__SCAN_IN), .A(n6131), 
        .B(n6130), .ZN(n6132) );
  OAI21_X1 U7240 ( .B1(n6137), .B2(n6583), .A(n6132), .ZN(U3050) );
  NOR2_X1 U7241 ( .A1(n6460), .A2(n6501), .ZN(n6135) );
  OAI22_X1 U7242 ( .A1(n6133), .A2(n6546), .B1(n6545), .B2(n6453), .ZN(n6134)
         );
  AOI211_X1 U7243 ( .C1(n6457), .C2(INSTQUEUE_REG_3__7__SCAN_IN), .A(n6135), 
        .B(n6134), .ZN(n6136) );
  OAI21_X1 U7244 ( .B1(n6137), .B2(n6590), .A(n6136), .ZN(U3051) );
  NAND2_X1 U7245 ( .A1(n6138), .A2(n6145), .ZN(n6142) );
  OR2_X1 U7246 ( .A1(n6140), .A2(n6139), .ZN(n6141) );
  NAND2_X1 U7247 ( .A1(n6142), .A2(n6141), .ZN(n6190) );
  NAND2_X1 U7248 ( .A1(n6143), .A2(n6463), .ZN(n6187) );
  INV_X1 U7249 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n6153) );
  AOI21_X1 U7250 ( .B1(n6145), .B2(n6144), .A(n6672), .ZN(n6149) );
  INV_X1 U7251 ( .A(n6703), .ZN(n6548) );
  OAI21_X1 U7252 ( .B1(n6147), .B2(n6548), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6148) );
  AOI22_X1 U7253 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6187), .B1(n6149), .B2(
        n6148), .ZN(n6151) );
  OAI22_X1 U7254 ( .A1(n6506), .A2(n6187), .B1(n6153), .B2(n6185), .ZN(n6155)
         );
  NOR2_X1 U7255 ( .A1(n6703), .A2(n6507), .ZN(n6154) );
  AOI211_X1 U7256 ( .C1(n6468), .C2(n6190), .A(n6155), .B(n6154), .ZN(n6156)
         );
  OAI21_X1 U7257 ( .B1(n6481), .B2(n6192), .A(n6156), .ZN(U3084) );
  INV_X1 U7258 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n6157) );
  OAI22_X1 U7259 ( .A1(n6699), .A2(n6187), .B1(n6157), .B2(n6185), .ZN(n6159)
         );
  NOR2_X1 U7260 ( .A1(n6703), .A2(n6701), .ZN(n6158) );
  AOI211_X1 U7261 ( .C1(n6593), .C2(n6190), .A(n6159), .B(n6158), .ZN(n6160)
         );
  OAI21_X1 U7262 ( .B1(n6704), .B2(n6192), .A(n6160), .ZN(U3085) );
  INV_X1 U7263 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6161) );
  OAI22_X1 U7264 ( .A1(n6519), .A2(n6187), .B1(n6161), .B2(n6185), .ZN(n6164)
         );
  NOR2_X1 U7265 ( .A1(n6703), .A2(n6162), .ZN(n6163) );
  AOI211_X1 U7266 ( .C1(n6601), .C2(n6190), .A(n6164), .B(n6163), .ZN(n6165)
         );
  OAI21_X1 U7267 ( .B1(n6520), .B2(n6192), .A(n6165), .ZN(U3086) );
  INV_X1 U7268 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n6166) );
  OAI22_X1 U7269 ( .A1(n6524), .A2(n6187), .B1(n6166), .B2(n6185), .ZN(n6169)
         );
  NOR2_X1 U7270 ( .A1(n6703), .A2(n6167), .ZN(n6168) );
  AOI211_X1 U7271 ( .C1(n6608), .C2(n6190), .A(n6169), .B(n6168), .ZN(n6170)
         );
  OAI21_X1 U7272 ( .B1(n6525), .B2(n6192), .A(n6170), .ZN(U3087) );
  INV_X1 U7273 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6171) );
  OAI22_X1 U7274 ( .A1(n6529), .A2(n6187), .B1(n6171), .B2(n6185), .ZN(n6174)
         );
  NOR2_X1 U7275 ( .A1(n6703), .A2(n6172), .ZN(n6173) );
  AOI211_X1 U7276 ( .C1(n6615), .C2(n6190), .A(n6174), .B(n6173), .ZN(n6175)
         );
  OAI21_X1 U7277 ( .B1(n6530), .B2(n6192), .A(n6175), .ZN(U3088) );
  INV_X1 U7278 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n6176) );
  OAI22_X1 U7279 ( .A1(n6534), .A2(n6187), .B1(n6176), .B2(n6185), .ZN(n6178)
         );
  NOR2_X1 U7280 ( .A1(n6703), .A2(n6535), .ZN(n6177) );
  AOI211_X1 U7281 ( .C1(n6622), .C2(n6190), .A(n6178), .B(n6177), .ZN(n6179)
         );
  OAI21_X1 U7282 ( .B1(n6492), .B2(n6192), .A(n6179), .ZN(U3089) );
  INV_X1 U7283 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n6180) );
  OAI22_X1 U7284 ( .A1(n6539), .A2(n6187), .B1(n6180), .B2(n6185), .ZN(n6183)
         );
  NOR2_X1 U7285 ( .A1(n6703), .A2(n6181), .ZN(n6182) );
  AOI211_X1 U7286 ( .C1(n6629), .C2(n6190), .A(n6183), .B(n6182), .ZN(n6184)
         );
  OAI21_X1 U7287 ( .B1(n6540), .B2(n6192), .A(n6184), .ZN(U3090) );
  INV_X1 U7288 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n6186) );
  OAI22_X1 U7289 ( .A1(n6545), .A2(n6187), .B1(n6186), .B2(n6185), .ZN(n6189)
         );
  NOR2_X1 U7290 ( .A1(n6703), .A2(n6546), .ZN(n6188) );
  AOI211_X1 U7291 ( .C1(n6637), .C2(n6190), .A(n6189), .B(n6188), .ZN(n6191)
         );
  OAI21_X1 U7292 ( .B1(n6501), .B2(n6192), .A(n6191), .ZN(U3091) );
  INV_X1 U7293 ( .A(n6193), .ZN(n6217) );
  INV_X1 U7294 ( .A(n6194), .ZN(n6203) );
  AOI211_X1 U7295 ( .C1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n6196), .A(n6463), .B(n6195), .ZN(n6199) );
  NAND2_X1 U7296 ( .A1(n6199), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6201) );
  OAI22_X1 U7297 ( .A1(n6199), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n6198), .B2(n6197), .ZN(n6200) );
  NAND2_X1 U7298 ( .A1(n6201), .A2(n6200), .ZN(n6202) );
  AOI222_X1 U7299 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6203), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6202), .C1(n6203), .C2(n6202), 
        .ZN(n6204) );
  OR2_X1 U7300 ( .A1(n6204), .A2(n6681), .ZN(n6205) );
  AOI22_X1 U7301 ( .A1(n6206), .A2(n6205), .B1(n6204), .B2(n6681), .ZN(n6214)
         );
  OAI21_X1 U7302 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6207), 
        .ZN(n6208) );
  AND4_X1 U7303 ( .A1(n6211), .A2(n6210), .A3(n6209), .A4(n6208), .ZN(n6213)
         );
  OAI211_X1 U7304 ( .C1(n6214), .C2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n6213), .B(n6212), .ZN(n6650) );
  INV_X1 U7305 ( .A(n6650), .ZN(n6215) );
  AOI22_X1 U7306 ( .A1(n6215), .A2(n6654), .B1(n6331), .B2(READY_N), .ZN(n6216) );
  AOI21_X1 U7307 ( .B1(n6218), .B2(n6217), .A(n6216), .ZN(n6663) );
  OAI21_X1 U7308 ( .B1(n6663), .B2(n6747), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n6219) );
  NAND2_X1 U7309 ( .A1(n6219), .A2(n6665), .ZN(U3453) );
  MUX2_X1 U7310 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n2966), .Z(U3448) );
  MUX2_X1 U7311 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n2966), .Z(U3447) );
  MUX2_X1 U7312 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n2966), .Z(U3446) );
  MUX2_X1 U7313 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n2966), .Z(U3445) );
  AND2_X1 U7314 ( .A1(n6330), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U7315 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n6221), .A(n6220), .ZN(
        n6222) );
  INV_X1 U7316 ( .A(n6222), .ZN(U2788) );
  NAND2_X1 U7317 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6694), .ZN(n6226) );
  OAI21_X1 U7318 ( .B1(n6224), .B2(n6223), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6225) );
  OAI21_X1 U7319 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6226), .A(n6225), .ZN(
        U2790) );
  INV_X1 U7320 ( .A(n6227), .ZN(n6229) );
  OAI21_X1 U7321 ( .B1(n6229), .B2(n6228), .A(n6345), .ZN(U2793) );
  NOR4_X1 U7322 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(n6230) );
  OAI21_X1 U7323 ( .B1(n6244), .B2(n6231), .A(n6230), .ZN(n6240) );
  NOR3_X1 U7324 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6725)
         );
  NOR4_X1 U7325 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n6233) );
  NOR2_X1 U7326 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n6232) );
  NAND3_X1 U7327 ( .A1(n6725), .A2(n6233), .A3(n6232), .ZN(n6239) );
  NOR4_X1 U7328 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6237)
         );
  NOR4_X1 U7329 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n6236) );
  NOR4_X1 U7330 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(
        DATAWIDTH_REG_26__SCAN_IN), .A3(DATAWIDTH_REG_28__SCAN_IN), .A4(
        DATAWIDTH_REG_30__SCAN_IN), .ZN(n6235) );
  NOR4_X1 U7331 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6234) );
  NAND4_X1 U7332 ( .A1(n6237), .A2(n6236), .A3(n6235), .A4(n6234), .ZN(n6238)
         );
  NOR4_X2 U7333 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6240), .A3(n6239), .A4(
        n6238), .ZN(n6686) );
  INV_X1 U7334 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6242) );
  NOR3_X1 U7335 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6243) );
  OAI21_X1 U7336 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6243), .A(n6686), .ZN(n6241)
         );
  OAI21_X1 U7337 ( .B1(n6686), .B2(n6242), .A(n6241), .ZN(U2794) );
  AOI21_X1 U7338 ( .B1(n6815), .B2(n6244), .A(n6243), .ZN(n6246) );
  INV_X1 U7339 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6245) );
  INV_X1 U7340 ( .A(n6686), .ZN(n6688) );
  AOI22_X1 U7341 ( .A1(n6686), .A2(n6246), .B1(n6245), .B2(n6688), .ZN(U2795)
         );
  NAND3_X1 U7342 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        n6257), .ZN(n6256) );
  INV_X1 U7343 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6777) );
  INV_X1 U7344 ( .A(n6294), .ZN(n6248) );
  AOI22_X1 U7345 ( .A1(n6279), .A2(n6248), .B1(REIP_REG_11__SCAN_IN), .B2(
        n6247), .ZN(n6250) );
  OAI211_X1 U7346 ( .C1(n6251), .C2(n6777), .A(n6250), .B(n6249), .ZN(n6252)
         );
  AOI21_X1 U7347 ( .B1(n6260), .B2(EBX_REG_11__SCAN_IN), .A(n6252), .ZN(n6255)
         );
  OAI22_X1 U7348 ( .A1(n6341), .A2(n6282), .B1(n6340), .B2(n6280), .ZN(n6253)
         );
  INV_X1 U7349 ( .A(n6253), .ZN(n6254) );
  OAI211_X1 U7350 ( .C1(REIP_REG_11__SCAN_IN), .C2(n6256), .A(n6255), .B(n6254), .ZN(U2816) );
  INV_X1 U7351 ( .A(n6257), .ZN(n6270) );
  AOI21_X1 U7352 ( .B1(n6259), .B2(n4982), .A(n6258), .ZN(n6388) );
  AOI22_X1 U7353 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6260), .B1(n6279), .B2(n6388), 
        .ZN(n6261) );
  OAI21_X1 U7354 ( .B1(n6262), .B2(n6287), .A(n6261), .ZN(n6263) );
  AOI211_X1 U7355 ( .C1(n6273), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6272), 
        .B(n6263), .ZN(n6269) );
  INV_X1 U7356 ( .A(n6264), .ZN(n6300) );
  AOI22_X1 U7357 ( .A1(n6300), .A2(n6267), .B1(n6266), .B2(n6265), .ZN(n6268)
         );
  OAI211_X1 U7358 ( .C1(REIP_REG_9__SCAN_IN), .C2(n6270), .A(n6269), .B(n6268), 
        .ZN(U2818) );
  AOI21_X1 U7359 ( .B1(REIP_REG_7__SCAN_IN), .B2(n6271), .A(
        REIP_REG_8__SCAN_IN), .ZN(n6288) );
  AOI21_X1 U7360 ( .B1(n6273), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6272), 
        .ZN(n6274) );
  OAI21_X1 U7361 ( .B1(n6276), .B2(n6275), .A(n6274), .ZN(n6277) );
  AOI21_X1 U7362 ( .B1(n6279), .B2(n6278), .A(n6277), .ZN(n6286) );
  OAI22_X1 U7363 ( .A1(n6283), .A2(n6282), .B1(n6281), .B2(n6280), .ZN(n6284)
         );
  INV_X1 U7364 ( .A(n6284), .ZN(n6285) );
  OAI211_X1 U7365 ( .C1(n6288), .C2(n6287), .A(n6286), .B(n6285), .ZN(U2819)
         );
  NOR2_X1 U7366 ( .A1(n6289), .A2(n6295), .ZN(n6290) );
  AOI21_X1 U7367 ( .B1(n6291), .B2(n6299), .A(n6290), .ZN(n6292) );
  OAI21_X1 U7368 ( .B1(n6293), .B2(n6302), .A(n6292), .ZN(U2846) );
  OAI22_X1 U7369 ( .A1(n6341), .A2(n5588), .B1(n6295), .B2(n6294), .ZN(n6296)
         );
  INV_X1 U7370 ( .A(n6296), .ZN(n6297) );
  OAI21_X1 U7371 ( .B1(n6298), .B2(n6302), .A(n6297), .ZN(U2848) );
  INV_X1 U7372 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6303) );
  AOI22_X1 U7373 ( .A1(n6300), .A2(n6299), .B1(n4196), .B2(n6388), .ZN(n6301)
         );
  OAI21_X1 U7374 ( .B1(n6303), .B2(n6302), .A(n6301), .ZN(U2850) );
  AOI22_X1 U7375 ( .A1(n6330), .A2(DATAO_REG_26__SCAN_IN), .B1(n6306), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n6304) );
  OAI21_X1 U7376 ( .B1(n6335), .B2(n6781), .A(n6304), .ZN(U2897) );
  AOI22_X1 U7377 ( .A1(n6330), .A2(DATAO_REG_25__SCAN_IN), .B1(n6306), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6305) );
  OAI21_X1 U7378 ( .B1(n6335), .B2(n6816), .A(n6305), .ZN(U2898) );
  INV_X1 U7379 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n6769) );
  AOI22_X1 U7380 ( .A1(n6306), .A2(EAX_REG_19__SCAN_IN), .B1(n6331), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n6307) );
  OAI21_X1 U7381 ( .B1(n6769), .B2(n6337), .A(n6307), .ZN(U2904) );
  AOI22_X1 U7382 ( .A1(n6331), .A2(LWORD_REG_15__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6308) );
  OAI21_X1 U7383 ( .B1(n6309), .B2(n6336), .A(n6308), .ZN(U2908) );
  INV_X1 U7384 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n6803) );
  AOI22_X1 U7385 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6321), .B1(n6330), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6310) );
  OAI21_X1 U7386 ( .B1(n6335), .B2(n6803), .A(n6310), .ZN(U2909) );
  AOI22_X1 U7387 ( .A1(n6331), .A2(LWORD_REG_13__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6311) );
  OAI21_X1 U7388 ( .B1(n6804), .B2(n6336), .A(n6311), .ZN(U2910) );
  AOI22_X1 U7389 ( .A1(n6331), .A2(LWORD_REG_12__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6312) );
  OAI21_X1 U7390 ( .B1(n6738), .B2(n6336), .A(n6312), .ZN(U2911) );
  INV_X1 U7391 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6314) );
  AOI22_X1 U7392 ( .A1(n6331), .A2(LWORD_REG_11__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6313) );
  OAI21_X1 U7393 ( .B1(n6314), .B2(n6336), .A(n6313), .ZN(U2912) );
  AOI22_X1 U7394 ( .A1(n6331), .A2(LWORD_REG_10__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6315) );
  OAI21_X1 U7395 ( .B1(n6316), .B2(n6336), .A(n6315), .ZN(U2913) );
  AOI22_X1 U7396 ( .A1(n6331), .A2(LWORD_REG_9__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6317) );
  OAI21_X1 U7397 ( .B1(n6318), .B2(n6336), .A(n6317), .ZN(U2914) );
  AOI22_X1 U7398 ( .A1(n6331), .A2(LWORD_REG_8__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6319) );
  OAI21_X1 U7399 ( .B1(n6826), .B2(n6336), .A(n6319), .ZN(U2915) );
  AOI22_X1 U7400 ( .A1(n6331), .A2(LWORD_REG_7__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6320) );
  OAI21_X1 U7401 ( .B1(n4995), .B2(n6336), .A(n6320), .ZN(U2916) );
  INV_X1 U7402 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n6801) );
  AOI22_X1 U7403 ( .A1(EAX_REG_6__SCAN_IN), .A2(n6321), .B1(n6331), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n6322) );
  OAI21_X1 U7404 ( .B1(n6801), .B2(n6337), .A(n6322), .ZN(U2917) );
  INV_X1 U7405 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n6847) );
  INV_X1 U7406 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n6323) );
  OAI222_X1 U7407 ( .A1(n6337), .A2(n6847), .B1(n6336), .B2(n6324), .C1(n6335), 
        .C2(n6323), .ZN(U2918) );
  INV_X1 U7408 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n6734) );
  INV_X1 U7409 ( .A(LWORD_REG_4__SCAN_IN), .ZN(n6732) );
  OAI222_X1 U7410 ( .A1(n6337), .A2(n6734), .B1(n6336), .B2(n6325), .C1(n6335), 
        .C2(n6732), .ZN(U2919) );
  AOI22_X1 U7411 ( .A1(n6331), .A2(LWORD_REG_3__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6326) );
  OAI21_X1 U7412 ( .B1(n6327), .B2(n6336), .A(n6326), .ZN(U2920) );
  AOI22_X1 U7413 ( .A1(n6331), .A2(LWORD_REG_2__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6328) );
  OAI21_X1 U7414 ( .B1(n6329), .B2(n6336), .A(n6328), .ZN(U2921) );
  AOI22_X1 U7415 ( .A1(n6331), .A2(LWORD_REG_1__SCAN_IN), .B1(n6330), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6332) );
  OAI21_X1 U7416 ( .B1(n6333), .B2(n6336), .A(n6332), .ZN(U2922) );
  INV_X1 U7417 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n6841) );
  INV_X1 U7418 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n6334) );
  OAI222_X1 U7419 ( .A1(n6337), .A2(n6841), .B1(n6336), .B2(n6746), .C1(n6335), 
        .C2(n6334), .ZN(U2923) );
  INV_X1 U7420 ( .A(n6338), .ZN(n6339) );
  AOI21_X1 U7421 ( .B1(n6365), .B2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6339), 
        .ZN(n6344) );
  OAI22_X1 U7422 ( .A1(n6341), .A2(n6358), .B1(n6340), .B2(n6375), .ZN(n6342)
         );
  INV_X1 U7423 ( .A(n6342), .ZN(n6343) );
  OAI211_X1 U7424 ( .C1(n6346), .C2(n6345), .A(n6344), .B(n6343), .ZN(U2975)
         );
  AOI21_X1 U7425 ( .B1(n6365), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6347), 
        .ZN(n6352) );
  OAI22_X1 U7426 ( .A1(n6349), .A2(n6345), .B1(n6348), .B2(n6358), .ZN(n6350)
         );
  INV_X1 U7427 ( .A(n6350), .ZN(n6351) );
  OAI211_X1 U7428 ( .C1(n6375), .C2(n6353), .A(n6352), .B(n6351), .ZN(U2980)
         );
  AOI22_X1 U7429 ( .A1(n6365), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6364), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n6362) );
  OR2_X1 U7430 ( .A1(n6355), .A2(n6354), .ZN(n6356) );
  NAND2_X1 U7431 ( .A1(n6357), .A2(n6356), .ZN(n6416) );
  OAI22_X1 U7432 ( .A1(n6416), .A2(n6345), .B1(n6359), .B2(n6358), .ZN(n6360)
         );
  INV_X1 U7433 ( .A(n6360), .ZN(n6361) );
  OAI211_X1 U7434 ( .C1(n6375), .C2(n6363), .A(n6362), .B(n6361), .ZN(U2982)
         );
  AND2_X1 U7435 ( .A1(n6364), .A2(REIP_REG_2__SCAN_IN), .ZN(n6431) );
  AOI21_X1 U7436 ( .B1(n6365), .B2(PHYADDRPOINTER_REG_2__SCAN_IN), .A(n6431), 
        .ZN(n6373) );
  XNOR2_X1 U7437 ( .A(n6366), .B(n6440), .ZN(n6368) );
  XNOR2_X1 U7438 ( .A(n6368), .B(n6367), .ZN(n6439) );
  AOI22_X1 U7439 ( .A1(n6371), .A2(n6370), .B1(n6439), .B2(n6369), .ZN(n6372)
         );
  OAI211_X1 U7440 ( .C1(n6375), .C2(n6374), .A(n6373), .B(n6372), .ZN(U2984)
         );
  NAND2_X1 U7441 ( .A1(n6379), .A2(n6397), .ZN(n6393) );
  AOI22_X1 U7442 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n5805), .B1(
        INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6376), .ZN(n6385) );
  AOI21_X1 U7443 ( .B1(n6378), .B2(n6433), .A(n6377), .ZN(n6384) );
  OAI21_X1 U7444 ( .B1(n6380), .B2(n6379), .A(n6401), .ZN(n6390) );
  INV_X1 U7445 ( .A(n6381), .ZN(n6438) );
  AOI22_X1 U7446 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n6390), .B1(n6382), .B2(n6438), .ZN(n6383) );
  OAI211_X1 U7447 ( .C1(n6393), .C2(n6385), .A(n6384), .B(n6383), .ZN(U3008)
         );
  INV_X1 U7448 ( .A(n6386), .ZN(n6387) );
  AOI21_X1 U7449 ( .B1(n6388), .B2(n6433), .A(n6387), .ZN(n6392) );
  AOI22_X1 U7450 ( .A1(n6390), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .B1(n6438), 
        .B2(n6389), .ZN(n6391) );
  OAI211_X1 U7451 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6393), .A(n6392), 
        .B(n6391), .ZN(U3009) );
  AOI21_X1 U7452 ( .B1(n6395), .B2(n6433), .A(n6394), .ZN(n6399) );
  AOI22_X1 U7453 ( .A1(n6397), .A2(n6400), .B1(n6396), .B2(n6438), .ZN(n6398)
         );
  OAI211_X1 U7454 ( .C1(n6401), .C2(n6400), .A(n6399), .B(n6398), .ZN(U3011)
         );
  INV_X1 U7455 ( .A(n6425), .ZN(n6402) );
  AOI21_X1 U7456 ( .B1(n6410), .B2(n6402), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .ZN(n6408) );
  INV_X1 U7457 ( .A(n6403), .ZN(n6405) );
  AOI22_X1 U7458 ( .A1(n6405), .A2(n6438), .B1(n6433), .B2(n6404), .ZN(n6407)
         );
  OAI211_X1 U7459 ( .C1(n6409), .C2(n6408), .A(n6407), .B(n6406), .ZN(U3013)
         );
  AOI211_X1 U7460 ( .C1(n6429), .C2(n6420), .A(n6425), .B(n6410), .ZN(n6418)
         );
  NOR2_X1 U7461 ( .A1(n6412), .A2(n6411), .ZN(n6413) );
  AOI21_X1 U7462 ( .B1(n6433), .B2(n6414), .A(n6413), .ZN(n6415) );
  OAI21_X1 U7463 ( .B1(n6416), .B2(n6381), .A(n6415), .ZN(n6417) );
  NOR2_X1 U7464 ( .A1(n6418), .A2(n6417), .ZN(n6419) );
  OAI21_X1 U7465 ( .B1(n6430), .B2(n6420), .A(n6419), .ZN(U3014) );
  INV_X1 U7466 ( .A(n6421), .ZN(n6422) );
  AOI21_X1 U7467 ( .B1(n6433), .B2(n6423), .A(n6422), .ZN(n6428) );
  OAI22_X1 U7468 ( .A1(n6425), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .B1(n6424), 
        .B2(n6381), .ZN(n6426) );
  INV_X1 U7469 ( .A(n6426), .ZN(n6427) );
  OAI211_X1 U7470 ( .C1(n6430), .C2(n6429), .A(n6428), .B(n6427), .ZN(U3015)
         );
  AOI21_X1 U7471 ( .B1(n6433), .B2(n6432), .A(n6431), .ZN(n6445) );
  OAI221_X1 U7472 ( .B1(n6436), .B2(n6435), .C1(n6436), .C2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(n6434), .ZN(n6444) );
  AOI22_X1 U7473 ( .A1(n6439), .A2(n6438), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n6437), .ZN(n6443) );
  NAND3_X1 U7474 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6441), .A3(n6440), 
        .ZN(n6442) );
  NAND4_X1 U7475 ( .A1(n6445), .A2(n6444), .A3(n6443), .A4(n6442), .ZN(U3016)
         );
  NOR2_X1 U7476 ( .A1(n6446), .A2(n6682), .ZN(U3019) );
  NOR2_X1 U7477 ( .A1(n6519), .A2(n6453), .ZN(n6447) );
  AOI21_X1 U7478 ( .B1(n6455), .B2(n6603), .A(n6447), .ZN(n6449) );
  AOI22_X1 U7479 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6457), .B1(n6601), 
        .B2(n6456), .ZN(n6448) );
  OAI211_X1 U7480 ( .C1(n6520), .C2(n6460), .A(n6449), .B(n6448), .ZN(U3046)
         );
  NOR2_X1 U7481 ( .A1(n6524), .A2(n6453), .ZN(n6450) );
  AOI21_X1 U7482 ( .B1(n6455), .B2(n6610), .A(n6450), .ZN(n6452) );
  AOI22_X1 U7483 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6457), .B1(n6608), 
        .B2(n6456), .ZN(n6451) );
  OAI211_X1 U7484 ( .C1(n6525), .C2(n6460), .A(n6452), .B(n6451), .ZN(U3047)
         );
  NOR2_X1 U7485 ( .A1(n6529), .A2(n6453), .ZN(n6454) );
  AOI21_X1 U7486 ( .B1(n6455), .B2(n6617), .A(n6454), .ZN(n6459) );
  AOI22_X1 U7487 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6457), .B1(n6615), 
        .B2(n6456), .ZN(n6458) );
  OAI211_X1 U7488 ( .C1(n6530), .C2(n6460), .A(n6459), .B(n6458), .ZN(U3048)
         );
  NAND2_X1 U7489 ( .A1(n6516), .A2(n6463), .ZN(n6474) );
  INV_X1 U7490 ( .A(n6474), .ZN(n6496) );
  NAND3_X1 U7491 ( .A1(n6675), .A2(n6472), .A3(n6515), .ZN(n6467) );
  NAND3_X1 U7492 ( .A1(n6465), .A2(n6464), .A3(n6681), .ZN(n6466) );
  NAND2_X1 U7493 ( .A1(n6467), .A2(n6466), .ZN(n6495) );
  AOI22_X1 U7494 ( .A1(n6557), .A2(n6496), .B1(n6468), .B2(n6495), .ZN(n6480)
         );
  AOI21_X1 U7495 ( .B1(n6702), .B2(n6470), .A(n6469), .ZN(n6478) );
  NAND2_X1 U7496 ( .A1(n6472), .A2(n6471), .ZN(n6502) );
  NAND2_X1 U7497 ( .A1(n6502), .A2(n6515), .ZN(n6477) );
  AOI21_X1 U7498 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6474), .A(n6473), .ZN(
        n6475) );
  OAI211_X1 U7499 ( .C1(n6478), .C2(n6477), .A(n6476), .B(n6475), .ZN(n6498)
         );
  AOI22_X1 U7500 ( .A1(n6498), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6558), 
        .B2(n6497), .ZN(n6479) );
  OAI211_X1 U7501 ( .C1(n6481), .C2(n6702), .A(n6480), .B(n6479), .ZN(U3068)
         );
  AOI22_X1 U7502 ( .A1(n6592), .A2(n6496), .B1(n6593), .B2(n6495), .ZN(n6483)
         );
  AOI22_X1 U7503 ( .A1(n6498), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6596), 
        .B2(n6497), .ZN(n6482) );
  OAI211_X1 U7504 ( .C1(n6704), .C2(n6702), .A(n6483), .B(n6482), .ZN(U3069)
         );
  AOI22_X1 U7505 ( .A1(n6600), .A2(n6496), .B1(n6601), .B2(n6495), .ZN(n6485)
         );
  AOI22_X1 U7506 ( .A1(n6498), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6603), 
        .B2(n6497), .ZN(n6484) );
  OAI211_X1 U7507 ( .C1(n6520), .C2(n6702), .A(n6485), .B(n6484), .ZN(U3070)
         );
  AOI22_X1 U7508 ( .A1(n6607), .A2(n6496), .B1(n6608), .B2(n6495), .ZN(n6487)
         );
  AOI22_X1 U7509 ( .A1(n6498), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6610), 
        .B2(n6497), .ZN(n6486) );
  OAI211_X1 U7510 ( .C1(n6525), .C2(n6702), .A(n6487), .B(n6486), .ZN(U3071)
         );
  AOI22_X1 U7511 ( .A1(n6614), .A2(n6496), .B1(n6615), .B2(n6495), .ZN(n6489)
         );
  AOI22_X1 U7512 ( .A1(n6498), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6617), 
        .B2(n6497), .ZN(n6488) );
  OAI211_X1 U7513 ( .C1(n6530), .C2(n6702), .A(n6489), .B(n6488), .ZN(U3072)
         );
  AOI22_X1 U7514 ( .A1(n6621), .A2(n6496), .B1(n6622), .B2(n6495), .ZN(n6491)
         );
  AOI22_X1 U7515 ( .A1(n6498), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6624), 
        .B2(n6497), .ZN(n6490) );
  OAI211_X1 U7516 ( .C1(n6492), .C2(n6702), .A(n6491), .B(n6490), .ZN(U3073)
         );
  AOI22_X1 U7517 ( .A1(n6628), .A2(n6496), .B1(n6629), .B2(n6495), .ZN(n6494)
         );
  AOI22_X1 U7518 ( .A1(n6498), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6631), 
        .B2(n6497), .ZN(n6493) );
  OAI211_X1 U7519 ( .C1(n6540), .C2(n6702), .A(n6494), .B(n6493), .ZN(U3074)
         );
  AOI22_X1 U7520 ( .A1(n6635), .A2(n6496), .B1(n6637), .B2(n6495), .ZN(n6500)
         );
  AOI22_X1 U7521 ( .A1(n6498), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6641), 
        .B2(n6497), .ZN(n6499) );
  OAI211_X1 U7522 ( .C1(n6501), .C2(n6702), .A(n6500), .B(n6499), .ZN(U3075)
         );
  INV_X1 U7523 ( .A(n6502), .ZN(n6504) );
  INV_X1 U7524 ( .A(n6700), .ZN(n6503) );
  AOI21_X1 U7525 ( .B1(n6504), .B2(n6552), .A(n6503), .ZN(n6511) );
  NOR2_X1 U7526 ( .A1(n6511), .A2(n6672), .ZN(n6505) );
  OAI22_X1 U7527 ( .A1(n6702), .A2(n6507), .B1(n6700), .B2(n6506), .ZN(n6508)
         );
  INV_X1 U7528 ( .A(n6508), .ZN(n6518) );
  NOR2_X1 U7529 ( .A1(n6510), .A2(n6509), .ZN(n6668) );
  INV_X1 U7530 ( .A(n6668), .ZN(n6512) );
  NAND3_X1 U7531 ( .A1(n6512), .A2(n6515), .A3(n6511), .ZN(n6514) );
  OAI211_X1 U7532 ( .C1(n6516), .C2(n6515), .A(n6514), .B(n6513), .ZN(n6709)
         );
  AOI22_X1 U7533 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6709), .B1(n6563), 
        .B2(n6548), .ZN(n6517) );
  OAI211_X1 U7534 ( .C1(n6706), .C2(n6566), .A(n6518), .B(n6517), .ZN(U3076)
         );
  OAI22_X1 U7535 ( .A1(n6703), .A2(n6520), .B1(n6700), .B2(n6519), .ZN(n6521)
         );
  INV_X1 U7536 ( .A(n6521), .ZN(n6523) );
  INV_X1 U7537 ( .A(n6702), .ZN(n6542) );
  AOI22_X1 U7538 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6709), .B1(n6603), 
        .B2(n6542), .ZN(n6522) );
  OAI211_X1 U7539 ( .C1(n6706), .C2(n6571), .A(n6523), .B(n6522), .ZN(U3078)
         );
  OAI22_X1 U7540 ( .A1(n6703), .A2(n6525), .B1(n6700), .B2(n6524), .ZN(n6526)
         );
  INV_X1 U7541 ( .A(n6526), .ZN(n6528) );
  AOI22_X1 U7542 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6709), .B1(n6610), 
        .B2(n6542), .ZN(n6527) );
  OAI211_X1 U7543 ( .C1(n6706), .C2(n6574), .A(n6528), .B(n6527), .ZN(U3079)
         );
  OAI22_X1 U7544 ( .A1(n6703), .A2(n6530), .B1(n6700), .B2(n6529), .ZN(n6531)
         );
  INV_X1 U7545 ( .A(n6531), .ZN(n6533) );
  AOI22_X1 U7546 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6709), .B1(n6617), 
        .B2(n6542), .ZN(n6532) );
  OAI211_X1 U7547 ( .C1(n6706), .C2(n6577), .A(n6533), .B(n6532), .ZN(U3080)
         );
  OAI22_X1 U7548 ( .A1(n6702), .A2(n6535), .B1(n6700), .B2(n6534), .ZN(n6536)
         );
  INV_X1 U7549 ( .A(n6536), .ZN(n6538) );
  AOI22_X1 U7550 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6709), .B1(n6623), 
        .B2(n6548), .ZN(n6537) );
  OAI211_X1 U7551 ( .C1(n6706), .C2(n6580), .A(n6538), .B(n6537), .ZN(U3081)
         );
  OAI22_X1 U7552 ( .A1(n6703), .A2(n6540), .B1(n6700), .B2(n6539), .ZN(n6541)
         );
  INV_X1 U7553 ( .A(n6541), .ZN(n6544) );
  AOI22_X1 U7554 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6709), .B1(n6631), 
        .B2(n6542), .ZN(n6543) );
  OAI211_X1 U7555 ( .C1(n6706), .C2(n6583), .A(n6544), .B(n6543), .ZN(U3082)
         );
  OAI22_X1 U7556 ( .A1(n6702), .A2(n6546), .B1(n6700), .B2(n6545), .ZN(n6547)
         );
  INV_X1 U7557 ( .A(n6547), .ZN(n6550) );
  AOI22_X1 U7558 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6709), .B1(n6639), 
        .B2(n6548), .ZN(n6549) );
  OAI211_X1 U7559 ( .C1(n6706), .C2(n6590), .A(n6550), .B(n6549), .ZN(U3083)
         );
  OR2_X1 U7560 ( .A1(n6551), .A2(n6677), .ZN(n6559) );
  NAND2_X1 U7561 ( .A1(n6553), .A2(n6552), .ZN(n6555) );
  INV_X1 U7562 ( .A(n6584), .ZN(n6554) );
  NAND2_X1 U7563 ( .A1(n6555), .A2(n6554), .ZN(n6561) );
  AOI22_X1 U7564 ( .A1(n6585), .A2(n6558), .B1(n6557), .B2(n6584), .ZN(n6565)
         );
  INV_X1 U7565 ( .A(n6559), .ZN(n6562) );
  AOI22_X1 U7566 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6587), .B1(n6563), 
        .B2(n6586), .ZN(n6564) );
  OAI211_X1 U7567 ( .C1(n6591), .C2(n6566), .A(n6565), .B(n6564), .ZN(U3108)
         );
  AOI22_X1 U7568 ( .A1(n6585), .A2(n6596), .B1(n6592), .B2(n6584), .ZN(n6568)
         );
  AOI22_X1 U7569 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6587), .B1(n6595), 
        .B2(n6586), .ZN(n6567) );
  OAI211_X1 U7570 ( .C1(n6591), .C2(n6705), .A(n6568), .B(n6567), .ZN(U3109)
         );
  AOI22_X1 U7571 ( .A1(n6586), .A2(n6602), .B1(n6600), .B2(n6584), .ZN(n6570)
         );
  AOI22_X1 U7572 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6587), .B1(n6603), 
        .B2(n6585), .ZN(n6569) );
  OAI211_X1 U7573 ( .C1(n6591), .C2(n6571), .A(n6570), .B(n6569), .ZN(U3110)
         );
  AOI22_X1 U7574 ( .A1(n6586), .A2(n6609), .B1(n6607), .B2(n6584), .ZN(n6573)
         );
  AOI22_X1 U7575 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6587), .B1(n6610), 
        .B2(n6585), .ZN(n6572) );
  OAI211_X1 U7576 ( .C1(n6591), .C2(n6574), .A(n6573), .B(n6572), .ZN(U3111)
         );
  AOI22_X1 U7577 ( .A1(n6585), .A2(n6617), .B1(n6614), .B2(n6584), .ZN(n6576)
         );
  AOI22_X1 U7578 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6587), .B1(n6616), 
        .B2(n6586), .ZN(n6575) );
  OAI211_X1 U7579 ( .C1(n6591), .C2(n6577), .A(n6576), .B(n6575), .ZN(U3112)
         );
  AOI22_X1 U7580 ( .A1(n6585), .A2(n6624), .B1(n6621), .B2(n6584), .ZN(n6579)
         );
  AOI22_X1 U7581 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6587), .B1(n6623), 
        .B2(n6586), .ZN(n6578) );
  OAI211_X1 U7582 ( .C1(n6591), .C2(n6580), .A(n6579), .B(n6578), .ZN(U3113)
         );
  AOI22_X1 U7583 ( .A1(n6586), .A2(n6630), .B1(n6628), .B2(n6584), .ZN(n6582)
         );
  AOI22_X1 U7584 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6587), .B1(n6631), 
        .B2(n6585), .ZN(n6581) );
  OAI211_X1 U7585 ( .C1(n6591), .C2(n6583), .A(n6582), .B(n6581), .ZN(U3114)
         );
  AOI22_X1 U7586 ( .A1(n6585), .A2(n6641), .B1(n6635), .B2(n6584), .ZN(n6589)
         );
  AOI22_X1 U7587 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6587), .B1(n6639), 
        .B2(n6586), .ZN(n6588) );
  OAI211_X1 U7588 ( .C1(n6591), .C2(n6590), .A(n6589), .B(n6588), .ZN(U3115)
         );
  INV_X1 U7589 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6599) );
  AOI22_X1 U7590 ( .A1(n6638), .A2(n6593), .B1(n6636), .B2(n6592), .ZN(n6598)
         );
  AOI22_X1 U7591 ( .A1(n6642), .A2(n6596), .B1(n6640), .B2(n6595), .ZN(n6597)
         );
  OAI211_X1 U7592 ( .C1(n6646), .C2(n6599), .A(n6598), .B(n6597), .ZN(U3141)
         );
  INV_X1 U7593 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n6606) );
  AOI22_X1 U7594 ( .A1(n6638), .A2(n6601), .B1(n6636), .B2(n6600), .ZN(n6605)
         );
  AOI22_X1 U7595 ( .A1(n6642), .A2(n6603), .B1(n6640), .B2(n6602), .ZN(n6604)
         );
  OAI211_X1 U7596 ( .C1(n6646), .C2(n6606), .A(n6605), .B(n6604), .ZN(U3142)
         );
  INV_X1 U7597 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n6613) );
  AOI22_X1 U7598 ( .A1(n6638), .A2(n6608), .B1(n6636), .B2(n6607), .ZN(n6612)
         );
  AOI22_X1 U7599 ( .A1(n6642), .A2(n6610), .B1(n6640), .B2(n6609), .ZN(n6611)
         );
  OAI211_X1 U7600 ( .C1(n6646), .C2(n6613), .A(n6612), .B(n6611), .ZN(U3143)
         );
  INV_X1 U7601 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n6620) );
  AOI22_X1 U7602 ( .A1(n6638), .A2(n6615), .B1(n6636), .B2(n6614), .ZN(n6619)
         );
  AOI22_X1 U7603 ( .A1(n6642), .A2(n6617), .B1(n6640), .B2(n6616), .ZN(n6618)
         );
  OAI211_X1 U7604 ( .C1(n6646), .C2(n6620), .A(n6619), .B(n6618), .ZN(U3144)
         );
  INV_X1 U7605 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6627) );
  AOI22_X1 U7606 ( .A1(n6638), .A2(n6622), .B1(n6636), .B2(n6621), .ZN(n6626)
         );
  AOI22_X1 U7607 ( .A1(n6642), .A2(n6624), .B1(n6640), .B2(n6623), .ZN(n6625)
         );
  OAI211_X1 U7608 ( .C1(n6646), .C2(n6627), .A(n6626), .B(n6625), .ZN(U3145)
         );
  INV_X1 U7609 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n6634) );
  AOI22_X1 U7610 ( .A1(n6638), .A2(n6629), .B1(n6636), .B2(n6628), .ZN(n6633)
         );
  AOI22_X1 U7611 ( .A1(n6642), .A2(n6631), .B1(n6640), .B2(n6630), .ZN(n6632)
         );
  OAI211_X1 U7612 ( .C1(n6646), .C2(n6634), .A(n6633), .B(n6632), .ZN(U3146)
         );
  INV_X1 U7613 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n6645) );
  AOI22_X1 U7614 ( .A1(n6638), .A2(n6637), .B1(n6636), .B2(n6635), .ZN(n6644)
         );
  AOI22_X1 U7615 ( .A1(n6642), .A2(n6641), .B1(n6640), .B2(n6639), .ZN(n6643)
         );
  OAI211_X1 U7616 ( .C1(n6646), .C2(n6645), .A(n6644), .B(n6643), .ZN(U3147)
         );
  AOI21_X1 U7617 ( .B1(READY_N), .B2(n6657), .A(n6663), .ZN(n6656) );
  AOI211_X1 U7618 ( .C1(n6694), .C2(n6647), .A(STATE2_REG_0__SCAN_IN), .B(
        n6663), .ZN(n6648) );
  AOI211_X1 U7619 ( .C1(n6654), .C2(n6650), .A(n6649), .B(n6648), .ZN(n6651)
         );
  OAI221_X1 U7620 ( .B1(n6747), .B2(n6656), .C1(n6747), .C2(n6652), .A(n6651), 
        .ZN(U3148) );
  INV_X1 U7621 ( .A(n6653), .ZN(n6655) );
  AOI21_X1 U7622 ( .B1(n6655), .B2(n6692), .A(n6654), .ZN(n6662) );
  INV_X1 U7623 ( .A(n6656), .ZN(n6658) );
  NAND2_X1 U7624 ( .A1(n6747), .A2(n6657), .ZN(n6664) );
  NAND3_X1 U7625 ( .A1(n6658), .A2(STATE2_REG_1__SCAN_IN), .A3(n6664), .ZN(
        n6660) );
  AND2_X1 U7626 ( .A1(n6660), .A2(n6659), .ZN(n6661) );
  OAI21_X1 U7627 ( .B1(n6663), .B2(n6662), .A(n6661), .ZN(U3149) );
  OAI211_X1 U7628 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6692), .A(n6665), .B(
        n6664), .ZN(n6667) );
  OAI21_X1 U7629 ( .B1(n6694), .B2(n6667), .A(n6666), .ZN(U3150) );
  AOI211_X1 U7630 ( .C1(n6671), .C2(n6670), .A(n6669), .B(n6668), .ZN(n6673)
         );
  NOR2_X1 U7631 ( .A1(n6673), .A2(n6672), .ZN(n6679) );
  OAI22_X1 U7632 ( .A1(n6677), .A2(n6676), .B1(n6675), .B2(n6674), .ZN(n6678)
         );
  OAI21_X1 U7633 ( .B1(n6679), .B2(n6678), .A(n6682), .ZN(n6680) );
  OAI21_X1 U7634 ( .B1(n6682), .B2(n6681), .A(n6680), .ZN(U3462) );
  AOI21_X1 U7635 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6683) );
  AOI22_X1 U7636 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6683), .B2(n6815), .ZN(n6685) );
  INV_X1 U7637 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6684) );
  AOI22_X1 U7638 ( .A1(n6686), .A2(n6685), .B1(n6684), .B2(n6688), .ZN(U3468)
         );
  INV_X1 U7639 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6689) );
  NOR2_X1 U7640 ( .A1(n6688), .A2(REIP_REG_1__SCAN_IN), .ZN(n6687) );
  AOI22_X1 U7641 ( .A1(n6689), .A2(n6688), .B1(n6797), .B2(n6687), .ZN(U3469)
         );
  AOI211_X1 U7642 ( .C1(n6331), .C2(n6692), .A(n6691), .B(n6690), .ZN(n6698)
         );
  OAI211_X1 U7643 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4071), .A(n6693), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6695) );
  AOI21_X1 U7644 ( .B1(n6695), .B2(STATE2_REG_0__SCAN_IN), .A(n6694), .ZN(
        n6697) );
  NAND2_X1 U7645 ( .A1(n6698), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6696) );
  OAI21_X1 U7646 ( .B1(n6698), .B2(n6697), .A(n6696), .ZN(U3472) );
  OAI22_X1 U7647 ( .A1(n6702), .A2(n6701), .B1(n6700), .B2(n6699), .ZN(n6708)
         );
  OAI22_X1 U7648 ( .A1(n6706), .A2(n6705), .B1(n6704), .B2(n6703), .ZN(n6707)
         );
  AOI211_X1 U7649 ( .C1(INSTQUEUE_REG_7__1__SCAN_IN), .C2(n6709), .A(n6708), 
        .B(n6707), .ZN(n6862) );
  NAND4_X1 U7650 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(
        INSTQUEUE_REG_5__7__SCAN_IN), .A3(INSTQUEUE_REG_7__7__SCAN_IN), .A4(
        INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6719) );
  NOR4_X1 U7651 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(
        INSTQUEUE_REG_15__0__SCAN_IN), .A3(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .A4(ADDRESS_REG_28__SCAN_IN), .ZN(n6712) );
  NOR3_X1 U7652 ( .A1(DATAI_11_), .A2(DATAO_REG_4__SCAN_IN), .A3(n6738), .ZN(
        n6711) );
  INV_X1 U7653 ( .A(DATAI_14_), .ZN(n6762) );
  NOR4_X1 U7654 ( .A1(EAX_REG_0__SCAN_IN), .A2(ADDRESS_REG_3__SCAN_IN), .A3(
        n6754), .A4(n6762), .ZN(n6710) );
  NAND4_X1 U7655 ( .A1(n6712), .A2(LWORD_REG_4__SCAN_IN), .A3(n6711), .A4(
        n6710), .ZN(n6718) );
  NAND4_X1 U7656 ( .A1(EAX_REG_21__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        UWORD_REG_5__SCAN_IN), .A4(DATAO_REG_19__SCAN_IN), .ZN(n6717) );
  NOR4_X1 U7657 ( .A1(EBX_REG_24__SCAN_IN), .A2(EBX_REG_19__SCAN_IN), .A3(
        DATAO_REG_27__SCAN_IN), .A4(n6777), .ZN(n6715) );
  NOR3_X1 U7658 ( .A1(DATAI_31_), .A2(ADDRESS_REG_25__SCAN_IN), .A3(n6780), 
        .ZN(n6714) );
  NOR4_X1 U7659 ( .A1(EBX_REG_20__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        n6816), .A4(n6797), .ZN(n6713) );
  NAND4_X1 U7660 ( .A1(n6715), .A2(UWORD_REG_10__SCAN_IN), .A3(n6714), .A4(
        n6713), .ZN(n6716) );
  NOR4_X1 U7661 ( .A1(n6719), .A2(n6718), .A3(n6717), .A4(n6716), .ZN(n6860)
         );
  INV_X1 U7662 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n6832) );
  NAND4_X1 U7663 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(
        INSTQUEUE_REG_5__5__SCAN_IN), .A3(INSTQUEUE_REG_14__5__SCAN_IN), .A4(
        n6832), .ZN(n6720) );
  NOR4_X1 U7664 ( .A1(n6157), .A2(n6752), .A3(n6721), .A4(n6720), .ZN(n6724)
         );
  INV_X1 U7665 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n6775) );
  NOR4_X1 U7666 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(
        INSTQUEUE_REG_3__4__SCAN_IN), .A3(INSTQUEUE_REG_2__1__SCAN_IN), .A4(
        n6775), .ZN(n6722) );
  NAND4_X1 U7667 ( .A1(n6724), .A2(n6723), .A3(n6722), .A4(n6831), .ZN(n6730)
         );
  NAND4_X1 U7668 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(DATAO_REG_0__SCAN_IN), 
        .A3(n6800), .A4(n6844), .ZN(n6729) );
  NAND4_X1 U7669 ( .A1(EAX_REG_27__SCAN_IN), .A2(DATAI_15_), .A3(n4969), .A4(
        n6847), .ZN(n6728) );
  NOR4_X1 U7670 ( .A1(LWORD_REG_14__SCAN_IN), .A2(EAX_REG_13__SCAN_IN), .A3(
        DATAO_REG_6__SCAN_IN), .A4(n6795), .ZN(n6726) );
  NAND4_X1 U7671 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6726), .A3(ADS_N_REG_SCAN_IN), 
        .A4(n6725), .ZN(n6727) );
  NOR4_X1 U7672 ( .A1(n6730), .A2(n6729), .A3(n6728), .A4(n6727), .ZN(n6859)
         );
  AOI22_X1 U7673 ( .A1(n6732), .A2(keyinput59), .B1(n4877), .B2(keyinput52), 
        .ZN(n6731) );
  OAI221_X1 U7674 ( .B1(n6732), .B2(keyinput59), .C1(n4877), .C2(keyinput52), 
        .A(n6731), .ZN(n6744) );
  INV_X1 U7675 ( .A(DATAI_11_), .ZN(n6735) );
  AOI22_X1 U7676 ( .A1(n6735), .A2(keyinput3), .B1(keyinput10), .B2(n6734), 
        .ZN(n6733) );
  OAI221_X1 U7677 ( .B1(n6735), .B2(keyinput3), .C1(n6734), .C2(keyinput10), 
        .A(n6733), .ZN(n6743) );
  AOI22_X1 U7678 ( .A1(n6737), .A2(keyinput49), .B1(n3060), .B2(keyinput37), 
        .ZN(n6736) );
  OAI221_X1 U7679 ( .B1(n6737), .B2(keyinput49), .C1(n3060), .C2(keyinput37), 
        .A(n6736), .ZN(n6742) );
  XOR2_X1 U7680 ( .A(n6738), .B(keyinput55), .Z(n6740) );
  XNOR2_X1 U7681 ( .A(INSTQUEUE_REG_3__4__SCAN_IN), .B(keyinput18), .ZN(n6739)
         );
  NAND2_X1 U7682 ( .A1(n6740), .A2(n6739), .ZN(n6741) );
  NOR4_X1 U7683 ( .A1(n6744), .A2(n6743), .A3(n6742), .A4(n6741), .ZN(n6792)
         );
  AOI22_X1 U7684 ( .A1(n6747), .A2(keyinput33), .B1(keyinput63), .B2(n6746), 
        .ZN(n6745) );
  OAI221_X1 U7685 ( .B1(n6747), .B2(keyinput33), .C1(n6746), .C2(keyinput63), 
        .A(n6745), .ZN(n6759) );
  AOI22_X1 U7686 ( .A1(n6157), .A2(keyinput2), .B1(keyinput8), .B2(n6749), 
        .ZN(n6748) );
  OAI221_X1 U7687 ( .B1(n6157), .B2(keyinput2), .C1(n6749), .C2(keyinput8), 
        .A(n6748), .ZN(n6758) );
  INV_X1 U7688 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6751) );
  AOI22_X1 U7689 ( .A1(n6752), .A2(keyinput6), .B1(n6751), .B2(keyinput56), 
        .ZN(n6750) );
  OAI221_X1 U7690 ( .B1(n6752), .B2(keyinput6), .C1(n6751), .C2(keyinput56), 
        .A(n6750), .ZN(n6757) );
  INV_X1 U7691 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6755) );
  AOI22_X1 U7692 ( .A1(n6755), .A2(keyinput1), .B1(keyinput28), .B2(n6754), 
        .ZN(n6753) );
  OAI221_X1 U7693 ( .B1(n6755), .B2(keyinput1), .C1(n6754), .C2(keyinput28), 
        .A(n6753), .ZN(n6756) );
  NOR4_X1 U7694 ( .A1(n6759), .A2(n6758), .A3(n6757), .A4(n6756), .ZN(n6791)
         );
  INV_X1 U7695 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n6761) );
  AOI22_X1 U7696 ( .A1(n6762), .A2(keyinput30), .B1(keyinput35), .B2(n6761), 
        .ZN(n6760) );
  OAI221_X1 U7697 ( .B1(n6762), .B2(keyinput30), .C1(n6761), .C2(keyinput35), 
        .A(n6760), .ZN(n6773) );
  INV_X1 U7698 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6764) );
  AOI22_X1 U7699 ( .A1(n6764), .A2(keyinput15), .B1(n4900), .B2(keyinput23), 
        .ZN(n6763) );
  OAI221_X1 U7700 ( .B1(n6764), .B2(keyinput15), .C1(n4900), .C2(keyinput23), 
        .A(n6763), .ZN(n6772) );
  AOI22_X1 U7701 ( .A1(n4881), .A2(keyinput43), .B1(keyinput27), .B2(n6766), 
        .ZN(n6765) );
  OAI221_X1 U7702 ( .B1(n4881), .B2(keyinput43), .C1(n6766), .C2(keyinput27), 
        .A(n6765), .ZN(n6771) );
  AOI22_X1 U7703 ( .A1(n6769), .A2(keyinput29), .B1(n6768), .B2(keyinput62), 
        .ZN(n6767) );
  OAI221_X1 U7704 ( .B1(n6769), .B2(keyinput29), .C1(n6768), .C2(keyinput62), 
        .A(n6767), .ZN(n6770) );
  NOR4_X1 U7705 ( .A1(n6773), .A2(n6772), .A3(n6771), .A4(n6770), .ZN(n6790)
         );
  AOI22_X1 U7706 ( .A1(n6775), .A2(keyinput7), .B1(keyinput5), .B2(n4922), 
        .ZN(n6774) );
  OAI221_X1 U7707 ( .B1(n6775), .B2(keyinput7), .C1(n4922), .C2(keyinput5), 
        .A(n6774), .ZN(n6788) );
  AOI22_X1 U7708 ( .A1(n6778), .A2(keyinput42), .B1(keyinput46), .B2(n6777), 
        .ZN(n6776) );
  OAI221_X1 U7709 ( .B1(n6778), .B2(keyinput42), .C1(n6777), .C2(keyinput46), 
        .A(n6776), .ZN(n6787) );
  AOI22_X1 U7710 ( .A1(n6781), .A2(keyinput20), .B1(n6780), .B2(keyinput13), 
        .ZN(n6779) );
  OAI221_X1 U7711 ( .B1(n6781), .B2(keyinput20), .C1(n6780), .C2(keyinput13), 
        .A(n6779), .ZN(n6786) );
  AOI22_X1 U7712 ( .A1(n6784), .A2(keyinput50), .B1(keyinput16), .B2(n6783), 
        .ZN(n6782) );
  OAI221_X1 U7713 ( .B1(n6784), .B2(keyinput50), .C1(n6783), .C2(keyinput16), 
        .A(n6782), .ZN(n6785) );
  NOR4_X1 U7714 ( .A1(n6788), .A2(n6787), .A3(n6786), .A4(n6785), .ZN(n6789)
         );
  NAND4_X1 U7715 ( .A1(n6792), .A2(n6791), .A3(n6790), .A4(n6789), .ZN(n6858)
         );
  INV_X1 U7716 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n6794) );
  AOI22_X1 U7717 ( .A1(n6795), .A2(keyinput26), .B1(n6794), .B2(keyinput41), 
        .ZN(n6793) );
  OAI221_X1 U7718 ( .B1(n6795), .B2(keyinput26), .C1(n6794), .C2(keyinput41), 
        .A(n6793), .ZN(n6808) );
  AOI22_X1 U7719 ( .A1(n6798), .A2(keyinput47), .B1(keyinput0), .B2(n6797), 
        .ZN(n6796) );
  OAI221_X1 U7720 ( .B1(n6798), .B2(keyinput47), .C1(n6797), .C2(keyinput0), 
        .A(n6796), .ZN(n6807) );
  AOI22_X1 U7721 ( .A1(n6801), .A2(keyinput9), .B1(n6800), .B2(keyinput32), 
        .ZN(n6799) );
  OAI221_X1 U7722 ( .B1(n6801), .B2(keyinput9), .C1(n6800), .C2(keyinput32), 
        .A(n6799), .ZN(n6806) );
  AOI22_X1 U7723 ( .A1(n6804), .A2(keyinput31), .B1(keyinput36), .B2(n6803), 
        .ZN(n6802) );
  OAI221_X1 U7724 ( .B1(n6804), .B2(keyinput31), .C1(n6803), .C2(keyinput36), 
        .A(n6802), .ZN(n6805) );
  NOR4_X1 U7725 ( .A1(n6808), .A2(n6807), .A3(n6806), .A4(n6805), .ZN(n6856)
         );
  INV_X1 U7726 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n6810) );
  AOI22_X1 U7727 ( .A1(n6810), .A2(keyinput17), .B1(keyinput40), .B2(n4370), 
        .ZN(n6809) );
  OAI221_X1 U7728 ( .B1(n6810), .B2(keyinput17), .C1(n4370), .C2(keyinput40), 
        .A(n6809), .ZN(n6823) );
  AOI22_X1 U7729 ( .A1(n6813), .A2(keyinput53), .B1(keyinput51), .B2(n6812), 
        .ZN(n6811) );
  OAI221_X1 U7730 ( .B1(n6813), .B2(keyinput53), .C1(n6812), .C2(keyinput51), 
        .A(n6811), .ZN(n6822) );
  AOI22_X1 U7731 ( .A1(n6816), .A2(keyinput60), .B1(n6815), .B2(keyinput61), 
        .ZN(n6814) );
  OAI221_X1 U7732 ( .B1(n6816), .B2(keyinput60), .C1(n6815), .C2(keyinput61), 
        .A(n6814), .ZN(n6821) );
  AOI22_X1 U7733 ( .A1(n6819), .A2(keyinput38), .B1(n6818), .B2(keyinput48), 
        .ZN(n6817) );
  OAI221_X1 U7734 ( .B1(n6819), .B2(keyinput38), .C1(n6818), .C2(keyinput48), 
        .A(n6817), .ZN(n6820) );
  NOR4_X1 U7735 ( .A1(n6823), .A2(n6822), .A3(n6821), .A4(n6820), .ZN(n6855)
         );
  INV_X1 U7736 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6825) );
  AOI22_X1 U7737 ( .A1(n6826), .A2(keyinput44), .B1(n6825), .B2(keyinput54), 
        .ZN(n6824) );
  OAI221_X1 U7738 ( .B1(n6826), .B2(keyinput44), .C1(n6825), .C2(keyinput54), 
        .A(n6824), .ZN(n6838) );
  INV_X1 U7739 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n6829) );
  AOI22_X1 U7740 ( .A1(n6829), .A2(keyinput34), .B1(keyinput12), .B2(n6828), 
        .ZN(n6827) );
  OAI221_X1 U7741 ( .B1(n6829), .B2(keyinput34), .C1(n6828), .C2(keyinput12), 
        .A(n6827), .ZN(n6837) );
  AOI22_X1 U7742 ( .A1(n6832), .A2(keyinput4), .B1(keyinput11), .B2(n6831), 
        .ZN(n6830) );
  OAI221_X1 U7743 ( .B1(n6832), .B2(keyinput4), .C1(n6831), .C2(keyinput11), 
        .A(n6830), .ZN(n6836) );
  XNOR2_X1 U7744 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .B(keyinput14), .ZN(n6834) );
  XNOR2_X1 U7745 ( .A(STATE2_REG_1__SCAN_IN), .B(keyinput19), .ZN(n6833) );
  NAND2_X1 U7746 ( .A1(n6834), .A2(n6833), .ZN(n6835) );
  NOR4_X1 U7747 ( .A1(n6838), .A2(n6837), .A3(n6836), .A4(n6835), .ZN(n6854)
         );
  AOI22_X1 U7748 ( .A1(n6841), .A2(keyinput45), .B1(n6840), .B2(keyinput24), 
        .ZN(n6839) );
  OAI221_X1 U7749 ( .B1(n6841), .B2(keyinput45), .C1(n6840), .C2(keyinput24), 
        .A(n6839), .ZN(n6852) );
  AOI22_X1 U7750 ( .A1(n6844), .A2(keyinput21), .B1(keyinput58), .B2(n6843), 
        .ZN(n6842) );
  OAI221_X1 U7751 ( .B1(n6844), .B2(keyinput21), .C1(n6843), .C2(keyinput58), 
        .A(n6842), .ZN(n6851) );
  AOI22_X1 U7752 ( .A1(n3911), .A2(keyinput22), .B1(n4969), .B2(keyinput25), 
        .ZN(n6845) );
  OAI221_X1 U7753 ( .B1(n3911), .B2(keyinput22), .C1(n4969), .C2(keyinput25), 
        .A(n6845), .ZN(n6850) );
  AOI22_X1 U7754 ( .A1(n6848), .A2(keyinput57), .B1(keyinput39), .B2(n6847), 
        .ZN(n6846) );
  OAI221_X1 U7755 ( .B1(n6848), .B2(keyinput57), .C1(n6847), .C2(keyinput39), 
        .A(n6846), .ZN(n6849) );
  NOR4_X1 U7756 ( .A1(n6852), .A2(n6851), .A3(n6850), .A4(n6849), .ZN(n6853)
         );
  NAND4_X1 U7757 ( .A1(n6856), .A2(n6855), .A3(n6854), .A4(n6853), .ZN(n6857)
         );
  AOI211_X1 U7758 ( .C1(n6860), .C2(n6859), .A(n6858), .B(n6857), .ZN(n6861)
         );
  XNOR2_X1 U7759 ( .A(n6862), .B(n6861), .ZN(U3077) );
  AND4_X1 U4286 ( .A1(n3190), .A2(n3189), .A3(n3188), .A4(n3187), .ZN(n3201)
         );
  NAND2_X1 U4441 ( .A1(n3404), .A2(n3403), .ZN(n3490) );
  AND2_X2 U5100 ( .A1(n3328), .A2(n3322), .ZN(n4527) );
  NAND2_X1 U4087 ( .A1(n5779), .A2(n3125), .ZN(n3121) );
  AND4_X1 U4290 ( .A1(n3194), .A2(n3193), .A3(n3192), .A4(n3191), .ZN(n3200)
         );
  AND2_X2 U3512 ( .A1(n4506), .A2(n4719), .ZN(n3263) );
  CLKBUF_X1 U3692 ( .A(n3282), .Z(n3986) );
  CLKBUF_X1 U3807 ( .A(n4245), .Z(n6671) );
endmodule

