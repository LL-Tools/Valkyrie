

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4402, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9920, n9921, n9922, n9923, n9924, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10615;

  AOI211_X1 U4907 ( .C1(n9161), .C2(n9148), .A(n8454), .B(n8453), .ZN(n8455)
         );
  AND2_X1 U4908 ( .A1(n9567), .A2(n9566), .ZN(n9793) );
  NAND2_X1 U4909 ( .A1(n9594), .A2(n9585), .ZN(n8356) );
  AOI21_X1 U4910 ( .B1(n8959), .B2(n5834), .A(n5751), .ZN(n8735) );
  OR2_X2 U4911 ( .A1(n9177), .A2(n8964), .ZN(n8730) );
  AND2_X1 U4912 ( .A1(n5739), .A2(n5738), .ZN(n8964) );
  INV_X1 U4913 ( .A(n6901), .ZN(n6916) );
  BUF_X2 U4914 ( .A(n4411), .Z(n6901) );
  AND4_X1 U4915 ( .A1(n5974), .A2(n5973), .A3(n5972), .A4(n5971), .ZN(n10139)
         );
  XNOR2_X1 U4916 ( .A(n6711), .B(n7768), .ZN(n6564) );
  INV_X1 U4917 ( .A(n6012), .ZN(n6106) );
  BUF_X2 U4918 ( .A(n5294), .Z(n8398) );
  XNOR2_X1 U4919 ( .A(n5794), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8765) );
  NAND2_X1 U4920 ( .A1(n5330), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5382) );
  NAND2_X1 U4921 ( .A1(n5228), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5300) );
  INV_X1 U4922 ( .A(n9284), .ZN(n4402) );
  INV_X2 U4923 ( .A(n4402), .ZN(P2_U3152) );
  INV_X1 U4924 ( .A(P2_STATE_REG_SCAN_IN), .ZN(n9284) );
  INV_X2 U4926 ( .A(n10615), .ZN(n4405) );
  INV_X1 U4928 ( .A(n8746), .ZN(n8755) );
  NAND2_X1 U4929 ( .A1(n5588), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U4930 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5229) );
  NOR2_X1 U4931 ( .A1(n7616), .A2(n6953), .ZN(n6722) );
  INV_X2 U4932 ( .A(n4413), .ZN(n6910) );
  INV_X1 U4933 ( .A(n9917), .ZN(n5872) );
  INV_X1 U4934 ( .A(n6467), .ZN(n6114) );
  NAND2_X1 U4935 ( .A1(n7922), .A2(n6376), .ZN(n8032) );
  INV_X1 U4936 ( .A(n8608), .ZN(n8600) );
  AND2_X1 U4937 ( .A1(n5731), .A2(n5713), .ZN(n8993) );
  OR3_X2 U4938 ( .A1(n5772), .A2(n5771), .A3(n5770), .ZN(n8451) );
  NAND2_X1 U4939 ( .A1(n8730), .A2(n8731), .ZN(n8982) );
  INV_X1 U4940 ( .A(n9008), .ZN(n9048) );
  INV_X1 U4941 ( .A(n8765), .ZN(n5811) );
  INV_X1 U4942 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9271) );
  INV_X2 U4943 ( .A(n7366), .ZN(n8568) );
  AND4_X1 U4944 ( .A1(n5367), .A2(n5366), .A3(n5365), .A4(n5364), .ZN(n7884)
         );
  INV_X1 U4945 ( .A(n5122), .ZN(n8591) );
  INV_X1 U4946 ( .A(n10222), .ZN(n7263) );
  NAND2_X1 U4947 ( .A1(n6170), .A2(n6169), .ZN(n6260) );
  AND4_X1 U4948 ( .A1(n5986), .A2(n5985), .A3(n5984), .A4(n5983), .ZN(n9730)
         );
  NAND4_X1 U4949 ( .A1(n5209), .A2(n5208), .A3(n5207), .A4(n5206), .ZN(n8790)
         );
  AND2_X1 U4950 ( .A1(n5223), .A2(n5222), .ZN(n10227) );
  INV_X2 U4951 ( .A(n5064), .ZN(n9711) );
  CLKBUF_X3 U4952 ( .A(n6742), .Z(n4411) );
  OR2_X2 U4953 ( .A1(n5451), .A2(n5450), .ZN(n5453) );
  NAND2_X2 U4954 ( .A1(n4907), .A2(n7567), .ZN(n7647) );
  NAND2_X2 U4955 ( .A1(n6821), .A2(n9288), .ZN(n9329) );
  NAND2_X2 U4956 ( .A1(n6820), .A2(n6819), .ZN(n9288) );
  XNOR2_X2 U4957 ( .A(n5869), .B(n4549), .ZN(n9917) );
  INV_X2 U4958 ( .A(n5731), .ZN(n5730) );
  INV_X2 U4959 ( .A(n5935), .ZN(n6469) );
  NAND2_X1 U4960 ( .A1(n6729), .A2(n10078), .ZN(n10055) );
  AND2_X2 U4961 ( .A1(n5097), .A2(n5099), .ZN(n5194) );
  XNOR2_X2 U4962 ( .A(n5095), .B(n5094), .ZN(n5099) );
  AOI21_X1 U4963 ( .B1(n6402), .B2(n4421), .A(n4476), .ZN(n4690) );
  NAND2_X4 U4964 ( .A1(n4572), .A2(n4570), .ZN(n5244) );
  NAND3_X2 U4965 ( .A1(n9478), .A2(n4574), .A3(n4573), .ZN(n4572) );
  INV_X1 U4966 ( .A(n5193), .ZN(n4406) );
  NAND2_X2 U4967 ( .A1(n5730), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5772) );
  NAND2_X2 U4968 ( .A1(n9272), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5093) );
  NAND2_X2 U4969 ( .A1(n9027), .A2(n9026), .ZN(n9025) );
  NOR2_X2 U4970 ( .A1(n6476), .A2(n6475), .ZN(n6481) );
  NAND2_X2 U4971 ( .A1(n5685), .A2(n5684), .ZN(n5704) );
  OR2_X2 U4974 ( .A1(n6486), .A2(n6483), .ZN(n6622) );
  AND2_X2 U4975 ( .A1(n8002), .A2(n5042), .ZN(n9739) );
  OAI21_X2 U4976 ( .B1(n10027), .B2(n10035), .A(n5938), .ZN(n7618) );
  OR2_X2 U4977 ( .A1(n6287), .A2(n6046), .ZN(n6244) );
  NOR2_X2 U4978 ( .A1(n6238), .A2(P1_IR_REG_19__SCAN_IN), .ZN(n6287) );
  NAND2_X2 U4979 ( .A1(n9089), .A2(n8420), .ZN(n9072) );
  NAND2_X2 U4980 ( .A1(n4909), .A2(n4908), .ZN(n9089) );
  OR2_X2 U4981 ( .A1(n5975), .A2(n10139), .ZN(n7922) );
  AOI21_X2 U4982 ( .B1(n8943), .B2(n9138), .A(n8942), .ZN(n9170) );
  NAND2_X2 U4983 ( .A1(n8426), .A2(n8424), .ZN(n8428) );
  AND2_X2 U4984 ( .A1(n7356), .A2(n7412), .ZN(n7871) );
  OAI21_X2 U4985 ( .B1(n5075), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5794) );
  AND2_X2 U4986 ( .A1(n6243), .A2(n6242), .ZN(n6264) );
  NOR2_X2 U4987 ( .A1(n8789), .A2(n7412), .ZN(n8616) );
  NAND2_X2 U4988 ( .A1(n5587), .A2(n5586), .ZN(n9211) );
  NAND2_X2 U4989 ( .A1(n6023), .A2(n6022), .ZN(n9880) );
  NAND2_X2 U4990 ( .A1(n8088), .A2(n8087), .ZN(n8132) );
  NAND2_X2 U4991 ( .A1(n7788), .A2(n4426), .ZN(n8088) );
  OAI21_X4 U4992 ( .B1(n7470), .B2(n7471), .A(n6760), .ZN(n7475) );
  NAND2_X2 U4993 ( .A1(n4946), .A2(n4945), .ZN(n7470) );
  NOR3_X2 U4994 ( .A1(n9043), .A2(n9006), .A3(n9057), .ZN(n9045) );
  XNOR2_X2 U4995 ( .A(n8435), .B(n4937), .ZN(n9165) );
  NAND2_X2 U4996 ( .A1(n8944), .A2(n8433), .ZN(n8435) );
  OR2_X1 U4997 ( .A1(n9321), .A2(n9319), .ZN(n4962) );
  XNOR2_X1 U4998 ( .A(n5698), .B(n5696), .ZN(n8513) );
  OAI21_X1 U4999 ( .B1(n8523), .B2(n4536), .A(n4533), .ZN(n5698) );
  AND3_X1 U5000 ( .A1(n7871), .A2(n4843), .A3(n4842), .ZN(n7564) );
  INV_X2 U5001 ( .A(n9144), .ZN(n4407) );
  NAND2_X1 U5002 ( .A1(n9116), .A2(n9115), .ZN(n7349) );
  AND2_X1 U5003 ( .A1(n6363), .A2(n6580), .ZN(n10035) );
  OAI22_X1 U5004 ( .A1(n10043), .A2(n4413), .B1(n7632), .B2(n6748), .ZN(n6749)
         );
  AND2_X1 U5005 ( .A1(n4948), .A2(n4951), .ZN(n6958) );
  NAND2_X2 U5006 ( .A1(n8624), .A2(n8628), .ZN(n7345) );
  INV_X1 U5007 ( .A(n10082), .ZN(n7721) );
  INV_X1 U5008 ( .A(n5926), .ZN(n10096) );
  AND4_X1 U5009 ( .A1(n6018), .A2(n6017), .A3(n6016), .A4(n6015), .ZN(n9876)
         );
  INV_X1 U5010 ( .A(n8790), .ZN(n4906) );
  INV_X1 U5011 ( .A(n6722), .ZN(n6753) );
  CLKBUF_X2 U5012 ( .A(n5204), .Z(n7049) );
  NAND2_X2 U5013 ( .A1(n5811), .A2(n8600), .ZN(n8595) );
  NAND2_X1 U5014 ( .A1(n5868), .A2(n5867), .ZN(n8413) );
  BUF_X1 U5015 ( .A(n6267), .Z(n4412) );
  XNOR2_X1 U5016 ( .A(n5027), .B(P1_IR_REG_27__SCAN_IN), .ZN(n6616) );
  CLKBUF_X2 U5017 ( .A(n5318), .Z(n6344) );
  INV_X2 U5018 ( .A(n5244), .ZN(n5291) );
  INV_X2 U5019 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5134) );
  NOR2_X1 U5020 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5854) );
  OAI211_X1 U5021 ( .C1(n8340), .C2(n6236), .A(n9764), .B(n4468), .ZN(n8404)
         );
  NAND2_X1 U5022 ( .A1(n4793), .A2(n6235), .ZN(n9764) );
  NOR2_X1 U5023 ( .A1(n8382), .A2(n8381), .ZN(n9299) );
  NAND2_X1 U5024 ( .A1(n4624), .A2(n4623), .ZN(n8382) );
  NAND2_X1 U5025 ( .A1(n4967), .A2(n4965), .ZN(n4624) );
  NAND2_X1 U5026 ( .A1(n4962), .A2(n4961), .ZN(n4623) );
  AND2_X1 U5027 ( .A1(n4651), .A2(n4650), .ZN(n9009) );
  NAND2_X1 U5028 ( .A1(n4542), .A2(n4541), .ZN(n9591) );
  AND2_X1 U5029 ( .A1(n9541), .A2(n6440), .ZN(n8361) );
  AND2_X1 U5030 ( .A1(n9015), .A2(n4855), .ZN(n4854) );
  NAND2_X1 U5031 ( .A1(n6127), .A2(n6126), .ZN(n9620) );
  NAND2_X1 U5032 ( .A1(n9515), .A2(n9520), .ZN(n9517) );
  NAND2_X1 U5033 ( .A1(n8317), .A2(n4927), .ZN(n4924) );
  NAND2_X1 U5034 ( .A1(n5014), .A2(n5011), .ZN(n9593) );
  NAND2_X1 U5035 ( .A1(n6213), .A2(n6212), .ZN(n8350) );
  NAND2_X1 U5036 ( .A1(n9637), .A2(n5007), .ZN(n5014) );
  NAND2_X1 U5037 ( .A1(n4779), .A2(n4778), .ZN(n9634) );
  NAND2_X1 U5038 ( .A1(n5729), .A2(n5728), .ZN(n9177) );
  AOI21_X1 U5039 ( .B1(n5013), .B2(n5016), .A(n5012), .ZN(n5011) );
  OR2_X1 U5040 ( .A1(n8978), .A2(n5733), .ZN(n5739) );
  OAI21_X1 U5041 ( .B1(n9694), .B2(n4579), .A(n4575), .ZN(n9637) );
  AND2_X1 U5042 ( .A1(n9658), .A2(n4482), .ZN(n9610) );
  NAND2_X2 U5043 ( .A1(n8319), .A2(n8323), .ZN(n8393) );
  INV_X1 U5044 ( .A(n6415), .ZN(n5012) );
  XNOR2_X1 U5045 ( .A(n5704), .B(n5699), .ZN(n6158) );
  AND2_X1 U5046 ( .A1(n5663), .A2(n5662), .ZN(n9036) );
  INV_X1 U5047 ( .A(n6859), .ZN(n9823) );
  OR2_X1 U5048 ( .A1(n9716), .A2(n9689), .ZN(n5059) );
  NAND2_X1 U5049 ( .A1(n5623), .A2(n5622), .ZN(n9201) );
  NAND2_X1 U5050 ( .A1(n4616), .A2(n4420), .ZN(n4618) );
  NAND2_X1 U5051 ( .A1(n4531), .A2(n4530), .ZN(n7441) );
  NAND2_X1 U5052 ( .A1(n6140), .A2(n6139), .ZN(n9817) );
  NOR2_X1 U5053 ( .A1(n4968), .A2(n4617), .ZN(n4615) );
  OAI21_X1 U5054 ( .B1(n5656), .B2(n5655), .A(n5654), .ZN(n5683) );
  AOI21_X1 U5055 ( .B1(n8068), .B2(n6019), .A(n4437), .ZN(n8051) );
  OAI21_X1 U5056 ( .B1(n7998), .B2(n6255), .A(n6254), .ZN(n7923) );
  NAND2_X1 U5057 ( .A1(n5470), .A2(n5469), .ZN(n9226) );
  OR2_X1 U5058 ( .A1(n5046), .A2(n6253), .ZN(n6254) );
  NAND2_X1 U5059 ( .A1(n5506), .A2(n5505), .ZN(n8279) );
  NAND2_X1 U5060 ( .A1(n6052), .A2(n6051), .ZN(n9864) );
  NAND2_X1 U5061 ( .A1(n10036), .A2(n6363), .ZN(n7621) );
  NAND2_X1 U5062 ( .A1(n6064), .A2(n6063), .ZN(n9856) );
  OAI21_X1 U5063 ( .B1(n10034), .B2(n4996), .A(n4994), .ZN(n7998) );
  NAND2_X1 U5064 ( .A1(n5520), .A2(n5519), .ZN(n8127) );
  NAND2_X1 U5065 ( .A1(n10034), .A2(n10035), .ZN(n10036) );
  NAND2_X2 U5066 ( .A1(n7601), .A2(n9124), .ZN(n9144) );
  INV_X1 U5067 ( .A(n5589), .ZN(n5588) );
  NAND2_X1 U5068 ( .A1(n6011), .A2(n6010), .ZN(n9888) );
  NAND2_X1 U5069 ( .A1(n4701), .A2(n4700), .ZN(n9245) );
  AOI21_X1 U5070 ( .B1(n7920), .B2(n7994), .A(n5963), .ZN(n8029) );
  NOR2_X2 U5071 ( .A1(n10030), .A2(n7625), .ZN(n8002) );
  AND2_X1 U5072 ( .A1(n6741), .A2(n6739), .ZN(n7283) );
  NAND2_X1 U5073 ( .A1(n5967), .A2(n5966), .ZN(n5975) );
  AND2_X1 U5074 ( .A1(n6378), .A2(n6375), .ZN(n7924) );
  NAND2_X1 U5075 ( .A1(n5507), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5548) );
  XNOR2_X1 U5076 ( .A(n5323), .B(n5322), .ZN(n7028) );
  OR2_X1 U5077 ( .A1(n9730), .A2(n10144), .ZN(n6378) );
  NAND2_X1 U5078 ( .A1(n6958), .A2(n6960), .ZN(n6959) );
  AND2_X1 U5079 ( .A1(n4551), .A2(n4550), .ZN(n7632) );
  AND2_X2 U5080 ( .A1(n10179), .A2(n10178), .ZN(n10195) );
  INV_X1 U5081 ( .A(n5523), .ZN(n5507) );
  CLKBUF_X1 U5082 ( .A(n7265), .Z(n8791) );
  AND4_X1 U5083 ( .A1(n5933), .A2(n5932), .A3(n5931), .A4(n5930), .ZN(n7542)
         );
  NAND4_X2 U5084 ( .A1(n5876), .A2(n5875), .A3(n5874), .A4(n5873), .ZN(n9444)
         );
  AND2_X1 U5085 ( .A1(n7034), .A2(n4410), .ZN(n4949) );
  INV_X2 U5086 ( .A(n4432), .ZN(n6913) );
  NAND4_X1 U5087 ( .A1(n5172), .A2(n5171), .A3(n5170), .A4(n5169), .ZN(n7265)
         );
  AND2_X2 U5088 ( .A1(n4950), .A2(n6743), .ZN(n4432) );
  BUF_X2 U5089 ( .A(n6753), .Z(n4413) );
  AND3_X1 U5090 ( .A1(n5102), .A2(n5101), .A3(n5100), .ZN(n5103) );
  AND4_X1 U5091 ( .A1(n5898), .A2(n5897), .A3(n5896), .A4(n5895), .ZN(n6721)
         );
  AND3_X1 U5092 ( .A1(n5916), .A2(n5915), .A3(n5914), .ZN(n5918) );
  CLKBUF_X1 U5093 ( .A(n6722), .Z(n6756) );
  AOI21_X1 U5094 ( .B1(n5908), .B2(P2_DATAO_REG_1__SCAN_IN), .A(n5907), .ZN(
        n5028) );
  AND2_X2 U5095 ( .A1(n5811), .A2(n8601), .ZN(n8746) );
  BUF_X2 U5096 ( .A(n5194), .Z(n7047) );
  CLKBUF_X1 U5097 ( .A(n5913), .Z(n6349) );
  XNOR2_X1 U5098 ( .A(n6240), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U5099 ( .A1(n5319), .A2(SI_8_), .ZN(n5347) );
  BUF_X4 U5100 ( .A(n5251), .Z(n4408) );
  XNOR2_X1 U5101 ( .A(n5076), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8608) );
  AND2_X1 U5102 ( .A1(n6244), .A2(n6239), .ZN(n6241) );
  NAND2_X1 U5103 ( .A1(n5868), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5869) );
  OAI21_X1 U5104 ( .B1(n5263), .B2(n5317), .A(n4805), .ZN(n5319) );
  MUX2_X1 U5105 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5866), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5867) );
  XNOR2_X1 U5106 ( .A(n5487), .B(SI_14_), .ZN(n5486) );
  INV_X1 U5107 ( .A(n5331), .ZN(n5330) );
  NAND2_X1 U5108 ( .A1(n5178), .A2(SI_3_), .ZN(n5238) );
  NAND2_X1 U5109 ( .A1(n5302), .A2(n5301), .ZN(n5331) );
  NAND2_X1 U5110 ( .A1(n4522), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6295) );
  AND2_X1 U5111 ( .A1(n4997), .A2(n5864), .ZN(n4786) );
  INV_X1 U5112 ( .A(n5300), .ZN(n5302) );
  NOR3_X1 U5113 ( .A1(n4999), .A2(P1_IR_REG_24__SCAN_IN), .A3(
        P1_IR_REG_28__SCAN_IN), .ZN(n4997) );
  INV_X1 U5114 ( .A(n5229), .ZN(n5228) );
  NAND4_X1 U5115 ( .A1(n5854), .A2(n5948), .A3(n5853), .A4(n10426), .ZN(n5987)
         );
  INV_X1 U5116 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5159) );
  NOR2_X1 U5117 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6072) );
  AND2_X1 U5118 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_7__SCAN_IN), 
        .ZN(n5301) );
  INV_X1 U5119 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5853) );
  NOR2_X1 U5120 ( .A1(P2_IR_REG_13__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5465) );
  INV_X1 U5121 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9478) );
  INV_X1 U5122 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6289) );
  INV_X1 U5123 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n5948) );
  NOR2_X1 U5124 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5852) );
  NOR2_X1 U5125 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n5850) );
  NOR2_X1 U5126 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5084) );
  NOR2_X1 U5127 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), .ZN(
        n5085) );
  INV_X1 U5128 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5272) );
  NOR2_X1 U5129 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n5086) );
  INV_X1 U5130 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4573) );
  INV_X4 U5131 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U5132 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n10423) );
  NAND2_X1 U5133 ( .A1(n8413), .A2(n9917), .ZN(n6271) );
  AOI21_X4 U5134 ( .B1(n9072), .B2(n8422), .A(n8421), .ZN(n9058) );
  AOI21_X2 U5135 ( .B1(n9246), .B2(n9162), .A(n9161), .ZN(n9163) );
  BUF_X1 U5136 ( .A(n9195), .Z(n4409) );
  NAND2_X1 U5137 ( .A1(n5946), .A2(n6998), .ZN(n5935) );
  NAND2_X4 U5138 ( .A1(n6267), .A2(n6616), .ZN(n5946) );
  OR2_X2 U5139 ( .A1(n5472), .A2(n5471), .ZN(n5521) );
  NAND2_X1 U5140 ( .A1(n4856), .A2(n4854), .ZN(n8947) );
  BUF_X4 U5141 ( .A(n6743), .Z(n4410) );
  AND2_X2 U5142 ( .A1(n7616), .A2(n6719), .ZN(n6743) );
  INV_X4 U5143 ( .A(n6012), .ZN(n6353) );
  NAND2_X2 U5144 ( .A1(n6264), .A2(n6279), .ZN(n7616) );
  AND2_X2 U5145 ( .A1(n6645), .A2(n6344), .ZN(n5251) );
  XNOR2_X1 U5146 ( .A(n4614), .B(n5878), .ZN(n6267) );
  NAND2_X2 U5147 ( .A1(n6245), .A2(n9568), .ZN(n6712) );
  BUF_X1 U5148 ( .A(n4411), .Z(n4414) );
  XNOR2_X1 U5149 ( .A(n6747), .B(n6745), .ZN(n9359) );
  INV_X1 U5150 ( .A(n5516), .ZN(n4809) );
  NAND2_X1 U5151 ( .A1(n5493), .A2(n5492), .ZN(n5496) );
  NOR2_X1 U5152 ( .A1(n5489), .A2(n4814), .ZN(n4813) );
  INV_X1 U5153 ( .A(n5464), .ZN(n4814) );
  NAND2_X1 U5154 ( .A1(n4438), .A2(n4535), .ZN(n4534) );
  NAND2_X1 U5155 ( .A1(n4643), .A2(n4644), .ZN(n8559) );
  AOI21_X1 U5156 ( .B1(n4648), .B2(n8739), .A(n4645), .ZN(n4644) );
  INV_X1 U5157 ( .A(n8945), .ZN(n4648) );
  OR2_X1 U5158 ( .A1(n9520), .A2(n9515), .ZN(n6488) );
  NAND3_X1 U5159 ( .A1(n4632), .A2(n5542), .A3(n4630), .ZN(n5561) );
  NAND2_X1 U5160 ( .A1(n4631), .A2(n5056), .ZN(n4630) );
  NAND2_X1 U5161 ( .A1(n5119), .A2(n5118), .ZN(n6645) );
  NAND2_X1 U5162 ( .A1(n8418), .A2(n4913), .ZN(n4909) );
  NOR2_X1 U5163 ( .A1(n8419), .A2(n4914), .ZN(n4913) );
  INV_X1 U5164 ( .A(n8416), .ZN(n4914) );
  INV_X1 U5165 ( .A(n5250), .ZN(n5294) );
  NAND2_X1 U5166 ( .A1(n9396), .A2(n4629), .ZN(n4627) );
  OR2_X1 U5167 ( .A1(n9394), .A2(n9393), .ZN(n4629) );
  OR2_X1 U5168 ( .A1(n6227), .A2(n6226), .ZN(n6268) );
  INV_X1 U5169 ( .A(n6205), .ZN(n6217) );
  AOI21_X1 U5170 ( .B1(n8713), .B2(n8701), .A(n8711), .ZN(n8703) );
  OR4_X1 U5171 ( .A1(n6359), .A2(n6477), .A3(n6358), .A4(n9776), .ZN(n6361) );
  NOR2_X1 U5172 ( .A1(n4436), .A2(n4966), .ZN(n4965) );
  INV_X1 U5173 ( .A(n9380), .ZN(n4966) );
  NAND2_X1 U5174 ( .A1(n5498), .A2(n5497), .ZN(n5542) );
  NAND2_X1 U5175 ( .A1(n5426), .A2(n5425), .ZN(n5429) );
  INV_X1 U5176 ( .A(SI_12_), .ZN(n5425) );
  NAND2_X1 U5177 ( .A1(n5344), .A2(SI_7_), .ZN(n4802) );
  NAND2_X1 U5178 ( .A1(n5264), .A2(SI_6_), .ZN(n5340) );
  NAND2_X1 U5179 ( .A1(n4662), .A2(n8596), .ZN(n4661) );
  AND2_X1 U5180 ( .A1(n8595), .A2(n8600), .ZN(n4662) );
  AND2_X1 U5181 ( .A1(n4931), .A2(n4647), .ZN(n4646) );
  INV_X1 U5182 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5077) );
  AND2_X1 U5183 ( .A1(n5070), .A2(n5069), .ZN(n5071) );
  NOR2_X1 U5184 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n5070) );
  NOR2_X1 U5185 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n5069) );
  INV_X1 U5186 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5068) );
  AND2_X1 U5187 ( .A1(n5067), .A2(n5066), .ZN(n4672) );
  NOR2_X1 U5188 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n5066) );
  INV_X1 U5189 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4699) );
  NAND2_X1 U5190 ( .A1(n7798), .A2(n7797), .ZN(n6775) );
  INV_X1 U5191 ( .A(n4965), .ZN(n4959) );
  NAND2_X1 U5192 ( .A1(n4431), .A2(n4958), .ZN(n4957) );
  NOR2_X1 U5193 ( .A1(n8386), .A2(n4960), .ZN(n4958) );
  INV_X1 U5194 ( .A(n4961), .ZN(n4960) );
  NAND2_X1 U5195 ( .A1(n4431), .A2(n4964), .ZN(n4963) );
  NAND2_X1 U5196 ( .A1(n4567), .A2(n7698), .ZN(n6607) );
  AND2_X1 U5197 ( .A1(n6569), .A2(n6234), .ZN(n6235) );
  NAND2_X1 U5198 ( .A1(n6262), .A2(n6596), .ZN(n5026) );
  NAND2_X1 U5199 ( .A1(n6161), .A2(n4658), .ZN(n6215) );
  AND2_X1 U5200 ( .A1(n4659), .A2(n4508), .ZN(n4658) );
  OR2_X1 U5201 ( .A1(n9545), .A2(n9792), .ZN(n6542) );
  INV_X1 U5202 ( .A(n6515), .ZN(n4580) );
  NAND2_X1 U5203 ( .A1(n10042), .A2(n7724), .ZN(n6577) );
  NOR2_X1 U5204 ( .A1(n4791), .A2(n4796), .ZN(n4789) );
  INV_X1 U5205 ( .A(n4792), .ZN(n4791) );
  NOR2_X1 U5206 ( .A1(n9734), .A2(n4528), .ZN(n4527) );
  INV_X1 U5207 ( .A(n5994), .ZN(n4528) );
  AND2_X1 U5208 ( .A1(n6279), .A2(n9568), .ZN(n6925) );
  NAND2_X1 U5209 ( .A1(n6306), .A2(n6300), .ZN(n6719) );
  NAND2_X1 U5210 ( .A1(n6341), .A2(n6340), .ZN(n6456) );
  NAND2_X1 U5211 ( .A1(n4822), .A2(n4827), .ZN(n6332) );
  AND2_X1 U5212 ( .A1(n5760), .A2(n5727), .ZN(n5758) );
  INV_X1 U5213 ( .A(n5599), .ZN(n4640) );
  AND2_X1 U5214 ( .A1(n5620), .A2(n5605), .ZN(n5618) );
  INV_X1 U5215 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n6044) );
  INV_X1 U5216 ( .A(n5577), .ZN(n5578) );
  NAND2_X1 U5217 ( .A1(n6072), .A2(n10487), .ZN(n4990) );
  AOI21_X1 U5218 ( .B1(n4810), .B2(n4448), .A(n4807), .ZN(n4806) );
  INV_X1 U5219 ( .A(n5496), .ZN(n4807) );
  AND2_X1 U5220 ( .A1(n4810), .A2(n4809), .ZN(n4808) );
  NOR2_X2 U5221 ( .A1(n5855), .A2(n5987), .ZN(n6045) );
  NAND2_X1 U5222 ( .A1(n5290), .A2(n5340), .ZN(n5314) );
  INV_X1 U5223 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4571) );
  NOR2_X1 U5224 ( .A1(n5617), .A2(n5616), .ZN(n4535) );
  AND2_X1 U5225 ( .A1(n7550), .A2(n5122), .ZN(n8761) );
  INV_X1 U5226 ( .A(n7049), .ZN(n7019) );
  INV_X1 U5227 ( .A(n5733), .ZN(n5834) );
  INV_X1 U5228 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4707) );
  NOR2_X2 U5229 ( .A1(n8947), .A2(n9162), .ZN(n8935) );
  NOR2_X1 U5230 ( .A1(n8445), .A2(n8444), .ZN(n4928) );
  AND2_X1 U5231 ( .A1(n4646), .A2(n4929), .ZN(n8961) );
  NOR2_X1 U5232 ( .A1(n9078), .A2(n4911), .ZN(n4908) );
  OR2_X1 U5233 ( .A1(n7269), .A2(n6704), .ZN(n9100) );
  NAND2_X1 U5234 ( .A1(n5565), .A2(n5564), .ZN(n9218) );
  NOR2_X1 U5235 ( .A1(n9312), .A2(n4626), .ZN(n4625) );
  INV_X1 U5236 ( .A(n4628), .ZN(n4626) );
  NAND2_X1 U5237 ( .A1(n9464), .A2(n9465), .ZN(n9463) );
  XNOR2_X1 U5238 ( .A(n4755), .B(n10293), .ZN(n9499) );
  NOR2_X1 U5239 ( .A1(n10009), .A2(n4756), .ZN(n4755) );
  AND2_X1 U5240 ( .A1(n9495), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4756) );
  OR2_X1 U5241 ( .A1(n9520), .A2(n10138), .ZN(n9523) );
  AND2_X1 U5242 ( .A1(n6274), .A2(n6273), .ZN(n9758) );
  NAND2_X1 U5243 ( .A1(n9591), .A2(n6157), .ZN(n9536) );
  AND2_X1 U5244 ( .A1(n9807), .A2(n9581), .ZN(n6593) );
  AOI21_X1 U5245 ( .B1(n4774), .B2(n4773), .A(n4464), .ZN(n4772) );
  INV_X1 U5246 ( .A(n6042), .ZN(n4773) );
  OAI211_X1 U5247 ( .C1(n5006), .C2(n5003), .A(n5001), .B(n6507), .ZN(n9702)
         );
  NAND2_X1 U5248 ( .A1(n5002), .A2(n5004), .ZN(n5001) );
  NOR2_X1 U5249 ( .A1(n8192), .A2(n6496), .ZN(n5004) );
  OR2_X1 U5250 ( .A1(n7628), .A2(n6925), .ZN(n10130) );
  AND2_X1 U5251 ( .A1(n5813), .A2(n9124), .ZN(n8558) );
  AND2_X1 U5252 ( .A1(n6923), .A2(n9408), .ZN(n4985) );
  NAND2_X1 U5253 ( .A1(n6225), .A2(n6224), .ZN(n9515) );
  NAND2_X1 U5254 ( .A1(n6223), .A2(n6469), .ZN(n6225) );
  AND2_X1 U5255 ( .A1(n6222), .A2(n6221), .ZN(n9413) );
  OR2_X1 U5256 ( .A1(n8348), .A2(n6217), .ZN(n6222) );
  OAI21_X1 U5257 ( .B1(n4713), .B2(n4714), .A(n8755), .ZN(n4711) );
  NAND2_X1 U5258 ( .A1(n8624), .A2(n4907), .ZN(n4714) );
  OAI21_X1 U5259 ( .B1(n8612), .B2(n8611), .A(n8622), .ZN(n8613) );
  NAND2_X1 U5260 ( .A1(n8626), .A2(n8638), .ZN(n4713) );
  INV_X1 U5261 ( .A(n8633), .ZN(n4709) );
  NAND2_X1 U5262 ( .A1(n4716), .A2(n4715), .ZN(n8632) );
  AOI21_X1 U5263 ( .B1(n8645), .B2(n8755), .A(n8652), .ZN(n4730) );
  NAND2_X1 U5264 ( .A1(n8281), .A2(n4736), .ZN(n4735) );
  INV_X1 U5265 ( .A(n8686), .ZN(n4736) );
  OAI21_X1 U5266 ( .B1(n4690), .B2(n4689), .A(n4686), .ZN(n6418) );
  NAND2_X1 U5267 ( .A1(n9671), .A2(n6406), .ZN(n4689) );
  NOR2_X1 U5268 ( .A1(n4688), .A2(n4687), .ZN(n4686) );
  AND2_X1 U5269 ( .A1(n9734), .A2(n6563), .ZN(n4563) );
  AND2_X1 U5270 ( .A1(n6247), .A2(n7924), .ZN(n4560) );
  AND2_X1 U5271 ( .A1(n4562), .A2(n10035), .ZN(n4561) );
  OR2_X1 U5272 ( .A1(n8709), .A2(n8755), .ZN(n4721) );
  OR3_X1 U5273 ( .A1(n8720), .A2(n8746), .A3(n8719), .ZN(n8721) );
  NOR2_X1 U5274 ( .A1(n9038), .A2(n4720), .ZN(n4719) );
  NOR2_X1 U5275 ( .A1(n8710), .A2(n8746), .ZN(n4720) );
  NOR2_X1 U5276 ( .A1(n4554), .A2(n9605), .ZN(n4553) );
  OR2_X1 U5277 ( .A1(n9578), .A2(n4555), .ZN(n4554) );
  NOR2_X1 U5278 ( .A1(n6566), .A2(n4557), .ZN(n4556) );
  INV_X1 U5279 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5827) );
  AND2_X1 U5280 ( .A1(n9318), .A2(n9379), .ZN(n4961) );
  OR2_X1 U5281 ( .A1(n6329), .A2(n6328), .ZN(n6333) );
  AOI21_X1 U5282 ( .B1(n5703), .B2(n4829), .A(n4828), .ZN(n4827) );
  INV_X1 U5283 ( .A(n5720), .ZN(n4828) );
  AND2_X1 U5284 ( .A1(n4635), .A2(n4478), .ZN(n4634) );
  NAND2_X1 U5285 ( .A1(n4638), .A2(n4640), .ZN(n4635) );
  OR2_X1 U5286 ( .A1(n5680), .A2(n5681), .ZN(n4697) );
  INV_X1 U5287 ( .A(n5680), .ZN(n4865) );
  NAND2_X1 U5288 ( .A1(n4941), .A2(n4940), .ZN(n4939) );
  NOR2_X1 U5289 ( .A1(n8750), .A2(n8560), .ZN(n4940) );
  NAND2_X1 U5290 ( .A1(n4944), .A2(n8748), .ZN(n4943) );
  NAND2_X1 U5291 ( .A1(n8936), .A2(n8560), .ZN(n4944) );
  NAND2_X1 U5292 ( .A1(n5687), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n5712) );
  NAND2_X1 U5293 ( .A1(n8426), .A2(n8427), .ZN(n8726) );
  NAND2_X1 U5294 ( .A1(n4847), .A2(n9071), .ZN(n4846) );
  INV_X1 U5295 ( .A(n4848), .ZN(n4847) );
  OR2_X1 U5296 ( .A1(n9207), .A2(n9103), .ZN(n9005) );
  AND2_X1 U5297 ( .A1(n9005), .A2(n8717), .ZN(n9078) );
  OR2_X1 U5298 ( .A1(n9211), .A2(n8524), .ZN(n8714) );
  NAND2_X1 U5299 ( .A1(n8131), .A2(n4916), .ZN(n4902) );
  OR2_X1 U5300 ( .A1(n8324), .A2(n8283), .ZN(n8693) );
  AOI21_X1 U5301 ( .B1(n4918), .B2(n4921), .A(n4916), .ZN(n4915) );
  OAI21_X1 U5302 ( .B1(n7576), .B2(n8652), .A(n4922), .ZN(n8076) );
  AND2_X1 U5303 ( .A1(n7746), .A2(n4923), .ZN(n4922) );
  NAND2_X1 U5304 ( .A1(n7734), .A2(n8647), .ZN(n4923) );
  INV_X1 U5305 ( .A(n7345), .ZN(n8614) );
  NAND2_X1 U5306 ( .A1(n5795), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5806) );
  OAI21_X1 U5307 ( .B1(n5376), .B2(P2_IR_REG_9__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5398) );
  INV_X1 U5308 ( .A(n8249), .ZN(n6816) );
  NAND2_X1 U5309 ( .A1(n6831), .A2(n6837), .ZN(n4981) );
  OR2_X1 U5310 ( .A1(n9341), .A2(n9340), .ZN(n6842) );
  NOR2_X1 U5311 ( .A1(n6843), .A2(n4983), .ZN(n4982) );
  INV_X1 U5312 ( .A(n6837), .ZN(n4983) );
  NOR2_X1 U5313 ( .A1(n6035), .A2(n7297), .ZN(n4653) );
  NOR2_X1 U5314 ( .A1(n6013), .A2(n10553), .ZN(n6024) );
  OR2_X1 U5315 ( .A1(n7088), .A2(n6925), .ZN(n6930) );
  NOR2_X1 U5316 ( .A1(n9758), .A2(n6477), .ZN(n4694) );
  NOR2_X1 U5317 ( .A1(n4681), .A2(n4458), .ZN(n4680) );
  OR2_X1 U5318 ( .A1(n6182), .A2(n6181), .ZN(n6192) );
  NOR2_X1 U5319 ( .A1(n9823), .A2(n6853), .ZN(n5038) );
  OR2_X1 U5320 ( .A1(n9817), .A2(n9622), .ZN(n6415) );
  OR2_X1 U5321 ( .A1(n6782), .A2(n10140), .ZN(n8040) );
  NAND2_X1 U5322 ( .A1(n10160), .A2(n7632), .ZN(n6364) );
  AND2_X1 U5323 ( .A1(n6235), .A2(n4480), .ZN(n4792) );
  NAND2_X1 U5324 ( .A1(n9593), .A2(n6555), .ZN(n4591) );
  AND2_X1 U5325 ( .A1(n9655), .A2(n9656), .ZN(n9658) );
  NAND2_X1 U5326 ( .A1(n7919), .A2(n5993), .ZN(n4529) );
  AND2_X1 U5327 ( .A1(n5758), .A2(n5759), .ZN(n6330) );
  OR2_X1 U5328 ( .A1(n5761), .A2(n5760), .ZN(n6336) );
  INV_X1 U5329 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6290) );
  INV_X1 U5330 ( .A(n4639), .ZN(n4638) );
  OAI21_X1 U5331 ( .B1(n4641), .B2(n4640), .A(n5618), .ZN(n4639) );
  AND2_X1 U5332 ( .A1(n5580), .A2(n4642), .ZN(n4641) );
  INV_X1 U5333 ( .A(n5600), .ZN(n4642) );
  NAND2_X1 U5334 ( .A1(n5583), .A2(n5582), .ZN(n5599) );
  XNOR2_X1 U5335 ( .A(n5579), .B(SI_18_), .ZN(n5577) );
  OAI21_X1 U5336 ( .B1(n5561), .B2(n5560), .A(n5559), .ZN(n5562) );
  NAND2_X1 U5337 ( .A1(n5496), .A2(n5495), .ZN(n5516) );
  INV_X1 U5338 ( .A(n4813), .ZN(n4812) );
  AOI21_X1 U5339 ( .B1(n4811), .B2(n4813), .A(n4470), .ZN(n4810) );
  INV_X1 U5340 ( .A(n5055), .ZN(n4811) );
  NAND2_X1 U5341 ( .A1(n5430), .A2(n5429), .ZN(n5463) );
  NOR2_X1 U5342 ( .A1(n5446), .A2(n4818), .ZN(n4817) );
  INV_X1 U5343 ( .A(n5422), .ZN(n4818) );
  NAND2_X1 U5344 ( .A1(n5395), .A2(n4820), .ZN(n4819) );
  NOR2_X1 U5345 ( .A1(n5423), .A2(n4821), .ZN(n4820) );
  INV_X1 U5346 ( .A(n5394), .ZN(n4821) );
  NAND2_X1 U5347 ( .A1(n5371), .A2(n5370), .ZN(n5393) );
  NAND2_X1 U5348 ( .A1(n4804), .A2(n4803), .ZN(n5344) );
  NAND2_X1 U5349 ( .A1(n5269), .A2(n5268), .ZN(n5290) );
  AND2_X1 U5350 ( .A1(n5241), .A2(n5242), .ZN(n4679) );
  OR2_X1 U5351 ( .A1(n5155), .A2(n5154), .ZN(n4675) );
  NAND2_X1 U5352 ( .A1(n5291), .A2(n5106), .ZN(n4853) );
  NAND2_X1 U5353 ( .A1(n8458), .A2(n8457), .ZN(n4540) );
  OAI211_X1 U5354 ( .C1(n9133), .C2(n4661), .A(n4660), .B(n4875), .ZN(n5125)
         );
  NAND2_X1 U5355 ( .A1(n10214), .A2(n4876), .ZN(n4875) );
  BUF_X1 U5356 ( .A(n5304), .Z(n5736) );
  NAND2_X1 U5357 ( .A1(n8513), .A2(n8512), .ZN(n4696) );
  NAND2_X1 U5358 ( .A1(n5547), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5567) );
  INV_X1 U5359 ( .A(n5548), .ZN(n5547) );
  AND2_X1 U5360 ( .A1(n4863), .A2(n5540), .ZN(n4862) );
  NAND2_X1 U5361 ( .A1(n5534), .A2(n5483), .ZN(n4863) );
  INV_X1 U5362 ( .A(n5534), .ZN(n4864) );
  INV_X1 U5363 ( .A(n8550), .ZN(n4869) );
  NAND2_X1 U5364 ( .A1(n4871), .A2(n5718), .ZN(n4870) );
  NAND2_X1 U5365 ( .A1(n4874), .A2(n4873), .ZN(n4872) );
  INV_X1 U5366 ( .A(n8503), .ZN(n4873) );
  NAND2_X1 U5367 ( .A1(n5719), .A2(n4670), .ZN(n4874) );
  AND3_X1 U5368 ( .A1(n5514), .A2(n5513), .A3(n5512), .ZN(n8228) );
  CLKBUF_X1 U5369 ( .A(n5193), .Z(n7052) );
  INV_X1 U5370 ( .A(n5194), .ZN(n5304) );
  OR2_X1 U5371 ( .A1(n5193), .A2(n7241), .ZN(n5128) );
  NAND2_X1 U5372 ( .A1(n8792), .A2(n5050), .ZN(n8803) );
  OR2_X1 U5373 ( .A1(n8369), .A2(n6624), .ZN(n5050) );
  NAND2_X1 U5374 ( .A1(n8845), .A2(n4739), .ZN(n8860) );
  NAND2_X1 U5375 ( .A1(n8849), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n4739) );
  NAND2_X1 U5376 ( .A1(n8860), .A2(n8861), .ZN(n8859) );
  AND2_X1 U5377 ( .A1(n4440), .A2(n10488), .ZN(n4698) );
  OR2_X1 U5378 ( .A1(n5326), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5376) );
  AND2_X1 U5379 ( .A1(n4753), .A2(n4751), .ZN(n4750) );
  OR2_X1 U5380 ( .A1(n6629), .A2(n6688), .ZN(n4753) );
  INV_X1 U5381 ( .A(n8893), .ZN(n4751) );
  AOI21_X1 U5382 ( .B1(n7085), .B2(n6628), .A(n7963), .ZN(n6629) );
  NOR2_X1 U5383 ( .A1(n4749), .A2(n4507), .ZN(n4746) );
  OR2_X1 U5384 ( .A1(n6633), .A2(n8920), .ZN(n4743) );
  INV_X1 U5385 ( .A(n7243), .ZN(n6702) );
  NAND2_X1 U5386 ( .A1(n4881), .A2(n4880), .ZN(n8946) );
  AOI21_X1 U5387 ( .B1(n4882), .B2(n4884), .A(n4465), .ZN(n4880) );
  OR2_X1 U5388 ( .A1(n9177), .A2(n8771), .ZN(n8431) );
  AND2_X1 U5389 ( .A1(n8963), .A2(n4883), .ZN(n4882) );
  NAND2_X1 U5390 ( .A1(n8588), .A2(n8431), .ZN(n4883) );
  INV_X1 U5391 ( .A(n8431), .ZN(n4884) );
  OR2_X1 U5392 ( .A1(n8995), .A2(n8444), .ZN(n4932) );
  NAND2_X1 U5393 ( .A1(n8972), .A2(n8982), .ZN(n8971) );
  INV_X1 U5394 ( .A(n4891), .ZN(n4890) );
  OAI22_X1 U5395 ( .A1(n4897), .A2(n4892), .B1(n9028), .B2(n8428), .ZN(n4891)
         );
  NAND2_X1 U5396 ( .A1(n9058), .A2(n9057), .ZN(n4899) );
  NAND2_X1 U5397 ( .A1(n8423), .A2(n8499), .ZN(n4898) );
  INV_X1 U5398 ( .A(n4899), .ZN(n4896) );
  OAI22_X1 U5399 ( .A1(n8419), .A2(n4912), .B1(n8775), .B2(n9211), .ZN(n4911)
         );
  AND2_X1 U5400 ( .A1(n4924), .A2(n4487), .ZN(n9079) );
  AND2_X1 U5401 ( .A1(n8714), .A2(n8700), .ZN(n9096) );
  AND3_X1 U5402 ( .A1(n5571), .A2(n5570), .A3(n5569), .ZN(n9101) );
  NAND2_X1 U5403 ( .A1(n8326), .A2(n8325), .ZN(n8418) );
  AND2_X1 U5404 ( .A1(n8316), .A2(n8693), .ZN(n8317) );
  NAND2_X1 U5405 ( .A1(n5400), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5451) );
  INV_X1 U5406 ( .A(n5401), .ZN(n5400) );
  NAND2_X1 U5407 ( .A1(n7274), .A2(n8614), .ZN(n7353) );
  INV_X1 U5408 ( .A(n9120), .ZN(n9102) );
  INV_X1 U5409 ( .A(n9138), .ZN(n9081) );
  NAND2_X1 U5410 ( .A1(n7594), .A2(n7593), .ZN(n7601) );
  AND2_X1 U5411 ( .A1(n7592), .A2(n7591), .ZN(n7593) );
  NAND2_X1 U5412 ( .A1(n8395), .A2(n8394), .ZN(n9162) );
  AOI21_X1 U5413 ( .B1(n8448), .B2(n9138), .A(n8447), .ZN(n9164) );
  NAND2_X1 U5414 ( .A1(n5449), .A2(n5448), .ZN(n9238) );
  AOI21_X1 U5415 ( .B1(n6682), .B2(n6695), .A(n4702), .ZN(n4701) );
  NAND2_X1 U5416 ( .A1(n7026), .A2(n8398), .ZN(n4700) );
  AND2_X1 U5417 ( .A1(n4408), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n4702) );
  AND2_X1 U5418 ( .A1(n5818), .A2(n10207), .ZN(n9246) );
  INV_X1 U5419 ( .A(n8595), .ZN(n10207) );
  NAND2_X1 U5420 ( .A1(n8331), .A2(n5798), .ZN(n10179) );
  OR2_X1 U5421 ( .A1(n8268), .A2(n5797), .ZN(n5798) );
  NAND2_X1 U5422 ( .A1(n4737), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U5423 ( .A1(n4934), .A2(n4423), .ZN(n4737) );
  NAND2_X1 U5424 ( .A1(n5806), .A2(n5805), .ZN(n5808) );
  INV_X1 U5425 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5081) );
  NAND2_X1 U5426 ( .A1(n4664), .A2(n4663), .ZN(n5082) );
  AOI21_X1 U5427 ( .B1(n4666), .B2(n9271), .A(n9271), .ZN(n4663) );
  INV_X1 U5428 ( .A(n4667), .ZN(n4666) );
  NAND2_X1 U5429 ( .A1(n4665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U5430 ( .A1(n4878), .A2(n5074), .ZN(n4665) );
  AND2_X1 U5431 ( .A1(n5071), .A2(n5073), .ZN(n4671) );
  INV_X1 U5432 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5073) );
  AND2_X1 U5433 ( .A1(n5465), .A2(n10423), .ZN(n5072) );
  NAND2_X1 U5434 ( .A1(n5273), .A2(n4440), .ZN(n5324) );
  NAND2_X1 U5435 ( .A1(n5028), .A2(n5909), .ZN(n6730) );
  OAI21_X1 U5436 ( .B1(n4963), .B2(n4959), .A(n4957), .ZN(n4953) );
  OAI22_X1 U5437 ( .A1(n4957), .A2(n6880), .B1(n4963), .B2(n4956), .ZN(n4955)
         );
  AND2_X1 U5438 ( .A1(n6890), .A2(n4494), .ZN(n4956) );
  NAND2_X1 U5439 ( .A1(n6077), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n6093) );
  INV_X1 U5440 ( .A(n6078), .ZN(n6077) );
  AND2_X1 U5441 ( .A1(n6930), .A2(n7614), .ZN(n7613) );
  AOI21_X1 U5442 ( .B1(n6722), .B2(n7666), .A(n6720), .ZN(n4951) );
  NAND2_X1 U5443 ( .A1(n4949), .A2(n4950), .ZN(n4948) );
  INV_X1 U5444 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U5445 ( .A1(n6024), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U5446 ( .A1(n6024), .A2(n4653), .ZN(n6054) );
  OAI21_X1 U5447 ( .B1(n4970), .B2(n4969), .A(n4466), .ZN(n4968) );
  INV_X1 U5448 ( .A(n7692), .ZN(n4969) );
  INV_X1 U5449 ( .A(n7475), .ZN(n4616) );
  INV_X1 U5450 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n10553) );
  OR2_X1 U5451 ( .A1(n6000), .A2(n5999), .ZN(n6013) );
  NAND2_X1 U5452 ( .A1(n5913), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5901) );
  NOR2_X1 U5453 ( .A1(n9406), .A2(n4987), .ZN(n9403) );
  OR2_X1 U5454 ( .A1(n9404), .A2(n9405), .ZN(n4987) );
  OR2_X1 U5455 ( .A1(n6066), .A2(n6065), .ZN(n6078) );
  OAI21_X1 U5456 ( .B1(n6615), .B2(n6610), .A(n6618), .ZN(n6611) );
  OR3_X1 U5457 ( .A1(n6607), .A2(n6279), .A3(n10052), .ZN(n4566) );
  NAND2_X1 U5458 ( .A1(n6615), .A2(n6925), .ZN(n4565) );
  OR2_X1 U5459 ( .A1(n6606), .A2(n10052), .ZN(n6609) );
  NAND2_X1 U5460 ( .A1(n4433), .A2(n7174), .ZN(n7173) );
  NAND2_X1 U5461 ( .A1(n7206), .A2(n4606), .ZN(n4605) );
  NAND2_X1 U5462 ( .A1(n7068), .A2(n7102), .ZN(n4606) );
  INV_X1 U5463 ( .A(n4763), .ZN(n4762) );
  OAI21_X1 U5464 ( .B1(n4765), .B2(n4764), .A(n7183), .ZN(n4763) );
  INV_X1 U5465 ( .A(n7184), .ZN(n4764) );
  AOI21_X1 U5466 ( .B1(n4758), .B2(n4428), .A(n4503), .ZN(n7301) );
  INV_X1 U5467 ( .A(n7229), .ZN(n4758) );
  NAND2_X1 U5468 ( .A1(n7301), .A2(n7300), .ZN(n7447) );
  NOR2_X1 U5469 ( .A1(n7457), .A2(n7456), .ZN(n7824) );
  AOI21_X1 U5470 ( .B1(n5025), .B2(n6568), .A(n5024), .ZN(n5023) );
  INV_X1 U5471 ( .A(n9517), .ZN(n5024) );
  NAND2_X1 U5472 ( .A1(n6458), .A2(n6457), .ZN(n9757) );
  NAND2_X1 U5473 ( .A1(n9517), .A2(n6488), .ZN(n6569) );
  INV_X1 U5474 ( .A(n6569), .ZN(n6262) );
  NAND2_X1 U5475 ( .A1(n6214), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n6227) );
  INV_X1 U5476 ( .A(n6215), .ZN(n6214) );
  AOI21_X1 U5477 ( .B1(n8405), .B2(n6205), .A(n6233), .ZN(n9520) );
  AND2_X1 U5478 ( .A1(n6204), .A2(n6215), .ZN(n9411) );
  AND2_X1 U5479 ( .A1(n6197), .A2(n6196), .ZN(n6198) );
  OR2_X1 U5480 ( .A1(n9542), .A2(n9538), .ZN(n6197) );
  NAND2_X1 U5481 ( .A1(n6543), .A2(n6548), .ZN(n8360) );
  AND2_X1 U5482 ( .A1(n6168), .A2(n6167), .ZN(n9547) );
  OR2_X1 U5483 ( .A1(n9570), .A2(n6217), .ZN(n6168) );
  NAND2_X1 U5484 ( .A1(n5019), .A2(n5020), .ZN(n5018) );
  NAND2_X1 U5485 ( .A1(n5017), .A2(n5020), .ZN(n5016) );
  NAND2_X1 U5486 ( .A1(n6412), .A2(n6586), .ZN(n5017) );
  AND2_X1 U5487 ( .A1(n9605), .A2(n6137), .ZN(n4543) );
  AND2_X1 U5488 ( .A1(n6129), .A2(n6128), .ZN(n6859) );
  NAND2_X1 U5489 ( .A1(n6103), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U5490 ( .A1(n6103), .A2(n4654), .ZN(n6130) );
  AND2_X1 U5491 ( .A1(n4581), .A2(n4576), .ZN(n4575) );
  NAND2_X1 U5492 ( .A1(n4582), .A2(n6416), .ZN(n4581) );
  NAND2_X1 U5493 ( .A1(n4578), .A2(n4577), .ZN(n4576) );
  AOI21_X1 U5494 ( .B1(n4780), .B2(n6098), .A(n4456), .ZN(n4778) );
  NAND2_X1 U5495 ( .A1(n4784), .A2(n9834), .ZN(n4783) );
  OR2_X1 U5496 ( .A1(n9669), .A2(n6098), .ZN(n4782) );
  NAND2_X1 U5497 ( .A1(n6076), .A2(n6075), .ZN(n9689) );
  INV_X1 U5498 ( .A(n6043), .ZN(n4776) );
  INV_X1 U5499 ( .A(n5002), .ZN(n5005) );
  OAI21_X1 U5500 ( .B1(n7919), .B2(n4526), .A(n4524), .ZN(n8068) );
  INV_X1 U5501 ( .A(n4527), .ZN(n4526) );
  AOI21_X1 U5502 ( .B1(n4527), .B2(n4525), .A(n4457), .ZN(n4524) );
  AND2_X1 U5503 ( .A1(n5044), .A2(n5043), .ZN(n5042) );
  INV_X1 U5504 ( .A(n7632), .ZN(n7625) );
  NAND2_X1 U5505 ( .A1(n7986), .A2(n5029), .ZN(n10030) );
  NOR2_X1 U5506 ( .A1(n5926), .A2(n5030), .ZN(n5029) );
  NAND2_X1 U5507 ( .A1(n4548), .A2(n4547), .ZN(n10027) );
  AOI21_X1 U5508 ( .B1(n7719), .B2(n7714), .A(n5894), .ZN(n4547) );
  INV_X1 U5509 ( .A(n8404), .ZN(n4523) );
  NAND2_X1 U5510 ( .A1(n6201), .A2(n6200), .ZN(n9776) );
  AND4_X1 U5511 ( .A1(n6059), .A2(n6058), .A3(n6057), .A4(n6056), .ZN(n9868)
         );
  AND2_X1 U5512 ( .A1(n6304), .A2(n6306), .ZN(n7037) );
  INV_X1 U5513 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5864) );
  XNOR2_X1 U5514 ( .A(n6466), .B(n6465), .ZN(n9270) );
  OAI21_X1 U5515 ( .B1(n6456), .B2(n4833), .A(n4831), .ZN(n6466) );
  XNOR2_X1 U5516 ( .A(n6461), .B(n6345), .ZN(n9275) );
  NAND2_X1 U5517 ( .A1(n4836), .A2(n4839), .ZN(n6461) );
  INV_X1 U5518 ( .A(n4990), .ZN(n4988) );
  XNOR2_X1 U5519 ( .A(n5463), .B(n5055), .ZN(n7054) );
  OR2_X1 U5520 ( .A1(n5988), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5947) );
  NAND2_X1 U5521 ( .A1(n5905), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U5522 ( .A1(n5919), .A2(n10392), .ZN(n5920) );
  NOR2_X1 U5523 ( .A1(n9938), .A2(n9937), .ZN(n9939) );
  NAND2_X1 U5524 ( .A1(n9942), .A2(n9943), .ZN(n9944) );
  INV_X1 U5525 ( .A(n9036), .ZN(n9192) );
  INV_X1 U5526 ( .A(n4535), .ZN(n4532) );
  AND2_X1 U5527 ( .A1(n5254), .A2(n5253), .ZN(n7412) );
  INV_X1 U5528 ( .A(n8324), .ZN(n8305) );
  NAND2_X1 U5529 ( .A1(n7272), .A2(n10206), .ZN(n9137) );
  NAND2_X1 U5530 ( .A1(n8374), .A2(n9145), .ZN(n8618) );
  NAND2_X1 U5531 ( .A1(n7441), .A2(n5285), .ZN(n7440) );
  INV_X1 U5532 ( .A(n8517), .ZN(n8553) );
  AOI21_X1 U5533 ( .B1(n4706), .B2(n8550), .A(n8549), .ZN(n4705) );
  NAND2_X1 U5534 ( .A1(n4872), .A2(n4870), .ZN(n4706) );
  AND4_X1 U5535 ( .A1(n4941), .A2(n8590), .A3(n8757), .A4(n8750), .ZN(n8592)
         );
  NAND2_X1 U5536 ( .A1(n4726), .A2(n7550), .ZN(n4725) );
  NAND2_X1 U5537 ( .A1(n4727), .A2(n8759), .ZN(n4726) );
  OAI21_X1 U5538 ( .B1(n8768), .B2(n8767), .A(n8766), .ZN(n4723) );
  NAND2_X1 U5539 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n5120) );
  OAI21_X1 U5540 ( .B1(n7889), .B2(n7029), .A(n8873), .ZN(n7398) );
  NAND2_X1 U5541 ( .A1(n7398), .A2(n7399), .ZN(n7397) );
  NAND2_X1 U5542 ( .A1(n7388), .A2(n7389), .ZN(n7387) );
  NOR2_X1 U5543 ( .A1(n7313), .A2(n4738), .ZN(n7420) );
  NOR2_X1 U5544 ( .A1(n6682), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4738) );
  NAND2_X1 U5545 ( .A1(n7420), .A2(n7419), .ZN(n7418) );
  NOR2_X1 U5546 ( .A1(n7504), .A2(n7505), .ZN(n7503) );
  NAND2_X1 U5547 ( .A1(n4753), .A2(n4747), .ZN(n8270) );
  NAND2_X1 U5548 ( .A1(n6629), .A2(n6688), .ZN(n4747) );
  NOR2_X1 U5549 ( .A1(n4743), .A2(n6634), .ZN(n8918) );
  INV_X1 U5550 ( .A(n9177), .ZN(n8981) );
  NAND2_X1 U5551 ( .A1(n10178), .A2(n5812), .ZN(n9124) );
  NOR2_X1 U5552 ( .A1(n6463), .A2(n5135), .ZN(n5136) );
  INV_X1 U5553 ( .A(n9444), .ZN(n10042) );
  NOR2_X1 U5554 ( .A1(n9403), .A2(n4986), .ZN(n6946) );
  OR2_X1 U5555 ( .A1(n6942), .A2(n6943), .ZN(n4986) );
  NOR2_X1 U5556 ( .A1(n9370), .A2(n4975), .ZN(n4974) );
  INV_X1 U5557 ( .A(n6857), .ZN(n4975) );
  AND2_X1 U5558 ( .A1(n6149), .A2(n6148), .ZN(n9807) );
  OR2_X1 U5559 ( .A1(n7543), .A2(n4412), .ZN(n9384) );
  AND3_X1 U5560 ( .A1(n6921), .A2(n10130), .A3(n6927), .ZN(n9408) );
  INV_X1 U5561 ( .A(n9408), .ZN(n9432) );
  INV_X1 U5562 ( .A(n9547), .ZN(n9782) );
  INV_X1 U5563 ( .A(n9791), .ZN(n9804) );
  OAI21_X1 U5564 ( .B1(n9387), .B2(n6217), .A(n6156), .ZN(n9581) );
  INV_X1 U5565 ( .A(n9877), .ZN(n9439) );
  NAND2_X1 U5566 ( .A1(n4608), .A2(n4607), .ZN(n7103) );
  INV_X1 U5567 ( .A(n7068), .ZN(n4607) );
  INV_X1 U5568 ( .A(n7067), .ZN(n4608) );
  NAND2_X1 U5569 ( .A1(n7111), .A2(n7110), .ZN(n7210) );
  NAND2_X1 U5570 ( .A1(n9463), .A2(n4498), .ZN(n7296) );
  OAI22_X1 U5571 ( .A1(n9498), .A2(n10023), .B1(n9994), .B2(n9499), .ZN(n4754)
         );
  NOR2_X1 U5572 ( .A1(n10026), .A2(n9478), .ZN(n4612) );
  XNOR2_X1 U5573 ( .A(n9757), .B(n9758), .ZN(n9754) );
  AOI21_X1 U5574 ( .B1(n10161), .B2(n6276), .A(n6275), .ZN(n6277) );
  NOR2_X1 U5575 ( .A1(n9758), .A2(n10141), .ZN(n6275) );
  OR3_X1 U5576 ( .A1(n9526), .A2(n6282), .A3(n10132), .ZN(n8408) );
  AOI21_X1 U5577 ( .B1(n4588), .B2(n10168), .A(n4585), .ZN(n9779) );
  NAND2_X1 U5578 ( .A1(n4587), .A2(n4586), .ZN(n4585) );
  XNOR2_X1 U5579 ( .A(n8361), .B(n8360), .ZN(n4588) );
  NAND2_X1 U5580 ( .A1(n9435), .A2(n10161), .ZN(n4586) );
  OR2_X1 U5581 ( .A1(n10089), .A2(n7615), .ZN(n9728) );
  NAND2_X1 U5582 ( .A1(n9711), .A2(n10050), .ZN(n9725) );
  AND2_X1 U5583 ( .A1(n9711), .A2(n7629), .ZN(n9718) );
  NOR2_X1 U5584 ( .A1(n10289), .A2(n4510), .ZN(n10288) );
  NOR2_X1 U5585 ( .A1(n10288), .A2(n10287), .ZN(n10286) );
  OAI21_X1 U5586 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10268), .ZN(n10597) );
  AOI21_X1 U5587 ( .B1(n4473), .B2(n8746), .A(n4709), .ZN(n4708) );
  AND2_X1 U5588 ( .A1(n4713), .A2(n8755), .ZN(n4712) );
  NAND2_X1 U5589 ( .A1(n4728), .A2(n4732), .ZN(n8671) );
  AOI21_X1 U5590 ( .B1(n8661), .B2(n8755), .A(n4733), .ZN(n4732) );
  NOR2_X1 U5591 ( .A1(n6362), .A2(n6473), .ZN(n4687) );
  NOR2_X1 U5592 ( .A1(n6531), .A2(n6477), .ZN(n4688) );
  NAND2_X1 U5593 ( .A1(n4734), .A2(n8698), .ZN(n8713) );
  AOI21_X1 U5594 ( .B1(n6418), .B2(n6417), .A(n6534), .ZN(n6419) );
  NOR2_X1 U5595 ( .A1(n9670), .A2(n8192), .ZN(n4558) );
  NOR2_X1 U5596 ( .A1(n6031), .A2(n4559), .ZN(n6565) );
  OAI21_X1 U5597 ( .B1(n5318), .B2(n5262), .A(n5261), .ZN(n5264) );
  NAND2_X1 U5598 ( .A1(n5263), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n5261) );
  INV_X1 U5599 ( .A(n7674), .ZN(n5459) );
  NAND2_X1 U5600 ( .A1(n8729), .A2(n8728), .ZN(n4717) );
  AND2_X1 U5601 ( .A1(n5627), .A2(n5626), .ZN(n5645) );
  OR2_X1 U5602 ( .A1(n8791), .A2(n7263), .ZN(n7347) );
  NAND2_X1 U5603 ( .A1(n9137), .A2(n8619), .ZN(n8611) );
  AND2_X1 U5604 ( .A1(n6436), .A2(n4684), .ZN(n4683) );
  NAND2_X1 U5605 ( .A1(n4685), .A2(n6477), .ZN(n4684) );
  INV_X1 U5606 ( .A(n6542), .ZN(n4685) );
  INV_X1 U5607 ( .A(n6452), .ZN(n4681) );
  NAND2_X1 U5608 ( .A1(n9542), .A2(n4442), .ZN(n6567) );
  INV_X1 U5609 ( .A(n9592), .ZN(n4552) );
  AND2_X1 U5610 ( .A1(n6424), .A2(n9561), .ZN(n6427) );
  INV_X1 U5611 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10506) );
  AND2_X1 U5612 ( .A1(n6331), .A2(n4824), .ZN(n4823) );
  NAND2_X1 U5613 ( .A1(n4827), .A2(n4825), .ZN(n4824) );
  INV_X1 U5614 ( .A(n4829), .ZN(n4825) );
  INV_X1 U5615 ( .A(n4827), .ZN(n4826) );
  NOR2_X1 U5616 ( .A1(n5721), .A2(n4830), .ZN(n4829) );
  INV_X1 U5617 ( .A(n5702), .ZN(n4830) );
  NOR2_X1 U5618 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5849) );
  NOR2_X1 U5619 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5851) );
  NAND2_X1 U5620 ( .A1(n5318), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n4805) );
  OAI21_X1 U5621 ( .B1(n5244), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n5216), .ZN(
        n5218) );
  OAI21_X1 U5622 ( .B1(n5244), .B2(n5177), .A(n5176), .ZN(n5178) );
  NAND2_X1 U5623 ( .A1(n5244), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5176) );
  OR2_X1 U5624 ( .A1(n5733), .A2(n5167), .ZN(n5170) );
  NAND2_X1 U5625 ( .A1(n4406), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5101) );
  OR2_X1 U5626 ( .A1(n5204), .A2(n6651), .ZN(n5100) );
  AND2_X1 U5627 ( .A1(n4858), .A2(n4857), .ZN(n4856) );
  NOR2_X1 U5628 ( .A1(n9177), .A2(n9182), .ZN(n4858) );
  NAND2_X1 U5629 ( .A1(n5062), .A2(n9010), .ZN(n4892) );
  AND2_X1 U5630 ( .A1(n4889), .A2(n9010), .ZN(n4888) );
  NOR2_X1 U5631 ( .A1(n4893), .A2(n4894), .ZN(n4889) );
  NAND2_X1 U5632 ( .A1(n9044), .A2(n9008), .ZN(n8438) );
  NAND2_X1 U5633 ( .A1(n6158), .A2(n8398), .ZN(n8426) );
  OR2_X1 U5634 ( .A1(n5664), .A2(n10329), .ZN(n5689) );
  AND2_X1 U5635 ( .A1(n8423), .A2(n9066), .ZN(n9007) );
  NAND2_X1 U5636 ( .A1(n5645), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5664) );
  INV_X1 U5637 ( .A(n9007), .ZN(n8710) );
  OR2_X1 U5638 ( .A1(n9207), .A2(n9211), .ZN(n4848) );
  NAND2_X1 U5639 ( .A1(n9096), .A2(n4926), .ZN(n4925) );
  INV_X1 U5640 ( .A(n8699), .ZN(n4926) );
  AND2_X1 U5641 ( .A1(n5057), .A2(n9096), .ZN(n4927) );
  AOI21_X1 U5642 ( .B1(n4920), .B2(n8129), .A(n4919), .ZN(n4918) );
  AND2_X1 U5643 ( .A1(n8644), .A2(n8642), .ZN(n8655) );
  NOR2_X1 U5644 ( .A1(n10237), .A2(n7876), .ZN(n4843) );
  AND2_X1 U5645 ( .A1(n8641), .A2(n8653), .ZN(n8639) );
  AND2_X1 U5646 ( .A1(n4907), .A2(n8624), .ZN(n4935) );
  AND2_X1 U5647 ( .A1(n8611), .A2(n8610), .ZN(n9118) );
  OR2_X1 U5648 ( .A1(n10179), .A2(P2_D_REG_1__SCAN_IN), .ZN(n5802) );
  INV_X1 U5649 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5829) );
  NAND2_X1 U5650 ( .A1(n5117), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5828) );
  OAI21_X1 U5651 ( .B1(n5074), .B2(n9271), .A(n5077), .ZN(n4667) );
  INV_X1 U5652 ( .A(n6764), .ZN(n4972) );
  INV_X1 U5653 ( .A(n6741), .ZN(n4947) );
  OR2_X1 U5654 ( .A1(n9321), .A2(n6872), .ZN(n4967) );
  NAND2_X1 U5655 ( .A1(n7475), .A2(n6764), .ZN(n7795) );
  NAND2_X1 U5656 ( .A1(n6714), .A2(n6925), .ZN(n4950) );
  NOR2_X1 U5657 ( .A1(n7211), .A2(n4766), .ZN(n4765) );
  INV_X1 U5658 ( .A(n7110), .ZN(n4766) );
  INV_X1 U5659 ( .A(n6719), .ZN(n6953) );
  INV_X1 U5660 ( .A(n5026), .ZN(n5025) );
  NAND2_X1 U5661 ( .A1(n9770), .A2(n5036), .ZN(n5035) );
  INV_X1 U5662 ( .A(n6280), .ZN(n5036) );
  NOR2_X1 U5663 ( .A1(n6162), .A2(n6171), .ZN(n4659) );
  INV_X1 U5664 ( .A(n6172), .ZN(n6161) );
  AND2_X1 U5665 ( .A1(n6261), .A2(n9782), .ZN(n6541) );
  NAND2_X1 U5666 ( .A1(n6427), .A2(n4593), .ZN(n4592) );
  NAND2_X1 U5667 ( .A1(n4461), .A2(n4594), .ZN(n4593) );
  NOR2_X1 U5668 ( .A1(n6411), .A2(n5008), .ZN(n5007) );
  INV_X1 U5669 ( .A(n5016), .ZN(n5008) );
  NOR2_X1 U5670 ( .A1(n6411), .A2(n5009), .ZN(n5013) );
  INV_X1 U5671 ( .A(n5018), .ZN(n5009) );
  NOR2_X1 U5672 ( .A1(n6117), .A2(n4655), .ZN(n4654) );
  AND2_X1 U5673 ( .A1(n6091), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6103) );
  INV_X1 U5674 ( .A(n6093), .ZN(n6091) );
  INV_X1 U5675 ( .A(n6531), .ZN(n4582) );
  NAND2_X1 U5676 ( .A1(n4419), .A2(n5000), .ZN(n5002) );
  AND2_X1 U5677 ( .A1(n8183), .A2(n8175), .ZN(n5000) );
  NOR2_X1 U5678 ( .A1(n9880), .A2(n9888), .ZN(n5041) );
  INV_X1 U5679 ( .A(n5993), .ZN(n4525) );
  INV_X1 U5680 ( .A(n5956), .ZN(n4657) );
  NOR2_X1 U5681 ( .A1(n5975), .A2(n10162), .ZN(n5044) );
  NAND2_X1 U5682 ( .A1(n6373), .A2(n8018), .ZN(n7920) );
  AOI22_X1 U5683 ( .A1(n4427), .A2(n4841), .B1(n4832), .B2(n6462), .ZN(n4831)
         );
  INV_X1 U5684 ( .A(n4837), .ZN(n4832) );
  AOI21_X1 U5685 ( .B1(n4841), .B2(n4839), .A(SI_30_), .ZN(n4837) );
  NOR2_X1 U5686 ( .A1(n4427), .A2(n4834), .ZN(n4833) );
  NOR2_X1 U5687 ( .A1(n4838), .A2(n4835), .ZN(n4834) );
  INV_X1 U5688 ( .A(n6462), .ZN(n4835) );
  INV_X1 U5689 ( .A(n4839), .ZN(n4838) );
  NAND2_X1 U5690 ( .A1(n6454), .A2(n6343), .ZN(n4839) );
  INV_X1 U5691 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U5692 ( .A1(n4636), .A2(n4634), .ZN(n5639) );
  NAND2_X1 U5693 ( .A1(n5654), .A2(n5644), .ZN(n5655) );
  OAI21_X1 U5694 ( .B1(n5314), .B2(SI_7_), .A(n5344), .ZN(n5316) );
  NAND2_X1 U5695 ( .A1(n4678), .A2(n4677), .ZN(n5343) );
  NAND2_X1 U5696 ( .A1(n8458), .A2(n4868), .ZN(n4867) );
  INV_X1 U5697 ( .A(n5741), .ZN(n4868) );
  NAND2_X1 U5698 ( .A1(n5485), .A2(n5484), .ZN(n8103) );
  NAND2_X1 U5699 ( .A1(n4438), .A2(n4537), .ZN(n4536) );
  AND2_X1 U5700 ( .A1(n4697), .A2(n4534), .ZN(n4533) );
  INV_X1 U5701 ( .A(n8522), .ZN(n4537) );
  NAND2_X1 U5702 ( .A1(n5414), .A2(n4669), .ZN(n7498) );
  INV_X1 U5703 ( .A(n5415), .ZN(n4669) );
  AND3_X1 U5704 ( .A1(n7530), .A2(n5413), .A3(n7498), .ZN(n7522) );
  INV_X1 U5705 ( .A(n7702), .ZN(n4703) );
  NAND2_X1 U5706 ( .A1(n7705), .A2(n4704), .ZN(n5416) );
  INV_X1 U5707 ( .A(n7817), .ZN(n4704) );
  INV_X1 U5708 ( .A(n7705), .ZN(n5419) );
  NAND2_X1 U5709 ( .A1(n4668), .A2(n5410), .ZN(n7704) );
  INV_X1 U5710 ( .A(n7522), .ZN(n4668) );
  NAND2_X1 U5711 ( .A1(n7440), .A2(n5289), .ZN(n4879) );
  NOR2_X1 U5712 ( .A1(n8569), .A2(n4943), .ZN(n4942) );
  NAND2_X1 U5713 ( .A1(n4939), .A2(n8757), .ZN(n4938) );
  NAND2_X1 U5714 ( .A1(n4475), .A2(n4939), .ZN(n4936) );
  AND3_X1 U5715 ( .A1(n5552), .A2(n5551), .A3(n5550), .ZN(n8283) );
  AND2_X1 U5716 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n8793) );
  NAND2_X1 U5717 ( .A1(n8794), .A2(n8793), .ZN(n8792) );
  NAND2_X1 U5718 ( .A1(n5159), .A2(n5134), .ZN(n5210) );
  OAI21_X1 U5719 ( .B1(n6999), .B2(n6625), .A(n8802), .ZN(n8817) );
  NAND2_X1 U5720 ( .A1(n7370), .A2(n4454), .ZN(n8846) );
  NAND2_X1 U5721 ( .A1(n8846), .A2(n8847), .ZN(n8845) );
  NAND2_X1 U5722 ( .A1(n8859), .A2(n4435), .ZN(n8875) );
  NAND2_X1 U5723 ( .A1(n7387), .A2(n4499), .ZN(n7314) );
  OR2_X1 U5724 ( .A1(n5090), .A2(n9271), .ZN(n5467) );
  AND2_X1 U5725 ( .A1(n4743), .A2(n4742), .ZN(n6635) );
  NAND2_X1 U5726 ( .A1(n8397), .A2(n8396), .ZN(n8936) );
  NAND2_X1 U5727 ( .A1(n4856), .A2(n9015), .ZN(n8957) );
  NAND2_X1 U5728 ( .A1(n9015), .A2(n4858), .ZN(n8975) );
  AND2_X1 U5729 ( .A1(n9015), .A2(n8429), .ZN(n8974) );
  INV_X1 U5730 ( .A(n4846), .ZN(n4844) );
  AND2_X1 U5731 ( .A1(n5633), .A2(n5632), .ZN(n9047) );
  NOR2_X1 U5732 ( .A1(n8393), .A2(n4848), .ZN(n9085) );
  NAND2_X1 U5733 ( .A1(n4924), .A2(n4925), .ZN(n9099) );
  NAND2_X1 U5734 ( .A1(n8436), .A2(n8699), .ZN(n9097) );
  NAND2_X1 U5735 ( .A1(n8317), .A2(n5057), .ZN(n8436) );
  NAND2_X1 U5736 ( .A1(n4415), .A2(n8280), .ZN(n4901) );
  NAND2_X1 U5737 ( .A1(n4903), .A2(n8131), .ZN(n8282) );
  NAND2_X1 U5738 ( .A1(n4904), .A2(n4415), .ZN(n4903) );
  NAND2_X1 U5739 ( .A1(n8128), .A2(n8684), .ZN(n8677) );
  OR2_X1 U5740 ( .A1(n9226), .A2(n8112), .ZN(n8679) );
  INV_X1 U5741 ( .A(n8129), .ZN(n8081) );
  AND4_X1 U5742 ( .A1(n5529), .A2(n5528), .A3(n5527), .A4(n5526), .ZN(n8155)
         );
  NAND2_X1 U5743 ( .A1(n8082), .A2(n8081), .ZN(n8133) );
  NAND2_X1 U5744 ( .A1(n8679), .A2(n8678), .ZN(n8129) );
  NAND2_X1 U5745 ( .A1(n5440), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n5472) );
  INV_X1 U5746 ( .A(n5453), .ZN(n5440) );
  AND2_X1 U5747 ( .A1(n7656), .A2(n4425), .ZN(n8142) );
  NOR2_X1 U5748 ( .A1(n7915), .A2(n9245), .ZN(n4851) );
  NAND2_X1 U5749 ( .A1(n7656), .A2(n4416), .ZN(n7784) );
  AND2_X1 U5750 ( .A1(n8672), .A2(n8670), .ZN(n8583) );
  NAND2_X1 U5751 ( .A1(n7656), .A2(n7657), .ZN(n7757) );
  CLKBUF_X1 U5752 ( .A(n7731), .Z(n7944) );
  CLKBUF_X1 U5753 ( .A(n7564), .Z(n7891) );
  NAND2_X1 U5754 ( .A1(n7576), .A2(n8576), .ZN(n7658) );
  AND4_X1 U5755 ( .A1(n5388), .A2(n5387), .A3(n5386), .A4(n5385), .ZN(n7654)
         );
  NAND2_X1 U5756 ( .A1(n7871), .A2(n4843), .ZN(n7890) );
  NAND2_X1 U5757 ( .A1(n7871), .A2(n10232), .ZN(n7873) );
  INV_X1 U5758 ( .A(n8639), .ZN(n7848) );
  NOR2_X1 U5759 ( .A1(n7644), .A2(n4905), .ZN(n7356) );
  AND2_X1 U5760 ( .A1(n6696), .A2(n6704), .ZN(n9120) );
  INV_X1 U5761 ( .A(n9100), .ZN(n9121) );
  NAND2_X1 U5762 ( .A1(n7268), .A2(n7604), .ZN(n7644) );
  NOR2_X1 U5763 ( .A1(n10206), .A2(n9133), .ZN(n9146) );
  CLKBUF_X1 U5764 ( .A(n8570), .Z(n9136) );
  NAND2_X1 U5765 ( .A1(n4801), .A2(n8399), .ZN(n9153) );
  NAND2_X1 U5766 ( .A1(n9270), .A2(n8398), .ZN(n4801) );
  INV_X1 U5767 ( .A(n10246), .ZN(n9239) );
  OR2_X1 U5768 ( .A1(n8595), .A2(n8758), .ZN(n10246) );
  INV_X1 U5769 ( .A(n9246), .ZN(n10245) );
  NAND2_X1 U5770 ( .A1(n10201), .A2(n5801), .ZN(n7592) );
  OR2_X1 U5771 ( .A1(n10179), .A2(P2_D_REG_0__SCAN_IN), .ZN(n5801) );
  OR2_X1 U5772 ( .A1(n7256), .A2(n7255), .ZN(n7589) );
  AND2_X1 U5773 ( .A1(n5049), .A2(n5074), .ZN(n4877) );
  INV_X1 U5774 ( .A(n4695), .ZN(n5399) );
  AOI21_X1 U5775 ( .B1(n5398), .B2(n5397), .A(n9271), .ZN(n4695) );
  OR2_X1 U5776 ( .A1(n6150), .A2(n9383), .ZN(n6172) );
  NAND2_X1 U5777 ( .A1(n7796), .A2(n6774), .ZN(n4622) );
  INV_X1 U5778 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5999) );
  NAND2_X1 U5779 ( .A1(n9394), .A2(n9393), .ZN(n4628) );
  OR2_X1 U5780 ( .A1(n6141), .A2(n9323), .ZN(n6150) );
  INV_X1 U5781 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5980) );
  OR2_X1 U5782 ( .A1(n5981), .A2(n5980), .ZN(n6000) );
  INV_X1 U5783 ( .A(n4980), .ZN(n4979) );
  OAI21_X1 U5784 ( .B1(n6843), .B2(n4981), .A(n6842), .ZN(n4980) );
  NAND2_X1 U5785 ( .A1(n5939), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5956) );
  INV_X1 U5786 ( .A(n5954), .ZN(n5939) );
  AND2_X1 U5787 ( .A1(n4653), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n4652) );
  OAI21_X1 U5788 ( .B1(n6459), .B2(n9757), .A(n4463), .ZN(n4692) );
  AOI21_X1 U5789 ( .B1(n9757), .B2(n6477), .A(n4694), .ZN(n4693) );
  AND4_X1 U5790 ( .A1(n5945), .A2(n5944), .A3(n5943), .A4(n5942), .ZN(n6754)
         );
  INV_X1 U5791 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7161) );
  OR2_X1 U5792 ( .A1(n5961), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n5964) );
  NAND2_X1 U5793 ( .A1(n7111), .A2(n4765), .ZN(n7208) );
  OAI21_X1 U5794 ( .B1(n7218), .B2(n7217), .A(n4598), .ZN(n9464) );
  NAND2_X1 U5795 ( .A1(n4600), .A2(n4599), .ZN(n4598) );
  INV_X1 U5796 ( .A(n7221), .ZN(n4600) );
  NAND2_X1 U5797 ( .A1(n7447), .A2(n7446), .ZN(n9971) );
  NOR2_X1 U5798 ( .A1(n7824), .A2(n4602), .ZN(n9480) );
  AND2_X1 U5799 ( .A1(n7825), .A2(n7826), .ZN(n4602) );
  NOR2_X1 U5800 ( .A1(n9487), .A2(n4761), .ZN(n9984) );
  OR2_X1 U5801 ( .A1(n9984), .A2(n9983), .ZN(n4760) );
  AND2_X1 U5802 ( .A1(n4760), .A2(n4759), .ZN(n9997) );
  NAND2_X1 U5803 ( .A1(n9987), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4759) );
  NOR2_X1 U5804 ( .A1(n9997), .A2(n9996), .ZN(n9995) );
  NAND2_X1 U5805 ( .A1(n4798), .A2(n4794), .ZN(n4793) );
  OR2_X1 U5806 ( .A1(n8341), .A2(n5026), .ZN(n9518) );
  NAND2_X1 U5807 ( .A1(n4439), .A2(n6569), .ZN(n6263) );
  AND2_X1 U5808 ( .A1(n9594), .A2(n5033), .ZN(n9526) );
  NOR2_X1 U5809 ( .A1(n5035), .A2(n5034), .ZN(n5033) );
  OR2_X1 U5810 ( .A1(n9515), .A2(n6260), .ZN(n5034) );
  NOR2_X1 U5811 ( .A1(n8356), .A2(n5035), .ZN(n8345) );
  NAND2_X1 U5812 ( .A1(n6276), .A2(n10159), .ZN(n4587) );
  NOR2_X1 U5813 ( .A1(n8356), .A2(n8357), .ZN(n9544) );
  OAI21_X1 U5814 ( .B1(n9593), .B2(n4590), .A(n4589), .ZN(n9543) );
  NAND2_X1 U5815 ( .A1(n4461), .A2(n4597), .ZN(n4590) );
  NAND2_X1 U5816 ( .A1(n4592), .A2(n4597), .ZN(n4589) );
  INV_X1 U5817 ( .A(n6541), .ZN(n4597) );
  NAND2_X1 U5818 ( .A1(n9543), .A2(n9542), .ZN(n9541) );
  OR2_X1 U5819 ( .A1(n6195), .A2(n6194), .ZN(n9538) );
  OR2_X1 U5820 ( .A1(n6593), .A2(n4594), .ZN(n9592) );
  AOI21_X1 U5821 ( .B1(n4543), .B2(n6138), .A(n4451), .ZN(n4541) );
  NAND2_X1 U5822 ( .A1(n9620), .A2(n4543), .ZN(n4542) );
  INV_X1 U5823 ( .A(n9817), .ZN(n5037) );
  NAND2_X1 U5824 ( .A1(n9658), .A2(n5038), .ZN(n9625) );
  OR2_X1 U5825 ( .A1(n9637), .A2(n9636), .ZN(n5021) );
  NOR2_X1 U5826 ( .A1(n9664), .A2(n4781), .ZN(n4780) );
  INV_X1 U5827 ( .A(n4783), .ZN(n4781) );
  NAND2_X1 U5828 ( .A1(n9694), .A2(n9693), .ZN(n9692) );
  AOI21_X1 U5829 ( .B1(n4418), .B2(n4775), .A(n4769), .ZN(n4768) );
  INV_X1 U5830 ( .A(n6403), .ZN(n4769) );
  NAND2_X1 U5831 ( .A1(n8058), .A2(n8060), .ZN(n8059) );
  NAND2_X1 U5832 ( .A1(n4657), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U5833 ( .A1(n8002), .A2(n5044), .ZN(n8026) );
  NAND2_X1 U5834 ( .A1(n8002), .A2(n8001), .ZN(n8025) );
  INV_X1 U5835 ( .A(n4995), .ZN(n4994) );
  OAI21_X1 U5836 ( .B1(n10035), .B2(n4996), .A(n6364), .ZN(n4995) );
  INV_X1 U5837 ( .A(n6584), .ZN(n4996) );
  NAND3_X1 U5838 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U5839 ( .A1(n7986), .A2(n10096), .ZN(n7988) );
  NAND2_X1 U5840 ( .A1(n5031), .A2(n7986), .ZN(n10028) );
  NOR2_X1 U5841 ( .A1(n5926), .A2(n7724), .ZN(n5031) );
  NOR2_X1 U5842 ( .A1(n4993), .A2(n4992), .ZN(n4991) );
  INV_X1 U5843 ( .A(n6249), .ZN(n4992) );
  NAND2_X1 U5844 ( .A1(n10082), .A2(n10096), .ZN(n7717) );
  NAND2_X1 U5845 ( .A1(n7774), .A2(n6249), .ZN(n6576) );
  NAND2_X1 U5846 ( .A1(n10061), .A2(n10055), .ZN(n7772) );
  NAND2_X1 U5847 ( .A1(n4788), .A2(n4790), .ZN(n9765) );
  AOI21_X1 U5848 ( .B1(n4792), .B2(n4797), .A(n4459), .ZN(n4790) );
  NAND2_X1 U5849 ( .A1(n4591), .A2(n4461), .ZN(n9562) );
  AND2_X1 U5850 ( .A1(n6189), .A2(n6188), .ZN(n9792) );
  AND2_X1 U5851 ( .A1(n6111), .A2(n6110), .ZN(n9844) );
  AND3_X1 U5852 ( .A1(n6082), .A2(n6081), .A3(n6080), .ZN(n9843) );
  AND4_X1 U5853 ( .A1(n6030), .A2(n6029), .A3(n6028), .A4(n6027), .ZN(n9884)
         );
  NAND2_X1 U5854 ( .A1(n4529), .A2(n4527), .ZN(n9737) );
  NAND2_X1 U5855 ( .A1(n4529), .A2(n5994), .ZN(n9735) );
  INV_X1 U5856 ( .A(n10159), .ZN(n10141) );
  AOI21_X1 U5857 ( .B1(n6957), .B2(n7221), .A(n4621), .ZN(n4620) );
  NOR2_X1 U5858 ( .A1(n6467), .A2(n5355), .ZN(n4621) );
  INV_X1 U5859 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5856) );
  INV_X1 U5860 ( .A(n10130), .ZN(n10163) );
  INV_X1 U5861 ( .A(n10117), .ZN(n10132) );
  INV_X1 U5862 ( .A(n4997), .ZN(n4785) );
  XNOR2_X1 U5863 ( .A(n6456), .B(n6455), .ZN(n8412) );
  XNOR2_X1 U5864 ( .A(n5767), .B(n6328), .ZN(n6223) );
  NAND2_X1 U5865 ( .A1(n6295), .A2(n5877), .ZN(n5027) );
  XNOR2_X1 U5866 ( .A(n5744), .B(n5759), .ZN(n8336) );
  NAND2_X1 U5867 ( .A1(n5742), .A2(n5760), .ZN(n5744) );
  XNOR2_X1 U5868 ( .A(n6298), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6306) );
  XNOR2_X1 U5869 ( .A(n5722), .B(n5721), .ZN(n8267) );
  OAI21_X1 U5870 ( .B1(n5704), .B2(n5703), .A(n5702), .ZN(n5722) );
  AND2_X1 U5871 ( .A1(n5684), .A2(n5661), .ZN(n5682) );
  NAND2_X1 U5872 ( .A1(n6242), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6240) );
  XNOR2_X1 U5873 ( .A(n5656), .B(n5655), .ZN(n7940) );
  NAND2_X1 U5874 ( .A1(n4816), .A2(n5620), .ZN(n5634) );
  NAND2_X1 U5875 ( .A1(n4637), .A2(n5599), .ZN(n5619) );
  NOR2_X1 U5876 ( .A1(n4990), .A2(n4469), .ZN(n4989) );
  NAND2_X1 U5877 ( .A1(n4633), .A2(n4806), .ZN(n5541) );
  NAND2_X1 U5878 ( .A1(n4808), .A2(n5463), .ZN(n4633) );
  OAI21_X1 U5879 ( .B1(n5463), .B2(n4812), .A(n4810), .ZN(n5515) );
  XNOR2_X1 U5880 ( .A(n5490), .B(n5486), .ZN(n7083) );
  NAND2_X1 U5881 ( .A1(n4815), .A2(n5464), .ZN(n5490) );
  NAND2_X1 U5882 ( .A1(n5463), .A2(n5055), .ZN(n4815) );
  NAND2_X1 U5883 ( .A1(n4819), .A2(n5422), .ZN(n5447) );
  NAND2_X1 U5884 ( .A1(n5395), .A2(n5394), .ZN(n5424) );
  OR2_X1 U5885 ( .A1(n5995), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n6006) );
  XNOR2_X1 U5886 ( .A(n5314), .B(n5293), .ZN(n7015) );
  AOI21_X1 U5887 ( .B1(n4675), .B2(n5244), .A(n4674), .ZN(n5156) );
  NOR2_X1 U5888 ( .A1(SI_0_), .A2(SI_1_), .ZN(n4674) );
  NAND2_X1 U5889 ( .A1(n5244), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5138) );
  INV_X1 U5890 ( .A(n5108), .ZN(n5107) );
  NAND2_X1 U5891 ( .A1(n7161), .A2(n5879), .ZN(n5905) );
  INV_X1 U5892 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5879) );
  NOR2_X1 U5893 ( .A1(n9940), .A2(n10594), .ZN(n9941) );
  NAND2_X1 U5894 ( .A1(n9945), .A2(n9946), .ZN(n9947) );
  AND4_X1 U5895 ( .A1(n5337), .A2(n5336), .A3(n5335), .A4(n5334), .ZN(n7577)
         );
  AND2_X1 U5896 ( .A1(n4866), .A2(n4867), .ZN(n8461) );
  NAND2_X1 U5897 ( .A1(n4539), .A2(n4452), .ZN(n4538) );
  AND2_X1 U5898 ( .A1(n5695), .A2(n5694), .ZN(n8505) );
  AND2_X1 U5899 ( .A1(n5613), .A2(n5612), .ZN(n9103) );
  AND4_X1 U5900 ( .A1(n5309), .A2(n5308), .A3(n5307), .A4(n5306), .ZN(n7883)
         );
  INV_X1 U5901 ( .A(n5414), .ZN(n7494) );
  INV_X1 U5902 ( .A(n5125), .ZN(n5124) );
  XNOR2_X1 U5903 ( .A(n9245), .B(n5780), .ZN(n7674) );
  AND4_X1 U5904 ( .A1(n5407), .A2(n5406), .A3(n5405), .A4(n5404), .ZN(n7820)
         );
  NAND2_X1 U5905 ( .A1(n4861), .A2(n4859), .ZN(n8210) );
  AOI21_X1 U5906 ( .B1(n4862), .B2(n4864), .A(n4860), .ZN(n4859) );
  INV_X1 U5907 ( .A(n8121), .ZN(n4860) );
  XNOR2_X1 U5908 ( .A(n5412), .B(n5411), .ZN(n7530) );
  AND4_X1 U5909 ( .A1(n5457), .A2(n5456), .A3(n5455), .A4(n5454), .ZN(n8116)
         );
  NAND2_X1 U5910 ( .A1(n8493), .A2(n8494), .ZN(n8532) );
  INV_X1 U5911 ( .A(n8473), .ZN(n8535) );
  OAI21_X1 U5912 ( .B1(n8372), .B2(n8371), .A(n5137), .ZN(n7362) );
  AND2_X1 U5913 ( .A1(n5595), .A2(n5594), .ZN(n8524) );
  OR2_X1 U5914 ( .A1(n7403), .A2(n9102), .ZN(n8498) );
  INV_X1 U5915 ( .A(n7408), .ZN(n4530) );
  INV_X1 U5916 ( .A(n7407), .ZN(n4531) );
  INV_X1 U5917 ( .A(n8498), .ZN(n8541) );
  INV_X1 U5918 ( .A(n8558), .ZN(n8545) );
  INV_X1 U5919 ( .A(n8505), .ZN(n9028) );
  OR2_X1 U5920 ( .A1(n6637), .A2(n10203), .ZN(n8773) );
  NOR2_X1 U5921 ( .A1(n5204), .A2(n7240), .ZN(n5130) );
  AND2_X1 U5922 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(
        n6652) );
  AND2_X1 U5923 ( .A1(n5327), .A2(n5376), .ZN(n8879) );
  NAND2_X1 U5924 ( .A1(n7397), .A2(n4502), .ZN(n7388) );
  NAND2_X1 U5925 ( .A1(n7418), .A2(n4501), .ZN(n7504) );
  AND2_X1 U5926 ( .A1(n6698), .A2(n6697), .ZN(n7967) );
  AOI21_X1 U5927 ( .B1(n7055), .B2(n7759), .A(n7503), .ZN(n7964) );
  NAND2_X1 U5928 ( .A1(n4752), .A2(n4753), .ZN(n8894) );
  OR2_X1 U5929 ( .A1(n6629), .A2(n4746), .ZN(n4745) );
  NAND2_X1 U5930 ( .A1(n6647), .A2(n6646), .ZN(n8928) );
  INV_X1 U5931 ( .A(n9153), .ZN(n8562) );
  XNOR2_X1 U5932 ( .A(n9157), .B(n9153), .ZN(n9155) );
  INV_X1 U5933 ( .A(n8936), .ZN(n9160) );
  NAND2_X1 U5934 ( .A1(n4929), .A2(n4931), .ZN(n8962) );
  OAI21_X1 U5935 ( .B1(n8972), .B2(n4884), .A(n4882), .ZN(n8954) );
  NAND2_X1 U5936 ( .A1(n8971), .A2(n8431), .ZN(n8955) );
  INV_X1 U5937 ( .A(n4932), .ZN(n8983) );
  OAI21_X1 U5938 ( .B1(n4886), .B2(n9058), .A(n4885), .ZN(n9003) );
  INV_X1 U5939 ( .A(n4897), .ZN(n4886) );
  AOI21_X1 U5940 ( .B1(n4897), .B2(n4894), .A(n4893), .ZN(n4885) );
  NAND2_X1 U5941 ( .A1(n4899), .A2(n4897), .ZN(n9037) );
  NOR2_X1 U5942 ( .A1(n4896), .A2(n4895), .ZN(n9039) );
  INV_X1 U5943 ( .A(n4898), .ZN(n4895) );
  INV_X1 U5944 ( .A(n4911), .ZN(n4910) );
  OAI21_X1 U5945 ( .B1(n8418), .B2(n8417), .A(n8416), .ZN(n9094) );
  NAND2_X1 U5946 ( .A1(n5546), .A2(n5545), .ZN(n8324) );
  NAND2_X1 U5947 ( .A1(n7788), .A2(n7742), .ZN(n7745) );
  INV_X1 U5948 ( .A(n9238), .ZN(n7758) );
  NAND2_X1 U5949 ( .A1(n7353), .A2(n8624), .ZN(n7648) );
  NAND2_X1 U5950 ( .A1(n9144), .A2(n7603), .ZN(n9088) );
  AND2_X1 U5951 ( .A1(n7602), .A2(n5122), .ZN(n9148) );
  INV_X1 U5952 ( .A(n9088), .ZN(n9134) );
  INV_X1 U5953 ( .A(n9021), .ZN(n9076) );
  NAND2_X1 U5954 ( .A1(n9166), .A2(n10243), .ZN(n4511) );
  INV_X2 U5955 ( .A(n10253), .ZN(n10254) );
  NAND2_X1 U5956 ( .A1(n4934), .A2(n4933), .ZN(n9272) );
  AND2_X1 U5957 ( .A1(n4423), .A2(n5094), .ZN(n4933) );
  XNOR2_X1 U5958 ( .A(n5796), .B(P2_IR_REG_24__SCAN_IN), .ZN(n8152) );
  INV_X1 U5959 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10434) );
  INV_X1 U5960 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7430) );
  AND2_X1 U5961 ( .A1(n5090), .A2(n5072), .ZN(n5501) );
  INV_X1 U5962 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10567) );
  INV_X1 U5963 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7086) );
  INV_X1 U5964 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10316) );
  INV_X1 U5965 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7045) );
  INV_X1 U5966 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n7025) );
  NAND2_X1 U5967 ( .A1(n5273), .A2(n5272), .ZN(n5275) );
  INV_X1 U5968 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5139) );
  NAND2_X1 U5969 ( .A1(n4627), .A2(n4628), .ZN(n9311) );
  AND2_X1 U5970 ( .A1(n6211), .A2(n6210), .ZN(n9548) );
  INV_X1 U5971 ( .A(n4955), .ZN(n4954) );
  NAND2_X1 U5972 ( .A1(n9321), .A2(n4953), .ZN(n4952) );
  NAND2_X1 U5973 ( .A1(n4978), .A2(n6837), .ZN(n9343) );
  OR2_X1 U5974 ( .A1(n9329), .A2(n6831), .ZN(n4978) );
  AND2_X1 U5975 ( .A1(n6924), .A2(n7613), .ZN(n9365) );
  NAND2_X1 U5976 ( .A1(n9309), .A2(n6857), .ZN(n4976) );
  AND2_X1 U5977 ( .A1(n4962), .A2(n9318), .ZN(n9382) );
  AND4_X1 U5978 ( .A1(n6005), .A2(n6004), .A3(n6003), .A4(n6002), .ZN(n10140)
         );
  INV_X1 U5979 ( .A(n7956), .ZN(n4617) );
  AND2_X1 U5980 ( .A1(n4618), .A2(n4619), .ZN(n7957) );
  INV_X1 U5981 ( .A(n4968), .ZN(n4619) );
  AND4_X2 U5982 ( .A1(n5903), .A2(n5900), .A3(n5901), .A4(n5902), .ZN(n7765)
         );
  INV_X1 U5983 ( .A(n9425), .ZN(n9386) );
  AND2_X1 U5984 ( .A1(n6124), .A2(n6123), .ZN(n9835) );
  INV_X1 U5985 ( .A(n9429), .ZN(n9410) );
  OR2_X1 U5986 ( .A1(n7543), .A2(n7159), .ZN(n9425) );
  AND2_X1 U5987 ( .A1(n6827), .A2(n6826), .ZN(n9422) );
  OR4_X1 U5988 ( .A1(n6603), .A2(n6246), .A3(n6482), .A4(n8015), .ZN(n6483) );
  NOR2_X1 U5989 ( .A1(n6614), .A2(n4564), .ZN(n6620) );
  NAND2_X1 U5990 ( .A1(n4566), .A2(n4565), .ZN(n4564) );
  INV_X1 U5991 ( .A(n9622), .ZN(n9803) );
  INV_X1 U5992 ( .A(n9835), .ZN(n9436) );
  NAND2_X1 U5993 ( .A1(n5913), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5873) );
  AND2_X1 U5994 ( .A1(n7173), .A2(n7063), .ZN(n9457) );
  INV_X1 U5995 ( .A(n4604), .ZN(n4603) );
  OAI21_X1 U5996 ( .B1(n4605), .B2(n7102), .A(n7105), .ZN(n4604) );
  AND2_X1 U5997 ( .A1(n7192), .A2(n7191), .ZN(n7194) );
  AND2_X1 U5998 ( .A1(n7187), .A2(n7115), .ZN(n7117) );
  AND2_X1 U5999 ( .A1(n7225), .A2(n7159), .ZN(n10013) );
  OAI21_X1 U6000 ( .B1(n7296), .B2(n7295), .A(n7294), .ZN(n7453) );
  XNOR2_X1 U6001 ( .A(n9480), .B(n4601), .ZN(n9479) );
  INV_X1 U6002 ( .A(n9488), .ZN(n4601) );
  INV_X1 U6003 ( .A(n10017), .ZN(n10001) );
  INV_X1 U6004 ( .A(n9501), .ZN(n4611) );
  AOI21_X1 U6005 ( .B1(n9270), .B2(n6469), .A(n6468), .ZN(n9508) );
  NAND2_X1 U6006 ( .A1(n6347), .A2(n6346), .ZN(n9750) );
  AND2_X1 U6007 ( .A1(n9523), .A2(n5065), .ZN(n9524) );
  AND2_X1 U6008 ( .A1(n6268), .A2(n6228), .ZN(n8405) );
  AND2_X1 U6009 ( .A1(n6179), .A2(n6178), .ZN(n9791) );
  OR2_X1 U6010 ( .A1(n9583), .A2(n6217), .ZN(n6179) );
  NAND2_X1 U6011 ( .A1(n4595), .A2(n6555), .ZN(n9579) );
  OR2_X1 U6012 ( .A1(n9593), .A2(n6593), .ZN(n4595) );
  INV_X1 U6013 ( .A(n9581), .ZN(n9814) );
  NAND2_X1 U6014 ( .A1(n5010), .A2(n5016), .ZN(n9607) );
  OR2_X1 U6015 ( .A1(n9637), .A2(n5018), .ZN(n5010) );
  NAND2_X1 U6016 ( .A1(n4544), .A2(n4543), .ZN(n9604) );
  OR2_X1 U6017 ( .A1(n9620), .A2(n6138), .ZN(n4544) );
  NAND2_X1 U6018 ( .A1(n6102), .A2(n6101), .ZN(n9662) );
  NAND2_X1 U6019 ( .A1(n4782), .A2(n4783), .ZN(n9665) );
  OR2_X1 U6020 ( .A1(n8182), .A2(n4775), .ZN(n4771) );
  NAND2_X1 U6021 ( .A1(n8182), .A2(n6042), .ZN(n4777) );
  NAND2_X1 U6022 ( .A1(n8173), .A2(n6504), .ZN(n8186) );
  NAND2_X1 U6023 ( .A1(n7054), .A2(n6469), .ZN(n4569) );
  AND4_X1 U6024 ( .A1(n6041), .A2(n6040), .A3(n6039), .A4(n6038), .ZN(n9877)
         );
  INV_X1 U6025 ( .A(n9718), .ZN(n9659) );
  NAND2_X1 U6026 ( .A1(n6114), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n4551) );
  AOI21_X1 U6027 ( .B1(n6469), .B2(n6992), .A(n4443), .ZN(n4550) );
  INV_X1 U6028 ( .A(n6284), .ZN(n6285) );
  NAND2_X1 U6029 ( .A1(n4523), .A2(n10128), .ZN(n5060) );
  AND2_X2 U6030 ( .A1(n6322), .A2(n6321), .ZN(n10588) );
  AND2_X1 U6031 ( .A1(n6932), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7614) );
  INV_X1 U6032 ( .A(n4998), .ZN(n4787) );
  INV_X1 U6033 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5878) );
  OAI21_X1 U6034 ( .B1(n4998), .B2(n4460), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4614) );
  CLKBUF_X1 U6035 ( .A(n6616), .Z(n9504) );
  INV_X1 U6036 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7700) );
  INV_X1 U6037 ( .A(n6264), .ZN(n7698) );
  INV_X1 U6038 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7533) );
  INV_X1 U6039 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7432) );
  AND2_X1 U6040 ( .A1(n6088), .A2(n6099), .ZN(n10000) );
  INV_X1 U6041 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10437) );
  INV_X1 U6042 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10514) );
  INV_X1 U6043 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10446) );
  NAND2_X1 U6044 ( .A1(n4676), .A2(n5248), .ZN(n5260) );
  XNOR2_X1 U6045 ( .A(n4767), .B(n5891), .ZN(n7143) );
  NAND2_X1 U6046 ( .A1(n5920), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4767) );
  NAND2_X1 U6047 ( .A1(n5920), .A2(n4609), .ZN(n7057) );
  OR2_X1 U6048 ( .A1(n5919), .A2(n10392), .ZN(n4609) );
  OAI21_X1 U6049 ( .B1(n10264), .B2(n9932), .A(n10266), .ZN(n10607) );
  AND2_X1 U6050 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9939), .ZN(n10593) );
  XNOR2_X1 U6051 ( .A(n9941), .B(n4521), .ZN(n10592) );
  INV_X1 U6052 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n4521) );
  XNOR2_X1 U6053 ( .A(n9944), .B(n4519), .ZN(n10606) );
  INV_X1 U6054 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n4519) );
  XNOR2_X1 U6055 ( .A(n9947), .B(n4520), .ZN(n10604) );
  NOR2_X1 U6056 ( .A1(n9951), .A2(n10600), .ZN(n10291) );
  NOR2_X1 U6057 ( .A1(n10286), .A2(n4509), .ZN(n10285) );
  NAND2_X1 U6058 ( .A1(n10285), .A2(n10284), .ZN(n10283) );
  OAI21_X1 U6059 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10283), .ZN(n10281) );
  NAND2_X1 U6060 ( .A1(n10281), .A2(n10282), .ZN(n10280) );
  NAND2_X1 U6061 ( .A1(n10280), .A2(n4513), .ZN(n10278) );
  NAND2_X1 U6062 ( .A1(n4515), .A2(n4514), .ZN(n4513) );
  OAI21_X1 U6063 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10277), .ZN(n10275) );
  OAI21_X1 U6064 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n10274), .ZN(n10272) );
  NAND2_X1 U6065 ( .A1(n10272), .A2(n10273), .ZN(n10271) );
  NAND2_X1 U6066 ( .A1(n10271), .A2(n4516), .ZN(n10269) );
  NAND2_X1 U6067 ( .A1(n4518), .A2(n4517), .ZN(n4516) );
  INV_X1 U6068 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n4518) );
  NAND2_X1 U6069 ( .A1(n4472), .A2(n4705), .ZN(n8557) );
  INV_X1 U6070 ( .A(n4723), .ZN(n4722) );
  NAND2_X1 U6071 ( .A1(n4725), .A2(n4441), .ZN(n4724) );
  NAND2_X1 U6072 ( .A1(n4742), .A2(n4744), .ZN(n8919) );
  NAND2_X1 U6073 ( .A1(n4741), .A2(n4740), .ZN(P2_U3358) );
  NAND2_X1 U6074 ( .A1(P2_STATE_REG_SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4740) );
  NAND2_X1 U6075 ( .A1(n9285), .A2(P2_U3152), .ZN(n4741) );
  OAI211_X1 U6076 ( .C1(n6946), .C2(n6922), .A(n4984), .B(n6941), .ZN(P1_U3218) );
  NAND2_X1 U6077 ( .A1(n6946), .A2(n4985), .ZN(n4984) );
  NAND2_X1 U6078 ( .A1(n7103), .A2(n7102), .ZN(n7207) );
  NOR2_X1 U6079 ( .A1(n4612), .A2(n4611), .ZN(n4610) );
  NAND2_X1 U6080 ( .A1(n9500), .A2(n10052), .ZN(n4757) );
  NAND2_X1 U6081 ( .A1(n4754), .A2(n9568), .ZN(n4613) );
  OR2_X1 U6082 ( .A1(n9779), .A2(n5064), .ZN(n4584) );
  AOI21_X1 U6083 ( .B1(n9777), .B2(n9718), .A(n8362), .ZN(n4583) );
  OAI21_X1 U6084 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9955), .A(n10596), .ZN(
        n9957) );
  AOI21_X1 U6085 ( .B1(n7940), .B2(n8398), .A(n5054), .ZN(n8423) );
  INV_X1 U6086 ( .A(n5718), .ZN(n4670) );
  AND2_X1 U6087 ( .A1(n8677), .A2(n8129), .ZN(n4415) );
  AND2_X1 U6088 ( .A1(n4851), .A2(n7758), .ZN(n4416) );
  INV_X1 U6089 ( .A(n9693), .ZN(n4577) );
  OR2_X1 U6090 ( .A1(n9418), .A2(n9548), .ZN(n4417) );
  AND2_X1 U6091 ( .A1(n4772), .A2(n6259), .ZN(n4418) );
  INV_X1 U6092 ( .A(n9636), .ZN(n5019) );
  INV_X1 U6093 ( .A(n8281), .ZN(n4916) );
  INV_X1 U6094 ( .A(n6573), .ZN(n4568) );
  OR2_X1 U6095 ( .A1(n6256), .A2(n8040), .ZN(n4419) );
  AND2_X1 U6096 ( .A1(n6773), .A2(n7692), .ZN(n4420) );
  AND2_X1 U6097 ( .A1(n6401), .A2(n9704), .ZN(n4421) );
  INV_X1 U6098 ( .A(n4797), .ZN(n4794) );
  NAND2_X1 U6099 ( .A1(n6568), .A2(n4417), .ZN(n4797) );
  AND2_X1 U6100 ( .A1(n4474), .A2(n8494), .ZN(n4422) );
  NAND2_X1 U6101 ( .A1(n4696), .A2(n4493), .ZN(n5719) );
  AND2_X1 U6102 ( .A1(n5092), .A2(n4484), .ZN(n4423) );
  INV_X1 U6103 ( .A(n9515), .ZN(n6283) );
  AND2_X1 U6104 ( .A1(n5041), .A2(n5040), .ZN(n4424) );
  AND2_X1 U6105 ( .A1(n4416), .A2(n4850), .ZN(n4425) );
  AND2_X1 U6106 ( .A1(n7743), .A2(n7742), .ZN(n4426) );
  AND2_X1 U6107 ( .A1(n4839), .A2(SI_30_), .ZN(n4427) );
  AND3_X1 U6108 ( .A1(n6097), .A2(n6096), .A3(n6095), .ZN(n9834) );
  NAND2_X1 U6109 ( .A1(n7234), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4428) );
  INV_X1 U6110 ( .A(n4749), .ZN(n4748) );
  NOR2_X1 U6111 ( .A1(n4429), .A2(n4505), .ZN(n4749) );
  AND2_X1 U6112 ( .A1(n4751), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4429) );
  OR2_X1 U6113 ( .A1(n4748), .A2(n4506), .ZN(n4430) );
  AND2_X2 U6114 ( .A1(n7927), .A2(n9728), .ZN(n5064) );
  OR3_X1 U6115 ( .A1(n8383), .A2(n8380), .A3(n8381), .ZN(n4431) );
  INV_X1 U6116 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5039) );
  AND2_X1 U6117 ( .A1(n7130), .A2(n7061), .ZN(n4433) );
  INV_X1 U6118 ( .A(n5912), .ZN(n6012) );
  NAND2_X1 U6119 ( .A1(n7658), .A2(n8647), .ZN(n7747) );
  INV_X2 U6120 ( .A(n5193), .ZN(n5166) );
  OR2_X1 U6121 ( .A1(n8393), .A2(n9211), .ZN(n4434) );
  OR2_X1 U6122 ( .A1(n7016), .A2(n6626), .ZN(n4435) );
  AND3_X1 U6123 ( .A1(n5192), .A2(n5191), .A3(n5190), .ZN(n7604) );
  NAND2_X1 U6124 ( .A1(n5429), .A2(n5428), .ZN(n5446) );
  NOR2_X1 U6125 ( .A1(n9379), .A2(n9318), .ZN(n4436) );
  INV_X1 U6126 ( .A(n6555), .ZN(n4594) );
  INV_X1 U6127 ( .A(n9057), .ZN(n4894) );
  NAND2_X1 U6128 ( .A1(n7535), .A2(n6751), .ZN(n7471) );
  INV_X1 U6129 ( .A(n9133), .ZN(n10214) );
  NOR2_X1 U6130 ( .A1(n9888), .A2(n9960), .ZN(n4437) );
  AND2_X1 U6131 ( .A1(n4865), .A2(n4422), .ZN(n4438) );
  OR2_X1 U6132 ( .A1(n8341), .A2(n6549), .ZN(n4439) );
  XNOR2_X1 U6133 ( .A(n9172), .B(n8735), .ZN(n8963) );
  OAI21_X1 U6134 ( .B1(n8523), .B2(n8522), .A(n4532), .ZN(n8493) );
  INV_X1 U6135 ( .A(n4775), .ZN(n4774) );
  OR2_X1 U6136 ( .A1(n6060), .A2(n4776), .ZN(n4775) );
  AND2_X1 U6137 ( .A1(n5272), .A2(n4699), .ZN(n4440) );
  INV_X1 U6138 ( .A(n4921), .ZN(n4920) );
  NAND2_X1 U6139 ( .A1(n8128), .A2(n8679), .ZN(n4921) );
  NAND2_X1 U6140 ( .A1(n8133), .A2(n8679), .ZN(n8196) );
  NAND2_X1 U6141 ( .A1(n4771), .A2(n4772), .ZN(n9703) );
  NAND2_X1 U6142 ( .A1(n9692), .A2(n6515), .ZN(n9646) );
  AND2_X1 U6143 ( .A1(n8594), .A2(n8597), .ZN(n4441) );
  AND3_X1 U6144 ( .A1(n4553), .A2(n4552), .A3(n9563), .ZN(n4442) );
  AND2_X1 U6145 ( .A1(n6957), .A2(n7109), .ZN(n4443) );
  NAND2_X1 U6146 ( .A1(n6116), .A2(n6115), .ZN(n6853) );
  AND2_X1 U6147 ( .A1(n6045), .A2(n6044), .ZN(n6073) );
  NAND2_X1 U6148 ( .A1(n4787), .A2(n4786), .ZN(n5868) );
  AOI21_X1 U6149 ( .B1(n8993), .B2(n5834), .A(n5717), .ZN(n9012) );
  AND2_X1 U6150 ( .A1(n6542), .A2(n6440), .ZN(n9542) );
  INV_X1 U6151 ( .A(n4930), .ZN(n8995) );
  NAND2_X1 U6152 ( .A1(n8747), .A2(n8748), .ZN(n8742) );
  INV_X1 U6153 ( .A(n8742), .ZN(n4937) );
  AND2_X1 U6154 ( .A1(n5251), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4444) );
  NOR2_X1 U6155 ( .A1(n6814), .A2(n6818), .ZN(n4445) );
  OR2_X1 U6156 ( .A1(n9776), .A2(n9783), .ZN(n4446) );
  NAND2_X1 U6157 ( .A1(n6073), .A2(n6072), .ZN(n6085) );
  AND2_X1 U6158 ( .A1(n9872), .A2(n9877), .ZN(n6496) );
  NOR2_X1 U6159 ( .A1(n8356), .A2(n6280), .ZN(n4447) );
  INV_X1 U6160 ( .A(n6596), .ZN(n6549) );
  OR2_X1 U6161 ( .A1(n8350), .A2(n9413), .ZN(n6596) );
  AND2_X1 U6162 ( .A1(n5278), .A2(n5277), .ZN(n10232) );
  AND2_X1 U6163 ( .A1(n4812), .A2(n4809), .ZN(n4448) );
  AND2_X1 U6164 ( .A1(n4909), .A2(n4910), .ZN(n4449) );
  AND2_X1 U6165 ( .A1(n4544), .A2(n6137), .ZN(n4450) );
  AND2_X1 U6166 ( .A1(n9817), .A2(n9803), .ZN(n4451) );
  AND2_X1 U6167 ( .A1(n4540), .A2(n8460), .ZN(n4452) );
  AND2_X1 U6168 ( .A1(n4932), .A2(n8588), .ZN(n4453) );
  INV_X1 U6169 ( .A(n6558), .ZN(n5020) );
  OR2_X1 U6170 ( .A1(n7381), .A2(n7809), .ZN(n4454) );
  NAND2_X1 U6171 ( .A1(n5711), .A2(n5710), .ZN(n9182) );
  OR2_X1 U6172 ( .A1(n9168), .A2(n8965), .ZN(n8740) );
  INV_X1 U6173 ( .A(n8740), .ZN(n4645) );
  AND2_X1 U6174 ( .A1(n4752), .A2(n4750), .ZN(n4455) );
  INV_X1 U6175 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10487) );
  AND2_X1 U6176 ( .A1(n9817), .A2(n9622), .ZN(n6411) );
  AND2_X1 U6177 ( .A1(n8040), .A2(n6379), .ZN(n9734) );
  AND2_X1 U6178 ( .A1(n9662), .A2(n9437), .ZN(n4456) );
  NOR2_X1 U6179 ( .A1(n6782), .A2(n9441), .ZN(n4457) );
  NAND2_X1 U6180 ( .A1(n4627), .A2(n4625), .ZN(n9309) );
  NAND2_X1 U6181 ( .A1(n6438), .A2(n6437), .ZN(n4458) );
  AND2_X1 U6182 ( .A1(n9763), .A2(n9762), .ZN(n4459) );
  AND2_X1 U6183 ( .A1(n6407), .A2(n6416), .ZN(n9664) );
  OR2_X1 U6184 ( .A1(n4999), .A2(P1_IR_REG_24__SCAN_IN), .ZN(n4460) );
  AND2_X1 U6185 ( .A1(n6556), .A2(n4596), .ZN(n4461) );
  AND3_X1 U6186 ( .A1(n4799), .A2(n5888), .A3(n5889), .ZN(n4462) );
  AND2_X1 U6187 ( .A1(n6605), .A2(n4693), .ZN(n4463) );
  NOR2_X1 U6188 ( .A1(n9864), .A2(n9438), .ZN(n4464) );
  NOR2_X1 U6189 ( .A1(n9172), .A2(n8770), .ZN(n4465) );
  NAND2_X1 U6190 ( .A1(n6785), .A2(n6784), .ZN(n4466) );
  OR2_X1 U6191 ( .A1(n9182), .A2(n9012), .ZN(n8605) );
  NAND2_X1 U6192 ( .A1(n6073), .A2(n4988), .ZN(n4467) );
  NAND2_X1 U6193 ( .A1(n6262), .A2(n6237), .ZN(n4468) );
  NAND2_X1 U6194 ( .A1(n5769), .A2(n5768), .ZN(n9168) );
  INV_X1 U6195 ( .A(n9168), .ZN(n4855) );
  AND2_X1 U6196 ( .A1(n9038), .A2(n4898), .ZN(n4897) );
  AND2_X1 U6197 ( .A1(n8650), .A2(n8647), .ZN(n8576) );
  INV_X1 U6198 ( .A(n4796), .ZN(n4795) );
  NAND2_X1 U6199 ( .A1(n6198), .A2(n4446), .ZN(n4796) );
  OR2_X1 U6200 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4469) );
  NAND2_X1 U6201 ( .A1(n4782), .A2(n4780), .ZN(n9663) );
  INV_X1 U6202 ( .A(n8684), .ZN(n4919) );
  AND2_X1 U6203 ( .A1(n5488), .A2(SI_14_), .ZN(n4470) );
  AND4_X1 U6204 ( .A1(n4563), .A2(n4561), .A3(n6561), .A4(n4560), .ZN(n4471)
         );
  AND2_X1 U6205 ( .A1(n8689), .A2(n8690), .ZN(n8281) );
  INV_X1 U6206 ( .A(n4579), .ZN(n4578) );
  OR2_X1 U6207 ( .A1(n6518), .A2(n4580), .ZN(n4579) );
  NOR2_X1 U6208 ( .A1(n4846), .A2(n8393), .ZN(n9051) );
  NAND3_X1 U6209 ( .A1(n4872), .A2(n4869), .A3(n4870), .ZN(n4472) );
  NAND2_X1 U6210 ( .A1(n8623), .A2(n7273), .ZN(n4473) );
  NAND2_X1 U6211 ( .A1(n5671), .A2(n8537), .ZN(n4474) );
  AND2_X1 U6212 ( .A1(n8757), .A2(n4937), .ZN(n4475) );
  INV_X1 U6213 ( .A(n5062), .ZN(n4893) );
  INV_X1 U6214 ( .A(n6568), .ZN(n6544) );
  NAND2_X1 U6215 ( .A1(n6596), .A2(n6546), .ZN(n6568) );
  NAND2_X1 U6216 ( .A1(n9693), .A2(n6405), .ZN(n4476) );
  INV_X1 U6217 ( .A(n6773), .ZN(n4973) );
  AND2_X1 U6218 ( .A1(n4622), .A2(n6775), .ZN(n6773) );
  OR2_X1 U6219 ( .A1(n5416), .A2(n4703), .ZN(n4477) );
  AND2_X1 U6220 ( .A1(n5635), .A2(n5620), .ZN(n4478) );
  AND2_X1 U6221 ( .A1(n6747), .A2(n6746), .ZN(n4479) );
  AND2_X1 U6222 ( .A1(n9755), .A2(n10128), .ZN(n4480) );
  NAND2_X1 U6223 ( .A1(n9658), .A2(n9643), .ZN(n9624) );
  OR2_X1 U6224 ( .A1(n5937), .A2(n5936), .ZN(n10031) );
  INV_X1 U6225 ( .A(n10031), .ZN(n5032) );
  AND2_X1 U6226 ( .A1(n5021), .A2(n6586), .ZN(n4481) );
  AND2_X1 U6227 ( .A1(n5038), .A2(n5037), .ZN(n4482) );
  AND2_X1 U6228 ( .A1(n8458), .A2(n4869), .ZN(n4483) );
  INV_X1 U6229 ( .A(n7595), .ZN(n4876) );
  NOR2_X1 U6230 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4484) );
  AND2_X1 U6231 ( .A1(n8725), .A2(n8724), .ZN(n4485) );
  AND2_X1 U6232 ( .A1(n6538), .A2(n6415), .ZN(n4486) );
  AND2_X1 U6233 ( .A1(n6512), .A2(n6515), .ZN(n9693) );
  AND2_X1 U6234 ( .A1(n6415), .A2(n5015), .ZN(n9606) );
  AND2_X1 U6235 ( .A1(n4925), .A2(n8700), .ZN(n4487) );
  AND2_X1 U6236 ( .A1(n4584), .A2(n4583), .ZN(n4488) );
  INV_X1 U6237 ( .A(n6260), .ZN(n9585) );
  AND2_X1 U6238 ( .A1(n9755), .A2(n6570), .ZN(n4489) );
  INV_X1 U6239 ( .A(n4907), .ZN(n8625) );
  NAND2_X1 U6240 ( .A1(n4906), .A2(n4905), .ZN(n4907) );
  NAND2_X1 U6241 ( .A1(n8615), .A2(n8614), .ZN(n4490) );
  AND2_X1 U6242 ( .A1(n8692), .A2(n8691), .ZN(n4491) );
  AND2_X1 U6243 ( .A1(n4867), .A2(n5757), .ZN(n4492) );
  NAND2_X1 U6244 ( .A1(n5698), .A2(n5697), .ZN(n4493) );
  INV_X1 U6245 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5094) );
  OR2_X1 U6246 ( .A1(n4959), .A2(n6877), .ZN(n4494) );
  AND2_X1 U6247 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_REG3_REG_8__SCAN_IN), 
        .ZN(n4495) );
  AND2_X1 U6248 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_27__SCAN_IN), .ZN(
        n4496) );
  INV_X1 U6249 ( .A(n4879), .ZN(n7465) );
  NAND2_X1 U6250 ( .A1(n5925), .A2(n5924), .ZN(n7713) );
  NAND2_X1 U6251 ( .A1(n5607), .A2(n5606), .ZN(n9207) );
  INV_X1 U6252 ( .A(n9207), .ZN(n4849) );
  NAND2_X1 U6253 ( .A1(n8039), .A2(n6257), .ZN(n5006) );
  NAND2_X1 U6254 ( .A1(n5746), .A2(n5745), .ZN(n9172) );
  AND2_X1 U6255 ( .A1(n8058), .A2(n5041), .ZN(n4497) );
  INV_X1 U6256 ( .A(n7673), .ZN(n7681) );
  OAI211_X1 U6257 ( .C1(n4879), .C2(n4477), .A(n5420), .B(n5417), .ZN(n7673)
         );
  XNOR2_X1 U6258 ( .A(n9232), .B(n8781), .ZN(n8667) );
  OR2_X1 U6259 ( .A1(n9469), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n4498) );
  NAND2_X1 U6260 ( .A1(n4770), .A2(n4768), .ZN(n9684) );
  OAI21_X1 U6261 ( .B1(n7475), .B2(n4973), .A(n4970), .ZN(n7691) );
  NAND2_X1 U6262 ( .A1(n4777), .A2(n6043), .ZN(n8191) );
  NAND2_X1 U6263 ( .A1(n4569), .A2(n6034), .ZN(n9872) );
  INV_X1 U6264 ( .A(n9872), .ZN(n5040) );
  AND2_X1 U6265 ( .A1(n5006), .A2(n4419), .ZN(n8174) );
  OR2_X1 U6266 ( .A1(n7384), .A2(n7911), .ZN(n4499) );
  NAND2_X1 U6267 ( .A1(n7656), .A2(n4851), .ZN(n4500) );
  OR2_X1 U6268 ( .A1(n7424), .A2(n6627), .ZN(n4501) );
  OR2_X1 U6269 ( .A1(n7395), .A2(n7900), .ZN(n4502) );
  INV_X1 U6270 ( .A(n8350), .ZN(n9770) );
  NOR2_X1 U6271 ( .A1(n8199), .A2(n8127), .ZN(n8143) );
  NOR2_X1 U6272 ( .A1(n7234), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4503) );
  AND2_X1 U6273 ( .A1(n4654), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n4504) );
  INV_X1 U6274 ( .A(n5503), .ZN(n4878) );
  INV_X1 U6275 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n4656) );
  NAND2_X1 U6276 ( .A1(n5439), .A2(n5438), .ZN(n9232) );
  INV_X1 U6277 ( .A(n9232), .ZN(n4850) );
  NAND2_X1 U6278 ( .A1(n5992), .A2(n4620), .ZN(n10144) );
  INV_X1 U6279 ( .A(n10144), .ZN(n5043) );
  AND2_X1 U6280 ( .A1(n7581), .A2(n9237), .ZN(n9250) );
  INV_X1 U6281 ( .A(n10128), .ZN(n10172) );
  AND2_X1 U6282 ( .A1(n6630), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4505) );
  NAND2_X1 U6283 ( .A1(n6714), .A2(n10052), .ZN(n6473) );
  NAND2_X1 U6284 ( .A1(n6090), .A2(n6089), .ZN(n9847) );
  AND2_X1 U6285 ( .A1(n4751), .A2(n6688), .ZN(n4506) );
  NAND2_X1 U6286 ( .A1(n5329), .A2(n5328), .ZN(n10244) );
  INV_X1 U6287 ( .A(n10244), .ZN(n4842) );
  INV_X1 U6288 ( .A(n6721), .ZN(n7034) );
  INV_X1 U6289 ( .A(n8032), .ZN(n4562) );
  NAND2_X1 U6290 ( .A1(n7286), .A2(n6741), .ZN(n9357) );
  INV_X1 U6291 ( .A(n4841), .ZN(n4840) );
  NOR2_X1 U6292 ( .A1(n6454), .A2(n6343), .ZN(n4841) );
  INV_X1 U6293 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n4655) );
  AND3_X1 U6294 ( .A1(n5886), .A2(n5885), .A3(n5884), .ZN(n9364) );
  NOR2_X1 U6295 ( .A1(n4505), .A2(n6688), .ZN(n4507) );
  NAND2_X1 U6296 ( .A1(n7283), .A2(n6740), .ZN(n7286) );
  NAND2_X1 U6297 ( .A1(n7717), .A2(n6578), .ZN(n7985) );
  AND2_X1 U6298 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(P1_REG3_REG_25__SCAN_IN), 
        .ZN(n4508) );
  XNOR2_X1 U6299 ( .A(n6113), .B(n6112), .ZN(n9568) );
  INV_X1 U6300 ( .A(n9568), .ZN(n10052) );
  INV_X1 U6301 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5079) );
  XNOR2_X1 U6302 ( .A(n5080), .B(n5079), .ZN(n7550) );
  INV_X1 U6303 ( .A(n5099), .ZN(n9278) );
  AND2_X1 U6305 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n4509) );
  AND2_X1 U6306 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n4510) );
  INV_X1 U6307 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n4514) );
  INV_X1 U6308 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n4517) );
  INV_X1 U6309 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5177) );
  INV_X1 U6310 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n4520) );
  INV_X1 U6311 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n4515) );
  INV_X1 U6312 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n4549) );
  INV_X1 U6313 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n4800) );
  INV_X1 U6314 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n4599) );
  NAND2_X1 U6315 ( .A1(n8753), .A2(n8754), .ZN(n4727) );
  NAND2_X2 U6316 ( .A1(n5133), .A2(n5132), .ZN(n8374) );
  AOI21_X1 U6317 ( .B1(n4718), .B2(n4485), .A(n4717), .ZN(n8733) );
  OAI21_X1 U6318 ( .B1(n8687), .B2(n4735), .A(n4491), .ZN(n4734) );
  OAI211_X1 U6319 ( .C1(n4725), .C2(n8760), .A(n4724), .B(n4722), .ZN(P2_U3244) );
  NAND2_X1 U6320 ( .A1(n4490), .A2(n4711), .ZN(n4710) );
  OAI211_X1 U6321 ( .C1(n8632), .C2(n4712), .A(n4710), .B(n4708), .ZN(n8637)
         );
  NAND3_X1 U6322 ( .A1(n9170), .A2(n9169), .A3(n4511), .ZN(n9254) );
  NAND2_X1 U6323 ( .A1(n9004), .A2(n8442), .ZN(n4651) );
  INV_X1 U6324 ( .A(n5291), .ZN(n5263) );
  NAND2_X1 U6325 ( .A1(n4649), .A2(n8729), .ZN(n4930) );
  NOR2_X1 U6326 ( .A1(n9009), .A2(n8443), .ZN(n8997) );
  NOR2_X1 U6327 ( .A1(n8961), .A2(n8739), .ZN(n8941) );
  NAND2_X1 U6328 ( .A1(n5342), .A2(n5343), .ZN(n5354) );
  NAND2_X1 U6329 ( .A1(n10053), .A2(n10056), .ZN(n10061) );
  NAND2_X1 U6330 ( .A1(n6372), .A2(n4512), .ZN(n6374) );
  AND2_X1 U6331 ( .A1(n6525), .A2(n8018), .ZN(n4512) );
  NAND2_X1 U6332 ( .A1(n6250), .A2(n6577), .ZN(n10034) );
  OAI21_X1 U6333 ( .B1(n6445), .B2(n9783), .A(n4683), .ZN(n4682) );
  NAND2_X4 U6334 ( .A1(n5946), .A2(n5291), .ZN(n6467) );
  NAND2_X1 U6335 ( .A1(n7774), .A2(n4991), .ZN(n7716) );
  NAND2_X1 U6336 ( .A1(n4692), .A2(n6471), .ZN(n4691) );
  OAI21_X1 U6337 ( .B1(n6410), .B2(n6411), .A(n4486), .ZN(n6421) );
  INV_X2 U6338 ( .A(n6730), .ZN(n10078) );
  NAND2_X1 U6339 ( .A1(n7741), .A2(n7740), .ZN(n7788) );
  NAND2_X1 U6340 ( .A1(n7639), .A2(n7352), .ZN(n7552) );
  NAND2_X1 U6341 ( .A1(n4890), .A2(n4887), .ZN(n8990) );
  NAND2_X1 U6342 ( .A1(n8284), .A2(n8688), .ZN(n8326) );
  NAND2_X2 U6343 ( .A1(n8989), .A2(n8430), .ZN(n8972) );
  NOR2_X1 U6344 ( .A1(n8365), .A2(n5250), .ZN(n4546) );
  OAI21_X1 U6345 ( .B1(n7879), .B2(n8655), .A(n7561), .ZN(n7731) );
  NAND3_X1 U6346 ( .A1(n6045), .A2(n5039), .A3(n5862), .ZN(n4522) );
  NAND2_X1 U6347 ( .A1(n6430), .A2(n6431), .ZN(n6432) );
  NAND2_X1 U6348 ( .A1(n6730), .A2(n7765), .ZN(n10053) );
  MUX2_X2 U6349 ( .A(n6435), .B(n6434), .S(n6477), .Z(n6445) );
  OR3_X1 U6350 ( .A1(n6394), .A2(n6393), .A3(n6392), .ZN(n6402) );
  AOI22_X1 U6351 ( .A1(n6481), .A2(n6480), .B1(n6599), .B2(n4691), .ZN(n6486)
         );
  NAND2_X1 U6352 ( .A1(n8461), .A2(n4538), .ZN(n8465) );
  NAND4_X1 U6353 ( .A1(n4872), .A2(n4870), .A3(n8457), .A4(n4869), .ZN(n4539)
         );
  NAND3_X1 U6354 ( .A1(n4661), .A2(n9133), .A3(n7595), .ZN(n4660) );
  NAND2_X2 U6355 ( .A1(n5121), .A2(n4545), .ZN(n9133) );
  NOR2_X2 U6356 ( .A1(n4444), .A2(n4546), .ZN(n4545) );
  NAND3_X1 U6357 ( .A1(n7713), .A2(n7985), .A3(n7719), .ZN(n4548) );
  NAND2_X1 U6358 ( .A1(n6577), .A2(n6579), .ZN(n7719) );
  INV_X2 U6359 ( .A(n6271), .ZN(n5913) );
  NAND3_X1 U6360 ( .A1(n5091), .A2(n5090), .A3(n4484), .ZN(n5117) );
  AND3_X2 U6361 ( .A1(n4672), .A2(n4673), .A3(n5071), .ZN(n5090) );
  AND4_X2 U6362 ( .A1(n5068), .A2(n5134), .A3(n5159), .A4(n5272), .ZN(n4673)
         );
  NAND3_X1 U6363 ( .A1(n9621), .A2(n5019), .A3(n4556), .ZN(n4555) );
  NAND3_X1 U6364 ( .A1(n9693), .A2(n9664), .A3(n4558), .ZN(n4557) );
  NAND4_X1 U6365 ( .A1(n6562), .A2(n4471), .A3(n7999), .A4(n8067), .ZN(n4559)
         );
  NAND4_X1 U6366 ( .A1(n6571), .A2(n6572), .A3(n4489), .A4(n4568), .ZN(n4567)
         );
  MUX2_X1 U6367 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n5244), .Z(n5245) );
  NAND3_X1 U6368 ( .A1(n4571), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4570) );
  INV_X1 U6369 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4574) );
  NAND2_X1 U6370 ( .A1(n6555), .A2(n6593), .ZN(n4596) );
  NAND2_X1 U6371 ( .A1(n7131), .A2(n7132), .ZN(n7130) );
  OAI21_X1 U6372 ( .B1(n7067), .B2(n4605), .A(n4603), .ZN(n7192) );
  NAND3_X1 U6373 ( .A1(n4613), .A2(n4757), .A3(n4610), .ZN(P1_U3260) );
  NAND2_X1 U6374 ( .A1(n4618), .A2(n4615), .ZN(n7955) );
  INV_X1 U6375 ( .A(n4806), .ZN(n4631) );
  NAND3_X1 U6376 ( .A1(n4808), .A2(n5056), .A3(n5463), .ZN(n4632) );
  OAI21_X1 U6377 ( .B1(n5581), .B2(n4640), .A(n4638), .ZN(n4816) );
  NAND2_X1 U6378 ( .A1(n5581), .A2(n4638), .ZN(n4636) );
  NAND2_X1 U6379 ( .A1(n5581), .A2(n4641), .ZN(n4637) );
  NAND2_X1 U6380 ( .A1(n5581), .A2(n5580), .ZN(n5601) );
  INV_X1 U6381 ( .A(n8963), .ZN(n4647) );
  NAND3_X1 U6382 ( .A1(n4646), .A2(n4648), .A3(n4929), .ZN(n4643) );
  INV_X1 U6383 ( .A(n8997), .ZN(n4649) );
  NOR2_X1 U6384 ( .A1(n8441), .A2(n9010), .ZN(n4650) );
  NAND2_X1 U6385 ( .A1(n6024), .A2(n4652), .ZN(n6066) );
  NAND2_X1 U6386 ( .A1(n6103), .A2(n4504), .ZN(n6141) );
  NAND2_X1 U6387 ( .A1(n4657), .A2(n4495), .ZN(n5981) );
  NAND2_X1 U6388 ( .A1(n6161), .A2(n4659), .ZN(n6203) );
  NAND2_X1 U6389 ( .A1(n6161), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6174) );
  NAND2_X2 U6390 ( .A1(n4661), .A2(n7595), .ZN(n5747) );
  NAND2_X1 U6391 ( .A1(n4878), .A2(n4666), .ZN(n4664) );
  NAND4_X1 U6392 ( .A1(n4671), .A2(n5072), .A3(n4673), .A4(n4672), .ZN(n5503)
         );
  NAND2_X1 U6393 ( .A1(n4679), .A2(n5243), .ZN(n5248) );
  INV_X1 U6394 ( .A(n5247), .ZN(n4676) );
  NAND3_X1 U6395 ( .A1(n4679), .A2(n5259), .A3(n5243), .ZN(n4677) );
  NAND2_X1 U6396 ( .A1(n5247), .A2(n5259), .ZN(n4678) );
  NAND3_X1 U6397 ( .A1(n4682), .A2(n6453), .A3(n4680), .ZN(n6470) );
  NAND2_X1 U6398 ( .A1(n5273), .A2(n4698), .ZN(n5326) );
  NAND3_X1 U6399 ( .A1(n5134), .A2(n5211), .A3(n5159), .ZN(n5213) );
  NAND4_X1 U6400 ( .A1(n5134), .A2(n5211), .A3(n5159), .A4(n4707), .ZN(n5271)
         );
  NAND2_X1 U6401 ( .A1(n8629), .A2(n8755), .ZN(n4715) );
  NAND2_X1 U6402 ( .A1(n8617), .A2(n8746), .ZN(n4716) );
  NAND3_X1 U6403 ( .A1(n4721), .A2(n8721), .A3(n4719), .ZN(n4718) );
  NAND2_X1 U6404 ( .A1(n8671), .A2(n8662), .ZN(n8663) );
  NAND2_X1 U6405 ( .A1(n4729), .A2(n8654), .ZN(n4728) );
  NAND2_X1 U6406 ( .A1(n4731), .A2(n4730), .ZN(n4729) );
  NAND2_X1 U6407 ( .A1(n8646), .A2(n8746), .ZN(n4731) );
  AND2_X1 U6408 ( .A1(n8660), .A2(n8746), .ZN(n4733) );
  AND2_X2 U6409 ( .A1(n5091), .A2(n5090), .ZN(n4934) );
  MUX2_X1 U6410 ( .A(n7244), .B(n7245), .S(n5134), .Z(n7248) );
  INV_X1 U6411 ( .A(n6634), .ZN(n4742) );
  INV_X1 U6412 ( .A(n6633), .ZN(n4744) );
  NAND2_X1 U6413 ( .A1(n4745), .A2(n4430), .ZN(n8904) );
  OR2_X1 U6414 ( .A1(n8270), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n4752) );
  INV_X1 U6415 ( .A(n4760), .ZN(n9982) );
  AND2_X1 U6416 ( .A1(n9489), .A2(n9488), .ZN(n4761) );
  OAI21_X1 U6417 ( .B1(n7111), .B2(n4764), .A(n4762), .ZN(n7187) );
  NAND2_X1 U6418 ( .A1(n8182), .A2(n4418), .ZN(n4770) );
  NAND2_X1 U6419 ( .A1(n9669), .A2(n4780), .ZN(n4779) );
  INV_X1 U6420 ( .A(n9847), .ZN(n4784) );
  NOR2_X1 U6421 ( .A1(n4998), .A2(n4785), .ZN(n5865) );
  NAND2_X1 U6422 ( .A1(n6045), .A2(n5862), .ZN(n4998) );
  NAND2_X1 U6423 ( .A1(n6199), .A2(n4795), .ZN(n4798) );
  NAND2_X1 U6424 ( .A1(n6199), .A2(n4789), .ZN(n4788) );
  NAND2_X1 U6425 ( .A1(n6199), .A2(n6198), .ZN(n8355) );
  NAND2_X1 U6426 ( .A1(n4798), .A2(n4417), .ZN(n8340) );
  NAND2_X2 U6427 ( .A1(n4462), .A2(n5890), .ZN(n10082) );
  OR2_X1 U6428 ( .A1(n6271), .A2(n4800), .ZN(n4799) );
  AND2_X1 U6429 ( .A1(n9768), .A2(n9767), .ZN(n5061) );
  AOI21_X1 U6430 ( .B1(n9766), .B2(n10117), .A(n9765), .ZN(n9767) );
  NAND2_X1 U6431 ( .A1(n6708), .A2(n8591), .ZN(n6709) );
  NOR2_X2 U6432 ( .A1(n8413), .A2(n5872), .ZN(n5912) );
  NAND2_X1 U6433 ( .A1(n5952), .A2(n5951), .ZN(n10162) );
  AND2_X1 U6434 ( .A1(n9153), .A2(n8564), .ZN(n8599) );
  INV_X4 U6435 ( .A(n5291), .ZN(n6998) );
  NAND2_X1 U6436 ( .A1(n5347), .A2(n4802), .ZN(n5351) );
  NAND2_X1 U6437 ( .A1(n5291), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n4803) );
  NAND2_X1 U6438 ( .A1(n5318), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4804) );
  NAND2_X1 U6439 ( .A1(n4819), .A2(n4817), .ZN(n5430) );
  NAND2_X1 U6440 ( .A1(n5704), .A2(n4829), .ZN(n4822) );
  OAI21_X1 U6441 ( .B1(n5704), .B2(n4826), .A(n4823), .ZN(n6341) );
  NAND2_X1 U6442 ( .A1(n6456), .A2(n4840), .ZN(n4836) );
  NAND2_X1 U6443 ( .A1(n5144), .A2(n5114), .ZN(n8365) );
  INV_X1 U6444 ( .A(n8393), .ZN(n4845) );
  NAND3_X1 U6445 ( .A1(n4845), .A2(n4844), .A3(n8423), .ZN(n9030) );
  NAND2_X1 U6446 ( .A1(n4853), .A2(n4852), .ZN(n5108) );
  AOI21_X1 U6447 ( .B1(n5244), .B2(n5105), .A(n5135), .ZN(n4852) );
  INV_X1 U6448 ( .A(n9172), .ZN(n4857) );
  NAND2_X1 U6449 ( .A1(n5485), .A2(n4862), .ZN(n4861) );
  OAI21_X1 U6450 ( .B1(n5485), .B2(n4864), .A(n4862), .ZN(n8120) );
  NAND2_X1 U6451 ( .A1(n8493), .A2(n4422), .ZN(n8470) );
  NAND2_X1 U6452 ( .A1(n4866), .A2(n4492), .ZN(n5823) );
  NAND3_X1 U6453 ( .A1(n4872), .A2(n4870), .A3(n4483), .ZN(n4866) );
  INV_X1 U6454 ( .A(n5719), .ZN(n4871) );
  NAND2_X1 U6455 ( .A1(n4878), .A2(n4877), .ZN(n5075) );
  INV_X1 U6456 ( .A(n4934), .ZN(n5789) );
  NAND2_X1 U6457 ( .A1(n8972), .A2(n4882), .ZN(n4881) );
  NAND2_X1 U6458 ( .A1(n9058), .A2(n4888), .ZN(n4887) );
  INV_X1 U6459 ( .A(n8132), .ZN(n4904) );
  OAI21_X2 U6460 ( .B1(n8132), .B2(n4901), .A(n4900), .ZN(n8284) );
  NAND2_X1 U6461 ( .A1(n4902), .A2(n8280), .ZN(n4900) );
  INV_X2 U6462 ( .A(n10227), .ZN(n4905) );
  NAND2_X1 U6463 ( .A1(n8417), .A2(n8416), .ZN(n4912) );
  NAND2_X1 U6464 ( .A1(n5117), .A2(n4496), .ZN(n6643) );
  NAND2_X1 U6465 ( .A1(n8082), .A2(n4918), .ZN(n4917) );
  NAND2_X1 U6466 ( .A1(n4917), .A2(n4915), .ZN(n8289) );
  OAI21_X1 U6467 ( .B1(n8082), .B2(n4921), .A(n4918), .ZN(n8134) );
  NAND2_X1 U6468 ( .A1(n8076), .A2(n8075), .ZN(n8079) );
  NAND2_X1 U6469 ( .A1(n8730), .A2(n8982), .ZN(n4931) );
  NAND2_X1 U6470 ( .A1(n4930), .A2(n4928), .ZN(n4929) );
  NAND2_X1 U6471 ( .A1(n7353), .A2(n4935), .ZN(n7569) );
  INV_X1 U6472 ( .A(n8569), .ZN(n4941) );
  OAI22_X1 U6473 ( .A1(n8559), .A2(n4936), .B1(n4938), .B2(n4942), .ZN(n8565)
         );
  NAND3_X1 U6474 ( .A1(n7283), .A2(n6740), .A3(n9359), .ZN(n4946) );
  AOI21_X1 U6475 ( .B1(n4947), .B2(n9359), .A(n4479), .ZN(n4945) );
  NAND2_X1 U6476 ( .A1(n9357), .A2(n9359), .ZN(n9358) );
  INV_X1 U6477 ( .A(n8386), .ZN(n4964) );
  NAND2_X1 U6478 ( .A1(n4954), .A2(n4952), .ZN(n6895) );
  NAND2_X1 U6479 ( .A1(n6773), .A2(n4972), .ZN(n4971) );
  AND2_X1 U6480 ( .A1(n6778), .A2(n4971), .ZN(n4970) );
  NAND2_X1 U6481 ( .A1(n9309), .A2(n4974), .ZN(n6866) );
  XNOR2_X1 U6482 ( .A(n4976), .B(n9373), .ZN(n9378) );
  NAND2_X1 U6483 ( .A1(n9329), .A2(n4982), .ZN(n4977) );
  NAND2_X1 U6484 ( .A1(n4977), .A2(n4979), .ZN(n9396) );
  NAND3_X1 U6485 ( .A1(n6045), .A2(n6044), .A3(n4989), .ZN(n6238) );
  INV_X2 U6486 ( .A(n7765), .ZN(n6729) );
  INV_X1 U6487 ( .A(n6578), .ZN(n4993) );
  XNOR2_X1 U6488 ( .A(n6576), .B(n6561), .ZN(n7983) );
  INV_X1 U6489 ( .A(n5863), .ZN(n4999) );
  NAND2_X1 U6490 ( .A1(n5006), .A2(n5005), .ZN(n8173) );
  INV_X1 U6491 ( .A(n5004), .ZN(n5003) );
  INV_X1 U6492 ( .A(n6411), .ZN(n5015) );
  INV_X1 U6493 ( .A(n5021), .ZN(n9635) );
  NAND2_X1 U6494 ( .A1(n5022), .A2(n5023), .ZN(n9519) );
  NAND2_X1 U6495 ( .A1(n8342), .A2(n5025), .ZN(n5022) );
  NOR2_X1 U6496 ( .A1(n8342), .A2(n6568), .ZN(n8341) );
  NAND2_X1 U6497 ( .A1(n10078), .A2(n10049), .ZN(n10048) );
  NAND2_X1 U6498 ( .A1(n9364), .A2(n5032), .ZN(n5030) );
  NAND2_X1 U6499 ( .A1(n8058), .A2(n4424), .ZN(n8188) );
  AOI21_X2 U6500 ( .B1(n9302), .B2(n9300), .A(n9299), .ZN(n9351) );
  NAND2_X1 U6501 ( .A1(n6246), .A2(n6264), .ZN(n7088) );
  NAND2_X1 U6502 ( .A1(n8946), .A2(n8945), .ZN(n8944) );
  NOR2_X1 U6503 ( .A1(n5131), .A2(n5130), .ZN(n5133) );
  OR2_X2 U6504 ( .A1(n8356), .A2(n9795), .ZN(n9566) );
  NAND2_X1 U6505 ( .A1(n5104), .A2(n5103), .ZN(n7261) );
  CLKBUF_X1 U6506 ( .A(n8289), .Z(n8285) );
  INV_X1 U6507 ( .A(n8413), .ZN(n5870) );
  INV_X1 U6508 ( .A(n5098), .ZN(n5097) );
  NAND2_X1 U6509 ( .A1(n5098), .A2(n5099), .ZN(n5193) );
  INV_X1 U6510 ( .A(n9004), .ZN(n9080) );
  NAND2_X1 U6511 ( .A1(n9759), .A2(n9526), .ZN(n9529) );
  INV_X1 U6512 ( .A(n6467), .ZN(n5908) );
  INV_X1 U6513 ( .A(n8042), .ZN(n6031) );
  AND2_X1 U6514 ( .A1(n8095), .A2(n8092), .ZN(n5045) );
  NOR2_X1 U6515 ( .A1(n6251), .A2(n7922), .ZN(n5046) );
  OR2_X1 U6516 ( .A1(n8755), .A2(n8638), .ZN(n5047) );
  NAND2_X1 U6517 ( .A1(n7351), .A2(n7350), .ZN(n7639) );
  AND2_X1 U6518 ( .A1(n6803), .A2(n6802), .ZN(n5048) );
  AND3_X1 U6519 ( .A1(n5079), .A2(n5081), .A3(n5077), .ZN(n5049) );
  AND2_X1 U6520 ( .A1(n8143), .A2(n8145), .ZN(n5051) );
  INV_X1 U6521 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n5317) );
  INV_X1 U6522 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n5292) );
  AND2_X1 U6523 ( .A1(n5394), .A2(n5375), .ZN(n5052) );
  AND2_X1 U6524 ( .A1(n5370), .A2(n5359), .ZN(n5053) );
  INV_X1 U6525 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5262) );
  AND2_X1 U6526 ( .A1(n4408), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n5054) );
  MUX2_X1 U6527 ( .A(n5134), .B(n9283), .S(n6645), .Z(n9145) );
  NOR2_X2 U6528 ( .A1(n5059), .A2(n9847), .ZN(n9655) );
  AND2_X1 U6529 ( .A1(n5464), .A2(n5434), .ZN(n5055) );
  INV_X1 U6530 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5805) );
  AND2_X1 U6531 ( .A1(n5542), .A2(n5500), .ZN(n5056) );
  OR2_X1 U6532 ( .A1(n7088), .A2(n4412), .ZN(n10138) );
  AND2_X1 U6533 ( .A1(n8701), .A2(n8699), .ZN(n5057) );
  NOR2_X1 U6534 ( .A1(n6620), .A2(n6619), .ZN(n5058) );
  NAND2_X1 U6535 ( .A1(n5838), .A2(n5819), .ZN(n8549) );
  INV_X1 U6536 ( .A(n9413), .ZN(n6276) );
  OR2_X1 U6537 ( .A1(n9036), .A2(n9048), .ZN(n5062) );
  INV_X1 U6538 ( .A(n10237), .ZN(n7563) );
  AND2_X1 U6539 ( .A1(n8639), .A2(n5047), .ZN(n5063) );
  NAND2_X1 U6540 ( .A1(n9146), .A2(n10222), .ZN(n9127) );
  OR2_X1 U6541 ( .A1(n9522), .A2(n9521), .ZN(n5065) );
  AND2_X1 U6542 ( .A1(n8629), .A2(n8633), .ZN(n7568) );
  AND2_X1 U6543 ( .A1(n7571), .A2(n8638), .ZN(n7572) );
  INV_X1 U6544 ( .A(n6743), .ZN(n6748) );
  OR2_X1 U6545 ( .A1(n6046), .A2(n6289), .ZN(n6239) );
  AOI21_X1 U6546 ( .B1(n8738), .B2(n8737), .A(n4645), .ZN(n8745) );
  INV_X1 U6547 ( .A(n5689), .ZN(n5687) );
  NAND2_X1 U6548 ( .A1(n5244), .A2(n6990), .ZN(n5216) );
  INV_X1 U6549 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5450) );
  INV_X1 U6550 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n10488) );
  INV_X1 U6551 ( .A(n6611), .ZN(n6612) );
  INV_X1 U6552 ( .A(n6564), .ZN(n6247) );
  OR2_X1 U6553 ( .A1(n6241), .A2(n6290), .ZN(n6243) );
  INV_X1 U6554 ( .A(n5486), .ZN(n5489) );
  INV_X1 U6555 ( .A(n8549), .ZN(n8457) );
  AND2_X1 U6556 ( .A1(n7366), .A2(n9122), .ZN(n5123) );
  AND2_X1 U6557 ( .A1(n6632), .A2(n8931), .ZN(n6633) );
  OR2_X1 U6558 ( .A1(n7000), .A2(n5250), .ZN(n5165) );
  OR2_X1 U6559 ( .A1(n6738), .A2(n6737), .ZN(n6741) );
  AND2_X1 U6560 ( .A1(n6862), .A2(n6863), .ZN(n9370) );
  INV_X1 U6561 ( .A(n9318), .ZN(n6879) );
  INV_X1 U6562 ( .A(n6348), .ZN(n6231) );
  INV_X1 U6563 ( .A(n9807), .ZN(n9600) );
  OR2_X1 U6564 ( .A1(n6339), .A2(n6338), .ZN(n6340) );
  INV_X1 U6565 ( .A(n5699), .ZN(n5703) );
  NAND2_X1 U6566 ( .A1(n5642), .A2(n5641), .ZN(n5654) );
  NAND2_X1 U6567 ( .A1(n5432), .A2(n5431), .ZN(n5464) );
  NAND2_X1 U6568 ( .A1(n5218), .A2(n5217), .ZN(n5239) );
  OR2_X1 U6569 ( .A1(n5174), .A2(n5173), .ZN(n5175) );
  NAND2_X1 U6570 ( .A1(n5843), .A2(n5842), .ZN(n8517) );
  OR2_X1 U6571 ( .A1(n7944), .A2(n8576), .ZN(n7653) );
  NAND2_X1 U6572 ( .A1(n5808), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5796) );
  AND2_X1 U6573 ( .A1(n6905), .A2(n6904), .ZN(n6943) );
  AND2_X1 U6574 ( .A1(n6889), .A2(n6888), .ZN(n8386) );
  AND3_X1 U6575 ( .A1(n6996), .A2(n7611), .A3(n7608), .ZN(n6927) );
  NAND2_X1 U6576 ( .A1(n6348), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5917) );
  AND2_X1 U6577 ( .A1(n7160), .A2(n6973), .ZN(n7225) );
  INV_X1 U6578 ( .A(n9757), .ZN(n9759) );
  INV_X1 U6579 ( .A(n6853), .ZN(n9643) );
  AND2_X1 U6580 ( .A1(n6928), .A2(n4412), .ZN(n10159) );
  AND2_X1 U6581 ( .A1(n6281), .A2(n6279), .ZN(n10117) );
  NAND2_X1 U6582 ( .A1(n6714), .A2(n7698), .ZN(n7628) );
  OR2_X1 U6583 ( .A1(n5865), .A2(n6046), .ZN(n5866) );
  INV_X1 U6584 ( .A(n5248), .ZN(n5246) );
  NOR2_X1 U6585 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10593), .ZN(n9940) );
  OAI21_X1 U6586 ( .B1(n7362), .B2(n7361), .A(n5175), .ZN(n7326) );
  NOR2_X1 U6587 ( .A1(n5841), .A2(n5810), .ZN(n5838) );
  INV_X1 U6588 ( .A(n8543), .ZN(n8495) );
  AND4_X1 U6589 ( .A1(n5477), .A2(n5476), .A3(n5475), .A4(n5474), .ZN(n8112)
         );
  OR2_X1 U6590 ( .A1(n5204), .A2(n6658), .ZN(n5208) );
  NAND2_X1 U6591 ( .A1(n8803), .A2(n8804), .ZN(n8802) );
  OR2_X1 U6592 ( .A1(P2_U3966), .A2(n6641), .ZN(n6705) );
  NAND2_X1 U6593 ( .A1(n8875), .A2(n8876), .ZN(n8873) );
  INV_X1 U6594 ( .A(n8917), .ZN(n8874) );
  INV_X1 U6595 ( .A(n8932), .ZN(n8878) );
  NAND2_X1 U6596 ( .A1(n8566), .A2(n8596), .ZN(n9138) );
  OR2_X1 U6597 ( .A1(n7592), .A2(n7307), .ZN(n7308) );
  AND3_X1 U6598 ( .A1(n7550), .A2(n8591), .A3(n5811), .ZN(n10249) );
  INV_X1 U6599 ( .A(n9250), .ZN(n10243) );
  AND2_X1 U6600 ( .A1(n6637), .A2(n5809), .ZN(n10178) );
  INV_X1 U6601 ( .A(n9417), .ZN(n6949) );
  INV_X1 U6602 ( .A(n9384), .ZN(n9427) );
  AND2_X1 U6603 ( .A1(n6147), .A2(n6146), .ZN(n9622) );
  NOR2_X1 U6604 ( .A1(n6967), .A2(P1_U3084), .ZN(n7160) );
  INV_X1 U6605 ( .A(n10023), .ZN(n10003) );
  INV_X1 U6606 ( .A(n10138), .ZN(n10161) );
  INV_X1 U6607 ( .A(n10040), .ZN(n10168) );
  INV_X1 U6608 ( .A(n9691), .ZN(n9741) );
  INV_X1 U6609 ( .A(n9725), .ZN(n9713) );
  AOI21_X1 U6610 ( .B1(n7037), .B2(n7039), .A(n7040), .ZN(n7611) );
  AND2_X1 U6611 ( .A1(n6265), .A2(n6482), .ZN(n10040) );
  OR2_X1 U6612 ( .A1(n6473), .A2(n6608), .ZN(n10089) );
  AND3_X1 U6613 ( .A1(n7613), .A2(n6320), .A3(n6319), .ZN(n6322) );
  AND2_X1 U6614 ( .A1(n6954), .A2(n6719), .ZN(n6932) );
  AND2_X1 U6615 ( .A1(n6050), .A2(n6061), .ZN(n7829) );
  INV_X1 U6616 ( .A(n7967), .ZN(n8922) );
  INV_X1 U6617 ( .A(n5846), .ZN(n5847) );
  OR2_X1 U6618 ( .A1(n8549), .A2(n8568), .ZN(n8473) );
  OR2_X1 U6619 ( .A1(n7403), .A2(n9100), .ZN(n8543) );
  INV_X1 U6620 ( .A(n8964), .ZN(n8771) );
  NAND2_X1 U6621 ( .A1(n6702), .A2(n6644), .ZN(n8917) );
  OR2_X1 U6622 ( .A1(n7589), .A2(n7308), .ZN(n10261) );
  INV_X2 U6623 ( .A(n10261), .ZN(n10263) );
  OR2_X1 U6624 ( .A1(n9216), .A2(n9215), .ZN(n9263) );
  OR2_X1 U6625 ( .A1(n7589), .A2(n7259), .ZN(n10253) );
  INV_X1 U6626 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10526) );
  CLKBUF_X1 U6627 ( .A(n8366), .Z(n9281) );
  INV_X1 U6628 ( .A(n9279), .ZN(n8368) );
  NAND2_X1 U6629 ( .A1(n6934), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9429) );
  NAND2_X1 U6630 ( .A1(n9365), .A2(n10163), .ZN(n9417) );
  INV_X1 U6631 ( .A(n9548), .ZN(n9783) );
  INV_X1 U6632 ( .A(n9792), .ZN(n9435) );
  INV_X1 U6633 ( .A(n9834), .ZN(n9695) );
  OR2_X1 U6634 ( .A1(n7165), .A2(n7159), .ZN(n10017) );
  INV_X1 U6635 ( .A(n10013), .ZN(n9994) );
  OR2_X1 U6636 ( .A1(P1_U3083), .A2(n6964), .ZN(n10026) );
  AND2_X1 U6637 ( .A1(n7996), .A2(n7619), .ZN(n10120) );
  NAND2_X1 U6638 ( .A1(n9711), .A2(n10045), .ZN(n9738) );
  NAND2_X1 U6639 ( .A1(n10175), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6324) );
  INV_X1 U6640 ( .A(n10177), .ZN(n10175) );
  AND2_X2 U6641 ( .A1(n6322), .A2(n7611), .ZN(n10177) );
  INV_X1 U6642 ( .A(n10588), .ZN(n10586) );
  NAND2_X1 U6643 ( .A1(n7614), .A2(n7038), .ZN(n10073) );
  AND2_X1 U6644 ( .A1(n8335), .A2(n8235), .ZN(n7040) );
  INV_X1 U6645 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n10566) );
  INV_X1 U6646 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7979) );
  INV_X1 U6647 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7238) );
  INV_X1 U6648 ( .A(n8013), .ZN(n9923) );
  NOR2_X1 U6649 ( .A1(n10602), .A2(n10601), .ZN(n10600) );
  NOR2_X1 U6650 ( .A1(n10291), .A2(n10290), .ZN(n10289) );
  INV_X2 U6651 ( .A(n8773), .ZN(P2_U3966) );
  NAND2_X1 U6652 ( .A1(n6710), .A2(n6709), .ZN(P2_U3264) );
  INV_X1 U6653 ( .A(n9445), .ZN(P1_U4006) );
  MUX2_X1 U6654 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n6323), .S(n10588), .Z(
        P1_U3519) );
  NOR2_X1 U6655 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n5067) );
  INV_X1 U6656 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5074) );
  NAND2_X1 U6657 ( .A1(n5075), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5076) );
  NAND2_X1 U6658 ( .A1(n5082), .A2(n5081), .ZN(n5078) );
  NAND2_X1 U6659 ( .A1(n5078), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5080) );
  XNOR2_X1 U6660 ( .A(n5082), .B(n5081), .ZN(n5122) );
  NAND2_X2 U6661 ( .A1(n10207), .A2(n8761), .ZN(n7366) );
  INV_X1 U6662 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5083) );
  NAND3_X1 U6663 ( .A1(n10423), .A2(n5465), .A3(n5083), .ZN(n5089) );
  NOR2_X1 U6664 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n5087) );
  NAND4_X1 U6665 ( .A1(n5087), .A2(n5086), .A3(n5085), .A4(n5084), .ZN(n5088)
         );
  NOR2_X1 U6666 ( .A1(n5089), .A2(n5088), .ZN(n5091) );
  NAND2_X1 U6667 ( .A1(n5829), .A2(n5827), .ZN(n5115) );
  INV_X1 U6668 ( .A(n5115), .ZN(n5092) );
  XNOR2_X2 U6669 ( .A(n5093), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5098) );
  BUF_X2 U6670 ( .A(n5098), .Z(n9276) );
  NAND2_X4 U6671 ( .A1(n9276), .A2(n9278), .ZN(n5733) );
  INV_X1 U6672 ( .A(n5733), .ZN(n5096) );
  NAND2_X1 U6673 ( .A1(n5096), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5104) );
  NAND2_X1 U6674 ( .A1(n5194), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5102) );
  OR2_X2 U6675 ( .A1(n5099), .A2(n5098), .ZN(n5204) );
  INV_X1 U6676 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6651) );
  INV_X2 U6677 ( .A(n5291), .ZN(n5318) );
  MUX2_X1 U6678 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n5318), .Z(n5112) );
  INV_X1 U6679 ( .A(n5112), .ZN(n5110) );
  INV_X1 U6680 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5106) );
  INV_X1 U6681 ( .A(SI_0_), .ZN(n5135) );
  INV_X1 U6682 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5105) );
  NAND2_X1 U6683 ( .A1(n5107), .A2(SI_1_), .ZN(n5142) );
  INV_X1 U6684 ( .A(SI_1_), .ZN(n5147) );
  NAND2_X1 U6685 ( .A1(n5108), .A2(n5147), .ZN(n5109) );
  NAND2_X1 U6686 ( .A1(n5142), .A2(n5109), .ZN(n5111) );
  NAND2_X1 U6687 ( .A1(n5110), .A2(n5111), .ZN(n5114) );
  INV_X1 U6688 ( .A(n5111), .ZN(n5113) );
  NAND2_X1 U6689 ( .A1(n5113), .A2(n5112), .ZN(n5144) );
  NAND2_X1 U6690 ( .A1(n6643), .A2(n5115), .ZN(n5119) );
  NOR2_X1 U6691 ( .A1(n9271), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n5116) );
  NAND2_X1 U6692 ( .A1(n5117), .A2(n5116), .ZN(n5118) );
  NAND2_X1 U6693 ( .A1(n6645), .A2(n5291), .ZN(n5250) );
  INV_X2 U6694 ( .A(n6645), .ZN(n6695) );
  XNOR2_X1 U6695 ( .A(n5120), .B(P2_IR_REG_1__SCAN_IN), .ZN(n8795) );
  NAND2_X1 U6696 ( .A1(n6695), .A2(n8795), .ZN(n5121) );
  NAND2_X1 U6697 ( .A1(n8765), .A2(n8591), .ZN(n8596) );
  NAND2_X1 U6698 ( .A1(n7550), .A2(n8608), .ZN(n7595) );
  NAND2_X1 U6699 ( .A1(n5123), .A2(n5124), .ZN(n5127) );
  INV_X1 U6700 ( .A(n5123), .ZN(n5126) );
  NAND2_X1 U6701 ( .A1(n5126), .A2(n5125), .ZN(n5137) );
  NAND2_X1 U6702 ( .A1(n5127), .A2(n5137), .ZN(n8372) );
  NAND2_X1 U6703 ( .A1(n5194), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5129) );
  INV_X1 U6704 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n7241) );
  NAND2_X1 U6705 ( .A1(n5129), .A2(n5128), .ZN(n5131) );
  INV_X1 U6706 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n7240) );
  NAND2_X1 U6707 ( .A1(n5096), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5132) );
  XNOR2_X1 U6708 ( .A(n5136), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9283) );
  INV_X1 U6709 ( .A(n9145), .ZN(n10206) );
  NAND2_X1 U6710 ( .A1(n8374), .A2(n10206), .ZN(n9132) );
  OAI22_X1 U6711 ( .A1(n9132), .A2(n8568), .B1(n10206), .B2(n5747), .ZN(n8371)
         );
  OAI21_X1 U6712 ( .B1(n5244), .B2(n5139), .A(n5138), .ZN(n5140) );
  NAND2_X1 U6713 ( .A1(n5140), .A2(SI_2_), .ZN(n5181) );
  OAI21_X1 U6714 ( .B1(n5140), .B2(SI_2_), .A(n5181), .ZN(n5141) );
  AND2_X1 U6715 ( .A1(n5142), .A2(n5141), .ZN(n5143) );
  NAND2_X1 U6716 ( .A1(n5144), .A2(n5143), .ZN(n5158) );
  XNOR2_X1 U6717 ( .A(n5139), .B(SI_2_), .ZN(n5150) );
  INV_X1 U6718 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8367) );
  NAND2_X1 U6719 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5145) );
  NAND2_X1 U6720 ( .A1(n8367), .A2(n5145), .ZN(n5149) );
  NAND2_X1 U6721 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(P1_DATAO_REG_1__SCAN_IN), 
        .ZN(n5146) );
  NAND2_X1 U6722 ( .A1(n5147), .A2(n5146), .ZN(n5148) );
  NAND3_X1 U6723 ( .A1(n5150), .A2(n5149), .A3(n5148), .ZN(n5151) );
  NAND2_X1 U6724 ( .A1(n5291), .A2(n5151), .ZN(n5157) );
  INV_X1 U6725 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8363) );
  NAND2_X1 U6726 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n5152) );
  NAND2_X1 U6727 ( .A1(n8363), .A2(n5152), .ZN(n5153) );
  AOI22_X1 U6728 ( .A1(n5153), .A2(SI_1_), .B1(P2_DATAO_REG_1__SCAN_IN), .B2(
        P2_DATAO_REG_0__SCAN_IN), .ZN(n5155) );
  XNOR2_X1 U6729 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(SI_2_), .ZN(n5154) );
  NAND2_X1 U6730 ( .A1(n5157), .A2(n5156), .ZN(n5182) );
  NAND2_X1 U6731 ( .A1(n5158), .A2(n5182), .ZN(n7000) );
  NAND2_X1 U6732 ( .A1(n5210), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5161) );
  INV_X1 U6733 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5160) );
  OR2_X1 U6734 ( .A1(n5161), .A2(n5160), .ZN(n5162) );
  NAND2_X1 U6735 ( .A1(n5161), .A2(n5160), .ZN(n5188) );
  AND2_X1 U6736 ( .A1(n5162), .A2(n5188), .ZN(n8805) );
  NAND2_X1 U6737 ( .A1(n6695), .A2(n8805), .ZN(n5164) );
  NAND2_X1 U6738 ( .A1(n5251), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5163) );
  AND3_X2 U6739 ( .A1(n5165), .A2(n5164), .A3(n5163), .ZN(n10222) );
  XNOR2_X1 U6740 ( .A(n5747), .B(n10222), .ZN(n5173) );
  NAND2_X1 U6741 ( .A1(n5166), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5172) );
  INV_X1 U6742 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6650) );
  OR2_X1 U6743 ( .A1(n5204), .A2(n6650), .ZN(n5171) );
  INV_X1 U6744 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5167) );
  INV_X1 U6745 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5168) );
  OR2_X1 U6746 ( .A1(n5304), .A2(n5168), .ZN(n5169) );
  NAND2_X1 U6747 ( .A1(n7366), .A2(n8791), .ZN(n5174) );
  XNOR2_X1 U6748 ( .A(n5173), .B(n5174), .ZN(n7361) );
  INV_X1 U6749 ( .A(n5178), .ZN(n5180) );
  INV_X1 U6750 ( .A(SI_3_), .ZN(n5179) );
  NAND2_X1 U6751 ( .A1(n5180), .A2(n5179), .ZN(n5236) );
  NAND2_X1 U6752 ( .A1(n5238), .A2(n5236), .ZN(n5184) );
  INV_X1 U6753 ( .A(n5184), .ZN(n5183) );
  NAND2_X1 U6754 ( .A1(n5182), .A2(n5181), .ZN(n5237) );
  NAND2_X1 U6755 ( .A1(n5183), .A2(n5237), .ZN(n5215) );
  INV_X1 U6756 ( .A(n5237), .ZN(n5185) );
  NAND2_X1 U6757 ( .A1(n5185), .A2(n5184), .ZN(n5186) );
  NAND2_X1 U6758 ( .A1(n5215), .A2(n5186), .ZN(n7012) );
  INV_X1 U6759 ( .A(n7012), .ZN(n5187) );
  NAND2_X1 U6760 ( .A1(n5294), .A2(n5187), .ZN(n5192) );
  NAND2_X1 U6761 ( .A1(n5251), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n5191) );
  NAND2_X1 U6762 ( .A1(n5188), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5189) );
  XNOR2_X1 U6763 ( .A(n5189), .B(P2_IR_REG_3__SCAN_IN), .ZN(n8821) );
  NAND2_X1 U6764 ( .A1(n6695), .A2(n8821), .ZN(n5190) );
  INV_X1 U6765 ( .A(n7604), .ZN(n7342) );
  XNOR2_X1 U6766 ( .A(n7342), .B(n5747), .ZN(n5199) );
  NAND2_X1 U6767 ( .A1(n5166), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5198) );
  INV_X1 U6768 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6657) );
  OR2_X1 U6769 ( .A1(n7049), .A2(n6657), .ZN(n5197) );
  OR2_X1 U6770 ( .A1(n5733), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5196) );
  NAND2_X1 U6771 ( .A1(n7047), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5195) );
  NAND4_X2 U6772 ( .A1(n5198), .A2(n5197), .A3(n5196), .A4(n5195), .ZN(n7343)
         );
  NAND2_X1 U6773 ( .A1(n7366), .A2(n7343), .ZN(n5201) );
  XNOR2_X1 U6774 ( .A(n5199), .B(n5201), .ZN(n7325) );
  NAND2_X1 U6775 ( .A1(n7326), .A2(n7325), .ZN(n5203) );
  INV_X1 U6776 ( .A(n5199), .ZN(n5200) );
  OR2_X1 U6777 ( .A1(n5201), .A2(n5200), .ZN(n5202) );
  NAND2_X1 U6778 ( .A1(n5203), .A2(n5202), .ZN(n7335) );
  NAND2_X1 U6779 ( .A1(n5166), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5209) );
  INV_X1 U6780 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6658) );
  OAI21_X1 U6781 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5229), .ZN(n7641) );
  OR2_X1 U6782 ( .A1(n5733), .A2(n7641), .ZN(n5207) );
  INV_X1 U6783 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n5205) );
  OR2_X1 U6784 ( .A1(n5304), .A2(n5205), .ZN(n5206) );
  AND2_X1 U6785 ( .A1(n7366), .A2(n8790), .ZN(n5225) );
  INV_X2 U6786 ( .A(n5747), .ZN(n5780) );
  NOR2_X1 U6787 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5211) );
  NAND2_X1 U6788 ( .A1(n5213), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5212) );
  MUX2_X1 U6789 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5212), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5214) );
  AND2_X1 U6790 ( .A1(n5214), .A2(n5271), .ZN(n8834) );
  AOI22_X1 U6791 ( .A1(n4408), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6695), .B2(
        n8834), .ZN(n5223) );
  NAND2_X1 U6792 ( .A1(n5215), .A2(n5238), .ZN(n5221) );
  INV_X1 U6793 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7008) );
  INV_X1 U6794 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6990) );
  INV_X1 U6795 ( .A(SI_4_), .ZN(n5217) );
  INV_X1 U6796 ( .A(n5218), .ZN(n5219) );
  NAND2_X1 U6797 ( .A1(n5219), .A2(SI_4_), .ZN(n5242) );
  NAND2_X1 U6798 ( .A1(n5239), .A2(n5242), .ZN(n5220) );
  XNOR2_X1 U6799 ( .A(n5221), .B(n5220), .ZN(n6989) );
  NAND2_X1 U6800 ( .A1(n6989), .A2(n5294), .ZN(n5222) );
  XNOR2_X1 U6801 ( .A(n5780), .B(n10227), .ZN(n5224) );
  AND2_X1 U6802 ( .A1(n5225), .A2(n5224), .ZN(n7333) );
  INV_X1 U6803 ( .A(n5224), .ZN(n5227) );
  INV_X1 U6804 ( .A(n5225), .ZN(n5226) );
  NAND2_X1 U6805 ( .A1(n5227), .A2(n5226), .ZN(n7331) );
  OAI21_X1 U6806 ( .B1(n7335), .B2(n7333), .A(n7331), .ZN(n7407) );
  NAND2_X1 U6807 ( .A1(n5166), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5235) );
  INV_X1 U6808 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6661) );
  OR2_X1 U6809 ( .A1(n7049), .A2(n6661), .ZN(n5234) );
  INV_X1 U6810 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10418) );
  NAND2_X1 U6811 ( .A1(n5229), .A2(n10418), .ZN(n5230) );
  NAND2_X1 U6812 ( .A1(n5300), .A2(n5230), .ZN(n7808) );
  OR2_X1 U6813 ( .A1(n5733), .A2(n7808), .ZN(n5233) );
  INV_X1 U6814 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5231) );
  OR2_X1 U6815 ( .A1(n5304), .A2(n5231), .ZN(n5232) );
  NAND4_X1 U6816 ( .A1(n5235), .A2(n5234), .A3(n5233), .A4(n5232), .ZN(n8789)
         );
  AND2_X1 U6817 ( .A1(n7366), .A2(n8789), .ZN(n5255) );
  NAND3_X1 U6818 ( .A1(n5237), .A2(n5239), .A3(n5236), .ZN(n5243) );
  INV_X1 U6819 ( .A(n5238), .ZN(n5240) );
  NAND2_X1 U6820 ( .A1(n5240), .A2(n5239), .ZN(n5241) );
  NAND2_X1 U6821 ( .A1(n5245), .A2(SI_5_), .ZN(n5259) );
  OAI21_X1 U6822 ( .B1(n5245), .B2(SI_5_), .A(n5259), .ZN(n5247) );
  NAND2_X1 U6823 ( .A1(n5246), .A2(n5247), .ZN(n5249) );
  NAND2_X1 U6824 ( .A1(n5249), .A2(n5260), .ZN(n7009) );
  OR2_X1 U6825 ( .A1(n7009), .A2(n5250), .ZN(n5254) );
  NAND2_X1 U6826 ( .A1(n5271), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5252) );
  XNOR2_X1 U6827 ( .A(n5252), .B(P2_IR_REG_5__SCAN_IN), .ZN(n7373) );
  AOI22_X1 U6828 ( .A1(n4408), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6695), .B2(
        n7373), .ZN(n5253) );
  XNOR2_X1 U6829 ( .A(n5780), .B(n7412), .ZN(n7435) );
  NAND2_X1 U6830 ( .A1(n5255), .A2(n7435), .ZN(n5284) );
  INV_X1 U6831 ( .A(n7435), .ZN(n5257) );
  INV_X1 U6832 ( .A(n5255), .ZN(n5256) );
  NAND2_X1 U6833 ( .A1(n5257), .A2(n5256), .ZN(n5258) );
  NAND2_X1 U6834 ( .A1(n5284), .A2(n5258), .ZN(n7408) );
  INV_X1 U6835 ( .A(n5264), .ZN(n5266) );
  INV_X1 U6836 ( .A(SI_6_), .ZN(n5265) );
  NAND2_X1 U6837 ( .A1(n5266), .A2(n5265), .ZN(n5350) );
  NAND2_X1 U6838 ( .A1(n5340), .A2(n5350), .ZN(n5267) );
  NAND2_X1 U6839 ( .A1(n5343), .A2(n5267), .ZN(n5270) );
  INV_X1 U6840 ( .A(n5343), .ZN(n5269) );
  INV_X1 U6841 ( .A(n5267), .ZN(n5268) );
  AND2_X1 U6842 ( .A1(n5270), .A2(n5290), .ZN(n6992) );
  NAND2_X1 U6843 ( .A1(n6992), .A2(n8398), .ZN(n5278) );
  INV_X1 U6844 ( .A(n5271), .ZN(n5273) );
  NAND2_X1 U6845 ( .A1(n5275), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5274) );
  MUX2_X1 U6846 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5274), .S(
        P2_IR_REG_6__SCAN_IN), .Z(n5276) );
  AND2_X1 U6847 ( .A1(n5276), .A2(n5324), .ZN(n8849) );
  AOI22_X1 U6848 ( .A1(n4408), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6695), .B2(
        n8849), .ZN(n5277) );
  XNOR2_X1 U6849 ( .A(n10232), .B(n5780), .ZN(n5286) );
  NAND2_X1 U6850 ( .A1(n5166), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5283) );
  INV_X1 U6851 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6664) );
  OR2_X1 U6852 ( .A1(n7049), .A2(n6664), .ZN(n5282) );
  INV_X1 U6853 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5299) );
  XNOR2_X1 U6854 ( .A(n5300), .B(n5299), .ZN(n7874) );
  OR2_X1 U6855 ( .A1(n5733), .A2(n7874), .ZN(n5281) );
  INV_X1 U6856 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n5279) );
  OR2_X1 U6857 ( .A1(n5304), .A2(n5279), .ZN(n5280) );
  NAND4_X1 U6858 ( .A1(n5283), .A2(n5282), .A3(n5281), .A4(n5280), .ZN(n8788)
         );
  NAND2_X1 U6859 ( .A1(n7366), .A2(n8788), .ZN(n5287) );
  XNOR2_X1 U6860 ( .A(n5286), .B(n5287), .ZN(n7442) );
  AND2_X1 U6861 ( .A1(n7442), .A2(n5284), .ZN(n5285) );
  INV_X1 U6862 ( .A(n5286), .ZN(n5288) );
  NAND2_X1 U6863 ( .A1(n5288), .A2(n5287), .ZN(n5289) );
  XNOR2_X1 U6864 ( .A(n5344), .B(SI_7_), .ZN(n5293) );
  NAND2_X1 U6865 ( .A1(n7015), .A2(n5294), .ZN(n5297) );
  NAND2_X1 U6866 ( .A1(n5324), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5295) );
  XNOR2_X1 U6867 ( .A(n5295), .B(P2_IR_REG_7__SCAN_IN), .ZN(n8863) );
  AOI22_X1 U6868 ( .A1(n4408), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6695), .B2(
        n8863), .ZN(n5296) );
  NAND2_X1 U6869 ( .A1(n5297), .A2(n5296), .ZN(n10237) );
  XNOR2_X1 U6870 ( .A(n10237), .B(n5747), .ZN(n5310) );
  NAND2_X1 U6871 ( .A1(n5166), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5309) );
  INV_X1 U6872 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6667) );
  OR2_X1 U6873 ( .A1(n7049), .A2(n6667), .ZN(n5308) );
  INV_X1 U6874 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5298) );
  OAI21_X1 U6875 ( .B1(n5300), .B2(n5299), .A(n5298), .ZN(n5303) );
  NAND2_X1 U6876 ( .A1(n5303), .A2(n5331), .ZN(n7843) );
  OR2_X1 U6877 ( .A1(n5733), .A2(n7843), .ZN(n5307) );
  INV_X1 U6878 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n5305) );
  OR2_X1 U6879 ( .A1(n5736), .A2(n5305), .ZN(n5306) );
  NOR2_X1 U6880 ( .A1(n7883), .A2(n8568), .ZN(n5311) );
  NAND2_X1 U6881 ( .A1(n5310), .A2(n5311), .ZN(n5415) );
  INV_X1 U6882 ( .A(n5310), .ZN(n7496) );
  INV_X1 U6883 ( .A(n5311), .ZN(n5312) );
  NAND2_X1 U6884 ( .A1(n7496), .A2(n5312), .ZN(n5313) );
  AND2_X1 U6885 ( .A1(n5415), .A2(n5313), .ZN(n7466) );
  NAND2_X1 U6886 ( .A1(n5314), .A2(SI_7_), .ZN(n5315) );
  NAND2_X1 U6887 ( .A1(n5316), .A2(n5315), .ZN(n5323) );
  INV_X1 U6888 ( .A(n5319), .ZN(n5321) );
  INV_X1 U6889 ( .A(SI_8_), .ZN(n5320) );
  NAND2_X1 U6890 ( .A1(n5321), .A2(n5320), .ZN(n5349) );
  NAND2_X1 U6891 ( .A1(n5347), .A2(n5349), .ZN(n5322) );
  NAND2_X1 U6892 ( .A1(n7028), .A2(n8398), .ZN(n5329) );
  NAND2_X1 U6893 ( .A1(n5326), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5325) );
  MUX2_X1 U6894 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5325), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5327) );
  AOI22_X1 U6895 ( .A1(n4408), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6695), .B2(
        n8879), .ZN(n5328) );
  XNOR2_X1 U6896 ( .A(n10244), .B(n5747), .ZN(n7517) );
  NAND2_X1 U6897 ( .A1(n5166), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5337) );
  INV_X1 U6898 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6670) );
  OR2_X1 U6899 ( .A1(n7049), .A2(n6670), .ZN(n5336) );
  INV_X1 U6900 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10344) );
  NAND2_X1 U6901 ( .A1(n5331), .A2(n10344), .ZN(n5332) );
  NAND2_X1 U6902 ( .A1(n5382), .A2(n5332), .ZN(n7893) );
  OR2_X1 U6903 ( .A1(n5733), .A2(n7893), .ZN(n5335) );
  INV_X1 U6904 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5333) );
  OR2_X1 U6905 ( .A1(n5736), .A2(n5333), .ZN(n5334) );
  NOR2_X1 U6906 ( .A1(n7577), .A2(n8568), .ZN(n5338) );
  NAND2_X1 U6907 ( .A1(n7517), .A2(n5338), .ZN(n5413) );
  OR2_X1 U6908 ( .A1(n7517), .A2(n5338), .ZN(n5339) );
  AND2_X1 U6909 ( .A1(n5413), .A2(n5339), .ZN(n5414) );
  AND2_X1 U6910 ( .A1(n7466), .A2(n5414), .ZN(n7497) );
  INV_X1 U6911 ( .A(n5340), .ZN(n5341) );
  NOR2_X1 U6912 ( .A1(n5351), .A2(n5341), .ZN(n5342) );
  INV_X1 U6913 ( .A(n5344), .ZN(n5346) );
  INV_X1 U6914 ( .A(SI_7_), .ZN(n5345) );
  NAND3_X1 U6915 ( .A1(n5347), .A2(n5346), .A3(n5345), .ZN(n5348) );
  OAI211_X1 U6916 ( .C1(n5351), .C2(n5350), .A(n5349), .B(n5348), .ZN(n5352)
         );
  INV_X1 U6917 ( .A(n5352), .ZN(n5353) );
  NAND2_X1 U6918 ( .A1(n5354), .A2(n5353), .ZN(n5369) );
  INV_X1 U6919 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n7004) );
  INV_X1 U6920 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5355) );
  MUX2_X1 U6921 ( .A(n7004), .B(n5355), .S(n6998), .Z(n5357) );
  INV_X1 U6922 ( .A(SI_9_), .ZN(n5356) );
  NAND2_X1 U6923 ( .A1(n5357), .A2(n5356), .ZN(n5370) );
  INV_X1 U6924 ( .A(n5357), .ZN(n5358) );
  NAND2_X1 U6925 ( .A1(n5358), .A2(SI_9_), .ZN(n5359) );
  XNOR2_X1 U6926 ( .A(n5369), .B(n5053), .ZN(n6994) );
  NAND2_X1 U6927 ( .A1(n6994), .A2(n8398), .ZN(n5362) );
  NAND2_X1 U6928 ( .A1(n5376), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5360) );
  XNOR2_X1 U6929 ( .A(n5360), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6675) );
  AOI22_X1 U6930 ( .A1(n4408), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6675), .B2(
        n6695), .ZN(n5361) );
  NAND2_X1 U6931 ( .A1(n5362), .A2(n5361), .ZN(n7904) );
  XNOR2_X1 U6932 ( .A(n7904), .B(n5780), .ZN(n5412) );
  NAND2_X1 U6933 ( .A1(n5166), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5367) );
  INV_X1 U6934 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6674) );
  OR2_X1 U6935 ( .A1(n7049), .A2(n6674), .ZN(n5366) );
  INV_X1 U6936 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5380) );
  XNOR2_X1 U6937 ( .A(n5382), .B(n5380), .ZN(n7899) );
  OR2_X1 U6938 ( .A1(n5733), .A2(n7899), .ZN(n5365) );
  INV_X1 U6939 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5363) );
  OR2_X1 U6940 ( .A1(n5736), .A2(n5363), .ZN(n5364) );
  NOR2_X1 U6941 ( .A1(n7884), .A2(n8568), .ZN(n5411) );
  INV_X1 U6942 ( .A(n5411), .ZN(n5368) );
  NAND2_X1 U6943 ( .A1(n5412), .A2(n5368), .ZN(n5410) );
  AND2_X1 U6944 ( .A1(n7497), .A2(n5410), .ZN(n7702) );
  NAND2_X1 U6945 ( .A1(n5369), .A2(n5053), .ZN(n5371) );
  MUX2_X1 U6946 ( .A(n7025), .B(n10506), .S(n6998), .Z(n5373) );
  INV_X1 U6947 ( .A(SI_10_), .ZN(n5372) );
  NAND2_X1 U6948 ( .A1(n5373), .A2(n5372), .ZN(n5394) );
  INV_X1 U6949 ( .A(n5373), .ZN(n5374) );
  NAND2_X1 U6950 ( .A1(n5374), .A2(SI_10_), .ZN(n5375) );
  XNOR2_X1 U6951 ( .A(n5393), .B(n5052), .ZN(n7013) );
  NAND2_X1 U6952 ( .A1(n7013), .A2(n8398), .ZN(n5378) );
  XNOR2_X1 U6953 ( .A(n5398), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6678) );
  AOI22_X1 U6954 ( .A1(n6695), .A2(n6678), .B1(n4408), .B2(
        P1_DATAO_REG_10__SCAN_IN), .ZN(n5377) );
  NAND2_X1 U6955 ( .A1(n5378), .A2(n5377), .ZN(n7915) );
  XNOR2_X1 U6956 ( .A(n7915), .B(n5747), .ZN(n7701) );
  NAND2_X1 U6957 ( .A1(n5166), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5388) );
  INV_X1 U6958 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10524) );
  OR2_X1 U6959 ( .A1(n7049), .A2(n10524), .ZN(n5387) );
  INV_X1 U6960 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n5379) );
  OAI21_X1 U6961 ( .B1(n5382), .B2(n5380), .A(n5379), .ZN(n5383) );
  NAND2_X1 U6962 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n5381) );
  OR2_X2 U6963 ( .A1(n5382), .A2(n5381), .ZN(n5401) );
  NAND2_X1 U6964 ( .A1(n5383), .A2(n5401), .ZN(n7910) );
  OR2_X1 U6965 ( .A1(n5733), .A2(n7910), .ZN(n5386) );
  INV_X1 U6966 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5384) );
  OR2_X1 U6967 ( .A1(n5736), .A2(n5384), .ZN(n5385) );
  NOR2_X1 U6968 ( .A1(n7654), .A2(n8568), .ZN(n5389) );
  NAND2_X1 U6969 ( .A1(n7701), .A2(n5389), .ZN(n5418) );
  INV_X1 U6970 ( .A(n7701), .ZN(n5391) );
  INV_X1 U6971 ( .A(n5389), .ZN(n5390) );
  NAND2_X1 U6972 ( .A1(n5391), .A2(n5390), .ZN(n5392) );
  NAND2_X1 U6973 ( .A1(n5418), .A2(n5392), .ZN(n7817) );
  NAND2_X1 U6974 ( .A1(n5393), .A2(n5052), .ZN(n5395) );
  MUX2_X1 U6975 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6998), .Z(n5421) );
  XNOR2_X1 U6976 ( .A(n5421), .B(SI_11_), .ZN(n5423) );
  INV_X1 U6977 ( .A(n5423), .ZN(n5396) );
  XNOR2_X1 U6978 ( .A(n5424), .B(n5396), .ZN(n7026) );
  INV_X1 U6979 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5397) );
  XNOR2_X1 U6980 ( .A(n5399), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6682) );
  NAND2_X1 U6981 ( .A1(n7019), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5407) );
  INV_X1 U6982 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7948) );
  OR2_X1 U6983 ( .A1(n7052), .A2(n7948), .ZN(n5406) );
  INV_X1 U6984 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7317) );
  NAND2_X1 U6985 ( .A1(n5401), .A2(n7317), .ZN(n5402) );
  NAND2_X1 U6986 ( .A1(n5451), .A2(n5402), .ZN(n7950) );
  OR2_X1 U6987 ( .A1(n5733), .A2(n7950), .ZN(n5405) );
  INV_X1 U6988 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n5403) );
  OR2_X1 U6989 ( .A1(n5736), .A2(n5403), .ZN(n5404) );
  NOR2_X1 U6990 ( .A1(n7820), .A2(n8568), .ZN(n5408) );
  NAND2_X1 U6991 ( .A1(n5459), .A2(n5408), .ZN(n7679) );
  INV_X1 U6992 ( .A(n5408), .ZN(n5458) );
  NAND2_X1 U6993 ( .A1(n7674), .A2(n5458), .ZN(n5409) );
  AND2_X1 U6994 ( .A1(n7679), .A2(n5409), .ZN(n7705) );
  OR2_X1 U6995 ( .A1(n5416), .A2(n7704), .ZN(n5417) );
  OR2_X1 U6996 ( .A1(n5419), .A2(n5418), .ZN(n5420) );
  NAND2_X1 U6997 ( .A1(n5421), .A2(SI_11_), .ZN(n5422) );
  MUX2_X1 U6998 ( .A(n7045), .B(n10446), .S(n6998), .Z(n5426) );
  INV_X1 U6999 ( .A(n5426), .ZN(n5427) );
  NAND2_X1 U7000 ( .A1(n5427), .A2(SI_12_), .ZN(n5428) );
  MUX2_X1 U7001 ( .A(n10316), .B(n10514), .S(n6998), .Z(n5432) );
  INV_X1 U7002 ( .A(SI_13_), .ZN(n5431) );
  INV_X1 U7003 ( .A(n5432), .ZN(n5433) );
  NAND2_X1 U7004 ( .A1(n5433), .A2(SI_13_), .ZN(n5434) );
  NAND2_X1 U7005 ( .A1(n7054), .A2(n8398), .ZN(n5439) );
  INV_X1 U7006 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5435) );
  NAND2_X1 U7007 ( .A1(n5467), .A2(n5435), .ZN(n5436) );
  NAND2_X1 U7008 ( .A1(n5436), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5437) );
  XNOR2_X1 U7009 ( .A(n5437), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7513) );
  AOI22_X1 U7010 ( .A1(n4408), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6695), .B2(
        n7513), .ZN(n5438) );
  XNOR2_X1 U7011 ( .A(n9232), .B(n5780), .ZN(n8096) );
  NAND2_X1 U7012 ( .A1(n7047), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5445) );
  INV_X1 U7013 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7759) );
  OR2_X1 U7014 ( .A1(n7052), .A2(n7759), .ZN(n5444) );
  INV_X1 U7015 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10527) );
  OR2_X1 U7016 ( .A1(n7049), .A2(n10527), .ZN(n5443) );
  INV_X1 U7017 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10570) );
  NAND2_X1 U7018 ( .A1(n5453), .A2(n10570), .ZN(n5441) );
  NAND2_X1 U7019 ( .A1(n5472), .A2(n5441), .ZN(n8115) );
  OR2_X1 U7020 ( .A1(n5733), .A2(n8115), .ZN(n5442) );
  NAND4_X1 U7021 ( .A1(n5445), .A2(n5444), .A3(n5443), .A4(n5442), .ZN(n8781)
         );
  NAND2_X1 U7022 ( .A1(n7366), .A2(n8781), .ZN(n5478) );
  NAND2_X1 U7023 ( .A1(n8096), .A2(n5478), .ZN(n8095) );
  XNOR2_X1 U7024 ( .A(n5447), .B(n5446), .ZN(n7042) );
  NAND2_X1 U7025 ( .A1(n7042), .A2(n8398), .ZN(n5449) );
  XNOR2_X1 U7026 ( .A(n5467), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6683) );
  AOI22_X1 U7027 ( .A1(n4408), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6695), .B2(
        n6683), .ZN(n5448) );
  XNOR2_X1 U7028 ( .A(n9238), .B(n5780), .ZN(n7678) );
  NAND2_X1 U7029 ( .A1(n5166), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5457) );
  INV_X1 U7030 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10435) );
  OR2_X1 U7031 ( .A1(n7049), .A2(n10435), .ZN(n5456) );
  NAND2_X1 U7032 ( .A1(n5451), .A2(n5450), .ZN(n5452) );
  NAND2_X1 U7033 ( .A1(n5453), .A2(n5452), .ZN(n7682) );
  OR2_X1 U7034 ( .A1(n5733), .A2(n7682), .ZN(n5455) );
  INV_X1 U7035 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10504) );
  OR2_X1 U7036 ( .A1(n5736), .A2(n10504), .ZN(n5454) );
  OR2_X1 U7037 ( .A1(n8116), .A2(n8568), .ZN(n7676) );
  NAND2_X1 U7038 ( .A1(n7678), .A2(n7676), .ZN(n8092) );
  NAND2_X1 U7039 ( .A1(n7673), .A2(n5045), .ZN(n5485) );
  INV_X1 U7040 ( .A(n8095), .ZN(n5482) );
  INV_X1 U7041 ( .A(n7678), .ZN(n5462) );
  NAND2_X1 U7042 ( .A1(n7679), .A2(n7676), .ZN(n5461) );
  NOR2_X1 U7043 ( .A1(n7676), .A2(n5458), .ZN(n5460) );
  AOI22_X1 U7044 ( .A1(n5462), .A2(n5461), .B1(n5460), .B2(n5459), .ZN(n5481)
         );
  MUX2_X1 U7045 ( .A(n7086), .B(n10437), .S(n6998), .Z(n5487) );
  NAND2_X1 U7046 ( .A1(n7083), .A2(n8398), .ZN(n5470) );
  OR2_X1 U7047 ( .A1(n5465), .A2(n9271), .ZN(n5466) );
  NAND2_X1 U7048 ( .A1(n5467), .A2(n5466), .ZN(n5517) );
  INV_X1 U7049 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5468) );
  XNOR2_X1 U7050 ( .A(n5517), .B(n5468), .ZN(n7975) );
  AOI22_X1 U7051 ( .A1(n4408), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6695), .B2(
        n7975), .ZN(n5469) );
  XNOR2_X1 U7052 ( .A(n9226), .B(n5780), .ZN(n5532) );
  NAND2_X1 U7053 ( .A1(n7019), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5477) );
  INV_X1 U7054 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6628) );
  OR2_X1 U7055 ( .A1(n7052), .A2(n6628), .ZN(n5476) );
  INV_X1 U7056 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U7057 ( .A1(n5472), .A2(n5471), .ZN(n5473) );
  NAND2_X1 U7058 ( .A1(n5521), .A2(n5473), .ZN(n8099) );
  OR2_X1 U7059 ( .A1(n5733), .A2(n8099), .ZN(n5475) );
  INV_X1 U7060 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10436) );
  OR2_X1 U7061 ( .A1(n5736), .A2(n10436), .ZN(n5474) );
  NOR2_X1 U7062 ( .A1(n8112), .A2(n8568), .ZN(n5530) );
  XNOR2_X1 U7063 ( .A(n5532), .B(n5530), .ZN(n8107) );
  INV_X1 U7064 ( .A(n8096), .ZN(n5480) );
  INV_X1 U7065 ( .A(n5478), .ZN(n5479) );
  NAND2_X1 U7066 ( .A1(n5480), .A2(n5479), .ZN(n8094) );
  OAI211_X1 U7067 ( .C1(n5482), .C2(n5481), .A(n8107), .B(n8094), .ZN(n5483)
         );
  INV_X1 U7068 ( .A(n5483), .ZN(n5484) );
  INV_X1 U7069 ( .A(n5487), .ZN(n5488) );
  INV_X1 U7070 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n5491) );
  MUX2_X1 U7071 ( .A(n10567), .B(n5491), .S(n6344), .Z(n5493) );
  INV_X1 U7072 ( .A(SI_15_), .ZN(n5492) );
  INV_X1 U7073 ( .A(n5493), .ZN(n5494) );
  NAND2_X1 U7074 ( .A1(n5494), .A2(SI_15_), .ZN(n5495) );
  MUX2_X1 U7075 ( .A(n10526), .B(n7238), .S(n6998), .Z(n5498) );
  INV_X1 U7076 ( .A(SI_16_), .ZN(n5497) );
  INV_X1 U7077 ( .A(n5498), .ZN(n5499) );
  NAND2_X1 U7078 ( .A1(n5499), .A2(SI_16_), .ZN(n5500) );
  XNOR2_X1 U7079 ( .A(n5541), .B(n5056), .ZN(n7237) );
  NAND2_X1 U7080 ( .A1(n7237), .A2(n8398), .ZN(n5506) );
  NOR2_X1 U7081 ( .A1(n5501), .A2(n9271), .ZN(n5502) );
  MUX2_X1 U7082 ( .A(n9271), .B(n5502), .S(P2_IR_REG_16__SCAN_IN), .Z(n5504)
         );
  OR2_X1 U7083 ( .A1(n5504), .A2(n4878), .ZN(n8896) );
  INV_X1 U7084 ( .A(n8896), .ZN(n6630) );
  AOI22_X1 U7085 ( .A1(n4408), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6695), .B2(
        n6630), .ZN(n5505) );
  XNOR2_X1 U7086 ( .A(n8279), .B(n5780), .ZN(n8159) );
  INV_X1 U7087 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8224) );
  OR2_X2 U7088 ( .A1(n5521), .A2(n8224), .ZN(n5523) );
  INV_X1 U7089 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U7090 ( .A1(n5523), .A2(n5508), .ZN(n5509) );
  NAND2_X1 U7091 ( .A1(n5548), .A2(n5509), .ZN(n8164) );
  OR2_X1 U7092 ( .A1(n8164), .A2(n5733), .ZN(n5514) );
  INV_X1 U7093 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8146) );
  OR2_X1 U7094 ( .A1(n7052), .A2(n8146), .ZN(n5511) );
  INV_X1 U7095 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8262) );
  OR2_X1 U7096 ( .A1(n7049), .A2(n8262), .ZN(n5510) );
  AND2_X1 U7097 ( .A1(n5511), .A2(n5510), .ZN(n5513) );
  NAND2_X1 U7098 ( .A1(n7047), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5512) );
  INV_X1 U7099 ( .A(n8228), .ZN(n8778) );
  NAND2_X1 U7100 ( .A1(n8778), .A2(n7366), .ZN(n5535) );
  XNOR2_X1 U7101 ( .A(n5515), .B(n5516), .ZN(n7144) );
  NAND2_X1 U7102 ( .A1(n7144), .A2(n8398), .ZN(n5520) );
  OAI21_X1 U7103 ( .B1(n5517), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5518) );
  XNOR2_X1 U7104 ( .A(n5518), .B(P2_IR_REG_15__SCAN_IN), .ZN(n6688) );
  AOI22_X1 U7105 ( .A1(n4408), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6695), .B2(
        n6688), .ZN(n5519) );
  XNOR2_X1 U7106 ( .A(n8127), .B(n5747), .ZN(n5536) );
  NAND2_X1 U7107 ( .A1(n5521), .A2(n8224), .ZN(n5522) );
  AND2_X1 U7108 ( .A1(n5523), .A2(n5522), .ZN(n8225) );
  NAND2_X1 U7109 ( .A1(n5834), .A2(n8225), .ZN(n5529) );
  INV_X1 U7110 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n6690) );
  OR2_X1 U7111 ( .A1(n7049), .A2(n6690), .ZN(n5528) );
  INV_X1 U7112 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5524) );
  OR2_X1 U7113 ( .A1(n7052), .A2(n5524), .ZN(n5527) );
  INV_X1 U7114 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n5525) );
  OR2_X1 U7115 ( .A1(n5736), .A2(n5525), .ZN(n5526) );
  NOR2_X1 U7116 ( .A1(n8155), .A2(n8568), .ZN(n8161) );
  INV_X1 U7117 ( .A(n5530), .ZN(n5531) );
  NAND2_X1 U7118 ( .A1(n5532), .A2(n5531), .ZN(n8154) );
  OAI21_X1 U7119 ( .B1(n5536), .B2(n8161), .A(n8154), .ZN(n5533) );
  AOI21_X1 U7120 ( .B1(n8159), .B2(n5535), .A(n5533), .ZN(n5534) );
  INV_X1 U7121 ( .A(n8159), .ZN(n5539) );
  INV_X1 U7122 ( .A(n5536), .ZN(n8156) );
  INV_X1 U7123 ( .A(n8161), .ZN(n8223) );
  OAI21_X1 U7124 ( .B1(n8156), .B2(n8223), .A(n5535), .ZN(n5538) );
  INV_X1 U7125 ( .A(n5535), .ZN(n8158) );
  AND3_X1 U7126 ( .A1(n5536), .A2(n8161), .A3(n8158), .ZN(n5537) );
  AOI21_X1 U7127 ( .B1(n5539), .B2(n5538), .A(n5537), .ZN(n5540) );
  MUX2_X1 U7128 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n6998), .Z(n5558) );
  XNOR2_X1 U7129 ( .A(n5558), .B(SI_17_), .ZN(n5560) );
  INV_X1 U7130 ( .A(n5560), .ZN(n5543) );
  XNOR2_X1 U7131 ( .A(n5561), .B(n5543), .ZN(n7249) );
  NAND2_X1 U7132 ( .A1(n7249), .A2(n8398), .ZN(n5546) );
  NAND2_X1 U7133 ( .A1(n5503), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5544) );
  XNOR2_X1 U7134 ( .A(n5544), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8905) );
  AOI22_X1 U7135 ( .A1(n4408), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6695), .B2(
        n8905), .ZN(n5545) );
  XNOR2_X1 U7136 ( .A(n8324), .B(n5747), .ZN(n5553) );
  INV_X1 U7137 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n8906) );
  NAND2_X1 U7138 ( .A1(n5548), .A2(n8906), .ZN(n5549) );
  NAND2_X1 U7139 ( .A1(n5567), .A2(n5549), .ZN(n8294) );
  OR2_X1 U7140 ( .A1(n8294), .A2(n5733), .ZN(n5552) );
  AOI22_X1 U7141 ( .A1(n5166), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n7019), .B2(
        P2_REG1_REG_17__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U7142 ( .A1(n7047), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5550) );
  NOR2_X1 U7143 ( .A1(n8283), .A2(n8568), .ZN(n5554) );
  NAND2_X1 U7144 ( .A1(n5553), .A2(n5554), .ZN(n5557) );
  INV_X1 U7145 ( .A(n5553), .ZN(n8211) );
  INV_X1 U7146 ( .A(n5554), .ZN(n5555) );
  NAND2_X1 U7147 ( .A1(n8211), .A2(n5555), .ZN(n5556) );
  AND2_X1 U7148 ( .A1(n5557), .A2(n5556), .ZN(n8121) );
  NAND2_X1 U7149 ( .A1(n8210), .A2(n5557), .ZN(n5572) );
  NAND2_X1 U7150 ( .A1(n5558), .A2(SI_17_), .ZN(n5559) );
  MUX2_X1 U7151 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6344), .Z(n5579) );
  XNOR2_X1 U7152 ( .A(n5562), .B(n5577), .ZN(n7416) );
  NAND2_X1 U7153 ( .A1(n7416), .A2(n8398), .ZN(n5565) );
  XNOR2_X1 U7154 ( .A(n5563), .B(P2_IR_REG_18__SCAN_IN), .ZN(n6648) );
  AOI22_X1 U7155 ( .A1(n4408), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6695), .B2(
        n6648), .ZN(n5564) );
  XNOR2_X1 U7156 ( .A(n9218), .B(n5780), .ZN(n5573) );
  INV_X1 U7157 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5566) );
  OR2_X2 U7158 ( .A1(n5567), .A2(n5566), .ZN(n5589) );
  NAND2_X1 U7159 ( .A1(n5567), .A2(n5566), .ZN(n5568) );
  AND2_X1 U7160 ( .A1(n5589), .A2(n5568), .ZN(n8321) );
  NAND2_X1 U7161 ( .A1(n8321), .A2(n5834), .ZN(n5571) );
  AOI22_X1 U7162 ( .A1(n5166), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n7019), .B2(
        P2_REG1_REG_18__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7163 ( .A1(n7047), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5569) );
  NOR2_X1 U7164 ( .A1(n9101), .A2(n8568), .ZN(n5574) );
  XNOR2_X1 U7165 ( .A(n5573), .B(n5574), .ZN(n8208) );
  NAND2_X1 U7166 ( .A1(n5572), .A2(n8208), .ZN(n8212) );
  INV_X1 U7167 ( .A(n5573), .ZN(n5575) );
  NAND2_X1 U7168 ( .A1(n5575), .A2(n5574), .ZN(n5576) );
  NAND2_X1 U7169 ( .A1(n8212), .A2(n5576), .ZN(n8487) );
  NAND2_X1 U7170 ( .A1(n5562), .A2(n5578), .ZN(n5581) );
  NAND2_X1 U7171 ( .A1(n5579), .A2(SI_18_), .ZN(n5580) );
  MUX2_X1 U7172 ( .A(n7430), .B(n7432), .S(n6998), .Z(n5583) );
  INV_X1 U7173 ( .A(SI_19_), .ZN(n5582) );
  INV_X1 U7174 ( .A(n5583), .ZN(n5584) );
  NAND2_X1 U7175 ( .A1(n5584), .A2(SI_19_), .ZN(n5585) );
  NAND2_X1 U7176 ( .A1(n5599), .A2(n5585), .ZN(n5600) );
  XNOR2_X1 U7177 ( .A(n5601), .B(n5600), .ZN(n7429) );
  NAND2_X1 U7178 ( .A1(n7429), .A2(n8398), .ZN(n5587) );
  AOI22_X1 U7179 ( .A1(n4408), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8591), .B2(
        n6695), .ZN(n5586) );
  XNOR2_X1 U7180 ( .A(n9211), .B(n5747), .ZN(n8484) );
  INV_X1 U7181 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10538) );
  NAND2_X1 U7182 ( .A1(n5589), .A2(n10538), .ZN(n5590) );
  NAND2_X1 U7183 ( .A1(n5625), .A2(n5590), .ZN(n9107) );
  OR2_X1 U7184 ( .A1(n9107), .A2(n5733), .ZN(n5595) );
  INV_X1 U7185 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n10482) );
  NAND2_X1 U7186 ( .A1(n7019), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5592) );
  INV_X1 U7187 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n10564) );
  OR2_X1 U7188 ( .A1(n5736), .A2(n10564), .ZN(n5591) );
  OAI211_X1 U7189 ( .C1(n7052), .C2(n10482), .A(n5592), .B(n5591), .ZN(n5593)
         );
  INV_X1 U7190 ( .A(n5593), .ZN(n5594) );
  NOR2_X1 U7191 ( .A1(n8524), .A2(n8568), .ZN(n5596) );
  AND2_X1 U7192 ( .A1(n8484), .A2(n5596), .ZN(n8482) );
  INV_X1 U7193 ( .A(n8484), .ZN(n5598) );
  INV_X1 U7194 ( .A(n5596), .ZN(n5597) );
  NAND2_X1 U7195 ( .A1(n5598), .A2(n5597), .ZN(n8486) );
  OAI21_X1 U7196 ( .B1(n8487), .B2(n8482), .A(n8486), .ZN(n8523) );
  MUX2_X1 U7197 ( .A(n10434), .B(n7533), .S(n6344), .Z(n5603) );
  INV_X1 U7198 ( .A(SI_20_), .ZN(n5602) );
  NAND2_X1 U7199 ( .A1(n5603), .A2(n5602), .ZN(n5620) );
  INV_X1 U7200 ( .A(n5603), .ZN(n5604) );
  NAND2_X1 U7201 ( .A1(n5604), .A2(SI_20_), .ZN(n5605) );
  XNOR2_X1 U7202 ( .A(n5619), .B(n5618), .ZN(n7532) );
  NAND2_X1 U7203 ( .A1(n7532), .A2(n8398), .ZN(n5607) );
  NAND2_X1 U7204 ( .A1(n4408), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n5606) );
  XNOR2_X1 U7205 ( .A(n9207), .B(n5747), .ZN(n5614) );
  XNOR2_X1 U7206 ( .A(n5625), .B(P2_REG3_REG_20__SCAN_IN), .ZN(n9086) );
  NAND2_X1 U7207 ( .A1(n9086), .A2(n5834), .ZN(n5613) );
  INV_X1 U7208 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U7209 ( .A1(n7047), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7210 ( .A1(n7019), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5608) );
  OAI211_X1 U7211 ( .C1(n7052), .C2(n5610), .A(n5609), .B(n5608), .ZN(n5611)
         );
  INV_X1 U7212 ( .A(n5611), .ZN(n5612) );
  NOR2_X1 U7213 ( .A1(n9103), .A2(n8568), .ZN(n5615) );
  XNOR2_X1 U7214 ( .A(n5614), .B(n5615), .ZN(n8522) );
  INV_X1 U7215 ( .A(n5614), .ZN(n5617) );
  INV_X1 U7216 ( .A(n5615), .ZN(n5616) );
  INV_X1 U7217 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n5621) );
  MUX2_X1 U7218 ( .A(n5621), .B(n7700), .S(n6344), .Z(n5636) );
  XNOR2_X1 U7219 ( .A(n5636), .B(SI_21_), .ZN(n5635) );
  XNOR2_X1 U7220 ( .A(n5634), .B(n5635), .ZN(n7587) );
  NAND2_X1 U7221 ( .A1(n7587), .A2(n8398), .ZN(n5623) );
  NAND2_X1 U7222 ( .A1(n4408), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n5622) );
  XNOR2_X1 U7223 ( .A(n9201), .B(n5780), .ZN(n5672) );
  INV_X1 U7224 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8525) );
  INV_X1 U7225 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5624) );
  OAI21_X1 U7226 ( .B1(n5625), .B2(n8525), .A(n5624), .ZN(n5628) );
  INV_X1 U7227 ( .A(n5625), .ZN(n5627) );
  AND2_X1 U7228 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_20__SCAN_IN), 
        .ZN(n5626) );
  INV_X1 U7229 ( .A(n5645), .ZN(n5646) );
  AND2_X1 U7230 ( .A1(n5628), .A2(n5646), .ZN(n9069) );
  NAND2_X1 U7231 ( .A1(n9069), .A2(n5834), .ZN(n5633) );
  INV_X1 U7232 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n10503) );
  NAND2_X1 U7233 ( .A1(n7019), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U7234 ( .A1(n5166), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5629) );
  OAI211_X1 U7235 ( .C1(n10503), .C2(n5736), .A(n5630), .B(n5629), .ZN(n5631)
         );
  INV_X1 U7236 ( .A(n5631), .ZN(n5632) );
  NOR2_X1 U7237 ( .A1(n9047), .A2(n8568), .ZN(n5674) );
  XNOR2_X1 U7238 ( .A(n5672), .B(n5674), .ZN(n8494) );
  INV_X1 U7239 ( .A(n5636), .ZN(n5637) );
  NAND2_X1 U7240 ( .A1(n5637), .A2(SI_21_), .ZN(n5638) );
  NAND2_X1 U7241 ( .A1(n5639), .A2(n5638), .ZN(n5656) );
  INV_X1 U7242 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n5640) );
  MUX2_X1 U7243 ( .A(n5640), .B(n7979), .S(n6344), .Z(n5642) );
  INV_X1 U7244 ( .A(SI_22_), .ZN(n5641) );
  INV_X1 U7245 ( .A(n5642), .ZN(n5643) );
  NAND2_X1 U7246 ( .A1(n5643), .A2(SI_22_), .ZN(n5644) );
  XNOR2_X1 U7247 ( .A(n8423), .B(n5747), .ZN(n5671) );
  INV_X1 U7248 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10296) );
  NAND2_X1 U7249 ( .A1(n5646), .A2(n10296), .ZN(n5647) );
  NAND2_X1 U7250 ( .A1(n5664), .A2(n5647), .ZN(n9054) );
  OR2_X1 U7251 ( .A1(n9054), .A2(n5733), .ZN(n5653) );
  INV_X1 U7252 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7253 ( .A1(n7019), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U7254 ( .A1(n7047), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5648) );
  OAI211_X1 U7255 ( .C1(n7052), .C2(n5650), .A(n5649), .B(n5648), .ZN(n5651)
         );
  INV_X1 U7256 ( .A(n5651), .ZN(n5652) );
  NAND2_X1 U7257 ( .A1(n5653), .A2(n5652), .ZN(n9066) );
  NAND2_X1 U7258 ( .A1(n9066), .A2(n7366), .ZN(n8537) );
  INV_X1 U7259 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n5657) );
  INV_X1 U7260 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8017) );
  MUX2_X1 U7261 ( .A(n5657), .B(n8017), .S(n6998), .Z(n5659) );
  INV_X1 U7262 ( .A(SI_23_), .ZN(n5658) );
  NAND2_X1 U7263 ( .A1(n5659), .A2(n5658), .ZN(n5684) );
  INV_X1 U7264 ( .A(n5659), .ZN(n5660) );
  NAND2_X1 U7265 ( .A1(n5660), .A2(SI_23_), .ZN(n5661) );
  XNOR2_X1 U7266 ( .A(n5683), .B(n5682), .ZN(n8014) );
  NAND2_X1 U7267 ( .A1(n8014), .A2(n8398), .ZN(n5663) );
  NAND2_X1 U7268 ( .A1(n4408), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n5662) );
  XNOR2_X1 U7269 ( .A(n9036), .B(n5780), .ZN(n5678) );
  INV_X1 U7270 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10329) );
  NAND2_X1 U7271 ( .A1(n5664), .A2(n10329), .ZN(n5665) );
  NAND2_X1 U7272 ( .A1(n5689), .A2(n5665), .ZN(n9033) );
  OR2_X1 U7273 ( .A1(n9033), .A2(n5733), .ZN(n5670) );
  INV_X1 U7274 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n10479) );
  NAND2_X1 U7275 ( .A1(n5166), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5667) );
  INV_X1 U7276 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n10381) );
  OR2_X1 U7277 ( .A1(n5736), .A2(n10381), .ZN(n5666) );
  OAI211_X1 U7278 ( .C1(n7049), .C2(n10479), .A(n5667), .B(n5666), .ZN(n5668)
         );
  INV_X1 U7279 ( .A(n5668), .ZN(n5669) );
  NAND2_X1 U7280 ( .A1(n5670), .A2(n5669), .ZN(n9008) );
  AND2_X1 U7281 ( .A1(n9008), .A2(n7366), .ZN(n5679) );
  INV_X1 U7282 ( .A(n5671), .ZN(n8533) );
  INV_X1 U7283 ( .A(n5672), .ZN(n5675) );
  NAND2_X1 U7284 ( .A1(n5675), .A2(n5674), .ZN(n8531) );
  NAND2_X1 U7285 ( .A1(n8531), .A2(n8537), .ZN(n5673) );
  NAND2_X1 U7286 ( .A1(n8533), .A2(n5673), .ZN(n5677) );
  NAND3_X1 U7287 ( .A1(n5675), .A2(n5674), .A3(n9066), .ZN(n5676) );
  NAND2_X1 U7288 ( .A1(n5677), .A2(n5676), .ZN(n8468) );
  AOI21_X1 U7289 ( .B1(n5678), .B2(n5679), .A(n8468), .ZN(n5681) );
  INV_X1 U7290 ( .A(n5678), .ZN(n8471) );
  INV_X1 U7291 ( .A(n5679), .ZN(n8476) );
  AND2_X1 U7292 ( .A1(n8471), .A2(n8476), .ZN(n5680) );
  NAND2_X1 U7293 ( .A1(n5683), .A2(n5682), .ZN(n5685) );
  INV_X1 U7294 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n5686) );
  MUX2_X1 U7295 ( .A(n5686), .B(n10566), .S(n6344), .Z(n5700) );
  XNOR2_X1 U7296 ( .A(n5700), .B(SI_24_), .ZN(n5699) );
  NAND2_X1 U7297 ( .A1(n4408), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n8424) );
  XOR2_X1 U7298 ( .A(n8428), .B(n5747), .Z(n5696) );
  INV_X1 U7299 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5688) );
  NAND2_X1 U7300 ( .A1(n5689), .A2(n5688), .ZN(n5690) );
  NAND2_X1 U7301 ( .A1(n5712), .A2(n5690), .ZN(n9017) );
  OR2_X1 U7302 ( .A1(n9017), .A2(n5733), .ZN(n5695) );
  INV_X1 U7303 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n10554) );
  NAND2_X1 U7304 ( .A1(n7047), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5692) );
  NAND2_X1 U7305 ( .A1(n4406), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5691) );
  OAI211_X1 U7306 ( .C1(n7049), .C2(n10554), .A(n5692), .B(n5691), .ZN(n5693)
         );
  INV_X1 U7307 ( .A(n5693), .ZN(n5694) );
  NOR2_X1 U7308 ( .A1(n8505), .A2(n8568), .ZN(n8512) );
  INV_X1 U7309 ( .A(n5696), .ZN(n5697) );
  INV_X1 U7310 ( .A(n5700), .ZN(n5701) );
  NAND2_X1 U7311 ( .A1(n5701), .A2(SI_24_), .ZN(n5702) );
  INV_X1 U7312 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n5705) );
  INV_X1 U7313 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8315) );
  MUX2_X1 U7314 ( .A(n5705), .B(n8315), .S(n6463), .Z(n5707) );
  INV_X1 U7315 ( .A(SI_25_), .ZN(n5706) );
  NAND2_X1 U7316 ( .A1(n5707), .A2(n5706), .ZN(n5720) );
  INV_X1 U7317 ( .A(n5707), .ZN(n5708) );
  NAND2_X1 U7318 ( .A1(n5708), .A2(SI_25_), .ZN(n5709) );
  NAND2_X1 U7319 ( .A1(n5720), .A2(n5709), .ZN(n5721) );
  NAND2_X1 U7320 ( .A1(n8267), .A2(n8398), .ZN(n5711) );
  NAND2_X1 U7321 ( .A1(n4408), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n5710) );
  XNOR2_X1 U7322 ( .A(n8429), .B(n5747), .ZN(n5718) );
  INV_X1 U7323 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8506) );
  OR2_X2 U7324 ( .A1(n5712), .A2(n8506), .ZN(n5731) );
  NAND2_X1 U7325 ( .A1(n5712), .A2(n8506), .ZN(n5713) );
  INV_X1 U7326 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n5716) );
  NAND2_X1 U7327 ( .A1(n5166), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5715) );
  NAND2_X1 U7328 ( .A1(n7019), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n5714) );
  OAI211_X1 U7329 ( .C1(n5716), .C2(n5736), .A(n5715), .B(n5714), .ZN(n5717)
         );
  NOR2_X1 U7330 ( .A1(n9012), .A2(n8568), .ZN(n8503) );
  INV_X1 U7331 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n5723) );
  INV_X1 U7332 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8333) );
  MUX2_X1 U7333 ( .A(n5723), .B(n8333), .S(n6344), .Z(n5725) );
  INV_X1 U7334 ( .A(SI_26_), .ZN(n5724) );
  NAND2_X1 U7335 ( .A1(n5725), .A2(n5724), .ZN(n5760) );
  INV_X1 U7336 ( .A(n5725), .ZN(n5726) );
  NAND2_X1 U7337 ( .A1(n5726), .A2(SI_26_), .ZN(n5727) );
  XNOR2_X1 U7338 ( .A(n6332), .B(n5758), .ZN(n8330) );
  NAND2_X1 U7339 ( .A1(n8330), .A2(n8398), .ZN(n5729) );
  NAND2_X1 U7340 ( .A1(n4408), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n5728) );
  XNOR2_X1 U7341 ( .A(n9177), .B(n5747), .ZN(n8459) );
  INV_X1 U7342 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10562) );
  NAND2_X1 U7343 ( .A1(n5731), .A2(n10562), .ZN(n5732) );
  NAND2_X1 U7344 ( .A1(n5772), .A2(n5732), .ZN(n8978) );
  INV_X1 U7345 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n10327) );
  NAND2_X1 U7346 ( .A1(n5166), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5735) );
  NAND2_X1 U7347 ( .A1(n7019), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5734) );
  OAI211_X1 U7348 ( .C1(n10327), .C2(n5736), .A(n5735), .B(n5734), .ZN(n5737)
         );
  INV_X1 U7349 ( .A(n5737), .ZN(n5738) );
  NOR2_X1 U7350 ( .A1(n8964), .A2(n8568), .ZN(n5740) );
  NAND2_X1 U7351 ( .A1(n8459), .A2(n5740), .ZN(n5741) );
  OAI21_X1 U7352 ( .B1(n8459), .B2(n5740), .A(n5741), .ZN(n8550) );
  NAND2_X1 U7353 ( .A1(n6332), .A2(n5758), .ZN(n5742) );
  INV_X1 U7354 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n5743) );
  INV_X1 U7355 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8415) );
  MUX2_X1 U7356 ( .A(n5743), .B(n8415), .S(n6463), .Z(n5763) );
  XNOR2_X1 U7357 ( .A(n5763), .B(SI_27_), .ZN(n5759) );
  NAND2_X1 U7358 ( .A1(n8336), .A2(n8398), .ZN(n5746) );
  NAND2_X1 U7359 ( .A1(n4408), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n5745) );
  XNOR2_X1 U7360 ( .A(n9172), .B(n5747), .ZN(n5752) );
  XNOR2_X1 U7361 ( .A(n5772), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8959) );
  INV_X1 U7362 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n5750) );
  NAND2_X1 U7363 ( .A1(n7019), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5749) );
  NAND2_X1 U7364 ( .A1(n7047), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5748) );
  OAI211_X1 U7365 ( .C1(n5750), .C2(n7052), .A(n5749), .B(n5748), .ZN(n5751)
         );
  NOR2_X1 U7366 ( .A1(n8735), .A2(n8568), .ZN(n5753) );
  NAND2_X1 U7367 ( .A1(n5752), .A2(n5753), .ZN(n5757) );
  INV_X1 U7368 ( .A(n5752), .ZN(n5755) );
  INV_X1 U7369 ( .A(n5753), .ZN(n5754) );
  NAND2_X1 U7370 ( .A1(n5755), .A2(n5754), .ZN(n5756) );
  AND2_X1 U7371 ( .A1(n5757), .A2(n5756), .ZN(n8458) );
  INV_X1 U7372 ( .A(n5823), .ZN(n5817) );
  NAND2_X1 U7373 ( .A1(n6332), .A2(n6330), .ZN(n5765) );
  INV_X1 U7374 ( .A(n5759), .ZN(n5761) );
  INV_X1 U7375 ( .A(SI_27_), .ZN(n5762) );
  NAND2_X1 U7376 ( .A1(n5763), .A2(n5762), .ZN(n6335) );
  AND2_X1 U7377 ( .A1(n6336), .A2(n6335), .ZN(n5764) );
  NAND2_X1 U7378 ( .A1(n5765), .A2(n5764), .ZN(n5767) );
  INV_X1 U7379 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n5766) );
  INV_X1 U7380 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9924) );
  MUX2_X1 U7381 ( .A(n5766), .B(n9924), .S(n6344), .Z(n6327) );
  XNOR2_X1 U7382 ( .A(n6327), .B(SI_28_), .ZN(n6328) );
  NAND2_X1 U7383 ( .A1(n6223), .A2(n8398), .ZN(n5769) );
  NAND2_X1 U7384 ( .A1(n5251), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n5768) );
  INV_X1 U7385 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5771) );
  INV_X1 U7386 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5770) );
  OAI21_X1 U7387 ( .B1(n5772), .B2(n5771), .A(n5770), .ZN(n5773) );
  AND2_X2 U7388 ( .A1(n5773), .A2(n8451), .ZN(n8949) );
  NAND2_X1 U7389 ( .A1(n8949), .A2(n5834), .ZN(n5779) );
  INV_X1 U7390 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U7391 ( .A1(n7047), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5775) );
  NAND2_X1 U7392 ( .A1(n7019), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5774) );
  OAI211_X1 U7393 ( .C1(n7052), .C2(n5776), .A(n5775), .B(n5774), .ZN(n5777)
         );
  INV_X1 U7394 ( .A(n5777), .ZN(n5778) );
  AND2_X2 U7395 ( .A1(n5779), .A2(n5778), .ZN(n8965) );
  NOR2_X1 U7396 ( .A1(n8965), .A2(n8568), .ZN(n5781) );
  XNOR2_X1 U7397 ( .A(n5781), .B(n5780), .ZN(n5821) );
  NOR4_X1 U7398 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_7__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5785) );
  NOR4_X1 U7399 ( .A1(P2_D_REG_8__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_2__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n5784) );
  NOR4_X1 U7400 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_18__SCAN_IN), .A3(
        P2_D_REG_19__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n5783) );
  NOR4_X1 U7401 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n5782) );
  AND4_X1 U7402 ( .A1(n5785), .A2(n5784), .A3(n5783), .A4(n5782), .ZN(n5800)
         );
  INV_X1 U7403 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10181) );
  INV_X1 U7404 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n10180) );
  INV_X1 U7405 ( .A(P2_D_REG_21__SCAN_IN), .ZN(n10339) );
  INV_X1 U7406 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10347) );
  NAND4_X1 U7407 ( .A1(n10181), .A2(n10180), .A3(n10339), .A4(n10347), .ZN(
        n5788) );
  NOR4_X1 U7408 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_29__SCAN_IN), .A3(
        P2_D_REG_31__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n5786) );
  INV_X1 U7409 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10476) );
  NAND2_X1 U7410 ( .A1(n5786), .A2(n10476), .ZN(n10406) );
  INV_X1 U7411 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10182) );
  INV_X1 U7412 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n10184) );
  INV_X1 U7413 ( .A(P2_D_REG_20__SCAN_IN), .ZN(n10187) );
  INV_X1 U7414 ( .A(P2_D_REG_22__SCAN_IN), .ZN(n10186) );
  NAND4_X1 U7415 ( .A1(n10182), .A2(n10184), .A3(n10187), .A4(n10186), .ZN(
        n5787) );
  NOR4_X1 U7416 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n5788), .A3(n10406), .A4(
        n5787), .ZN(n5799) );
  OR2_X1 U7417 ( .A1(n5789), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n5790) );
  NAND2_X1 U7418 ( .A1(n5790), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5791) );
  XNOR2_X1 U7419 ( .A(n5791), .B(P2_IR_REG_26__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U7420 ( .A1(n5789), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5792) );
  XNOR2_X1 U7421 ( .A(n5792), .B(P2_IR_REG_25__SCAN_IN), .ZN(n8268) );
  INV_X1 U7422 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5793) );
  NAND2_X1 U7423 ( .A1(n5794), .A2(n5793), .ZN(n5795) );
  XNOR2_X1 U7424 ( .A(n8152), .B(P2_B_REG_SCAN_IN), .ZN(n5797) );
  AOI21_X1 U7425 ( .B1(n5800), .B2(n5799), .A(n10179), .ZN(n7256) );
  OR2_X1 U7426 ( .A1(n8152), .A2(n8331), .ZN(n10201) );
  OR2_X1 U7427 ( .A1(n8331), .A2(n8268), .ZN(n10204) );
  NAND2_X1 U7428 ( .A1(n5802), .A2(n10204), .ZN(n7590) );
  OR2_X1 U7429 ( .A1(n7592), .A2(n7590), .ZN(n5803) );
  OR2_X1 U7430 ( .A1(n7256), .A2(n5803), .ZN(n5841) );
  AND2_X1 U7431 ( .A1(n8331), .A2(n8268), .ZN(n5804) );
  NAND2_X1 U7432 ( .A1(n8152), .A2(n5804), .ZN(n6637) );
  OR2_X1 U7433 ( .A1(n5806), .A2(n5805), .ZN(n5807) );
  NAND2_X1 U7434 ( .A1(n5808), .A2(n5807), .ZN(n6636) );
  AND2_X1 U7435 ( .A1(n6636), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5809) );
  INV_X1 U7436 ( .A(n10178), .ZN(n5810) );
  NOR2_X1 U7437 ( .A1(n8595), .A2(n7550), .ZN(n7603) );
  NAND2_X1 U7438 ( .A1(n5838), .A2(n7603), .ZN(n5813) );
  NAND2_X1 U7439 ( .A1(n10249), .A2(n8600), .ZN(n7257) );
  INV_X1 U7440 ( .A(n7257), .ZN(n5812) );
  NOR3_X1 U7441 ( .A1(n4855), .A2(n5821), .A3(n8545), .ZN(n5814) );
  AOI21_X1 U7442 ( .B1(n4855), .B2(n5821), .A(n5814), .ZN(n5815) );
  INV_X1 U7443 ( .A(n5815), .ZN(n5816) );
  NAND2_X1 U7444 ( .A1(n5817), .A2(n5816), .ZN(n5826) );
  INV_X1 U7445 ( .A(n8761), .ZN(n5818) );
  NAND2_X1 U7446 ( .A1(n8765), .A2(n8608), .ZN(n7269) );
  INV_X1 U7447 ( .A(n7269), .ZN(n6696) );
  NOR2_X1 U7448 ( .A1(n9246), .A2(n6696), .ZN(n5819) );
  OAI21_X1 U7449 ( .B1(n4855), .B2(n8558), .A(n8549), .ZN(n5825) );
  NAND3_X1 U7450 ( .A1(n9168), .A2(n8558), .A3(n5821), .ZN(n5820) );
  OAI21_X1 U7451 ( .B1(n9168), .B2(n5821), .A(n5820), .ZN(n5822) );
  NAND2_X1 U7452 ( .A1(n5823), .A2(n5822), .ZN(n5824) );
  NAND3_X1 U7453 ( .A1(n5826), .A2(n5825), .A3(n5824), .ZN(n5848) );
  NAND2_X1 U7454 ( .A1(n5828), .A2(n5827), .ZN(n6642) );
  NAND2_X1 U7455 ( .A1(n6642), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5830) );
  XNOR2_X1 U7456 ( .A(n5830), .B(n5829), .ZN(n6704) );
  OR2_X1 U7457 ( .A1(n8735), .A2(n9100), .ZN(n5837) );
  INV_X1 U7458 ( .A(n8451), .ZN(n5835) );
  INV_X1 U7459 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8452) );
  NAND2_X1 U7460 ( .A1(n7019), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5832) );
  NAND2_X1 U7461 ( .A1(n7047), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5831) );
  OAI211_X1 U7462 ( .C1(n8452), .C2(n7052), .A(n5832), .B(n5831), .ZN(n5833)
         );
  AOI21_X1 U7463 ( .B1(n5835), .B2(n5834), .A(n5833), .ZN(n8434) );
  OR2_X1 U7464 ( .A1(n8434), .A2(n9102), .ZN(n5836) );
  NAND2_X1 U7465 ( .A1(n5837), .A2(n5836), .ZN(n8942) );
  INV_X1 U7466 ( .A(n8942), .ZN(n5845) );
  NAND2_X1 U7467 ( .A1(n5838), .A2(n8761), .ZN(n7403) );
  NAND2_X1 U7468 ( .A1(n10178), .A2(n7603), .ZN(n5839) );
  OAI21_X1 U7469 ( .B1(n9246), .B2(P2_U3152), .A(n5839), .ZN(n5840) );
  NAND2_X1 U7470 ( .A1(n5841), .A2(n5840), .ZN(n5843) );
  OAI211_X1 U7471 ( .C1(n8761), .C2(n7269), .A(n6637), .B(n6636), .ZN(n7254)
         );
  NAND2_X1 U7472 ( .A1(n7254), .A2(P2_STATE_REG_SCAN_IN), .ZN(n5842) );
  AOI22_X1 U7473 ( .A1(n8949), .A2(n8517), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n5844) );
  OAI21_X1 U7474 ( .B1(n5845), .B2(n7403), .A(n5844), .ZN(n5846) );
  NAND2_X1 U7475 ( .A1(n5848), .A2(n5847), .ZN(P2_U3222) );
  NAND4_X1 U7476 ( .A1(n5852), .A2(n5851), .A3(n5850), .A4(n5849), .ZN(n5855)
         );
  INV_X2 U7477 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10426) );
  NOR2_X1 U7478 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5859) );
  NOR2_X1 U7479 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n5858) );
  NOR2_X1 U7480 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n5857) );
  NAND4_X1 U7481 ( .A1(n5859), .A2(n5858), .A3(n5857), .A4(n5856), .ZN(n5861)
         );
  NAND4_X1 U7482 ( .A1(n6289), .A2(n10487), .A3(n6044), .A4(n6293), .ZN(n5860)
         );
  NOR2_X1 U7483 ( .A1(n5861), .A2(n5860), .ZN(n5862) );
  NOR3_X1 U7484 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .A3(
        P1_IR_REG_26__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U7485 ( .A1(n6106), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5876) );
  AND2_X4 U7486 ( .A1(n5872), .A2(n5870), .ZN(n6205) );
  INV_X1 U7487 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5871) );
  XNOR2_X1 U7488 ( .A(n5871), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n9363) );
  NAND2_X1 U7489 ( .A1(n6205), .A2(n9363), .ZN(n5875) );
  AND2_X4 U7490 ( .A1(n5872), .A2(n8413), .ZN(n6348) );
  NAND2_X1 U7491 ( .A1(n6348), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5874) );
  OAI21_X1 U7492 ( .B1(P1_IR_REG_25__SCAN_IN), .B2(P1_IR_REG_26__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5877) );
  NAND2_X1 U7493 ( .A1(n6989), .A2(n6469), .ZN(n5886) );
  OR2_X1 U7494 ( .A1(n6467), .A2(n6990), .ZN(n5885) );
  INV_X1 U7495 ( .A(n5905), .ZN(n5881) );
  NOR2_X1 U7496 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n5880) );
  NAND2_X1 U7497 ( .A1(n5881), .A2(n5880), .ZN(n5988) );
  NAND2_X1 U7498 ( .A1(n5988), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5882) );
  MUX2_X1 U7499 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5882), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5883) );
  NAND2_X1 U7500 ( .A1(n5883), .A2(n5947), .ZN(n7172) );
  OR2_X1 U7501 ( .A1(n5946), .A2(n7172), .ZN(n5884) );
  NAND3_X1 U7502 ( .A1(n5886), .A2(n5885), .A3(n5884), .ZN(n7724) );
  NAND2_X1 U7503 ( .A1(n9444), .A2(n9364), .ZN(n6579) );
  NAND2_X1 U7504 ( .A1(n6106), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5890) );
  INV_X1 U7505 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5887) );
  NAND2_X1 U7506 ( .A1(n6205), .A2(n5887), .ZN(n5889) );
  NAND2_X1 U7507 ( .A1(n6348), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5888) );
  INV_X1 U7508 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n10392) );
  INV_X1 U7509 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5891) );
  INV_X1 U7510 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n7011) );
  OR2_X1 U7511 ( .A1(n6467), .A2(n7011), .ZN(n5893) );
  OR2_X1 U7512 ( .A1(n5935), .A2(n7012), .ZN(n5892) );
  OAI211_X1 U7513 ( .C1(n5946), .C2(n7143), .A(n5893), .B(n5892), .ZN(n5926)
         );
  NOR2_X1 U7514 ( .A1(n10082), .A2(n5926), .ZN(n7714) );
  NOR2_X1 U7515 ( .A1(n9444), .A2(n7724), .ZN(n5894) );
  NAND2_X1 U7516 ( .A1(n6348), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5898) );
  NAND2_X1 U7517 ( .A1(n5912), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5897) );
  NAND2_X1 U7518 ( .A1(n6205), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5896) );
  NAND2_X1 U7519 ( .A1(n5913), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5895) );
  NAND2_X1 U7520 ( .A1(n6998), .A2(SI_0_), .ZN(n5899) );
  XNOR2_X1 U7521 ( .A(n5899), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n9926) );
  MUX2_X1 U7522 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9926), .S(n5946), .Z(n7666) );
  NAND2_X1 U7523 ( .A1(n7034), .A2(n7666), .ZN(n10054) );
  NAND2_X1 U7524 ( .A1(n6348), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5903) );
  NAND2_X1 U7525 ( .A1(n5912), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5902) );
  NAND2_X1 U7526 ( .A1(n6205), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5900) );
  OR2_X1 U7527 ( .A1(n8365), .A2(n5935), .ZN(n5909) );
  NAND2_X1 U7528 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5904) );
  MUX2_X1 U7529 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5904), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n5906) );
  NAND2_X1 U7530 ( .A1(n5906), .A2(n5905), .ZN(n8364) );
  NOR2_X1 U7531 ( .A1(n5946), .A2(n8364), .ZN(n5907) );
  OAI21_X1 U7532 ( .B1(n10054), .B2(n7765), .A(n10078), .ZN(n5911) );
  NAND2_X1 U7533 ( .A1(n10054), .A2(n7765), .ZN(n5910) );
  NAND2_X1 U7534 ( .A1(n5911), .A2(n5910), .ZN(n7764) );
  NAND2_X1 U7535 ( .A1(n6205), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5916) );
  NAND2_X1 U7536 ( .A1(n5912), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5915) );
  NAND2_X1 U7537 ( .A1(n5913), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5914) );
  NAND2_X2 U7538 ( .A1(n5918), .A2(n5917), .ZN(n6711) );
  INV_X1 U7539 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6988) );
  OR2_X1 U7540 ( .A1(n6467), .A2(n6988), .ZN(n5923) );
  OR2_X1 U7541 ( .A1(n5946), .A2(n7057), .ZN(n5922) );
  OR2_X1 U7542 ( .A1(n7000), .A2(n5935), .ZN(n5921) );
  NAND3_X2 U7543 ( .A1(n5923), .A2(n5922), .A3(n5921), .ZN(n6715) );
  INV_X2 U7544 ( .A(n6715), .ZN(n7768) );
  NAND2_X1 U7545 ( .A1(n7764), .A2(n6564), .ZN(n5925) );
  INV_X1 U7546 ( .A(n6711), .ZN(n7981) );
  NAND2_X1 U7547 ( .A1(n7981), .A2(n7768), .ZN(n5924) );
  NAND2_X1 U7548 ( .A1(n7721), .A2(n5926), .ZN(n6578) );
  NAND2_X1 U7549 ( .A1(n6353), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5933) );
  INV_X1 U7550 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U7551 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5927) );
  NAND2_X1 U7552 ( .A1(n5928), .A2(n5927), .ZN(n5929) );
  AND2_X1 U7553 ( .A1(n5954), .A2(n5929), .ZN(n10032) );
  NAND2_X1 U7554 ( .A1(n6205), .A2(n10032), .ZN(n5932) );
  NAND2_X1 U7555 ( .A1(n5913), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n5931) );
  NAND2_X1 U7556 ( .A1(n6348), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5930) );
  INV_X1 U7557 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6991) );
  NAND2_X1 U7558 ( .A1(n5947), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5934) );
  XNOR2_X1 U7559 ( .A(n5934), .B(n5948), .ZN(n9446) );
  OAI22_X1 U7560 ( .A1(n6467), .A2(n6991), .B1(n5946), .B2(n9446), .ZN(n5937)
         );
  NOR2_X1 U7561 ( .A1(n7009), .A2(n5935), .ZN(n5936) );
  NAND2_X1 U7562 ( .A1(n7542), .A2(n10031), .ZN(n6363) );
  INV_X1 U7563 ( .A(n7542), .ZN(n9443) );
  NAND2_X1 U7564 ( .A1(n9443), .A2(n5032), .ZN(n6580) );
  NAND2_X1 U7565 ( .A1(n9443), .A2(n10031), .ZN(n5938) );
  NAND2_X1 U7566 ( .A1(n6106), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n5945) );
  INV_X1 U7567 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U7568 ( .A1(n5956), .A2(n5940), .ZN(n5941) );
  AND2_X1 U7569 ( .A1(n5969), .A2(n5941), .ZN(n7469) );
  NAND2_X1 U7570 ( .A1(n6205), .A2(n7469), .ZN(n5944) );
  NAND2_X1 U7571 ( .A1(n5913), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U7572 ( .A1(n6348), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5942) );
  NAND2_X1 U7573 ( .A1(n7015), .A2(n6469), .ZN(n5952) );
  INV_X2 U7574 ( .A(n5946), .ZN(n6957) );
  INV_X1 U7575 ( .A(n5947), .ZN(n5949) );
  NAND2_X1 U7576 ( .A1(n5949), .A2(n5948), .ZN(n5961) );
  NAND2_X1 U7577 ( .A1(n5964), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5950) );
  XNOR2_X1 U7578 ( .A(n5950), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7112) );
  AOI22_X1 U7579 ( .A1(n6114), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6957), .B2(
        n7112), .ZN(n5951) );
  OR2_X1 U7580 ( .A1(n6754), .A2(n10162), .ZN(n6373) );
  NAND2_X1 U7581 ( .A1(n10162), .A2(n6754), .ZN(n8018) );
  NAND2_X1 U7582 ( .A1(n6353), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5960) );
  INV_X1 U7583 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U7584 ( .A1(n5954), .A2(n5953), .ZN(n5955) );
  AND2_X1 U7585 ( .A1(n5956), .A2(n5955), .ZN(n7630) );
  NAND2_X1 U7586 ( .A1(n6205), .A2(n7630), .ZN(n5959) );
  NAND2_X1 U7587 ( .A1(n5913), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n5958) );
  NAND2_X1 U7588 ( .A1(n6348), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5957) );
  AND4_X2 U7589 ( .A1(n5960), .A2(n5959), .A3(n5958), .A4(n5957), .ZN(n10043)
         );
  INV_X1 U7590 ( .A(n10043), .ZN(n10160) );
  NAND2_X1 U7591 ( .A1(n5961), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5962) );
  XNOR2_X1 U7592 ( .A(n5962), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7109) );
  NOR2_X1 U7593 ( .A1(n10160), .A2(n7625), .ZN(n7994) );
  INV_X1 U7594 ( .A(n6754), .ZN(n9442) );
  NOR2_X1 U7595 ( .A1(n10162), .A2(n9442), .ZN(n5963) );
  NAND2_X1 U7596 ( .A1(n7028), .A2(n6469), .ZN(n5967) );
  OAI21_X1 U7597 ( .B1(n5964), .B2(P1_IR_REG_7__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5965) );
  XNOR2_X1 U7598 ( .A(n5965), .B(P1_IR_REG_8__SCAN_IN), .ZN(n7190) );
  AOI22_X1 U7599 ( .A1(n6114), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6957), .B2(
        n7190), .ZN(n5966) );
  NAND2_X1 U7600 ( .A1(n6353), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5974) );
  INV_X1 U7601 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5968) );
  NAND2_X1 U7602 ( .A1(n5969), .A2(n5968), .ZN(n5970) );
  AND2_X1 U7603 ( .A1(n5981), .A2(n5970), .ZN(n8034) );
  NAND2_X1 U7604 ( .A1(n6205), .A2(n8034), .ZN(n5973) );
  NAND2_X1 U7605 ( .A1(n5913), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7606 ( .A1(n6348), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5971) );
  NAND2_X1 U7607 ( .A1(n5975), .A2(n10139), .ZN(n6376) );
  NAND3_X1 U7608 ( .A1(n7618), .A2(n8029), .A3(n8032), .ZN(n5979) );
  NAND2_X1 U7609 ( .A1(n10043), .A2(n7625), .ZN(n6525) );
  NAND2_X1 U7610 ( .A1(n6525), .A2(n6364), .ZN(n6560) );
  NAND2_X1 U7611 ( .A1(n7920), .A2(n6560), .ZN(n8028) );
  NAND3_X1 U7612 ( .A1(n8032), .A2(n8029), .A3(n8028), .ZN(n5977) );
  INV_X1 U7613 ( .A(n10139), .ZN(n10158) );
  NAND2_X1 U7614 ( .A1(n5975), .A2(n10158), .ZN(n5976) );
  AND2_X1 U7615 ( .A1(n5977), .A2(n5976), .ZN(n5978) );
  NAND2_X1 U7616 ( .A1(n5979), .A2(n5978), .ZN(n7919) );
  NAND2_X1 U7617 ( .A1(n6353), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n5986) );
  NAND2_X1 U7618 ( .A1(n5981), .A2(n5980), .ZN(n5982) );
  AND2_X1 U7619 ( .A1(n6000), .A2(n5982), .ZN(n7929) );
  NAND2_X1 U7620 ( .A1(n6205), .A2(n7929), .ZN(n5985) );
  NAND2_X1 U7621 ( .A1(n5913), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5984) );
  NAND2_X1 U7622 ( .A1(n6348), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5983) );
  INV_X1 U7623 ( .A(n9730), .ZN(n9959) );
  NAND2_X1 U7624 ( .A1(n6994), .A2(n6469), .ZN(n5992) );
  INV_X1 U7625 ( .A(n5987), .ZN(n5990) );
  INV_X1 U7626 ( .A(n5988), .ZN(n5989) );
  NAND2_X1 U7627 ( .A1(n5990), .A2(n5989), .ZN(n5995) );
  NAND2_X1 U7628 ( .A1(n5995), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5991) );
  XNOR2_X1 U7629 ( .A(n5991), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7221) );
  OR2_X1 U7630 ( .A1(n9959), .A2(n10144), .ZN(n5993) );
  NAND2_X1 U7631 ( .A1(n10144), .A2(n9959), .ZN(n5994) );
  NAND2_X1 U7632 ( .A1(n7013), .A2(n6469), .ZN(n5998) );
  NAND2_X1 U7633 ( .A1(n6006), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5996) );
  XNOR2_X1 U7634 ( .A(n5996), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9469) );
  AOI22_X1 U7635 ( .A1(n6114), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6957), .B2(
        n9469), .ZN(n5997) );
  NAND2_X1 U7636 ( .A1(n5998), .A2(n5997), .ZN(n6782) );
  NAND2_X1 U7637 ( .A1(n6000), .A2(n5999), .ZN(n6001) );
  AND2_X1 U7638 ( .A1(n6013), .A2(n6001), .ZN(n9727) );
  NAND2_X1 U7639 ( .A1(n6205), .A2(n9727), .ZN(n6005) );
  NAND2_X1 U7640 ( .A1(n6106), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U7641 ( .A1(n6348), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U7642 ( .A1(n5913), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n6002) );
  NAND2_X1 U7643 ( .A1(n6782), .A2(n10140), .ZN(n6379) );
  INV_X1 U7644 ( .A(n10140), .ZN(n9441) );
  NAND2_X1 U7645 ( .A1(n7026), .A2(n6469), .ZN(n6011) );
  INV_X1 U7646 ( .A(n6006), .ZN(n6008) );
  INV_X1 U7647 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6007) );
  NAND2_X1 U7648 ( .A1(n6008), .A2(n6007), .ZN(n6020) );
  NAND2_X1 U7649 ( .A1(n6020), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6009) );
  XNOR2_X1 U7650 ( .A(n6009), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7234) );
  AOI22_X1 U7651 ( .A1(n6114), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6957), .B2(
        n7234), .ZN(n6010) );
  NAND2_X1 U7652 ( .A1(n6353), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6018) );
  INV_X1 U7653 ( .A(n6024), .ZN(n6025) );
  NAND2_X1 U7654 ( .A1(n6013), .A2(n10553), .ZN(n6014) );
  AND2_X1 U7655 ( .A1(n6025), .A2(n6014), .ZN(n8061) );
  NAND2_X1 U7656 ( .A1(n6205), .A2(n8061), .ZN(n6017) );
  NAND2_X1 U7657 ( .A1(n6349), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n6016) );
  NAND2_X1 U7658 ( .A1(n6348), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6015) );
  INV_X1 U7659 ( .A(n9876), .ZN(n9960) );
  NAND2_X1 U7660 ( .A1(n9888), .A2(n9960), .ZN(n6019) );
  NAND2_X1 U7661 ( .A1(n7042), .A2(n6469), .ZN(n6023) );
  OAI21_X1 U7662 ( .B1(n6020), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6021) );
  XNOR2_X1 U7663 ( .A(n6021), .B(P1_IR_REG_12__SCAN_IN), .ZN(n7451) );
  AOI22_X1 U7664 ( .A1(n6114), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n6957), .B2(
        n7451), .ZN(n6022) );
  NAND2_X1 U7665 ( .A1(n6353), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n6030) );
  INV_X1 U7666 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7297) );
  NAND2_X1 U7667 ( .A1(n6025), .A2(n7297), .ZN(n6026) );
  AND2_X1 U7668 ( .A1(n6036), .A2(n6026), .ZN(n8251) );
  NAND2_X1 U7669 ( .A1(n6205), .A2(n8251), .ZN(n6029) );
  NAND2_X1 U7670 ( .A1(n6348), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7671 ( .A1(n5913), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6027) );
  OR2_X1 U7672 ( .A1(n9880), .A2(n9884), .ZN(n6368) );
  NAND2_X1 U7673 ( .A1(n9880), .A2(n9884), .ZN(n6380) );
  AND2_X1 U7674 ( .A1(n6368), .A2(n6380), .ZN(n8042) );
  NAND2_X1 U7675 ( .A1(n8051), .A2(n6031), .ZN(n8050) );
  INV_X1 U7676 ( .A(n9884), .ZN(n9440) );
  NAND2_X1 U7677 ( .A1(n9880), .A2(n9440), .ZN(n6032) );
  NAND2_X1 U7678 ( .A1(n8050), .A2(n6032), .ZN(n8182) );
  INV_X1 U7679 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6046) );
  OR2_X1 U7680 ( .A1(n6045), .A2(n6046), .ZN(n6033) );
  XNOR2_X1 U7681 ( .A(n6033), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7454) );
  AOI22_X1 U7682 ( .A1(n6114), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n6957), .B2(
        n7454), .ZN(n6034) );
  NAND2_X1 U7683 ( .A1(n6106), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n6041) );
  NAND2_X1 U7684 ( .A1(n6036), .A2(n6035), .ZN(n6037) );
  AND2_X1 U7685 ( .A1(n6054), .A2(n6037), .ZN(n8243) );
  NAND2_X1 U7686 ( .A1(n6205), .A2(n8243), .ZN(n6040) );
  NAND2_X1 U7687 ( .A1(n6349), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6039) );
  NAND2_X1 U7688 ( .A1(n6348), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6038) );
  OR2_X1 U7689 ( .A1(n9872), .A2(n9439), .ZN(n6042) );
  NAND2_X1 U7690 ( .A1(n9872), .A2(n9439), .ZN(n6043) );
  NAND2_X1 U7691 ( .A1(n7083), .A2(n6469), .ZN(n6052) );
  NOR2_X1 U7692 ( .A1(n6073), .A2(n6046), .ZN(n6047) );
  NAND2_X1 U7693 ( .A1(n6047), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6050) );
  INV_X1 U7694 ( .A(n6047), .ZN(n6049) );
  INV_X1 U7695 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U7696 ( .A1(n6049), .A2(n6048), .ZN(n6061) );
  AOI22_X1 U7697 ( .A1(n6114), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6957), .B2(
        n7829), .ZN(n6051) );
  NAND2_X1 U7698 ( .A1(n6353), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n6059) );
  INV_X1 U7699 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7700 ( .A1(n6054), .A2(n6053), .ZN(n6055) );
  AND2_X1 U7701 ( .A1(n6066), .A2(n6055), .ZN(n9295) );
  NAND2_X1 U7702 ( .A1(n6205), .A2(n9295), .ZN(n6058) );
  NAND2_X1 U7703 ( .A1(n5913), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7704 ( .A1(n6348), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6056) );
  INV_X1 U7705 ( .A(n9868), .ZN(n9438) );
  AND2_X1 U7706 ( .A1(n9864), .A2(n9438), .ZN(n6060) );
  NAND2_X1 U7707 ( .A1(n7144), .A2(n6469), .ZN(n6064) );
  NAND2_X1 U7708 ( .A1(n6061), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6062) );
  XNOR2_X1 U7709 ( .A(n6062), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9488) );
  AOI22_X1 U7710 ( .A1(n6114), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6957), .B2(
        n9488), .ZN(n6063) );
  INV_X1 U7711 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6065) );
  NAND2_X1 U7712 ( .A1(n6066), .A2(n6065), .ZN(n6067) );
  NAND2_X1 U7713 ( .A1(n6078), .A2(n6067), .ZN(n9710) );
  NAND2_X1 U7714 ( .A1(n6353), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n6069) );
  NAND2_X1 U7715 ( .A1(n6349), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6068) );
  AND2_X1 U7716 ( .A1(n6069), .A2(n6068), .ZN(n6071) );
  NAND2_X1 U7717 ( .A1(n6348), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n6070) );
  OAI211_X1 U7718 ( .C1(n9710), .C2(n6217), .A(n6071), .B(n6070), .ZN(n9696)
         );
  OR2_X1 U7719 ( .A1(n9856), .A2(n9696), .ZN(n6259) );
  NAND2_X1 U7720 ( .A1(n9856), .A2(n9696), .ZN(n6403) );
  NAND2_X1 U7721 ( .A1(n7237), .A2(n6469), .ZN(n6076) );
  NAND2_X1 U7722 ( .A1(n6085), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6074) );
  XNOR2_X1 U7723 ( .A(n6074), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9987) );
  AOI22_X1 U7724 ( .A1(n6114), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6957), .B2(
        n9987), .ZN(n6075) );
  INV_X1 U7725 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n10445) );
  NAND2_X1 U7726 ( .A1(n6078), .A2(n10445), .ZN(n6079) );
  NAND2_X1 U7727 ( .A1(n6093), .A2(n6079), .ZN(n9686) );
  OR2_X1 U7728 ( .A1(n9686), .A2(n6217), .ZN(n6082) );
  AOI22_X1 U7729 ( .A1(n6353), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n6348), .B2(
        P1_REG2_REG_16__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U7730 ( .A1(n6349), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n6080) );
  OR2_X1 U7731 ( .A1(n9689), .A2(n9843), .ZN(n6512) );
  NAND2_X1 U7732 ( .A1(n9689), .A2(n9843), .ZN(n6515) );
  NAND2_X1 U7733 ( .A1(n9684), .A2(n4577), .ZN(n6084) );
  INV_X1 U7734 ( .A(n9843), .ZN(n9676) );
  NAND2_X1 U7735 ( .A1(n9689), .A2(n9676), .ZN(n6083) );
  NAND2_X1 U7736 ( .A1(n6084), .A2(n6083), .ZN(n9669) );
  NAND2_X1 U7737 ( .A1(n7249), .A2(n6469), .ZN(n6090) );
  NAND2_X1 U7738 ( .A1(n4467), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6087) );
  INV_X1 U7739 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6086) );
  OR2_X1 U7740 ( .A1(n6087), .A2(n6086), .ZN(n6088) );
  NAND2_X1 U7741 ( .A1(n6087), .A2(n6086), .ZN(n6099) );
  AOI22_X1 U7742 ( .A1(n6114), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6957), .B2(
        n10000), .ZN(n6089) );
  INV_X1 U7743 ( .A(n6103), .ZN(n6104) );
  INV_X1 U7744 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6092) );
  NAND2_X1 U7745 ( .A1(n6093), .A2(n6092), .ZN(n6094) );
  AND2_X1 U7746 ( .A1(n6104), .A2(n6094), .ZN(n9675) );
  NAND2_X1 U7747 ( .A1(n9675), .A2(n6205), .ZN(n6097) );
  AOI22_X1 U7748 ( .A1(n6353), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n6349), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n6096) );
  NAND2_X1 U7749 ( .A1(n6348), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n6095) );
  AND2_X1 U7750 ( .A1(n9847), .A2(n9695), .ZN(n6098) );
  NAND2_X1 U7751 ( .A1(n7416), .A2(n6469), .ZN(n6102) );
  NAND2_X1 U7752 ( .A1(n6099), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6100) );
  XNOR2_X1 U7753 ( .A(n6100), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9495) );
  AOI22_X1 U7754 ( .A1(n6114), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n9495), .B2(
        n6957), .ZN(n6101) );
  NAND2_X1 U7755 ( .A1(n6104), .A2(n4655), .ZN(n6105) );
  NAND2_X1 U7756 ( .A1(n6118), .A2(n6105), .ZN(n9651) );
  OR2_X1 U7757 ( .A1(n9651), .A2(n6217), .ZN(n6111) );
  INV_X1 U7758 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9484) );
  NAND2_X1 U7759 ( .A1(n6349), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7760 ( .A1(n6348), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n6107) );
  OAI211_X1 U7761 ( .C1(n6012), .C2(n9484), .A(n6108), .B(n6107), .ZN(n6109)
         );
  INV_X1 U7762 ( .A(n6109), .ZN(n6110) );
  OR2_X1 U7763 ( .A1(n9662), .A2(n9844), .ZN(n6407) );
  NAND2_X1 U7764 ( .A1(n9662), .A2(n9844), .ZN(n6416) );
  INV_X1 U7765 ( .A(n9844), .ZN(n9437) );
  NAND2_X1 U7766 ( .A1(n7429), .A2(n6469), .ZN(n6116) );
  NAND2_X1 U7767 ( .A1(n6238), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6113) );
  INV_X1 U7768 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6112) );
  AOI22_X1 U7769 ( .A1(n6114), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10052), 
        .B2(n6957), .ZN(n6115) );
  INV_X1 U7770 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7771 ( .A1(n6118), .A2(n6117), .ZN(n6119) );
  AND2_X1 U7772 ( .A1(n6130), .A2(n6119), .ZN(n9640) );
  NAND2_X1 U7773 ( .A1(n9640), .A2(n6205), .ZN(n6124) );
  INV_X1 U7774 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9485) );
  NAND2_X1 U7775 ( .A1(n6349), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7776 ( .A1(n6348), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6120) );
  OAI211_X1 U7777 ( .C1(n6012), .C2(n9485), .A(n6121), .B(n6120), .ZN(n6122)
         );
  INV_X1 U7778 ( .A(n6122), .ZN(n6123) );
  OR2_X1 U7779 ( .A1(n6853), .A2(n9436), .ZN(n6125) );
  NAND2_X1 U7780 ( .A1(n9634), .A2(n6125), .ZN(n6127) );
  NAND2_X1 U7781 ( .A1(n6853), .A2(n9436), .ZN(n6126) );
  NAND2_X1 U7782 ( .A1(n7532), .A2(n6469), .ZN(n6129) );
  OR2_X1 U7783 ( .A1(n6467), .A2(n7533), .ZN(n6128) );
  NAND2_X1 U7784 ( .A1(n6130), .A2(n4656), .ZN(n6131) );
  NAND2_X1 U7785 ( .A1(n6141), .A2(n6131), .ZN(n9628) );
  OR2_X1 U7786 ( .A1(n9628), .A2(n6217), .ZN(n6136) );
  INV_X1 U7787 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n10295) );
  NAND2_X1 U7788 ( .A1(n6349), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6133) );
  NAND2_X1 U7789 ( .A1(n6348), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6132) );
  OAI211_X1 U7790 ( .C1(n6012), .C2(n10295), .A(n6133), .B(n6132), .ZN(n6134)
         );
  INV_X1 U7791 ( .A(n6134), .ZN(n6135) );
  NAND2_X1 U7792 ( .A1(n6136), .A2(n6135), .ZN(n9614) );
  AND2_X1 U7793 ( .A1(n9823), .A2(n9614), .ZN(n6138) );
  OR2_X1 U7794 ( .A1(n9823), .A2(n9614), .ZN(n6137) );
  NAND2_X1 U7795 ( .A1(n7587), .A2(n6469), .ZN(n6140) );
  OR2_X1 U7796 ( .A1(n6467), .A2(n7700), .ZN(n6139) );
  INV_X1 U7797 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9323) );
  NAND2_X1 U7798 ( .A1(n6141), .A2(n9323), .ZN(n6142) );
  NAND2_X1 U7799 ( .A1(n6150), .A2(n6142), .ZN(n9612) );
  OR2_X1 U7800 ( .A1(n9612), .A2(n6217), .ZN(n6147) );
  INV_X1 U7801 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n9611) );
  NAND2_X1 U7802 ( .A1(n6353), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7803 ( .A1(n6349), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6143) );
  OAI211_X1 U7804 ( .C1(n9611), .C2(n6231), .A(n6144), .B(n6143), .ZN(n6145)
         );
  INV_X1 U7805 ( .A(n6145), .ZN(n6146) );
  NAND2_X1 U7806 ( .A1(n7940), .A2(n6469), .ZN(n6149) );
  OR2_X1 U7807 ( .A1(n6467), .A2(n7979), .ZN(n6148) );
  INV_X1 U7808 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9383) );
  NAND2_X1 U7809 ( .A1(n6150), .A2(n9383), .ZN(n6151) );
  NAND2_X1 U7810 ( .A1(n6172), .A2(n6151), .ZN(n9387) );
  INV_X1 U7811 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7812 ( .A1(n6353), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7813 ( .A1(n6349), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n6152) );
  OAI211_X1 U7814 ( .C1(n6154), .C2(n6231), .A(n6153), .B(n6152), .ZN(n6155)
         );
  INV_X1 U7815 ( .A(n6155), .ZN(n6156) );
  NAND2_X1 U7816 ( .A1(n9807), .A2(n9814), .ZN(n6157) );
  NAND2_X1 U7817 ( .A1(n9600), .A2(n9581), .ZN(n9556) );
  NAND2_X1 U7818 ( .A1(n6158), .A2(n6469), .ZN(n6160) );
  OR2_X1 U7819 ( .A1(n6467), .A2(n10566), .ZN(n6159) );
  NAND2_X2 U7820 ( .A1(n6160), .A2(n6159), .ZN(n9795) );
  INV_X1 U7821 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6162) );
  NAND2_X1 U7822 ( .A1(n6174), .A2(n6162), .ZN(n6163) );
  NAND2_X1 U7823 ( .A1(n6203), .A2(n6163), .ZN(n9570) );
  INV_X1 U7824 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n9572) );
  NAND2_X1 U7825 ( .A1(n6353), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7826 ( .A1(n6349), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n6164) );
  OAI211_X1 U7827 ( .C1(n6231), .C2(n9572), .A(n6165), .B(n6164), .ZN(n6166)
         );
  INV_X1 U7828 ( .A(n6166), .ZN(n6167) );
  OR2_X1 U7829 ( .A1(n9795), .A2(n9782), .ZN(n6193) );
  INV_X1 U7830 ( .A(n6193), .ZN(n6182) );
  NAND2_X1 U7831 ( .A1(n9795), .A2(n9782), .ZN(n6180) );
  NAND2_X1 U7832 ( .A1(n8014), .A2(n6469), .ZN(n6170) );
  OR2_X1 U7833 ( .A1(n6467), .A2(n8017), .ZN(n6169) );
  INV_X1 U7834 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7835 ( .A1(n6172), .A2(n6171), .ZN(n6173) );
  NAND2_X1 U7836 ( .A1(n6174), .A2(n6173), .ZN(n9583) );
  INV_X1 U7837 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n9582) );
  NAND2_X1 U7838 ( .A1(n6353), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6176) );
  NAND2_X1 U7839 ( .A1(n6349), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6175) );
  OAI211_X1 U7840 ( .C1(n9582), .C2(n6231), .A(n6176), .B(n6175), .ZN(n6177)
         );
  INV_X1 U7841 ( .A(n6177), .ZN(n6178) );
  NAND2_X1 U7842 ( .A1(n6260), .A2(n9804), .ZN(n9558) );
  AND2_X1 U7843 ( .A1(n6180), .A2(n9558), .ZN(n6181) );
  AND2_X1 U7844 ( .A1(n9556), .A2(n6192), .ZN(n9537) );
  NAND2_X1 U7845 ( .A1(n8267), .A2(n6469), .ZN(n6184) );
  OR2_X1 U7846 ( .A1(n6467), .A2(n8315), .ZN(n6183) );
  XNOR2_X1 U7847 ( .A(n6203), .B(P1_REG3_REG_25__SCAN_IN), .ZN(n9551) );
  NAND2_X1 U7848 ( .A1(n9551), .A2(n6205), .ZN(n6189) );
  INV_X1 U7849 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n9546) );
  NAND2_X1 U7850 ( .A1(n6353), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n6186) );
  NAND2_X1 U7851 ( .A1(n6349), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6185) );
  OAI211_X1 U7852 ( .C1(n9546), .C2(n6231), .A(n6186), .B(n6185), .ZN(n6187)
         );
  INV_X1 U7853 ( .A(n6187), .ZN(n6188) );
  NAND2_X1 U7854 ( .A1(n9545), .A2(n9792), .ZN(n6440) );
  INV_X1 U7855 ( .A(n9542), .ZN(n6191) );
  AND2_X1 U7856 ( .A1(n9537), .A2(n6191), .ZN(n6190) );
  NAND2_X1 U7857 ( .A1(n9536), .A2(n6190), .ZN(n6199) );
  INV_X1 U7858 ( .A(n6192), .ZN(n6195) );
  OR2_X1 U7859 ( .A1(n6260), .A2(n9804), .ZN(n9557) );
  AND2_X1 U7860 ( .A1(n9557), .A2(n6193), .ZN(n6194) );
  OR2_X1 U7861 ( .A1(n9545), .A2(n9435), .ZN(n6196) );
  NAND2_X1 U7862 ( .A1(n8330), .A2(n6469), .ZN(n6201) );
  OR2_X1 U7863 ( .A1(n6467), .A2(n8333), .ZN(n6200) );
  INV_X1 U7864 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8388) );
  INV_X1 U7865 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6202) );
  OAI21_X1 U7866 ( .B1(n6203), .B2(n8388), .A(n6202), .ZN(n6204) );
  NAND2_X1 U7867 ( .A1(n9411), .A2(n6205), .ZN(n6211) );
  INV_X1 U7868 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n6208) );
  NAND2_X1 U7869 ( .A1(n6353), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7870 ( .A1(n6349), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n6206) );
  OAI211_X1 U7871 ( .C1(n6208), .C2(n6231), .A(n6207), .B(n6206), .ZN(n6209)
         );
  INV_X1 U7872 ( .A(n6209), .ZN(n6210) );
  INV_X1 U7873 ( .A(n9776), .ZN(n9418) );
  NAND2_X1 U7874 ( .A1(n8336), .A2(n6469), .ZN(n6213) );
  OR2_X1 U7875 ( .A1(n6467), .A2(n8415), .ZN(n6212) );
  INV_X1 U7876 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n10569) );
  NAND2_X1 U7877 ( .A1(n6215), .A2(n10569), .ZN(n6216) );
  NAND2_X1 U7878 ( .A1(n6227), .A2(n6216), .ZN(n8348) );
  INV_X1 U7879 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n8347) );
  NAND2_X1 U7880 ( .A1(n6353), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n6219) );
  NAND2_X1 U7881 ( .A1(n6349), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6218) );
  OAI211_X1 U7882 ( .C1(n8347), .C2(n6231), .A(n6219), .B(n6218), .ZN(n6220)
         );
  INV_X1 U7883 ( .A(n6220), .ZN(n6221) );
  NAND2_X1 U7884 ( .A1(n8350), .A2(n9413), .ZN(n6546) );
  OR2_X1 U7885 ( .A1(n6467), .A2(n9924), .ZN(n6224) );
  INV_X1 U7886 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U7887 ( .A1(n6227), .A2(n6226), .ZN(n6228) );
  INV_X1 U7888 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n6232) );
  NAND2_X1 U7889 ( .A1(n6353), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n6230) );
  NAND2_X1 U7890 ( .A1(n6349), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6229) );
  OAI211_X1 U7891 ( .C1(n6232), .C2(n6231), .A(n6230), .B(n6229), .ZN(n6233)
         );
  AND2_X1 U7892 ( .A1(n9770), .A2(n9413), .ZN(n6237) );
  INV_X1 U7893 ( .A(n6237), .ZN(n6234) );
  OR2_X1 U7894 ( .A1(n6544), .A2(n6569), .ZN(n6236) );
  NAND2_X1 U7895 ( .A1(n6241), .A2(n6290), .ZN(n6242) );
  XNOR2_X1 U7896 ( .A(n6244), .B(n6289), .ZN(n6279) );
  XNOR2_X1 U7897 ( .A(n6246), .B(n7616), .ZN(n6245) );
  INV_X1 U7898 ( .A(n6279), .ZN(n6608) );
  NAND2_X1 U7899 ( .A1(n6712), .A2(n10089), .ZN(n10128) );
  NAND2_X1 U7900 ( .A1(n6721), .A2(n7666), .ZN(n10056) );
  INV_X1 U7901 ( .A(n7772), .ZN(n6248) );
  NAND2_X1 U7902 ( .A1(n6248), .A2(n6247), .ZN(n7774) );
  NAND2_X1 U7903 ( .A1(n7981), .A2(n6715), .ZN(n6249) );
  AND2_X1 U7904 ( .A1(n6579), .A2(n7717), .ZN(n6575) );
  NAND2_X1 U7905 ( .A1(n7716), .A2(n6575), .ZN(n6250) );
  AND2_X1 U7906 ( .A1(n6525), .A2(n6363), .ZN(n6584) );
  NAND2_X1 U7907 ( .A1(n10144), .A2(n9730), .ZN(n6375) );
  INV_X1 U7908 ( .A(n7924), .ZN(n6251) );
  OR2_X1 U7909 ( .A1(n7920), .A2(n5046), .ZN(n6255) );
  INV_X1 U7910 ( .A(n8018), .ZN(n6252) );
  NOR2_X1 U7911 ( .A1(n8032), .A2(n6252), .ZN(n7921) );
  AND2_X1 U7912 ( .A1(n7921), .A2(n7924), .ZN(n6253) );
  NAND2_X1 U7913 ( .A1(n7923), .A2(n6378), .ZN(n8039) );
  NAND2_X1 U7914 ( .A1(n9888), .A2(n9876), .ZN(n6385) );
  AND2_X1 U7915 ( .A1(n6380), .A2(n6385), .ZN(n6494) );
  AND2_X1 U7916 ( .A1(n9734), .A2(n6494), .ZN(n6257) );
  INV_X1 U7917 ( .A(n6494), .ZN(n6256) );
  NOR2_X1 U7918 ( .A1(n9888), .A2(n9876), .ZN(n8041) );
  NAND2_X1 U7919 ( .A1(n6380), .A2(n8041), .ZN(n6258) );
  AND2_X1 U7920 ( .A1(n6258), .A2(n6368), .ZN(n8175) );
  NOR2_X1 U7921 ( .A1(n9872), .A2(n9877), .ZN(n6395) );
  NOR2_X1 U7922 ( .A1(n6395), .A2(n6496), .ZN(n8183) );
  INV_X1 U7923 ( .A(n6496), .ZN(n6504) );
  XNOR2_X1 U7924 ( .A(n9864), .B(n9868), .ZN(n8192) );
  OR2_X1 U7925 ( .A1(n9864), .A2(n9868), .ZN(n6507) );
  NAND2_X1 U7926 ( .A1(n6259), .A2(n6403), .ZN(n9704) );
  INV_X1 U7927 ( .A(n9696), .ZN(n9861) );
  NOR2_X1 U7928 ( .A1(n9856), .A2(n9861), .ZN(n6510) );
  AOI21_X2 U7929 ( .B1(n9702), .B2(n9704), .A(n6510), .ZN(n9694) );
  NAND2_X1 U7930 ( .A1(n9847), .A2(n9834), .ZN(n9647) );
  NAND2_X1 U7931 ( .A1(n6416), .A2(n9647), .ZN(n6518) );
  OR2_X1 U7932 ( .A1(n9847), .A2(n9834), .ZN(n9648) );
  AND2_X1 U7933 ( .A1(n6407), .A2(n9648), .ZN(n6531) );
  OR2_X1 U7934 ( .A1(n6853), .A2(n9835), .ZN(n6414) );
  NAND2_X1 U7935 ( .A1(n6853), .A2(n9835), .ZN(n6586) );
  NAND2_X1 U7936 ( .A1(n6414), .A2(n6586), .ZN(n9636) );
  INV_X1 U7937 ( .A(n6586), .ZN(n6528) );
  INV_X1 U7938 ( .A(n9614), .ZN(n9813) );
  NAND2_X1 U7939 ( .A1(n9823), .A2(n9813), .ZN(n6412) );
  AND2_X1 U7940 ( .A1(n6859), .A2(n9614), .ZN(n6558) );
  NAND2_X1 U7941 ( .A1(n9600), .A2(n9814), .ZN(n6555) );
  OR2_X1 U7942 ( .A1(n6260), .A2(n9791), .ZN(n6556) );
  NAND2_X1 U7943 ( .A1(n9795), .A2(n9547), .ZN(n6424) );
  NAND2_X1 U7944 ( .A1(n6260), .A2(n9791), .ZN(n9561) );
  INV_X1 U7945 ( .A(n9795), .ZN(n6261) );
  OR2_X1 U7946 ( .A1(n9776), .A2(n9548), .ZN(n6543) );
  NAND2_X1 U7947 ( .A1(n9776), .A2(n9548), .ZN(n6548) );
  OAI21_X2 U7948 ( .B1(n8361), .B2(n8360), .A(n6548), .ZN(n8342) );
  NAND2_X1 U7949 ( .A1(n6263), .A2(n9518), .ZN(n6266) );
  NAND2_X1 U7950 ( .A1(n6246), .A2(n10052), .ZN(n6265) );
  NAND2_X1 U7951 ( .A1(n6264), .A2(n6608), .ZN(n6482) );
  NAND2_X1 U7952 ( .A1(n6266), .A2(n10168), .ZN(n6278) );
  INV_X1 U7953 ( .A(n6268), .ZN(n9530) );
  NAND2_X1 U7954 ( .A1(n9530), .A2(n6205), .ZN(n6274) );
  INV_X1 U7955 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n10397) );
  NAND2_X1 U7956 ( .A1(n6353), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7957 ( .A1(n6348), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6269) );
  OAI211_X1 U7958 ( .C1(n6271), .C2(n10397), .A(n6270), .B(n6269), .ZN(n6272)
         );
  INV_X1 U7959 ( .A(n6272), .ZN(n6273) );
  INV_X1 U7960 ( .A(n7088), .ZN(n6928) );
  NAND2_X1 U7961 ( .A1(n6278), .A2(n6277), .ZN(n8410) );
  INV_X1 U7962 ( .A(n8410), .ZN(n6286) );
  INV_X1 U7963 ( .A(n7666), .ZN(n10049) );
  NOR2_X2 U7964 ( .A1(n10048), .A2(n6715), .ZN(n7986) );
  INV_X1 U7965 ( .A(n10162), .ZN(n8001) );
  INV_X1 U7966 ( .A(n6782), .ZN(n9963) );
  AND2_X2 U7967 ( .A1(n9739), .A2(n9963), .ZN(n8058) );
  INV_X1 U7968 ( .A(n9888), .ZN(n8060) );
  NOR2_X2 U7969 ( .A1(n8188), .A2(n9864), .ZN(n9715) );
  INV_X1 U7970 ( .A(n9856), .ZN(n9714) );
  NAND2_X1 U7971 ( .A1(n9715), .A2(n9714), .ZN(n9716) );
  INV_X1 U7972 ( .A(n9662), .ZN(n9656) );
  AND2_X2 U7973 ( .A1(n9610), .A2(n9807), .ZN(n9594) );
  OR2_X1 U7974 ( .A1(n9545), .A2(n9795), .ZN(n8357) );
  OR2_X1 U7975 ( .A1(n8357), .A2(n9776), .ZN(n6280) );
  NOR2_X1 U7976 ( .A1(n6283), .A2(n8345), .ZN(n6282) );
  INV_X1 U7977 ( .A(n7628), .ZN(n6281) );
  OAI21_X1 U7978 ( .B1(n6283), .B2(n10130), .A(n8408), .ZN(n6284) );
  NAND3_X1 U7979 ( .A1(n5060), .A2(n6286), .A3(n6285), .ZN(n6323) );
  INV_X1 U7980 ( .A(n6287), .ZN(n6292) );
  INV_X1 U7981 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6288) );
  NAND3_X1 U7982 ( .A1(n6290), .A2(n6289), .A3(n6288), .ZN(n6291) );
  OAI21_X1 U7983 ( .B1(n6292), .B2(n6291), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n6294) );
  XNOR2_X1 U7984 ( .A(n6294), .B(n6293), .ZN(n6954) );
  INV_X1 U7985 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6296) );
  NAND2_X1 U7986 ( .A1(n6295), .A2(n6296), .ZN(n6297) );
  NAND2_X1 U7987 ( .A1(n6297), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6298) );
  XNOR2_X1 U7988 ( .A(n6295), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7989 ( .A1(n4998), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6299) );
  XNOR2_X1 U7990 ( .A(n6299), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6302) );
  AND2_X1 U7991 ( .A1(n6301), .A2(n6302), .ZN(n6300) );
  INV_X1 U7992 ( .A(n6301), .ZN(n8313) );
  NAND2_X1 U7993 ( .A1(n8313), .A2(P1_B_REG_SCAN_IN), .ZN(n6303) );
  INV_X1 U7994 ( .A(n6302), .ZN(n8235) );
  MUX2_X1 U7995 ( .A(P1_B_REG_SCAN_IN), .B(n6303), .S(n8235), .Z(n6304) );
  INV_X1 U7996 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U7997 ( .A1(n7037), .A2(n6305), .ZN(n6308) );
  INV_X1 U7998 ( .A(n6306), .ZN(n8335) );
  NAND2_X1 U7999 ( .A1(n8335), .A2(n8313), .ZN(n6307) );
  NAND2_X1 U8000 ( .A1(n6308), .A2(n6307), .ZN(n7609) );
  NOR2_X1 U8001 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_2__SCAN_IN), .ZN(
        n10429) );
  NOR4_X1 U8002 ( .A1(P1_D_REG_30__SCAN_IN), .A2(P1_D_REG_31__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6311) );
  NOR4_X1 U8003 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n6310) );
  NOR4_X1 U8004 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_6__SCAN_IN), .ZN(n6309) );
  AND4_X1 U8005 ( .A1(n10429), .A2(n6311), .A3(n6310), .A4(n6309), .ZN(n6317)
         );
  NOR4_X1 U8006 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n6315) );
  NOR4_X1 U8007 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_15__SCAN_IN), .ZN(n6314) );
  NOR4_X1 U8008 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n6313) );
  NOR4_X1 U8009 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6312) );
  AND4_X1 U8010 ( .A1(n6315), .A2(n6314), .A3(n6313), .A4(n6312), .ZN(n6316)
         );
  NAND2_X1 U8011 ( .A1(n6317), .A2(n6316), .ZN(n6318) );
  NAND2_X1 U8012 ( .A1(n7037), .A2(n6318), .ZN(n7608) );
  AND2_X1 U8013 ( .A1(n7609), .A2(n7608), .ZN(n6320) );
  OR2_X1 U8014 ( .A1(n10089), .A2(n6264), .ZN(n6319) );
  INV_X1 U8015 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n7039) );
  INV_X1 U8016 ( .A(n7611), .ZN(n6321) );
  NAND2_X1 U8017 ( .A1(n6323), .A2(n10177), .ZN(n6325) );
  NAND2_X1 U8018 ( .A1(n6325), .A2(n6324), .ZN(P1_U3551) );
  INV_X1 U8019 ( .A(SI_28_), .ZN(n6326) );
  NAND2_X1 U8020 ( .A1(n6327), .A2(n6326), .ZN(n6334) );
  INV_X1 U8021 ( .A(n6334), .ZN(n6329) );
  AND2_X1 U8022 ( .A1(n6330), .A2(n6333), .ZN(n6331) );
  INV_X1 U8023 ( .A(n6333), .ZN(n6339) );
  AND2_X1 U8024 ( .A1(n6335), .A2(n6334), .ZN(n6337) );
  AND2_X1 U8025 ( .A1(n6337), .A2(n6336), .ZN(n6338) );
  INV_X1 U8026 ( .A(SI_29_), .ZN(n6343) );
  INV_X1 U8027 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n6342) );
  INV_X1 U8028 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10444) );
  MUX2_X1 U8029 ( .A(n6342), .B(n10444), .S(n6344), .Z(n6454) );
  MUX2_X1 U8030 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n6344), .Z(n6462) );
  INV_X1 U8031 ( .A(SI_30_), .ZN(n6460) );
  XNOR2_X1 U8032 ( .A(n6462), .B(n6460), .ZN(n6345) );
  NAND2_X1 U8033 ( .A1(n9275), .A2(n6469), .ZN(n6347) );
  INV_X1 U8034 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n9918) );
  OR2_X1 U8035 ( .A1(n6467), .A2(n9918), .ZN(n6346) );
  NAND2_X1 U8036 ( .A1(n6353), .A2(P1_REG1_REG_30__SCAN_IN), .ZN(n6352) );
  NAND2_X1 U8037 ( .A1(n6348), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6351) );
  NAND2_X1 U8038 ( .A1(n6349), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6350) );
  AND3_X1 U8039 ( .A1(n6352), .A2(n6351), .A3(n6350), .ZN(n9521) );
  INV_X1 U8040 ( .A(n9521), .ZN(n9434) );
  NAND2_X1 U8041 ( .A1(n6349), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6356) );
  NAND2_X1 U8042 ( .A1(n6353), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U8043 ( .A1(n6348), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6354) );
  NAND3_X1 U8044 ( .A1(n6356), .A2(n6355), .A3(n6354), .ZN(n9505) );
  NAND2_X1 U8045 ( .A1(n9434), .A2(n9505), .ZN(n6357) );
  NAND2_X1 U8046 ( .A1(n9750), .A2(n6357), .ZN(n6599) );
  INV_X1 U8047 ( .A(n6473), .ZN(n6477) );
  NAND2_X1 U8048 ( .A1(n9517), .A2(n6546), .ZN(n6359) );
  NOR2_X1 U8049 ( .A1(n6440), .A2(n9783), .ZN(n6358) );
  AND2_X1 U8050 ( .A1(n9548), .A2(n6477), .ZN(n6447) );
  NAND3_X1 U8051 ( .A1(n6488), .A2(n6447), .A3(n6596), .ZN(n6360) );
  NAND2_X1 U8052 ( .A1(n6361), .A2(n6360), .ZN(n6436) );
  INV_X1 U8053 ( .A(n6518), .ZN(n6362) );
  AND2_X1 U8054 ( .A1(n6373), .A2(n6364), .ZN(n6519) );
  OAI21_X1 U8055 ( .B1(n7621), .B2(n6560), .A(n6519), .ZN(n6366) );
  NAND2_X1 U8056 ( .A1(n6376), .A2(n8018), .ZN(n6495) );
  INV_X1 U8057 ( .A(n6495), .ZN(n6365) );
  NAND2_X1 U8058 ( .A1(n6366), .A2(n6365), .ZN(n6367) );
  NAND3_X1 U8059 ( .A1(n6367), .A2(n6378), .A3(n7922), .ZN(n6371) );
  NAND2_X1 U8060 ( .A1(n6379), .A2(n6375), .ZN(n6492) );
  INV_X1 U8061 ( .A(n6492), .ZN(n6370) );
  XNOR2_X1 U8062 ( .A(n9888), .B(n9876), .ZN(n8055) );
  INV_X1 U8063 ( .A(n8055), .ZN(n8067) );
  NAND4_X1 U8064 ( .A1(n6368), .A2(n6477), .A3(n8040), .A4(n8067), .ZN(n6369)
         );
  AOI21_X1 U8065 ( .B1(n6371), .B2(n6370), .A(n6369), .ZN(n6394) );
  INV_X1 U8066 ( .A(n6560), .ZN(n7620) );
  NAND2_X1 U8067 ( .A1(n7621), .A2(n7620), .ZN(n6372) );
  NAND3_X1 U8068 ( .A1(n6374), .A2(n7922), .A3(n6373), .ZN(n6377) );
  NAND3_X1 U8069 ( .A1(n6377), .A2(n6376), .A3(n6375), .ZN(n6383) );
  NAND2_X1 U8070 ( .A1(n8040), .A2(n6378), .ZN(n6500) );
  INV_X1 U8071 ( .A(n6500), .ZN(n6382) );
  NAND4_X1 U8072 ( .A1(n6380), .A2(n6379), .A3(n6473), .A4(n8067), .ZN(n6381)
         );
  AOI21_X1 U8073 ( .B1(n6383), .B2(n6382), .A(n6381), .ZN(n6393) );
  INV_X1 U8074 ( .A(n8175), .ZN(n6384) );
  OR2_X1 U8075 ( .A1(n6384), .A2(n6395), .ZN(n6506) );
  NAND2_X1 U8076 ( .A1(n6506), .A2(n6473), .ZN(n6391) );
  NOR2_X1 U8077 ( .A1(n6385), .A2(n9440), .ZN(n6387) );
  AOI21_X1 U8078 ( .B1(n6385), .B2(n9440), .A(n6473), .ZN(n6386) );
  OAI21_X1 U8079 ( .B1(n6387), .B2(n9880), .A(n6386), .ZN(n6388) );
  INV_X1 U8080 ( .A(n6388), .ZN(n6389) );
  NOR2_X1 U8081 ( .A1(n6496), .A2(n6389), .ZN(n6390) );
  NAND2_X1 U8082 ( .A1(n9864), .A2(n9868), .ZN(n6490) );
  NAND4_X1 U8083 ( .A1(n6391), .A2(n6390), .A3(n6507), .A4(n6490), .ZN(n6392)
         );
  INV_X1 U8084 ( .A(n6395), .ZN(n6396) );
  NAND2_X1 U8085 ( .A1(n6396), .A2(n6507), .ZN(n6397) );
  NAND2_X1 U8086 ( .A1(n6397), .A2(n6490), .ZN(n6400) );
  NAND2_X1 U8087 ( .A1(n6490), .A2(n6504), .ZN(n6398) );
  NAND2_X1 U8088 ( .A1(n6398), .A2(n6507), .ZN(n6399) );
  MUX2_X1 U8089 ( .A(n6400), .B(n6399), .S(n6473), .Z(n6401) );
  MUX2_X1 U8090 ( .A(n9856), .B(n9696), .S(n6473), .Z(n6404) );
  NAND2_X1 U8091 ( .A1(n6404), .A2(n6403), .ZN(n6405) );
  NAND2_X1 U8092 ( .A1(n9648), .A2(n9647), .ZN(n9670) );
  INV_X1 U8093 ( .A(n9670), .ZN(n9671) );
  MUX2_X1 U8094 ( .A(n6512), .B(n6515), .S(n6473), .Z(n6406) );
  NAND3_X1 U8095 ( .A1(n6418), .A2(n6407), .A3(n6414), .ZN(n6409) );
  AND2_X1 U8096 ( .A1(n6412), .A2(n6586), .ZN(n6408) );
  AOI21_X1 U8097 ( .B1(n6409), .B2(n6408), .A(n6558), .ZN(n6410) );
  INV_X1 U8098 ( .A(n6593), .ZN(n6538) );
  INV_X1 U8099 ( .A(n6412), .ZN(n6557) );
  NAND2_X1 U8100 ( .A1(n6415), .A2(n6557), .ZN(n6413) );
  NAND3_X1 U8101 ( .A1(n6555), .A2(n5015), .A3(n6413), .ZN(n6589) );
  NAND3_X1 U8102 ( .A1(n5020), .A2(n6415), .A3(n6414), .ZN(n6534) );
  NAND2_X1 U8103 ( .A1(n6586), .A2(n6416), .ZN(n6532) );
  INV_X1 U8104 ( .A(n6532), .ZN(n6417) );
  OR2_X1 U8105 ( .A1(n6589), .A2(n6419), .ZN(n6420) );
  MUX2_X1 U8106 ( .A(n6421), .B(n6420), .S(n6473), .Z(n6429) );
  NAND2_X1 U8107 ( .A1(n6429), .A2(n6538), .ZN(n6422) );
  NAND2_X1 U8108 ( .A1(n6422), .A2(n6427), .ZN(n6426) );
  INV_X1 U8109 ( .A(n6556), .ZN(n6423) );
  OR2_X1 U8110 ( .A1(n6541), .A2(n6423), .ZN(n6594) );
  NAND2_X1 U8111 ( .A1(n6594), .A2(n6424), .ZN(n6425) );
  NAND3_X1 U8112 ( .A1(n6426), .A2(n6425), .A3(n6542), .ZN(n6435) );
  OR2_X1 U8113 ( .A1(n6427), .A2(n6541), .ZN(n6428) );
  NAND2_X1 U8114 ( .A1(n6428), .A2(n6440), .ZN(n6597) );
  INV_X1 U8115 ( .A(n6597), .ZN(n6433) );
  INV_X1 U8116 ( .A(n6594), .ZN(n6431) );
  NAND2_X1 U8117 ( .A1(n6429), .A2(n6555), .ZN(n6430) );
  NAND2_X1 U8118 ( .A1(n6433), .A2(n6432), .ZN(n6434) );
  OR2_X1 U8119 ( .A1(n9517), .A2(n6473), .ZN(n6438) );
  NAND3_X1 U8120 ( .A1(n9517), .A2(n6549), .A3(n6473), .ZN(n6437) );
  AND2_X1 U8121 ( .A1(n9776), .A2(n6542), .ZN(n6439) );
  MUX2_X1 U8122 ( .A(n6439), .B(n9783), .S(n6473), .Z(n6441) );
  NAND4_X1 U8123 ( .A1(n6488), .A2(n6477), .A3(n6596), .A4(n6441), .ZN(n6444)
         );
  AND2_X1 U8124 ( .A1(n6440), .A2(n6473), .ZN(n6442) );
  NAND4_X1 U8125 ( .A1(n9517), .A2(n6442), .A3(n6546), .A4(n6441), .ZN(n6443)
         );
  NAND2_X1 U8126 ( .A1(n6444), .A2(n6443), .ZN(n6446) );
  NAND2_X1 U8127 ( .A1(n6446), .A2(n6445), .ZN(n6453) );
  INV_X1 U8128 ( .A(n6447), .ZN(n6448) );
  OAI22_X1 U8129 ( .A1(n6546), .A2(n6473), .B1(n9418), .B2(n6448), .ZN(n6449)
         );
  NAND2_X1 U8130 ( .A1(n6449), .A2(n6596), .ZN(n6450) );
  NAND2_X1 U8131 ( .A1(n6450), .A2(n6488), .ZN(n6451) );
  OAI21_X1 U8132 ( .B1(n6473), .B2(n6488), .A(n6451), .ZN(n6452) );
  NAND2_X1 U8133 ( .A1(n6470), .A2(n9758), .ZN(n6459) );
  XNOR2_X1 U8134 ( .A(n6454), .B(SI_29_), .ZN(n6455) );
  NAND2_X1 U8135 ( .A1(n8412), .A2(n6469), .ZN(n6458) );
  OR2_X1 U8136 ( .A1(n6467), .A2(n10444), .ZN(n6457) );
  OR2_X1 U8137 ( .A1(n9750), .A2(n9521), .ZN(n6487) );
  NAND2_X1 U8138 ( .A1(n6487), .A2(n9505), .ZN(n6474) );
  MUX2_X1 U8139 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n6463), .Z(n6464) );
  XNOR2_X1 U8140 ( .A(n6464), .B(SI_31_), .ZN(n6465) );
  INV_X1 U8141 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n9912) );
  NOR2_X1 U8142 ( .A1(n6467), .A2(n9912), .ZN(n6468) );
  INV_X1 U8143 ( .A(n9508), .ZN(n9746) );
  NAND2_X1 U8144 ( .A1(n6474), .A2(n9746), .ZN(n6605) );
  INV_X1 U8145 ( .A(n6470), .ZN(n6472) );
  INV_X1 U8146 ( .A(n9758), .ZN(n9760) );
  NAND3_X1 U8147 ( .A1(n6472), .A2(n6477), .A3(n9760), .ZN(n6471) );
  NAND2_X1 U8148 ( .A1(n6599), .A2(n6473), .ZN(n6478) );
  AOI21_X1 U8149 ( .B1(n6472), .B2(n9757), .A(n6478), .ZN(n6476) );
  AOI21_X1 U8150 ( .B1(n6474), .B2(n9746), .A(n6473), .ZN(n6475) );
  OAI22_X1 U8151 ( .A1(n6478), .A2(n6487), .B1(n6477), .B2(n9505), .ZN(n6479)
         );
  NAND2_X1 U8152 ( .A1(n6479), .A2(n9746), .ZN(n6480) );
  AND2_X1 U8153 ( .A1(n9508), .A2(n9505), .ZN(n6603) );
  OR2_X1 U8154 ( .A1(n6954), .A2(P1_U3084), .ZN(n8015) );
  NAND2_X1 U8155 ( .A1(n6608), .A2(n10052), .ZN(n6484) );
  NOR4_X1 U8156 ( .A1(n6603), .A2(n7088), .A3(n8015), .A4(n6484), .ZN(n6485)
         );
  NAND2_X1 U8157 ( .A1(n6486), .A2(n6485), .ZN(n6621) );
  OAI21_X1 U8158 ( .B1(n9508), .B2(n9505), .A(n6487), .ZN(n6573) );
  OR2_X1 U8159 ( .A1(n9757), .A2(n9758), .ZN(n6489) );
  AND2_X1 U8160 ( .A1(n6489), .A2(n6488), .ZN(n6552) );
  INV_X1 U8161 ( .A(n6552), .ZN(n6602) );
  NAND2_X1 U8162 ( .A1(n9856), .A2(n9861), .ZN(n6491) );
  AND2_X1 U8163 ( .A1(n6491), .A2(n6490), .ZN(n6509) );
  NAND2_X1 U8164 ( .A1(n6492), .A2(n8040), .ZN(n6493) );
  AND2_X1 U8165 ( .A1(n6494), .A2(n6493), .ZN(n6499) );
  NOR2_X1 U8166 ( .A1(n6496), .A2(n6495), .ZN(n6497) );
  NAND4_X1 U8167 ( .A1(n6515), .A2(n6509), .A3(n6499), .A4(n6497), .ZN(n6498)
         );
  NOR2_X1 U8168 ( .A1(n6518), .A2(n6498), .ZN(n6585) );
  INV_X1 U8169 ( .A(n6585), .ZN(n6520) );
  INV_X1 U8170 ( .A(n6499), .ZN(n6503) );
  INV_X1 U8171 ( .A(n7922), .ZN(n6501) );
  NOR2_X1 U8172 ( .A1(n6501), .A2(n6500), .ZN(n6502) );
  NOR2_X1 U8173 ( .A1(n6503), .A2(n6502), .ZN(n6505) );
  OAI21_X1 U8174 ( .B1(n6506), .B2(n6505), .A(n6504), .ZN(n6508) );
  AND2_X1 U8175 ( .A1(n6508), .A2(n6507), .ZN(n6514) );
  INV_X1 U8176 ( .A(n6509), .ZN(n6513) );
  INV_X1 U8177 ( .A(n6510), .ZN(n6511) );
  OAI211_X1 U8178 ( .C1(n6514), .C2(n6513), .A(n6512), .B(n6511), .ZN(n6516)
         );
  NAND2_X1 U8179 ( .A1(n6516), .A2(n6515), .ZN(n6517) );
  OAI22_X1 U8180 ( .A1(n6520), .A2(n6519), .B1(n6518), .B2(n6517), .ZN(n6587)
         );
  INV_X1 U8181 ( .A(n6587), .ZN(n6530) );
  OR2_X1 U8182 ( .A1(n6721), .A2(n7666), .ZN(n7087) );
  NAND2_X1 U8183 ( .A1(n7087), .A2(n10055), .ZN(n6559) );
  INV_X1 U8184 ( .A(n6559), .ZN(n6522) );
  AOI21_X1 U8185 ( .B1(n6711), .B2(n7768), .A(n7698), .ZN(n6521) );
  NAND3_X1 U8186 ( .A1(n6522), .A2(n6575), .A3(n6521), .ZN(n6523) );
  NAND2_X1 U8187 ( .A1(n6523), .A2(n6584), .ZN(n6526) );
  INV_X1 U8188 ( .A(n6580), .ZN(n6524) );
  NAND2_X1 U8189 ( .A1(n6525), .A2(n6524), .ZN(n6574) );
  OAI21_X1 U8190 ( .B1(n10034), .B2(n6526), .A(n6574), .ZN(n6527) );
  NAND2_X1 U8191 ( .A1(n6585), .A2(n6527), .ZN(n6529) );
  AOI21_X1 U8192 ( .B1(n6530), .B2(n6529), .A(n6528), .ZN(n6537) );
  NOR2_X1 U8193 ( .A1(n6532), .A2(n6531), .ZN(n6533) );
  NOR2_X1 U8194 ( .A1(n6534), .A2(n6533), .ZN(n6591) );
  INV_X1 U8195 ( .A(n6591), .ZN(n6536) );
  INV_X1 U8196 ( .A(n6589), .ZN(n6535) );
  OAI21_X1 U8197 ( .B1(n6537), .B2(n6536), .A(n6535), .ZN(n6539) );
  NAND3_X1 U8198 ( .A1(n6539), .A2(n6556), .A3(n6538), .ZN(n6540) );
  NOR2_X1 U8199 ( .A1(n6541), .A2(n6540), .ZN(n6545) );
  AND2_X1 U8200 ( .A1(n6543), .A2(n6542), .ZN(n6595) );
  OAI211_X1 U8201 ( .C1(n6545), .C2(n6597), .A(n6544), .B(n6595), .ZN(n6553)
         );
  AND2_X1 U8202 ( .A1(n9517), .A2(n6546), .ZN(n6547) );
  OAI21_X1 U8203 ( .B1(n6549), .B2(n6548), .A(n6547), .ZN(n6551) );
  AND2_X1 U8204 ( .A1(n9757), .A2(n9758), .ZN(n6550) );
  AOI21_X1 U8205 ( .B1(n6552), .B2(n6551), .A(n6550), .ZN(n6600) );
  NAND2_X1 U8206 ( .A1(n9750), .A2(n9521), .ZN(n6570) );
  OAI211_X1 U8207 ( .C1(n6602), .C2(n6553), .A(n6600), .B(n6570), .ZN(n6554)
         );
  AOI21_X1 U8208 ( .B1(n4568), .B2(n6554), .A(n6603), .ZN(n6615) );
  INV_X1 U8209 ( .A(n6603), .ZN(n6572) );
  INV_X1 U8210 ( .A(n9606), .ZN(n9605) );
  NAND2_X1 U8211 ( .A1(n6556), .A2(n9561), .ZN(n9578) );
  NOR2_X1 U8212 ( .A1(n6558), .A2(n6557), .ZN(n9621) );
  NOR2_X1 U8213 ( .A1(n10061), .A2(n6559), .ZN(n6563) );
  NOR2_X1 U8214 ( .A1(n6560), .A2(n7719), .ZN(n6562) );
  INV_X1 U8215 ( .A(n7985), .ZN(n6561) );
  INV_X1 U8216 ( .A(n7920), .ZN(n7999) );
  NAND3_X1 U8217 ( .A1(n9704), .A2(n8183), .A3(n6565), .ZN(n6566) );
  XNOR2_X1 U8218 ( .A(n9795), .B(n9782), .ZN(n9563) );
  NOR4_X1 U8219 ( .A1(n6569), .A2(n8360), .A3(n6568), .A4(n6567), .ZN(n6571)
         );
  INV_X1 U8220 ( .A(n9754), .ZN(n9755) );
  NAND3_X1 U8221 ( .A1(n6576), .A2(n6575), .A3(n6574), .ZN(n6583) );
  INV_X1 U8222 ( .A(n6577), .ZN(n6581) );
  OAI211_X1 U8223 ( .C1(n6581), .C2(n4993), .A(n6580), .B(n6579), .ZN(n6582)
         );
  AND4_X1 U8224 ( .A1(n6585), .A2(n6584), .A3(n6583), .A4(n6582), .ZN(n6588)
         );
  OAI21_X1 U8225 ( .B1(n6588), .B2(n6587), .A(n6586), .ZN(n6590) );
  AOI21_X1 U8226 ( .B1(n6591), .B2(n6590), .A(n6589), .ZN(n6592) );
  NOR3_X1 U8227 ( .A1(n6594), .A2(n6593), .A3(n6592), .ZN(n6598) );
  OAI211_X1 U8228 ( .C1(n6598), .C2(n6597), .A(n6596), .B(n6595), .ZN(n6601)
         );
  OAI211_X1 U8229 ( .C1(n6602), .C2(n6601), .A(n6600), .B(n6599), .ZN(n6604)
         );
  AOI211_X1 U8230 ( .C1(n6605), .C2(n6604), .A(n7698), .B(n6603), .ZN(n6606)
         );
  NAND3_X1 U8231 ( .A1(n6609), .A2(n6608), .A3(n6607), .ZN(n6613) );
  NAND2_X1 U8232 ( .A1(n6279), .A2(n10052), .ZN(n6610) );
  INV_X1 U8233 ( .A(n8015), .ZN(n6618) );
  NAND2_X1 U8234 ( .A1(n6613), .A2(n6612), .ZN(n6614) );
  INV_X1 U8235 ( .A(P1_B_REG_SCAN_IN), .ZN(n9503) );
  INV_X1 U8236 ( .A(n7614), .ZN(n7097) );
  INV_X1 U8237 ( .A(n6925), .ZN(n7627) );
  NOR4_X1 U8238 ( .A1(n10138), .A2(n7097), .A3(n9504), .A4(n7627), .ZN(n6617)
         );
  AOI211_X1 U8239 ( .C1(n6618), .C2(n6714), .A(n9503), .B(n6617), .ZN(n6619)
         );
  NAND3_X1 U8240 ( .A1(n6622), .A2(n6621), .A3(n5058), .ZN(P1_U3240) );
  NAND2_X1 U8241 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6636), .ZN(n10203) );
  NAND2_X1 U8242 ( .A1(n6630), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n6623) );
  OAI21_X1 U8243 ( .B1(n6630), .B2(P2_REG2_REG_16__SCAN_IN), .A(n6623), .ZN(
        n8893) );
  INV_X1 U8244 ( .A(n7975), .ZN(n7085) );
  INV_X1 U8245 ( .A(n7513), .ZN(n7055) );
  INV_X1 U8246 ( .A(n6683), .ZN(n7424) );
  INV_X1 U8247 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n6627) );
  INV_X1 U8248 ( .A(n6682), .ZN(n7320) );
  INV_X1 U8249 ( .A(n6678), .ZN(n7384) );
  INV_X1 U8250 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7911) );
  INV_X1 U8251 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7900) );
  INV_X1 U8252 ( .A(n6675), .ZN(n7395) );
  INV_X1 U8253 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7889) );
  INV_X1 U8254 ( .A(n8879), .ZN(n7029) );
  INV_X1 U8255 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n7870) );
  INV_X1 U8256 ( .A(n8849), .ZN(n7001) );
  INV_X1 U8257 ( .A(n7373), .ZN(n7381) );
  INV_X1 U8258 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7809) );
  INV_X1 U8259 ( .A(n8834), .ZN(n7006) );
  INV_X1 U8260 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7642) );
  INV_X1 U8261 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7600) );
  INV_X1 U8262 ( .A(n8821), .ZN(n7005) );
  INV_X1 U8263 ( .A(n8805), .ZN(n6999) );
  INV_X1 U8264 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6625) );
  XOR2_X1 U8265 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n8795), .Z(n8794) );
  INV_X1 U8266 ( .A(n8795), .ZN(n8369) );
  INV_X1 U8267 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6624) );
  XOR2_X1 U8268 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n8805), .Z(n8804) );
  XOR2_X1 U8269 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n8821), .Z(n8818) );
  NAND2_X1 U8270 ( .A1(n8817), .A2(n8818), .ZN(n8816) );
  OAI21_X1 U8271 ( .B1(n7600), .B2(n7005), .A(n8816), .ZN(n8830) );
  XOR2_X1 U8272 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n8834), .Z(n8831) );
  NAND2_X1 U8273 ( .A1(n8830), .A2(n8831), .ZN(n8829) );
  OAI21_X1 U8274 ( .B1(n7006), .B2(n7642), .A(n8829), .ZN(n7371) );
  XOR2_X1 U8275 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7373), .Z(n7372) );
  NAND2_X1 U8276 ( .A1(n7371), .A2(n7372), .ZN(n7370) );
  MUX2_X1 U8277 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n7870), .S(n8849), .Z(n8847)
         );
  XOR2_X1 U8278 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n8863), .Z(n8861) );
  INV_X1 U8279 ( .A(n8863), .ZN(n7016) );
  INV_X1 U8280 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6626) );
  MUX2_X1 U8281 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7889), .S(n8879), .Z(n8876)
         );
  XOR2_X1 U8282 ( .A(n6675), .B(P2_REG2_REG_9__SCAN_IN), .Z(n7399) );
  XNOR2_X1 U8283 ( .A(n6678), .B(n7911), .ZN(n7389) );
  MUX2_X1 U8284 ( .A(n7948), .B(P2_REG2_REG_11__SCAN_IN), .S(n6682), .Z(n7315)
         );
  NOR2_X1 U8285 ( .A1(n7314), .A2(n7315), .ZN(n7313) );
  XOR2_X1 U8286 ( .A(n6683), .B(P2_REG2_REG_12__SCAN_IN), .Z(n7419) );
  XNOR2_X1 U8287 ( .A(n7513), .B(P2_REG2_REG_13__SCAN_IN), .ZN(n7505) );
  MUX2_X1 U8288 ( .A(n6628), .B(P2_REG2_REG_14__SCAN_IN), .S(n7975), .Z(n7965)
         );
  NOR2_X1 U8289 ( .A1(n7964), .A2(n7965), .ZN(n7963) );
  NAND2_X1 U8290 ( .A1(n8905), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n6631) );
  OAI21_X1 U8291 ( .B1(n8905), .B2(P2_REG2_REG_17__SCAN_IN), .A(n6631), .ZN(
        n8903) );
  NOR2_X1 U8292 ( .A1(n8904), .A2(n8903), .ZN(n8902) );
  AOI21_X1 U8293 ( .B1(n8905), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8902), .ZN(
        n6632) );
  INV_X1 U8294 ( .A(n6648), .ZN(n8931) );
  NOR2_X1 U8295 ( .A1(n6632), .A2(n8931), .ZN(n6634) );
  INV_X1 U8296 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8920) );
  XNOR2_X1 U8297 ( .A(n6635), .B(n10482), .ZN(n6703) );
  NAND2_X1 U8298 ( .A1(n10178), .A2(n7269), .ZN(n6640) );
  OR2_X1 U8299 ( .A1(n6704), .A2(P2_U3152), .ZN(n8339) );
  NOR2_X1 U8300 ( .A1(n6636), .A2(P2_U3152), .ZN(n8597) );
  INV_X1 U8301 ( .A(n8597), .ZN(n8764) );
  OAI21_X1 U8302 ( .B1(n6637), .B2(n8339), .A(n8764), .ZN(n6638) );
  INV_X1 U8303 ( .A(n6638), .ZN(n6639) );
  NAND2_X1 U8304 ( .A1(n6640), .A2(n6639), .ZN(n6647) );
  AND2_X1 U8305 ( .A1(n6647), .A2(n6645), .ZN(n6641) );
  NAND2_X1 U8306 ( .A1(n6643), .A2(n6642), .ZN(n8401) );
  INV_X1 U8307 ( .A(n8401), .ZN(n8762) );
  NAND2_X1 U8308 ( .A1(n6705), .A2(n8762), .ZN(n7243) );
  INV_X1 U8309 ( .A(n6704), .ZN(n6644) );
  AND2_X1 U8310 ( .A1(n6645), .A2(n8401), .ZN(n6646) );
  OR2_X1 U8311 ( .A1(n6648), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6692) );
  NAND2_X1 U8312 ( .A1(n6648), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6649) );
  AND2_X1 U8313 ( .A1(n6692), .A2(n6649), .ZN(n8925) );
  INV_X1 U8314 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8311) );
  XNOR2_X1 U8315 ( .A(n8905), .B(n8311), .ZN(n8910) );
  XNOR2_X1 U8316 ( .A(n8896), .B(n8262), .ZN(n8891) );
  MUX2_X1 U8317 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6650), .S(n8805), .Z(n6655)
         );
  MUX2_X1 U8318 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6651), .S(n8795), .Z(n6653)
         );
  NAND2_X1 U8319 ( .A1(n6653), .A2(n6652), .ZN(n8807) );
  NAND2_X1 U8320 ( .A1(n8795), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8806) );
  NAND2_X1 U8321 ( .A1(n8807), .A2(n8806), .ZN(n6654) );
  NAND2_X1 U8322 ( .A1(n6655), .A2(n6654), .ZN(n8810) );
  NAND2_X1 U8323 ( .A1(n8805), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6656) );
  NAND2_X1 U8324 ( .A1(n8810), .A2(n6656), .ZN(n8822) );
  MUX2_X1 U8325 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6657), .S(n8821), .Z(n8823)
         );
  NAND2_X1 U8326 ( .A1(n8822), .A2(n8823), .ZN(n8837) );
  NAND2_X1 U8327 ( .A1(n8821), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n8836) );
  NAND2_X1 U8328 ( .A1(n8837), .A2(n8836), .ZN(n6660) );
  MUX2_X1 U8329 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6658), .S(n8834), .Z(n6659)
         );
  NAND2_X1 U8330 ( .A1(n6660), .A2(n6659), .ZN(n8839) );
  NAND2_X1 U8331 ( .A1(n8834), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7375) );
  NAND2_X1 U8332 ( .A1(n8839), .A2(n7375), .ZN(n6663) );
  MUX2_X1 U8333 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6661), .S(n7373), .Z(n6662)
         );
  NAND2_X1 U8334 ( .A1(n6663), .A2(n6662), .ZN(n8852) );
  NAND2_X1 U8335 ( .A1(n7373), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n8851) );
  NAND2_X1 U8336 ( .A1(n8852), .A2(n8851), .ZN(n6666) );
  MUX2_X1 U8337 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6664), .S(n8849), .Z(n6665)
         );
  NAND2_X1 U8338 ( .A1(n6666), .A2(n6665), .ZN(n8866) );
  NAND2_X1 U8339 ( .A1(n8849), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n8865) );
  NAND2_X1 U8340 ( .A1(n8866), .A2(n8865), .ZN(n6669) );
  MUX2_X1 U8341 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6667), .S(n8863), .Z(n6668)
         );
  NAND2_X1 U8342 ( .A1(n6669), .A2(n6668), .ZN(n8882) );
  NAND2_X1 U8343 ( .A1(n8863), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8881) );
  NAND2_X1 U8344 ( .A1(n8882), .A2(n8881), .ZN(n6672) );
  MUX2_X1 U8345 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6670), .S(n8879), .Z(n6671)
         );
  NAND2_X1 U8346 ( .A1(n6672), .A2(n6671), .ZN(n8884) );
  NAND2_X1 U8347 ( .A1(n8879), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6673) );
  NAND2_X1 U8348 ( .A1(n8884), .A2(n6673), .ZN(n7394) );
  XNOR2_X1 U8349 ( .A(n6675), .B(n6674), .ZN(n7393) );
  NAND2_X1 U8350 ( .A1(n7394), .A2(n7393), .ZN(n6677) );
  NAND2_X1 U8351 ( .A1(n6675), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6676) );
  NAND2_X1 U8352 ( .A1(n6677), .A2(n6676), .ZN(n7383) );
  XNOR2_X1 U8353 ( .A(n6678), .B(n10524), .ZN(n7382) );
  NAND2_X1 U8354 ( .A1(n7383), .A2(n7382), .ZN(n6680) );
  NAND2_X1 U8355 ( .A1(n6678), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6679) );
  NAND2_X1 U8356 ( .A1(n6680), .A2(n6679), .ZN(n7312) );
  INV_X1 U8357 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6681) );
  XNOR2_X1 U8358 ( .A(n6682), .B(n6681), .ZN(n7311) );
  AOI22_X1 U8359 ( .A1(n7312), .A2(n7311), .B1(P2_REG1_REG_11__SCAN_IN), .B2(
        n6682), .ZN(n7421) );
  NOR2_X1 U8360 ( .A1(n6683), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6684) );
  AOI21_X1 U8361 ( .B1(n6683), .B2(P2_REG1_REG_12__SCAN_IN), .A(n6684), .ZN(
        n7422) );
  NAND2_X1 U8362 ( .A1(n7421), .A2(n7422), .ZN(n7508) );
  INV_X1 U8363 ( .A(n6684), .ZN(n7507) );
  OR2_X1 U8364 ( .A1(n7513), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6686) );
  NAND2_X1 U8365 ( .A1(n7513), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n6685) );
  NAND2_X1 U8366 ( .A1(n6686), .A2(n6685), .ZN(n7506) );
  AOI21_X1 U8367 ( .B1(n7508), .B2(n7507), .A(n7506), .ZN(n7970) );
  INV_X1 U8368 ( .A(n6686), .ZN(n7969) );
  INV_X1 U8369 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n6687) );
  XNOR2_X1 U8370 ( .A(n7975), .B(n6687), .ZN(n7968) );
  OAI21_X1 U8371 ( .B1(n7970), .B2(n7969), .A(n7968), .ZN(n7972) );
  OAI21_X1 U8372 ( .B1(P2_REG1_REG_14__SCAN_IN), .B2(n7975), .A(n7972), .ZN(
        n6689) );
  XOR2_X1 U8373 ( .A(n6688), .B(n6689), .Z(n8271) );
  INV_X1 U8374 ( .A(n6688), .ZN(n8274) );
  OAI22_X1 U8375 ( .A1(n8271), .A2(n6690), .B1(n8274), .B2(n6689), .ZN(n8892)
         );
  NOR2_X1 U8376 ( .A1(n8891), .A2(n8892), .ZN(n8890) );
  AOI21_X1 U8377 ( .B1(n8896), .B2(n8262), .A(n8890), .ZN(n8909) );
  NAND2_X1 U8378 ( .A1(n8910), .A2(n8909), .ZN(n8908) );
  INV_X1 U8379 ( .A(n8908), .ZN(n6691) );
  AOI21_X1 U8380 ( .B1(n8905), .B2(P2_REG1_REG_17__SCAN_IN), .A(n6691), .ZN(
        n8924) );
  NAND2_X1 U8381 ( .A1(n8925), .A2(n8924), .ZN(n8923) );
  NAND2_X1 U8382 ( .A1(n8923), .A2(n6692), .ZN(n6693) );
  XNOR2_X1 U8383 ( .A(n6693), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n6707) );
  INV_X1 U8384 ( .A(n6707), .ZN(n6694) );
  OAI22_X1 U8385 ( .A1(n6703), .A2(n8917), .B1(n8928), .B2(n6694), .ZN(n6701)
         );
  OAI21_X1 U8386 ( .B1(n10178), .B2(n8597), .A(n6695), .ZN(n6698) );
  NAND2_X1 U8387 ( .A1(n10178), .A2(n6696), .ZN(n6697) );
  NAND2_X1 U8388 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n6699) );
  OAI21_X1 U8389 ( .B1(n7967), .B2(n4574), .A(n6699), .ZN(n6700) );
  AOI21_X1 U8390 ( .B1(n6701), .B2(n5122), .A(n6700), .ZN(n6710) );
  NAND2_X1 U8391 ( .A1(n6703), .A2(n6702), .ZN(n6706) );
  NAND2_X1 U8392 ( .A1(n6705), .A2(n6704), .ZN(n8932) );
  OAI211_X1 U8393 ( .C1(n6707), .C2(n8928), .A(n6706), .B(n8932), .ZN(n6708)
         );
  AOI22_X1 U8394 ( .A1(n6722), .A2(n6711), .B1(n4410), .B2(n6715), .ZN(n6713)
         );
  NAND2_X1 U8395 ( .A1(n6712), .A2(n7616), .ZN(n6742) );
  XNOR2_X1 U8396 ( .A(n6713), .B(n4411), .ZN(n6717) );
  INV_X1 U8397 ( .A(n6246), .ZN(n6714) );
  AOI22_X1 U8398 ( .A1(n4432), .A2(n6711), .B1(n6756), .B2(n6715), .ZN(n6716)
         );
  NAND2_X1 U8399 ( .A1(n6717), .A2(n6716), .ZN(n7282) );
  OR2_X1 U8400 ( .A1(n6717), .A2(n6716), .ZN(n6718) );
  AND2_X1 U8401 ( .A1(n7282), .A2(n6718), .ZN(n7200) );
  NOR2_X1 U8402 ( .A1(n6719), .A2(n7161), .ZN(n6720) );
  INV_X1 U8403 ( .A(n6721), .ZN(n6723) );
  NAND2_X1 U8404 ( .A1(n6723), .A2(n6722), .ZN(n6725) );
  AOI22_X1 U8405 ( .A1(n6743), .A2(n7666), .B1(P1_REG1_REG_0__SCAN_IN), .B2(
        n6953), .ZN(n6724) );
  NAND2_X1 U8406 ( .A1(n6725), .A2(n6724), .ZN(n6960) );
  INV_X1 U8407 ( .A(n6960), .ZN(n6726) );
  NAND2_X1 U8408 ( .A1(n6726), .A2(n4411), .ZN(n6727) );
  AND2_X1 U8409 ( .A1(n6959), .A2(n6727), .ZN(n6731) );
  OAI22_X1 U8410 ( .A1(n7765), .A2(n6753), .B1(n10078), .B2(n6748), .ZN(n6728)
         );
  XNOR2_X1 U8411 ( .A(n6728), .B(n4411), .ZN(n6732) );
  NAND2_X1 U8412 ( .A1(n6731), .A2(n6732), .ZN(n7121) );
  AOI22_X1 U8413 ( .A1(n6729), .A2(n4432), .B1(n6756), .B2(n6730), .ZN(n7123)
         );
  NAND2_X1 U8414 ( .A1(n7121), .A2(n7123), .ZN(n6735) );
  INV_X1 U8415 ( .A(n6731), .ZN(n6734) );
  INV_X1 U8416 ( .A(n6732), .ZN(n6733) );
  NAND2_X1 U8417 ( .A1(n6734), .A2(n6733), .ZN(n7122) );
  NAND2_X1 U8418 ( .A1(n6735), .A2(n7122), .ZN(n7199) );
  NAND2_X1 U8419 ( .A1(n7200), .A2(n7199), .ZN(n7198) );
  NAND2_X1 U8420 ( .A1(n7198), .A2(n7282), .ZN(n6740) );
  OAI22_X1 U8421 ( .A1(n7721), .A2(n4413), .B1(n10096), .B2(n6748), .ZN(n6736)
         );
  XNOR2_X1 U8422 ( .A(n4411), .B(n6736), .ZN(n6738) );
  OAI22_X1 U8423 ( .A1(n6913), .A2(n7721), .B1(n4413), .B2(n10096), .ZN(n6737)
         );
  NAND2_X1 U8424 ( .A1(n6738), .A2(n6737), .ZN(n6739) );
  AOI22_X1 U8425 ( .A1(n6756), .A2(n9444), .B1(n4410), .B2(n7724), .ZN(n6744)
         );
  XNOR2_X1 U8426 ( .A(n4411), .B(n6744), .ZN(n6747) );
  OAI22_X1 U8427 ( .A1(n6913), .A2(n10042), .B1(n4413), .B2(n9364), .ZN(n6745)
         );
  INV_X1 U8428 ( .A(n6745), .ZN(n6746) );
  XNOR2_X1 U8429 ( .A(n4414), .B(n6749), .ZN(n6758) );
  OAI22_X1 U8430 ( .A1(n6913), .A2(n10043), .B1(n4413), .B2(n7632), .ZN(n6757)
         );
  OR2_X1 U8431 ( .A1(n6758), .A2(n6757), .ZN(n7535) );
  OAI22_X1 U8432 ( .A1(n7542), .A2(n4413), .B1(n5032), .B2(n6748), .ZN(n6750)
         );
  XNOR2_X1 U8433 ( .A(n4414), .B(n6750), .ZN(n7483) );
  OAI22_X1 U8434 ( .A1(n6913), .A2(n7542), .B1(n4413), .B2(n5032), .ZN(n7486)
         );
  OR2_X1 U8435 ( .A1(n7483), .A2(n7486), .ZN(n6751) );
  NAND2_X1 U8436 ( .A1(n7483), .A2(n7486), .ZN(n7472) );
  NAND2_X1 U8437 ( .A1(n10162), .A2(n4410), .ZN(n6752) );
  OAI21_X1 U8438 ( .B1(n6754), .B2(n4413), .A(n6752), .ZN(n6755) );
  XNOR2_X1 U8439 ( .A(n6901), .B(n6755), .ZN(n6761) );
  AOI22_X1 U8440 ( .A1(n9442), .A2(n4432), .B1(n6756), .B2(n10162), .ZN(n6762)
         );
  XNOR2_X1 U8441 ( .A(n6761), .B(n6762), .ZN(n7476) );
  NAND2_X1 U8442 ( .A1(n6758), .A2(n6757), .ZN(n7534) );
  OAI211_X1 U8443 ( .C1(n7471), .C2(n7472), .A(n7476), .B(n7534), .ZN(n6759)
         );
  INV_X1 U8444 ( .A(n6759), .ZN(n6760) );
  INV_X1 U8445 ( .A(n6761), .ZN(n6763) );
  NAND2_X1 U8446 ( .A1(n6763), .A2(n6762), .ZN(n6764) );
  NAND2_X1 U8447 ( .A1(n5975), .A2(n6910), .ZN(n6766) );
  NAND2_X1 U8448 ( .A1(n10158), .A2(n4432), .ZN(n6765) );
  NAND2_X1 U8449 ( .A1(n6766), .A2(n6765), .ZN(n6774) );
  NAND2_X1 U8450 ( .A1(n5975), .A2(n4410), .ZN(n6768) );
  OR2_X1 U8451 ( .A1(n10139), .A2(n4413), .ZN(n6767) );
  NAND2_X1 U8452 ( .A1(n6768), .A2(n6767), .ZN(n6769) );
  XNOR2_X1 U8453 ( .A(n6769), .B(n4414), .ZN(n7796) );
  NAND2_X1 U8454 ( .A1(n10144), .A2(n4410), .ZN(n6770) );
  OAI21_X1 U8455 ( .B1(n9730), .B2(n4413), .A(n6770), .ZN(n6771) );
  XNOR2_X1 U8456 ( .A(n6771), .B(n4414), .ZN(n7798) );
  NAND2_X1 U8457 ( .A1(n10144), .A2(n6756), .ZN(n6772) );
  OAI21_X1 U8458 ( .B1(n6913), .B2(n9730), .A(n6772), .ZN(n7797) );
  INV_X1 U8459 ( .A(n7796), .ZN(n7854) );
  INV_X1 U8460 ( .A(n6774), .ZN(n7794) );
  NAND3_X1 U8461 ( .A1(n7854), .A2(n7794), .A3(n6775), .ZN(n6777) );
  OR2_X1 U8462 ( .A1(n7798), .A2(n7797), .ZN(n6776) );
  AND2_X1 U8463 ( .A1(n6777), .A2(n6776), .ZN(n6778) );
  NAND2_X1 U8464 ( .A1(n6782), .A2(n4410), .ZN(n6780) );
  OR2_X1 U8465 ( .A1(n10140), .A2(n4413), .ZN(n6779) );
  NAND2_X1 U8466 ( .A1(n6780), .A2(n6779), .ZN(n6781) );
  XNOR2_X1 U8467 ( .A(n6781), .B(n6901), .ZN(n6783) );
  AOI22_X1 U8468 ( .A1(n6782), .A2(n6910), .B1(n4432), .B2(n9441), .ZN(n6784)
         );
  XNOR2_X1 U8469 ( .A(n6783), .B(n6784), .ZN(n7692) );
  INV_X1 U8470 ( .A(n6783), .ZN(n6785) );
  NAND2_X1 U8471 ( .A1(n9888), .A2(n4410), .ZN(n6787) );
  OR2_X1 U8472 ( .A1(n9876), .A2(n4413), .ZN(n6786) );
  NAND2_X1 U8473 ( .A1(n6787), .A2(n6786), .ZN(n6788) );
  XNOR2_X1 U8474 ( .A(n6788), .B(n6901), .ZN(n6790) );
  NOR2_X1 U8475 ( .A1(n6913), .A2(n9876), .ZN(n6789) );
  AOI21_X1 U8476 ( .B1(n9888), .B2(n6910), .A(n6789), .ZN(n6791) );
  XNOR2_X1 U8477 ( .A(n6790), .B(n6791), .ZN(n7956) );
  INV_X1 U8478 ( .A(n6791), .ZN(n6792) );
  NAND2_X1 U8479 ( .A1(n6790), .A2(n6792), .ZN(n6793) );
  NAND2_X1 U8480 ( .A1(n7955), .A2(n6793), .ZN(n8249) );
  NAND2_X1 U8481 ( .A1(n9880), .A2(n4410), .ZN(n6795) );
  OR2_X1 U8482 ( .A1(n9884), .A2(n4413), .ZN(n6794) );
  NAND2_X1 U8483 ( .A1(n6795), .A2(n6794), .ZN(n6796) );
  XNOR2_X1 U8484 ( .A(n6796), .B(n6916), .ZN(n6808) );
  NOR2_X1 U8485 ( .A1(n6913), .A2(n9884), .ZN(n6797) );
  AOI21_X1 U8486 ( .B1(n9880), .B2(n6910), .A(n6797), .ZN(n6807) );
  XNOR2_X1 U8487 ( .A(n6808), .B(n6807), .ZN(n8250) );
  NAND2_X1 U8488 ( .A1(n9872), .A2(n4410), .ZN(n6799) );
  OR2_X1 U8489 ( .A1(n9877), .A2(n4413), .ZN(n6798) );
  NAND2_X1 U8490 ( .A1(n6799), .A2(n6798), .ZN(n6800) );
  XNOR2_X1 U8491 ( .A(n6800), .B(n6916), .ZN(n8238) );
  INV_X1 U8492 ( .A(n8238), .ZN(n6803) );
  NOR2_X1 U8493 ( .A1(n6913), .A2(n9877), .ZN(n6801) );
  AOI21_X1 U8494 ( .B1(n9872), .B2(n6910), .A(n6801), .ZN(n8237) );
  INV_X1 U8495 ( .A(n8237), .ZN(n6802) );
  OR2_X1 U8496 ( .A1(n8250), .A2(n5048), .ZN(n6814) );
  NAND2_X1 U8497 ( .A1(n9864), .A2(n4410), .ZN(n6805) );
  OR2_X1 U8498 ( .A1(n9868), .A2(n4413), .ZN(n6804) );
  NAND2_X1 U8499 ( .A1(n6805), .A2(n6804), .ZN(n6806) );
  XNOR2_X1 U8500 ( .A(n6806), .B(n6901), .ZN(n6818) );
  NAND2_X1 U8501 ( .A1(n6816), .A2(n4445), .ZN(n9287) );
  NAND2_X1 U8502 ( .A1(n8238), .A2(n8237), .ZN(n6809) );
  NAND2_X1 U8503 ( .A1(n6808), .A2(n6807), .ZN(n8236) );
  AND2_X1 U8504 ( .A1(n6809), .A2(n8236), .ZN(n6810) );
  OR2_X1 U8505 ( .A1(n5048), .A2(n6810), .ZN(n6817) );
  OR2_X1 U8506 ( .A1(n6818), .A2(n6817), .ZN(n9286) );
  NAND2_X1 U8507 ( .A1(n9864), .A2(n6910), .ZN(n6812) );
  NAND2_X1 U8508 ( .A1(n9438), .A2(n4432), .ZN(n6811) );
  NAND2_X1 U8509 ( .A1(n6812), .A2(n6811), .ZN(n9291) );
  AND2_X1 U8510 ( .A1(n9286), .A2(n9291), .ZN(n6813) );
  NAND2_X1 U8511 ( .A1(n9287), .A2(n6813), .ZN(n6821) );
  INV_X1 U8512 ( .A(n6814), .ZN(n6815) );
  NAND2_X1 U8513 ( .A1(n6816), .A2(n6815), .ZN(n6820) );
  AND2_X1 U8514 ( .A1(n6818), .A2(n6817), .ZN(n6819) );
  NAND2_X1 U8515 ( .A1(n9689), .A2(n4410), .ZN(n6823) );
  NAND2_X1 U8516 ( .A1(n9676), .A2(n6910), .ZN(n6822) );
  NAND2_X1 U8517 ( .A1(n6823), .A2(n6822), .ZN(n6824) );
  XNOR2_X1 U8518 ( .A(n6824), .B(n6916), .ZN(n9332) );
  NOR2_X1 U8519 ( .A1(n9843), .A2(n6913), .ZN(n6825) );
  AOI21_X1 U8520 ( .B1(n9689), .B2(n6910), .A(n6825), .ZN(n9331) );
  NAND2_X1 U8521 ( .A1(n9856), .A2(n6910), .ZN(n6827) );
  NAND2_X1 U8522 ( .A1(n4432), .A2(n9696), .ZN(n6826) );
  NAND2_X1 U8523 ( .A1(n9856), .A2(n4410), .ZN(n6829) );
  NAND2_X1 U8524 ( .A1(n9696), .A2(n6910), .ZN(n6828) );
  NAND2_X1 U8525 ( .A1(n6829), .A2(n6828), .ZN(n6830) );
  XNOR2_X1 U8526 ( .A(n6830), .B(n6916), .ZN(n6834) );
  OAI22_X1 U8527 ( .A1(n9332), .A2(n9331), .B1(n9422), .B2(n6834), .ZN(n6831)
         );
  INV_X1 U8528 ( .A(n6834), .ZN(n9330) );
  INV_X1 U8529 ( .A(n9422), .ZN(n6832) );
  INV_X1 U8530 ( .A(n9331), .ZN(n6833) );
  OAI21_X1 U8531 ( .B1(n9330), .B2(n6832), .A(n6833), .ZN(n6836) );
  NOR2_X1 U8532 ( .A1(n6833), .A2(n6832), .ZN(n6835) );
  AOI22_X1 U8533 ( .A1(n9332), .A2(n6836), .B1(n6835), .B2(n6834), .ZN(n6837)
         );
  NAND2_X1 U8534 ( .A1(n9847), .A2(n4410), .ZN(n6839) );
  OR2_X1 U8535 ( .A1(n9834), .A2(n4413), .ZN(n6838) );
  NAND2_X1 U8536 ( .A1(n6839), .A2(n6838), .ZN(n6840) );
  XNOR2_X1 U8537 ( .A(n6840), .B(n6916), .ZN(n9341) );
  NOR2_X1 U8538 ( .A1(n9834), .A2(n6913), .ZN(n6841) );
  AOI21_X1 U8539 ( .B1(n9847), .B2(n6910), .A(n6841), .ZN(n9340) );
  AND2_X1 U8540 ( .A1(n9341), .A2(n9340), .ZN(n6843) );
  NAND2_X1 U8541 ( .A1(n9662), .A2(n6910), .ZN(n6845) );
  NAND2_X1 U8542 ( .A1(n9437), .A2(n4432), .ZN(n6844) );
  NAND2_X1 U8543 ( .A1(n6845), .A2(n6844), .ZN(n9393) );
  NAND2_X1 U8544 ( .A1(n9662), .A2(n4410), .ZN(n6847) );
  NAND2_X1 U8545 ( .A1(n9437), .A2(n6910), .ZN(n6846) );
  NAND2_X1 U8546 ( .A1(n6847), .A2(n6846), .ZN(n6848) );
  XNOR2_X1 U8547 ( .A(n6848), .B(n6901), .ZN(n9394) );
  NAND2_X1 U8548 ( .A1(n6853), .A2(n4410), .ZN(n6850) );
  NAND2_X1 U8549 ( .A1(n9436), .A2(n6910), .ZN(n6849) );
  NAND2_X1 U8550 ( .A1(n6850), .A2(n6849), .ZN(n6851) );
  XNOR2_X1 U8551 ( .A(n6851), .B(n6916), .ZN(n6855) );
  NOR2_X1 U8552 ( .A1(n9835), .A2(n6913), .ZN(n6852) );
  AOI21_X1 U8553 ( .B1(n6853), .B2(n6910), .A(n6852), .ZN(n6854) );
  NAND2_X1 U8554 ( .A1(n6855), .A2(n6854), .ZN(n6857) );
  OR2_X1 U8555 ( .A1(n6855), .A2(n6854), .ZN(n6856) );
  NAND2_X1 U8556 ( .A1(n6857), .A2(n6856), .ZN(n9312) );
  OAI22_X1 U8557 ( .A1(n6859), .A2(n6748), .B1(n9813), .B2(n4413), .ZN(n6858)
         );
  XNOR2_X1 U8558 ( .A(n6858), .B(n6916), .ZN(n6862) );
  OR2_X1 U8559 ( .A1(n6859), .A2(n4413), .ZN(n6861) );
  NAND2_X1 U8560 ( .A1(n9614), .A2(n4432), .ZN(n6860) );
  AND2_X1 U8561 ( .A1(n6861), .A2(n6860), .ZN(n6863) );
  INV_X1 U8562 ( .A(n6862), .ZN(n6865) );
  INV_X1 U8563 ( .A(n6863), .ZN(n6864) );
  NAND2_X1 U8564 ( .A1(n6865), .A2(n6864), .ZN(n9371) );
  NAND2_X1 U8565 ( .A1(n6866), .A2(n9371), .ZN(n9321) );
  NAND2_X1 U8566 ( .A1(n9817), .A2(n4410), .ZN(n6868) );
  NAND2_X1 U8567 ( .A1(n9803), .A2(n6910), .ZN(n6867) );
  NAND2_X1 U8568 ( .A1(n6868), .A2(n6867), .ZN(n6869) );
  XNOR2_X1 U8569 ( .A(n6869), .B(n6901), .ZN(n6873) );
  NAND2_X1 U8570 ( .A1(n9817), .A2(n6910), .ZN(n6871) );
  NAND2_X1 U8571 ( .A1(n9803), .A2(n4432), .ZN(n6870) );
  NAND2_X1 U8572 ( .A1(n6871), .A2(n6870), .ZN(n6874) );
  AND2_X1 U8573 ( .A1(n6873), .A2(n6874), .ZN(n9319) );
  OAI22_X1 U8574 ( .A1(n9807), .A2(n4413), .B1(n9814), .B2(n6913), .ZN(n9379)
         );
  OR2_X1 U8575 ( .A1(n9319), .A2(n9379), .ZN(n6872) );
  INV_X1 U8576 ( .A(n6872), .ZN(n6877) );
  INV_X1 U8577 ( .A(n6873), .ZN(n6876) );
  INV_X1 U8578 ( .A(n6874), .ZN(n6875) );
  NAND2_X1 U8579 ( .A1(n6876), .A2(n6875), .ZN(n9318) );
  OAI22_X1 U8580 ( .A1(n9807), .A2(n6748), .B1(n9814), .B2(n4413), .ZN(n6878)
         );
  XNOR2_X1 U8581 ( .A(n6878), .B(n6901), .ZN(n9380) );
  INV_X1 U8582 ( .A(n9319), .ZN(n6880) );
  OAI22_X1 U8583 ( .A1(n9585), .A2(n4413), .B1(n9791), .B2(n6913), .ZN(n8380)
         );
  NAND2_X1 U8584 ( .A1(n6260), .A2(n4410), .ZN(n6882) );
  NAND2_X1 U8585 ( .A1(n9804), .A2(n6910), .ZN(n6881) );
  NAND2_X1 U8586 ( .A1(n6882), .A2(n6881), .ZN(n6883) );
  XNOR2_X1 U8587 ( .A(n6883), .B(n6901), .ZN(n8381) );
  NAND2_X1 U8588 ( .A1(n9795), .A2(n4410), .ZN(n6885) );
  NAND2_X1 U8589 ( .A1(n9782), .A2(n6910), .ZN(n6884) );
  NAND2_X1 U8590 ( .A1(n6885), .A2(n6884), .ZN(n6886) );
  XNOR2_X1 U8591 ( .A(n6886), .B(n6916), .ZN(n6889) );
  NOR2_X1 U8592 ( .A1(n9547), .A2(n6913), .ZN(n6887) );
  AOI21_X1 U8593 ( .B1(n9795), .B2(n6910), .A(n6887), .ZN(n6888) );
  NOR2_X1 U8594 ( .A1(n6889), .A2(n6888), .ZN(n8383) );
  AOI21_X1 U8595 ( .B1(n8380), .B2(n8381), .A(n8383), .ZN(n6890) );
  NAND2_X1 U8596 ( .A1(n9545), .A2(n4410), .ZN(n6892) );
  OR2_X1 U8597 ( .A1(n9792), .A2(n4413), .ZN(n6891) );
  NAND2_X1 U8598 ( .A1(n6892), .A2(n6891), .ZN(n6893) );
  XNOR2_X1 U8599 ( .A(n6893), .B(n6916), .ZN(n6897) );
  NOR2_X1 U8600 ( .A1(n9792), .A2(n6913), .ZN(n6894) );
  AOI21_X1 U8601 ( .B1(n9545), .B2(n6756), .A(n6894), .ZN(n6896) );
  XNOR2_X1 U8602 ( .A(n6897), .B(n6896), .ZN(n8384) );
  NOR2_X1 U8603 ( .A1(n6895), .A2(n8384), .ZN(n9406) );
  AND2_X1 U8604 ( .A1(n6897), .A2(n6896), .ZN(n9405) );
  NOR2_X1 U8605 ( .A1(n9548), .A2(n6913), .ZN(n6898) );
  AOI21_X1 U8606 ( .B1(n9776), .B2(n6910), .A(n6898), .ZN(n6903) );
  NAND2_X1 U8607 ( .A1(n9776), .A2(n4410), .ZN(n6900) );
  NAND2_X1 U8608 ( .A1(n9783), .A2(n6910), .ZN(n6899) );
  NAND2_X1 U8609 ( .A1(n6900), .A2(n6899), .ZN(n6902) );
  XNOR2_X1 U8610 ( .A(n6902), .B(n6901), .ZN(n6905) );
  XOR2_X1 U8611 ( .A(n6903), .B(n6905), .Z(n9404) );
  INV_X1 U8612 ( .A(n6903), .ZN(n6904) );
  NAND2_X1 U8613 ( .A1(n8350), .A2(n4410), .ZN(n6907) );
  NAND2_X1 U8614 ( .A1(n6276), .A2(n6910), .ZN(n6906) );
  NAND2_X1 U8615 ( .A1(n6907), .A2(n6906), .ZN(n6908) );
  XNOR2_X1 U8616 ( .A(n6908), .B(n6916), .ZN(n6912) );
  NOR2_X1 U8617 ( .A1(n9413), .A2(n6913), .ZN(n6909) );
  AOI21_X1 U8618 ( .B1(n8350), .B2(n6910), .A(n6909), .ZN(n6911) );
  NAND2_X1 U8619 ( .A1(n6912), .A2(n6911), .ZN(n6937) );
  OAI21_X1 U8620 ( .B1(n6912), .B2(n6911), .A(n6937), .ZN(n6942) );
  NAND2_X1 U8621 ( .A1(n9515), .A2(n6910), .ZN(n6915) );
  OR2_X1 U8622 ( .A1(n9520), .A2(n6913), .ZN(n6914) );
  NAND2_X1 U8623 ( .A1(n6915), .A2(n6914), .ZN(n6917) );
  XNOR2_X1 U8624 ( .A(n6917), .B(n6916), .ZN(n6920) );
  NAND2_X1 U8625 ( .A1(n9515), .A2(n4410), .ZN(n6918) );
  OAI21_X1 U8626 ( .B1(n9520), .B2(n4413), .A(n6918), .ZN(n6919) );
  XNOR2_X1 U8627 ( .A(n6920), .B(n6919), .ZN(n6923) );
  INV_X1 U8628 ( .A(n6923), .ZN(n6938) );
  AND2_X1 U8629 ( .A1(n7088), .A2(n7614), .ZN(n6921) );
  INV_X1 U8630 ( .A(n7609), .ZN(n6996) );
  NAND3_X1 U8631 ( .A1(n6938), .A2(n9408), .A3(n6937), .ZN(n6922) );
  NOR2_X1 U8632 ( .A1(n7628), .A2(n6279), .ZN(n10050) );
  INV_X1 U8633 ( .A(n6927), .ZN(n6929) );
  NAND2_X1 U8634 ( .A1(n10050), .A2(n6929), .ZN(n6924) );
  AND2_X1 U8635 ( .A1(n7614), .A2(n6925), .ZN(n6926) );
  NAND3_X1 U8636 ( .A1(n6928), .A2(n6927), .A3(n6926), .ZN(n7543) );
  INV_X1 U8637 ( .A(n4412), .ZN(n7159) );
  NAND2_X1 U8638 ( .A1(n9760), .A2(n9386), .ZN(n6936) );
  OAI21_X1 U8639 ( .B1(n10050), .B2(n10130), .A(n6929), .ZN(n6931) );
  NAND2_X1 U8640 ( .A1(n6931), .A2(n6930), .ZN(n7098) );
  INV_X1 U8641 ( .A(n6932), .ZN(n6933) );
  OR2_X1 U8642 ( .A1(n7098), .A2(n6933), .ZN(n6934) );
  AOI22_X1 U8643 ( .A1(n8405), .A2(n9410), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6935) );
  OAI211_X1 U8644 ( .C1(n9413), .C2(n9384), .A(n6936), .B(n6935), .ZN(n6940)
         );
  NOR3_X1 U8645 ( .A1(n6938), .A2(n9432), .A3(n6937), .ZN(n6939) );
  AOI211_X1 U8646 ( .C1(n6949), .C2(n9515), .A(n6940), .B(n6939), .ZN(n6941)
         );
  OAI21_X1 U8647 ( .B1(n9403), .B2(n6943), .A(n6942), .ZN(n6944) );
  INV_X1 U8648 ( .A(n6944), .ZN(n6945) );
  OAI21_X1 U8649 ( .B1(n6946), .B2(n6945), .A(n9408), .ZN(n6952) );
  INV_X1 U8650 ( .A(n9520), .ZN(n9514) );
  NOR2_X1 U8651 ( .A1(n9548), .A2(n9384), .ZN(n6948) );
  OAI22_X1 U8652 ( .A1(n8348), .A2(n9429), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10569), .ZN(n6947) );
  AOI211_X1 U8653 ( .C1(n9514), .C2(n9386), .A(n6948), .B(n6947), .ZN(n6951)
         );
  NAND2_X1 U8654 ( .A1(n8350), .A2(n6949), .ZN(n6950) );
  NAND3_X1 U8655 ( .A1(n6952), .A2(n6951), .A3(n6950), .ZN(P1_U3212) );
  NAND2_X1 U8656 ( .A1(n6954), .A2(n6953), .ZN(n6963) );
  OR2_X2 U8657 ( .A1(n6963), .A2(P1_U3084), .ZN(n9445) );
  INV_X1 U8658 ( .A(n6954), .ZN(n6955) );
  OR2_X1 U8659 ( .A1(n7088), .A2(n6955), .ZN(n6956) );
  NAND2_X1 U8660 ( .A1(n6956), .A2(n6963), .ZN(n6967) );
  OAI21_X1 U8661 ( .B1(n6967), .B2(n6957), .A(P1_STATE_REG_SCAN_IN), .ZN(
        P1_U3083) );
  AND2_X1 U8662 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n6975) );
  INV_X1 U8663 ( .A(n6975), .ZN(n7152) );
  OAI21_X1 U8664 ( .B1(n6958), .B2(n6960), .A(n6959), .ZN(n7099) );
  MUX2_X1 U8665 ( .A(n7152), .B(n7099), .S(n9504), .Z(n6962) );
  OAI21_X1 U8666 ( .B1(n9504), .B2(P1_REG2_REG_0__SCAN_IN), .A(n7159), .ZN(
        n7162) );
  AOI21_X1 U8667 ( .B1(n7161), .B2(n7162), .A(n9445), .ZN(n6961) );
  OAI21_X1 U8668 ( .B1(n6962), .B2(n4412), .A(n6961), .ZN(n7181) );
  INV_X1 U8669 ( .A(n7181), .ZN(n6987) );
  INV_X1 U8670 ( .A(n6963), .ZN(n6964) );
  INV_X1 U8671 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6965) );
  NOR2_X1 U8672 ( .A1(n10026), .A2(n6965), .ZN(n6986) );
  INV_X1 U8673 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6972) );
  INV_X1 U8674 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10152) );
  MUX2_X1 U8675 ( .A(n10152), .B(P1_REG1_REG_2__SCAN_IN), .S(n7057), .Z(n6970)
         );
  INV_X1 U8676 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10150) );
  MUX2_X1 U8677 ( .A(n10150), .B(P1_REG1_REG_1__SCAN_IN), .S(n8364), .Z(n7148)
         );
  AND2_X1 U8678 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n7147) );
  NAND2_X1 U8679 ( .A1(n7148), .A2(n7147), .ZN(n7146) );
  INV_X1 U8680 ( .A(n8364), .ZN(n6977) );
  NAND2_X1 U8681 ( .A1(n6977), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6966) );
  NAND2_X1 U8682 ( .A1(n7146), .A2(n6966), .ZN(n6969) );
  INV_X1 U8683 ( .A(n9504), .ZN(n6973) );
  NOR2_X1 U8684 ( .A1(n6973), .A2(n4412), .ZN(n6968) );
  NAND2_X1 U8685 ( .A1(n7160), .A2(n6968), .ZN(n10023) );
  NAND2_X1 U8686 ( .A1(n6969), .A2(n6970), .ZN(n7059) );
  OAI211_X1 U8687 ( .C1(n6970), .C2(n6969), .A(n10003), .B(n7059), .ZN(n6971)
         );
  OAI21_X1 U8688 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6972), .A(n6971), .ZN(n6985) );
  INV_X1 U8689 ( .A(n7225), .ZN(n7165) );
  INV_X1 U8690 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6974) );
  MUX2_X1 U8691 ( .A(n6974), .B(P1_REG2_REG_1__SCAN_IN), .S(n8364), .Z(n6976)
         );
  NAND2_X1 U8692 ( .A1(n6976), .A2(n6975), .ZN(n7155) );
  NAND2_X1 U8693 ( .A1(n6977), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6981) );
  NAND2_X1 U8694 ( .A1(n7155), .A2(n6981), .ZN(n6979) );
  INV_X1 U8695 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7776) );
  MUX2_X1 U8696 ( .A(n7776), .B(P1_REG2_REG_2__SCAN_IN), .S(n7057), .Z(n6978)
         );
  NAND2_X1 U8697 ( .A1(n6979), .A2(n6978), .ZN(n7138) );
  MUX2_X1 U8698 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n7776), .S(n7057), .Z(n6980)
         );
  NAND3_X1 U8699 ( .A1(n7155), .A2(n6981), .A3(n6980), .ZN(n6982) );
  NAND3_X1 U8700 ( .A1(n10013), .A2(n7138), .A3(n6982), .ZN(n6983) );
  OAI21_X1 U8701 ( .B1(n10017), .B2(n7057), .A(n6983), .ZN(n6984) );
  OR4_X1 U8702 ( .A1(n6987), .A2(n6986), .A3(n6985), .A4(n6984), .ZN(P1_U3243)
         );
  NAND2_X1 U8703 ( .A1(n6998), .A2(P1_U3084), .ZN(n9921) );
  OAI222_X1 U8704 ( .A1(P1_U3084), .A2(n7057), .B1(n9921), .B2(n7000), .C1(
        n6988), .C2(n4405), .ZN(P1_U3351) );
  INV_X1 U8705 ( .A(n6989), .ZN(n7007) );
  OAI222_X1 U8706 ( .A1(n4405), .A2(n6990), .B1(n9921), .B2(n7007), .C1(
        P1_U3084), .C2(n7172), .ZN(P1_U3349) );
  OAI222_X1 U8707 ( .A1(P1_U3084), .A2(n9446), .B1(n9921), .B2(n7009), .C1(
        n6991), .C2(n4405), .ZN(P1_U3348) );
  INV_X1 U8708 ( .A(n7109), .ZN(n7082) );
  INV_X1 U8709 ( .A(n6992), .ZN(n7002) );
  INV_X1 U8710 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6993) );
  OAI222_X1 U8711 ( .A1(P1_U3084), .A2(n7082), .B1(n9921), .B2(n7002), .C1(
        n6993), .C2(n4405), .ZN(P1_U3347) );
  INV_X1 U8712 ( .A(n6994), .ZN(n7003) );
  AOI22_X1 U8714 ( .A1(n7221), .A2(P1_STATE_REG_SCAN_IN), .B1(n10615), .B2(
        P2_DATAO_REG_9__SCAN_IN), .ZN(n6995) );
  OAI21_X1 U8715 ( .B1(n7003), .B2(n9921), .A(n6995), .ZN(P1_U3344) );
  NAND2_X1 U8716 ( .A1(n7614), .A2(n6996), .ZN(n6997) );
  OAI21_X1 U8717 ( .B1(n7614), .B2(n6305), .A(n6997), .ZN(P1_U3441) );
  AND2_X1 U8718 ( .A1(n6998), .A2(P2_U3152), .ZN(n9279) );
  NAND2_X1 U8719 ( .A1(n5291), .A2(P2_U3152), .ZN(n8366) );
  OAI222_X1 U8720 ( .A1(n8368), .A2(n5139), .B1(n9281), .B2(n7000), .C1(n6999), 
        .C2(P2_U3152), .ZN(P2_U3356) );
  OAI222_X1 U8721 ( .A1(n8368), .A2(n5262), .B1(n9281), .B2(n7002), .C1(n7001), 
        .C2(P2_U3152), .ZN(P2_U3352) );
  OAI222_X1 U8722 ( .A1(n8368), .A2(n7004), .B1(n9281), .B2(n7003), .C1(n7395), 
        .C2(P2_U3152), .ZN(P2_U3349) );
  OAI222_X1 U8723 ( .A1(n8368), .A2(n5177), .B1(n9281), .B2(n7012), .C1(n7005), 
        .C2(P2_U3152), .ZN(P2_U3355) );
  OAI222_X1 U8724 ( .A1(n8368), .A2(n7008), .B1(n9281), .B2(n7007), .C1(
        P2_U3152), .C2(n7006), .ZN(P2_U3354) );
  INV_X1 U8725 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7010) );
  OAI222_X1 U8726 ( .A1(n8368), .A2(n7010), .B1(n9281), .B2(n7009), .C1(n7381), 
        .C2(P2_U3152), .ZN(P2_U3353) );
  INV_X1 U8727 ( .A(n9921), .ZN(n8013) );
  OAI222_X1 U8728 ( .A1(P1_U3084), .A2(n7143), .B1(n9923), .B2(n7012), .C1(
        n7011), .C2(n4405), .ZN(P1_U3350) );
  INV_X1 U8729 ( .A(n7013), .ZN(n7024) );
  AOI22_X1 U8730 ( .A1(n9469), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10615), .ZN(n7014) );
  OAI21_X1 U8731 ( .B1(n7024), .B2(n9923), .A(n7014), .ZN(P1_U3343) );
  INV_X1 U8732 ( .A(n7015), .ZN(n7017) );
  OAI222_X1 U8733 ( .A1(n8368), .A2(n5292), .B1(n9281), .B2(n7017), .C1(
        P2_U3152), .C2(n7016), .ZN(P2_U3351) );
  INV_X1 U8734 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n7018) );
  INV_X1 U8735 ( .A(n7112), .ZN(n7212) );
  OAI222_X1 U8736 ( .A1(n4405), .A2(n7018), .B1(n9923), .B2(n7017), .C1(
        P1_U3084), .C2(n7212), .ZN(P1_U3346) );
  NAND2_X1 U8737 ( .A1(n4406), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n7022) );
  NAND2_X1 U8738 ( .A1(n7019), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n7021) );
  NAND2_X1 U8739 ( .A1(n7047), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n7020) );
  AND3_X1 U8740 ( .A1(n7022), .A2(n7021), .A3(n7020), .ZN(n8563) );
  NAND2_X1 U8741 ( .A1(n8773), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n7023) );
  OAI21_X1 U8742 ( .B1(n8773), .B2(n8563), .A(n7023), .ZN(P2_U3582) );
  OAI222_X1 U8743 ( .A1(n8368), .A2(n7025), .B1(n9281), .B2(n7024), .C1(n7384), 
        .C2(P2_U3152), .ZN(P2_U3348) );
  INV_X1 U8744 ( .A(n7026), .ZN(n7032) );
  AOI22_X1 U8745 ( .A1(n7234), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10615), .ZN(n7027) );
  OAI21_X1 U8746 ( .B1(n7032), .B2(n9921), .A(n7027), .ZN(P1_U3342) );
  INV_X1 U8747 ( .A(n7028), .ZN(n7030) );
  OAI222_X1 U8748 ( .A1(n8368), .A2(n5317), .B1(n9281), .B2(n7030), .C1(
        P2_U3152), .C2(n7029), .ZN(P2_U3350) );
  INV_X1 U8749 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n7031) );
  INV_X1 U8750 ( .A(n7190), .ZN(n7106) );
  OAI222_X1 U8751 ( .A1(n4405), .A2(n7031), .B1(n9921), .B2(n7030), .C1(
        P1_U3084), .C2(n7106), .ZN(P1_U3345) );
  INV_X1 U8752 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n7033) );
  OAI222_X1 U8753 ( .A1(n8368), .A2(n7033), .B1(n9281), .B2(n7032), .C1(n7320), 
        .C2(P2_U3152), .ZN(P2_U3347) );
  NAND2_X1 U8754 ( .A1(n6723), .A2(P1_U4006), .ZN(n7035) );
  OAI21_X1 U8755 ( .B1(P1_U4006), .B2(n5106), .A(n7035), .ZN(P1_U3555) );
  INV_X1 U8756 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n10398) );
  NAND2_X1 U8757 ( .A1(n9505), .A2(P1_U4006), .ZN(n7036) );
  OAI21_X1 U8758 ( .B1(P1_U4006), .B2(n10398), .A(n7036), .ZN(P1_U3586) );
  INV_X1 U8759 ( .A(n7037), .ZN(n7038) );
  INV_X1 U8760 ( .A(n10073), .ZN(n10074) );
  NOR2_X1 U8761 ( .A1(n10074), .A2(P1_D_REG_0__SCAN_IN), .ZN(n7041) );
  OAI22_X1 U8762 ( .A1(n7041), .A2(n7040), .B1(n7614), .B2(n7039), .ZN(
        P1_U3440) );
  INV_X1 U8763 ( .A(n7042), .ZN(n7044) );
  INV_X1 U8764 ( .A(n7451), .ZN(n7043) );
  OAI222_X1 U8765 ( .A1(n4405), .A2(n10446), .B1(n9921), .B2(n7044), .C1(
        P1_U3084), .C2(n7043), .ZN(P1_U3341) );
  OAI222_X1 U8766 ( .A1(n8368), .A2(n7045), .B1(n9281), .B2(n7044), .C1(
        P2_U3152), .C2(n7424), .ZN(P2_U3346) );
  NOR2_X1 U8767 ( .A1(P2_U3966), .A2(n8922), .ZN(P2_U3151) );
  NAND2_X1 U8768 ( .A1(P2_U3966), .A2(n8374), .ZN(n7046) );
  OAI21_X1 U8769 ( .B1(P2_U3966), .B2(n5105), .A(n7046), .ZN(P2_U3552) );
  INV_X1 U8770 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n10481) );
  NAND2_X1 U8771 ( .A1(n7047), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7051) );
  INV_X1 U8772 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7048) );
  OR2_X1 U8773 ( .A1(n7049), .A2(n7048), .ZN(n7050) );
  OAI211_X1 U8774 ( .C1(n7052), .C2(n10481), .A(n7051), .B(n7050), .ZN(n8561)
         );
  NAND2_X1 U8775 ( .A1(P2_U3966), .A2(n8561), .ZN(n7053) );
  OAI21_X1 U8776 ( .B1(P2_U3966), .B2(n9912), .A(n7053), .ZN(P2_U3583) );
  INV_X1 U8777 ( .A(n7054), .ZN(n7056) );
  OAI222_X1 U8778 ( .A1(n8368), .A2(n10316), .B1(n9281), .B2(n7056), .C1(n7055), .C2(P2_U3152), .ZN(P2_U3345) );
  INV_X1 U8779 ( .A(n7454), .ZN(n9974) );
  OAI222_X1 U8780 ( .A1(P1_U3084), .A2(n9974), .B1(n9923), .B2(n7056), .C1(
        n10514), .C2(n4405), .ZN(P1_U3340) );
  INV_X1 U8781 ( .A(n10026), .ZN(n9455) );
  INV_X1 U8782 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10433) );
  MUX2_X1 U8783 ( .A(n10433), .B(P1_REG1_REG_6__SCAN_IN), .S(n7109), .Z(n7068)
         );
  INV_X1 U8784 ( .A(n7057), .ZN(n7071) );
  NAND2_X1 U8785 ( .A1(n7071), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n7058) );
  NAND2_X1 U8786 ( .A1(n7059), .A2(n7058), .ZN(n7131) );
  XNOR2_X1 U8787 ( .A(n7143), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n7132) );
  INV_X1 U8788 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n7060) );
  OR2_X1 U8789 ( .A1(n7143), .A2(n7060), .ZN(n7061) );
  XNOR2_X1 U8790 ( .A(n7172), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n7174) );
  INV_X1 U8791 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n7062) );
  NAND2_X1 U8792 ( .A1(n7172), .A2(n7062), .ZN(n7063) );
  XNOR2_X1 U8793 ( .A(n9446), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n9458) );
  NAND2_X1 U8794 ( .A1(n9457), .A2(n9458), .ZN(n9456) );
  INV_X1 U8795 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7064) );
  OR2_X1 U8796 ( .A1(n9446), .A2(n7064), .ZN(n7065) );
  NAND2_X1 U8797 ( .A1(n9456), .A2(n7065), .ZN(n7067) );
  INV_X1 U8798 ( .A(n7103), .ZN(n7066) );
  AOI21_X1 U8799 ( .B1(n7068), .B2(n7067), .A(n7066), .ZN(n7069) );
  NAND2_X1 U8800 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7545) );
  OAI21_X1 U8801 ( .B1(n10023), .B2(n7069), .A(n7545), .ZN(n7070) );
  AOI21_X1 U8802 ( .B1(n9455), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n7070), .ZN(
        n7081) );
  NAND2_X1 U8803 ( .A1(n7071), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n7137) );
  NAND2_X1 U8804 ( .A1(n7138), .A2(n7137), .ZN(n7073) );
  INV_X1 U8805 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7984) );
  MUX2_X1 U8806 ( .A(n7984), .B(P1_REG2_REG_3__SCAN_IN), .S(n7143), .Z(n7072)
         );
  NAND2_X1 U8807 ( .A1(n7073), .A2(n7072), .ZN(n7140) );
  OR2_X1 U8808 ( .A1(n7143), .A2(n7984), .ZN(n7074) );
  AND2_X1 U8809 ( .A1(n7140), .A2(n7074), .ZN(n7170) );
  INV_X1 U8810 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n10464) );
  NAND2_X1 U8811 ( .A1(n7172), .A2(n10464), .ZN(n9448) );
  OAI21_X1 U8812 ( .B1(n7172), .B2(n10464), .A(n9448), .ZN(n7075) );
  INV_X1 U8813 ( .A(n7075), .ZN(n7171) );
  NAND2_X1 U8814 ( .A1(n7170), .A2(n7171), .ZN(n9450) );
  NAND2_X1 U8815 ( .A1(n9450), .A2(n9448), .ZN(n7076) );
  INV_X1 U8816 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10047) );
  MUX2_X1 U8817 ( .A(n10047), .B(P1_REG2_REG_5__SCAN_IN), .S(n9446), .Z(n9447)
         );
  NAND2_X1 U8818 ( .A1(n7076), .A2(n9447), .ZN(n9452) );
  NAND2_X1 U8819 ( .A1(n9446), .A2(n10047), .ZN(n7077) );
  AND2_X1 U8820 ( .A1(n9452), .A2(n7077), .ZN(n7079) );
  INV_X1 U8821 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7624) );
  MUX2_X1 U8822 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7624), .S(n7109), .Z(n7078)
         );
  NAND2_X1 U8823 ( .A1(n7079), .A2(n7078), .ZN(n7111) );
  OAI211_X1 U8824 ( .C1(n7079), .C2(n7078), .A(n10013), .B(n7111), .ZN(n7080)
         );
  OAI211_X1 U8825 ( .C1(n10017), .C2(n7082), .A(n7081), .B(n7080), .ZN(
        P1_U3247) );
  INV_X1 U8826 ( .A(n7829), .ZN(n7825) );
  INV_X1 U8827 ( .A(n7083), .ZN(n7084) );
  OAI222_X1 U8828 ( .A1(P1_U3084), .A2(n7825), .B1(n9923), .B2(n7084), .C1(
        n10437), .C2(n4405), .ZN(P1_U3339) );
  OAI222_X1 U8829 ( .A1(n8368), .A2(n7086), .B1(P2_U3152), .B2(n7085), .C1(
        n7084), .C2(n8366), .ZN(P2_U3344) );
  INV_X1 U8830 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n7158) );
  NAND2_X1 U8831 ( .A1(n7087), .A2(n10056), .ZN(n7089) );
  NAND3_X1 U8832 ( .A1(n7089), .A2(n7088), .A3(n7628), .ZN(n7091) );
  NAND2_X1 U8833 ( .A1(n10159), .A2(n6729), .ZN(n7090) );
  NAND2_X1 U8834 ( .A1(n7091), .A2(n7090), .ZN(n7669) );
  INV_X1 U8835 ( .A(n7669), .ZN(n7092) );
  OAI21_X1 U8836 ( .B1(n10049), .B2(n7628), .A(n7092), .ZN(n7094) );
  NAND2_X1 U8837 ( .A1(n7094), .A2(n10177), .ZN(n7093) );
  OAI21_X1 U8838 ( .B1(n10177), .B2(n7158), .A(n7093), .ZN(P1_U3523) );
  INV_X1 U8839 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n7096) );
  NAND2_X1 U8840 ( .A1(n7094), .A2(n10588), .ZN(n7095) );
  OAI21_X1 U8841 ( .B1(n10588), .B2(n7096), .A(n7095), .ZN(P1_U3454) );
  NOR2_X1 U8842 ( .A1(n7098), .A2(n7097), .ZN(n7205) );
  INV_X1 U8843 ( .A(n7205), .ZN(n7127) );
  AOI22_X1 U8844 ( .A1(n7127), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9408), .B2(
        n7099), .ZN(n7101) );
  AOI22_X1 U8845 ( .A1(n6949), .A2(n7666), .B1(n9386), .B2(n6729), .ZN(n7100)
         );
  NAND2_X1 U8846 ( .A1(n7101), .A2(n7100), .ZN(P1_U3230) );
  XNOR2_X1 U8847 ( .A(n7221), .B(P1_REG1_REG_9__SCAN_IN), .ZN(n7217) );
  INV_X1 U8848 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7107) );
  OR2_X1 U8849 ( .A1(n7109), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7102) );
  INV_X1 U8850 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7104) );
  XNOR2_X1 U8851 ( .A(n7112), .B(n7104), .ZN(n7206) );
  OR2_X1 U8852 ( .A1(n7112), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7105) );
  MUX2_X1 U8853 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n7107), .S(n7190), .Z(n7191)
         );
  AOI21_X1 U8854 ( .B1(n7107), .B2(n7106), .A(n7194), .ZN(n7218) );
  XOR2_X1 U8855 ( .A(n7217), .B(n7218), .Z(n7120) );
  AND2_X1 U8856 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7802) );
  INV_X1 U8857 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10602) );
  NOR2_X1 U8858 ( .A1(n10026), .A2(n10602), .ZN(n7108) );
  AOI211_X1 U8859 ( .C1(n10001), .C2(n7221), .A(n7802), .B(n7108), .ZN(n7119)
         );
  NAND2_X1 U8860 ( .A1(n7109), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n7110) );
  OR2_X1 U8861 ( .A1(n7112), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7184) );
  NAND2_X1 U8862 ( .A1(n7112), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n7113) );
  NAND2_X1 U8863 ( .A1(n7184), .A2(n7113), .ZN(n7211) );
  INV_X1 U8864 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7114) );
  MUX2_X1 U8865 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n7114), .S(n7190), .Z(n7183)
         );
  OR2_X1 U8866 ( .A1(n7190), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n7115) );
  INV_X1 U8867 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7926) );
  MUX2_X1 U8868 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n7926), .S(n7221), .Z(n7116)
         );
  NAND2_X1 U8869 ( .A1(n7117), .A2(n7116), .ZN(n9472) );
  OAI211_X1 U8870 ( .C1(n7117), .C2(n7116), .A(n10013), .B(n9472), .ZN(n7118)
         );
  OAI211_X1 U8871 ( .C1(n7120), .C2(n10023), .A(n7119), .B(n7118), .ZN(
        P1_U3250) );
  NAND2_X1 U8872 ( .A1(n7121), .A2(n7122), .ZN(n7124) );
  XNOR2_X1 U8873 ( .A(n7124), .B(n7123), .ZN(n7129) );
  AOI22_X1 U8874 ( .A1(n9427), .A2(n6723), .B1(n9386), .B2(n6711), .ZN(n7125)
         );
  OAI21_X1 U8875 ( .B1(n10078), .B2(n9417), .A(n7125), .ZN(n7126) );
  AOI21_X1 U8876 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n7127), .A(n7126), .ZN(
        n7128) );
  OAI21_X1 U8877 ( .B1(n7129), .B2(n9432), .A(n7128), .ZN(P1_U3220) );
  OAI211_X1 U8878 ( .C1(n7132), .C2(n7131), .A(n10003), .B(n7130), .ZN(n7134)
         );
  NOR2_X1 U8879 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n5887), .ZN(n7290) );
  INV_X1 U8880 ( .A(n7290), .ZN(n7133) );
  NAND2_X1 U8881 ( .A1(n7134), .A2(n7133), .ZN(n7135) );
  AOI21_X1 U8882 ( .B1(n9455), .B2(P1_ADDR_REG_3__SCAN_IN), .A(n7135), .ZN(
        n7142) );
  MUX2_X1 U8883 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n7984), .S(n7143), .Z(n7136)
         );
  NAND3_X1 U8884 ( .A1(n7138), .A2(n7137), .A3(n7136), .ZN(n7139) );
  NAND3_X1 U8885 ( .A1(n10013), .A2(n7140), .A3(n7139), .ZN(n7141) );
  OAI211_X1 U8886 ( .C1(n10017), .C2(n7143), .A(n7142), .B(n7141), .ZN(
        P1_U3244) );
  INV_X1 U8887 ( .A(n7144), .ZN(n7197) );
  AOI22_X1 U8888 ( .A1(n9488), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n10615), .ZN(n7145) );
  OAI21_X1 U8889 ( .B1(n7197), .B2(n9921), .A(n7145), .ZN(P1_U3338) );
  INV_X1 U8890 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10541) );
  INV_X1 U8891 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7150) );
  OAI211_X1 U8892 ( .C1(n7148), .C2(n7147), .A(n10003), .B(n7146), .ZN(n7149)
         );
  OAI21_X1 U8893 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7150), .A(n7149), .ZN(n7151) );
  AOI21_X1 U8894 ( .B1(n9455), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n7151), .ZN(
        n7157) );
  MUX2_X1 U8895 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n6974), .S(n8364), .Z(n7153)
         );
  NAND2_X1 U8896 ( .A1(n7153), .A2(n7152), .ZN(n7154) );
  NAND3_X1 U8897 ( .A1(n10013), .A2(n7155), .A3(n7154), .ZN(n7156) );
  OAI211_X1 U8898 ( .C1(n10017), .C2(n8364), .A(n7157), .B(n7156), .ZN(
        P1_U3242) );
  INV_X1 U8899 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7169) );
  AND3_X1 U8900 ( .A1(n10003), .A2(P1_IR_REG_0__SCAN_IN), .A3(n7158), .ZN(
        n7167) );
  NAND3_X1 U8901 ( .A1(n7160), .A2(n7159), .A3(P1_REG1_REG_0__SCAN_IN), .ZN(
        n7164) );
  XNOR2_X1 U8902 ( .A(n7162), .B(n7161), .ZN(n7163) );
  AOI21_X1 U8903 ( .B1(n7165), .B2(n7164), .A(n7163), .ZN(n7166) );
  AOI211_X1 U8904 ( .C1(P1_REG3_REG_0__SCAN_IN), .C2(P1_U3084), .A(n7167), .B(
        n7166), .ZN(n7168) );
  OAI21_X1 U8905 ( .B1(n10026), .B2(n7169), .A(n7168), .ZN(P1_U3241) );
  OAI21_X1 U8906 ( .B1(n7171), .B2(n7170), .A(n9450), .ZN(n7180) );
  NOR2_X1 U8907 ( .A1(n10017), .A2(n7172), .ZN(n7179) );
  INV_X1 U8908 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10475) );
  OAI21_X1 U8909 ( .B1(n7174), .B2(n4433), .A(n7173), .ZN(n7175) );
  NAND2_X1 U8910 ( .A1(n10003), .A2(n7175), .ZN(n7177) );
  NAND2_X1 U8911 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3084), .ZN(n7176) );
  OAI211_X1 U8912 ( .C1(n10475), .C2(n10026), .A(n7177), .B(n7176), .ZN(n7178)
         );
  AOI211_X1 U8913 ( .C1(n10013), .C2(n7180), .A(n7179), .B(n7178), .ZN(n7182)
         );
  NAND2_X1 U8914 ( .A1(n7182), .A2(n7181), .ZN(P1_U3245) );
  NAND2_X1 U8915 ( .A1(P1_U3084), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7856) );
  OAI21_X1 U8916 ( .B1(n10026), .B2(n4520), .A(n7856), .ZN(n7189) );
  INV_X1 U8917 ( .A(n7183), .ZN(n7185) );
  NAND3_X1 U8918 ( .A1(n7208), .A2(n7185), .A3(n7184), .ZN(n7186) );
  AOI21_X1 U8919 ( .B1(n7187), .B2(n7186), .A(n9994), .ZN(n7188) );
  AOI211_X1 U8920 ( .C1(n10001), .C2(n7190), .A(n7189), .B(n7188), .ZN(n7196)
         );
  NOR2_X1 U8921 ( .A1(n7192), .A2(n7191), .ZN(n7193) );
  OAI21_X1 U8922 ( .B1(n7194), .B2(n7193), .A(n10003), .ZN(n7195) );
  NAND2_X1 U8923 ( .A1(n7196), .A2(n7195), .ZN(P1_U3249) );
  OAI222_X1 U8924 ( .A1(n8368), .A2(n10567), .B1(n9281), .B2(n7197), .C1(
        P2_U3152), .C2(n8274), .ZN(P2_U3343) );
  OAI21_X1 U8925 ( .B1(n7200), .B2(n7199), .A(n7198), .ZN(n7201) );
  NAND2_X1 U8926 ( .A1(n7201), .A2(n9408), .ZN(n7204) );
  INV_X1 U8927 ( .A(n9365), .ZN(n9402) );
  OR2_X1 U8928 ( .A1(n10130), .A2(n7768), .ZN(n10083) );
  OAI22_X1 U8929 ( .A1(n9402), .A2(n10083), .B1(n7765), .B2(n9384), .ZN(n7202)
         );
  AOI21_X1 U8930 ( .B1(n9386), .B2(n10082), .A(n7202), .ZN(n7203) );
  OAI211_X1 U8931 ( .C1(n7205), .C2(n6972), .A(n7204), .B(n7203), .ZN(P1_U3235) );
  XOR2_X1 U8932 ( .A(n7207), .B(n7206), .Z(n7216) );
  AND2_X1 U8933 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7480) );
  INV_X1 U8934 ( .A(n7208), .ZN(n7209) );
  AOI21_X1 U8935 ( .B1(n7211), .B2(n7210), .A(n7209), .ZN(n7213) );
  OAI22_X1 U8936 ( .A1(n9994), .A2(n7213), .B1(n7212), .B2(n10017), .ZN(n7214)
         );
  AOI211_X1 U8937 ( .C1(n9455), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n7480), .B(
        n7214), .ZN(n7215) );
  OAI21_X1 U8938 ( .B1(n10023), .B2(n7216), .A(n7215), .ZN(P1_U3248) );
  OR2_X1 U8939 ( .A1(n7234), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7293) );
  NAND2_X1 U8940 ( .A1(n7234), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7294) );
  NAND2_X1 U8941 ( .A1(n7293), .A2(n7294), .ZN(n7220) );
  INV_X1 U8942 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n7219) );
  MUX2_X1 U8943 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n7219), .S(n9469), .Z(n9465)
         );
  MUX2_X1 U8944 ( .A(n7293), .B(n7220), .S(n7296), .Z(n7236) );
  NAND2_X1 U8945 ( .A1(n10003), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7227) );
  NAND2_X1 U8946 ( .A1(n7221), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9471) );
  NAND2_X1 U8947 ( .A1(n9472), .A2(n9471), .ZN(n7223) );
  INV_X1 U8948 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n9724) );
  MUX2_X1 U8949 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n9724), .S(n9469), .Z(n7222)
         );
  NAND2_X1 U8950 ( .A1(n7223), .A2(n7222), .ZN(n9474) );
  NAND2_X1 U8951 ( .A1(n9469), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n7224) );
  NAND2_X1 U8952 ( .A1(n9474), .A2(n7224), .ZN(n7229) );
  NAND3_X1 U8953 ( .A1(n7229), .A2(n7225), .A3(P1_REG2_REG_11__SCAN_IN), .ZN(
        n7226) );
  OAI211_X1 U8954 ( .C1(n7296), .C2(n7227), .A(n10017), .B(n7226), .ZN(n7233)
         );
  INV_X1 U8955 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n7228) );
  NAND2_X1 U8956 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7958) );
  OAI21_X1 U8957 ( .B1(n10026), .B2(n7228), .A(n7958), .ZN(n7232) );
  NOR3_X1 U8958 ( .A1(n7229), .A2(n7234), .A3(P1_REG2_REG_11__SCAN_IN), .ZN(
        n7230) );
  NOR3_X1 U8959 ( .A1(n7301), .A2(n7230), .A3(n9994), .ZN(n7231) );
  AOI211_X1 U8960 ( .C1(n7234), .C2(n7233), .A(n7232), .B(n7231), .ZN(n7235)
         );
  OAI21_X1 U8961 ( .B1(n7236), .B2(n10023), .A(n7235), .ZN(P1_U3252) );
  INV_X1 U8962 ( .A(n7237), .ZN(n7239) );
  INV_X1 U8963 ( .A(n9987), .ZN(n9481) );
  OAI222_X1 U8964 ( .A1(n4405), .A2(n7238), .B1(n9923), .B2(n7239), .C1(n9481), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  OAI222_X1 U8965 ( .A1(n8368), .A2(n10526), .B1(n8366), .B2(n7239), .C1(n8896), .C2(P2_U3152), .ZN(P2_U3342) );
  OAI22_X1 U8966 ( .A1(n8917), .A2(n7241), .B1(n7240), .B2(n8928), .ZN(n7245)
         );
  OR2_X1 U8967 ( .A1(n8928), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n7242) );
  OAI211_X1 U8968 ( .C1(n7243), .C2(P2_REG2_REG_0__SCAN_IN), .A(n7242), .B(
        n8932), .ZN(n7244) );
  INV_X1 U8969 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n7246) );
  INV_X1 U8970 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7935) );
  OAI22_X1 U8971 ( .A1(n7967), .A2(n7246), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7935), .ZN(n7247) );
  OR2_X1 U8972 ( .A1(n7248), .A2(n7247), .ZN(P2_U3245) );
  INV_X1 U8973 ( .A(n7249), .ZN(n7253) );
  AOI22_X1 U8974 ( .A1(n10000), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10615), .ZN(n7251) );
  OAI21_X1 U8975 ( .B1(n7253), .B2(n9921), .A(n7251), .ZN(P1_U3336) );
  AOI22_X1 U8976 ( .A1(n8905), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n9279), .ZN(n7252) );
  OAI21_X1 U8977 ( .B1(n7253), .B2(n8366), .A(n7252), .ZN(P2_U3341) );
  OR2_X1 U8978 ( .A1(n7254), .A2(P2_U3152), .ZN(n7255) );
  NAND2_X1 U8979 ( .A1(n7257), .A2(n7590), .ZN(n7307) );
  INV_X1 U8980 ( .A(n7307), .ZN(n7258) );
  NAND2_X1 U8981 ( .A1(n7592), .A2(n7258), .ZN(n7259) );
  INV_X1 U8982 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7281) );
  INV_X1 U8983 ( .A(n7261), .ZN(n7260) );
  NAND2_X1 U8984 ( .A1(n7260), .A2(n9133), .ZN(n8619) );
  NAND2_X1 U8985 ( .A1(n7261), .A2(n10214), .ZN(n8610) );
  NAND2_X1 U8986 ( .A1(n8619), .A2(n8610), .ZN(n8570) );
  NAND2_X1 U8987 ( .A1(n8570), .A2(n9132), .ZN(n9131) );
  OR2_X1 U8988 ( .A1(n9122), .A2(n9133), .ZN(n7262) );
  NAND2_X1 U8989 ( .A1(n9131), .A2(n7262), .ZN(n9116) );
  INV_X1 U8990 ( .A(n7265), .ZN(n7264) );
  NAND2_X2 U8991 ( .A1(n7264), .A2(n7263), .ZN(n7273) );
  NAND2_X1 U8992 ( .A1(n7265), .A2(n10222), .ZN(n8609) );
  AND2_X1 U8993 ( .A1(n7273), .A2(n8609), .ZN(n9119) );
  INV_X1 U8994 ( .A(n9119), .ZN(n9115) );
  NAND2_X1 U8995 ( .A1(n7349), .A2(n7347), .ZN(n7266) );
  OR2_X2 U8996 ( .A1(n7343), .A2(n7604), .ZN(n8624) );
  NAND2_X1 U8997 ( .A1(n7343), .A2(n7604), .ZN(n8628) );
  NAND2_X1 U8998 ( .A1(n7266), .A2(n7345), .ZN(n7638) );
  OR2_X1 U8999 ( .A1(n7266), .A2(n7345), .ZN(n7267) );
  NAND2_X1 U9000 ( .A1(n7638), .A2(n7267), .ZN(n7596) );
  INV_X1 U9001 ( .A(n9127), .ZN(n7268) );
  OAI21_X1 U9002 ( .B1(n7268), .B2(n7604), .A(n7644), .ZN(n7605) );
  INV_X1 U9003 ( .A(n7550), .ZN(n8758) );
  OAI22_X1 U9004 ( .A1(n7605), .A2(n10246), .B1(n7604), .B2(n10245), .ZN(n7279) );
  AND2_X1 U9005 ( .A1(n7269), .A2(n5122), .ZN(n7271) );
  NAND2_X1 U9006 ( .A1(n7595), .A2(n5811), .ZN(n7270) );
  NAND2_X1 U9007 ( .A1(n7271), .A2(n7270), .ZN(n7581) );
  INV_X1 U9008 ( .A(n7581), .ZN(n8137) );
  NAND2_X1 U9009 ( .A1(n7596), .A2(n8137), .ZN(n7278) );
  AOI22_X1 U9010 ( .A1(n9120), .A2(n8790), .B1(n8791), .B2(n9121), .ZN(n7277)
         );
  INV_X1 U9011 ( .A(n8374), .ZN(n7272) );
  NAND2_X1 U9012 ( .A1(n9118), .A2(n9119), .ZN(n9117) );
  NAND2_X1 U9013 ( .A1(n9117), .A2(n7273), .ZN(n7274) );
  OAI21_X1 U9014 ( .B1(n8614), .B2(n7274), .A(n7353), .ZN(n7275) );
  NAND2_X1 U9015 ( .A1(n8758), .A2(n8608), .ZN(n8566) );
  NAND2_X1 U9016 ( .A1(n7275), .A2(n9138), .ZN(n7276) );
  NAND3_X1 U9017 ( .A1(n7278), .A2(n7277), .A3(n7276), .ZN(n7597) );
  AOI211_X1 U9018 ( .C1(n10249), .C2(n7596), .A(n7279), .B(n7597), .ZN(n7309)
         );
  OR2_X1 U9019 ( .A1(n7309), .A2(n10253), .ZN(n7280) );
  OAI21_X1 U9020 ( .B1(n10254), .B2(n7281), .A(n7280), .ZN(P2_U3460) );
  INV_X1 U9021 ( .A(n7198), .ZN(n7285) );
  INV_X1 U9022 ( .A(n7282), .ZN(n7284) );
  NOR3_X1 U9023 ( .A1(n7285), .A2(n7284), .A3(n7283), .ZN(n7288) );
  INV_X1 U9024 ( .A(n7286), .ZN(n7287) );
  OAI21_X1 U9025 ( .B1(n7288), .B2(n7287), .A(n9408), .ZN(n7292) );
  OAI22_X1 U9026 ( .A1(n9417), .A2(n10096), .B1(n10042), .B2(n9425), .ZN(n7289) );
  AOI211_X1 U9027 ( .C1(n9427), .C2(n6711), .A(n7290), .B(n7289), .ZN(n7291)
         );
  OAI211_X1 U9028 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9429), .A(n7292), .B(
        n7291), .ZN(P1_U3216) );
  INV_X1 U9029 ( .A(n7293), .ZN(n7295) );
  XOR2_X1 U9030 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n7451), .Z(n7452) );
  XNOR2_X1 U9031 ( .A(n7453), .B(n7452), .ZN(n7306) );
  INV_X1 U9032 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7299) );
  OR2_X1 U9033 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7297), .ZN(n7298) );
  OAI21_X1 U9034 ( .B1(n10026), .B2(n7299), .A(n7298), .ZN(n7304) );
  INV_X1 U9035 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n8046) );
  XNOR2_X1 U9036 ( .A(n7451), .B(n8046), .ZN(n7300) );
  OAI211_X1 U9037 ( .C1(n7301), .C2(n7300), .A(n7447), .B(n10013), .ZN(n7302)
         );
  INV_X1 U9038 ( .A(n7302), .ZN(n7303) );
  AOI211_X1 U9039 ( .C1(n10001), .C2(n7451), .A(n7304), .B(n7303), .ZN(n7305)
         );
  OAI21_X1 U9040 ( .B1(n7306), .B2(n10023), .A(n7305), .ZN(P1_U3253) );
  OR2_X1 U9041 ( .A1(n7309), .A2(n10261), .ZN(n7310) );
  OAI21_X1 U9042 ( .B1(n10263), .B2(n6657), .A(n7310), .ZN(P2_U3523) );
  XNOR2_X1 U9043 ( .A(n7312), .B(n7311), .ZN(n7324) );
  AOI21_X1 U9044 ( .B1(n7315), .B2(n7314), .A(n7313), .ZN(n7316) );
  OR2_X1 U9045 ( .A1(n7316), .A2(n8917), .ZN(n7323) );
  NOR2_X1 U9046 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7317), .ZN(n7318) );
  AOI21_X1 U9047 ( .B1(n8922), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7318), .ZN(
        n7319) );
  OAI21_X1 U9048 ( .B1(n8932), .B2(n7320), .A(n7319), .ZN(n7321) );
  INV_X1 U9049 ( .A(n7321), .ZN(n7322) );
  OAI211_X1 U9050 ( .C1(n7324), .C2(n8928), .A(n7323), .B(n7322), .ZN(P2_U3256) );
  XNOR2_X1 U9051 ( .A(n7326), .B(n7325), .ZN(n7330) );
  AOI22_X1 U9052 ( .A1(n8541), .A2(n8790), .B1(n8495), .B2(n8791), .ZN(n7329)
         );
  INV_X1 U9053 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n8819) );
  MUX2_X1 U9054 ( .A(P2_U3152), .B(n8517), .S(n8819), .Z(n7327) );
  AOI21_X1 U9055 ( .B1(n8545), .B2(n7342), .A(n7327), .ZN(n7328) );
  OAI211_X1 U9056 ( .C1(n8549), .C2(n7330), .A(n7329), .B(n7328), .ZN(P2_U3220) );
  INV_X1 U9057 ( .A(n7331), .ZN(n7332) );
  NOR2_X1 U9058 ( .A1(n7333), .A2(n7332), .ZN(n7334) );
  XNOR2_X1 U9059 ( .A(n7335), .B(n7334), .ZN(n7341) );
  INV_X1 U9060 ( .A(n7641), .ZN(n7336) );
  NAND2_X1 U9061 ( .A1(n8517), .A2(n7336), .ZN(n7337) );
  NAND2_X1 U9062 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n8832) );
  NAND2_X1 U9063 ( .A1(n7337), .A2(n8832), .ZN(n7339) );
  INV_X1 U9064 ( .A(n7343), .ZN(n7650) );
  INV_X1 U9065 ( .A(n8789), .ZN(n7868) );
  OAI22_X1 U9066 ( .A1(n7650), .A2(n8543), .B1(n8498), .B2(n7868), .ZN(n7338)
         );
  AOI211_X1 U9067 ( .C1(n4905), .C2(n8545), .A(n7339), .B(n7338), .ZN(n7340)
         );
  OAI21_X1 U9068 ( .B1(n7341), .B2(n8549), .A(n7340), .ZN(P2_U3232) );
  INV_X1 U9069 ( .A(n10249), .ZN(n9237) );
  OR2_X1 U9070 ( .A1(n7343), .A2(n7342), .ZN(n7637) );
  INV_X1 U9071 ( .A(n7637), .ZN(n7344) );
  NAND2_X1 U9072 ( .A1(n8790), .A2(n10227), .ZN(n7567) );
  OAI21_X1 U9073 ( .B1(n7345), .B2(n7344), .A(n7647), .ZN(n7346) );
  INV_X1 U9074 ( .A(n7346), .ZN(n7351) );
  AND2_X1 U9075 ( .A1(n7347), .A2(n7637), .ZN(n7348) );
  NAND2_X1 U9076 ( .A1(n7349), .A2(n7348), .ZN(n7350) );
  OR2_X1 U9077 ( .A1(n8790), .A2(n4905), .ZN(n7352) );
  INV_X1 U9078 ( .A(n8616), .ZN(n8626) );
  NAND2_X1 U9079 ( .A1(n8789), .A2(n7412), .ZN(n8627) );
  NAND2_X1 U9080 ( .A1(n8626), .A2(n8627), .ZN(n8575) );
  NAND2_X1 U9081 ( .A1(n7552), .A2(n8575), .ZN(n7863) );
  OAI21_X1 U9082 ( .B1(n7552), .B2(n8575), .A(n7863), .ZN(n7807) );
  INV_X1 U9083 ( .A(n7807), .ZN(n7359) );
  NAND2_X1 U9084 ( .A1(n7569), .A2(n7567), .ZN(n7354) );
  XNOR2_X1 U9085 ( .A(n7354), .B(n8575), .ZN(n7355) );
  INV_X1 U9086 ( .A(n8788), .ZN(n7570) );
  OAI22_X1 U9087 ( .A1(n7570), .A2(n9102), .B1(n4906), .B2(n9100), .ZN(n7406)
         );
  AOI21_X1 U9088 ( .B1(n7355), .B2(n9138), .A(n7406), .ZN(n7814) );
  INV_X1 U9089 ( .A(n7412), .ZN(n7811) );
  OAI21_X1 U9090 ( .B1(n7356), .B2(n7412), .A(n9239), .ZN(n7357) );
  NOR2_X1 U9091 ( .A1(n7357), .A2(n7871), .ZN(n7806) );
  AOI21_X1 U9092 ( .B1(n9246), .B2(n7811), .A(n7806), .ZN(n7358) );
  OAI211_X1 U9093 ( .C1(n9250), .C2(n7359), .A(n7814), .B(n7358), .ZN(n7413)
         );
  NAND2_X1 U9094 ( .A1(n7413), .A2(n10254), .ZN(n7360) );
  OAI21_X1 U9095 ( .B1(n10254), .B2(n5231), .A(n7360), .ZN(P2_U3466) );
  AOI22_X1 U9096 ( .A1(n7263), .A2(n8545), .B1(n8541), .B2(n7343), .ZN(n7365)
         );
  XOR2_X1 U9097 ( .A(n7362), .B(n7361), .Z(n7363) );
  NAND2_X1 U9098 ( .A1(n8553), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8373) );
  AOI22_X1 U9099 ( .A1(n8457), .A2(n7363), .B1(n8373), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n7364) );
  OAI211_X1 U9100 ( .C1(n7260), .C2(n8543), .A(n7365), .B(n7364), .ZN(P2_U3239) );
  AOI22_X1 U9101 ( .A1(n10206), .A2(n8545), .B1(n8541), .B2(n9122), .ZN(n7369)
         );
  OAI21_X1 U9102 ( .B1(n7366), .B2(n9145), .A(n9137), .ZN(n7367) );
  AOI22_X1 U9103 ( .A1(n8457), .A2(n7367), .B1(n8373), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n7368) );
  OAI211_X1 U9104 ( .C1(n8618), .C2(n8473), .A(n7369), .B(n7368), .ZN(P2_U3234) );
  OAI211_X1 U9105 ( .C1(n7372), .C2(n7371), .A(n8874), .B(n7370), .ZN(n7380)
         );
  NAND2_X1 U9106 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n7404) );
  INV_X1 U9107 ( .A(n7404), .ZN(n7378) );
  INV_X1 U9108 ( .A(n8928), .ZN(n8811) );
  MUX2_X1 U9109 ( .A(n6661), .B(P2_REG1_REG_5__SCAN_IN), .S(n7373), .Z(n7374)
         );
  NAND3_X1 U9110 ( .A1(n8839), .A2(n7375), .A3(n7374), .ZN(n7376) );
  AND3_X1 U9111 ( .A1(n8811), .A2(n8852), .A3(n7376), .ZN(n7377) );
  AOI211_X1 U9112 ( .C1(P2_ADDR_REG_5__SCAN_IN), .C2(n8922), .A(n7378), .B(
        n7377), .ZN(n7379) );
  OAI211_X1 U9113 ( .C1(n8932), .C2(n7381), .A(n7380), .B(n7379), .ZN(P2_U3250) );
  XNOR2_X1 U9114 ( .A(n7383), .B(n7382), .ZN(n7392) );
  NAND2_X1 U9115 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n7818) );
  INV_X1 U9116 ( .A(n7818), .ZN(n7386) );
  NOR2_X1 U9117 ( .A1(n8932), .A2(n7384), .ZN(n7385) );
  AOI211_X1 U9118 ( .C1(P2_ADDR_REG_10__SCAN_IN), .C2(n8922), .A(n7386), .B(
        n7385), .ZN(n7391) );
  OAI211_X1 U9119 ( .C1(n7389), .C2(n7388), .A(n8874), .B(n7387), .ZN(n7390)
         );
  OAI211_X1 U9120 ( .C1(n7392), .C2(n8928), .A(n7391), .B(n7390), .ZN(P2_U3255) );
  XNOR2_X1 U9121 ( .A(n7394), .B(n7393), .ZN(n7402) );
  AND2_X1 U9122 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n7523) );
  NOR2_X1 U9123 ( .A1(n8932), .A2(n7395), .ZN(n7396) );
  AOI211_X1 U9124 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n8922), .A(n7523), .B(
        n7396), .ZN(n7401) );
  OAI211_X1 U9125 ( .C1(n7399), .C2(n7398), .A(n8874), .B(n7397), .ZN(n7400)
         );
  OAI211_X1 U9126 ( .C1(n7402), .C2(n8928), .A(n7401), .B(n7400), .ZN(P2_U3254) );
  INV_X1 U9127 ( .A(n7403), .ZN(n8555) );
  OAI21_X1 U9128 ( .B1(n8553), .B2(n7808), .A(n7404), .ZN(n7405) );
  AOI21_X1 U9129 ( .B1(n8555), .B2(n7406), .A(n7405), .ZN(n7411) );
  AOI21_X1 U9130 ( .B1(n7408), .B2(n7407), .A(n8549), .ZN(n7409) );
  NAND2_X1 U9131 ( .A1(n7409), .A2(n7441), .ZN(n7410) );
  OAI211_X1 U9132 ( .C1(n7412), .C2(n8558), .A(n7411), .B(n7410), .ZN(P2_U3229) );
  NAND2_X1 U9133 ( .A1(n7413), .A2(n10263), .ZN(n7414) );
  OAI21_X1 U9134 ( .B1(n10263), .B2(n6661), .A(n7414), .ZN(P2_U3525) );
  NAND2_X1 U9135 ( .A1(n8773), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n7415) );
  OAI21_X1 U9136 ( .B1(n8434), .B2(n8773), .A(n7415), .ZN(P2_U3581) );
  INV_X1 U9137 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n10340) );
  INV_X1 U9138 ( .A(n7416), .ZN(n7417) );
  OAI222_X1 U9139 ( .A1(n8368), .A2(n10340), .B1(n8366), .B2(n7417), .C1(
        P2_U3152), .C2(n8931), .ZN(P2_U3340) );
  INV_X1 U9140 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n10550) );
  INV_X1 U9141 ( .A(n9495), .ZN(n10016) );
  OAI222_X1 U9142 ( .A1(n4405), .A2(n10550), .B1(n9923), .B2(n7417), .C1(
        P1_U3084), .C2(n10016), .ZN(P1_U3335) );
  OAI211_X1 U9143 ( .C1(n7420), .C2(n7419), .A(n7418), .B(n8874), .ZN(n7428)
         );
  OAI21_X1 U9144 ( .B1(n7422), .B2(n7421), .A(n7508), .ZN(n7426) );
  AND2_X1 U9145 ( .A1(P2_U3152), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n7683) );
  AOI21_X1 U9146 ( .B1(n8922), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n7683), .ZN(
        n7423) );
  OAI21_X1 U9147 ( .B1(n8932), .B2(n7424), .A(n7423), .ZN(n7425) );
  AOI21_X1 U9148 ( .B1(n8811), .B2(n7426), .A(n7425), .ZN(n7427) );
  NAND2_X1 U9149 ( .A1(n7428), .A2(n7427), .ZN(P2_U3257) );
  INV_X1 U9150 ( .A(n7429), .ZN(n7431) );
  OAI222_X1 U9151 ( .A1(n8368), .A2(n7430), .B1(n8366), .B2(n7431), .C1(n5122), 
        .C2(P2_U3152), .ZN(P2_U3339) );
  OAI222_X1 U9152 ( .A1(n4405), .A2(n7432), .B1(n9923), .B2(n7431), .C1(
        P1_U3084), .C2(n9568), .ZN(P1_U3334) );
  INV_X1 U9153 ( .A(n7883), .ZN(n8787) );
  INV_X1 U9154 ( .A(n7874), .ZN(n7433) );
  AND2_X1 U9155 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n8848) );
  AOI21_X1 U9156 ( .B1(n8517), .B2(n7433), .A(n8848), .ZN(n7434) );
  OAI21_X1 U9157 ( .B1(n8558), .B2(n10232), .A(n7434), .ZN(n7439) );
  INV_X1 U9158 ( .A(n7442), .ZN(n7436) );
  NAND3_X1 U9159 ( .A1(n8535), .A2(n7436), .A3(n7435), .ZN(n7437) );
  AOI21_X1 U9160 ( .B1(n7437), .B2(n8543), .A(n7868), .ZN(n7438) );
  AOI211_X1 U9161 ( .C1(n8541), .C2(n8787), .A(n7439), .B(n7438), .ZN(n7445)
         );
  OAI21_X1 U9162 ( .B1(n7442), .B2(n7441), .A(n7440), .ZN(n7443) );
  NAND2_X1 U9163 ( .A1(n7443), .A2(n8457), .ZN(n7444) );
  NAND2_X1 U9164 ( .A1(n7445), .A2(n7444), .ZN(P2_U3241) );
  INV_X1 U9165 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7832) );
  NAND2_X1 U9166 ( .A1(n7451), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7446) );
  INV_X1 U9167 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7448) );
  XNOR2_X1 U9168 ( .A(n7454), .B(n7448), .ZN(n9970) );
  NAND2_X1 U9169 ( .A1(n9971), .A2(n9970), .ZN(n9969) );
  NAND2_X1 U9170 ( .A1(n7454), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n7449) );
  NAND2_X1 U9171 ( .A1(n9969), .A2(n7449), .ZN(n7830) );
  XNOR2_X1 U9172 ( .A(n7830), .B(n7825), .ZN(n7833) );
  XOR2_X1 U9173 ( .A(n7832), .B(n7833), .Z(n7462) );
  INV_X1 U9174 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7450) );
  NAND2_X1 U9175 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9292) );
  OAI21_X1 U9176 ( .B1(n10026), .B2(n7450), .A(n9292), .ZN(n7460) );
  AOI22_X1 U9177 ( .A1(n7453), .A2(n7452), .B1(n7451), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n9977) );
  NOR2_X1 U9178 ( .A1(n7454), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7455) );
  AOI21_X1 U9179 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n7454), .A(n7455), .ZN(
        n9976) );
  AND2_X1 U9180 ( .A1(n9977), .A2(n9976), .ZN(n9978) );
  NOR2_X1 U9181 ( .A1(n9978), .A2(n7455), .ZN(n7457) );
  XNOR2_X1 U9182 ( .A(n7829), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7456) );
  AOI21_X1 U9183 ( .B1(n7457), .B2(n7456), .A(n7824), .ZN(n7458) );
  NOR2_X1 U9184 ( .A1(n7458), .A2(n10023), .ZN(n7459) );
  AOI211_X1 U9185 ( .C1(n10001), .C2(n7829), .A(n7460), .B(n7459), .ZN(n7461)
         );
  OAI21_X1 U9186 ( .B1(n9994), .B2(n7462), .A(n7461), .ZN(P1_U3255) );
  OAI22_X1 U9187 ( .A1(n8553), .A2(n7843), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5298), .ZN(n7464) );
  OAI22_X1 U9188 ( .A1(n7570), .A2(n8543), .B1(n8498), .B2(n7577), .ZN(n7463)
         );
  AOI211_X1 U9189 ( .C1(n10237), .C2(n8545), .A(n7464), .B(n7463), .ZN(n7468)
         );
  NAND2_X1 U9190 ( .A1(n7465), .A2(n7466), .ZN(n7495) );
  OAI211_X1 U9191 ( .C1(n7465), .C2(n7466), .A(n7495), .B(n8457), .ZN(n7467)
         );
  NAND2_X1 U9192 ( .A1(n7468), .A2(n7467), .ZN(P2_U3215) );
  INV_X1 U9193 ( .A(n7469), .ZN(n8003) );
  AOI21_X1 U9194 ( .B1(n7470), .B2(n7472), .A(n7471), .ZN(n7474) );
  INV_X1 U9195 ( .A(n7534), .ZN(n7473) );
  NOR2_X1 U9196 ( .A1(n7474), .A2(n7473), .ZN(n7477) );
  OAI21_X1 U9197 ( .B1(n7477), .B2(n7476), .A(n7475), .ZN(n7478) );
  NAND2_X1 U9198 ( .A1(n7478), .A2(n9408), .ZN(n7482) );
  OAI22_X1 U9199 ( .A1(n9417), .A2(n8001), .B1(n10043), .B2(n9384), .ZN(n7479)
         );
  AOI211_X1 U9200 ( .C1(n9386), .C2(n10158), .A(n7480), .B(n7479), .ZN(n7481)
         );
  OAI211_X1 U9201 ( .C1(n9429), .C2(n8003), .A(n7482), .B(n7481), .ZN(P1_U3211) );
  INV_X1 U9202 ( .A(n7483), .ZN(n7484) );
  NAND2_X1 U9203 ( .A1(n7470), .A2(n7484), .ZN(n7536) );
  OAI21_X1 U9204 ( .B1(n7470), .B2(n7484), .A(n7536), .ZN(n7485) );
  NOR2_X1 U9205 ( .A1(n7485), .A2(n7486), .ZN(n7538) );
  AOI21_X1 U9206 ( .B1(n7486), .B2(n7485), .A(n7538), .ZN(n7491) );
  NAND2_X1 U9207 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9461) );
  INV_X1 U9208 ( .A(n9461), .ZN(n7488) );
  OAI22_X1 U9209 ( .A1(n9417), .A2(n5032), .B1(n10043), .B2(n9425), .ZN(n7487)
         );
  AOI211_X1 U9210 ( .C1(n9427), .C2(n9444), .A(n7488), .B(n7487), .ZN(n7490)
         );
  NAND2_X1 U9211 ( .A1(n9410), .A2(n10032), .ZN(n7489) );
  OAI211_X1 U9212 ( .C1(n7491), .C2(n9432), .A(n7490), .B(n7489), .ZN(P1_U3225) );
  NAND2_X1 U9213 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n8877) );
  OAI21_X1 U9214 ( .B1(n8553), .B2(n7893), .A(n8877), .ZN(n7493) );
  OAI22_X1 U9215 ( .A1(n7884), .A2(n8498), .B1(n8543), .B2(n7883), .ZN(n7492)
         );
  AOI211_X1 U9216 ( .C1(n10244), .C2(n8545), .A(n7493), .B(n7492), .ZN(n7502)
         );
  AOI21_X1 U9217 ( .B1(n7495), .B2(n7494), .A(n8549), .ZN(n7500) );
  NOR3_X1 U9218 ( .A1(n8473), .A2(n7883), .A3(n7496), .ZN(n7499) );
  NAND2_X1 U9219 ( .A1(n7465), .A2(n7497), .ZN(n7521) );
  AND2_X1 U9220 ( .A1(n7498), .A2(n7521), .ZN(n7516) );
  OAI21_X1 U9221 ( .B1(n7500), .B2(n7499), .A(n7516), .ZN(n7501) );
  NAND2_X1 U9222 ( .A1(n7502), .A2(n7501), .ZN(P2_U3223) );
  AOI21_X1 U9223 ( .B1(n7505), .B2(n7504), .A(n7503), .ZN(n7515) );
  NAND2_X1 U9224 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8113) );
  OAI21_X1 U9225 ( .B1(n7967), .B2(n4515), .A(n8113), .ZN(n7512) );
  INV_X1 U9226 ( .A(n7970), .ZN(n7510) );
  NAND3_X1 U9227 ( .A1(n7508), .A2(n7507), .A3(n7506), .ZN(n7509) );
  AOI21_X1 U9228 ( .B1(n7510), .B2(n7509), .A(n8928), .ZN(n7511) );
  AOI211_X1 U9229 ( .C1(n8878), .C2(n7513), .A(n7512), .B(n7511), .ZN(n7514)
         );
  OAI21_X1 U9230 ( .B1(n7515), .B2(n8917), .A(n7514), .ZN(P2_U3258) );
  INV_X1 U9231 ( .A(n7516), .ZN(n7520) );
  INV_X1 U9232 ( .A(n7517), .ZN(n7518) );
  NOR3_X1 U9233 ( .A1(n8473), .A2(n7577), .A3(n7518), .ZN(n7519) );
  AOI21_X1 U9234 ( .B1(n7520), .B2(n8457), .A(n7519), .ZN(n7531) );
  AND2_X1 U9235 ( .A1(n7522), .A2(n7521), .ZN(n7528) );
  INV_X1 U9236 ( .A(n7904), .ZN(n7566) );
  INV_X1 U9237 ( .A(n7654), .ZN(n8784) );
  INV_X1 U9238 ( .A(n7577), .ZN(n8786) );
  AOI22_X1 U9239 ( .A1(n8541), .A2(n8784), .B1(n8495), .B2(n8786), .ZN(n7526)
         );
  INV_X1 U9240 ( .A(n7899), .ZN(n7524) );
  AOI21_X1 U9241 ( .B1(n8517), .B2(n7524), .A(n7523), .ZN(n7525) );
  OAI211_X1 U9242 ( .C1(n7566), .C2(n8558), .A(n7526), .B(n7525), .ZN(n7527)
         );
  AOI21_X1 U9243 ( .B1(n7528), .B2(n8457), .A(n7527), .ZN(n7529) );
  OAI21_X1 U9244 ( .B1(n7531), .B2(n7530), .A(n7529), .ZN(P2_U3233) );
  INV_X1 U9245 ( .A(n7532), .ZN(n7549) );
  OAI222_X1 U9246 ( .A1(n4405), .A2(n7533), .B1(n9923), .B2(n7549), .C1(n6279), 
        .C2(P1_U3084), .ZN(P1_U3333) );
  NAND2_X1 U9247 ( .A1(n7535), .A2(n7534), .ZN(n7540) );
  INV_X1 U9248 ( .A(n7536), .ZN(n7537) );
  NOR2_X1 U9249 ( .A1(n7538), .A2(n7537), .ZN(n7539) );
  XOR2_X1 U9250 ( .A(n7540), .B(n7539), .Z(n7548) );
  OR2_X1 U9251 ( .A1(n10130), .A2(n7632), .ZN(n10115) );
  NAND2_X1 U9252 ( .A1(n10159), .A2(n9442), .ZN(n7541) );
  OAI21_X1 U9253 ( .B1(n7542), .B2(n10138), .A(n7541), .ZN(n7622) );
  INV_X1 U9254 ( .A(n7543), .ZN(n9361) );
  NAND2_X1 U9255 ( .A1(n7622), .A2(n9361), .ZN(n7544) );
  OAI211_X1 U9256 ( .C1(n9402), .C2(n10115), .A(n7545), .B(n7544), .ZN(n7546)
         );
  AOI21_X1 U9257 ( .B1(n7630), .B2(n9410), .A(n7546), .ZN(n7547) );
  OAI21_X1 U9258 ( .B1(n7548), .B2(n9432), .A(n7547), .ZN(P1_U3237) );
  OAI222_X1 U9259 ( .A1(n8368), .A2(n10434), .B1(P2_U3152), .B2(n7550), .C1(
        n8366), .C2(n7549), .ZN(P2_U3338) );
  OR2_X1 U9260 ( .A1(n7904), .A2(n7884), .ZN(n8650) );
  NAND2_X1 U9261 ( .A1(n7904), .A2(n7884), .ZN(n8647) );
  INV_X1 U9262 ( .A(n10232), .ZN(n7876) );
  NAND2_X1 U9263 ( .A1(n7876), .A2(n8788), .ZN(n7553) );
  AND2_X1 U9264 ( .A1(n8575), .A2(n7553), .ZN(n7551) );
  NAND2_X1 U9265 ( .A1(n7552), .A2(n7551), .ZN(n7558) );
  INV_X1 U9266 ( .A(n7553), .ZN(n7556) );
  OR2_X1 U9267 ( .A1(n8789), .A2(n7811), .ZN(n7862) );
  OR2_X1 U9268 ( .A1(n8788), .A2(n7876), .ZN(n7554) );
  AND2_X1 U9269 ( .A1(n7862), .A2(n7554), .ZN(n7555) );
  OR2_X1 U9270 ( .A1(n7556), .A2(n7555), .ZN(n7557) );
  NAND2_X1 U9271 ( .A1(n7558), .A2(n7557), .ZN(n7847) );
  OR2_X1 U9272 ( .A1(n10237), .A2(n7883), .ZN(n8641) );
  NAND2_X1 U9273 ( .A1(n10237), .A2(n7883), .ZN(n8653) );
  NAND2_X1 U9274 ( .A1(n7847), .A2(n7848), .ZN(n7560) );
  OR2_X1 U9275 ( .A1(n10237), .A2(n8787), .ZN(n7559) );
  NAND2_X1 U9276 ( .A1(n7560), .A2(n7559), .ZN(n7879) );
  OR2_X1 U9277 ( .A1(n10244), .A2(n7577), .ZN(n8644) );
  NAND2_X1 U9278 ( .A1(n10244), .A2(n7577), .ZN(n8642) );
  NAND2_X1 U9279 ( .A1(n10244), .A2(n8786), .ZN(n7561) );
  INV_X1 U9280 ( .A(n7653), .ZN(n7562) );
  AOI21_X1 U9281 ( .B1(n8576), .B2(n7944), .A(n7562), .ZN(n7907) );
  INV_X1 U9282 ( .A(n7907), .ZN(n7583) );
  AND2_X2 U9283 ( .A1(n7564), .A2(n7566), .ZN(n7656) );
  INV_X1 U9284 ( .A(n7656), .ZN(n7565) );
  OAI21_X1 U9285 ( .B1(n7566), .B2(n7891), .A(n7565), .ZN(n7901) );
  OAI22_X1 U9286 ( .A1(n7901), .A2(n10246), .B1(n7566), .B2(n10245), .ZN(n7582) );
  AND2_X1 U9287 ( .A1(n8627), .A2(n7567), .ZN(n8629) );
  NAND2_X1 U9288 ( .A1(n10232), .A2(n8788), .ZN(n8633) );
  NAND2_X1 U9289 ( .A1(n7569), .A2(n7568), .ZN(n7573) );
  NAND2_X1 U9290 ( .A1(n8616), .A2(n8633), .ZN(n7571) );
  NAND2_X1 U9291 ( .A1(n7570), .A2(n7876), .ZN(n8638) );
  NAND2_X1 U9292 ( .A1(n7573), .A2(n7572), .ZN(n7574) );
  NAND2_X1 U9293 ( .A1(n7574), .A2(n8639), .ZN(n7840) );
  NAND2_X1 U9294 ( .A1(n7840), .A2(n8653), .ZN(n7575) );
  NAND2_X1 U9295 ( .A1(n7575), .A2(n8655), .ZN(n7882) );
  NAND2_X1 U9296 ( .A1(n7882), .A2(n8642), .ZN(n7576) );
  OAI21_X1 U9297 ( .B1(n8576), .B2(n7576), .A(n7658), .ZN(n7579) );
  OAI22_X1 U9298 ( .A1(n7654), .A2(n9102), .B1(n7577), .B2(n9100), .ZN(n7578)
         );
  AOI21_X1 U9299 ( .B1(n7579), .B2(n9138), .A(n7578), .ZN(n7580) );
  OAI21_X1 U9300 ( .B1(n7907), .B2(n7581), .A(n7580), .ZN(n7898) );
  AOI211_X1 U9301 ( .C1(n10249), .C2(n7583), .A(n7582), .B(n7898), .ZN(n7586)
         );
  NAND2_X1 U9302 ( .A1(n10261), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7584) );
  OAI21_X1 U9303 ( .B1(n7586), .B2(n10261), .A(n7584), .ZN(P2_U3529) );
  NAND2_X1 U9304 ( .A1(n10253), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n7585) );
  OAI21_X1 U9305 ( .B1(n7586), .B2(n10253), .A(n7585), .ZN(P2_U3478) );
  INV_X1 U9306 ( .A(n7587), .ZN(n7699) );
  AOI22_X1 U9307 ( .A1(n8608), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n9279), .ZN(n7588) );
  OAI21_X1 U9308 ( .B1(n7699), .B2(n9281), .A(n7588), .ZN(P2_U3337) );
  INV_X1 U9309 ( .A(n7589), .ZN(n7594) );
  INV_X1 U9310 ( .A(n7590), .ZN(n7591) );
  NOR2_X1 U9311 ( .A1(n7595), .A2(n5122), .ZN(n7636) );
  AND2_X1 U9312 ( .A1(n9144), .A2(n7636), .ZN(n7880) );
  NAND2_X1 U9313 ( .A1(n7880), .A2(n7596), .ZN(n7599) );
  INV_X1 U9314 ( .A(n9124), .ZN(n9143) );
  AOI22_X1 U9315 ( .A1(n9144), .A2(n7597), .B1(n9143), .B2(n8819), .ZN(n7598)
         );
  OAI211_X1 U9316 ( .C1(n9144), .C2(n7600), .A(n7599), .B(n7598), .ZN(n7607)
         );
  INV_X1 U9317 ( .A(n7601), .ZN(n7602) );
  NAND2_X1 U9318 ( .A1(n9148), .A2(n9239), .ZN(n9021) );
  OAI22_X1 U9319 ( .A1(n9021), .A2(n7605), .B1(n9088), .B2(n7604), .ZN(n7606)
         );
  OR2_X1 U9320 ( .A1(n7607), .A2(n7606), .ZN(P2_U3293) );
  INV_X1 U9321 ( .A(n7608), .ZN(n7610) );
  NOR3_X1 U9322 ( .A1(n7611), .A2(n7610), .A3(n7609), .ZN(n7612) );
  NAND2_X1 U9323 ( .A1(n7613), .A2(n7612), .ZN(n7927) );
  NAND2_X1 U9324 ( .A1(n7614), .A2(n7698), .ZN(n7615) );
  INV_X1 U9325 ( .A(n7616), .ZN(n7617) );
  NAND2_X1 U9326 ( .A1(n7617), .A2(n10052), .ZN(n9708) );
  NAND2_X1 U9327 ( .A1(n6712), .A2(n9708), .ZN(n10045) );
  OR2_X1 U9328 ( .A1(n7618), .A2(n7620), .ZN(n7996) );
  NAND2_X1 U9329 ( .A1(n7618), .A2(n7620), .ZN(n7619) );
  XNOR2_X1 U9330 ( .A(n7621), .B(n7620), .ZN(n7623) );
  AOI21_X1 U9331 ( .B1(n7623), .B2(n10168), .A(n7622), .ZN(n10121) );
  MUX2_X1 U9332 ( .A(n7624), .B(n10121), .S(n9711), .Z(n7635) );
  AND2_X1 U9333 ( .A1(n10030), .A2(n7625), .ZN(n7626) );
  NOR2_X1 U9334 ( .A1(n8002), .A2(n7626), .ZN(n10118) );
  NOR2_X1 U9335 ( .A1(n7628), .A2(n7627), .ZN(n7629) );
  INV_X1 U9336 ( .A(n7630), .ZN(n7631) );
  OAI22_X1 U9337 ( .A1(n9725), .A2(n7632), .B1(n9728), .B2(n7631), .ZN(n7633)
         );
  AOI21_X1 U9338 ( .B1(n10118), .B2(n9718), .A(n7633), .ZN(n7634) );
  OAI211_X1 U9339 ( .C1(n9738), .C2(n10120), .A(n7635), .B(n7634), .ZN(
        P1_U3285) );
  OAI21_X2 U9340 ( .B1(n8137), .B2(n7636), .A(n9144), .ZN(n9114) );
  INV_X1 U9341 ( .A(n9114), .ZN(n9135) );
  INV_X1 U9342 ( .A(n7647), .ZN(n8571) );
  NAND3_X1 U9343 ( .A1(n7638), .A2(n8571), .A3(n7637), .ZN(n7640) );
  NAND2_X1 U9344 ( .A1(n7640), .A2(n7639), .ZN(n10230) );
  OAI22_X1 U9345 ( .A1(n9144), .A2(n7642), .B1(n7641), .B2(n9124), .ZN(n7643)
         );
  AOI21_X1 U9346 ( .B1(n9135), .B2(n10230), .A(n7643), .ZN(n7652) );
  NAND2_X1 U9347 ( .A1(n7644), .A2(n4905), .ZN(n7645) );
  NAND2_X1 U9348 ( .A1(n7645), .A2(n9239), .ZN(n7646) );
  NOR2_X1 U9349 ( .A1(n7356), .A2(n7646), .ZN(n10225) );
  XNOR2_X1 U9350 ( .A(n7648), .B(n7647), .ZN(n7649) );
  OAI222_X1 U9351 ( .A1(n9102), .A2(n7868), .B1(n9100), .B2(n7650), .C1(n7649), 
        .C2(n9081), .ZN(n10228) );
  AOI22_X1 U9352 ( .A1(n10225), .A2(n9148), .B1(n10228), .B2(n9144), .ZN(n7651) );
  OAI211_X1 U9353 ( .C1(n10227), .C2(n9088), .A(n7652), .B(n7651), .ZN(
        P2_U3292) );
  INV_X1 U9354 ( .A(n7884), .ZN(n8785) );
  OR2_X1 U9355 ( .A1(n7904), .A2(n8785), .ZN(n7732) );
  NAND2_X1 U9356 ( .A1(n7653), .A2(n7732), .ZN(n7655) );
  OR2_X1 U9357 ( .A1(n7915), .A2(n7654), .ZN(n8657) );
  NAND2_X1 U9358 ( .A1(n7915), .A2(n7654), .ZN(n8648) );
  NAND2_X1 U9359 ( .A1(n8657), .A2(n8648), .ZN(n8578) );
  XNOR2_X1 U9360 ( .A(n7655), .B(n8578), .ZN(n7908) );
  INV_X1 U9361 ( .A(n7915), .ZN(n7657) );
  OAI21_X1 U9362 ( .B1(n7656), .B2(n7657), .A(n7757), .ZN(n7912) );
  OAI22_X1 U9363 ( .A1(n7912), .A2(n10246), .B1(n7657), .B2(n10245), .ZN(n7662) );
  XNOR2_X1 U9364 ( .A(n7747), .B(n8578), .ZN(n7661) );
  NAND2_X1 U9365 ( .A1(n7908), .A2(n8137), .ZN(n7660) );
  INV_X1 U9366 ( .A(n7820), .ZN(n8783) );
  AOI22_X1 U9367 ( .A1(n9121), .A2(n8785), .B1(n8783), .B2(n9120), .ZN(n7659)
         );
  OAI211_X1 U9368 ( .C1(n9081), .C2(n7661), .A(n7660), .B(n7659), .ZN(n7909)
         );
  AOI211_X1 U9369 ( .C1(n10249), .C2(n7908), .A(n7662), .B(n7909), .ZN(n7665)
         );
  NAND2_X1 U9370 ( .A1(n10253), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n7663) );
  OAI21_X1 U9371 ( .B1(n7665), .B2(n10253), .A(n7663), .ZN(P2_U3481) );
  NAND2_X1 U9372 ( .A1(n10261), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7664) );
  OAI21_X1 U9373 ( .B1(n7665), .B2(n10261), .A(n7664), .ZN(P2_U3530) );
  INV_X1 U9374 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7672) );
  OAI21_X1 U9375 ( .B1(n9713), .B2(n9718), .A(n7666), .ZN(n7671) );
  INV_X1 U9376 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7667) );
  NOR2_X1 U9377 ( .A1(n9728), .A2(n7667), .ZN(n7668) );
  OAI21_X1 U9378 ( .B1(n7669), .B2(n7668), .A(n9711), .ZN(n7670) );
  OAI211_X1 U9379 ( .C1(n7672), .C2(n9711), .A(n7671), .B(n7670), .ZN(P1_U3291) );
  NOR3_X1 U9380 ( .A1(n8473), .A2(n7820), .A3(n7674), .ZN(n7675) );
  AOI21_X1 U9381 ( .B1(n7673), .B2(n8457), .A(n7675), .ZN(n7690) );
  INV_X1 U9382 ( .A(n7676), .ZN(n7677) );
  XNOR2_X1 U9383 ( .A(n7678), .B(n7677), .ZN(n7689) );
  AND2_X1 U9384 ( .A1(n7689), .A2(n7679), .ZN(n7680) );
  NAND2_X1 U9385 ( .A1(n7681), .A2(n7680), .ZN(n8093) );
  INV_X1 U9386 ( .A(n8093), .ZN(n7687) );
  AOI22_X1 U9387 ( .A1(n8495), .A2(n8783), .B1(n8541), .B2(n8781), .ZN(n7685)
         );
  INV_X1 U9388 ( .A(n7682), .ZN(n7786) );
  AOI21_X1 U9389 ( .B1(n8517), .B2(n7786), .A(n7683), .ZN(n7684) );
  OAI211_X1 U9390 ( .C1(n7758), .C2(n8558), .A(n7685), .B(n7684), .ZN(n7686)
         );
  AOI21_X1 U9391 ( .B1(n7687), .B2(n8457), .A(n7686), .ZN(n7688) );
  OAI21_X1 U9392 ( .B1(n7690), .B2(n7689), .A(n7688), .ZN(P2_U3226) );
  XOR2_X1 U9393 ( .A(n7691), .B(n7692), .Z(n7697) );
  NAND2_X1 U9394 ( .A1(n9386), .A2(n9960), .ZN(n7693) );
  NAND2_X1 U9395 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9467) );
  OAI211_X1 U9396 ( .C1(n9730), .C2(n9384), .A(n7693), .B(n9467), .ZN(n7695)
         );
  NOR2_X1 U9397 ( .A1(n9417), .A2(n9963), .ZN(n7694) );
  AOI211_X1 U9398 ( .C1(n9410), .C2(n9727), .A(n7695), .B(n7694), .ZN(n7696)
         );
  OAI21_X1 U9399 ( .B1(n7697), .B2(n9432), .A(n7696), .ZN(P1_U3215) );
  OAI222_X1 U9400 ( .A1(n4405), .A2(n7700), .B1(n9923), .B2(n7699), .C1(n7698), 
        .C2(P1_U3084), .ZN(P1_U3332) );
  NAND3_X1 U9401 ( .A1(n8535), .A2(n8784), .A3(n7701), .ZN(n7707) );
  NAND2_X1 U9402 ( .A1(n7465), .A2(n7702), .ZN(n7703) );
  AND2_X1 U9403 ( .A1(n7704), .A2(n7703), .ZN(n7816) );
  NOR2_X1 U9404 ( .A1(n7816), .A2(n7817), .ZN(n7815) );
  OAI21_X1 U9405 ( .B1(n7815), .B2(n7705), .A(n8457), .ZN(n7706) );
  AOI21_X1 U9406 ( .B1(n7707), .B2(n7706), .A(n7673), .ZN(n7712) );
  INV_X1 U9407 ( .A(n9245), .ZN(n7951) );
  INV_X1 U9408 ( .A(n8116), .ZN(n8782) );
  AOI22_X1 U9409 ( .A1(n8495), .A2(n8784), .B1(n8541), .B2(n8782), .ZN(n7710)
         );
  INV_X1 U9410 ( .A(n7950), .ZN(n7708) );
  AOI22_X1 U9411 ( .A1(n8517), .A2(n7708), .B1(P2_REG3_REG_11__SCAN_IN), .B2(
        P2_U3152), .ZN(n7709) );
  OAI211_X1 U9412 ( .C1(n7951), .C2(n8558), .A(n7710), .B(n7709), .ZN(n7711)
         );
  OR2_X1 U9413 ( .A1(n7712), .A2(n7711), .ZN(P2_U3238) );
  AOI21_X1 U9414 ( .B1(n7713), .B2(n7985), .A(n7714), .ZN(n7715) );
  XOR2_X1 U9415 ( .A(n7719), .B(n7715), .Z(n10108) );
  INV_X1 U9416 ( .A(n10108), .ZN(n10105) );
  NAND2_X1 U9417 ( .A1(n7716), .A2(n7717), .ZN(n7718) );
  XOR2_X1 U9418 ( .A(n7719), .B(n7718), .Z(n7723) );
  NAND2_X1 U9419 ( .A1(n10159), .A2(n9443), .ZN(n7720) );
  OAI21_X1 U9420 ( .B1(n7721), .B2(n10138), .A(n7720), .ZN(n9362) );
  INV_X1 U9421 ( .A(n9362), .ZN(n7722) );
  OAI21_X1 U9422 ( .B1(n7723), .B2(n10040), .A(n7722), .ZN(n10106) );
  NAND2_X1 U9423 ( .A1(n10106), .A2(n9711), .ZN(n7730) );
  NAND2_X1 U9424 ( .A1(n7988), .A2(n7724), .ZN(n7725) );
  AND2_X1 U9425 ( .A1(n10028), .A2(n7725), .ZN(n10103) );
  INV_X1 U9426 ( .A(n9363), .ZN(n7726) );
  OAI22_X1 U9427 ( .A1(n9711), .A2(n10464), .B1(n7726), .B2(n9728), .ZN(n7728)
         );
  NOR2_X1 U9428 ( .A1(n9725), .A2(n9364), .ZN(n7727) );
  AOI211_X1 U9429 ( .C1(n10103), .C2(n9718), .A(n7728), .B(n7727), .ZN(n7729)
         );
  OAI211_X1 U9430 ( .C1(n9738), .C2(n10105), .A(n7730), .B(n7729), .ZN(
        P1_U3287) );
  AND2_X1 U9431 ( .A1(n8578), .A2(n7732), .ZN(n7943) );
  OR2_X1 U9432 ( .A1(n9245), .A2(n7820), .ZN(n8658) );
  AND2_X1 U9433 ( .A1(n9245), .A2(n7820), .ZN(n7780) );
  INV_X1 U9434 ( .A(n7780), .ZN(n8669) );
  NAND2_X1 U9435 ( .A1(n8658), .A2(n8669), .ZN(n8579) );
  NAND3_X1 U9436 ( .A1(n7731), .A2(n7943), .A3(n8579), .ZN(n7739) );
  INV_X1 U9437 ( .A(n8576), .ZN(n7734) );
  INV_X1 U9438 ( .A(n7732), .ZN(n7733) );
  NOR2_X1 U9439 ( .A1(n7734), .A2(n7733), .ZN(n7735) );
  NAND2_X1 U9440 ( .A1(n8578), .A2(n7735), .ZN(n7737) );
  NAND2_X1 U9441 ( .A1(n7915), .A2(n8784), .ZN(n7736) );
  NAND2_X1 U9442 ( .A1(n7737), .A2(n7736), .ZN(n7942) );
  AOI22_X1 U9443 ( .A1(n7942), .A2(n8579), .B1(n8783), .B2(n9245), .ZN(n7738)
         );
  NAND2_X1 U9444 ( .A1(n7739), .A2(n7738), .ZN(n7790) );
  INV_X1 U9445 ( .A(n7790), .ZN(n7741) );
  OR2_X1 U9446 ( .A1(n9238), .A2(n8116), .ZN(n8672) );
  NAND2_X1 U9447 ( .A1(n9238), .A2(n8116), .ZN(n8670) );
  INV_X1 U9448 ( .A(n8583), .ZN(n7740) );
  OR2_X1 U9449 ( .A1(n9238), .A2(n8782), .ZN(n7742) );
  INV_X1 U9450 ( .A(n8667), .ZN(n7743) );
  INV_X1 U9451 ( .A(n8088), .ZN(n7744) );
  AOI21_X1 U9452 ( .B1(n8667), .B2(n7745), .A(n7744), .ZN(n9231) );
  OAI22_X1 U9453 ( .A1(n8112), .A2(n9102), .B1(n8116), .B2(n9100), .ZN(n7756)
         );
  AND2_X1 U9454 ( .A1(n8672), .A2(n8658), .ZN(n8662) );
  AND2_X1 U9455 ( .A1(n8657), .A2(n8662), .ZN(n7746) );
  INV_X1 U9456 ( .A(n8662), .ZN(n7750) );
  INV_X1 U9457 ( .A(n8648), .ZN(n7748) );
  OR2_X1 U9458 ( .A1(n7780), .A2(n7748), .ZN(n8660) );
  INV_X1 U9459 ( .A(n8660), .ZN(n7749) );
  OR2_X1 U9460 ( .A1(n7750), .A2(n7749), .ZN(n8073) );
  AND2_X1 U9461 ( .A1(n8076), .A2(n8073), .ZN(n7752) );
  NAND2_X1 U9462 ( .A1(n7752), .A2(n8670), .ZN(n7751) );
  NAND2_X1 U9463 ( .A1(n7751), .A2(n8667), .ZN(n7754) );
  NAND3_X1 U9464 ( .A1(n7752), .A2(n7743), .A3(n8670), .ZN(n7753) );
  AOI21_X1 U9465 ( .B1(n7754), .B2(n7753), .A(n9081), .ZN(n7755) );
  AOI211_X1 U9466 ( .C1(n8137), .C2(n9231), .A(n7756), .B(n7755), .ZN(n9235)
         );
  AOI21_X1 U9467 ( .B1(n9232), .B2(n7784), .A(n8142), .ZN(n9233) );
  NOR2_X1 U9468 ( .A1(n9088), .A2(n4850), .ZN(n7761) );
  OAI22_X1 U9469 ( .A1(n9144), .A2(n7759), .B1(n8115), .B2(n9124), .ZN(n7760)
         );
  AOI211_X1 U9470 ( .C1(n9233), .C2(n9076), .A(n7761), .B(n7760), .ZN(n7763)
         );
  NAND2_X1 U9471 ( .A1(n9231), .A2(n7880), .ZN(n7762) );
  OAI211_X1 U9472 ( .C1(n9235), .C2(n4407), .A(n7763), .B(n7762), .ZN(P2_U3283) );
  XOR2_X1 U9473 ( .A(n7764), .B(n6564), .Z(n10090) );
  NAND2_X1 U9474 ( .A1(n9711), .A2(n10159), .ZN(n9726) );
  INV_X1 U9475 ( .A(n9726), .ZN(n7771) );
  NAND2_X1 U9476 ( .A1(n9711), .A2(n10161), .ZN(n9731) );
  OAI22_X1 U9477 ( .A1(n7765), .A2(n9731), .B1(n9725), .B2(n7768), .ZN(n7770)
         );
  INV_X1 U9478 ( .A(n10048), .ZN(n7767) );
  INV_X1 U9479 ( .A(n7986), .ZN(n7766) );
  OAI21_X1 U9480 ( .B1(n7768), .B2(n7767), .A(n7766), .ZN(n10085) );
  OAI22_X1 U9481 ( .A1(n9659), .A2(n10085), .B1(n6972), .B2(n9728), .ZN(n7769)
         );
  AOI211_X1 U9482 ( .C1(n7771), .C2(n10082), .A(n7770), .B(n7769), .ZN(n7778)
         );
  NAND2_X1 U9483 ( .A1(n7772), .A2(n6564), .ZN(n7773) );
  NAND2_X1 U9484 ( .A1(n7774), .A2(n7773), .ZN(n7775) );
  NAND2_X1 U9485 ( .A1(n7775), .A2(n10168), .ZN(n10087) );
  MUX2_X1 U9486 ( .A(n10087), .B(n7776), .S(n5064), .Z(n7777) );
  OAI211_X1 U9487 ( .C1(n9738), .C2(n10090), .A(n7778), .B(n7777), .ZN(
        P1_U3289) );
  NAND2_X1 U9488 ( .A1(n7747), .A2(n8657), .ZN(n7779) );
  NAND2_X1 U9489 ( .A1(n7779), .A2(n8648), .ZN(n7946) );
  OR2_X1 U9490 ( .A1(n7946), .A2(n7780), .ZN(n7781) );
  NAND2_X1 U9491 ( .A1(n7781), .A2(n8658), .ZN(n7782) );
  XOR2_X1 U9492 ( .A(n8583), .B(n7782), .Z(n7783) );
  AOI222_X1 U9493 ( .A1(n9138), .A2(n7783), .B1(n8781), .B2(n9120), .C1(n8783), 
        .C2(n9121), .ZN(n9242) );
  INV_X1 U9494 ( .A(n7784), .ZN(n7785) );
  AOI21_X1 U9495 ( .B1(n9238), .B2(n4500), .A(n7785), .ZN(n9240) );
  AOI22_X1 U9496 ( .A1(n4407), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7786), .B2(
        n9143), .ZN(n7787) );
  OAI21_X1 U9497 ( .B1(n7758), .B2(n9088), .A(n7787), .ZN(n7792) );
  INV_X1 U9498 ( .A(n7788), .ZN(n7789) );
  AOI21_X1 U9499 ( .B1(n8583), .B2(n7790), .A(n7789), .ZN(n9243) );
  NOR2_X1 U9500 ( .A1(n9243), .A2(n9114), .ZN(n7791) );
  AOI211_X1 U9501 ( .C1(n9240), .C2(n9076), .A(n7792), .B(n7791), .ZN(n7793)
         );
  OAI21_X1 U9502 ( .B1(n9242), .B2(n4407), .A(n7793), .ZN(P2_U3284) );
  NAND2_X1 U9503 ( .A1(n7795), .A2(n7794), .ZN(n7852) );
  NOR2_X1 U9504 ( .A1(n7795), .A2(n7794), .ZN(n7851) );
  AOI21_X1 U9505 ( .B1(n7796), .B2(n7852), .A(n7851), .ZN(n7800) );
  XNOR2_X1 U9506 ( .A(n7798), .B(n7797), .ZN(n7799) );
  XNOR2_X1 U9507 ( .A(n7800), .B(n7799), .ZN(n7805) );
  OAI22_X1 U9508 ( .A1(n9417), .A2(n5043), .B1(n10139), .B2(n9384), .ZN(n7801)
         );
  AOI211_X1 U9509 ( .C1(n9386), .C2(n9441), .A(n7802), .B(n7801), .ZN(n7804)
         );
  NAND2_X1 U9510 ( .A1(n9410), .A2(n7929), .ZN(n7803) );
  OAI211_X1 U9511 ( .C1(n7805), .C2(n9432), .A(n7804), .B(n7803), .ZN(P1_U3229) );
  AOI22_X1 U9512 ( .A1(n9135), .A2(n7807), .B1(n9148), .B2(n7806), .ZN(n7813)
         );
  OAI22_X1 U9513 ( .A1(n9144), .A2(n7809), .B1(n7808), .B2(n9124), .ZN(n7810)
         );
  AOI21_X1 U9514 ( .B1(n9134), .B2(n7811), .A(n7810), .ZN(n7812) );
  OAI211_X1 U9515 ( .C1(n4407), .C2(n7814), .A(n7813), .B(n7812), .ZN(P2_U3291) );
  AOI211_X1 U9516 ( .C1(n7817), .C2(n7816), .A(n8549), .B(n7815), .ZN(n7823)
         );
  NAND2_X1 U9517 ( .A1(n8545), .A2(n7915), .ZN(n7819) );
  OAI211_X1 U9518 ( .C1(n8553), .C2(n7910), .A(n7819), .B(n7818), .ZN(n7822)
         );
  OAI22_X1 U9519 ( .A1(n7884), .A2(n8543), .B1(n8498), .B2(n7820), .ZN(n7821)
         );
  OR3_X1 U9520 ( .A1(n7823), .A2(n7822), .A3(n7821), .ZN(P2_U3219) );
  INV_X1 U9521 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n7826) );
  XOR2_X1 U9522 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9479), .Z(n7838) );
  INV_X1 U9523 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7828) );
  NAND2_X1 U9524 ( .A1(n10001), .A2(n9488), .ZN(n7827) );
  NAND2_X1 U9525 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9424) );
  OAI211_X1 U9526 ( .C1(n7828), .C2(n10026), .A(n7827), .B(n9424), .ZN(n7837)
         );
  INV_X1 U9527 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7835) );
  NOR2_X1 U9528 ( .A1(n7830), .A2(n7829), .ZN(n7831) );
  AOI21_X1 U9529 ( .B1(n7833), .B2(n7832), .A(n7831), .ZN(n9489) );
  XNOR2_X1 U9530 ( .A(n9489), .B(n9488), .ZN(n7834) );
  NOR2_X1 U9531 ( .A1(n7834), .A2(n7835), .ZN(n9487) );
  AOI211_X1 U9532 ( .C1(n7835), .C2(n7834), .A(n9994), .B(n9487), .ZN(n7836)
         );
  AOI211_X1 U9533 ( .C1(n10003), .C2(n7838), .A(n7837), .B(n7836), .ZN(n7839)
         );
  INV_X1 U9534 ( .A(n7839), .ZN(P1_U3256) );
  AOI21_X1 U9535 ( .B1(n7569), .B2(n8629), .A(n8616), .ZN(n7866) );
  NAND2_X1 U9536 ( .A1(n8638), .A2(n8633), .ZN(n8573) );
  NOR2_X1 U9537 ( .A1(n7866), .A2(n8573), .ZN(n7865) );
  NAND2_X1 U9538 ( .A1(n7848), .A2(n8638), .ZN(n7841) );
  OAI21_X1 U9539 ( .B1(n7865), .B2(n7841), .A(n7840), .ZN(n7842) );
  AOI222_X1 U9540 ( .A1(n9138), .A2(n7842), .B1(n8786), .B2(n9120), .C1(n8788), 
        .C2(n9121), .ZN(n10239) );
  OAI22_X1 U9541 ( .A1(n9144), .A2(n6626), .B1(n7843), .B2(n9124), .ZN(n7846)
         );
  NAND2_X1 U9542 ( .A1(n7873), .A2(n10237), .ZN(n7844) );
  NAND2_X1 U9543 ( .A1(n7890), .A2(n7844), .ZN(n10238) );
  NOR2_X1 U9544 ( .A1(n9021), .A2(n10238), .ZN(n7845) );
  AOI211_X1 U9545 ( .C1(n9134), .C2(n10237), .A(n7846), .B(n7845), .ZN(n7850)
         );
  XNOR2_X1 U9546 ( .A(n7847), .B(n7848), .ZN(n10242) );
  NAND2_X1 U9547 ( .A1(n9135), .A2(n10242), .ZN(n7849) );
  OAI211_X1 U9548 ( .C1(n10239), .C2(n4407), .A(n7850), .B(n7849), .ZN(
        P2_U3289) );
  INV_X1 U9549 ( .A(n7851), .ZN(n7853) );
  NAND2_X1 U9550 ( .A1(n7853), .A2(n7852), .ZN(n7855) );
  XNOR2_X1 U9551 ( .A(n7855), .B(n7854), .ZN(n7861) );
  NAND2_X1 U9552 ( .A1(n9427), .A2(n9442), .ZN(n7857) );
  OAI211_X1 U9553 ( .C1(n9730), .C2(n9425), .A(n7857), .B(n7856), .ZN(n7858)
         );
  AOI21_X1 U9554 ( .B1(n9410), .B2(n8034), .A(n7858), .ZN(n7860) );
  NAND2_X1 U9555 ( .A1(n6949), .A2(n5975), .ZN(n7859) );
  OAI211_X1 U9556 ( .C1(n7861), .C2(n9432), .A(n7860), .B(n7859), .ZN(P1_U3219) );
  NAND2_X1 U9557 ( .A1(n7863), .A2(n7862), .ZN(n7864) );
  XOR2_X1 U9558 ( .A(n8573), .B(n7864), .Z(n10231) );
  AOI21_X1 U9559 ( .B1(n7866), .B2(n8573), .A(n7865), .ZN(n7867) );
  OAI222_X1 U9560 ( .A1(n9102), .A2(n7883), .B1(n9100), .B2(n7868), .C1(n9081), 
        .C2(n7867), .ZN(n10234) );
  INV_X1 U9561 ( .A(n10234), .ZN(n7869) );
  MUX2_X1 U9562 ( .A(n7870), .B(n7869), .S(n9144), .Z(n7878) );
  OR2_X1 U9563 ( .A1(n7871), .A2(n10232), .ZN(n7872) );
  NAND2_X1 U9564 ( .A1(n7873), .A2(n7872), .ZN(n10233) );
  OAI22_X1 U9565 ( .A1(n9021), .A2(n10233), .B1(n7874), .B2(n9124), .ZN(n7875)
         );
  AOI21_X1 U9566 ( .B1(n9134), .B2(n7876), .A(n7875), .ZN(n7877) );
  OAI211_X1 U9567 ( .C1(n10231), .C2(n9114), .A(n7878), .B(n7877), .ZN(
        P2_U3290) );
  INV_X1 U9568 ( .A(n8655), .ZN(n8580) );
  XNOR2_X1 U9569 ( .A(n7879), .B(n8580), .ZN(n10250) );
  INV_X1 U9570 ( .A(n10250), .ZN(n7897) );
  INV_X1 U9571 ( .A(n7880), .ZN(n8151) );
  NAND2_X1 U9572 ( .A1(n10250), .A2(n8137), .ZN(n7888) );
  NAND3_X1 U9573 ( .A1(n7840), .A2(n8580), .A3(n8653), .ZN(n7881) );
  NAND2_X1 U9574 ( .A1(n7882), .A2(n7881), .ZN(n7886) );
  OAI22_X1 U9575 ( .A1(n7884), .A2(n9102), .B1(n7883), .B2(n9100), .ZN(n7885)
         );
  AOI21_X1 U9576 ( .B1(n7886), .B2(n9138), .A(n7885), .ZN(n7887) );
  AND2_X1 U9577 ( .A1(n7888), .A2(n7887), .ZN(n10252) );
  MUX2_X1 U9578 ( .A(n10252), .B(n7889), .S(n4407), .Z(n7896) );
  AND2_X1 U9579 ( .A1(n7890), .A2(n10244), .ZN(n7892) );
  OR2_X1 U9580 ( .A1(n7892), .A2(n7891), .ZN(n10247) );
  OAI22_X1 U9581 ( .A1(n9021), .A2(n10247), .B1(n7893), .B2(n9124), .ZN(n7894)
         );
  AOI21_X1 U9582 ( .B1(n9134), .B2(n10244), .A(n7894), .ZN(n7895) );
  OAI211_X1 U9583 ( .C1(n7897), .C2(n8151), .A(n7896), .B(n7895), .ZN(P2_U3288) );
  NAND2_X1 U9584 ( .A1(n7898), .A2(n9144), .ZN(n7906) );
  OAI22_X1 U9585 ( .A1(n9144), .A2(n7900), .B1(n7899), .B2(n9124), .ZN(n7903)
         );
  NOR2_X1 U9586 ( .A1(n9021), .A2(n7901), .ZN(n7902) );
  AOI211_X1 U9587 ( .C1(n9134), .C2(n7904), .A(n7903), .B(n7902), .ZN(n7905)
         );
  OAI211_X1 U9588 ( .C1(n7907), .C2(n8151), .A(n7906), .B(n7905), .ZN(P2_U3287) );
  INV_X1 U9589 ( .A(n7908), .ZN(n7918) );
  NAND2_X1 U9590 ( .A1(n7909), .A2(n9144), .ZN(n7917) );
  OAI22_X1 U9591 ( .A1(n9144), .A2(n7911), .B1(n7910), .B2(n9124), .ZN(n7914)
         );
  NOR2_X1 U9592 ( .A1(n9021), .A2(n7912), .ZN(n7913) );
  AOI211_X1 U9593 ( .C1(n9134), .C2(n7915), .A(n7914), .B(n7913), .ZN(n7916)
         );
  OAI211_X1 U9594 ( .C1(n7918), .C2(n8151), .A(n7917), .B(n7916), .ZN(P2_U3286) );
  XOR2_X1 U9595 ( .A(n7919), .B(n7924), .Z(n10147) );
  OR2_X1 U9596 ( .A1(n7998), .A2(n7920), .ZN(n8019) );
  NAND2_X1 U9597 ( .A1(n8019), .A2(n7921), .ZN(n8021) );
  NAND2_X1 U9598 ( .A1(n8021), .A2(n7922), .ZN(n7925) );
  OAI211_X1 U9599 ( .C1(n7925), .C2(n7924), .A(n10168), .B(n7923), .ZN(n10145)
         );
  MUX2_X1 U9600 ( .A(n10145), .B(n7926), .S(n5064), .Z(n7934) );
  AOI211_X1 U9601 ( .C1(n10144), .C2(n8026), .A(n10132), .B(n9739), .ZN(n10142) );
  INV_X1 U9602 ( .A(n7927), .ZN(n7928) );
  NAND2_X1 U9603 ( .A1(n7928), .A2(n9568), .ZN(n9691) );
  INV_X1 U9604 ( .A(n7929), .ZN(n7930) );
  OAI22_X1 U9605 ( .A1(n9725), .A2(n5043), .B1(n9728), .B2(n7930), .ZN(n7932)
         );
  OAI22_X1 U9606 ( .A1(n10139), .A2(n9731), .B1(n9726), .B2(n10140), .ZN(n7931) );
  AOI211_X1 U9607 ( .C1(n10142), .C2(n9741), .A(n7932), .B(n7931), .ZN(n7933)
         );
  OAI211_X1 U9608 ( .C1(n9738), .C2(n10147), .A(n7934), .B(n7933), .ZN(
        P1_U3282) );
  NAND2_X1 U9609 ( .A1(n9137), .A2(n8618), .ZN(n10208) );
  INV_X1 U9610 ( .A(n10208), .ZN(n7939) );
  AOI22_X1 U9611 ( .A1(n10208), .A2(n9138), .B1(n9120), .B2(n9122), .ZN(n10210) );
  OAI22_X1 U9612 ( .A1(n4407), .A2(n10210), .B1(n7935), .B2(n9124), .ZN(n7936)
         );
  AOI21_X1 U9613 ( .B1(P2_REG2_REG_0__SCAN_IN), .B2(n4407), .A(n7936), .ZN(
        n7938) );
  OAI21_X1 U9614 ( .B1(n9076), .B2(n9134), .A(n10206), .ZN(n7937) );
  OAI211_X1 U9615 ( .C1(n7939), .C2(n9114), .A(n7938), .B(n7937), .ZN(P2_U3296) );
  INV_X1 U9616 ( .A(n7940), .ZN(n7978) );
  AOI22_X1 U9617 ( .A1(n8765), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n9279), .ZN(n7941) );
  OAI21_X1 U9618 ( .B1(n7978), .B2(n9281), .A(n7941), .ZN(P2_U3336) );
  AOI21_X1 U9619 ( .B1(n7944), .B2(n7943), .A(n7942), .ZN(n7945) );
  XOR2_X1 U9620 ( .A(n8579), .B(n7945), .Z(n9249) );
  XOR2_X1 U9621 ( .A(n8579), .B(n7946), .Z(n7947) );
  AOI222_X1 U9622 ( .A1(n9138), .A2(n7947), .B1(n8782), .B2(n9120), .C1(n8784), 
        .C2(n9121), .ZN(n9248) );
  MUX2_X1 U9623 ( .A(n7948), .B(n9248), .S(n9144), .Z(n7954) );
  XNOR2_X1 U9624 ( .A(n7757), .B(n9245), .ZN(n7949) );
  NOR2_X1 U9625 ( .A1(n7949), .A2(n10246), .ZN(n9244) );
  OAI22_X1 U9626 ( .A1(n9088), .A2(n7951), .B1(n7950), .B2(n9124), .ZN(n7952)
         );
  AOI21_X1 U9627 ( .B1(n9244), .B2(n9148), .A(n7952), .ZN(n7953) );
  OAI211_X1 U9628 ( .C1(n9114), .C2(n9249), .A(n7954), .B(n7953), .ZN(P2_U3285) );
  OAI211_X1 U9629 ( .C1(n7957), .C2(n7956), .A(n7955), .B(n9408), .ZN(n7962)
         );
  NAND2_X1 U9630 ( .A1(n9386), .A2(n9440), .ZN(n7959) );
  OAI211_X1 U9631 ( .C1(n10140), .C2(n9384), .A(n7959), .B(n7958), .ZN(n7960)
         );
  AOI21_X1 U9632 ( .B1(n9410), .B2(n8061), .A(n7960), .ZN(n7961) );
  OAI211_X1 U9633 ( .C1(n8060), .C2(n9417), .A(n7962), .B(n7961), .ZN(P1_U3234) );
  AOI21_X1 U9634 ( .B1(n7965), .B2(n7964), .A(n7963), .ZN(n7977) );
  INV_X1 U9635 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7966) );
  NAND2_X1 U9636 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n8098) );
  OAI21_X1 U9637 ( .B1(n7967), .B2(n7966), .A(n8098), .ZN(n7974) );
  OR3_X1 U9638 ( .A1(n7970), .A2(n7969), .A3(n7968), .ZN(n7971) );
  AOI21_X1 U9639 ( .B1(n7972), .B2(n7971), .A(n8928), .ZN(n7973) );
  AOI211_X1 U9640 ( .C1(n8878), .C2(n7975), .A(n7974), .B(n7973), .ZN(n7976)
         );
  OAI21_X1 U9641 ( .B1(n7977), .B2(n8917), .A(n7976), .ZN(P2_U3259) );
  OAI222_X1 U9642 ( .A1(n4405), .A2(n7979), .B1(n9923), .B2(n7978), .C1(
        P1_U3084), .C2(n6714), .ZN(P1_U3331) );
  NAND2_X1 U9643 ( .A1(n10159), .A2(n9444), .ZN(n7980) );
  OAI21_X1 U9644 ( .B1(n7981), .B2(n10138), .A(n7980), .ZN(n7982) );
  AOI21_X1 U9645 ( .B1(n7983), .B2(n10168), .A(n7982), .ZN(n10098) );
  MUX2_X1 U9646 ( .A(n10098), .B(n7984), .S(n5064), .Z(n7993) );
  XNOR2_X1 U9647 ( .A(n7713), .B(n7985), .ZN(n10101) );
  INV_X1 U9648 ( .A(n9738), .ZN(n9700) );
  NAND2_X1 U9649 ( .A1(n10101), .A2(n9700), .ZN(n7990) );
  OR2_X1 U9650 ( .A1(n7986), .A2(n10096), .ZN(n7987) );
  AND2_X1 U9651 ( .A1(n7988), .A2(n7987), .ZN(n10095) );
  INV_X1 U9652 ( .A(n9728), .ZN(n10067) );
  AOI22_X1 U9653 ( .A1(n9718), .A2(n10095), .B1(n10067), .B2(n5887), .ZN(n7989) );
  OAI211_X1 U9654 ( .C1(n10096), .C2(n9725), .A(n7990), .B(n7989), .ZN(n7991)
         );
  INV_X1 U9655 ( .A(n7991), .ZN(n7992) );
  NAND2_X1 U9656 ( .A1(n7993), .A2(n7992), .ZN(P1_U3288) );
  INV_X1 U9657 ( .A(n7994), .ZN(n7995) );
  NAND2_X1 U9658 ( .A1(n7996), .A2(n7995), .ZN(n7997) );
  XNOR2_X1 U9659 ( .A(n7997), .B(n7999), .ZN(n10171) );
  INV_X1 U9660 ( .A(n7998), .ZN(n8000) );
  OAI21_X1 U9661 ( .B1(n8000), .B2(n7999), .A(n8019), .ZN(n10169) );
  NOR2_X1 U9662 ( .A1(n5064), .A2(n10040), .ZN(n9672) );
  OAI211_X1 U9663 ( .C1(n8002), .C2(n8001), .A(n10117), .B(n8025), .ZN(n10166)
         );
  INV_X1 U9664 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n8004) );
  OAI22_X1 U9665 ( .A1(n9711), .A2(n8004), .B1(n8003), .B2(n9728), .ZN(n8005)
         );
  AOI21_X1 U9666 ( .B1(n9713), .B2(n10162), .A(n8005), .ZN(n8008) );
  OAI22_X1 U9667 ( .A1(n10043), .A2(n9731), .B1(n9726), .B2(n10139), .ZN(n8006) );
  INV_X1 U9668 ( .A(n8006), .ZN(n8007) );
  OAI211_X1 U9669 ( .C1(n10166), .C2(n9691), .A(n8008), .B(n8007), .ZN(n8009)
         );
  AOI21_X1 U9670 ( .B1(n10169), .B2(n9672), .A(n8009), .ZN(n8010) );
  OAI21_X1 U9671 ( .B1(n10171), .B2(n9738), .A(n8010), .ZN(P1_U3284) );
  INV_X1 U9672 ( .A(n8014), .ZN(n8012) );
  AOI21_X1 U9673 ( .B1(P1_DATAO_REG_23__SCAN_IN), .B2(n9279), .A(n8597), .ZN(
        n8011) );
  OAI21_X1 U9674 ( .B1(n8012), .B2(n8366), .A(n8011), .ZN(P2_U3335) );
  NAND2_X1 U9675 ( .A1(n8014), .A2(n8013), .ZN(n8016) );
  OAI211_X1 U9676 ( .C1(n8017), .C2(n4405), .A(n8016), .B(n8015), .ZN(P1_U3330) );
  NAND2_X1 U9677 ( .A1(n8019), .A2(n8018), .ZN(n8020) );
  NAND2_X1 U9678 ( .A1(n8020), .A2(n8032), .ZN(n8022) );
  NAND3_X1 U9679 ( .A1(n8022), .A2(n10168), .A3(n8021), .ZN(n8024) );
  AOI22_X1 U9680 ( .A1(n10161), .A2(n9442), .B1(n10159), .B2(n9959), .ZN(n8023) );
  NAND2_X1 U9681 ( .A1(n8024), .A2(n8023), .ZN(n10136) );
  MUX2_X1 U9682 ( .A(n10136), .B(P1_REG2_REG_8__SCAN_IN), .S(n5064), .Z(n8038)
         );
  INV_X1 U9683 ( .A(n8025), .ZN(n8027) );
  INV_X1 U9684 ( .A(n5975), .ZN(n10131) );
  OAI21_X1 U9685 ( .B1(n8027), .B2(n10131), .A(n8026), .ZN(n10133) );
  OR2_X1 U9686 ( .A1(n7618), .A2(n8028), .ZN(n8030) );
  AND2_X1 U9687 ( .A1(n8030), .A2(n8029), .ZN(n8031) );
  NAND2_X1 U9688 ( .A1(n8031), .A2(n8032), .ZN(n10129) );
  INV_X1 U9689 ( .A(n8031), .ZN(n8033) );
  NAND2_X1 U9690 ( .A1(n8033), .A2(n4562), .ZN(n10127) );
  NAND3_X1 U9691 ( .A1(n10129), .A2(n9700), .A3(n10127), .ZN(n8036) );
  AOI22_X1 U9692 ( .A1(n9713), .A2(n5975), .B1(n8034), .B2(n10067), .ZN(n8035)
         );
  OAI211_X1 U9693 ( .C1(n9659), .C2(n10133), .A(n8036), .B(n8035), .ZN(n8037)
         );
  OR2_X1 U9694 ( .A1(n8038), .A2(n8037), .ZN(P1_U3283) );
  NAND2_X1 U9695 ( .A1(n8039), .A2(n9734), .ZN(n9723) );
  NAND2_X1 U9696 ( .A1(n9723), .A2(n8040), .ZN(n8056) );
  AOI21_X1 U9697 ( .B1(n8056), .B2(n8067), .A(n8041), .ZN(n8043) );
  XNOR2_X1 U9698 ( .A(n8043), .B(n8042), .ZN(n8044) );
  NAND2_X1 U9699 ( .A1(n8044), .A2(n10168), .ZN(n9881) );
  AOI211_X1 U9700 ( .C1(n9880), .C2(n8059), .A(n10132), .B(n4497), .ZN(n9878)
         );
  INV_X1 U9701 ( .A(n9731), .ZN(n9677) );
  INV_X1 U9702 ( .A(n8251), .ZN(n8045) );
  OAI22_X1 U9703 ( .A1(n9711), .A2(n8046), .B1(n8045), .B2(n9728), .ZN(n8047)
         );
  AOI21_X1 U9704 ( .B1(n9677), .B2(n9960), .A(n8047), .ZN(n8049) );
  NAND2_X1 U9705 ( .A1(n9713), .A2(n9880), .ZN(n8048) );
  OAI211_X1 U9706 ( .C1(n9877), .C2(n9726), .A(n8049), .B(n8048), .ZN(n8053)
         );
  OAI21_X1 U9707 ( .B1(n8051), .B2(n6031), .A(n8050), .ZN(n9883) );
  NOR2_X1 U9708 ( .A1(n9883), .A2(n9738), .ZN(n8052) );
  AOI211_X1 U9709 ( .C1(n9878), .C2(n9741), .A(n8053), .B(n8052), .ZN(n8054)
         );
  OAI21_X1 U9710 ( .B1(n5064), .B2(n9881), .A(n8054), .ZN(P1_U3279) );
  XNOR2_X1 U9711 ( .A(n8056), .B(n8055), .ZN(n8057) );
  NAND2_X1 U9712 ( .A1(n8057), .A2(n10168), .ZN(n9890) );
  OAI21_X1 U9713 ( .B1(n8058), .B2(n8060), .A(n8059), .ZN(n9885) );
  INV_X1 U9714 ( .A(n9885), .ZN(n8071) );
  INV_X1 U9715 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n8063) );
  INV_X1 U9716 ( .A(n8061), .ZN(n8062) );
  OAI22_X1 U9717 ( .A1(n9711), .A2(n8063), .B1(n8062), .B2(n9728), .ZN(n8064)
         );
  AOI21_X1 U9718 ( .B1(n9677), .B2(n9441), .A(n8064), .ZN(n8066) );
  NAND2_X1 U9719 ( .A1(n9713), .A2(n9888), .ZN(n8065) );
  OAI211_X1 U9720 ( .C1(n9884), .C2(n9726), .A(n8066), .B(n8065), .ZN(n8070)
         );
  XNOR2_X1 U9721 ( .A(n8068), .B(n8067), .ZN(n9891) );
  NOR2_X1 U9722 ( .A1(n9891), .A2(n9738), .ZN(n8069) );
  AOI211_X1 U9723 ( .C1(n8071), .C2(n9718), .A(n8070), .B(n8069), .ZN(n8072)
         );
  OAI21_X1 U9724 ( .B1(n5064), .B2(n9890), .A(n8072), .ZN(P1_U3280) );
  INV_X1 U9725 ( .A(n8781), .ZN(n8102) );
  NAND2_X1 U9726 ( .A1(n9232), .A2(n8102), .ZN(n8674) );
  AND2_X1 U9727 ( .A1(n8670), .A2(n8674), .ZN(n8074) );
  AND2_X1 U9728 ( .A1(n8074), .A2(n8073), .ZN(n8075) );
  INV_X1 U9729 ( .A(n8674), .ZN(n8077) );
  OR2_X1 U9730 ( .A1(n8077), .A2(n8667), .ZN(n8078) );
  NAND2_X1 U9731 ( .A1(n8079), .A2(n8078), .ZN(n8082) );
  INV_X1 U9732 ( .A(n8082), .ZN(n8080) );
  NAND2_X1 U9733 ( .A1(n9226), .A2(n8112), .ZN(n8678) );
  AOI21_X1 U9734 ( .B1(n8080), .B2(n8129), .A(n9081), .ZN(n8084) );
  OAI22_X1 U9735 ( .A1(n8102), .A2(n9100), .B1(n8155), .B2(n9102), .ZN(n8083)
         );
  AOI21_X1 U9736 ( .B1(n8084), .B2(n8133), .A(n8083), .ZN(n9229) );
  XNOR2_X1 U9737 ( .A(n8142), .B(n9226), .ZN(n9227) );
  INV_X1 U9738 ( .A(n9226), .ZN(n8141) );
  INV_X1 U9739 ( .A(n8099), .ZN(n8085) );
  AOI22_X1 U9740 ( .A1(n4407), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8085), .B2(
        n9143), .ZN(n8086) );
  OAI21_X1 U9741 ( .B1(n8141), .B2(n9088), .A(n8086), .ZN(n8090) );
  NAND2_X1 U9742 ( .A1(n9232), .A2(n8781), .ZN(n8087) );
  NOR2_X1 U9743 ( .A1(n8132), .A2(n8081), .ZN(n8203) );
  AOI21_X1 U9744 ( .B1(n8081), .B2(n8132), .A(n8203), .ZN(n9230) );
  NOR2_X1 U9745 ( .A1(n9230), .A2(n9114), .ZN(n8089) );
  AOI211_X1 U9746 ( .C1(n9227), .C2(n9076), .A(n8090), .B(n8089), .ZN(n8091)
         );
  OAI21_X1 U9747 ( .B1(n4407), .B2(n9229), .A(n8091), .ZN(P2_U3282) );
  NAND2_X1 U9748 ( .A1(n8093), .A2(n8092), .ZN(n8111) );
  NAND2_X1 U9749 ( .A1(n8095), .A2(n8094), .ZN(n8110) );
  NOR2_X1 U9750 ( .A1(n8111), .A2(n8110), .ZN(n8109) );
  NOR3_X1 U9751 ( .A1(n8473), .A2(n8102), .A3(n8096), .ZN(n8097) );
  AOI21_X1 U9752 ( .B1(n8109), .B2(n8457), .A(n8097), .ZN(n8108) );
  INV_X1 U9753 ( .A(n8155), .ZN(n8779) );
  OAI21_X1 U9754 ( .B1(n8553), .B2(n8099), .A(n8098), .ZN(n8100) );
  AOI21_X1 U9755 ( .B1(n8541), .B2(n8779), .A(n8100), .ZN(n8101) );
  OAI21_X1 U9756 ( .B1(n8102), .B2(n8543), .A(n8101), .ZN(n8105) );
  NOR2_X1 U9757 ( .A1(n8103), .A2(n8549), .ZN(n8104) );
  AOI211_X1 U9758 ( .C1(n9226), .C2(n8545), .A(n8105), .B(n8104), .ZN(n8106)
         );
  OAI21_X1 U9759 ( .B1(n8108), .B2(n8107), .A(n8106), .ZN(P2_U3217) );
  AOI211_X1 U9760 ( .C1(n8111), .C2(n8110), .A(n8549), .B(n8109), .ZN(n8119)
         );
  INV_X1 U9761 ( .A(n8112), .ZN(n8780) );
  NAND2_X1 U9762 ( .A1(n8541), .A2(n8780), .ZN(n8114) );
  OAI211_X1 U9763 ( .C1(n8553), .C2(n8115), .A(n8114), .B(n8113), .ZN(n8118)
         );
  OAI22_X1 U9764 ( .A1(n4850), .A2(n8558), .B1(n8543), .B2(n8116), .ZN(n8117)
         );
  OR3_X1 U9765 ( .A1(n8119), .A2(n8118), .A3(n8117), .ZN(P2_U3236) );
  OAI211_X1 U9766 ( .C1(n8121), .C2(n8120), .A(n8210), .B(n8457), .ZN(n8126)
         );
  OR2_X1 U9767 ( .A1(n9101), .A2(n9102), .ZN(n8123) );
  NAND2_X1 U9768 ( .A1(n8778), .A2(n9121), .ZN(n8122) );
  NAND2_X1 U9769 ( .A1(n8123), .A2(n8122), .ZN(n8291) );
  OAI22_X1 U9770 ( .A1(n8553), .A2(n8294), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8906), .ZN(n8124) );
  AOI21_X1 U9771 ( .B1(n8555), .B2(n8291), .A(n8124), .ZN(n8125) );
  OAI211_X1 U9772 ( .C1(n8305), .C2(n8558), .A(n8126), .B(n8125), .ZN(P2_U3230) );
  NOR2_X1 U9773 ( .A1(n8127), .A2(n8155), .ZN(n8685) );
  INV_X1 U9774 ( .A(n8685), .ZN(n8128) );
  NAND2_X1 U9775 ( .A1(n8127), .A2(n8155), .ZN(n8684) );
  NOR2_X1 U9776 ( .A1(n9226), .A2(n8780), .ZN(n8202) );
  NOR2_X1 U9777 ( .A1(n8127), .A2(n8779), .ZN(n8130) );
  AOI21_X1 U9778 ( .B1(n8677), .B2(n8202), .A(n8130), .ZN(n8131) );
  OR2_X1 U9779 ( .A1(n8279), .A2(n8228), .ZN(n8689) );
  NAND2_X1 U9780 ( .A1(n8279), .A2(n8228), .ZN(n8690) );
  XNOR2_X1 U9781 ( .A(n8282), .B(n4916), .ZN(n8138) );
  INV_X1 U9782 ( .A(n8138), .ZN(n8259) );
  OAI21_X1 U9783 ( .B1(n8281), .B2(n8134), .A(n8285), .ZN(n8135) );
  NAND2_X1 U9784 ( .A1(n8135), .A2(n9138), .ZN(n8140) );
  OAI22_X1 U9785 ( .A1(n8283), .A2(n9102), .B1(n8155), .B2(n9100), .ZN(n8136)
         );
  AOI21_X1 U9786 ( .B1(n8138), .B2(n8137), .A(n8136), .ZN(n8139) );
  NAND2_X1 U9787 ( .A1(n8140), .A2(n8139), .ZN(n8261) );
  NAND2_X1 U9788 ( .A1(n8261), .A2(n9144), .ZN(n8150) );
  NAND2_X1 U9789 ( .A1(n8142), .A2(n8141), .ZN(n8199) );
  INV_X1 U9790 ( .A(n8143), .ZN(n8198) );
  AND2_X1 U9791 ( .A1(n8198), .A2(n8279), .ZN(n8144) );
  NOR2_X1 U9792 ( .A1(n5051), .A2(n8144), .ZN(n8257) );
  INV_X1 U9793 ( .A(n8279), .ZN(n8145) );
  NOR2_X1 U9794 ( .A1(n8145), .A2(n9088), .ZN(n8148) );
  OAI22_X1 U9795 ( .A1(n9144), .A2(n8146), .B1(n8164), .B2(n9124), .ZN(n8147)
         );
  AOI211_X1 U9796 ( .C1(n8257), .C2(n9076), .A(n8148), .B(n8147), .ZN(n8149)
         );
  OAI211_X1 U9797 ( .C1(n8259), .C2(n8151), .A(n8150), .B(n8149), .ZN(P2_U3280) );
  INV_X1 U9798 ( .A(n6158), .ZN(n8234) );
  AOI22_X1 U9799 ( .A1(n8152), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n9279), .ZN(n8153) );
  OAI21_X1 U9800 ( .B1(n8234), .B2(n8366), .A(n8153), .ZN(P2_U3334) );
  NAND2_X1 U9801 ( .A1(n8103), .A2(n8154), .ZN(n8157) );
  NOR2_X1 U9802 ( .A1(n8157), .A2(n8156), .ZN(n8221) );
  NOR2_X1 U9803 ( .A1(n8473), .A2(n8155), .ZN(n8222) );
  AOI21_X1 U9804 ( .B1(n8221), .B2(n8457), .A(n8222), .ZN(n8172) );
  NAND2_X1 U9805 ( .A1(n8157), .A2(n8156), .ZN(n8219) );
  XNOR2_X1 U9806 ( .A(n8159), .B(n8158), .ZN(n8162) );
  INV_X1 U9807 ( .A(n8162), .ZN(n8160) );
  NAND2_X1 U9808 ( .A1(n8219), .A2(n8160), .ZN(n8171) );
  OAI21_X1 U9809 ( .B1(n8221), .B2(n8161), .A(n8219), .ZN(n8163) );
  NAND3_X1 U9810 ( .A1(n8163), .A2(n8457), .A3(n8162), .ZN(n8170) );
  NAND2_X1 U9811 ( .A1(n8495), .A2(n8779), .ZN(n8167) );
  INV_X1 U9812 ( .A(n8164), .ZN(n8165) );
  AND2_X1 U9813 ( .A1(P2_U3152), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n8898) );
  AOI21_X1 U9814 ( .B1(n8517), .B2(n8165), .A(n8898), .ZN(n8166) );
  OAI211_X1 U9815 ( .C1(n8283), .C2(n8498), .A(n8167), .B(n8166), .ZN(n8168)
         );
  AOI21_X1 U9816 ( .B1(n8279), .B2(n8545), .A(n8168), .ZN(n8169) );
  OAI211_X1 U9817 ( .C1(n8172), .C2(n8171), .A(n8170), .B(n8169), .ZN(P2_U3228) );
  INV_X1 U9818 ( .A(n8173), .ZN(n8177) );
  AOI21_X1 U9819 ( .B1(n8174), .B2(n8175), .A(n8183), .ZN(n8176) );
  OAI21_X1 U9820 ( .B1(n8177), .B2(n8176), .A(n10168), .ZN(n9874) );
  AOI22_X1 U9821 ( .A1(n5064), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n8243), .B2(
        n10067), .ZN(n8179) );
  NAND2_X1 U9822 ( .A1(n9677), .A2(n9440), .ZN(n8178) );
  OAI211_X1 U9823 ( .C1(n9868), .C2(n9726), .A(n8179), .B(n8178), .ZN(n8181)
         );
  OAI21_X1 U9824 ( .B1(n4497), .B2(n5040), .A(n8188), .ZN(n9869) );
  NOR2_X1 U9825 ( .A1(n9869), .A2(n9659), .ZN(n8180) );
  AOI211_X1 U9826 ( .C1(n9713), .C2(n9872), .A(n8181), .B(n8180), .ZN(n8185)
         );
  XOR2_X1 U9827 ( .A(n8183), .B(n8182), .Z(n9875) );
  OR2_X1 U9828 ( .A1(n9875), .A2(n9738), .ZN(n8184) );
  OAI211_X1 U9829 ( .C1(n9874), .C2(n5064), .A(n8185), .B(n8184), .ZN(P1_U3278) );
  XOR2_X1 U9830 ( .A(n8186), .B(n8192), .Z(n8187) );
  AOI22_X1 U9831 ( .A1(n8187), .A2(n10168), .B1(n10161), .B2(n9439), .ZN(n9866) );
  AOI211_X1 U9832 ( .C1(n9864), .C2(n8188), .A(n10132), .B(n9715), .ZN(n9862)
         );
  NAND2_X1 U9833 ( .A1(n9864), .A2(n9713), .ZN(n8190) );
  AOI22_X1 U9834 ( .A1(n5064), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n9295), .B2(
        n10067), .ZN(n8189) );
  OAI211_X1 U9835 ( .C1(n9861), .C2(n9726), .A(n8190), .B(n8189), .ZN(n8194)
         );
  XNOR2_X1 U9836 ( .A(n8191), .B(n8192), .ZN(n9867) );
  NOR2_X1 U9837 ( .A1(n9867), .A2(n9738), .ZN(n8193) );
  AOI211_X1 U9838 ( .C1(n9741), .C2(n9862), .A(n8194), .B(n8193), .ZN(n8195)
         );
  OAI21_X1 U9839 ( .B1(n9866), .B2(n5064), .A(n8195), .ZN(P1_U3277) );
  XNOR2_X1 U9840 ( .A(n8196), .B(n8677), .ZN(n8197) );
  AOI222_X1 U9841 ( .A1(n9138), .A2(n8197), .B1(n8778), .B2(n9120), .C1(n8780), 
        .C2(n9121), .ZN(n9224) );
  AOI21_X1 U9842 ( .B1(n8127), .B2(n8199), .A(n8143), .ZN(n9222) );
  INV_X1 U9843 ( .A(n8127), .ZN(n8201) );
  AOI22_X1 U9844 ( .A1(n4407), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8225), .B2(
        n9143), .ZN(n8200) );
  OAI21_X1 U9845 ( .B1(n8201), .B2(n9088), .A(n8200), .ZN(n8206) );
  NOR2_X1 U9846 ( .A1(n8203), .A2(n8202), .ZN(n8204) );
  XNOR2_X1 U9847 ( .A(n8204), .B(n8677), .ZN(n9225) );
  NOR2_X1 U9848 ( .A1(n9225), .A2(n9114), .ZN(n8205) );
  AOI211_X1 U9849 ( .C1(n9222), .C2(n9076), .A(n8206), .B(n8205), .ZN(n8207)
         );
  OAI21_X1 U9850 ( .B1(n4407), .B2(n9224), .A(n8207), .ZN(P2_U3281) );
  INV_X1 U9851 ( .A(n9218), .ZN(n8323) );
  INV_X1 U9852 ( .A(n8208), .ZN(n8209) );
  AOI21_X1 U9853 ( .B1(n8210), .B2(n8209), .A(n8549), .ZN(n8214) );
  NOR3_X1 U9854 ( .A1(n8211), .A2(n8283), .A3(n8473), .ZN(n8213) );
  OAI21_X1 U9855 ( .B1(n8214), .B2(n8213), .A(n8212), .ZN(n8218) );
  INV_X1 U9856 ( .A(n8283), .ZN(n8777) );
  AOI22_X1 U9857 ( .A1(n8517), .A2(n8321), .B1(P2_REG3_REG_18__SCAN_IN), .B2(
        P2_U3152), .ZN(n8215) );
  OAI21_X1 U9858 ( .B1(n8498), .B2(n8524), .A(n8215), .ZN(n8216) );
  AOI21_X1 U9859 ( .B1(n8495), .B2(n8777), .A(n8216), .ZN(n8217) );
  OAI211_X1 U9860 ( .C1(n8323), .C2(n8558), .A(n8218), .B(n8217), .ZN(P2_U3240) );
  INV_X1 U9861 ( .A(n8219), .ZN(n8220) );
  NOR2_X1 U9862 ( .A1(n8221), .A2(n8220), .ZN(n8233) );
  INV_X1 U9863 ( .A(n8222), .ZN(n8232) );
  NAND3_X1 U9864 ( .A1(n8233), .A2(n8457), .A3(n8223), .ZN(n8231) );
  NAND2_X1 U9865 ( .A1(n8495), .A2(n8780), .ZN(n8227) );
  NOR2_X1 U9866 ( .A1(n8224), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8272) );
  AOI21_X1 U9867 ( .B1(n8517), .B2(n8225), .A(n8272), .ZN(n8226) );
  OAI211_X1 U9868 ( .C1(n8228), .C2(n8498), .A(n8227), .B(n8226), .ZN(n8229)
         );
  AOI21_X1 U9869 ( .B1(n8127), .B2(n8545), .A(n8229), .ZN(n8230) );
  OAI211_X1 U9870 ( .C1(n8233), .C2(n8232), .A(n8231), .B(n8230), .ZN(P2_U3243) );
  OAI222_X1 U9871 ( .A1(P1_U3084), .A2(n8235), .B1(n9923), .B2(n8234), .C1(
        n10566), .C2(n4405), .ZN(P1_U3329) );
  OR2_X1 U9872 ( .A1(n8249), .A2(n8250), .ZN(n8247) );
  NAND2_X1 U9873 ( .A1(n8247), .A2(n8236), .ZN(n8240) );
  XNOR2_X1 U9874 ( .A(n8238), .B(n8237), .ZN(n8239) );
  XNOR2_X1 U9875 ( .A(n8240), .B(n8239), .ZN(n8246) );
  NAND2_X1 U9876 ( .A1(n9427), .A2(n9440), .ZN(n8241) );
  NAND2_X1 U9877 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9972) );
  OAI211_X1 U9878 ( .C1(n9868), .C2(n9425), .A(n8241), .B(n9972), .ZN(n8242)
         );
  AOI21_X1 U9879 ( .B1(n9410), .B2(n8243), .A(n8242), .ZN(n8245) );
  NAND2_X1 U9880 ( .A1(n9872), .A2(n6949), .ZN(n8244) );
  OAI211_X1 U9881 ( .C1(n8246), .C2(n9432), .A(n8245), .B(n8244), .ZN(P1_U3232) );
  INV_X1 U9882 ( .A(n8247), .ZN(n8248) );
  AOI21_X1 U9883 ( .B1(n8250), .B2(n8249), .A(n8248), .ZN(n8256) );
  NAND2_X1 U9884 ( .A1(n9410), .A2(n8251), .ZN(n8253) );
  AOI22_X1 U9885 ( .A1(n9386), .A2(n9439), .B1(P1_REG3_REG_12__SCAN_IN), .B2(
        P1_U3084), .ZN(n8252) );
  OAI211_X1 U9886 ( .C1(n9876), .C2(n9384), .A(n8253), .B(n8252), .ZN(n8254)
         );
  AOI21_X1 U9887 ( .B1(n6949), .B2(n9880), .A(n8254), .ZN(n8255) );
  OAI21_X1 U9888 ( .B1(n8256), .B2(n9432), .A(n8255), .ZN(P1_U3222) );
  AOI22_X1 U9889 ( .A1(n8257), .A2(n9239), .B1(n9246), .B2(n8279), .ZN(n8258)
         );
  OAI21_X1 U9890 ( .B1(n8259), .B2(n9237), .A(n8258), .ZN(n8260) );
  NOR2_X1 U9891 ( .A1(n8261), .A2(n8260), .ZN(n8264) );
  MUX2_X1 U9892 ( .A(n8262), .B(n8264), .S(n10263), .Z(n8263) );
  INV_X1 U9893 ( .A(n8263), .ZN(P2_U3536) );
  INV_X1 U9894 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8265) );
  MUX2_X1 U9895 ( .A(n8265), .B(n8264), .S(n10254), .Z(n8266) );
  INV_X1 U9896 ( .A(n8266), .ZN(P2_U3499) );
  INV_X1 U9897 ( .A(n8267), .ZN(n8314) );
  AOI22_X1 U9898 ( .A1(n8268), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_25__SCAN_IN), .B2(n9279), .ZN(n8269) );
  OAI21_X1 U9899 ( .B1(n8314), .B2(n8366), .A(n8269), .ZN(P2_U3333) );
  XNOR2_X1 U9900 ( .A(n8270), .B(n5524), .ZN(n8278) );
  XNOR2_X1 U9901 ( .A(n8271), .B(P2_REG1_REG_15__SCAN_IN), .ZN(n8276) );
  AOI21_X1 U9902 ( .B1(n8922), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n8272), .ZN(
        n8273) );
  OAI21_X1 U9903 ( .B1(n8932), .B2(n8274), .A(n8273), .ZN(n8275) );
  AOI21_X1 U9904 ( .B1(n8276), .B2(n8811), .A(n8275), .ZN(n8277) );
  OAI21_X1 U9905 ( .B1(n8278), .B2(n8917), .A(n8277), .ZN(P2_U3260) );
  NAND2_X1 U9906 ( .A1(n8279), .A2(n8778), .ZN(n8280) );
  NAND2_X1 U9907 ( .A1(n8324), .A2(n8283), .ZN(n8694) );
  NAND2_X1 U9908 ( .A1(n8693), .A2(n8694), .ZN(n8688) );
  OAI21_X1 U9909 ( .B1(n8284), .B2(n8688), .A(n8326), .ZN(n8302) );
  INV_X1 U9910 ( .A(n8302), .ZN(n8301) );
  NAND2_X1 U9911 ( .A1(n8285), .A2(n8690), .ZN(n8286) );
  NAND2_X1 U9912 ( .A1(n8286), .A2(n8688), .ZN(n8290) );
  INV_X1 U9913 ( .A(n8690), .ZN(n8287) );
  NOR2_X1 U9914 ( .A1(n8688), .A2(n8287), .ZN(n8288) );
  NAND2_X1 U9915 ( .A1(n8289), .A2(n8288), .ZN(n8316) );
  NAND3_X1 U9916 ( .A1(n8290), .A2(n9138), .A3(n8316), .ZN(n8293) );
  INV_X1 U9917 ( .A(n8291), .ZN(n8292) );
  NAND2_X1 U9918 ( .A1(n8293), .A2(n8292), .ZN(n8307) );
  NAND2_X1 U9919 ( .A1(n8307), .A2(n9144), .ZN(n8300) );
  INV_X1 U9920 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8295) );
  OAI22_X1 U9921 ( .A1(n9144), .A2(n8295), .B1(n8294), .B2(n9124), .ZN(n8298)
         );
  AND2_X2 U9922 ( .A1(n5051), .A2(n8305), .ZN(n8319) );
  OAI21_X1 U9923 ( .B1(n5051), .B2(n8305), .A(n9239), .ZN(n8296) );
  OR2_X1 U9924 ( .A1(n8319), .A2(n8296), .ZN(n8303) );
  INV_X1 U9925 ( .A(n9148), .ZN(n9109) );
  NOR2_X1 U9926 ( .A1(n8303), .A2(n9109), .ZN(n8297) );
  AOI211_X1 U9927 ( .C1(n9134), .C2(n8324), .A(n8298), .B(n8297), .ZN(n8299)
         );
  OAI211_X1 U9928 ( .C1(n9114), .C2(n8301), .A(n8300), .B(n8299), .ZN(P2_U3279) );
  INV_X1 U9929 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8308) );
  NAND2_X1 U9930 ( .A1(n8302), .A2(n10243), .ZN(n8304) );
  OAI211_X1 U9931 ( .C1(n8305), .C2(n10245), .A(n8304), .B(n8303), .ZN(n8306)
         );
  NOR2_X1 U9932 ( .A1(n8307), .A2(n8306), .ZN(n8310) );
  MUX2_X1 U9933 ( .A(n8308), .B(n8310), .S(n10254), .Z(n8309) );
  INV_X1 U9934 ( .A(n8309), .ZN(P2_U3502) );
  MUX2_X1 U9935 ( .A(n8311), .B(n8310), .S(n10263), .Z(n8312) );
  INV_X1 U9936 ( .A(n8312), .ZN(P2_U3537) );
  OAI222_X1 U9937 ( .A1(n4405), .A2(n8315), .B1(n9923), .B2(n8314), .C1(
        P1_U3084), .C2(n8313), .ZN(P1_U3328) );
  OR2_X1 U9938 ( .A1(n9218), .A2(n9101), .ZN(n8701) );
  NAND2_X1 U9939 ( .A1(n9218), .A2(n9101), .ZN(n8699) );
  OAI21_X1 U9940 ( .B1(n8317), .B2(n5057), .A(n8436), .ZN(n8318) );
  INV_X1 U9941 ( .A(n8524), .ZN(n8775) );
  AOI222_X1 U9942 ( .A1(n9138), .A2(n8318), .B1(n8775), .B2(n9120), .C1(n8777), 
        .C2(n9121), .ZN(n9220) );
  INV_X1 U9943 ( .A(n8319), .ZN(n8320) );
  AOI211_X1 U9944 ( .C1(n9218), .C2(n8320), .A(n10246), .B(n4845), .ZN(n9217)
         );
  AOI22_X1 U9945 ( .A1(n4407), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8321), .B2(
        n9143), .ZN(n8322) );
  OAI21_X1 U9946 ( .B1(n8323), .B2(n9088), .A(n8322), .ZN(n8328) );
  OR2_X1 U9947 ( .A1(n8324), .A2(n8777), .ZN(n8325) );
  XNOR2_X1 U9948 ( .A(n8418), .B(n5057), .ZN(n9221) );
  NOR2_X1 U9949 ( .A1(n9221), .A2(n9114), .ZN(n8327) );
  AOI211_X1 U9950 ( .C1(n9217), .C2(n9148), .A(n8328), .B(n8327), .ZN(n8329)
         );
  OAI21_X1 U9951 ( .B1(n9220), .B2(n4407), .A(n8329), .ZN(P2_U3278) );
  INV_X1 U9952 ( .A(n8330), .ZN(n8334) );
  AOI22_X1 U9953 ( .A1(n8331), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n9279), .ZN(n8332) );
  OAI21_X1 U9954 ( .B1(n8334), .B2(n8366), .A(n8332), .ZN(P2_U3332) );
  OAI222_X1 U9955 ( .A1(P1_U3084), .A2(n8335), .B1(n9923), .B2(n8334), .C1(
        n8333), .C2(n4405), .ZN(P1_U3327) );
  INV_X1 U9956 ( .A(n8336), .ZN(n8414) );
  AOI22_X1 U9957 ( .A1(n8762), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n9279), .ZN(n8337) );
  OAI21_X1 U9958 ( .B1(n8414), .B2(n8366), .A(n8337), .ZN(P2_U3331) );
  INV_X1 U9959 ( .A(n6223), .ZN(n9922) );
  NAND2_X1 U9960 ( .A1(n9279), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n8338) );
  OAI211_X1 U9961 ( .C1(n9922), .C2(n9281), .A(n8339), .B(n8338), .ZN(P2_U3330) );
  XNOR2_X1 U9962 ( .A(n8340), .B(n6568), .ZN(n9775) );
  AOI211_X1 U9963 ( .C1(n8342), .C2(n6568), .A(n10040), .B(n8341), .ZN(n8344)
         );
  OAI22_X1 U9964 ( .A1(n9520), .A2(n10141), .B1(n9548), .B2(n10138), .ZN(n8343) );
  NOR2_X1 U9965 ( .A1(n8344), .A2(n8343), .ZN(n9774) );
  INV_X1 U9966 ( .A(n9774), .ZN(n8353) );
  NOR2_X1 U9967 ( .A1(n9770), .A2(n4447), .ZN(n8346) );
  OR2_X1 U9968 ( .A1(n8346), .A2(n8345), .ZN(n9771) );
  OAI22_X1 U9969 ( .A1(n8348), .A2(n9728), .B1(n8347), .B2(n9711), .ZN(n8349)
         );
  AOI21_X1 U9970 ( .B1(n8350), .B2(n9713), .A(n8349), .ZN(n8351) );
  OAI21_X1 U9971 ( .B1(n9771), .B2(n9659), .A(n8351), .ZN(n8352) );
  AOI21_X1 U9972 ( .B1(n8353), .B2(n9711), .A(n8352), .ZN(n8354) );
  OAI21_X1 U9973 ( .B1(n9775), .B2(n9738), .A(n8354), .ZN(P1_U3264) );
  XOR2_X1 U9974 ( .A(n8360), .B(n8355), .Z(n9780) );
  INV_X1 U9975 ( .A(n9544), .ZN(n8358) );
  AOI21_X1 U9976 ( .B1(n9776), .B2(n8358), .A(n4447), .ZN(n9777) );
  AOI22_X1 U9977 ( .A1(n9411), .A2(n10067), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n5064), .ZN(n8359) );
  OAI21_X1 U9978 ( .B1(n9418), .B2(n9725), .A(n8359), .ZN(n8362) );
  OAI21_X1 U9979 ( .B1(n9780), .B2(n9738), .A(n4488), .ZN(P1_U3265) );
  OAI222_X1 U9980 ( .A1(P1_U3084), .A2(n8364), .B1(n4405), .B2(n8363), .C1(
        n9921), .C2(n8365), .ZN(P1_U3352) );
  OAI222_X1 U9981 ( .A1(P2_U3152), .A2(n8369), .B1(n8368), .B2(n8367), .C1(
        n8366), .C2(n8365), .ZN(P2_U3357) );
  NOR2_X1 U9982 ( .A1(n8372), .A2(n8371), .ZN(n8370) );
  AOI21_X1 U9983 ( .B1(n8372), .B2(n8371), .A(n8370), .ZN(n8379) );
  AOI22_X1 U9984 ( .A1(n8545), .A2(n9133), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n8373), .ZN(n8378) );
  NAND2_X1 U9985 ( .A1(n8791), .A2(n9120), .ZN(n8376) );
  NAND2_X1 U9986 ( .A1(n8374), .A2(n9121), .ZN(n8375) );
  NAND2_X1 U9987 ( .A1(n8376), .A2(n8375), .ZN(n9140) );
  NAND2_X1 U9988 ( .A1(n8555), .A2(n9140), .ZN(n8377) );
  OAI211_X1 U9989 ( .C1(n8379), .C2(n8549), .A(n8378), .B(n8377), .ZN(P2_U3224) );
  INV_X1 U9990 ( .A(n9545), .ZN(n9786) );
  INV_X1 U9991 ( .A(n8380), .ZN(n9302) );
  NAND2_X1 U9992 ( .A1(n8382), .A2(n8381), .ZN(n9300) );
  OR2_X1 U9993 ( .A1(n8383), .A2(n8386), .ZN(n9350) );
  NOR2_X1 U9994 ( .A1(n9351), .A2(n9350), .ZN(n9349) );
  INV_X1 U9995 ( .A(n8384), .ZN(n8385) );
  NOR3_X1 U9996 ( .A1(n9349), .A2(n8386), .A3(n8385), .ZN(n8387) );
  OAI21_X1 U9997 ( .B1(n8387), .B2(n9406), .A(n9408), .ZN(n8392) );
  OAI22_X1 U9998 ( .A1(n9547), .A2(n9384), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8388), .ZN(n8390) );
  NOR2_X1 U9999 ( .A1(n9548), .A2(n9425), .ZN(n8389) );
  AOI211_X1 U10000 ( .C1(n9410), .C2(n9551), .A(n8390), .B(n8389), .ZN(n8391)
         );
  OAI211_X1 U10001 ( .C1(n9786), .C2(n9417), .A(n8392), .B(n8391), .ZN(
        P1_U3223) );
  INV_X1 U10002 ( .A(n9201), .ZN(n9071) );
  OR2_X2 U10003 ( .A1(n9030), .A2(n9192), .ZN(n9031) );
  NOR2_X4 U10004 ( .A1(n9031), .A2(n8428), .ZN(n9015) );
  NAND2_X1 U10005 ( .A1(n8412), .A2(n8398), .ZN(n8395) );
  NAND2_X1 U10006 ( .A1(n4408), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n8394) );
  NAND2_X1 U10007 ( .A1(n9275), .A2(n8398), .ZN(n8397) );
  NAND2_X1 U10008 ( .A1(n4408), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n8396) );
  NAND2_X1 U10009 ( .A1(n8935), .A2(n9160), .ZN(n9157) );
  NAND2_X1 U10010 ( .A1(n4408), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n8399) );
  INV_X1 U10011 ( .A(n8561), .ZN(n8564) );
  INV_X1 U10012 ( .A(P2_B_REG_SCAN_IN), .ZN(n8400) );
  OAI21_X1 U10013 ( .B1(n8401), .B2(n8400), .A(n9120), .ZN(n8446) );
  NOR2_X1 U10014 ( .A1(n8564), .A2(n8446), .ZN(n9152) );
  INV_X1 U10015 ( .A(n9152), .ZN(n9158) );
  NOR2_X1 U10016 ( .A1(n4407), .A2(n9158), .ZN(n8938) );
  NOR2_X1 U10017 ( .A1(n8562), .A2(n9088), .ZN(n8402) );
  AOI211_X1 U10018 ( .C1(n4407), .C2(P2_REG2_REG_31__SCAN_IN), .A(n8938), .B(
        n8402), .ZN(n8403) );
  OAI21_X1 U10019 ( .B1(n9155), .B2(n9021), .A(n8403), .ZN(P2_U3265) );
  AOI22_X1 U10020 ( .A1(n8405), .A2(n10067), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n5064), .ZN(n8407) );
  NAND2_X1 U10021 ( .A1(n9515), .A2(n9713), .ZN(n8406) );
  OAI211_X1 U10022 ( .C1(n8408), .C2(n9691), .A(n8407), .B(n8406), .ZN(n8409)
         );
  AOI21_X1 U10023 ( .B1(n8410), .B2(n9711), .A(n8409), .ZN(n8411) );
  OAI21_X1 U10024 ( .B1(n8404), .B2(n9738), .A(n8411), .ZN(P1_U3263) );
  INV_X1 U10025 ( .A(n8412), .ZN(n9282) );
  OAI222_X1 U10026 ( .A1(n4405), .A2(n10444), .B1(n9921), .B2(n9282), .C1(
        n8413), .C2(P1_U3084), .ZN(P1_U3324) );
  OAI222_X1 U10027 ( .A1(n4405), .A2(n8415), .B1(P1_U3084), .B2(n9504), .C1(
        n8414), .C2(n9921), .ZN(P1_U3326) );
  INV_X1 U10028 ( .A(n9101), .ZN(n8776) );
  NOR2_X1 U10029 ( .A1(n9218), .A2(n8776), .ZN(n8417) );
  NAND2_X1 U10030 ( .A1(n9218), .A2(n8776), .ZN(n8416) );
  AND2_X1 U10031 ( .A1(n9211), .A2(n8775), .ZN(n8419) );
  NAND2_X1 U10032 ( .A1(n9207), .A2(n9103), .ZN(n8717) );
  INV_X1 U10033 ( .A(n9103), .ZN(n9065) );
  NAND2_X1 U10034 ( .A1(n9207), .A2(n9065), .ZN(n8420) );
  INV_X1 U10035 ( .A(n9047), .ZN(n8774) );
  OR2_X1 U10036 ( .A1(n9201), .A2(n8774), .ZN(n8422) );
  AND2_X1 U10037 ( .A1(n9201), .A2(n8774), .ZN(n8421) );
  INV_X1 U10038 ( .A(n8423), .ZN(n8539) );
  INV_X1 U10039 ( .A(n9066), .ZN(n8499) );
  NAND2_X1 U10040 ( .A1(n8539), .A2(n8499), .ZN(n8437) );
  NAND2_X1 U10041 ( .A1(n8710), .A2(n8437), .ZN(n9057) );
  XNOR2_X1 U10042 ( .A(n9192), .B(n9048), .ZN(n9038) );
  INV_X1 U10043 ( .A(n8424), .ZN(n8425) );
  NOR2_X1 U10044 ( .A1(n8505), .A2(n8425), .ZN(n8427) );
  NAND2_X1 U10045 ( .A1(n8428), .A2(n8505), .ZN(n8727) );
  AND2_X1 U10046 ( .A1(n8726), .A2(n8727), .ZN(n8725) );
  NAND2_X1 U10047 ( .A1(n9182), .A2(n9012), .ZN(n8603) );
  NAND2_X1 U10048 ( .A1(n8605), .A2(n8603), .ZN(n8996) );
  NAND2_X1 U10049 ( .A1(n8990), .A2(n8996), .ZN(n8989) );
  INV_X1 U10050 ( .A(n9182), .ZN(n8429) );
  INV_X1 U10051 ( .A(n9012), .ZN(n8772) );
  NAND2_X1 U10052 ( .A1(n8429), .A2(n9012), .ZN(n8430) );
  NAND2_X1 U10053 ( .A1(n9177), .A2(n8964), .ZN(n8731) );
  INV_X1 U10054 ( .A(n8735), .ZN(n8770) );
  NAND2_X1 U10055 ( .A1(n9168), .A2(n8965), .ZN(n8432) );
  NAND2_X2 U10056 ( .A1(n8740), .A2(n8432), .ZN(n8945) );
  INV_X1 U10057 ( .A(n8965), .ZN(n8769) );
  NAND2_X1 U10058 ( .A1(n4855), .A2(n8965), .ZN(n8433) );
  OR2_X1 U10059 ( .A1(n9162), .A2(n8434), .ZN(n8747) );
  NAND2_X1 U10060 ( .A1(n9162), .A2(n8434), .ZN(n8748) );
  NAND2_X1 U10061 ( .A1(n9211), .A2(n8524), .ZN(n8700) );
  NAND2_X1 U10062 ( .A1(n9079), .A2(n9078), .ZN(n9004) );
  OR2_X1 U10063 ( .A1(n9201), .A2(n9047), .ZN(n8704) );
  NAND2_X1 U10064 ( .A1(n8704), .A2(n9005), .ZN(n8716) );
  AOI211_X1 U10065 ( .C1(n9036), .C2(n9008), .A(n8716), .B(n9007), .ZN(n8442)
         );
  NAND2_X1 U10066 ( .A1(n9201), .A2(n9047), .ZN(n9044) );
  NAND2_X1 U10067 ( .A1(n8437), .A2(n9044), .ZN(n8719) );
  NAND3_X1 U10068 ( .A1(n8719), .A2(n9048), .A3(n8710), .ZN(n8440) );
  INV_X1 U10069 ( .A(n8437), .ZN(n8706) );
  OAI22_X1 U10070 ( .A1(n8710), .A2(n9048), .B1(n8438), .B2(n8706), .ZN(n8439)
         );
  AOI21_X1 U10071 ( .B1(n9036), .B2(n8440), .A(n8439), .ZN(n8441) );
  NAND2_X1 U10072 ( .A1(n8726), .A2(n8727), .ZN(n9010) );
  INV_X1 U10073 ( .A(n8726), .ZN(n8443) );
  INV_X1 U10074 ( .A(n8605), .ZN(n8444) );
  INV_X1 U10075 ( .A(n8730), .ZN(n8445) );
  NOR2_X1 U10076 ( .A1(n9172), .A2(n8735), .ZN(n8739) );
  XNOR2_X1 U10077 ( .A(n8559), .B(n8742), .ZN(n8448) );
  OAI22_X1 U10078 ( .A1(n8965), .A2(n9100), .B1(n8563), .B2(n8446), .ZN(n8447)
         );
  INV_X1 U10079 ( .A(n9164), .ZN(n8449) );
  NAND2_X1 U10080 ( .A1(n8449), .A2(n9144), .ZN(n8456) );
  AOI211_X1 U10081 ( .C1(n9162), .C2(n8947), .A(n10246), .B(n8935), .ZN(n9161)
         );
  INV_X1 U10082 ( .A(n9162), .ZN(n8450) );
  NOR2_X1 U10083 ( .A1(n8450), .A2(n9088), .ZN(n8454) );
  OAI22_X1 U10084 ( .A1(n9144), .A2(n8452), .B1(n8451), .B2(n9124), .ZN(n8453)
         );
  OAI211_X1 U10085 ( .C1(n9165), .C2(n9114), .A(n8456), .B(n8455), .ZN(
        P2_U3267) );
  NAND3_X1 U10086 ( .A1(n8459), .A2(n8535), .A3(n8771), .ZN(n8460) );
  AOI22_X1 U10087 ( .A1(n8959), .A2(n8517), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8462) );
  OAI21_X1 U10088 ( .B1(n8965), .B2(n8498), .A(n8462), .ZN(n8463) );
  AOI21_X1 U10089 ( .B1(n8495), .B2(n8771), .A(n8463), .ZN(n8464) );
  OAI211_X1 U10090 ( .C1(n4857), .C2(n8558), .A(n8465), .B(n8464), .ZN(
        P2_U3216) );
  OAI22_X1 U10091 ( .A1(n8553), .A2(n9033), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10329), .ZN(n8466) );
  AOI21_X1 U10092 ( .B1(n8495), .B2(n9066), .A(n8466), .ZN(n8467) );
  OAI21_X1 U10093 ( .B1(n8505), .B2(n8498), .A(n8467), .ZN(n8475) );
  INV_X1 U10094 ( .A(n8468), .ZN(n8469) );
  NAND2_X1 U10095 ( .A1(n8470), .A2(n8469), .ZN(n8472) );
  XNOR2_X1 U10096 ( .A(n8472), .B(n8471), .ZN(n8477) );
  NOR3_X1 U10097 ( .A1(n8477), .A2(n9048), .A3(n8473), .ZN(n8474) );
  AOI211_X1 U10098 ( .C1(n9192), .C2(n8545), .A(n8475), .B(n8474), .ZN(n8479)
         );
  NAND3_X1 U10099 ( .A1(n8477), .A2(n8457), .A3(n8476), .ZN(n8478) );
  NAND2_X1 U10100 ( .A1(n8479), .A2(n8478), .ZN(P2_U3218) );
  OAI22_X1 U10101 ( .A1(n8553), .A2(n9107), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10538), .ZN(n8480) );
  AOI21_X1 U10102 ( .B1(n8495), .B2(n8776), .A(n8480), .ZN(n8481) );
  OAI21_X1 U10103 ( .B1(n9103), .B2(n8498), .A(n8481), .ZN(n8491) );
  INV_X1 U10104 ( .A(n8486), .ZN(n8483) );
  NOR3_X1 U10105 ( .A1(n8483), .A2(n8482), .A3(n8549), .ZN(n8489) );
  NAND3_X1 U10106 ( .A1(n8484), .A2(n8535), .A3(n8775), .ZN(n8485) );
  OAI21_X1 U10107 ( .B1(n8486), .B2(n8549), .A(n8485), .ZN(n8488) );
  MUX2_X1 U10108 ( .A(n8489), .B(n8488), .S(n8487), .Z(n8490) );
  AOI211_X1 U10109 ( .C1(n9211), .C2(n8545), .A(n8491), .B(n8490), .ZN(n8492)
         );
  INV_X1 U10110 ( .A(n8492), .ZN(P2_U3221) );
  XNOR2_X1 U10111 ( .A(n8493), .B(n8494), .ZN(n8502) );
  NAND2_X1 U10112 ( .A1(n8495), .A2(n9065), .ZN(n8497) );
  AOI22_X1 U10113 ( .A1(n8517), .A2(n9069), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8496) );
  OAI211_X1 U10114 ( .C1(n8499), .C2(n8498), .A(n8497), .B(n8496), .ZN(n8500)
         );
  AOI21_X1 U10115 ( .B1(n9201), .B2(n8545), .A(n8500), .ZN(n8501) );
  OAI21_X1 U10116 ( .B1(n8502), .B2(n8549), .A(n8501), .ZN(P2_U3225) );
  XNOR2_X1 U10117 ( .A(n4670), .B(n8503), .ZN(n8504) );
  XNOR2_X1 U10118 ( .A(n4871), .B(n8504), .ZN(n8511) );
  OAI22_X1 U10119 ( .A1(n8964), .A2(n9102), .B1(n8505), .B2(n9100), .ZN(n8998)
         );
  INV_X1 U10120 ( .A(n8993), .ZN(n8507) );
  OAI22_X1 U10121 ( .A1(n8553), .A2(n8507), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8506), .ZN(n8509) );
  NOR2_X1 U10122 ( .A1(n8429), .A2(n8558), .ZN(n8508) );
  AOI211_X1 U10123 ( .C1(n8555), .C2(n8998), .A(n8509), .B(n8508), .ZN(n8510)
         );
  OAI21_X1 U10124 ( .B1(n8511), .B2(n8549), .A(n8510), .ZN(P2_U3227) );
  INV_X1 U10125 ( .A(n8428), .ZN(n9186) );
  NAND2_X1 U10126 ( .A1(n8535), .A2(n9028), .ZN(n8515) );
  OR2_X1 U10127 ( .A1(n8549), .A2(n8512), .ZN(n8514) );
  MUX2_X1 U10128 ( .A(n8515), .B(n8514), .S(n8513), .Z(n8521) );
  INV_X1 U10129 ( .A(n9017), .ZN(n8516) );
  AOI22_X1 U10130 ( .A1(n8517), .A2(n8516), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8518) );
  OAI21_X1 U10131 ( .B1(n8543), .B2(n9048), .A(n8518), .ZN(n8519) );
  AOI21_X1 U10132 ( .B1(n8541), .B2(n8772), .A(n8519), .ZN(n8520) );
  OAI211_X1 U10133 ( .C1(n9186), .C2(n8558), .A(n8521), .B(n8520), .ZN(
        P2_U3231) );
  XNOR2_X1 U10134 ( .A(n8523), .B(n8522), .ZN(n8530) );
  OAI22_X1 U10135 ( .A1(n9047), .A2(n9102), .B1(n8524), .B2(n9100), .ZN(n9083)
         );
  INV_X1 U10136 ( .A(n9086), .ZN(n8526) );
  OAI22_X1 U10137 ( .A1(n8553), .A2(n8526), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8525), .ZN(n8528) );
  NOR2_X1 U10138 ( .A1(n4849), .A2(n8558), .ZN(n8527) );
  AOI211_X1 U10139 ( .C1(n8555), .C2(n9083), .A(n8528), .B(n8527), .ZN(n8529)
         );
  OAI21_X1 U10140 ( .B1(n8530), .B2(n8549), .A(n8529), .ZN(P2_U3235) );
  NAND2_X1 U10141 ( .A1(n8532), .A2(n8531), .ZN(n8534) );
  XNOR2_X1 U10142 ( .A(n8534), .B(n8533), .ZN(n8536) );
  NAND3_X1 U10143 ( .A1(n8536), .A2(n8535), .A3(n9066), .ZN(n8548) );
  INV_X1 U10144 ( .A(n8536), .ZN(n8538) );
  NAND3_X1 U10145 ( .A1(n8538), .A2(n8457), .A3(n8537), .ZN(n8547) );
  OAI22_X1 U10146 ( .A1(n8553), .A2(n9054), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10296), .ZN(n8540) );
  AOI21_X1 U10147 ( .B1(n8541), .B2(n9008), .A(n8540), .ZN(n8542) );
  OAI21_X1 U10148 ( .B1(n9047), .B2(n8543), .A(n8542), .ZN(n8544) );
  AOI21_X1 U10149 ( .B1(n8539), .B2(n8545), .A(n8544), .ZN(n8546) );
  NAND3_X1 U10150 ( .A1(n8548), .A2(n8547), .A3(n8546), .ZN(P2_U3237) );
  OR2_X1 U10151 ( .A1(n8735), .A2(n9102), .ZN(n8552) );
  OR2_X1 U10152 ( .A1(n9012), .A2(n9100), .ZN(n8551) );
  NAND2_X1 U10153 ( .A1(n8552), .A2(n8551), .ZN(n8984) );
  OAI22_X1 U10154 ( .A1(n8553), .A2(n8978), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10562), .ZN(n8554) );
  AOI21_X1 U10155 ( .B1(n8984), .B2(n8555), .A(n8554), .ZN(n8556) );
  OAI211_X1 U10156 ( .C1(n8981), .C2(n8558), .A(n8557), .B(n8556), .ZN(
        P2_U3242) );
  NOR2_X1 U10157 ( .A1(n8561), .A2(n8600), .ZN(n8560) );
  OR2_X1 U10158 ( .A1(n8936), .A2(n8563), .ZN(n8750) );
  NAND2_X1 U10159 ( .A1(n8562), .A2(n8561), .ZN(n8756) );
  NAND2_X1 U10160 ( .A1(n8936), .A2(n8563), .ZN(n8751) );
  NAND2_X1 U10161 ( .A1(n8756), .A2(n8751), .ZN(n8569) );
  XNOR2_X1 U10162 ( .A(n8565), .B(n8591), .ZN(n8768) );
  INV_X1 U10163 ( .A(n8566), .ZN(n8567) );
  OAI21_X1 U10164 ( .B1(n8568), .B2(n8567), .A(n8597), .ZN(n8767) );
  INV_X1 U10165 ( .A(n8982), .ZN(n8588) );
  INV_X1 U10166 ( .A(n8996), .ZN(n8729) );
  NAND2_X1 U10167 ( .A1(n8704), .A2(n9044), .ZN(n9073) );
  NOR2_X1 U10168 ( .A1(n9136), .A2(n9115), .ZN(n8572) );
  NAND4_X1 U10169 ( .A1(n8572), .A2(n8758), .A3(n8571), .A4(n8614), .ZN(n8574)
         );
  NOR4_X1 U10170 ( .A1(n8575), .A2(n8574), .A3(n8573), .A4(n10208), .ZN(n8577)
         );
  NAND3_X1 U10171 ( .A1(n8577), .A2(n8639), .A3(n8576), .ZN(n8581) );
  NOR4_X1 U10172 ( .A1(n8581), .A2(n8580), .A3(n8579), .A4(n8578), .ZN(n8582)
         );
  NAND4_X1 U10173 ( .A1(n8081), .A2(n8583), .A3(n8582), .A4(n8667), .ZN(n8584)
         );
  NOR4_X1 U10174 ( .A1(n4916), .A2(n8688), .A3(n8677), .A4(n8584), .ZN(n8585)
         );
  NAND4_X1 U10175 ( .A1(n9078), .A2(n5057), .A3(n9096), .A4(n8585), .ZN(n8586)
         );
  NOR4_X1 U10176 ( .A1(n9010), .A2(n9057), .A3(n9073), .A4(n8586), .ZN(n8587)
         );
  INV_X1 U10177 ( .A(n9038), .ZN(n9026) );
  NAND4_X1 U10178 ( .A1(n8588), .A2(n8729), .A3(n8587), .A4(n9026), .ZN(n8589)
         );
  NOR4_X1 U10179 ( .A1(n8742), .A2(n8945), .A3(n8963), .A4(n8589), .ZN(n8590)
         );
  INV_X1 U10180 ( .A(n8599), .ZN(n8757) );
  XNOR2_X1 U10181 ( .A(n8592), .B(n8591), .ZN(n8593) );
  OAI22_X1 U10182 ( .A1(n8593), .A2(n8608), .B1(n8758), .B2(n8596), .ZN(n8594)
         );
  NAND3_X1 U10183 ( .A1(n8597), .A2(n8596), .A3(n8595), .ZN(n8760) );
  INV_X1 U10184 ( .A(n8750), .ZN(n8598) );
  NOR2_X1 U10185 ( .A1(n8599), .A2(n8598), .ZN(n8602) );
  NOR2_X1 U10186 ( .A1(n8600), .A2(n5122), .ZN(n8601) );
  MUX2_X1 U10187 ( .A(n8602), .B(n4941), .S(n8746), .Z(n8754) );
  INV_X1 U10188 ( .A(n8603), .ZN(n8604) );
  OR2_X1 U10189 ( .A1(n8982), .A2(n8604), .ZN(n8607) );
  NAND2_X1 U10190 ( .A1(n8730), .A2(n8605), .ZN(n8606) );
  MUX2_X1 U10191 ( .A(n8607), .B(n8606), .S(n8746), .Z(n8734) );
  AND2_X1 U10192 ( .A1(n8618), .A2(n8608), .ZN(n8612) );
  AND2_X1 U10193 ( .A1(n8610), .A2(n8609), .ZN(n8622) );
  NAND3_X1 U10194 ( .A1(n8613), .A2(n7273), .A3(n8755), .ZN(n8615) );
  NOR2_X1 U10195 ( .A1(n8616), .A2(n8625), .ZN(n8617) );
  INV_X1 U10196 ( .A(n8618), .ZN(n8620) );
  NAND2_X1 U10197 ( .A1(n8620), .A2(n8619), .ZN(n8621) );
  NAND2_X1 U10198 ( .A1(n8622), .A2(n8621), .ZN(n8623) );
  INV_X1 U10199 ( .A(n8627), .ZN(n8631) );
  NAND2_X1 U10200 ( .A1(n8629), .A2(n8628), .ZN(n8630) );
  OAI21_X1 U10201 ( .B1(n8632), .B2(n8631), .A(n8630), .ZN(n8634) );
  NAND2_X1 U10202 ( .A1(n8634), .A2(n8633), .ZN(n8635) );
  NAND2_X1 U10203 ( .A1(n8635), .A2(n8746), .ZN(n8636) );
  NAND2_X1 U10204 ( .A1(n8637), .A2(n8636), .ZN(n8640) );
  NAND2_X1 U10205 ( .A1(n8640), .A2(n5063), .ZN(n8656) );
  NAND3_X1 U10206 ( .A1(n8656), .A2(n8655), .A3(n8641), .ZN(n8643) );
  NAND2_X1 U10207 ( .A1(n8643), .A2(n8642), .ZN(n8646) );
  NAND2_X1 U10208 ( .A1(n8644), .A2(n8650), .ZN(n8645) );
  INV_X1 U10209 ( .A(n8647), .ZN(n8652) );
  AND2_X1 U10210 ( .A1(n8648), .A2(n8647), .ZN(n8649) );
  MUX2_X1 U10211 ( .A(n8650), .B(n8649), .S(n8755), .Z(n8651) );
  AND2_X1 U10212 ( .A1(n8651), .A2(n8657), .ZN(n8654) );
  NAND4_X1 U10213 ( .A1(n8656), .A2(n8655), .A3(n8654), .A4(n8653), .ZN(n8659)
         );
  NAND3_X1 U10214 ( .A1(n8659), .A2(n8658), .A3(n8657), .ZN(n8661) );
  NAND2_X1 U10215 ( .A1(n8663), .A2(n8670), .ZN(n8664) );
  NAND2_X1 U10216 ( .A1(n8664), .A2(n8746), .ZN(n8668) );
  NAND2_X1 U10217 ( .A1(n8781), .A2(n8746), .ZN(n8665) );
  NOR2_X1 U10218 ( .A1(n9232), .A2(n8665), .ZN(n8666) );
  AOI21_X1 U10219 ( .B1(n8668), .B2(n8667), .A(n8666), .ZN(n8676) );
  NAND3_X1 U10220 ( .A1(n8671), .A2(n8670), .A3(n8669), .ZN(n8673) );
  AOI21_X1 U10221 ( .B1(n8673), .B2(n8672), .A(n8746), .ZN(n8675) );
  OAI22_X1 U10222 ( .A1(n8676), .A2(n8675), .B1(n8746), .B2(n8674), .ZN(n8683)
         );
  INV_X1 U10223 ( .A(n8677), .ZN(n8681) );
  MUX2_X1 U10224 ( .A(n8679), .B(n8678), .S(n8755), .Z(n8680) );
  NAND2_X1 U10225 ( .A1(n8681), .A2(n8680), .ZN(n8682) );
  AOI21_X1 U10226 ( .B1(n8683), .B2(n8081), .A(n8682), .ZN(n8687) );
  MUX2_X1 U10227 ( .A(n8685), .B(n4919), .S(n8746), .Z(n8686) );
  INV_X1 U10228 ( .A(n8688), .ZN(n8692) );
  MUX2_X1 U10229 ( .A(n8690), .B(n8689), .S(n8746), .Z(n8691) );
  NAND2_X1 U10230 ( .A1(n8701), .A2(n8693), .ZN(n8696) );
  INV_X1 U10231 ( .A(n8694), .ZN(n8695) );
  MUX2_X1 U10232 ( .A(n8696), .B(n8695), .S(n8746), .Z(n8697) );
  INV_X1 U10233 ( .A(n8697), .ZN(n8698) );
  NAND2_X1 U10234 ( .A1(n8700), .A2(n8699), .ZN(n8711) );
  NAND2_X1 U10235 ( .A1(n9005), .A2(n8714), .ZN(n8702) );
  OAI211_X1 U10236 ( .C1(n8703), .C2(n8702), .A(n8717), .B(n9044), .ZN(n8708)
         );
  INV_X1 U10237 ( .A(n8704), .ZN(n8705) );
  NOR2_X1 U10238 ( .A1(n9007), .A2(n8705), .ZN(n8707) );
  AOI21_X1 U10239 ( .B1(n8708), .B2(n8707), .A(n8706), .ZN(n8709) );
  INV_X1 U10240 ( .A(n8711), .ZN(n8712) );
  NAND2_X1 U10241 ( .A1(n8713), .A2(n8712), .ZN(n8715) );
  NAND2_X1 U10242 ( .A1(n8715), .A2(n8714), .ZN(n8718) );
  AOI21_X1 U10243 ( .B1(n8718), .B2(n8717), .A(n8716), .ZN(n8720) );
  NAND2_X1 U10244 ( .A1(n9048), .A2(n8755), .ZN(n8723) );
  NAND2_X1 U10245 ( .A1(n9008), .A2(n8746), .ZN(n8722) );
  MUX2_X1 U10246 ( .A(n8723), .B(n8722), .S(n9036), .Z(n8724) );
  MUX2_X1 U10247 ( .A(n8727), .B(n8726), .S(n8755), .Z(n8728) );
  MUX2_X1 U10248 ( .A(n8731), .B(n8730), .S(n8755), .Z(n8732) );
  OAI211_X1 U10249 ( .C1(n8734), .C2(n8733), .A(n4647), .B(n8732), .ZN(n8738)
         );
  AND2_X1 U10250 ( .A1(n9172), .A2(n8735), .ZN(n8736) );
  OAI21_X1 U10251 ( .B1(n8945), .B2(n8736), .A(n8755), .ZN(n8737) );
  INV_X1 U10252 ( .A(n8739), .ZN(n8741) );
  AOI21_X1 U10253 ( .B1(n8741), .B2(n8740), .A(n8755), .ZN(n8744) );
  NAND3_X1 U10254 ( .A1(n9168), .A2(n8965), .A3(n8746), .ZN(n8743) );
  OAI211_X1 U10255 ( .C1(n8745), .C2(n8744), .A(n4937), .B(n8743), .ZN(n8752)
         );
  MUX2_X1 U10256 ( .A(n8748), .B(n8747), .S(n8746), .Z(n8749) );
  NAND4_X1 U10257 ( .A1(n8752), .A2(n8751), .A3(n8750), .A4(n8749), .ZN(n8753)
         );
  MUX2_X1 U10258 ( .A(n8757), .B(n8756), .S(n8755), .Z(n8759) );
  NAND4_X1 U10259 ( .A1(n10178), .A2(n9121), .A3(n8762), .A4(n8761), .ZN(n8763) );
  OAI211_X1 U10260 ( .C1(n8765), .C2(n8764), .A(n8763), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8766) );
  MUX2_X1 U10261 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8769), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U10262 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8770), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10263 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8771), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U10264 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8772), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U10265 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9028), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U10266 ( .A(n9008), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8773), .Z(
        P2_U3575) );
  MUX2_X1 U10267 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9066), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10268 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8774), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10269 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n9065), .S(P2_U3966), .Z(
        P2_U3572) );
  MUX2_X1 U10270 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8775), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10271 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n8776), .S(P2_U3966), .Z(
        P2_U3570) );
  MUX2_X1 U10272 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8777), .S(P2_U3966), .Z(
        P2_U3569) );
  MUX2_X1 U10273 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8778), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10274 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8779), .S(P2_U3966), .Z(
        P2_U3567) );
  MUX2_X1 U10275 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n8780), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10276 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8781), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10277 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8782), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U10278 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n8783), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10279 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n8784), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10280 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n8785), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10281 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8786), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U10282 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8787), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U10283 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8788), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U10284 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8789), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U10285 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n8790), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U10286 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n7343), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U10287 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8791), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U10288 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n9122), .S(P2_U3966), .Z(
        P2_U3553) );
  OAI211_X1 U10289 ( .C1(n8794), .C2(n8793), .A(n8874), .B(n8792), .ZN(n8801)
         );
  AOI22_X1 U10290 ( .A1(n8922), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n8800) );
  NAND2_X1 U10291 ( .A1(n8878), .A2(n8795), .ZN(n8799) );
  MUX2_X1 U10292 ( .A(n6651), .B(P2_REG1_REG_1__SCAN_IN), .S(n8795), .Z(n8796)
         );
  OAI21_X1 U10293 ( .B1(n7240), .B2(n5134), .A(n8796), .ZN(n8797) );
  NAND3_X1 U10294 ( .A1(n8811), .A2(n8807), .A3(n8797), .ZN(n8798) );
  NAND4_X1 U10295 ( .A1(n8801), .A2(n8800), .A3(n8799), .A4(n8798), .ZN(
        P2_U3246) );
  OAI211_X1 U10296 ( .C1(n8804), .C2(n8803), .A(n8874), .B(n8802), .ZN(n8815)
         );
  AOI22_X1 U10297 ( .A1(n8922), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n8814) );
  NAND2_X1 U10298 ( .A1(n8878), .A2(n8805), .ZN(n8813) );
  MUX2_X1 U10299 ( .A(n6650), .B(P2_REG1_REG_2__SCAN_IN), .S(n8805), .Z(n8808)
         );
  NAND3_X1 U10300 ( .A1(n8808), .A2(n8807), .A3(n8806), .ZN(n8809) );
  NAND3_X1 U10301 ( .A1(n8811), .A2(n8810), .A3(n8809), .ZN(n8812) );
  NAND4_X1 U10302 ( .A1(n8815), .A2(n8814), .A3(n8813), .A4(n8812), .ZN(
        P2_U3247) );
  OAI211_X1 U10303 ( .C1(n8818), .C2(n8817), .A(n8874), .B(n8816), .ZN(n8828)
         );
  NOR2_X1 U10304 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8819), .ZN(n8820) );
  AOI21_X1 U10305 ( .B1(n8922), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n8820), .ZN(
        n8827) );
  NAND2_X1 U10306 ( .A1(n8878), .A2(n8821), .ZN(n8826) );
  OAI21_X1 U10307 ( .B1(n8823), .B2(n8822), .A(n8837), .ZN(n8824) );
  OR2_X1 U10308 ( .A1(n8928), .A2(n8824), .ZN(n8825) );
  NAND4_X1 U10309 ( .A1(n8828), .A2(n8827), .A3(n8826), .A4(n8825), .ZN(
        P2_U3248) );
  OAI211_X1 U10310 ( .C1(n8831), .C2(n8830), .A(n8874), .B(n8829), .ZN(n8844)
         );
  INV_X1 U10311 ( .A(n8832), .ZN(n8833) );
  AOI21_X1 U10312 ( .B1(n8922), .B2(P2_ADDR_REG_4__SCAN_IN), .A(n8833), .ZN(
        n8843) );
  NAND2_X1 U10313 ( .A1(n8878), .A2(n8834), .ZN(n8842) );
  MUX2_X1 U10314 ( .A(n6658), .B(P2_REG1_REG_4__SCAN_IN), .S(n8834), .Z(n8835)
         );
  NAND3_X1 U10315 ( .A1(n8837), .A2(n8836), .A3(n8835), .ZN(n8838) );
  NAND2_X1 U10316 ( .A1(n8839), .A2(n8838), .ZN(n8840) );
  OR2_X1 U10317 ( .A1(n8928), .A2(n8840), .ZN(n8841) );
  NAND4_X1 U10318 ( .A1(n8844), .A2(n8843), .A3(n8842), .A4(n8841), .ZN(
        P2_U3249) );
  OAI211_X1 U10319 ( .C1(n8847), .C2(n8846), .A(n8874), .B(n8845), .ZN(n8858)
         );
  AOI21_X1 U10320 ( .B1(n8922), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8848), .ZN(
        n8857) );
  NAND2_X1 U10321 ( .A1(n8878), .A2(n8849), .ZN(n8856) );
  MUX2_X1 U10322 ( .A(n6664), .B(P2_REG1_REG_6__SCAN_IN), .S(n8849), .Z(n8850)
         );
  NAND3_X1 U10323 ( .A1(n8852), .A2(n8851), .A3(n8850), .ZN(n8853) );
  NAND2_X1 U10324 ( .A1(n8866), .A2(n8853), .ZN(n8854) );
  OR2_X1 U10325 ( .A1(n8928), .A2(n8854), .ZN(n8855) );
  NAND4_X1 U10326 ( .A1(n8858), .A2(n8857), .A3(n8856), .A4(n8855), .ZN(
        P2_U3251) );
  OAI211_X1 U10327 ( .C1(n8861), .C2(n8860), .A(n8874), .B(n8859), .ZN(n8872)
         );
  NOR2_X1 U10328 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5298), .ZN(n8862) );
  AOI21_X1 U10329 ( .B1(n8922), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8862), .ZN(
        n8871) );
  NAND2_X1 U10330 ( .A1(n8878), .A2(n8863), .ZN(n8870) );
  MUX2_X1 U10331 ( .A(n6667), .B(P2_REG1_REG_7__SCAN_IN), .S(n8863), .Z(n8864)
         );
  NAND3_X1 U10332 ( .A1(n8866), .A2(n8865), .A3(n8864), .ZN(n8867) );
  NAND2_X1 U10333 ( .A1(n8882), .A2(n8867), .ZN(n8868) );
  OR2_X1 U10334 ( .A1(n8928), .A2(n8868), .ZN(n8869) );
  NAND4_X1 U10335 ( .A1(n8872), .A2(n8871), .A3(n8870), .A4(n8869), .ZN(
        P2_U3252) );
  OAI211_X1 U10336 ( .C1(n8876), .C2(n8875), .A(n8874), .B(n8873), .ZN(n8889)
         );
  INV_X1 U10337 ( .A(n8877), .ZN(n10424) );
  AOI21_X1 U10338 ( .B1(n8922), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n10424), .ZN(
        n8888) );
  NAND2_X1 U10339 ( .A1(n8878), .A2(n8879), .ZN(n8887) );
  MUX2_X1 U10340 ( .A(n6670), .B(P2_REG1_REG_8__SCAN_IN), .S(n8879), .Z(n8880)
         );
  NAND3_X1 U10341 ( .A1(n8882), .A2(n8881), .A3(n8880), .ZN(n8883) );
  NAND2_X1 U10342 ( .A1(n8884), .A2(n8883), .ZN(n8885) );
  OR2_X1 U10343 ( .A1(n8928), .A2(n8885), .ZN(n8886) );
  NAND4_X1 U10344 ( .A1(n8889), .A2(n8888), .A3(n8887), .A4(n8886), .ZN(
        P2_U3253) );
  AOI21_X1 U10345 ( .B1(n8892), .B2(n8891), .A(n8890), .ZN(n8901) );
  AOI211_X1 U10346 ( .C1(n8894), .C2(n8893), .A(n4455), .B(n8917), .ZN(n8895)
         );
  INV_X1 U10347 ( .A(n8895), .ZN(n8900) );
  NOR2_X1 U10348 ( .A1(n8932), .A2(n8896), .ZN(n8897) );
  AOI211_X1 U10349 ( .C1(P2_ADDR_REG_16__SCAN_IN), .C2(n8922), .A(n8898), .B(
        n8897), .ZN(n8899) );
  OAI211_X1 U10350 ( .C1(n8901), .C2(n8928), .A(n8900), .B(n8899), .ZN(
        P2_U3261) );
  AOI211_X1 U10351 ( .C1(n8904), .C2(n8903), .A(n8902), .B(n8917), .ZN(n8916)
         );
  INV_X1 U10352 ( .A(n8905), .ZN(n8914) );
  NOR2_X1 U10353 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8906), .ZN(n8907) );
  AOI21_X1 U10354 ( .B1(n8922), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8907), .ZN(
        n8913) );
  OAI21_X1 U10355 ( .B1(n8910), .B2(n8909), .A(n8908), .ZN(n8911) );
  OR2_X1 U10356 ( .A1(n8928), .A2(n8911), .ZN(n8912) );
  OAI211_X1 U10357 ( .C1(n8932), .C2(n8914), .A(n8913), .B(n8912), .ZN(n8915)
         );
  OR2_X1 U10358 ( .A1(n8916), .A2(n8915), .ZN(P2_U3262) );
  AOI211_X1 U10359 ( .C1(n8920), .C2(n8919), .A(n8918), .B(n8917), .ZN(n8934)
         );
  NOR2_X1 U10360 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5566), .ZN(n8921) );
  AOI21_X1 U10361 ( .B1(n8922), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n8921), .ZN(
        n8930) );
  OAI21_X1 U10362 ( .B1(n8925), .B2(n8924), .A(n8923), .ZN(n8926) );
  INV_X1 U10363 ( .A(n8926), .ZN(n8927) );
  OR2_X1 U10364 ( .A1(n8928), .A2(n8927), .ZN(n8929) );
  OAI211_X1 U10365 ( .C1(n8932), .C2(n8931), .A(n8930), .B(n8929), .ZN(n8933)
         );
  OR2_X1 U10366 ( .A1(n8934), .A2(n8933), .ZN(P2_U3263) );
  INV_X1 U10367 ( .A(n8935), .ZN(n8937) );
  NAND2_X1 U10368 ( .A1(n8937), .A2(n8936), .ZN(n9156) );
  NAND3_X1 U10369 ( .A1(n9157), .A2(n9076), .A3(n9156), .ZN(n8940) );
  AOI21_X1 U10370 ( .B1(n4407), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8938), .ZN(
        n8939) );
  OAI211_X1 U10371 ( .C1(n9160), .C2(n9088), .A(n8940), .B(n8939), .ZN(
        P2_U3266) );
  XOR2_X1 U10372 ( .A(n8941), .B(n8945), .Z(n8943) );
  OAI21_X1 U10373 ( .B1(n8946), .B2(n8945), .A(n8944), .ZN(n9166) );
  AOI21_X1 U10374 ( .B1(n9168), .B2(n8957), .A(n10246), .ZN(n8948) );
  AND2_X1 U10375 ( .A1(n8948), .A2(n8947), .ZN(n9167) );
  NAND2_X1 U10376 ( .A1(n9167), .A2(n9148), .ZN(n8951) );
  AOI22_X1 U10377 ( .A1(n4407), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8949), .B2(
        n9143), .ZN(n8950) );
  OAI211_X1 U10378 ( .C1(n4855), .C2(n9088), .A(n8951), .B(n8950), .ZN(n8952)
         );
  AOI21_X1 U10379 ( .B1(n9166), .B2(n9135), .A(n8952), .ZN(n8953) );
  OAI21_X1 U10380 ( .B1(n9170), .B2(n4407), .A(n8953), .ZN(P2_U3268) );
  OAI21_X1 U10381 ( .B1(n8955), .B2(n8963), .A(n8954), .ZN(n8956) );
  INV_X1 U10382 ( .A(n8956), .ZN(n9175) );
  INV_X1 U10383 ( .A(n8957), .ZN(n8958) );
  AOI211_X1 U10384 ( .C1(n9172), .C2(n8975), .A(n10246), .B(n8958), .ZN(n9171)
         );
  AOI22_X1 U10385 ( .A1(n4407), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8959), .B2(
        n9143), .ZN(n8960) );
  OAI21_X1 U10386 ( .B1(n4857), .B2(n9088), .A(n8960), .ZN(n8969) );
  AOI211_X1 U10387 ( .C1(n8963), .C2(n8962), .A(n9081), .B(n8961), .ZN(n8967)
         );
  OAI22_X1 U10388 ( .A1(n8965), .A2(n9102), .B1(n8964), .B2(n9100), .ZN(n8966)
         );
  NOR2_X1 U10389 ( .A1(n8967), .A2(n8966), .ZN(n9174) );
  NOR2_X1 U10390 ( .A1(n9174), .A2(n4407), .ZN(n8968) );
  AOI211_X1 U10391 ( .C1(n9171), .C2(n9148), .A(n8969), .B(n8968), .ZN(n8970)
         );
  OAI21_X1 U10392 ( .B1(n9175), .B2(n9114), .A(n8970), .ZN(P2_U3269) );
  OAI21_X1 U10393 ( .B1(n8972), .B2(n8982), .A(n8971), .ZN(n8973) );
  INV_X1 U10394 ( .A(n8973), .ZN(n9180) );
  INV_X1 U10395 ( .A(n8974), .ZN(n8977) );
  INV_X1 U10396 ( .A(n8975), .ZN(n8976) );
  AOI211_X1 U10397 ( .C1(n9177), .C2(n8977), .A(n10246), .B(n8976), .ZN(n9176)
         );
  INV_X1 U10398 ( .A(n8978), .ZN(n8979) );
  AOI22_X1 U10399 ( .A1(n4407), .A2(P2_REG2_REG_26__SCAN_IN), .B1(n8979), .B2(
        n9143), .ZN(n8980) );
  OAI21_X1 U10400 ( .B1(n8981), .B2(n9088), .A(n8980), .ZN(n8987) );
  AOI211_X1 U10401 ( .C1(n8983), .C2(n8982), .A(n9081), .B(n4453), .ZN(n8985)
         );
  NOR2_X1 U10402 ( .A1(n8985), .A2(n8984), .ZN(n9179) );
  NOR2_X1 U10403 ( .A1(n9179), .A2(n4407), .ZN(n8986) );
  AOI211_X1 U10404 ( .C1(n9176), .C2(n9148), .A(n8987), .B(n8986), .ZN(n8988)
         );
  OAI21_X1 U10405 ( .B1(n9180), .B2(n9114), .A(n8988), .ZN(P2_U3270) );
  OAI21_X1 U10406 ( .B1(n8990), .B2(n8996), .A(n8989), .ZN(n8991) );
  INV_X1 U10407 ( .A(n8991), .ZN(n9185) );
  INV_X1 U10408 ( .A(n9015), .ZN(n8992) );
  AOI211_X1 U10409 ( .C1(n9182), .C2(n8992), .A(n10246), .B(n8974), .ZN(n9181)
         );
  AOI22_X1 U10410 ( .A1(n4407), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8993), .B2(
        n9143), .ZN(n8994) );
  OAI21_X1 U10411 ( .B1(n8429), .B2(n9088), .A(n8994), .ZN(n9001) );
  AOI211_X1 U10412 ( .C1(n8997), .C2(n8996), .A(n9081), .B(n8995), .ZN(n8999)
         );
  NOR2_X1 U10413 ( .A1(n8999), .A2(n8998), .ZN(n9184) );
  NOR2_X1 U10414 ( .A1(n9184), .A2(n4407), .ZN(n9000) );
  AOI211_X1 U10415 ( .C1(n9148), .C2(n9181), .A(n9001), .B(n9000), .ZN(n9002)
         );
  OAI21_X1 U10416 ( .B1(n9185), .B2(n9114), .A(n9002), .ZN(P2_U3271) );
  XNOR2_X1 U10417 ( .A(n9003), .B(n9010), .ZN(n9191) );
  INV_X1 U10418 ( .A(n9005), .ZN(n9062) );
  NOR3_X1 U10419 ( .A1(n9080), .A2(n9062), .A3(n9073), .ZN(n9043) );
  INV_X1 U10420 ( .A(n9044), .ZN(n9006) );
  NOR2_X1 U10421 ( .A1(n9045), .A2(n9007), .ZN(n9027) );
  OAI21_X1 U10422 ( .B1(n9036), .B2(n9008), .A(n9025), .ZN(n9011) );
  AOI211_X1 U10423 ( .C1(n9011), .C2(n9010), .A(n9009), .B(n9081), .ZN(n9014)
         );
  OAI22_X1 U10424 ( .A1(n9012), .A2(n9102), .B1(n9048), .B2(n9100), .ZN(n9013)
         );
  NOR2_X1 U10425 ( .A1(n9014), .A2(n9013), .ZN(n9190) );
  INV_X1 U10426 ( .A(n9190), .ZN(n9023) );
  AND2_X1 U10427 ( .A1(n9031), .A2(n8428), .ZN(n9016) );
  OR2_X1 U10428 ( .A1(n9016), .A2(n9015), .ZN(n9187) );
  INV_X1 U10429 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n9018) );
  OAI22_X1 U10430 ( .A1(n9144), .A2(n9018), .B1(n9017), .B2(n9124), .ZN(n9019)
         );
  AOI21_X1 U10431 ( .B1(n8428), .B2(n9134), .A(n9019), .ZN(n9020) );
  OAI21_X1 U10432 ( .B1(n9187), .B2(n9021), .A(n9020), .ZN(n9022) );
  AOI21_X1 U10433 ( .B1(n9023), .B2(n9144), .A(n9022), .ZN(n9024) );
  OAI21_X1 U10434 ( .B1(n9114), .B2(n9191), .A(n9024), .ZN(P2_U3272) );
  OAI21_X1 U10435 ( .B1(n9027), .B2(n9026), .A(n9025), .ZN(n9029) );
  AOI222_X1 U10436 ( .A1(n9138), .A2(n9029), .B1(n9028), .B2(n9120), .C1(n9066), .C2(n9121), .ZN(n9195) );
  INV_X1 U10437 ( .A(n9031), .ZN(n9032) );
  AOI21_X1 U10438 ( .B1(n9192), .B2(n9030), .A(n9032), .ZN(n9193) );
  INV_X1 U10439 ( .A(n9033), .ZN(n9034) );
  AOI22_X1 U10440 ( .A1(n4407), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9034), .B2(
        n9143), .ZN(n9035) );
  OAI21_X1 U10441 ( .B1(n9036), .B2(n9088), .A(n9035), .ZN(n9041) );
  OAI21_X1 U10442 ( .B1(n9039), .B2(n9038), .A(n9037), .ZN(n9196) );
  NOR2_X1 U10443 ( .A1(n9196), .A2(n9114), .ZN(n9040) );
  AOI211_X1 U10444 ( .C1(n9193), .C2(n9076), .A(n9041), .B(n9040), .ZN(n9042)
         );
  OAI21_X1 U10445 ( .B1(n4409), .B2(n4407), .A(n9042), .ZN(P2_U3273) );
  INV_X1 U10446 ( .A(n9043), .ZN(n9064) );
  NAND2_X1 U10447 ( .A1(n9064), .A2(n9044), .ZN(n9046) );
  AOI211_X1 U10448 ( .C1(n9057), .C2(n9046), .A(n9081), .B(n9045), .ZN(n9050)
         );
  OAI22_X1 U10449 ( .A1(n9048), .A2(n9102), .B1(n9047), .B2(n9100), .ZN(n9049)
         );
  NOR2_X1 U10450 ( .A1(n9050), .A2(n9049), .ZN(n9199) );
  INV_X1 U10451 ( .A(n9051), .ZN(n9053) );
  INV_X1 U10452 ( .A(n9030), .ZN(n9052) );
  AOI211_X1 U10453 ( .C1(n8539), .C2(n9053), .A(n10246), .B(n9052), .ZN(n9197)
         );
  INV_X1 U10454 ( .A(n9054), .ZN(n9055) );
  AOI22_X1 U10455 ( .A1(n4407), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9055), .B2(
        n9143), .ZN(n9056) );
  OAI21_X1 U10456 ( .B1(n8423), .B2(n9088), .A(n9056), .ZN(n9060) );
  XNOR2_X1 U10457 ( .A(n9058), .B(n4894), .ZN(n9200) );
  NOR2_X1 U10458 ( .A1(n9200), .A2(n9114), .ZN(n9059) );
  AOI211_X1 U10459 ( .C1(n9197), .C2(n9148), .A(n9060), .B(n9059), .ZN(n9061)
         );
  OAI21_X1 U10460 ( .B1(n9199), .B2(n4407), .A(n9061), .ZN(P2_U3274) );
  OAI21_X1 U10461 ( .B1(n9080), .B2(n9062), .A(n9073), .ZN(n9063) );
  NAND2_X1 U10462 ( .A1(n9064), .A2(n9063), .ZN(n9067) );
  AOI222_X1 U10463 ( .A1(n9138), .A2(n9067), .B1(n9066), .B2(n9120), .C1(n9065), .C2(n9121), .ZN(n9204) );
  INV_X1 U10464 ( .A(n9085), .ZN(n9068) );
  AOI21_X1 U10465 ( .B1(n9201), .B2(n9068), .A(n9051), .ZN(n9202) );
  AOI22_X1 U10466 ( .A1(n4407), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9069), .B2(
        n9143), .ZN(n9070) );
  OAI21_X1 U10467 ( .B1(n9071), .B2(n9088), .A(n9070), .ZN(n9075) );
  XNOR2_X1 U10468 ( .A(n9072), .B(n9073), .ZN(n9205) );
  NOR2_X1 U10469 ( .A1(n9205), .A2(n9114), .ZN(n9074) );
  AOI211_X1 U10470 ( .C1(n9202), .C2(n9076), .A(n9075), .B(n9074), .ZN(n9077)
         );
  OAI21_X1 U10471 ( .B1(n9204), .B2(n4407), .A(n9077), .ZN(P2_U3275) );
  INV_X1 U10472 ( .A(n9078), .ZN(n9090) );
  INV_X1 U10473 ( .A(n9079), .ZN(n9082) );
  AOI211_X1 U10474 ( .C1(n9090), .C2(n9082), .A(n9081), .B(n9080), .ZN(n9084)
         );
  NOR2_X1 U10475 ( .A1(n9084), .A2(n9083), .ZN(n9209) );
  AOI211_X1 U10476 ( .C1(n9207), .C2(n4434), .A(n10246), .B(n9085), .ZN(n9206)
         );
  AOI22_X1 U10477 ( .A1(n4407), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9086), .B2(
        n9143), .ZN(n9087) );
  OAI21_X1 U10478 ( .B1(n4849), .B2(n9088), .A(n9087), .ZN(n9092) );
  OAI21_X1 U10479 ( .B1(n4449), .B2(n9090), .A(n9089), .ZN(n9210) );
  NOR2_X1 U10480 ( .A1(n9210), .A2(n9114), .ZN(n9091) );
  AOI211_X1 U10481 ( .C1(n9206), .C2(n9148), .A(n9092), .B(n9091), .ZN(n9093)
         );
  OAI21_X1 U10482 ( .B1(n9209), .B2(n4407), .A(n9093), .ZN(P2_U3276) );
  INV_X1 U10483 ( .A(n9096), .ZN(n9095) );
  XNOR2_X1 U10484 ( .A(n9094), .B(n9095), .ZN(n9214) );
  NOR2_X1 U10485 ( .A1(n9097), .A2(n9096), .ZN(n9098) );
  OAI21_X1 U10486 ( .B1(n9099), .B2(n9098), .A(n9138), .ZN(n9106) );
  OAI22_X1 U10487 ( .A1(n9103), .A2(n9102), .B1(n9101), .B2(n9100), .ZN(n9104)
         );
  INV_X1 U10488 ( .A(n9104), .ZN(n9105) );
  NAND2_X1 U10489 ( .A1(n9106), .A2(n9105), .ZN(n9216) );
  NAND2_X1 U10490 ( .A1(n9216), .A2(n9144), .ZN(n9113) );
  OAI22_X1 U10491 ( .A1(n9144), .A2(n10482), .B1(n9107), .B2(n9124), .ZN(n9111) );
  AOI21_X1 U10492 ( .B1(n8393), .B2(n9211), .A(n10246), .ZN(n9108) );
  NAND2_X1 U10493 ( .A1(n9108), .A2(n4434), .ZN(n9213) );
  NOR2_X1 U10494 ( .A1(n9213), .A2(n9109), .ZN(n9110) );
  AOI211_X1 U10495 ( .C1(n9134), .C2(n9211), .A(n9111), .B(n9110), .ZN(n9112)
         );
  OAI211_X1 U10496 ( .C1(n9114), .C2(n9214), .A(n9113), .B(n9112), .ZN(
        P2_U3277) );
  OAI21_X1 U10497 ( .B1(n9116), .B2(n9115), .A(n7349), .ZN(n10224) );
  AOI22_X1 U10498 ( .A1(n9135), .A2(n10224), .B1(n9134), .B2(n7263), .ZN(n9130) );
  OAI21_X1 U10499 ( .B1(n9119), .B2(n9118), .A(n9117), .ZN(n9123) );
  AOI222_X1 U10500 ( .A1(n9138), .A2(n9123), .B1(n9122), .B2(n9121), .C1(n7343), .C2(n9120), .ZN(n10221) );
  OAI22_X1 U10501 ( .A1(n4407), .A2(n10221), .B1(n5167), .B2(n9124), .ZN(n9125) );
  INV_X1 U10502 ( .A(n9125), .ZN(n9129) );
  OR2_X1 U10503 ( .A1(n10222), .A2(n9146), .ZN(n9126) );
  AND3_X1 U10504 ( .A1(n9127), .A2(n9239), .A3(n9126), .ZN(n10219) );
  AOI22_X1 U10505 ( .A1(n4407), .A2(P2_REG2_REG_2__SCAN_IN), .B1(n9148), .B2(
        n10219), .ZN(n9128) );
  NAND3_X1 U10506 ( .A1(n9130), .A2(n9129), .A3(n9128), .ZN(P2_U3294) );
  OAI21_X1 U10507 ( .B1(n9136), .B2(n9132), .A(n9131), .ZN(n10217) );
  AOI22_X1 U10508 ( .A1(n9135), .A2(n10217), .B1(n9134), .B2(n9133), .ZN(n9151) );
  XNOR2_X1 U10509 ( .A(n9137), .B(n9136), .ZN(n9139) );
  NAND2_X1 U10510 ( .A1(n9139), .A2(n9138), .ZN(n9142) );
  INV_X1 U10511 ( .A(n9140), .ZN(n9141) );
  NAND2_X1 U10512 ( .A1(n9142), .A2(n9141), .ZN(n10215) );
  AOI22_X1 U10513 ( .A1(n9144), .A2(n10215), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9143), .ZN(n9150) );
  OAI21_X1 U10514 ( .B1(n10214), .B2(n9145), .A(n9239), .ZN(n9147) );
  NOR2_X1 U10515 ( .A1(n9147), .A2(n9146), .ZN(n10212) );
  AOI22_X1 U10516 ( .A1(n4407), .A2(P2_REG2_REG_1__SCAN_IN), .B1(n9148), .B2(
        n10212), .ZN(n9149) );
  NAND3_X1 U10517 ( .A1(n9151), .A2(n9150), .A3(n9149), .ZN(P2_U3295) );
  AOI21_X1 U10518 ( .B1(n9153), .B2(n9246), .A(n9152), .ZN(n9154) );
  OAI21_X1 U10519 ( .B1(n9155), .B2(n10246), .A(n9154), .ZN(n9251) );
  MUX2_X1 U10520 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9251), .S(n10263), .Z(
        P2_U3551) );
  NAND3_X1 U10521 ( .A1(n9157), .A2(n9239), .A3(n9156), .ZN(n9159) );
  OAI211_X1 U10522 ( .C1(n9160), .C2(n10245), .A(n9159), .B(n9158), .ZN(n9252)
         );
  MUX2_X1 U10523 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9252), .S(n10263), .Z(
        P2_U3550) );
  OAI211_X1 U10524 ( .C1(n9165), .C2(n9250), .A(n9164), .B(n9163), .ZN(n9253)
         );
  MUX2_X1 U10525 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9253), .S(n10263), .Z(
        P2_U3549) );
  AOI21_X1 U10526 ( .B1(n9246), .B2(n9168), .A(n9167), .ZN(n9169) );
  MUX2_X1 U10527 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9254), .S(n10263), .Z(
        P2_U3548) );
  AOI21_X1 U10528 ( .B1(n9246), .B2(n9172), .A(n9171), .ZN(n9173) );
  OAI211_X1 U10529 ( .C1(n9250), .C2(n9175), .A(n9174), .B(n9173), .ZN(n9255)
         );
  MUX2_X1 U10530 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9255), .S(n10263), .Z(
        P2_U3547) );
  AOI21_X1 U10531 ( .B1(n9246), .B2(n9177), .A(n9176), .ZN(n9178) );
  OAI211_X1 U10532 ( .C1(n9250), .C2(n9180), .A(n9179), .B(n9178), .ZN(n9256)
         );
  MUX2_X1 U10533 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9256), .S(n10263), .Z(
        P2_U3546) );
  AOI21_X1 U10534 ( .B1(n9246), .B2(n9182), .A(n9181), .ZN(n9183) );
  OAI211_X1 U10535 ( .C1(n9250), .C2(n9185), .A(n9184), .B(n9183), .ZN(n9257)
         );
  MUX2_X1 U10536 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9257), .S(n10263), .Z(
        P2_U3545) );
  OAI22_X1 U10537 ( .A1(n9187), .A2(n10246), .B1(n9186), .B2(n10245), .ZN(
        n9188) );
  INV_X1 U10538 ( .A(n9188), .ZN(n9189) );
  OAI211_X1 U10539 ( .C1(n9250), .C2(n9191), .A(n9190), .B(n9189), .ZN(n9258)
         );
  MUX2_X1 U10540 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9258), .S(n10263), .Z(
        P2_U3544) );
  AOI22_X1 U10541 ( .A1(n9193), .A2(n9239), .B1(n9246), .B2(n9192), .ZN(n9194)
         );
  OAI211_X1 U10542 ( .C1(n9250), .C2(n9196), .A(n4409), .B(n9194), .ZN(n9259)
         );
  MUX2_X1 U10543 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9259), .S(n10263), .Z(
        P2_U3543) );
  AOI21_X1 U10544 ( .B1(n9246), .B2(n8539), .A(n9197), .ZN(n9198) );
  OAI211_X1 U10545 ( .C1(n9250), .C2(n9200), .A(n9199), .B(n9198), .ZN(n9260)
         );
  MUX2_X1 U10546 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9260), .S(n10263), .Z(
        P2_U3542) );
  AOI22_X1 U10547 ( .A1(n9202), .A2(n9239), .B1(n9246), .B2(n9201), .ZN(n9203)
         );
  OAI211_X1 U10548 ( .C1(n9250), .C2(n9205), .A(n9204), .B(n9203), .ZN(n9261)
         );
  MUX2_X1 U10549 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9261), .S(n10263), .Z(
        P2_U3541) );
  AOI21_X1 U10550 ( .B1(n9246), .B2(n9207), .A(n9206), .ZN(n9208) );
  OAI211_X1 U10551 ( .C1(n9250), .C2(n9210), .A(n9209), .B(n9208), .ZN(n9262)
         );
  MUX2_X1 U10552 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9262), .S(n10263), .Z(
        P2_U3540) );
  NAND2_X1 U10553 ( .A1(n9211), .A2(n9246), .ZN(n9212) );
  OAI211_X1 U10554 ( .C1(n9214), .C2(n9250), .A(n9213), .B(n9212), .ZN(n9215)
         );
  MUX2_X1 U10555 ( .A(n9263), .B(P2_REG1_REG_19__SCAN_IN), .S(n10261), .Z(
        P2_U3539) );
  AOI21_X1 U10556 ( .B1(n9246), .B2(n9218), .A(n9217), .ZN(n9219) );
  OAI211_X1 U10557 ( .C1(n9250), .C2(n9221), .A(n9220), .B(n9219), .ZN(n9264)
         );
  MUX2_X1 U10558 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9264), .S(n10263), .Z(
        P2_U3538) );
  AOI22_X1 U10559 ( .A1(n9222), .A2(n9239), .B1(n9246), .B2(n8127), .ZN(n9223)
         );
  OAI211_X1 U10560 ( .C1(n9250), .C2(n9225), .A(n9224), .B(n9223), .ZN(n9265)
         );
  MUX2_X1 U10561 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9265), .S(n10263), .Z(
        P2_U3535) );
  AOI22_X1 U10562 ( .A1(n9227), .A2(n9239), .B1(n9246), .B2(n9226), .ZN(n9228)
         );
  OAI211_X1 U10563 ( .C1(n9230), .C2(n9250), .A(n9229), .B(n9228), .ZN(n9266)
         );
  MUX2_X1 U10564 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n9266), .S(n10263), .Z(
        P2_U3534) );
  INV_X1 U10565 ( .A(n9231), .ZN(n9236) );
  AOI22_X1 U10566 ( .A1(n9233), .A2(n9239), .B1(n9246), .B2(n9232), .ZN(n9234)
         );
  OAI211_X1 U10567 ( .C1(n9237), .C2(n9236), .A(n9235), .B(n9234), .ZN(n9267)
         );
  MUX2_X1 U10568 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n9267), .S(n10263), .Z(
        P2_U3533) );
  AOI22_X1 U10569 ( .A1(n9240), .A2(n9239), .B1(n9246), .B2(n9238), .ZN(n9241)
         );
  OAI211_X1 U10570 ( .C1(n9250), .C2(n9243), .A(n9242), .B(n9241), .ZN(n9268)
         );
  MUX2_X1 U10571 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9268), .S(n10263), .Z(
        P2_U3532) );
  AOI21_X1 U10572 ( .B1(n9246), .B2(n9245), .A(n9244), .ZN(n9247) );
  OAI211_X1 U10573 ( .C1(n9250), .C2(n9249), .A(n9248), .B(n9247), .ZN(n9269)
         );
  MUX2_X1 U10574 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9269), .S(n10263), .Z(
        P2_U3531) );
  MUX2_X1 U10575 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9251), .S(n10254), .Z(
        P2_U3519) );
  MUX2_X1 U10576 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9252), .S(n10254), .Z(
        P2_U3518) );
  MUX2_X1 U10577 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9253), .S(n10254), .Z(
        P2_U3517) );
  MUX2_X1 U10578 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9254), .S(n10254), .Z(
        P2_U3516) );
  MUX2_X1 U10579 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9255), .S(n10254), .Z(
        P2_U3515) );
  MUX2_X1 U10580 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9256), .S(n10254), .Z(
        P2_U3514) );
  MUX2_X1 U10581 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9257), .S(n10254), .Z(
        P2_U3513) );
  MUX2_X1 U10582 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9258), .S(n10254), .Z(
        P2_U3512) );
  MUX2_X1 U10583 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9259), .S(n10254), .Z(
        P2_U3511) );
  MUX2_X1 U10584 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9260), .S(n10254), .Z(
        P2_U3510) );
  MUX2_X1 U10585 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9261), .S(n10254), .Z(
        P2_U3509) );
  MUX2_X1 U10586 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9262), .S(n10254), .Z(
        P2_U3508) );
  MUX2_X1 U10587 ( .A(n9263), .B(P2_REG0_REG_19__SCAN_IN), .S(n10253), .Z(
        P2_U3507) );
  MUX2_X1 U10588 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9264), .S(n10254), .Z(
        P2_U3505) );
  MUX2_X1 U10589 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9265), .S(n10254), .Z(
        P2_U3496) );
  MUX2_X1 U10590 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n9266), .S(n10254), .Z(
        P2_U3493) );
  MUX2_X1 U10591 ( .A(P2_REG0_REG_13__SCAN_IN), .B(n9267), .S(n10254), .Z(
        P2_U3490) );
  MUX2_X1 U10592 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n9268), .S(n10254), .Z(
        P2_U3487) );
  MUX2_X1 U10593 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n9269), .S(n10254), .Z(
        P2_U3484) );
  INV_X1 U10594 ( .A(n9270), .ZN(n9916) );
  NOR4_X1 U10595 ( .A1(n9272), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9271), .A4(
        P2_U3152), .ZN(n9273) );
  AOI21_X1 U10596 ( .B1(n9279), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9273), .ZN(
        n9274) );
  OAI21_X1 U10597 ( .B1(n9916), .B2(n9281), .A(n9274), .ZN(P2_U3327) );
  INV_X1 U10598 ( .A(n9275), .ZN(n9920) );
  AOI22_X1 U10599 ( .A1(n9276), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n9279), .ZN(n9277) );
  OAI21_X1 U10600 ( .B1(n9920), .B2(n9281), .A(n9277), .ZN(P2_U3328) );
  AOI22_X1 U10601 ( .A1(n9278), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_29__SCAN_IN), .B2(n9279), .ZN(n9280) );
  OAI21_X1 U10602 ( .B1(n9282), .B2(n9281), .A(n9280), .ZN(P2_U3329) );
  INV_X1 U10603 ( .A(n9283), .ZN(n9285) );
  AND2_X1 U10604 ( .A1(n9287), .A2(n9286), .ZN(n9289) );
  NAND2_X1 U10605 ( .A1(n9289), .A2(n9288), .ZN(n9290) );
  XOR2_X1 U10606 ( .A(n9291), .B(n9290), .Z(n9298) );
  NAND2_X1 U10607 ( .A1(n9427), .A2(n9439), .ZN(n9293) );
  OAI211_X1 U10608 ( .C1(n9861), .C2(n9425), .A(n9293), .B(n9292), .ZN(n9294)
         );
  AOI21_X1 U10609 ( .B1(n9410), .B2(n9295), .A(n9294), .ZN(n9297) );
  NAND2_X1 U10610 ( .A1(n9864), .A2(n6949), .ZN(n9296) );
  OAI211_X1 U10611 ( .C1(n9298), .C2(n9432), .A(n9297), .B(n9296), .ZN(
        P1_U3213) );
  INV_X1 U10612 ( .A(n9299), .ZN(n9301) );
  NAND2_X1 U10613 ( .A1(n9301), .A2(n9300), .ZN(n9303) );
  XNOR2_X1 U10614 ( .A(n9303), .B(n9302), .ZN(n9308) );
  NAND2_X1 U10615 ( .A1(n9782), .A2(n9386), .ZN(n9305) );
  AOI22_X1 U10616 ( .A1(n9581), .A2(n9427), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9304) );
  OAI211_X1 U10617 ( .C1(n9429), .C2(n9583), .A(n9305), .B(n9304), .ZN(n9306)
         );
  AOI21_X1 U10618 ( .B1(n6260), .B2(n6949), .A(n9306), .ZN(n9307) );
  OAI21_X1 U10619 ( .B1(n9308), .B2(n9432), .A(n9307), .ZN(P1_U3214) );
  INV_X1 U10620 ( .A(n9309), .ZN(n9310) );
  AOI21_X1 U10621 ( .B1(n9312), .B2(n9311), .A(n9310), .ZN(n9317) );
  NAND2_X1 U10622 ( .A1(n9614), .A2(n9386), .ZN(n9313) );
  NAND2_X1 U10623 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9501) );
  OAI211_X1 U10624 ( .C1(n9844), .C2(n9384), .A(n9313), .B(n9501), .ZN(n9314)
         );
  AOI21_X1 U10625 ( .B1(n9640), .B2(n9410), .A(n9314), .ZN(n9316) );
  NOR2_X1 U10626 ( .A1(n9643), .A2(n10130), .ZN(n9827) );
  NAND2_X1 U10627 ( .A1(n9827), .A2(n9365), .ZN(n9315) );
  OAI211_X1 U10628 ( .C1(n9317), .C2(n9432), .A(n9316), .B(n9315), .ZN(
        P1_U3217) );
  NOR2_X1 U10629 ( .A1(n6879), .A2(n9319), .ZN(n9320) );
  XNOR2_X1 U10630 ( .A(n9321), .B(n9320), .ZN(n9328) );
  NAND2_X1 U10631 ( .A1(n9614), .A2(n9427), .ZN(n9322) );
  OAI21_X1 U10632 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n9323), .A(n9322), .ZN(
        n9324) );
  AOI21_X1 U10633 ( .B1(n9581), .B2(n9386), .A(n9324), .ZN(n9325) );
  OAI21_X1 U10634 ( .B1(n9612), .B2(n9429), .A(n9325), .ZN(n9326) );
  AOI21_X1 U10635 ( .B1(n9817), .B2(n6949), .A(n9326), .ZN(n9327) );
  OAI21_X1 U10636 ( .B1(n9328), .B2(n9432), .A(n9327), .ZN(P1_U3221) );
  NAND2_X1 U10637 ( .A1(n9689), .A2(n10163), .ZN(n9854) );
  NOR2_X1 U10638 ( .A1(n9329), .A2(n9330), .ZN(n9419) );
  NAND2_X1 U10639 ( .A1(n9329), .A2(n9330), .ZN(n9420) );
  OAI21_X1 U10640 ( .B1(n9419), .B2(n9422), .A(n9420), .ZN(n9334) );
  XNOR2_X1 U10641 ( .A(n9332), .B(n9331), .ZN(n9333) );
  XNOR2_X1 U10642 ( .A(n9334), .B(n9333), .ZN(n9335) );
  NAND2_X1 U10643 ( .A1(n9335), .A2(n9408), .ZN(n9339) );
  OAI22_X1 U10644 ( .A1(n9834), .A2(n9425), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n10445), .ZN(n9337) );
  NOR2_X1 U10645 ( .A1(n9429), .A2(n9686), .ZN(n9336) );
  AOI211_X1 U10646 ( .C1(n9427), .C2(n9696), .A(n9337), .B(n9336), .ZN(n9338)
         );
  OAI211_X1 U10647 ( .C1(n9402), .C2(n9854), .A(n9339), .B(n9338), .ZN(
        P1_U3224) );
  XNOR2_X1 U10648 ( .A(n9341), .B(n9340), .ZN(n9342) );
  XNOR2_X1 U10649 ( .A(n9343), .B(n9342), .ZN(n9348) );
  NAND2_X1 U10650 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9993) );
  NAND2_X1 U10651 ( .A1(n9427), .A2(n9676), .ZN(n9344) );
  OAI211_X1 U10652 ( .C1(n9844), .C2(n9425), .A(n9993), .B(n9344), .ZN(n9345)
         );
  AOI21_X1 U10653 ( .B1(n9410), .B2(n9675), .A(n9345), .ZN(n9347) );
  NAND2_X1 U10654 ( .A1(n9847), .A2(n6949), .ZN(n9346) );
  OAI211_X1 U10655 ( .C1(n9348), .C2(n9432), .A(n9347), .B(n9346), .ZN(
        P1_U3226) );
  AOI21_X1 U10656 ( .B1(n9351), .B2(n9350), .A(n9349), .ZN(n9356) );
  NAND2_X1 U10657 ( .A1(n9435), .A2(n9386), .ZN(n9353) );
  AOI22_X1 U10658 ( .A1(n9804), .A2(n9427), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9352) );
  OAI211_X1 U10659 ( .C1(n9429), .C2(n9570), .A(n9353), .B(n9352), .ZN(n9354)
         );
  AOI21_X1 U10660 ( .B1(n9795), .B2(n6949), .A(n9354), .ZN(n9355) );
  OAI21_X1 U10661 ( .B1(n9356), .B2(n9432), .A(n9355), .ZN(P1_U3227) );
  OAI21_X1 U10662 ( .B1(n9359), .B2(n9357), .A(n9358), .ZN(n9360) );
  NAND2_X1 U10663 ( .A1(n9360), .A2(n9408), .ZN(n9369) );
  AOI22_X1 U10664 ( .A1(n9362), .A2(n9361), .B1(P1_REG3_REG_4__SCAN_IN), .B2(
        P1_U3084), .ZN(n9368) );
  NAND2_X1 U10665 ( .A1(n9410), .A2(n9363), .ZN(n9367) );
  NOR2_X1 U10666 ( .A1(n10130), .A2(n9364), .ZN(n10102) );
  NAND2_X1 U10667 ( .A1(n9365), .A2(n10102), .ZN(n9366) );
  NAND4_X1 U10668 ( .A1(n9369), .A2(n9368), .A3(n9367), .A4(n9366), .ZN(
        P1_U3228) );
  INV_X1 U10669 ( .A(n9370), .ZN(n9372) );
  NAND2_X1 U10670 ( .A1(n9372), .A2(n9371), .ZN(n9373) );
  OAI22_X1 U10671 ( .A1(n9835), .A2(n9384), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n4656), .ZN(n9374) );
  AOI21_X1 U10672 ( .B1(n9803), .B2(n9386), .A(n9374), .ZN(n9375) );
  OAI21_X1 U10673 ( .B1(n9628), .B2(n9429), .A(n9375), .ZN(n9376) );
  AOI21_X1 U10674 ( .B1(n9823), .B2(n6949), .A(n9376), .ZN(n9377) );
  OAI21_X1 U10675 ( .B1(n9378), .B2(n9432), .A(n9377), .ZN(P1_U3231) );
  XNOR2_X1 U10676 ( .A(n9380), .B(n9379), .ZN(n9381) );
  XNOR2_X1 U10677 ( .A(n9382), .B(n9381), .ZN(n9391) );
  OAI22_X1 U10678 ( .A1(n9622), .A2(n9384), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9383), .ZN(n9385) );
  AOI21_X1 U10679 ( .B1(n9804), .B2(n9386), .A(n9385), .ZN(n9389) );
  INV_X1 U10680 ( .A(n9387), .ZN(n9596) );
  NAND2_X1 U10681 ( .A1(n9596), .A2(n9410), .ZN(n9388) );
  OAI211_X1 U10682 ( .C1(n9807), .C2(n9417), .A(n9389), .B(n9388), .ZN(n9390)
         );
  AOI21_X1 U10683 ( .B1(n9391), .B2(n9408), .A(n9390), .ZN(n9392) );
  INV_X1 U10684 ( .A(n9392), .ZN(P1_U3233) );
  NAND2_X1 U10685 ( .A1(n9662), .A2(n10163), .ZN(n9832) );
  XNOR2_X1 U10686 ( .A(n9394), .B(n9393), .ZN(n9395) );
  XNOR2_X1 U10687 ( .A(n9396), .B(n9395), .ZN(n9397) );
  NAND2_X1 U10688 ( .A1(n9397), .A2(n9408), .ZN(n9401) );
  NAND2_X1 U10689 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10014)
         );
  OAI21_X1 U10690 ( .B1(n9835), .B2(n9425), .A(n10014), .ZN(n9399) );
  NOR2_X1 U10691 ( .A1(n9429), .A2(n9651), .ZN(n9398) );
  AOI211_X1 U10692 ( .C1(n9427), .C2(n9695), .A(n9399), .B(n9398), .ZN(n9400)
         );
  OAI211_X1 U10693 ( .C1(n9402), .C2(n9832), .A(n9401), .B(n9400), .ZN(
        P1_U3236) );
  INV_X1 U10694 ( .A(n9403), .ZN(n9409) );
  OAI21_X1 U10695 ( .B1(n9406), .B2(n9405), .A(n9404), .ZN(n9407) );
  NAND3_X1 U10696 ( .A1(n9409), .A2(n9408), .A3(n9407), .ZN(n9416) );
  AOI22_X1 U10697 ( .A1(n9411), .A2(n9410), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9412) );
  OAI21_X1 U10698 ( .B1(n9413), .B2(n9425), .A(n9412), .ZN(n9414) );
  AOI21_X1 U10699 ( .B1(n9427), .B2(n9435), .A(n9414), .ZN(n9415) );
  OAI211_X1 U10700 ( .C1(n9418), .C2(n9417), .A(n9416), .B(n9415), .ZN(
        P1_U3238) );
  INV_X1 U10701 ( .A(n9419), .ZN(n9421) );
  NAND2_X1 U10702 ( .A1(n9421), .A2(n9420), .ZN(n9423) );
  XNOR2_X1 U10703 ( .A(n9423), .B(n9422), .ZN(n9433) );
  OAI21_X1 U10704 ( .B1(n9425), .B2(n9843), .A(n9424), .ZN(n9426) );
  AOI21_X1 U10705 ( .B1(n9427), .B2(n9438), .A(n9426), .ZN(n9428) );
  OAI21_X1 U10706 ( .B1(n9710), .B2(n9429), .A(n9428), .ZN(n9430) );
  AOI21_X1 U10707 ( .B1(n9856), .B2(n6949), .A(n9430), .ZN(n9431) );
  OAI21_X1 U10708 ( .B1(n9433), .B2(n9432), .A(n9431), .ZN(P1_U3239) );
  MUX2_X1 U10709 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9434), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10710 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9760), .S(P1_U4006), .Z(
        P1_U3584) );
  MUX2_X1 U10711 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9514), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10712 ( .A(n6276), .B(P1_DATAO_REG_27__SCAN_IN), .S(n9445), .Z(
        P1_U3582) );
  MUX2_X1 U10713 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9783), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10714 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9435), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10715 ( .A(n9782), .B(P1_DATAO_REG_24__SCAN_IN), .S(n9445), .Z(
        P1_U3579) );
  MUX2_X1 U10716 ( .A(n9804), .B(P1_DATAO_REG_23__SCAN_IN), .S(n9445), .Z(
        P1_U3578) );
  MUX2_X1 U10717 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9581), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10718 ( .A(n9803), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9445), .Z(
        P1_U3576) );
  MUX2_X1 U10719 ( .A(n9614), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9445), .Z(
        P1_U3575) );
  MUX2_X1 U10720 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9436), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10721 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9437), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10722 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9695), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10723 ( .A(n9676), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9445), .Z(
        P1_U3571) );
  MUX2_X1 U10724 ( .A(n9696), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9445), .Z(
        P1_U3570) );
  MUX2_X1 U10725 ( .A(n9438), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9445), .Z(
        P1_U3569) );
  MUX2_X1 U10726 ( .A(n9439), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9445), .Z(
        P1_U3568) );
  MUX2_X1 U10727 ( .A(n9440), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9445), .Z(
        P1_U3567) );
  MUX2_X1 U10728 ( .A(n9960), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9445), .Z(
        P1_U3566) );
  MUX2_X1 U10729 ( .A(n9441), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9445), .Z(
        P1_U3565) );
  MUX2_X1 U10730 ( .A(n9959), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9445), .Z(
        P1_U3564) );
  MUX2_X1 U10731 ( .A(n10158), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9445), .Z(
        P1_U3563) );
  MUX2_X1 U10732 ( .A(n9442), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9445), .Z(
        P1_U3562) );
  MUX2_X1 U10733 ( .A(n10160), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9445), .Z(
        P1_U3561) );
  MUX2_X1 U10734 ( .A(n9443), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9445), .Z(
        P1_U3560) );
  MUX2_X1 U10735 ( .A(n9444), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9445), .Z(
        P1_U3559) );
  MUX2_X1 U10736 ( .A(n10082), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9445), .Z(
        P1_U3558) );
  MUX2_X1 U10737 ( .A(n6711), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9445), .Z(
        P1_U3557) );
  MUX2_X1 U10738 ( .A(n6729), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9445), .Z(
        P1_U3556) );
  INV_X1 U10739 ( .A(n9446), .ZN(n9454) );
  INV_X1 U10740 ( .A(n9447), .ZN(n9449) );
  NAND3_X1 U10741 ( .A1(n9450), .A2(n9449), .A3(n9448), .ZN(n9451) );
  AOI21_X1 U10742 ( .B1(n9452), .B2(n9451), .A(n9994), .ZN(n9453) );
  AOI21_X1 U10743 ( .B1(n10001), .B2(n9454), .A(n9453), .ZN(n9462) );
  NAND2_X1 U10744 ( .A1(n9455), .A2(P1_ADDR_REG_5__SCAN_IN), .ZN(n9460) );
  OAI211_X1 U10745 ( .C1(n9458), .C2(n9457), .A(n10003), .B(n9456), .ZN(n9459)
         );
  NAND4_X1 U10746 ( .A1(n9462), .A2(n9461), .A3(n9460), .A4(n9459), .ZN(
        P1_U3246) );
  OAI21_X1 U10747 ( .B1(n9465), .B2(n9464), .A(n9463), .ZN(n9466) );
  NAND2_X1 U10748 ( .A1(n9466), .A2(n10003), .ZN(n9477) );
  INV_X1 U10749 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n10342) );
  OAI21_X1 U10750 ( .B1(n10026), .B2(n10342), .A(n9467), .ZN(n9468) );
  AOI21_X1 U10751 ( .B1(n9469), .B2(n10001), .A(n9468), .ZN(n9476) );
  MUX2_X1 U10752 ( .A(n9724), .B(P1_REG2_REG_10__SCAN_IN), .S(n9469), .Z(n9470) );
  NAND3_X1 U10753 ( .A1(n9472), .A2(n9471), .A3(n9470), .ZN(n9473) );
  NAND3_X1 U10754 ( .A1(n10013), .A2(n9474), .A3(n9473), .ZN(n9475) );
  NAND3_X1 U10755 ( .A1(n9477), .A2(n9476), .A3(n9475), .ZN(P1_U3251) );
  XNOR2_X1 U10756 ( .A(n9495), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n10021) );
  INV_X1 U10757 ( .A(n10000), .ZN(n9483) );
  INV_X1 U10758 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9482) );
  XOR2_X1 U10759 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10000), .Z(n10004) );
  AOI22_X1 U10760 ( .A1(n9480), .A2(n9488), .B1(P1_REG1_REG_15__SCAN_IN), .B2(
        n9479), .ZN(n9988) );
  XNOR2_X1 U10761 ( .A(n9987), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n9989) );
  INV_X1 U10762 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n10346) );
  OAI22_X1 U10763 ( .A1(n9988), .A2(n9989), .B1(n10346), .B2(n9481), .ZN(
        n10005) );
  NAND2_X1 U10764 ( .A1(n10004), .A2(n10005), .ZN(n10002) );
  OAI21_X1 U10765 ( .B1(n9483), .B2(n9482), .A(n10002), .ZN(n10020) );
  NOR2_X1 U10766 ( .A1(n10021), .A2(n10020), .ZN(n10019) );
  AOI21_X1 U10767 ( .B1(n10016), .B2(n9484), .A(n10019), .ZN(n9486) );
  XNOR2_X1 U10768 ( .A(n9486), .B(n9485), .ZN(n9497) );
  NAND2_X1 U10769 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9987), .ZN(n9490) );
  OAI21_X1 U10770 ( .B1(n9987), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9490), .ZN(
        n9983) );
  NAND2_X1 U10771 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n10000), .ZN(n9491) );
  OAI21_X1 U10772 ( .B1(n10000), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9491), .ZN(
        n9996) );
  AOI21_X1 U10773 ( .B1(n10000), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9995), .ZN(
        n10010) );
  INV_X1 U10774 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9492) );
  OR2_X1 U10775 ( .A1(n9495), .A2(n9492), .ZN(n9494) );
  NAND2_X1 U10776 ( .A1(n9495), .A2(n9492), .ZN(n9493) );
  AND2_X1 U10777 ( .A1(n9494), .A2(n9493), .ZN(n10011) );
  NOR2_X1 U10778 ( .A1(n10010), .A2(n10011), .ZN(n10009) );
  NAND2_X1 U10779 ( .A1(n9499), .A2(n10013), .ZN(n9496) );
  OAI211_X1 U10780 ( .C1(n9497), .C2(n10023), .A(n9496), .B(n10017), .ZN(n9500) );
  INV_X1 U10781 ( .A(n9497), .ZN(n9498) );
  NOR2_X1 U10782 ( .A1(n9750), .A2(n9529), .ZN(n9502) );
  XNOR2_X1 U10783 ( .A(n9508), .B(n9502), .ZN(n9748) );
  OAI21_X1 U10784 ( .B1(n9504), .B2(n9503), .A(n10159), .ZN(n9522) );
  INV_X1 U10785 ( .A(n9505), .ZN(n9506) );
  NOR2_X1 U10786 ( .A1(n9522), .A2(n9506), .ZN(n9749) );
  INV_X1 U10787 ( .A(n9749), .ZN(n9507) );
  NOR2_X1 U10788 ( .A1(n9507), .A2(n5064), .ZN(n9511) );
  NOR2_X1 U10789 ( .A1(n9508), .A2(n9725), .ZN(n9509) );
  AOI211_X1 U10790 ( .C1(n5064), .C2(P1_REG2_REG_31__SCAN_IN), .A(n9511), .B(
        n9509), .ZN(n9510) );
  OAI21_X1 U10791 ( .B1(n9748), .B2(n9659), .A(n9510), .ZN(P1_U3261) );
  XNOR2_X1 U10792 ( .A(n9750), .B(n9529), .ZN(n9752) );
  AOI21_X1 U10793 ( .B1(n5064), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9511), .ZN(
        n9513) );
  NAND2_X1 U10794 ( .A1(n9750), .A2(n9713), .ZN(n9512) );
  OAI211_X1 U10795 ( .C1(n9752), .C2(n9659), .A(n9513), .B(n9512), .ZN(
        P1_U3262) );
  NAND2_X1 U10796 ( .A1(n9515), .A2(n9514), .ZN(n9756) );
  NAND2_X1 U10797 ( .A1(n9764), .A2(n9756), .ZN(n9516) );
  XNOR2_X1 U10798 ( .A(n9516), .B(n9754), .ZN(n9535) );
  XNOR2_X1 U10799 ( .A(n9519), .B(n9754), .ZN(n9525) );
  OAI21_X1 U10800 ( .B1(n9525), .B2(n10040), .A(n9524), .ZN(n9753) );
  NAND2_X1 U10801 ( .A1(n9753), .A2(n9711), .ZN(n9534) );
  INV_X1 U10802 ( .A(n9526), .ZN(n9527) );
  NAND2_X1 U10803 ( .A1(n9757), .A2(n9527), .ZN(n9528) );
  AND2_X1 U10804 ( .A1(n9529), .A2(n9528), .ZN(n9766) );
  AOI22_X1 U10805 ( .A1(n9530), .A2(n10067), .B1(P1_REG2_REG_29__SCAN_IN), 
        .B2(n5064), .ZN(n9531) );
  OAI21_X1 U10806 ( .B1(n9759), .B2(n9725), .A(n9531), .ZN(n9532) );
  AOI21_X1 U10807 ( .B1(n9766), .B2(n9718), .A(n9532), .ZN(n9533) );
  OAI211_X1 U10808 ( .C1(n9535), .C2(n9738), .A(n9534), .B(n9533), .ZN(
        P1_U3355) );
  NAND2_X1 U10809 ( .A1(n9536), .A2(n9537), .ZN(n9539) );
  NAND2_X1 U10810 ( .A1(n9539), .A2(n9538), .ZN(n9540) );
  XNOR2_X1 U10811 ( .A(n9540), .B(n9542), .ZN(n9790) );
  OAI21_X1 U10812 ( .B1(n9543), .B2(n9542), .A(n9541), .ZN(n9788) );
  AOI21_X1 U10813 ( .B1(n9545), .B2(n9566), .A(n9544), .ZN(n9781) );
  NAND2_X1 U10814 ( .A1(n9781), .A2(n9718), .ZN(n9553) );
  OAI22_X1 U10815 ( .A1(n9547), .A2(n9731), .B1(n9546), .B2(n9711), .ZN(n9550)
         );
  NOR2_X1 U10816 ( .A1(n9548), .A2(n9726), .ZN(n9549) );
  AOI211_X1 U10817 ( .C1(n10067), .C2(n9551), .A(n9550), .B(n9549), .ZN(n9552)
         );
  OAI211_X1 U10818 ( .C1(n9786), .C2(n9725), .A(n9553), .B(n9552), .ZN(n9554)
         );
  AOI21_X1 U10819 ( .B1(n9788), .B2(n9672), .A(n9554), .ZN(n9555) );
  OAI21_X1 U10820 ( .B1(n9790), .B2(n9738), .A(n9555), .ZN(P1_U3266) );
  NAND2_X1 U10821 ( .A1(n9536), .A2(n9556), .ZN(n9577) );
  NAND2_X1 U10822 ( .A1(n9577), .A2(n9557), .ZN(n9559) );
  NAND2_X1 U10823 ( .A1(n9559), .A2(n9558), .ZN(n9560) );
  XOR2_X1 U10824 ( .A(n9563), .B(n9560), .Z(n9798) );
  NAND2_X1 U10825 ( .A1(n9562), .A2(n9561), .ZN(n9564) );
  XNOR2_X1 U10826 ( .A(n9564), .B(n9563), .ZN(n9565) );
  NAND2_X1 U10827 ( .A1(n9565), .A2(n10168), .ZN(n9797) );
  AOI21_X1 U10828 ( .B1(n8356), .B2(n9795), .A(n10132), .ZN(n9567) );
  NAND2_X1 U10829 ( .A1(n9793), .A2(n9568), .ZN(n9569) );
  OAI211_X1 U10830 ( .C1(n9728), .C2(n9570), .A(n9797), .B(n9569), .ZN(n9571)
         );
  NAND2_X1 U10831 ( .A1(n9571), .A2(n9711), .ZN(n9576) );
  NOR2_X1 U10832 ( .A1(n9792), .A2(n9726), .ZN(n9574) );
  OAI22_X1 U10833 ( .A1(n9791), .A2(n9731), .B1(n9572), .B2(n9711), .ZN(n9573)
         );
  AOI211_X1 U10834 ( .C1(n9795), .C2(n9713), .A(n9574), .B(n9573), .ZN(n9575)
         );
  OAI211_X1 U10835 ( .C1(n9798), .C2(n9738), .A(n9576), .B(n9575), .ZN(
        P1_U3267) );
  XNOR2_X1 U10836 ( .A(n9577), .B(n9578), .ZN(n9802) );
  XOR2_X1 U10837 ( .A(n9579), .B(n9578), .Z(n9580) );
  AOI222_X1 U10838 ( .A1(n9581), .A2(n10161), .B1(n10168), .B2(n9580), .C1(
        n9782), .C2(n10159), .ZN(n9801) );
  OAI22_X1 U10839 ( .A1(n9583), .A2(n9728), .B1(n9582), .B2(n9711), .ZN(n9584)
         );
  AOI21_X1 U10840 ( .B1(n6260), .B2(n9713), .A(n9584), .ZN(n9588) );
  OR2_X1 U10841 ( .A1(n9594), .A2(n9585), .ZN(n9586) );
  AND2_X1 U10842 ( .A1(n8356), .A2(n9586), .ZN(n9799) );
  NAND2_X1 U10843 ( .A1(n9799), .A2(n9718), .ZN(n9587) );
  OAI211_X1 U10844 ( .C1(n9801), .C2(n5064), .A(n9588), .B(n9587), .ZN(n9589)
         );
  INV_X1 U10845 ( .A(n9589), .ZN(n9590) );
  OAI21_X1 U10846 ( .B1(n9738), .B2(n9802), .A(n9590), .ZN(P1_U3268) );
  XNOR2_X1 U10847 ( .A(n9591), .B(n9592), .ZN(n9811) );
  XNOR2_X1 U10848 ( .A(n9593), .B(n9592), .ZN(n9809) );
  INV_X1 U10849 ( .A(n9594), .ZN(n9595) );
  OAI211_X1 U10850 ( .C1(n9807), .C2(n9610), .A(n9595), .B(n10117), .ZN(n9806)
         );
  NOR2_X1 U10851 ( .A1(n9791), .A2(n9726), .ZN(n9599) );
  AOI22_X1 U10852 ( .A1(n9596), .A2(n10067), .B1(P1_REG2_REG_22__SCAN_IN), 
        .B2(n5064), .ZN(n9597) );
  OAI21_X1 U10853 ( .B1(n9622), .B2(n9731), .A(n9597), .ZN(n9598) );
  AOI211_X1 U10854 ( .C1(n9600), .C2(n9713), .A(n9599), .B(n9598), .ZN(n9601)
         );
  OAI21_X1 U10855 ( .B1(n9806), .B2(n9691), .A(n9601), .ZN(n9602) );
  AOI21_X1 U10856 ( .B1(n9809), .B2(n9672), .A(n9602), .ZN(n9603) );
  OAI21_X1 U10857 ( .B1(n9738), .B2(n9811), .A(n9603), .ZN(P1_U3269) );
  OAI21_X1 U10858 ( .B1(n4450), .B2(n9605), .A(n9604), .ZN(n9820) );
  XNOR2_X1 U10859 ( .A(n9607), .B(n9606), .ZN(n9812) );
  NAND2_X1 U10860 ( .A1(n9812), .A2(n9672), .ZN(n9619) );
  NAND2_X1 U10861 ( .A1(n9625), .A2(n9817), .ZN(n9608) );
  NAND2_X1 U10862 ( .A1(n9608), .A2(n10117), .ZN(n9609) );
  NOR2_X1 U10863 ( .A1(n9610), .A2(n9609), .ZN(n9815) );
  NAND2_X1 U10864 ( .A1(n9817), .A2(n9713), .ZN(n9616) );
  OAI22_X1 U10865 ( .A1(n9612), .A2(n9728), .B1(n9611), .B2(n9711), .ZN(n9613)
         );
  AOI21_X1 U10866 ( .B1(n9677), .B2(n9614), .A(n9613), .ZN(n9615) );
  OAI211_X1 U10867 ( .C1(n9814), .C2(n9726), .A(n9616), .B(n9615), .ZN(n9617)
         );
  AOI21_X1 U10868 ( .B1(n9815), .B2(n9741), .A(n9617), .ZN(n9618) );
  OAI211_X1 U10869 ( .C1(n9820), .C2(n9738), .A(n9619), .B(n9618), .ZN(
        P1_U3270) );
  XOR2_X1 U10870 ( .A(n9620), .B(n9621), .Z(n9825) );
  XNOR2_X1 U10871 ( .A(n4481), .B(n9621), .ZN(n9623) );
  OAI222_X1 U10872 ( .A1(n9623), .A2(n10040), .B1(n10141), .B2(n9622), .C1(
        n10138), .C2(n9835), .ZN(n9821) );
  AOI21_X1 U10873 ( .B1(n9624), .B2(n9823), .A(n10132), .ZN(n9626) );
  AND2_X1 U10874 ( .A1(n9626), .A2(n9625), .ZN(n9822) );
  NAND2_X1 U10875 ( .A1(n9822), .A2(n9741), .ZN(n9631) );
  INV_X1 U10876 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n9627) );
  OAI22_X1 U10877 ( .A1(n9628), .A2(n9728), .B1(n9711), .B2(n9627), .ZN(n9629)
         );
  AOI21_X1 U10878 ( .B1(n9823), .B2(n9713), .A(n9629), .ZN(n9630) );
  NAND2_X1 U10879 ( .A1(n9631), .A2(n9630), .ZN(n9632) );
  AOI21_X1 U10880 ( .B1(n9821), .B2(n9711), .A(n9632), .ZN(n9633) );
  OAI21_X1 U10881 ( .B1(n9738), .B2(n9825), .A(n9633), .ZN(P1_U3271) );
  XNOR2_X1 U10882 ( .A(n9634), .B(n9636), .ZN(n9830) );
  AOI21_X1 U10883 ( .B1(n9637), .B2(n9636), .A(n9635), .ZN(n9638) );
  OAI222_X1 U10884 ( .A1(n10141), .A2(n9813), .B1(n10138), .B2(n9844), .C1(
        n9638), .C2(n10040), .ZN(n9828) );
  OR2_X1 U10885 ( .A1(n9658), .A2(n9643), .ZN(n9639) );
  AND3_X1 U10886 ( .A1(n9624), .A2(n9639), .A3(n10117), .ZN(n9826) );
  NAND2_X1 U10887 ( .A1(n9826), .A2(n9741), .ZN(n9642) );
  AOI22_X1 U10888 ( .A1(n5064), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9640), .B2(
        n10067), .ZN(n9641) );
  OAI211_X1 U10889 ( .C1(n9643), .C2(n9725), .A(n9642), .B(n9641), .ZN(n9644)
         );
  AOI21_X1 U10890 ( .B1(n9828), .B2(n9711), .A(n9644), .ZN(n9645) );
  OAI21_X1 U10891 ( .B1(n9738), .B2(n9830), .A(n9645), .ZN(P1_U3272) );
  INV_X1 U10892 ( .A(n9647), .ZN(n9649) );
  OAI21_X1 U10893 ( .B1(n9646), .B2(n9649), .A(n9648), .ZN(n9650) );
  XNOR2_X1 U10894 ( .A(n9650), .B(n9664), .ZN(n9841) );
  INV_X1 U10895 ( .A(n9672), .ZN(n9668) );
  INV_X1 U10896 ( .A(n9651), .ZN(n9652) );
  AOI22_X1 U10897 ( .A1(n5064), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9652), .B2(
        n10067), .ZN(n9654) );
  NAND2_X1 U10898 ( .A1(n9677), .A2(n9695), .ZN(n9653) );
  OAI211_X1 U10899 ( .C1(n9835), .C2(n9726), .A(n9654), .B(n9653), .ZN(n9661)
         );
  NOR2_X1 U10900 ( .A1(n9655), .A2(n9656), .ZN(n9657) );
  OR2_X1 U10901 ( .A1(n9658), .A2(n9657), .ZN(n9833) );
  NOR2_X1 U10902 ( .A1(n9833), .A2(n9659), .ZN(n9660) );
  AOI211_X1 U10903 ( .C1(n9713), .C2(n9662), .A(n9661), .B(n9660), .ZN(n9667)
         );
  NAND2_X1 U10904 ( .A1(n9665), .A2(n9664), .ZN(n9831) );
  NAND3_X1 U10905 ( .A1(n9663), .A2(n9831), .A3(n9700), .ZN(n9666) );
  OAI211_X1 U10906 ( .C1(n9841), .C2(n9668), .A(n9667), .B(n9666), .ZN(
        P1_U3273) );
  XNOR2_X1 U10907 ( .A(n9669), .B(n9670), .ZN(n9850) );
  XNOR2_X1 U10908 ( .A(n9646), .B(n9671), .ZN(n9842) );
  NAND2_X1 U10909 ( .A1(n9842), .A2(n9672), .ZN(n9683) );
  NAND2_X1 U10910 ( .A1(n5059), .A2(n9847), .ZN(n9673) );
  NAND2_X1 U10911 ( .A1(n9673), .A2(n10117), .ZN(n9674) );
  NOR2_X1 U10912 ( .A1(n9655), .A2(n9674), .ZN(n9845) );
  NOR2_X1 U10913 ( .A1(n4784), .A2(n9725), .ZN(n9681) );
  AOI22_X1 U10914 ( .A1(n5064), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9675), .B2(
        n10067), .ZN(n9679) );
  NAND2_X1 U10915 ( .A1(n9677), .A2(n9676), .ZN(n9678) );
  OAI211_X1 U10916 ( .C1(n9844), .C2(n9726), .A(n9679), .B(n9678), .ZN(n9680)
         );
  AOI211_X1 U10917 ( .C1(n9845), .C2(n9741), .A(n9681), .B(n9680), .ZN(n9682)
         );
  OAI211_X1 U10918 ( .C1(n9850), .C2(n9738), .A(n9683), .B(n9682), .ZN(
        P1_U3274) );
  XNOR2_X1 U10919 ( .A(n9684), .B(n9693), .ZN(n9851) );
  AOI21_X1 U10920 ( .B1(n9716), .B2(n9689), .A(n10132), .ZN(n9685) );
  NAND2_X1 U10921 ( .A1(n9685), .A2(n5059), .ZN(n9852) );
  INV_X1 U10922 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9687) );
  OAI22_X1 U10923 ( .A1(n9711), .A2(n9687), .B1(n9686), .B2(n9728), .ZN(n9688)
         );
  AOI21_X1 U10924 ( .B1(n9689), .B2(n9713), .A(n9688), .ZN(n9690) );
  OAI21_X1 U10925 ( .B1(n9852), .B2(n9691), .A(n9690), .ZN(n9699) );
  OAI21_X1 U10926 ( .B1(n9694), .B2(n9693), .A(n9692), .ZN(n9697) );
  AOI222_X1 U10927 ( .A1(n9697), .A2(n10168), .B1(n9696), .B2(n10161), .C1(
        n9695), .C2(n10159), .ZN(n9855) );
  NOR2_X1 U10928 ( .A1(n9855), .A2(n5064), .ZN(n9698) );
  AOI211_X1 U10929 ( .C1(n9851), .C2(n9700), .A(n9699), .B(n9698), .ZN(n9701)
         );
  INV_X1 U10930 ( .A(n9701), .ZN(P1_U3275) );
  XOR2_X1 U10931 ( .A(n9702), .B(n9704), .Z(n9707) );
  OAI22_X1 U10932 ( .A1(n9843), .A2(n10141), .B1(n9868), .B2(n10138), .ZN(
        n9706) );
  XNOR2_X1 U10933 ( .A(n9703), .B(n9704), .ZN(n9860) );
  NOR2_X1 U10934 ( .A1(n9860), .A2(n6712), .ZN(n9705) );
  AOI211_X1 U10935 ( .C1(n9707), .C2(n10168), .A(n9706), .B(n9705), .ZN(n9859)
         );
  INV_X1 U10936 ( .A(n9708), .ZN(n9709) );
  NAND2_X1 U10937 ( .A1(n9711), .A2(n9709), .ZN(n10068) );
  OAI22_X1 U10938 ( .A1(n9711), .A2(n7835), .B1(n9710), .B2(n9728), .ZN(n9712)
         );
  AOI21_X1 U10939 ( .B1(n9856), .B2(n9713), .A(n9712), .ZN(n9720) );
  OR2_X1 U10940 ( .A1(n9715), .A2(n9714), .ZN(n9717) );
  AND2_X1 U10941 ( .A1(n9717), .A2(n9716), .ZN(n9857) );
  NAND2_X1 U10942 ( .A1(n9857), .A2(n9718), .ZN(n9719) );
  OAI211_X1 U10943 ( .C1(n9860), .C2(n10068), .A(n9720), .B(n9719), .ZN(n9721)
         );
  INV_X1 U10944 ( .A(n9721), .ZN(n9722) );
  OAI21_X1 U10945 ( .B1(n9859), .B2(n5064), .A(n9722), .ZN(P1_U3276) );
  OAI211_X1 U10946 ( .C1(n8039), .C2(n9734), .A(n10168), .B(n9723), .ZN(n9964)
         );
  MUX2_X1 U10947 ( .A(n9964), .B(n9724), .S(n5064), .Z(n9745) );
  OAI22_X1 U10948 ( .A1(n9876), .A2(n9726), .B1(n9725), .B2(n9963), .ZN(n9733)
         );
  INV_X1 U10949 ( .A(n9727), .ZN(n9729) );
  OAI22_X1 U10950 ( .A1(n9731), .A2(n9730), .B1(n9729), .B2(n9728), .ZN(n9732)
         );
  NOR2_X1 U10951 ( .A1(n9733), .A2(n9732), .ZN(n9744) );
  NAND2_X1 U10952 ( .A1(n9735), .A2(n9734), .ZN(n9736) );
  NAND2_X1 U10953 ( .A1(n9737), .A2(n9736), .ZN(n9967) );
  NAND2_X1 U10954 ( .A1(n9967), .A2(n9700), .ZN(n9743) );
  OAI21_X1 U10955 ( .B1(n9739), .B2(n9963), .A(n10117), .ZN(n9740) );
  NOR2_X1 U10956 ( .A1(n9740), .A2(n8058), .ZN(n9958) );
  NAND2_X1 U10957 ( .A1(n9958), .A2(n9741), .ZN(n9742) );
  NAND4_X1 U10958 ( .A1(n9745), .A2(n9744), .A3(n9743), .A4(n9742), .ZN(
        P1_U3281) );
  AOI21_X1 U10959 ( .B1(n9746), .B2(n10163), .A(n9749), .ZN(n9747) );
  OAI21_X1 U10960 ( .B1(n9748), .B2(n10132), .A(n9747), .ZN(n9892) );
  MUX2_X1 U10961 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9892), .S(n10177), .Z(
        P1_U3554) );
  AOI21_X1 U10962 ( .B1(n9750), .B2(n10163), .A(n9749), .ZN(n9751) );
  OAI21_X1 U10963 ( .B1(n9752), .B2(n10132), .A(n9751), .ZN(n9893) );
  MUX2_X1 U10964 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9893), .S(n10177), .Z(
        P1_U3553) );
  INV_X1 U10965 ( .A(n9753), .ZN(n9769) );
  NAND4_X1 U10966 ( .A1(n9764), .A2(n9754), .A3(n10128), .A4(n9756), .ZN(n9768) );
  OR2_X1 U10967 ( .A1(n9756), .A2(n10172), .ZN(n9761) );
  OAI211_X1 U10968 ( .C1(n9761), .C2(n9758), .A(n10130), .B(n9757), .ZN(n9763)
         );
  OAI21_X1 U10969 ( .B1(n9761), .B2(n9760), .A(n9759), .ZN(n9762) );
  NAND2_X1 U10970 ( .A1(n9769), .A2(n5061), .ZN(n9894) );
  MUX2_X1 U10971 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9894), .S(n10177), .Z(
        P1_U3552) );
  OAI22_X1 U10972 ( .A1(n9771), .A2(n10132), .B1(n9770), .B2(n10130), .ZN(
        n9772) );
  INV_X1 U10973 ( .A(n9772), .ZN(n9773) );
  OAI211_X1 U10974 ( .C1(n10172), .C2(n9775), .A(n9774), .B(n9773), .ZN(n9895)
         );
  MUX2_X1 U10975 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9895), .S(n10177), .Z(
        P1_U3550) );
  AOI22_X1 U10976 ( .A1(n9777), .A2(n10117), .B1(n10163), .B2(n9776), .ZN(
        n9778) );
  OAI211_X1 U10977 ( .C1(n10172), .C2(n9780), .A(n9779), .B(n9778), .ZN(n9896)
         );
  MUX2_X1 U10978 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9896), .S(n10177), .Z(
        P1_U3549) );
  NAND2_X1 U10979 ( .A1(n9781), .A2(n10117), .ZN(n9785) );
  AOI22_X1 U10980 ( .A1(n9783), .A2(n10159), .B1(n10161), .B2(n9782), .ZN(
        n9784) );
  OAI211_X1 U10981 ( .C1(n9786), .C2(n10130), .A(n9785), .B(n9784), .ZN(n9787)
         );
  AOI21_X1 U10982 ( .B1(n9788), .B2(n10168), .A(n9787), .ZN(n9789) );
  OAI21_X1 U10983 ( .B1(n10172), .B2(n9790), .A(n9789), .ZN(n9897) );
  MUX2_X1 U10984 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9897), .S(n10177), .Z(
        P1_U3548) );
  OAI22_X1 U10985 ( .A1(n9792), .A2(n10141), .B1(n9791), .B2(n10138), .ZN(
        n9794) );
  AOI211_X1 U10986 ( .C1(n10163), .C2(n9795), .A(n9794), .B(n9793), .ZN(n9796)
         );
  OAI211_X1 U10987 ( .C1(n10172), .C2(n9798), .A(n9797), .B(n9796), .ZN(n9898)
         );
  MUX2_X1 U10988 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9898), .S(n10177), .Z(
        P1_U3547) );
  AOI22_X1 U10989 ( .A1(n9799), .A2(n10117), .B1(n10163), .B2(n6260), .ZN(
        n9800) );
  OAI211_X1 U10990 ( .C1(n10172), .C2(n9802), .A(n9801), .B(n9800), .ZN(n9899)
         );
  MUX2_X1 U10991 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9899), .S(n10177), .Z(
        P1_U3546) );
  AOI22_X1 U10992 ( .A1(n9804), .A2(n10159), .B1(n10161), .B2(n9803), .ZN(
        n9805) );
  OAI211_X1 U10993 ( .C1(n9807), .C2(n10130), .A(n9806), .B(n9805), .ZN(n9808)
         );
  AOI21_X1 U10994 ( .B1(n9809), .B2(n10168), .A(n9808), .ZN(n9810) );
  OAI21_X1 U10995 ( .B1(n10172), .B2(n9811), .A(n9810), .ZN(n9900) );
  MUX2_X1 U10996 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9900), .S(n10177), .Z(
        P1_U3545) );
  NAND2_X1 U10997 ( .A1(n9812), .A2(n10168), .ZN(n9819) );
  OAI22_X1 U10998 ( .A1(n9814), .A2(n10141), .B1(n9813), .B2(n10138), .ZN(
        n9816) );
  AOI211_X1 U10999 ( .C1(n10163), .C2(n9817), .A(n9816), .B(n9815), .ZN(n9818)
         );
  OAI211_X1 U11000 ( .C1(n10172), .C2(n9820), .A(n9819), .B(n9818), .ZN(n9901)
         );
  MUX2_X1 U11001 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9901), .S(n10177), .Z(
        P1_U3544) );
  AOI211_X1 U11002 ( .C1(n10163), .C2(n9823), .A(n9822), .B(n9821), .ZN(n9824)
         );
  OAI21_X1 U11003 ( .B1(n10172), .B2(n9825), .A(n9824), .ZN(n9902) );
  MUX2_X1 U11004 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9902), .S(n10177), .Z(
        P1_U3543) );
  NOR3_X1 U11005 ( .A1(n9828), .A2(n9827), .A3(n9826), .ZN(n9829) );
  OAI21_X1 U11006 ( .B1(n10172), .B2(n9830), .A(n9829), .ZN(n9903) );
  MUX2_X1 U11007 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9903), .S(n10177), .Z(
        P1_U3542) );
  AND3_X1 U11008 ( .A1(n9663), .A2(n9831), .A3(n10128), .ZN(n9839) );
  INV_X1 U11009 ( .A(n9832), .ZN(n9838) );
  NOR2_X1 U11010 ( .A1(n9833), .A2(n10132), .ZN(n9837) );
  OAI22_X1 U11011 ( .A1(n9835), .A2(n10141), .B1(n9834), .B2(n10138), .ZN(
        n9836) );
  NOR4_X1 U11012 ( .A1(n9839), .A2(n9838), .A3(n9837), .A4(n9836), .ZN(n9840)
         );
  OAI21_X1 U11013 ( .B1(n9841), .B2(n10040), .A(n9840), .ZN(n9904) );
  MUX2_X1 U11014 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9904), .S(n10177), .Z(
        P1_U3541) );
  NAND2_X1 U11015 ( .A1(n9842), .A2(n10168), .ZN(n9849) );
  OAI22_X1 U11016 ( .A1(n9844), .A2(n10141), .B1(n9843), .B2(n10138), .ZN(
        n9846) );
  AOI211_X1 U11017 ( .C1(n10163), .C2(n9847), .A(n9846), .B(n9845), .ZN(n9848)
         );
  OAI211_X1 U11018 ( .C1(n10172), .C2(n9850), .A(n9849), .B(n9848), .ZN(n9905)
         );
  MUX2_X1 U11019 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9905), .S(n10177), .Z(
        P1_U3540) );
  NAND2_X1 U11020 ( .A1(n9851), .A2(n10128), .ZN(n9853) );
  NAND4_X1 U11021 ( .A1(n9855), .A2(n9854), .A3(n9853), .A4(n9852), .ZN(n9906)
         );
  MUX2_X1 U11022 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9906), .S(n10177), .Z(
        P1_U3539) );
  AOI22_X1 U11023 ( .A1(n9857), .A2(n10117), .B1(n10163), .B2(n9856), .ZN(
        n9858) );
  OAI211_X1 U11024 ( .C1(n10089), .C2(n9860), .A(n9859), .B(n9858), .ZN(n9907)
         );
  MUX2_X1 U11025 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9907), .S(n10177), .Z(
        P1_U3538) );
  NOR2_X1 U11026 ( .A1(n10141), .A2(n9861), .ZN(n9863) );
  AOI211_X1 U11027 ( .C1(n10163), .C2(n9864), .A(n9863), .B(n9862), .ZN(n9865)
         );
  OAI211_X1 U11028 ( .C1(n10172), .C2(n9867), .A(n9866), .B(n9865), .ZN(n9908)
         );
  MUX2_X1 U11029 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9908), .S(n10177), .Z(
        P1_U3537) );
  OAI22_X1 U11030 ( .A1(n10141), .A2(n9868), .B1(n9884), .B2(n10138), .ZN(
        n9871) );
  NOR2_X1 U11031 ( .A1(n9869), .A2(n10132), .ZN(n9870) );
  AOI211_X1 U11032 ( .C1(n10163), .C2(n9872), .A(n9871), .B(n9870), .ZN(n9873)
         );
  OAI211_X1 U11033 ( .C1(n10172), .C2(n9875), .A(n9874), .B(n9873), .ZN(n9909)
         );
  MUX2_X1 U11034 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9909), .S(n10177), .Z(
        P1_U3536) );
  OAI22_X1 U11035 ( .A1(n10141), .A2(n9877), .B1(n9876), .B2(n10138), .ZN(
        n9879) );
  AOI211_X1 U11036 ( .C1(n10163), .C2(n9880), .A(n9879), .B(n9878), .ZN(n9882)
         );
  OAI211_X1 U11037 ( .C1(n10172), .C2(n9883), .A(n9882), .B(n9881), .ZN(n9910)
         );
  MUX2_X1 U11038 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9910), .S(n10177), .Z(
        P1_U3535) );
  OAI22_X1 U11039 ( .A1(n10141), .A2(n9884), .B1(n10140), .B2(n10138), .ZN(
        n9887) );
  NOR2_X1 U11040 ( .A1(n9885), .A2(n10132), .ZN(n9886) );
  AOI211_X1 U11041 ( .C1(n10163), .C2(n9888), .A(n9887), .B(n9886), .ZN(n9889)
         );
  OAI211_X1 U11042 ( .C1(n10172), .C2(n9891), .A(n9890), .B(n9889), .ZN(n9911)
         );
  MUX2_X1 U11043 ( .A(n9911), .B(P1_REG1_REG_11__SCAN_IN), .S(n10175), .Z(
        P1_U3534) );
  MUX2_X1 U11044 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9892), .S(n10588), .Z(
        P1_U3522) );
  MUX2_X1 U11045 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9893), .S(n10588), .Z(
        P1_U3521) );
  MUX2_X1 U11046 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9894), .S(n10588), .Z(
        P1_U3520) );
  MUX2_X1 U11047 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9895), .S(n10588), .Z(
        P1_U3518) );
  MUX2_X1 U11048 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9896), .S(n10588), .Z(
        P1_U3517) );
  MUX2_X1 U11049 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9897), .S(n10588), .Z(
        P1_U3516) );
  MUX2_X1 U11050 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9898), .S(n10588), .Z(
        P1_U3515) );
  MUX2_X1 U11051 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9899), .S(n10588), .Z(
        P1_U3514) );
  MUX2_X1 U11052 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9900), .S(n10588), .Z(
        P1_U3513) );
  MUX2_X1 U11053 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9901), .S(n10588), .Z(
        P1_U3512) );
  MUX2_X1 U11054 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9902), .S(n10588), .Z(
        P1_U3511) );
  MUX2_X1 U11055 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9903), .S(n10588), .Z(
        P1_U3510) );
  MUX2_X1 U11056 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9904), .S(n10588), .Z(
        P1_U3508) );
  MUX2_X1 U11057 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9905), .S(n10588), .Z(
        P1_U3505) );
  MUX2_X1 U11058 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9906), .S(n10588), .Z(
        P1_U3502) );
  MUX2_X1 U11059 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9907), .S(n10588), .Z(
        P1_U3499) );
  MUX2_X1 U11060 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9908), .S(n10588), .Z(
        P1_U3496) );
  MUX2_X1 U11061 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9909), .S(n10588), .Z(
        P1_U3493) );
  MUX2_X1 U11062 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n9910), .S(n10588), .Z(
        P1_U3490) );
  MUX2_X1 U11063 ( .A(n9911), .B(P1_REG0_REG_11__SCAN_IN), .S(n10586), .Z(
        P1_U3487) );
  NAND3_X1 U11064 ( .A1(n4549), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n9913) );
  OAI22_X1 U11065 ( .A1(n5868), .A2(n9913), .B1(n9912), .B2(n4405), .ZN(n9914)
         );
  INV_X1 U11066 ( .A(n9914), .ZN(n9915) );
  OAI21_X1 U11067 ( .B1(n9916), .B2(n9921), .A(n9915), .ZN(P1_U3322) );
  OAI222_X1 U11068 ( .A1(n9921), .A2(n9920), .B1(P1_U3084), .B2(n9917), .C1(
        n9918), .C2(n4405), .ZN(P1_U3323) );
  OAI222_X1 U11069 ( .A1(n4405), .A2(n9924), .B1(n9923), .B2(n9922), .C1(n4412), .C2(P1_U3084), .ZN(P1_U3325) );
  MUX2_X1 U11070 ( .A(n9926), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  INV_X1 U11071 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10598) );
  NOR2_X1 U11072 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9927) );
  AOI21_X1 U11073 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9927), .ZN(n10270) );
  NOR2_X1 U11074 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9928) );
  AOI21_X1 U11075 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9928), .ZN(n10273) );
  NOR2_X1 U11076 ( .A1(P1_ADDR_REG_15__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .ZN(n9929) );
  AOI21_X1 U11077 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9929), .ZN(n10276) );
  NOR2_X1 U11078 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9930) );
  AOI21_X1 U11079 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9930), .ZN(n10279) );
  NOR2_X1 U11080 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9931) );
  AOI21_X1 U11081 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9931), .ZN(n10282) );
  NOR2_X1 U11082 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9938) );
  XNOR2_X1 U11083 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10612) );
  NAND2_X1 U11084 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9936) );
  XOR2_X1 U11085 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10610) );
  NAND2_X1 U11086 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9934) );
  XOR2_X1 U11087 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10608) );
  AOI21_X1 U11088 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10264) );
  INV_X1 U11089 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9932) );
  NAND3_X1 U11090 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10266) );
  NAND2_X1 U11091 ( .A1(n10608), .A2(n10607), .ZN(n9933) );
  NAND2_X1 U11092 ( .A1(n9934), .A2(n9933), .ZN(n10609) );
  NAND2_X1 U11093 ( .A1(n10610), .A2(n10609), .ZN(n9935) );
  NAND2_X1 U11094 ( .A1(n9936), .A2(n9935), .ZN(n10611) );
  NOR2_X1 U11095 ( .A1(n10612), .A2(n10611), .ZN(n9937) );
  NOR2_X1 U11096 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9939), .ZN(n10594) );
  NAND2_X1 U11097 ( .A1(n9941), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9943) );
  NAND2_X1 U11098 ( .A1(n10592), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9942) );
  NAND2_X1 U11099 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9944), .ZN(n9946) );
  NAND2_X1 U11100 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10606), .ZN(n9945) );
  NAND2_X1 U11101 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9947), .ZN(n9949) );
  NAND2_X1 U11102 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10604), .ZN(n9948) );
  NAND2_X1 U11103 ( .A1(n9949), .A2(n9948), .ZN(n9950) );
  AND2_X1 U11104 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9950), .ZN(n9951) );
  XNOR2_X1 U11105 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9950), .ZN(n10601) );
  NAND2_X1 U11106 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n9952) );
  OAI21_X1 U11107 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9952), .ZN(n10290) );
  NAND2_X1 U11108 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9953) );
  OAI21_X1 U11109 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9953), .ZN(n10287) );
  NOR2_X1 U11110 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9954) );
  AOI21_X1 U11111 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9954), .ZN(n10284) );
  NAND2_X1 U11112 ( .A1(n10279), .A2(n10278), .ZN(n10277) );
  NAND2_X1 U11113 ( .A1(n10276), .A2(n10275), .ZN(n10274) );
  NAND2_X1 U11114 ( .A1(n10270), .A2(n10269), .ZN(n10268) );
  NOR2_X1 U11115 ( .A1(n10598), .A2(n10597), .ZN(n9955) );
  NAND2_X1 U11116 ( .A1(n10598), .A2(n10597), .ZN(n10596) );
  XNOR2_X1 U11117 ( .A(n9478), .B(P2_ADDR_REG_19__SCAN_IN), .ZN(n9956) );
  XNOR2_X1 U11118 ( .A(n9957), .B(n9956), .ZN(ADD_1071_U4) );
  INV_X1 U11119 ( .A(n9958), .ZN(n9962) );
  AOI22_X1 U11120 ( .A1(n10159), .A2(n9960), .B1(n10161), .B2(n9959), .ZN(
        n9961) );
  OAI211_X1 U11121 ( .C1(n9963), .C2(n10130), .A(n9962), .B(n9961), .ZN(n9966)
         );
  INV_X1 U11122 ( .A(n9964), .ZN(n9965) );
  AOI211_X1 U11123 ( .C1(n10128), .C2(n9967), .A(n9966), .B(n9965), .ZN(n9968)
         );
  INV_X1 U11124 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n10497) );
  AOI22_X1 U11125 ( .A1(n10588), .A2(n9968), .B1(n10497), .B2(n10586), .ZN(
        P1_U3484) );
  AOI22_X1 U11126 ( .A1(n10177), .A2(n9968), .B1(n7219), .B2(n10175), .ZN(
        P1_U3533) );
  XNOR2_X1 U11127 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11128 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  OAI211_X1 U11129 ( .C1(n9971), .C2(n9970), .A(n9969), .B(n10013), .ZN(n9973)
         );
  OAI211_X1 U11130 ( .C1(n10017), .C2(n9974), .A(n9973), .B(n9972), .ZN(n9975)
         );
  INV_X1 U11131 ( .A(n9975), .ZN(n9981) );
  NOR2_X1 U11132 ( .A1(n9977), .A2(n9976), .ZN(n9979) );
  OAI21_X1 U11133 ( .B1(n9979), .B2(n9978), .A(n10003), .ZN(n9980) );
  OAI211_X1 U11134 ( .C1(n4514), .C2(n10026), .A(n9981), .B(n9980), .ZN(
        P1_U3254) );
  NOR2_X1 U11135 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10445), .ZN(n9986) );
  AOI211_X1 U11136 ( .C1(n9984), .C2(n9983), .A(n9994), .B(n9982), .ZN(n9985)
         );
  AOI211_X1 U11137 ( .C1(n10001), .C2(n9987), .A(n9986), .B(n9985), .ZN(n9992)
         );
  XOR2_X1 U11138 ( .A(n9989), .B(n9988), .Z(n9990) );
  NAND2_X1 U11139 ( .A1(n9990), .A2(n10003), .ZN(n9991) );
  OAI211_X1 U11140 ( .C1(n4517), .C2(n10026), .A(n9992), .B(n9991), .ZN(
        P1_U3257) );
  INV_X1 U11141 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10008) );
  INV_X1 U11142 ( .A(n9993), .ZN(n9999) );
  AOI211_X1 U11143 ( .C1(n9997), .C2(n9996), .A(n9995), .B(n9994), .ZN(n9998)
         );
  AOI211_X1 U11144 ( .C1(n10001), .C2(n10000), .A(n9999), .B(n9998), .ZN(
        n10007) );
  OAI211_X1 U11145 ( .C1(n10005), .C2(n10004), .A(n10003), .B(n10002), .ZN(
        n10006) );
  OAI211_X1 U11146 ( .C1(n10008), .C2(n10026), .A(n10007), .B(n10006), .ZN(
        P1_U3258) );
  INV_X1 U11147 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10512) );
  AOI21_X1 U11148 ( .B1(n10011), .B2(n10010), .A(n10009), .ZN(n10012) );
  NAND2_X1 U11149 ( .A1(n10013), .A2(n10012), .ZN(n10015) );
  OAI211_X1 U11150 ( .C1(n10017), .C2(n10016), .A(n10015), .B(n10014), .ZN(
        n10018) );
  INV_X1 U11151 ( .A(n10018), .ZN(n10025) );
  AOI21_X1 U11152 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(n10022) );
  OR2_X1 U11153 ( .A1(n10023), .A2(n10022), .ZN(n10024) );
  OAI211_X1 U11154 ( .C1(n10512), .C2(n10026), .A(n10025), .B(n10024), .ZN(
        P1_U3259) );
  XOR2_X1 U11155 ( .A(n10035), .B(n10027), .Z(n10113) );
  NAND2_X1 U11156 ( .A1(n10028), .A2(n10031), .ZN(n10029) );
  NAND3_X1 U11157 ( .A1(n10030), .A2(n10117), .A3(n10029), .ZN(n10110) );
  AOI22_X1 U11158 ( .A1(n10067), .A2(n10032), .B1(n10050), .B2(n10031), .ZN(
        n10033) );
  OAI21_X1 U11159 ( .B1(n10110), .B2(n10052), .A(n10033), .ZN(n10044) );
  INV_X1 U11160 ( .A(n10034), .ZN(n10039) );
  INV_X1 U11161 ( .A(n10035), .ZN(n10038) );
  INV_X1 U11162 ( .A(n10036), .ZN(n10037) );
  AOI21_X1 U11163 ( .B1(n10039), .B2(n10038), .A(n10037), .ZN(n10041) );
  OAI222_X1 U11164 ( .A1(n10141), .A2(n10043), .B1(n10138), .B2(n10042), .C1(
        n10041), .C2(n10040), .ZN(n10111) );
  AOI211_X1 U11165 ( .C1(n10045), .C2(n10113), .A(n10044), .B(n10111), .ZN(
        n10046) );
  AOI22_X1 U11166 ( .A1(n5064), .A2(n10047), .B1(n10046), .B2(n9711), .ZN(
        P1_U3286) );
  OAI211_X1 U11167 ( .C1(n10078), .C2(n10049), .A(n10117), .B(n10048), .ZN(
        n10076) );
  INV_X1 U11168 ( .A(n10050), .ZN(n10051) );
  OAI22_X1 U11169 ( .A1(n10052), .A2(n10076), .B1(n10051), .B2(n10078), .ZN(
        n10066) );
  NAND2_X1 U11170 ( .A1(n10053), .A2(n10055), .ZN(n10058) );
  XNOR2_X1 U11171 ( .A(n10058), .B(n10054), .ZN(n10075) );
  INV_X1 U11172 ( .A(n6712), .ZN(n10093) );
  NAND2_X1 U11173 ( .A1(n10075), .A2(n10093), .ZN(n10065) );
  INV_X1 U11174 ( .A(n10055), .ZN(n10060) );
  INV_X1 U11175 ( .A(n10056), .ZN(n10057) );
  NAND2_X1 U11176 ( .A1(n10058), .A2(n10057), .ZN(n10059) );
  OAI211_X1 U11177 ( .C1(n10061), .C2(n10060), .A(n10059), .B(n10168), .ZN(
        n10063) );
  AOI22_X1 U11178 ( .A1(n10161), .A2(n6723), .B1(n10159), .B2(n6711), .ZN(
        n10062) );
  AND2_X1 U11179 ( .A1(n10063), .A2(n10062), .ZN(n10064) );
  NAND2_X1 U11180 ( .A1(n10065), .A2(n10064), .ZN(n10080) );
  AOI211_X1 U11181 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n10067), .A(n10066), .B(
        n10080), .ZN(n10070) );
  INV_X1 U11182 ( .A(n10075), .ZN(n10069) );
  OAI22_X1 U11183 ( .A1(n10070), .A2(n5064), .B1(n10069), .B2(n10068), .ZN(
        n10071) );
  INV_X1 U11184 ( .A(n10071), .ZN(n10072) );
  OAI21_X1 U11185 ( .B1(n6974), .B2(n9711), .A(n10072), .ZN(P1_U3290) );
  AND2_X1 U11186 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10073), .ZN(P1_U3292) );
  AND2_X1 U11187 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10073), .ZN(P1_U3293) );
  AND2_X1 U11188 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10073), .ZN(P1_U3294) );
  AND2_X1 U11189 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10073), .ZN(P1_U3295) );
  AND2_X1 U11190 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10073), .ZN(P1_U3296) );
  AND2_X1 U11191 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10073), .ZN(P1_U3297) );
  AND2_X1 U11192 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10073), .ZN(P1_U3298) );
  AND2_X1 U11193 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10073), .ZN(P1_U3299) );
  AND2_X1 U11194 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10073), .ZN(P1_U3300) );
  AND2_X1 U11195 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10073), .ZN(P1_U3301) );
  AND2_X1 U11196 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10073), .ZN(P1_U3302) );
  AND2_X1 U11197 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10073), .ZN(P1_U3303) );
  INV_X1 U11198 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n10432) );
  NOR2_X1 U11199 ( .A1(n10074), .A2(n10432), .ZN(P1_U3304) );
  AND2_X1 U11200 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10073), .ZN(P1_U3305) );
  AND2_X1 U11201 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10073), .ZN(P1_U3306) );
  AND2_X1 U11202 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10073), .ZN(P1_U3307) );
  AND2_X1 U11203 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10073), .ZN(P1_U3308) );
  INV_X1 U11204 ( .A(P1_D_REG_14__SCAN_IN), .ZN(n10489) );
  NOR2_X1 U11205 ( .A1(n10074), .A2(n10489), .ZN(P1_U3309) );
  AND2_X1 U11206 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10073), .ZN(P1_U3310) );
  INV_X1 U11207 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10297) );
  NOR2_X1 U11208 ( .A1(n10074), .A2(n10297), .ZN(P1_U3311) );
  INV_X1 U11209 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n10379) );
  NOR2_X1 U11210 ( .A1(n10074), .A2(n10379), .ZN(P1_U3312) );
  AND2_X1 U11211 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10073), .ZN(P1_U3313) );
  AND2_X1 U11212 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10073), .ZN(P1_U3314) );
  INV_X1 U11213 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n10332) );
  NOR2_X1 U11214 ( .A1(n10074), .A2(n10332), .ZN(P1_U3315) );
  INV_X1 U11215 ( .A(P1_D_REG_7__SCAN_IN), .ZN(n10306) );
  NOR2_X1 U11216 ( .A1(n10074), .A2(n10306), .ZN(P1_U3316) );
  INV_X1 U11217 ( .A(P1_D_REG_6__SCAN_IN), .ZN(n10472) );
  NOR2_X1 U11218 ( .A1(n10074), .A2(n10472), .ZN(P1_U3317) );
  INV_X1 U11219 ( .A(P1_D_REG_5__SCAN_IN), .ZN(n10319) );
  NOR2_X1 U11220 ( .A1(n10074), .A2(n10319), .ZN(P1_U3318) );
  AND2_X1 U11221 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10073), .ZN(P1_U3319) );
  AND2_X1 U11222 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10073), .ZN(P1_U3320) );
  INV_X1 U11223 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10498) );
  NOR2_X1 U11224 ( .A1(n10074), .A2(n10498), .ZN(P1_U3321) );
  INV_X1 U11225 ( .A(n10089), .ZN(n10125) );
  NAND2_X1 U11226 ( .A1(n10075), .A2(n10125), .ZN(n10077) );
  OAI211_X1 U11227 ( .C1(n10078), .C2(n10130), .A(n10077), .B(n10076), .ZN(
        n10079) );
  NOR2_X1 U11228 ( .A1(n10080), .A2(n10079), .ZN(n10151) );
  INV_X1 U11229 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10081) );
  AOI22_X1 U11230 ( .A1(n10588), .A2(n10151), .B1(n10081), .B2(n10586), .ZN(
        P1_U3457) );
  INV_X1 U11231 ( .A(n10090), .ZN(n10092) );
  AOI22_X1 U11232 ( .A1(n10161), .A2(n6729), .B1(n10159), .B2(n10082), .ZN(
        n10084) );
  OAI211_X1 U11233 ( .C1(n10132), .C2(n10085), .A(n10084), .B(n10083), .ZN(
        n10086) );
  INV_X1 U11234 ( .A(n10086), .ZN(n10088) );
  OAI211_X1 U11235 ( .C1(n10090), .C2(n10089), .A(n10088), .B(n10087), .ZN(
        n10091) );
  AOI21_X1 U11236 ( .B1(n10093), .B2(n10092), .A(n10091), .ZN(n10153) );
  INV_X1 U11237 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10094) );
  AOI22_X1 U11238 ( .A1(n10588), .A2(n10153), .B1(n10094), .B2(n10586), .ZN(
        P1_U3460) );
  INV_X1 U11239 ( .A(n10095), .ZN(n10097) );
  OAI22_X1 U11240 ( .A1(n10097), .A2(n10132), .B1(n10096), .B2(n10130), .ZN(
        n10100) );
  INV_X1 U11241 ( .A(n10098), .ZN(n10099) );
  AOI211_X1 U11242 ( .C1(n10128), .C2(n10101), .A(n10100), .B(n10099), .ZN(
        n10154) );
  AOI22_X1 U11243 ( .A1(n10588), .A2(n10154), .B1(n4800), .B2(n10586), .ZN(
        P1_U3463) );
  AOI21_X1 U11244 ( .B1(n10103), .B2(n10117), .A(n10102), .ZN(n10104) );
  OAI21_X1 U11245 ( .B1(n10105), .B2(n6712), .A(n10104), .ZN(n10107) );
  AOI211_X1 U11246 ( .C1(n10125), .C2(n10108), .A(n10107), .B(n10106), .ZN(
        n10155) );
  INV_X1 U11247 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10109) );
  AOI22_X1 U11248 ( .A1(n10588), .A2(n10155), .B1(n10109), .B2(n10586), .ZN(
        P1_U3466) );
  OAI21_X1 U11249 ( .B1(n5032), .B2(n10130), .A(n10110), .ZN(n10112) );
  AOI211_X1 U11250 ( .C1(n10128), .C2(n10113), .A(n10112), .B(n10111), .ZN(
        n10156) );
  INV_X1 U11251 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10114) );
  AOI22_X1 U11252 ( .A1(n10588), .A2(n10156), .B1(n10114), .B2(n10586), .ZN(
        P1_U3469) );
  INV_X1 U11253 ( .A(n10120), .ZN(n10124) );
  INV_X1 U11254 ( .A(n10115), .ZN(n10116) );
  AOI21_X1 U11255 ( .B1(n10118), .B2(n10117), .A(n10116), .ZN(n10119) );
  OAI21_X1 U11256 ( .B1(n10120), .B2(n6712), .A(n10119), .ZN(n10123) );
  INV_X1 U11257 ( .A(n10121), .ZN(n10122) );
  AOI211_X1 U11258 ( .C1(n10125), .C2(n10124), .A(n10123), .B(n10122), .ZN(
        n10157) );
  INV_X1 U11259 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n10126) );
  AOI22_X1 U11260 ( .A1(n10588), .A2(n10157), .B1(n10126), .B2(n10586), .ZN(
        P1_U3472) );
  AND3_X1 U11261 ( .A1(n10129), .A2(n10128), .A3(n10127), .ZN(n10135) );
  OAI22_X1 U11262 ( .A1(n10133), .A2(n10132), .B1(n10131), .B2(n10130), .ZN(
        n10134) );
  NOR3_X1 U11263 ( .A1(n10136), .A2(n10135), .A3(n10134), .ZN(n10174) );
  INV_X1 U11264 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10137) );
  AOI22_X1 U11265 ( .A1(n10588), .A2(n10174), .B1(n10137), .B2(n10586), .ZN(
        P1_U3478) );
  OAI22_X1 U11266 ( .A1(n10141), .A2(n10140), .B1(n10139), .B2(n10138), .ZN(
        n10143) );
  AOI211_X1 U11267 ( .C1(n10163), .C2(n10144), .A(n10143), .B(n10142), .ZN(
        n10146) );
  OAI211_X1 U11268 ( .C1(n10172), .C2(n10147), .A(n10146), .B(n10145), .ZN(
        n10148) );
  INV_X1 U11269 ( .A(n10148), .ZN(n10176) );
  INV_X1 U11270 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U11271 ( .A1(n10588), .A2(n10176), .B1(n10149), .B2(n10586), .ZN(
        P1_U3481) );
  AOI22_X1 U11272 ( .A1(n10177), .A2(n10151), .B1(n10150), .B2(n10175), .ZN(
        P1_U3524) );
  AOI22_X1 U11273 ( .A1(n10177), .A2(n10153), .B1(n10152), .B2(n10175), .ZN(
        P1_U3525) );
  AOI22_X1 U11274 ( .A1(n10177), .A2(n10154), .B1(n7060), .B2(n10175), .ZN(
        P1_U3526) );
  AOI22_X1 U11275 ( .A1(n10177), .A2(n10155), .B1(n7062), .B2(n10175), .ZN(
        P1_U3527) );
  AOI22_X1 U11276 ( .A1(n10177), .A2(n10156), .B1(n7064), .B2(n10175), .ZN(
        P1_U3528) );
  AOI22_X1 U11277 ( .A1(n10177), .A2(n10157), .B1(n10433), .B2(n10175), .ZN(
        P1_U3529) );
  AOI22_X1 U11278 ( .A1(n10161), .A2(n10160), .B1(n10159), .B2(n10158), .ZN(
        n10165) );
  NAND2_X1 U11279 ( .A1(n10163), .A2(n10162), .ZN(n10164) );
  NAND3_X1 U11280 ( .A1(n10166), .A2(n10165), .A3(n10164), .ZN(n10167) );
  AOI21_X1 U11281 ( .B1(n10169), .B2(n10168), .A(n10167), .ZN(n10170) );
  OAI21_X1 U11282 ( .B1(n10172), .B2(n10171), .A(n10170), .ZN(n10587) );
  OAI22_X1 U11283 ( .A1(n10175), .A2(n10587), .B1(P1_REG1_REG_7__SCAN_IN), 
        .B2(n10177), .ZN(n10173) );
  INV_X1 U11284 ( .A(n10173), .ZN(P1_U3530) );
  AOI22_X1 U11285 ( .A1(n10177), .A2(n10174), .B1(n7107), .B2(n10175), .ZN(
        P1_U3531) );
  AOI22_X1 U11286 ( .A1(n10177), .A2(n10176), .B1(n4599), .B2(n10175), .ZN(
        P1_U3532) );
  INV_X1 U11287 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n10320) );
  NOR2_X1 U11288 ( .A1(n10195), .A2(n10320), .ZN(P2_U3297) );
  NOR2_X1 U11289 ( .A1(n10195), .A2(n10180), .ZN(P2_U3298) );
  INV_X1 U11290 ( .A(P2_D_REG_29__SCAN_IN), .ZN(n10549) );
  NOR2_X1 U11291 ( .A1(n10195), .A2(n10549), .ZN(P2_U3299) );
  NOR2_X1 U11292 ( .A1(n10195), .A2(n10181), .ZN(P2_U3300) );
  NOR2_X1 U11293 ( .A1(n10195), .A2(n10182), .ZN(P2_U3301) );
  INV_X1 U11294 ( .A(P2_D_REG_26__SCAN_IN), .ZN(n10183) );
  NOR2_X1 U11295 ( .A1(n10195), .A2(n10183), .ZN(P2_U3302) );
  NOR2_X1 U11296 ( .A1(n10195), .A2(n10184), .ZN(P2_U3303) );
  INV_X1 U11297 ( .A(P2_D_REG_24__SCAN_IN), .ZN(n10185) );
  NOR2_X1 U11298 ( .A1(n10195), .A2(n10185), .ZN(P2_U3304) );
  NOR2_X1 U11299 ( .A1(n10195), .A2(n10347), .ZN(P2_U3305) );
  NOR2_X1 U11300 ( .A1(n10195), .A2(n10186), .ZN(P2_U3306) );
  NOR2_X1 U11301 ( .A1(n10195), .A2(n10339), .ZN(P2_U3307) );
  NOR2_X1 U11302 ( .A1(n10195), .A2(n10187), .ZN(P2_U3308) );
  INV_X1 U11303 ( .A(P2_D_REG_19__SCAN_IN), .ZN(n10188) );
  NOR2_X1 U11304 ( .A1(n10195), .A2(n10188), .ZN(P2_U3309) );
  INV_X1 U11305 ( .A(P2_D_REG_18__SCAN_IN), .ZN(n10189) );
  NOR2_X1 U11306 ( .A1(n10195), .A2(n10189), .ZN(P2_U3310) );
  INV_X1 U11307 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10190) );
  NOR2_X1 U11308 ( .A1(n10195), .A2(n10190), .ZN(P2_U3311) );
  INV_X1 U11309 ( .A(P2_D_REG_16__SCAN_IN), .ZN(n10191) );
  NOR2_X1 U11310 ( .A1(n10195), .A2(n10191), .ZN(P2_U3312) );
  NOR2_X1 U11311 ( .A1(n10195), .A2(n10476), .ZN(P2_U3313) );
  INV_X1 U11312 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10192) );
  NOR2_X1 U11313 ( .A1(n10195), .A2(n10192), .ZN(P2_U3314) );
  INV_X1 U11314 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10193) );
  NOR2_X1 U11315 ( .A1(n10195), .A2(n10193), .ZN(P2_U3315) );
  INV_X1 U11316 ( .A(P2_D_REG_12__SCAN_IN), .ZN(n10194) );
  NOR2_X1 U11317 ( .A1(n10195), .A2(n10194), .ZN(P2_U3316) );
  INV_X1 U11318 ( .A(P2_D_REG_11__SCAN_IN), .ZN(n10196) );
  NOR2_X1 U11319 ( .A1(n10195), .A2(n10196), .ZN(P2_U3317) );
  INV_X1 U11320 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10197) );
  NOR2_X1 U11321 ( .A1(n10195), .A2(n10197), .ZN(P2_U3318) );
  INV_X1 U11322 ( .A(P2_D_REG_9__SCAN_IN), .ZN(n10198) );
  NOR2_X1 U11323 ( .A1(n10195), .A2(n10198), .ZN(P2_U3319) );
  INV_X1 U11324 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10461) );
  NOR2_X1 U11325 ( .A1(n10195), .A2(n10461), .ZN(P2_U3320) );
  INV_X1 U11326 ( .A(P2_D_REG_7__SCAN_IN), .ZN(n10199) );
  NOR2_X1 U11327 ( .A1(n10195), .A2(n10199), .ZN(P2_U3321) );
  INV_X1 U11328 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10458) );
  NOR2_X1 U11329 ( .A1(n10195), .A2(n10458), .ZN(P2_U3322) );
  INV_X1 U11330 ( .A(P2_D_REG_5__SCAN_IN), .ZN(n10535) );
  NOR2_X1 U11331 ( .A1(n10195), .A2(n10535), .ZN(P2_U3323) );
  INV_X1 U11332 ( .A(P2_D_REG_4__SCAN_IN), .ZN(n10200) );
  NOR2_X1 U11333 ( .A1(n10195), .A2(n10200), .ZN(P2_U3324) );
  INV_X1 U11334 ( .A(P2_D_REG_3__SCAN_IN), .ZN(n10478) );
  NOR2_X1 U11335 ( .A1(n10195), .A2(n10478), .ZN(P2_U3325) );
  INV_X1 U11336 ( .A(P2_D_REG_2__SCAN_IN), .ZN(n10505) );
  NOR2_X1 U11337 ( .A1(n10195), .A2(n10505), .ZN(P2_U3326) );
  OAI22_X1 U11338 ( .A1(P2_D_REG_0__SCAN_IN), .A2(n10195), .B1(n10201), .B2(
        n10203), .ZN(n10202) );
  INV_X1 U11339 ( .A(n10202), .ZN(P2_U3437) );
  OAI22_X1 U11340 ( .A1(P2_D_REG_1__SCAN_IN), .A2(n10195), .B1(n10204), .B2(
        n10203), .ZN(n10205) );
  INV_X1 U11341 ( .A(n10205), .ZN(P2_U3438) );
  AOI22_X1 U11342 ( .A1(n10208), .A2(n10243), .B1(n10207), .B2(n10206), .ZN(
        n10209) );
  AND2_X1 U11343 ( .A1(n10210), .A2(n10209), .ZN(n10255) );
  INV_X1 U11344 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10211) );
  AOI22_X1 U11345 ( .A1(n10254), .A2(n10255), .B1(n10211), .B2(n10253), .ZN(
        P2_U3451) );
  INV_X1 U11346 ( .A(n10212), .ZN(n10213) );
  OAI21_X1 U11347 ( .B1(n10214), .B2(n10245), .A(n10213), .ZN(n10216) );
  AOI211_X1 U11348 ( .C1(n10243), .C2(n10217), .A(n10216), .B(n10215), .ZN(
        n10256) );
  INV_X1 U11349 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10218) );
  AOI22_X1 U11350 ( .A1(n10254), .A2(n10256), .B1(n10218), .B2(n10253), .ZN(
        P2_U3454) );
  INV_X1 U11351 ( .A(n10219), .ZN(n10220) );
  OAI211_X1 U11352 ( .C1(n10222), .C2(n10245), .A(n10221), .B(n10220), .ZN(
        n10223) );
  AOI21_X1 U11353 ( .B1(n10243), .B2(n10224), .A(n10223), .ZN(n10257) );
  AOI22_X1 U11354 ( .A1(n10254), .A2(n10257), .B1(n5168), .B2(n10253), .ZN(
        P2_U3457) );
  INV_X1 U11355 ( .A(n10225), .ZN(n10226) );
  OAI21_X1 U11356 ( .B1(n10227), .B2(n10245), .A(n10226), .ZN(n10229) );
  AOI211_X1 U11357 ( .C1(n10243), .C2(n10230), .A(n10229), .B(n10228), .ZN(
        n10258) );
  AOI22_X1 U11358 ( .A1(n10254), .A2(n10258), .B1(n5205), .B2(n10253), .ZN(
        P2_U3463) );
  INV_X1 U11359 ( .A(n10231), .ZN(n10236) );
  OAI22_X1 U11360 ( .A1(n10233), .A2(n10246), .B1(n10232), .B2(n10245), .ZN(
        n10235) );
  AOI211_X1 U11361 ( .C1(n10243), .C2(n10236), .A(n10235), .B(n10234), .ZN(
        n10259) );
  AOI22_X1 U11362 ( .A1(n10254), .A2(n10259), .B1(n5279), .B2(n10253), .ZN(
        P2_U3469) );
  OAI22_X1 U11363 ( .A1(n10238), .A2(n10246), .B1(n7563), .B2(n10245), .ZN(
        n10241) );
  INV_X1 U11364 ( .A(n10239), .ZN(n10240) );
  AOI211_X1 U11365 ( .C1(n10243), .C2(n10242), .A(n10241), .B(n10240), .ZN(
        n10260) );
  AOI22_X1 U11366 ( .A1(n10254), .A2(n10260), .B1(n5305), .B2(n10253), .ZN(
        P2_U3472) );
  OAI22_X1 U11367 ( .A1(n10247), .A2(n10246), .B1(n4842), .B2(n10245), .ZN(
        n10248) );
  AOI21_X1 U11368 ( .B1(n10250), .B2(n10249), .A(n10248), .ZN(n10251) );
  AND2_X1 U11369 ( .A1(n10252), .A2(n10251), .ZN(n10262) );
  AOI22_X1 U11370 ( .A1(n10254), .A2(n10262), .B1(n5333), .B2(n10253), .ZN(
        P2_U3475) );
  AOI22_X1 U11371 ( .A1(n10263), .A2(n10255), .B1(n7240), .B2(n10261), .ZN(
        P2_U3520) );
  AOI22_X1 U11372 ( .A1(n10263), .A2(n10256), .B1(n6651), .B2(n10261), .ZN(
        P2_U3521) );
  AOI22_X1 U11373 ( .A1(n10263), .A2(n10257), .B1(n6650), .B2(n10261), .ZN(
        P2_U3522) );
  AOI22_X1 U11374 ( .A1(n10263), .A2(n10258), .B1(n6658), .B2(n10261), .ZN(
        P2_U3524) );
  AOI22_X1 U11375 ( .A1(n10263), .A2(n10259), .B1(n6664), .B2(n10261), .ZN(
        P2_U3526) );
  AOI22_X1 U11376 ( .A1(n10263), .A2(n10260), .B1(n6667), .B2(n10261), .ZN(
        P2_U3527) );
  AOI22_X1 U11377 ( .A1(n10263), .A2(n10262), .B1(n6670), .B2(n10261), .ZN(
        P2_U3528) );
  INV_X1 U11378 ( .A(n10264), .ZN(n10265) );
  NAND2_X1 U11379 ( .A1(n10266), .A2(n10265), .ZN(n10267) );
  XNOR2_X1 U11380 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10267), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11381 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11382 ( .B1(n10270), .B2(n10269), .A(n10268), .ZN(ADD_1071_U56) );
  OAI21_X1 U11383 ( .B1(n10273), .B2(n10272), .A(n10271), .ZN(ADD_1071_U57) );
  OAI21_X1 U11384 ( .B1(n10276), .B2(n10275), .A(n10274), .ZN(ADD_1071_U58) );
  OAI21_X1 U11385 ( .B1(n10279), .B2(n10278), .A(n10277), .ZN(ADD_1071_U59) );
  OAI21_X1 U11386 ( .B1(n10282), .B2(n10281), .A(n10280), .ZN(ADD_1071_U60) );
  OAI21_X1 U11387 ( .B1(n10285), .B2(n10284), .A(n10283), .ZN(ADD_1071_U61) );
  AOI21_X1 U11388 ( .B1(n10288), .B2(n10287), .A(n10286), .ZN(ADD_1071_U62) );
  AOI21_X1 U11389 ( .B1(n10291), .B2(n10290), .A(n10289), .ZN(ADD_1071_U63) );
  INV_X1 U11390 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10293) );
  AOI22_X1 U11391 ( .A1(n10293), .A2(keyinput51), .B1(n5856), .B2(keyinput47), 
        .ZN(n10292) );
  OAI221_X1 U11392 ( .B1(n10293), .B2(keyinput51), .C1(n5856), .C2(keyinput47), 
        .A(n10292), .ZN(n10304) );
  AOI22_X1 U11393 ( .A1(n10296), .A2(keyinput87), .B1(n10295), .B2(keyinput110), .ZN(n10294) );
  OAI221_X1 U11394 ( .B1(n10296), .B2(keyinput87), .C1(n10295), .C2(
        keyinput110), .A(n10294), .ZN(n10303) );
  XNOR2_X1 U11395 ( .A(n10297), .B(keyinput15), .ZN(n10302) );
  XNOR2_X1 U11396 ( .A(P2_IR_REG_2__SCAN_IN), .B(keyinput7), .ZN(n10300) );
  XNOR2_X1 U11397 ( .A(P1_IR_REG_11__SCAN_IN), .B(keyinput125), .ZN(n10299) );
  XNOR2_X1 U11398 ( .A(P1_REG0_REG_20__SCAN_IN), .B(keyinput40), .ZN(n10298)
         );
  NAND3_X1 U11399 ( .A1(n10300), .A2(n10299), .A3(n10298), .ZN(n10301) );
  NOR4_X1 U11400 ( .A1(n10304), .A2(n10303), .A3(n10302), .A4(n10301), .ZN(
        n10585) );
  AOI22_X1 U11401 ( .A1(n10306), .A2(keyinput39), .B1(keyinput12), .B2(n6154), 
        .ZN(n10305) );
  OAI221_X1 U11402 ( .B1(n10306), .B2(keyinput39), .C1(n6154), .C2(keyinput12), 
        .A(n10305), .ZN(n10314) );
  NAND2_X1 U11403 ( .A1(n6305), .A2(keyinput102), .ZN(n10307) );
  OAI221_X1 U11404 ( .B1(n5805), .B2(keyinput9), .C1(n6305), .C2(keyinput102), 
        .A(n10307), .ZN(n10313) );
  XOR2_X1 U11405 ( .A(n7911), .B(keyinput100), .Z(n10311) );
  XNOR2_X1 U11406 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput1), .ZN(n10310) );
  XNOR2_X1 U11407 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput76), .ZN(n10309) );
  XNOR2_X1 U11408 ( .A(P1_REG1_REG_15__SCAN_IN), .B(keyinput78), .ZN(n10308)
         );
  NAND4_X1 U11409 ( .A1(n10311), .A2(n10310), .A3(n10309), .A4(n10308), .ZN(
        n10312) );
  NOR3_X1 U11410 ( .A1(n10314), .A2(n10313), .A3(n10312), .ZN(n10584) );
  AOI22_X1 U11411 ( .A1(n10316), .A2(keyinput34), .B1(keyinput118), .B2(n9611), 
        .ZN(n10315) );
  OAI221_X1 U11412 ( .B1(n10316), .B2(keyinput34), .C1(n9611), .C2(keyinput118), .A(n10315), .ZN(n10325) );
  INV_X1 U11413 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n10438) );
  AOI22_X1 U11414 ( .A1(n10436), .A2(keyinput45), .B1(n10438), .B2(keyinput122), .ZN(n10317) );
  OAI221_X1 U11415 ( .B1(n10436), .B2(keyinput45), .C1(n10438), .C2(
        keyinput122), .A(n10317), .ZN(n10324) );
  AOI22_X1 U11416 ( .A1(n10320), .A2(keyinput3), .B1(n10319), .B2(keyinput82), 
        .ZN(n10318) );
  OAI221_X1 U11417 ( .B1(n10320), .B2(keyinput3), .C1(n10319), .C2(keyinput82), 
        .A(n10318), .ZN(n10323) );
  AOI22_X1 U11418 ( .A1(n10435), .A2(keyinput54), .B1(keyinput105), .B2(n6657), 
        .ZN(n10321) );
  OAI221_X1 U11419 ( .B1(n10435), .B2(keyinput54), .C1(n6657), .C2(keyinput105), .A(n10321), .ZN(n10322) );
  NOR4_X1 U11420 ( .A1(n10325), .A2(n10324), .A3(n10323), .A4(n10322), .ZN(
        n10391) );
  AOI22_X1 U11421 ( .A1(n10432), .A2(keyinput89), .B1(keyinput109), .B2(n10327), .ZN(n10326) );
  OAI221_X1 U11422 ( .B1(n10432), .B2(keyinput89), .C1(n10327), .C2(
        keyinput109), .A(n10326), .ZN(n10337) );
  INV_X1 U11423 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U11424 ( .A1(n10330), .A2(keyinput97), .B1(keyinput18), .B2(n10329), 
        .ZN(n10328) );
  OAI221_X1 U11425 ( .B1(n10330), .B2(keyinput97), .C1(n10329), .C2(keyinput18), .A(n10328), .ZN(n10336) );
  AOI22_X1 U11426 ( .A1(n10437), .A2(keyinput115), .B1(n10332), .B2(keyinput95), .ZN(n10331) );
  OAI221_X1 U11427 ( .B1(n10437), .B2(keyinput115), .C1(n10332), .C2(
        keyinput95), .A(n10331), .ZN(n10335) );
  INV_X1 U11428 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10431) );
  AOI22_X1 U11429 ( .A1(n10431), .A2(keyinput67), .B1(keyinput44), .B2(n5566), 
        .ZN(n10333) );
  OAI221_X1 U11430 ( .B1(n10431), .B2(keyinput67), .C1(n5566), .C2(keyinput44), 
        .A(n10333), .ZN(n10334) );
  NOR4_X1 U11431 ( .A1(n10337), .A2(n10336), .A3(n10335), .A4(n10334), .ZN(
        n10390) );
  AOI22_X1 U11432 ( .A1(n10340), .A2(keyinput99), .B1(keyinput120), .B2(n10339), .ZN(n10338) );
  OAI221_X1 U11433 ( .B1(n10340), .B2(keyinput99), .C1(n10339), .C2(
        keyinput120), .A(n10338), .ZN(n10351) );
  AOI22_X1 U11434 ( .A1(n7448), .A2(keyinput17), .B1(keyinput72), .B2(n10342), 
        .ZN(n10341) );
  OAI221_X1 U11435 ( .B1(n7448), .B2(keyinput17), .C1(n10342), .C2(keyinput72), 
        .A(n10341), .ZN(n10350) );
  AOI22_X1 U11436 ( .A1(n10398), .A2(keyinput119), .B1(n10344), .B2(keyinput4), 
        .ZN(n10343) );
  OAI221_X1 U11437 ( .B1(n10398), .B2(keyinput119), .C1(n10344), .C2(keyinput4), .A(n10343), .ZN(n10349) );
  AOI22_X1 U11438 ( .A1(n10347), .A2(keyinput5), .B1(n10346), .B2(keyinput38), 
        .ZN(n10345) );
  OAI221_X1 U11439 ( .B1(n10347), .B2(keyinput5), .C1(n10346), .C2(keyinput38), 
        .A(n10345), .ZN(n10348) );
  NOR4_X1 U11440 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        n10389) );
  INV_X1 U11441 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n10605) );
  OAI22_X1 U11442 ( .A1(n10446), .A2(keyinput104), .B1(n10605), .B2(keyinput8), 
        .ZN(n10352) );
  AOI221_X1 U11443 ( .B1(n10446), .B2(keyinput104), .C1(keyinput8), .C2(n10605), .A(n10352), .ZN(n10387) );
  AOI22_X1 U11444 ( .A1(n9492), .A2(keyinput94), .B1(n10445), .B2(keyinput53), 
        .ZN(n10353) );
  OAI221_X1 U11445 ( .B1(n9492), .B2(keyinput94), .C1(n10445), .C2(keyinput53), 
        .A(n10353), .ZN(n10354) );
  INV_X1 U11446 ( .A(n10354), .ZN(n10373) );
  XNOR2_X1 U11447 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput107), .ZN(n10358)
         );
  XNOR2_X1 U11448 ( .A(P1_IR_REG_28__SCAN_IN), .B(keyinput83), .ZN(n10357) );
  XNOR2_X1 U11449 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput43), .ZN(n10356) );
  XNOR2_X1 U11450 ( .A(P1_REG3_REG_6__SCAN_IN), .B(keyinput93), .ZN(n10355) );
  NAND4_X1 U11451 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10364) );
  XNOR2_X1 U11452 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(keyinput116), .ZN(n10362)
         );
  XNOR2_X1 U11453 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(keyinput73), .ZN(n10361)
         );
  XNOR2_X1 U11454 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(keyinput70), .ZN(n10360)
         );
  XNOR2_X1 U11455 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(keyinput84), .ZN(n10359)
         );
  NAND4_X1 U11456 ( .A1(n10362), .A2(n10361), .A3(n10360), .A4(n10359), .ZN(
        n10363) );
  NOR2_X1 U11457 ( .A1(n10364), .A2(n10363), .ZN(n10372) );
  INV_X1 U11458 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n10365) );
  XNOR2_X1 U11459 ( .A(keyinput114), .B(n10365), .ZN(n10367) );
  XNOR2_X1 U11460 ( .A(keyinput31), .B(n7870), .ZN(n10366) );
  NOR2_X1 U11461 ( .A1(n10367), .A2(n10366), .ZN(n10371) );
  XNOR2_X1 U11462 ( .A(keyinput68), .B(n6627), .ZN(n10369) );
  XNOR2_X1 U11463 ( .A(keyinput79), .B(n5079), .ZN(n10368) );
  NOR2_X1 U11464 ( .A1(n10369), .A2(n10368), .ZN(n10370) );
  AND4_X1 U11465 ( .A1(n10373), .A2(n10372), .A3(n10371), .A4(n10370), .ZN(
        n10386) );
  AOI22_X1 U11466 ( .A1(n8046), .A2(keyinput24), .B1(keyinput63), .B2(n5305), 
        .ZN(n10374) );
  OAI221_X1 U11467 ( .B1(n8046), .B2(keyinput24), .C1(n5305), .C2(keyinput63), 
        .A(n10374), .ZN(n10377) );
  AOI22_X1 U11468 ( .A1(n10397), .A2(keyinput19), .B1(keyinput28), .B2(n5650), 
        .ZN(n10375) );
  OAI221_X1 U11469 ( .B1(n10397), .B2(keyinput19), .C1(n5650), .C2(keyinput28), 
        .A(n10375), .ZN(n10376) );
  NOR2_X1 U11470 ( .A1(n10377), .A2(n10376), .ZN(n10385) );
  AOI22_X1 U11471 ( .A1(n10379), .A2(keyinput6), .B1(keyinput41), .B2(n6974), 
        .ZN(n10378) );
  OAI221_X1 U11472 ( .B1(n10379), .B2(keyinput6), .C1(n6974), .C2(keyinput41), 
        .A(n10378), .ZN(n10383) );
  AOI22_X1 U11473 ( .A1(n10381), .A2(keyinput126), .B1(n10433), .B2(keyinput69), .ZN(n10380) );
  OAI221_X1 U11474 ( .B1(n10381), .B2(keyinput126), .C1(n10433), .C2(
        keyinput69), .A(n10380), .ZN(n10382) );
  NOR2_X1 U11475 ( .A1(n10383), .A2(n10382), .ZN(n10384) );
  AND4_X1 U11476 ( .A1(n10387), .A2(n10386), .A3(n10385), .A4(n10384), .ZN(
        n10388) );
  AND4_X1 U11477 ( .A1(n10391), .A2(n10390), .A3(n10389), .A4(n10388), .ZN(
        n10583) );
  INV_X1 U11478 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n10459) );
  NAND4_X1 U11479 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_REG2_REG_31__SCAN_IN), 
        .A3(n10459), .A4(n10479), .ZN(n10396) );
  NAND4_X1 U11480 ( .A1(P1_REG0_REG_10__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), 
        .A3(P2_REG2_REG_19__SCAN_IN), .A4(P2_REG2_REG_31__SCAN_IN), .ZN(n10395) );
  NAND4_X1 U11481 ( .A1(n10392), .A2(P1_IR_REG_16__SCAN_IN), .A3(SI_14_), .A4(
        P1_IR_REG_29__SCAN_IN), .ZN(n10394) );
  NAND4_X1 U11482 ( .A1(n10488), .A2(P2_REG1_REG_7__SCAN_IN), .A3(
        P1_REG2_REG_4__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n10393) );
  NOR4_X1 U11483 ( .A1(n10396), .A2(n10395), .A3(n10394), .A4(n10393), .ZN(
        n10416) );
  NAND4_X1 U11484 ( .A1(P2_DATAO_REG_2__SCAN_IN), .A2(P1_REG2_REG_12__SCAN_IN), 
        .A3(P2_REG0_REG_7__SCAN_IN), .A4(P2_REG2_REG_6__SCAN_IN), .ZN(n10402)
         );
  NAND4_X1 U11485 ( .A1(P2_ADDR_REG_19__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), 
        .A3(n10397), .A4(n5650), .ZN(n10401) );
  NAND4_X1 U11486 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(P1_REG2_REG_20__SCAN_IN), 
        .A3(P2_D_REG_8__SCAN_IN), .A4(n10398), .ZN(n10400) );
  NAND4_X1 U11487 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), 
        .A3(P2_D_REG_23__SCAN_IN), .A4(n7448), .ZN(n10399) );
  NOR4_X1 U11488 ( .A1(n10402), .A2(n10401), .A3(n10400), .A4(n10399), .ZN(
        n10415) );
  NAND4_X1 U11489 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P2_REG0_REG_25__SCAN_IN), 
        .A3(n10562), .A4(n9912), .ZN(n10405) );
  NAND4_X1 U11490 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG0_REG_31__SCAN_IN), 
        .A3(n10550), .A4(n10554), .ZN(n10404) );
  NAND4_X1 U11491 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n10566), .A3(n10567), 
        .A4(n10564), .ZN(n10403) );
  NOR4_X1 U11492 ( .A1(n10406), .A2(n10405), .A3(n10404), .A4(n10403), .ZN(
        n10414) );
  INV_X1 U11493 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10540) );
  INV_X1 U11494 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n10407) );
  NAND4_X1 U11495 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(P2_REG3_REG_19__SCAN_IN), 
        .A3(n10540), .A4(n10407), .ZN(n10408) );
  NOR3_X1 U11496 ( .A1(n10503), .A2(P1_DATAO_REG_5__SCAN_IN), .A3(n10408), 
        .ZN(n10409) );
  NAND3_X1 U11497 ( .A1(n10409), .A2(P2_REG0_REG_12__SCAN_IN), .A3(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n10412) );
  NAND4_X1 U11498 ( .A1(n10526), .A2(n4656), .A3(n6661), .A4(n8452), .ZN(
        n10411) );
  NAND4_X1 U11499 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_DATAO_REG_10__SCAN_IN), 
        .A3(P2_REG1_REG_10__SCAN_IN), .A4(n10527), .ZN(n10410) );
  NOR3_X1 U11500 ( .A1(n10412), .A2(n10411), .A3(n10410), .ZN(n10413) );
  NAND4_X1 U11501 ( .A1(n10416), .A2(n10415), .A3(n10414), .A4(n10413), .ZN(
        n10456) );
  INV_X1 U11502 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10603) );
  NAND4_X1 U11503 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P2_ADDR_REG_6__SCAN_IN), 
        .A3(P1_ADDR_REG_18__SCAN_IN), .A4(n10603), .ZN(n10422) );
  NAND4_X1 U11504 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P2_ADDR_REG_15__SCAN_IN), 
        .A3(P1_ADDR_REG_10__SCAN_IN), .A4(n7911), .ZN(n10421) );
  NAND4_X1 U11505 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_REG2_REG_22__SCAN_IN), 
        .A3(P1_REG1_REG_20__SCAN_IN), .A4(P2_REG3_REG_22__SCAN_IN), .ZN(n10417) );
  NOR3_X1 U11506 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n10417), .A3(
        P1_D_REG_1__SCAN_IN), .ZN(n10419) );
  NAND3_X1 U11507 ( .A1(n10419), .A2(P1_D_REG_7__SCAN_IN), .A3(n10418), .ZN(
        n10420) );
  NOR3_X1 U11508 ( .A1(n10422), .A2(n10421), .A3(n10420), .ZN(n10454) );
  NAND4_X1 U11509 ( .A1(n10423), .A2(P2_REG3_REG_13__SCAN_IN), .A3(
        P1_ADDR_REG_1__SCAN_IN), .A4(P1_ADDR_REG_4__SCAN_IN), .ZN(n10428) );
  NOR2_X1 U11510 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .ZN(n10425) );
  NAND3_X1 U11511 ( .A1(n10426), .A2(n10425), .A3(n10424), .ZN(n10427) );
  NOR4_X1 U11512 ( .A1(n10428), .A2(n10427), .A3(P1_IR_REG_9__SCAN_IN), .A4(
        P1_REG3_REG_27__SCAN_IN), .ZN(n10430) );
  AND2_X1 U11513 ( .A1(n10430), .A2(n10429), .ZN(n10453) );
  NAND4_X1 U11514 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(P2_REG0_REG_26__SCAN_IN), 
        .A3(n10432), .A4(n10431), .ZN(n10442) );
  NAND4_X1 U11515 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG0_REG_23__SCAN_IN), 
        .A3(n10434), .A4(n10433), .ZN(n10441) );
  NAND4_X1 U11516 ( .A1(P1_REG2_REG_21__SCAN_IN), .A2(P1_DATAO_REG_13__SCAN_IN), .A3(n10435), .A4(n6657), .ZN(n10440) );
  NAND4_X1 U11517 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10438), .A3(n10437), .A4(
        n10436), .ZN(n10439) );
  NOR4_X1 U11518 ( .A1(n10442), .A2(n10441), .A3(n10440), .A4(n10439), .ZN(
        n10452) );
  NAND4_X1 U11519 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .A3(P1_REG2_REG_1__SCAN_IN), .A4(P2_IR_REG_20__SCAN_IN), .ZN(n10450)
         );
  INV_X1 U11520 ( .A(P1_REG0_REG_20__SCAN_IN), .ZN(n10443) );
  NAND4_X1 U11521 ( .A1(P1_REG2_REG_19__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), 
        .A3(n5856), .A4(n10443), .ZN(n10449) );
  NAND4_X1 U11522 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_REG3_REG_6__SCAN_IN), 
        .A3(n10445), .A4(n10444), .ZN(n10448) );
  NAND4_X1 U11523 ( .A1(P2_DATAO_REG_3__SCAN_IN), .A2(n10446), .A3(n9492), 
        .A4(n6627), .ZN(n10447) );
  NOR4_X1 U11524 ( .A1(n10450), .A2(n10449), .A3(n10448), .A4(n10447), .ZN(
        n10451) );
  NAND4_X1 U11525 ( .A1(n10454), .A2(n10453), .A3(n10452), .A4(n10451), .ZN(
        n10455) );
  OAI21_X1 U11526 ( .B1(n10456), .B2(n10455), .A(P2_IR_REG_23__SCAN_IN), .ZN(
        n10581) );
  AOI22_X1 U11527 ( .A1(n10459), .A2(keyinput57), .B1(n10458), .B2(keyinput96), 
        .ZN(n10457) );
  OAI221_X1 U11528 ( .B1(n10459), .B2(keyinput57), .C1(n10458), .C2(keyinput96), .A(n10457), .ZN(n10470) );
  AOI22_X1 U11529 ( .A1(n9627), .A2(keyinput86), .B1(keyinput124), .B2(n10461), 
        .ZN(n10460) );
  OAI221_X1 U11530 ( .B1(n9627), .B2(keyinput86), .C1(n10461), .C2(keyinput124), .A(n10460), .ZN(n10469) );
  INV_X1 U11531 ( .A(SI_14_), .ZN(n10463) );
  AOI22_X1 U11532 ( .A1(n10464), .A2(keyinput91), .B1(n10463), .B2(keyinput108), .ZN(n10462) );
  OAI221_X1 U11533 ( .B1(n10464), .B2(keyinput91), .C1(n10463), .C2(
        keyinput108), .A(n10462), .ZN(n10468) );
  XOR2_X1 U11534 ( .A(n5864), .B(keyinput32), .Z(n10466) );
  XNOR2_X1 U11535 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput80), .ZN(n10465) );
  NAND2_X1 U11536 ( .A1(n10466), .A2(n10465), .ZN(n10467) );
  NOR4_X1 U11537 ( .A1(n10470), .A2(n10469), .A3(n10468), .A4(n10467), .ZN(
        n10521) );
  INV_X1 U11538 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n10473) );
  AOI22_X1 U11539 ( .A1(n10473), .A2(keyinput127), .B1(n10472), .B2(keyinput50), .ZN(n10471) );
  OAI221_X1 U11540 ( .B1(n10473), .B2(keyinput127), .C1(n10472), .C2(
        keyinput50), .A(n10471), .ZN(n10486) );
  AOI22_X1 U11541 ( .A1(n10476), .A2(keyinput11), .B1(keyinput13), .B2(n10475), 
        .ZN(n10474) );
  OAI221_X1 U11542 ( .B1(n10476), .B2(keyinput11), .C1(n10475), .C2(keyinput13), .A(n10474), .ZN(n10485) );
  AOI22_X1 U11543 ( .A1(n10479), .A2(keyinput65), .B1(n10478), .B2(keyinput30), 
        .ZN(n10477) );
  OAI221_X1 U11544 ( .B1(n10479), .B2(keyinput65), .C1(n10478), .C2(keyinput30), .A(n10477), .ZN(n10484) );
  AOI22_X1 U11545 ( .A1(n10482), .A2(keyinput113), .B1(keyinput27), .B2(n10481), .ZN(n10480) );
  OAI221_X1 U11546 ( .B1(n10482), .B2(keyinput113), .C1(n10481), .C2(
        keyinput27), .A(n10480), .ZN(n10483) );
  NOR4_X1 U11547 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n10520) );
  XNOR2_X1 U11548 ( .A(n10487), .B(keyinput103), .ZN(n10492) );
  XNOR2_X1 U11549 ( .A(n10488), .B(keyinput71), .ZN(n10491) );
  XNOR2_X1 U11550 ( .A(keyinput81), .B(n10489), .ZN(n10490) );
  NOR3_X1 U11551 ( .A1(n10492), .A2(n10491), .A3(n10490), .ZN(n10495) );
  XOR2_X1 U11552 ( .A(n5468), .B(keyinput55), .Z(n10494) );
  XNOR2_X1 U11553 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(keyinput26), .ZN(n10493)
         );
  NAND3_X1 U11554 ( .A1(n10495), .A2(n10494), .A3(n10493), .ZN(n10501) );
  AOI22_X1 U11555 ( .A1(n10497), .A2(keyinput117), .B1(keyinput23), .B2(n6667), 
        .ZN(n10496) );
  OAI221_X1 U11556 ( .B1(n10497), .B2(keyinput117), .C1(n6667), .C2(keyinput23), .A(n10496), .ZN(n10500) );
  XNOR2_X1 U11557 ( .A(n10498), .B(keyinput14), .ZN(n10499) );
  NOR3_X1 U11558 ( .A1(n10501), .A2(n10500), .A3(n10499), .ZN(n10519) );
  AOI22_X1 U11559 ( .A1(n10504), .A2(keyinput106), .B1(n10503), .B2(
        keyinput112), .ZN(n10502) );
  OAI221_X1 U11560 ( .B1(n10504), .B2(keyinput106), .C1(n10503), .C2(
        keyinput112), .A(n10502), .ZN(n10509) );
  XNOR2_X1 U11561 ( .A(n10505), .B(keyinput98), .ZN(n10508) );
  XNOR2_X1 U11562 ( .A(n10506), .B(keyinput66), .ZN(n10507) );
  OR3_X1 U11563 ( .A1(n10509), .A2(n10508), .A3(n10507), .ZN(n10517) );
  INV_X1 U11564 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n10511) );
  AOI22_X1 U11565 ( .A1(n10512), .A2(keyinput0), .B1(n10511), .B2(keyinput62), 
        .ZN(n10510) );
  OAI221_X1 U11566 ( .B1(n10512), .B2(keyinput0), .C1(n10511), .C2(keyinput62), 
        .A(n10510), .ZN(n10516) );
  INV_X1 U11567 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n10591) );
  AOI22_X1 U11568 ( .A1(n10591), .A2(keyinput10), .B1(n10514), .B2(keyinput37), 
        .ZN(n10513) );
  OAI221_X1 U11569 ( .B1(n10591), .B2(keyinput10), .C1(n10514), .C2(keyinput37), .A(n10513), .ZN(n10515) );
  NOR3_X1 U11570 ( .A1(n10517), .A2(n10516), .A3(n10515), .ZN(n10518) );
  NAND4_X1 U11571 ( .A1(n10521), .A2(n10520), .A3(n10519), .A4(n10518), .ZN(
        n10580) );
  AOI22_X1 U11572 ( .A1(n8452), .A2(keyinput90), .B1(n6661), .B2(keyinput88), 
        .ZN(n10522) );
  OAI221_X1 U11573 ( .B1(n8452), .B2(keyinput90), .C1(n6661), .C2(keyinput88), 
        .A(n10522), .ZN(n10533) );
  AOI22_X1 U11574 ( .A1(n10524), .A2(keyinput85), .B1(P2_U3152), .B2(keyinput2), .ZN(n10523) );
  OAI221_X1 U11575 ( .B1(n10524), .B2(keyinput85), .C1(P2_U3152), .C2(
        keyinput2), .A(n10523), .ZN(n10532) );
  AOI22_X1 U11576 ( .A1(n10527), .A2(keyinput74), .B1(n10526), .B2(keyinput25), 
        .ZN(n10525) );
  OAI221_X1 U11577 ( .B1(n10527), .B2(keyinput74), .C1(n10526), .C2(keyinput25), .A(n10525), .ZN(n10531) );
  XNOR2_X1 U11578 ( .A(P1_REG3_REG_20__SCAN_IN), .B(keyinput61), .ZN(n10529)
         );
  XNOR2_X1 U11579 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput60), .ZN(n10528) );
  NAND2_X1 U11580 ( .A1(n10529), .A2(n10528), .ZN(n10530) );
  NOR4_X1 U11581 ( .A1(n10533), .A2(n10532), .A3(n10531), .A4(n10530), .ZN(
        n10578) );
  INV_X1 U11582 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U11583 ( .A1(n10536), .A2(keyinput29), .B1(n10535), .B2(keyinput101), .ZN(n10534) );
  OAI221_X1 U11584 ( .B1(n10536), .B2(keyinput29), .C1(n10535), .C2(
        keyinput101), .A(n10534), .ZN(n10547) );
  AOI22_X1 U11585 ( .A1(n10603), .A2(keyinput77), .B1(n10538), .B2(keyinput58), 
        .ZN(n10537) );
  OAI221_X1 U11586 ( .B1(n10603), .B2(keyinput77), .C1(n10538), .C2(keyinput58), .A(n10537), .ZN(n10546) );
  AOI22_X1 U11587 ( .A1(n10541), .A2(keyinput35), .B1(n10540), .B2(keyinput111), .ZN(n10539) );
  OAI221_X1 U11588 ( .B1(n10541), .B2(keyinput35), .C1(n10540), .C2(
        keyinput111), .A(n10539), .ZN(n10545) );
  XNOR2_X1 U11589 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(keyinput123), .ZN(n10543)
         );
  XNOR2_X1 U11590 ( .A(P1_REG1_REG_30__SCAN_IN), .B(keyinput42), .ZN(n10542)
         );
  NAND2_X1 U11591 ( .A1(n10543), .A2(n10542), .ZN(n10544) );
  NOR4_X1 U11592 ( .A1(n10547), .A2(n10546), .A3(n10545), .A4(n10544), .ZN(
        n10577) );
  AOI22_X1 U11593 ( .A1(n10550), .A2(keyinput20), .B1(keyinput75), .B2(n10549), 
        .ZN(n10548) );
  OAI221_X1 U11594 ( .B1(n10550), .B2(keyinput20), .C1(n10549), .C2(keyinput75), .A(n10548), .ZN(n10560) );
  AOI22_X1 U11595 ( .A1(n10426), .A2(keyinput92), .B1(keyinput64), .B2(n6112), 
        .ZN(n10551) );
  OAI221_X1 U11596 ( .B1(n10426), .B2(keyinput92), .C1(n6112), .C2(keyinput64), 
        .A(n10551), .ZN(n10559) );
  AOI22_X1 U11597 ( .A1(n10554), .A2(keyinput56), .B1(n10553), .B2(keyinput36), 
        .ZN(n10552) );
  OAI221_X1 U11598 ( .B1(n10554), .B2(keyinput56), .C1(n10553), .C2(keyinput36), .A(n10552), .ZN(n10558) );
  XNOR2_X1 U11599 ( .A(P2_REG0_REG_25__SCAN_IN), .B(keyinput22), .ZN(n10556)
         );
  XNOR2_X1 U11600 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput46), .ZN(n10555) );
  NAND2_X1 U11601 ( .A1(n10556), .A2(n10555), .ZN(n10557) );
  NOR4_X1 U11602 ( .A1(n10560), .A2(n10559), .A3(n10558), .A4(n10557), .ZN(
        n10576) );
  AOI22_X1 U11603 ( .A1(n10562), .A2(keyinput121), .B1(keyinput33), .B2(n9912), 
        .ZN(n10561) );
  OAI221_X1 U11604 ( .B1(n10562), .B2(keyinput121), .C1(n9912), .C2(keyinput33), .A(n10561), .ZN(n10574) );
  AOI22_X1 U11605 ( .A1(n9687), .A2(keyinput49), .B1(keyinput48), .B2(n10564), 
        .ZN(n10563) );
  OAI221_X1 U11606 ( .B1(n9687), .B2(keyinput49), .C1(n10564), .C2(keyinput48), 
        .A(n10563), .ZN(n10573) );
  AOI22_X1 U11607 ( .A1(n10567), .A2(keyinput21), .B1(n10566), .B2(keyinput59), 
        .ZN(n10565) );
  OAI221_X1 U11608 ( .B1(n10567), .B2(keyinput21), .C1(n10566), .C2(keyinput59), .A(n10565), .ZN(n10572) );
  AOI22_X1 U11609 ( .A1(n10570), .A2(keyinput16), .B1(n10569), .B2(keyinput52), 
        .ZN(n10568) );
  OAI221_X1 U11610 ( .B1(n10570), .B2(keyinput16), .C1(n10569), .C2(keyinput52), .A(n10568), .ZN(n10571) );
  NOR4_X1 U11611 ( .A1(n10574), .A2(n10573), .A3(n10572), .A4(n10571), .ZN(
        n10575) );
  NAND4_X1 U11612 ( .A1(n10578), .A2(n10577), .A3(n10576), .A4(n10575), .ZN(
        n10579) );
  AOI211_X1 U11613 ( .C1(keyinput9), .C2(n10581), .A(n10580), .B(n10579), .ZN(
        n10582) );
  NAND4_X1 U11614 ( .A1(n10585), .A2(n10584), .A3(n10583), .A4(n10582), .ZN(
        n10590) );
  AOI22_X1 U11615 ( .A1(n10588), .A2(n10587), .B1(P1_REG0_REG_7__SCAN_IN), 
        .B2(n10586), .ZN(n10589) );
  XOR2_X1 U11616 ( .A(n10590), .B(n10589), .Z(P1_U3475) );
  XNOR2_X1 U11617 ( .A(n10592), .B(n10591), .ZN(ADD_1071_U50) );
  NOR2_X1 U11618 ( .A1(n10594), .A2(n10593), .ZN(n10595) );
  XOR2_X1 U11619 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10595), .Z(ADD_1071_U51) );
  OAI21_X1 U11620 ( .B1(n10598), .B2(n10597), .A(n10596), .ZN(n10599) );
  XNOR2_X1 U11621 ( .A(n10599), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11622 ( .B1(n10602), .B2(n10601), .A(n10600), .ZN(ADD_1071_U47) );
  XNOR2_X1 U11623 ( .A(n10604), .B(n10603), .ZN(ADD_1071_U48) );
  XNOR2_X1 U11624 ( .A(n10606), .B(n10605), .ZN(ADD_1071_U49) );
  XOR2_X1 U11625 ( .A(n10608), .B(n10607), .Z(ADD_1071_U54) );
  XOR2_X1 U11626 ( .A(n10609), .B(n10610), .Z(ADD_1071_U53) );
  XNOR2_X1 U11627 ( .A(n10612), .B(n10611), .ZN(ADD_1071_U52) );
  CLKBUF_X1 U4925 ( .A(n5263), .Z(n6463) );
  NAND2_X1 U4927 ( .A1(n6184), .A2(n6183), .ZN(n9545) );
  CLKBUF_X1 U4972 ( .A(n7261), .Z(n9122) );
  AND2_X1 U4973 ( .A1(n5291), .A2(P1_U3084), .ZN(n10615) );
endmodule

