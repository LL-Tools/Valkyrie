

module b15_C_AntiSAT_k_128_1 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2996, n2997, n2999, n3000, n3001, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3034, n3035, n3036, n3037, n3038,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788;

  INV_X1 U3443 ( .A(n6294), .ZN(n6276) );
  NOR2_X1 U3444 ( .A1(n5516), .A2(n3704), .ZN(n3060) );
  NAND2_X1 U34450 ( .A1(n3998), .A2(n3997), .ZN(n5295) );
  AOI21_X1 U34460 ( .B1(n3815), .B2(n3817), .A(n4723), .ZN(n4384) );
  AND2_X1 U34470 ( .A1(n3424), .A2(n4408), .ZN(n4448) );
  AND2_X1 U34480 ( .A1(n4442), .A2(n3421), .ZN(n4410) );
  CLKBUF_X1 U3450 ( .A(n3034), .Z(n4127) );
  CLKBUF_X2 U34510 ( .A(n3026), .Z(n3038) );
  CLKBUF_X1 U34520 ( .A(n3311), .Z(n3312) );
  OAI21_X1 U34530 ( .B1(n3221), .B2(n3219), .A(n3220), .ZN(n4344) );
  INV_X1 U34550 ( .A(n3606), .ZN(n4528) );
  AND2_X2 U34560 ( .A1(n3216), .A2(n3606), .ZN(n5139) );
  INV_X1 U3457 ( .A(n3251), .ZN(n3075) );
  AND4_X1 U3458 ( .A1(n3128), .A2(n3127), .A3(n3126), .A4(n3125), .ZN(n3129)
         );
  AND2_X2 U34600 ( .A1(n4357), .A2(n4585), .ZN(n4222) );
  AND2_X2 U34610 ( .A1(n4578), .A2(n4351), .ZN(n3032) );
  AND2_X2 U34620 ( .A1(n3113), .A2(n4585), .ZN(n3037) );
  AND2_X1 U34630 ( .A1(n4573), .A2(n4352), .ZN(n3313) );
  NAND2_X1 U34650 ( .A1(n3818), .A2(n6479), .ZN(n3409) );
  AND4_X1 U3466 ( .A1(n3156), .A2(n3155), .A3(n3154), .A4(n3153), .ZN(n3157)
         );
  AND2_X1 U3467 ( .A1(n3219), .A2(n3546), .ZN(n3566) );
  NAND2_X1 U34680 ( .A1(n3355), .A2(n3354), .ZN(n4589) );
  NAND2_X2 U34690 ( .A1(n3158), .A2(n3157), .ZN(n3219) );
  NAND2_X1 U34700 ( .A1(n3611), .A2(n3610), .ZN(n3613) );
  NAND2_X1 U34720 ( .A1(n3410), .A2(n3411), .ZN(n3415) );
  INV_X1 U34730 ( .A(n3001), .ZN(n4773) );
  INV_X1 U34740 ( .A(n6151), .ZN(n6143) );
  INV_X1 U3475 ( .A(n6161), .ZN(n6180) );
  OR2_X2 U3476 ( .A1(n5531), .A2(n5514), .ZN(n5516) );
  INV_X1 U3477 ( .A(n6303), .ZN(n6287) );
  AOI21_X1 U3478 ( .B1(n5413), .B2(n5423), .A(n5412), .ZN(n5414) );
  AND2_X2 U3479 ( .A1(n4354), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4357)
         );
  NAND2_X1 U3480 ( .A1(n3415), .A2(n3414), .ZN(n3815) );
  AND2_X1 U3481 ( .A1(n3579), .A2(n3578), .ZN(n6481) );
  AOI211_X1 U3482 ( .C1(n5553), .C2(n6158), .A(n5469), .B(n5468), .ZN(n5470)
         );
  NOR3_X4 U3483 ( .A1(n5516), .A2(n3704), .A3(n3051), .ZN(n5418) );
  NAND2_X2 U3484 ( .A1(n5673), .A2(n3520), .ZN(n5660) );
  NAND2_X2 U3485 ( .A1(n5675), .A2(n5674), .ZN(n5673) );
  NAND2_X2 U3486 ( .A1(n3244), .A2(n3243), .ZN(n3580) );
  AOI211_X2 U3487 ( .C1(n5933), .C2(REIP_REG_24__SCAN_IN), .A(n5925), .B(n5924), .ZN(n5926) );
  BUF_X4 U3489 ( .A(n3313), .Z(n2996) );
  INV_X2 U3490 ( .A(n3517), .ZN(n5718) );
  NOR2_X1 U3491 ( .A1(n5438), .A2(n5491), .ZN(n4282) );
  NAND2_X1 U3492 ( .A1(n5295), .A2(n3069), .ZN(n5593) );
  NAND2_X1 U3493 ( .A1(n3402), .A2(n3401), .ZN(n4804) );
  NAND2_X1 U3494 ( .A1(n3420), .A2(n3419), .ZN(n4463) );
  AOI211_X1 U3495 ( .C1(n4490), .C2(n6448), .A(n4583), .B(n4582), .ZN(n5867)
         );
  XNOR2_X1 U3496 ( .A(n3288), .B(n3287), .ZN(n3393) );
  NAND2_X1 U3497 ( .A1(n3260), .A2(n3259), .ZN(n3329) );
  OAI21_X1 U3498 ( .B1(n3240), .B2(n3224), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3226) );
  NOR2_X2 U3500 ( .A1(n3816), .A2(n3270), .ZN(n3234) );
  OR2_X1 U3501 ( .A1(n3213), .A2(n3212), .ZN(n3246) );
  INV_X2 U3502 ( .A(n3222), .ZN(n3242) );
  AND4_X1 U3503 ( .A1(n3124), .A2(n3123), .A3(n3122), .A4(n3121), .ZN(n3130)
         );
  BUF_X2 U3505 ( .A(n3276), .Z(n3035) );
  CLKBUF_X2 U3506 ( .A(n3292), .Z(n4244) );
  CLKBUF_X2 U3507 ( .A(n3203), .Z(n4246) );
  BUF_X2 U3509 ( .A(n3310), .Z(n4236) );
  AND2_X2 U3510 ( .A1(n4351), .A2(n4585), .ZN(n3367) );
  AND2_X1 U3512 ( .A1(n5675), .A2(n3049), .ZN(n5652) );
  OR2_X1 U3513 ( .A1(n5620), .A2(n6151), .ZN(n3053) );
  INV_X1 U3514 ( .A(n5472), .ZN(n5620) );
  AOI221_X1 U3515 ( .B1(REIP_REG_23__SCAN_IN), .B2(n5933), .C1(n5932), .C2(
        n5933), .A(n5931), .ZN(n5934) );
  XOR2_X1 U3516 ( .A(n5429), .B(n5428), .Z(n5472) );
  NAND2_X1 U3517 ( .A1(n4282), .A2(n4283), .ZN(n5428) );
  NAND2_X1 U3518 ( .A1(n5440), .A2(n5438), .ZN(n5627) );
  OAI21_X1 U3519 ( .B1(n5573), .B2(n5574), .A(n5564), .ZN(n5930) );
  AND2_X1 U3520 ( .A1(n3090), .A2(n3510), .ZN(n5729) );
  NAND2_X1 U3521 ( .A1(n3018), .A2(n3022), .ZN(n5564) );
  NOR2_X1 U3522 ( .A1(n5578), .A2(n5579), .ZN(n5573) );
  AND2_X1 U3523 ( .A1(n3011), .A2(n3012), .ZN(n5511) );
  AND2_X1 U3524 ( .A1(n4074), .A2(n4073), .ZN(n3018) );
  AND2_X1 U3525 ( .A1(n4074), .A2(n4073), .ZN(n3011) );
  INV_X1 U3526 ( .A(n5593), .ZN(n4074) );
  NAND2_X1 U3527 ( .A1(n3021), .A2(n3504), .ZN(n5197) );
  NAND2_X1 U3528 ( .A1(n5163), .A2(n5164), .ZN(n3021) );
  INV_X1 U3529 ( .A(n3088), .ZN(n3083) );
  NAND2_X1 U3530 ( .A1(n3087), .A2(n5736), .ZN(n3086) );
  AND2_X1 U3531 ( .A1(n3041), .A2(n5736), .ZN(n3088) );
  AND2_X1 U3532 ( .A1(n3495), .A2(n3019), .ZN(n3010) );
  NAND2_X1 U3533 ( .A1(n3047), .A2(n3513), .ZN(n3089) );
  AND2_X1 U3534 ( .A1(n3060), .A2(n3059), .ZN(n5495) );
  AND2_X1 U3535 ( .A1(n5393), .A2(n3509), .ZN(n3512) );
  NAND2_X1 U3536 ( .A1(n5727), .A2(n6000), .ZN(n3513) );
  OR2_X1 U3537 ( .A1(n3498), .A2(n3497), .ZN(n3508) );
  OR2_X1 U3538 ( .A1(n3498), .A2(n3497), .ZN(n3007) );
  AND3_X1 U3539 ( .A1(n3826), .A2(n4617), .A3(n4432), .ZN(n4650) );
  NAND2_X1 U3540 ( .A1(n3832), .A2(n3831), .ZN(n4652) );
  OAI21_X1 U3541 ( .B1(n3458), .B2(n3560), .A(n3457), .ZN(n3459) );
  NOR2_X1 U3542 ( .A1(n4616), .A2(n4457), .ZN(n4617) );
  XNOR2_X1 U3543 ( .A(n3486), .B(n3485), .ZN(n3840) );
  AOI21_X1 U3544 ( .B1(n3775), .B2(n3949), .A(n3783), .ZN(n4616) );
  AND2_X1 U3545 ( .A1(n3450), .A2(n3389), .ZN(n3775) );
  AND2_X1 U3546 ( .A1(n3067), .A2(n3066), .ZN(n3065) );
  OR2_X1 U3547 ( .A1(n4804), .A2(n3939), .ZN(n3814) );
  XNOR2_X1 U3548 ( .A(n3393), .B(n3392), .ZN(n3805) );
  NAND2_X1 U3549 ( .A1(n4463), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4462)
         );
  NAND2_X1 U3550 ( .A1(n3352), .A2(n3351), .ZN(n3402) );
  NAND2_X1 U3551 ( .A1(n3398), .A2(n3400), .ZN(n3351) );
  NAND2_X2 U3552 ( .A1(n3722), .A2(n3605), .ZN(n6307) );
  NOR2_X1 U3553 ( .A1(n3023), .A2(n5579), .ZN(n3022) );
  NAND2_X1 U3554 ( .A1(n3269), .A2(n3268), .ZN(n3354) );
  AND2_X1 U3555 ( .A1(n4413), .A2(n4412), .ZN(n4452) );
  OR2_X1 U3556 ( .A1(n4346), .A2(n3776), .ZN(n3706) );
  AND2_X1 U3557 ( .A1(n5596), .A2(n3751), .ZN(n3756) );
  INV_X1 U3558 ( .A(n5139), .ZN(n6591) );
  OR2_X1 U3559 ( .A1(n3159), .A2(n3234), .ZN(n3249) );
  INV_X2 U3560 ( .A(n5541), .ZN(n5596) );
  INV_X1 U3561 ( .A(n3246), .ZN(n4521) );
  AND2_X2 U3562 ( .A1(n3600), .A2(n3606), .ZN(n5134) );
  OR2_X1 U3563 ( .A1(n3302), .A2(n3301), .ZN(n3500) );
  NAND3_X2 U3564 ( .A1(n3180), .A2(n3179), .A3(n3178), .ZN(n3600) );
  INV_X2 U3565 ( .A(n3106), .ZN(n2997) );
  AND2_X1 U3566 ( .A1(n3606), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3546) );
  OR2_X1 U3567 ( .A1(n3319), .A2(n3318), .ZN(n3417) );
  AND2_X2 U3568 ( .A1(n3120), .A2(n3119), .ZN(n3222) );
  AND4_X1 U3569 ( .A1(n3173), .A2(n3172), .A3(n3171), .A4(n3170), .ZN(n3179)
         );
  NAND2_X2 U3570 ( .A1(n3130), .A2(n3129), .ZN(n3251) );
  AND2_X1 U3571 ( .A1(n3169), .A2(n3168), .ZN(n3180) );
  AND4_X1 U3572 ( .A1(n3163), .A2(n3162), .A3(n3161), .A4(n3160), .ZN(n3169)
         );
  AND4_X1 U3573 ( .A1(n3112), .A2(n3111), .A3(n3110), .A4(n3109), .ZN(n3120)
         );
  AND4_X1 U3574 ( .A1(n3189), .A2(n3188), .A3(n3187), .A4(n3186), .ZN(n3200)
         );
  AND4_X1 U3575 ( .A1(n3185), .A2(n3184), .A3(n3183), .A4(n3182), .ZN(n3201)
         );
  AND4_X1 U3576 ( .A1(n3152), .A2(n3151), .A3(n3150), .A4(n3149), .ZN(n3158)
         );
  AND4_X1 U3577 ( .A1(n3116), .A2(n3117), .A3(n3118), .A4(n3115), .ZN(n3119)
         );
  AND4_X1 U3578 ( .A1(n3193), .A2(n3192), .A3(n3191), .A4(n3190), .ZN(n3199)
         );
  AND4_X1 U3579 ( .A1(n3197), .A2(n3196), .A3(n3195), .A4(n3194), .ZN(n3198)
         );
  AND4_X1 U3580 ( .A1(n3167), .A2(n3166), .A3(n3165), .A4(n3164), .ZN(n3168)
         );
  AND4_X1 U3581 ( .A1(n3177), .A2(n3176), .A3(n3175), .A4(n3174), .ZN(n3178)
         );
  BUF_X2 U3582 ( .A(n3275), .Z(n4247) );
  NAND2_X2 U3583 ( .A1(n4268), .A2(n6350), .ZN(n6303) );
  AND2_X2 U3584 ( .A1(n3114), .A2(n4357), .ZN(n3292) );
  INV_X2 U3585 ( .A(n6559), .ZN(n6597) );
  AND2_X2 U3586 ( .A1(n4573), .A2(n4351), .ZN(n4183) );
  AND2_X2 U3587 ( .A1(n4573), .A2(n4351), .ZN(n3028) );
  NOR2_X1 U3588 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4596), .ZN(n6239) );
  INV_X2 U3589 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6479) );
  OR2_X1 U3590 ( .A1(n3594), .A2(n3600), .ZN(n2999) );
  OR2_X1 U3591 ( .A1(n3594), .A2(n3600), .ZN(n3602) );
  NOR2_X2 U3592 ( .A1(n5320), .A2(n5321), .ZN(n5378) );
  NOR2_X2 U3593 ( .A1(n5223), .A2(n5224), .ZN(n3062) );
  XNOR2_X2 U3594 ( .A(n3761), .B(n3760), .ZN(n5553) );
  NAND2_X2 U3595 ( .A1(n3222), .A2(n3251), .ZN(n4376) );
  BUF_X1 U3596 ( .A(n5717), .Z(n3000) );
  NAND2_X1 U3597 ( .A1(n3427), .A2(n3794), .ZN(n3001) );
  NAND2_X1 U3598 ( .A1(n3427), .A2(n3794), .ZN(n3784) );
  AND2_X2 U3599 ( .A1(n4578), .A2(n4352), .ZN(n3275) );
  INV_X1 U3600 ( .A(n3794), .ZN(n3064) );
  NAND2_X1 U3601 ( .A1(n5151), .A2(n5152), .ZN(n3003) );
  AND2_X1 U3602 ( .A1(n5439), .A2(n3012), .ZN(n3004) );
  OR2_X1 U3603 ( .A1(n5190), .A2(n5119), .ZN(n3005) );
  OR2_X1 U3604 ( .A1(n4921), .A2(n5119), .ZN(n5116) );
  NAND2_X1 U3605 ( .A1(n3019), .A2(n3006), .ZN(n3009) );
  NAND2_X1 U3606 ( .A1(n5164), .A2(n3098), .ZN(n3006) );
  NAND2_X1 U3607 ( .A1(n3486), .A2(n3548), .ZN(n3498) );
  NOR3_X2 U3608 ( .A1(n5310), .A2(n3055), .A3(n5586), .ZN(n3057) );
  OR2_X2 U3609 ( .A1(n3020), .A2(n3504), .ZN(n3019) );
  AOI21_X1 U3610 ( .B1(n3098), .B2(n3505), .A(n3096), .ZN(n3095) );
  AND2_X2 U3611 ( .A1(n4357), .A2(n4578), .ZN(n3276) );
  NAND2_X1 U3612 ( .A1(n3496), .A2(n3010), .ZN(n3008) );
  NAND2_X1 U3613 ( .A1(n3008), .A2(n3009), .ZN(n3097) );
  AND2_X1 U3614 ( .A1(n3065), .A2(n3022), .ZN(n3012) );
  CLKBUF_X1 U3615 ( .A(n5273), .Z(n3013) );
  NAND2_X1 U3616 ( .A1(n3097), .A2(n3017), .ZN(n3014) );
  AND2_X2 U3617 ( .A1(n3014), .A2(n3015), .ZN(n5273) );
  OR2_X1 U3618 ( .A1(n3016), .A2(n5255), .ZN(n3015) );
  INV_X1 U3619 ( .A(n5256), .ZN(n3016) );
  AND2_X1 U3620 ( .A1(n3095), .A2(n5256), .ZN(n3017) );
  INV_X1 U3621 ( .A(n3098), .ZN(n3020) );
  INV_X1 U3622 ( .A(n5574), .ZN(n3023) );
  NOR2_X1 U3623 ( .A1(n5428), .A2(n5429), .ZN(n4267) );
  CLKBUF_X1 U3624 ( .A(n4906), .Z(n3024) );
  AND2_X4 U3625 ( .A1(n3107), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4578)
         );
  BUF_X2 U3626 ( .A(n3304), .Z(n3025) );
  AND2_X1 U3628 ( .A1(n4573), .A2(n4351), .ZN(n3027) );
  AND2_X1 U3629 ( .A1(n3113), .A2(n4578), .ZN(n3304) );
  AND2_X1 U3630 ( .A1(n4357), .A2(n4585), .ZN(n3029) );
  AND2_X2 U3631 ( .A1(n4357), .A2(n4585), .ZN(n3030) );
  NAND2_X2 U3632 ( .A1(n5706), .A2(n5705), .ZN(n5704) );
  AOI22_X2 U3633 ( .A1(n5711), .A2(n5712), .B1(n3506), .B2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5706) );
  NAND2_X2 U3634 ( .A1(n3064), .A2(n3040), .ZN(n3791) );
  AND2_X2 U3635 ( .A1(n3747), .A2(n3052), .ZN(n5412) );
  NOR2_X4 U3636 ( .A1(n5660), .A2(n5661), .ZN(n3747) );
  OAI21_X2 U3637 ( .B1(n3506), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5704), 
        .ZN(n5700) );
  AND2_X4 U3638 ( .A1(n4352), .A2(n4585), .ZN(n3277) );
  AND2_X4 U3639 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4585) );
  OR2_X2 U3640 ( .A1(n3580), .A2(n4528), .ZN(n4288) );
  INV_X1 U3641 ( .A(n3007), .ZN(n3031) );
  NAND2_X2 U3642 ( .A1(n3425), .A2(n4488), .ZN(n3794) );
  OR2_X1 U3643 ( .A1(n3815), .A2(n3560), .ZN(n3420) );
  AND2_X2 U3644 ( .A1(n4376), .A2(n3270), .ZN(n3045) );
  INV_X2 U3645 ( .A(n3219), .ZN(n3270) );
  BUF_X4 U3646 ( .A(n3276), .Z(n3034) );
  AND2_X4 U3647 ( .A1(n3114), .A2(n4351), .ZN(n3331) );
  AND2_X4 U3648 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4351) );
  NAND2_X2 U3649 ( .A1(n5975), .A2(n5974), .ZN(n5392) );
  OAI21_X2 U3650 ( .B1(n5273), .B2(n5271), .A(n5269), .ZN(n5975) );
  OAI21_X1 U3651 ( .B1(n3784), .B2(n3560), .A(n3430), .ZN(n3432) );
  AOI211_X2 U3652 ( .C1(n5797), .C2(n6322), .A(n5796), .B(n5795), .ZN(n5798)
         );
  XNOR2_X2 U3653 ( .A(n5686), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5797)
         );
  NOR2_X2 U3654 ( .A1(n3005), .A2(n4921), .ZN(n5191) );
  OAI21_X2 U3655 ( .B1(n3990), .B2(n3994), .A(n5312), .ZN(n5265) );
  AND2_X4 U3656 ( .A1(n3113), .A2(n4585), .ZN(n4245) );
  AND2_X1 U3657 ( .A1(n3387), .A2(n3386), .ZN(n3792) );
  OR2_X1 U3658 ( .A1(n3342), .A2(n3341), .ZN(n3404) );
  INV_X1 U3659 ( .A(n3474), .ZN(n3475) );
  INV_X1 U3660 ( .A(n3791), .ZN(n3476) );
  NAND2_X1 U3661 ( .A1(n3791), .A2(n3474), .ZN(n3827) );
  INV_X1 U3662 ( .A(n3548), .ZN(n3560) );
  OAI21_X1 U3663 ( .B1(n5392), .B2(n3084), .A(n3082), .ZN(n5679) );
  INV_X1 U3664 ( .A(n3086), .ZN(n3084) );
  AOI21_X1 U3665 ( .B1(n3083), .B2(n3086), .A(n3046), .ZN(n3082) );
  NAND2_X1 U3666 ( .A1(n3362), .A2(n3361), .ZN(n3572) );
  AND2_X1 U3667 ( .A1(n3242), .A2(n3600), .ZN(n3548) );
  AND2_X1 U3668 ( .A1(n3473), .A2(n3472), .ZN(n3474) );
  OR2_X1 U3669 ( .A1(n3447), .A2(n3446), .ZN(n3455) );
  INV_X1 U3670 ( .A(n3285), .ZN(n3394) );
  NAND3_X1 U3671 ( .A1(n3254), .A2(n3256), .A3(n3255), .ZN(n3260) );
  NAND2_X1 U3672 ( .A1(n3328), .A2(n3497), .ZN(n3350) );
  OR2_X1 U3673 ( .A1(n3362), .A2(n3344), .ZN(n3343) );
  AND2_X1 U3674 ( .A1(n4051), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4052)
         );
  OR2_X1 U3675 ( .A1(n5445), .A2(n4723), .ZN(n3106) );
  INV_X1 U3676 ( .A(n3048), .ZN(n3063) );
  AND2_X1 U3677 ( .A1(n5737), .A2(n3514), .ZN(n3515) );
  NOR2_X1 U3678 ( .A1(n5210), .A2(n3099), .ZN(n3098) );
  INV_X1 U3679 ( .A(n3507), .ZN(n3099) );
  INV_X1 U3680 ( .A(n3750), .ZN(n3757) );
  OR2_X1 U3681 ( .A1(n3327), .A2(n6479), .ZN(n3497) );
  NAND2_X1 U3682 ( .A1(n5596), .A2(n5134), .ZN(n3702) );
  NAND2_X1 U3683 ( .A1(n4514), .A2(n3246), .ZN(n3710) );
  NAND2_X1 U3684 ( .A1(n3241), .A2(n3713), .ZN(n3289) );
  AND4_X1 U3685 ( .A1(n3230), .A2(n3239), .A3(n4579), .A4(n3238), .ZN(n3241)
         );
  INV_X1 U3686 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6453) );
  INV_X1 U3687 ( .A(n5180), .ZN(n5175) );
  INV_X1 U3688 ( .A(n4122), .ZN(n4265) );
  OR2_X1 U3689 ( .A1(n4262), .A2(n5484), .ZN(n4273) );
  NAND2_X1 U3690 ( .A1(n4196), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4262)
         );
  INV_X1 U3691 ( .A(n5565), .ZN(n3066) );
  NOR2_X1 U3692 ( .A1(n5512), .A2(n3068), .ZN(n3067) );
  NAND2_X1 U3693 ( .A1(n5525), .A2(n5527), .ZN(n5526) );
  AND2_X1 U3694 ( .A1(n4120), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4157)
         );
  NAND2_X1 U3695 ( .A1(n3994), .A2(n3990), .ZN(n5312) );
  INV_X1 U3696 ( .A(n5662), .ZN(n3093) );
  NOR2_X1 U3697 ( .A1(n5300), .A2(n3058), .ZN(n3056) );
  NAND2_X1 U3698 ( .A1(n5392), .A2(n3088), .ZN(n3081) );
  NAND2_X1 U3699 ( .A1(n5392), .A2(n3041), .ZN(n3085) );
  OR2_X1 U3700 ( .A1(n5379), .A2(n5308), .ZN(n5310) );
  NAND2_X1 U3701 ( .A1(n5378), .A2(n5377), .ZN(n5379) );
  OR2_X1 U3702 ( .A1(n5197), .A2(n3505), .ZN(n3100) );
  NOR2_X2 U3703 ( .A1(n5054), .A2(n4924), .ZN(n5137) );
  INV_X1 U3704 ( .A(n3374), .ZN(n3375) );
  AND2_X1 U3705 ( .A1(n5325), .A2(n6350), .ZN(n5332) );
  AND2_X1 U3706 ( .A1(n4761), .A2(n4490), .ZN(n5329) );
  AND2_X1 U3707 ( .A1(n3532), .A2(n3539), .ZN(n3575) );
  OR2_X1 U3708 ( .A1(n3540), .A2(n3531), .ZN(n3532) );
  NAND2_X1 U3709 ( .A1(n3566), .A2(n3548), .ZN(n3577) );
  AND2_X2 U3710 ( .A1(n4382), .A2(n4424), .ZN(n6195) );
  AND2_X1 U3711 ( .A1(n5613), .A2(n5444), .ZN(n6202) );
  AND2_X1 U3712 ( .A1(n5613), .A2(n5446), .ZN(n6206) );
  INV_X1 U3713 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6357) );
  NOR2_X1 U3714 ( .A1(n6567), .A2(n6481), .ZN(n5400) );
  INV_X1 U3715 ( .A(n3792), .ZN(n3388) );
  OR2_X1 U3716 ( .A1(n3385), .A2(n3384), .ZN(n3452) );
  INV_X1 U3717 ( .A(n4514), .ZN(n3708) );
  AND2_X2 U3718 ( .A1(n3076), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3113)
         );
  AOI22_X1 U3719 ( .A1(n3203), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3125) );
  NAND2_X1 U3720 ( .A1(n3270), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3362) );
  NAND2_X1 U3721 ( .A1(n4528), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3361) );
  AOI22_X1 U3722 ( .A1(n4239), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3146) );
  NAND2_X1 U3723 ( .A1(n4222), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3193)
         );
  NAND2_X1 U3724 ( .A1(n4140), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3190) );
  INV_X1 U3725 ( .A(n5527), .ZN(n3068) );
  AND2_X1 U3726 ( .A1(n3071), .A2(n4021), .ZN(n3070) );
  INV_X1 U3727 ( .A(n5545), .ZN(n3071) );
  NOR2_X1 U3728 ( .A1(n4013), .A2(n6063), .ZN(n4014) );
  NAND2_X1 U3729 ( .A1(n3064), .A2(n3388), .ZN(n3450) );
  NAND2_X1 U3730 ( .A1(n3075), .A2(n5445), .ZN(n3816) );
  INV_X1 U3731 ( .A(n5492), .ZN(n3059) );
  INV_X1 U3732 ( .A(n3089), .ZN(n3087) );
  NAND2_X1 U3733 ( .A1(n3840), .A2(n3548), .ZN(n3492) );
  OAI21_X1 U3734 ( .B1(n3479), .B2(n3498), .A(n3478), .ZN(n3480) );
  NAND2_X1 U3735 ( .A1(n3397), .A2(n3396), .ZN(n3422) );
  AOI22_X1 U3736 ( .A1(n4183), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3153) );
  AOI22_X1 U3737 ( .A1(n3030), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3154) );
  OR2_X1 U3738 ( .A1(n3373), .A2(n3372), .ZN(n3429) );
  AND2_X1 U3739 ( .A1(n3270), .A2(n3242), .ZN(n4343) );
  NAND2_X1 U3740 ( .A1(n3566), .A2(n4429), .ZN(n3225) );
  INV_X1 U3741 ( .A(n3600), .ZN(n3216) );
  AOI22_X1 U3742 ( .A1(n3026), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3117) );
  AOI21_X1 U3743 ( .B1(n5121), .B2(n4596), .A(n5400), .ZN(n4494) );
  INV_X1 U3744 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6458) );
  INV_X1 U3745 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n5235) );
  NAND2_X1 U3746 ( .A1(n5569), .A2(n5529), .ZN(n5531) );
  NAND2_X1 U3747 ( .A1(n3682), .A2(n3056), .ZN(n3055) );
  AND2_X1 U3748 ( .A1(n3663), .A2(n3662), .ZN(n5321) );
  AND2_X1 U3749 ( .A1(n3653), .A2(n3652), .ZN(n5194) );
  AND2_X1 U3750 ( .A1(n4362), .A2(n3721), .ZN(n4375) );
  OR2_X1 U3751 ( .A1(n3824), .A2(n3823), .ZN(n4435) );
  AND2_X1 U3752 ( .A1(n4388), .A2(n4387), .ZN(n6209) );
  AND2_X1 U3753 ( .A1(n4195), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4196)
         );
  AND2_X1 U3754 ( .A1(n4157), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4158)
         );
  NAND2_X1 U3755 ( .A1(n4158), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4194)
         );
  NOR2_X1 U3756 ( .A1(n4119), .A2(n5936), .ZN(n4120) );
  AOI211_X1 U3757 ( .C1(n2997), .C2(EAX_REG_24__SCAN_IN), .A(n4138), .B(n4137), 
        .ZN(n5565) );
  INV_X1 U3758 ( .A(n4075), .ZN(n4076) );
  NAND2_X1 U3759 ( .A1(n4077), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4119)
         );
  NAND2_X1 U3760 ( .A1(n4052), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4075)
         );
  INV_X1 U3761 ( .A(n5584), .ZN(n4073) );
  AND2_X1 U3762 ( .A1(n5590), .A2(n3070), .ZN(n3069) );
  AND2_X1 U3763 ( .A1(n5295), .A2(n3070), .ZN(n5591) );
  AND2_X1 U3764 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n4014), .ZN(n4051)
         );
  NAND2_X1 U3765 ( .A1(n5295), .A2(n4021), .ZN(n5604) );
  NAND2_X1 U3766 ( .A1(n3973), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4013)
         );
  INV_X1 U3767 ( .A(n5295), .ZN(n5602) );
  AND2_X1 U3768 ( .A1(n3956), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3973)
         );
  NAND2_X1 U3769 ( .A1(n5392), .A2(n3512), .ZN(n3090) );
  NOR2_X1 U3770 ( .A1(n6757), .A2(n3936), .ZN(n3956) );
  AND2_X1 U3771 ( .A1(n3899), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3772)
         );
  NAND2_X1 U3772 ( .A1(n3869), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3884)
         );
  INV_X1 U3773 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3885) );
  NOR2_X1 U3774 ( .A1(n3856), .A2(n6114), .ZN(n3869) );
  NAND2_X1 U3775 ( .A1(n3852), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3856)
         );
  CLKBUF_X1 U3776 ( .A(n4921), .Z(n5118) );
  AND3_X1 U3777 ( .A1(n3855), .A2(n3854), .A3(n3853), .ZN(n5047) );
  AOI21_X1 U3778 ( .B1(n3840), .B2(n3949), .A(n3839), .ZN(n5002) );
  NAND2_X1 U3779 ( .A1(n3827), .A2(n3949), .ZN(n3832) );
  NOR2_X1 U3780 ( .A1(n3797), .A2(n6283), .ZN(n3828) );
  AOI21_X1 U3781 ( .B1(n3791), .B2(n3804), .A(n3803), .ZN(n4847) );
  INV_X1 U3782 ( .A(n3802), .ZN(n3803) );
  NAND2_X1 U3783 ( .A1(n3785), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3797)
         );
  NOR2_X1 U3784 ( .A1(n3807), .A2(n5235), .ZN(n3785) );
  NAND2_X1 U3785 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3807) );
  OAI21_X1 U3786 ( .B1(n4804), .B2(n3560), .A(n3408), .ZN(n4440) );
  NOR2_X1 U3787 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3079) );
  NAND2_X1 U3788 ( .A1(n3759), .A2(n3758), .ZN(n5449) );
  INV_X1 U3789 ( .A(n5418), .ZN(n5416) );
  INV_X1 U3790 ( .A(n3060), .ZN(n5493) );
  NAND2_X1 U3791 ( .A1(n3518), .A2(n5727), .ZN(n3092) );
  NOR2_X1 U3792 ( .A1(n3519), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3094)
         );
  NOR2_X1 U3793 ( .A1(n5310), .A2(n5300), .ZN(n5607) );
  NAND2_X1 U3794 ( .A1(n3062), .A2(n3061), .ZN(n5320) );
  NAND2_X1 U3795 ( .A1(n5195), .A2(n5194), .ZN(n5224) );
  INV_X1 U3796 ( .A(n5211), .ZN(n3096) );
  OR2_X1 U3797 ( .A1(n6575), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4269) );
  AND2_X1 U3798 ( .A1(n3645), .A2(n3644), .ZN(n5051) );
  AND2_X1 U3799 ( .A1(n3640), .A2(n3639), .ZN(n5004) );
  NAND2_X1 U3800 ( .A1(n3633), .A2(n3632), .ZN(n4914) );
  INV_X1 U3801 ( .A(n4911), .ZN(n3632) );
  INV_X1 U3802 ( .A(n4912), .ZN(n3633) );
  AND2_X1 U3803 ( .A1(n3626), .A2(n3625), .ZN(n4609) );
  NAND2_X1 U3804 ( .A1(n3628), .A2(n3627), .ZN(n4912) );
  INV_X1 U3805 ( .A(n4609), .ZN(n3627) );
  NOR2_X1 U3806 ( .A1(n3710), .A2(n3242), .ZN(n3243) );
  INV_X1 U3807 ( .A(n5134), .ZN(n4379) );
  INV_X1 U3808 ( .A(n3756), .ZN(n4374) );
  AND2_X1 U3809 ( .A1(n3599), .A2(n4424), .ZN(n3722) );
  CLKBUF_X1 U3810 ( .A(n4491), .Z(n5183) );
  INV_X1 U3811 ( .A(n3289), .ZN(n3290) );
  INV_X1 U3812 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4354) );
  AND2_X1 U3813 ( .A1(n4805), .A2(n4804), .ZN(n4811) );
  OR2_X1 U3814 ( .A1(n4490), .A2(n4966), .ZN(n6349) );
  AND2_X1 U3815 ( .A1(n5860), .A2(n4601), .ZN(n4805) );
  OR2_X1 U3816 ( .A1(n6565), .A2(n4494), .ZN(n4549) );
  AND2_X1 U3817 ( .A1(n5860), .A2(n4602), .ZN(n4635) );
  NOR2_X1 U3818 ( .A1(n4804), .A2(n4810), .ZN(n4674) );
  INV_X1 U3819 ( .A(n6177), .ZN(n6160) );
  NAND2_X1 U3820 ( .A1(n5175), .A2(n5128), .ZN(n6185) );
  INV_X1 U3821 ( .A(n5547), .ZN(n6138) );
  AND2_X1 U3822 ( .A1(n5176), .A2(n6151), .ZN(n6157) );
  INV_X1 U3823 ( .A(n6172), .ZN(n6169) );
  INV_X1 U3824 ( .A(n5608), .ZN(n6191) );
  INV_X1 U3825 ( .A(n5288), .ZN(n5233) );
  NAND2_X1 U3826 ( .A1(n4428), .A2(n4427), .ZN(n5613) );
  BUF_X1 U3828 ( .A(n6238), .Z(n6229) );
  INV_X1 U3829 ( .A(n4428), .ZN(n6260) );
  OR2_X1 U3830 ( .A1(n4273), .A2(n5432), .ZN(n4275) );
  NAND2_X1 U3831 ( .A1(n5428), .A2(n4284), .ZN(n5443) );
  OR2_X1 U3832 ( .A1(n4282), .A2(n4283), .ZN(n4284) );
  OR2_X1 U3833 ( .A1(n5511), .A2(n5439), .ZN(n5440) );
  AND2_X1 U3834 ( .A1(n5313), .A2(n5267), .ZN(n6100) );
  INV_X1 U3835 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U3836 ( .A1(n6282), .A2(n6299), .ZN(n6294) );
  INV_X1 U3837 ( .A(n6282), .ZN(n6300) );
  XNOR2_X1 U3838 ( .A(n3077), .B(n4356), .ZN(n3771) );
  NAND2_X1 U3839 ( .A1(n3080), .A2(n3078), .ZN(n3077) );
  NAND2_X1 U3840 ( .A1(n5413), .A2(n3079), .ZN(n3078) );
  NAND2_X1 U3841 ( .A1(n5412), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3080) );
  AND2_X1 U3842 ( .A1(n5787), .A2(n3742), .ZN(n5763) );
  AND2_X1 U3843 ( .A1(n5841), .A2(n3741), .ZN(n5787) );
  AND2_X1 U3844 ( .A1(n5799), .A2(n3729), .ZN(n5791) );
  NOR2_X1 U3845 ( .A1(n5310), .A2(n3054), .ZN(n5594) );
  INV_X1 U3846 ( .A(n3056), .ZN(n3054) );
  NAND2_X1 U3847 ( .A1(n3085), .A2(n3089), .ZN(n5739) );
  NAND2_X1 U3848 ( .A1(n3100), .A2(n3507), .ZN(n5214) );
  OR2_X1 U3849 ( .A1(n5150), .A2(n5149), .ZN(n6312) );
  INV_X1 U3850 ( .A(n6333), .ZN(n6309) );
  INV_X1 U3851 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n4930) );
  CLKBUF_X1 U3852 ( .A(n4341), .Z(n4342) );
  INV_X1 U3853 ( .A(n4804), .ZN(n5856) );
  CLKBUF_X1 U3854 ( .A(n3805), .Z(n5860) );
  INV_X1 U3855 ( .A(n4490), .ZN(n5877) );
  INV_X1 U3856 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6738) );
  NOR2_X1 U3857 ( .A1(n4496), .A2(n3815), .ZN(n4751) );
  AOI22_X1 U3858 ( .A1(n5332), .A2(n5329), .B1(n6344), .B2(n5327), .ZN(n5371)
         );
  OR2_X1 U3859 ( .A1(n3577), .A2(n3576), .ZN(n3578) );
  OAI21_X1 U3860 ( .B1(n5627), .B2(n6303), .A(n3072), .ZN(U2959) );
  INV_X1 U3861 ( .A(n3073), .ZN(n3072) );
  OAI21_X1 U3862 ( .B1(n5442), .B2(n6297), .A(n3074), .ZN(n3073) );
  AOI21_X1 U3863 ( .B1(n6276), .B2(n5504), .A(n5441), .ZN(n3074) );
  CLKBUF_X3 U3864 ( .A(n4140), .Z(n4237) );
  INV_X1 U3865 ( .A(n3510), .ZN(n3511) );
  AND2_X1 U3866 ( .A1(n3388), .A2(n3063), .ZN(n3040) );
  NAND2_X1 U3867 ( .A1(n4650), .A2(n4652), .ZN(n4651) );
  INV_X1 U3868 ( .A(n5445), .ZN(n5612) );
  NOR2_X1 U3869 ( .A1(n5564), .A2(n5565), .ZN(n5525) );
  NAND2_X1 U3870 ( .A1(n3081), .A2(n3086), .ZN(n5726) );
  AND2_X1 U3871 ( .A1(n3512), .A2(n3513), .ZN(n3041) );
  INV_X2 U3872 ( .A(n3007), .ZN(n3506) );
  AND3_X1 U3873 ( .A1(n3137), .A2(n3136), .A3(n3135), .ZN(n3042) );
  OR2_X1 U3874 ( .A1(n5443), .A2(n6303), .ZN(n3043) );
  AND2_X1 U3875 ( .A1(n3218), .A2(n3217), .ZN(n3230) );
  AND2_X1 U3876 ( .A1(n3506), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3044)
         );
  AND2_X1 U3877 ( .A1(n5727), .A2(n3740), .ZN(n3046) );
  OR2_X1 U3878 ( .A1(n3511), .A2(n3044), .ZN(n3047) );
  NAND2_X1 U3879 ( .A1(n3097), .A2(n3095), .ZN(n5257) );
  AND2_X1 U3880 ( .A1(n3449), .A2(n3448), .ZN(n3048) );
  AND2_X1 U3881 ( .A1(n5674), .A2(n3093), .ZN(n3049) );
  OR2_X1 U3882 ( .A1(n5310), .A2(n3055), .ZN(n3050) );
  INV_X1 U3883 ( .A(n6307), .ZN(n6322) );
  INV_X1 U3884 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3107) );
  NAND2_X1 U3885 ( .A1(n4385), .A2(n3770), .ZN(n6297) );
  INV_X1 U3886 ( .A(n6297), .ZN(n6289) );
  AND2_X1 U3887 ( .A1(n3825), .A2(n4435), .ZN(n4432) );
  INV_X1 U3888 ( .A(n3062), .ZN(n5291) );
  INV_X1 U3889 ( .A(n5292), .ZN(n3061) );
  NAND2_X1 U3890 ( .A1(n4452), .A2(n3621), .ZN(n4610) );
  INV_X1 U3891 ( .A(n4610), .ZN(n3628) );
  NAND2_X1 U3892 ( .A1(n3059), .A2(n5451), .ZN(n3051) );
  AND2_X1 U3893 ( .A1(n3746), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3052)
         );
  AOI21_X2 U3894 ( .B1(n5250), .B2(n5134), .A(n3614), .ZN(n4413) );
  NAND2_X1 U3895 ( .A1(n5479), .A2(n3053), .ZN(U2797) );
  INV_X1 U3896 ( .A(n3057), .ZN(n5588) );
  INV_X1 U3897 ( .A(n5544), .ZN(n3058) );
  NAND3_X1 U3898 ( .A1(n4650), .A2(n4652), .A3(n3841), .ZN(n5000) );
  NAND2_X1 U3899 ( .A1(n3242), .A2(n3075), .ZN(n3221) );
  NOR2_X1 U3900 ( .A1(n4549), .A2(n3075), .ZN(n6409) );
  INV_X1 U3901 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3076) );
  AND2_X2 U3902 ( .A1(n4573), .A2(n3113), .ZN(n3203) );
  NOR2_X4 U3903 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4573) );
  NAND2_X1 U3904 ( .A1(n5718), .A2(n3094), .ZN(n3091) );
  NAND2_X1 U3905 ( .A1(n3092), .A2(n3091), .ZN(n5675) );
  NAND2_X1 U3906 ( .A1(n5718), .A2(n3516), .ZN(n5717) );
  NAND2_X1 U3907 ( .A1(n3101), .A2(n3391), .ZN(n3435) );
  NAND3_X1 U3908 ( .A1(n3450), .A2(n3548), .A3(n3389), .ZN(n3101) );
  INV_X1 U3909 ( .A(n3422), .ZN(n3423) );
  NAND2_X1 U3910 ( .A1(n5679), .A2(n3515), .ZN(n3517) );
  NAND2_X1 U3911 ( .A1(n3004), .A2(n3011), .ZN(n5438) );
  NOR2_X1 U3912 ( .A1(n3247), .A2(n3104), .ZN(n3248) );
  NAND2_X1 U3913 ( .A1(n3476), .A2(n3475), .ZN(n3486) );
  INV_X1 U3914 ( .A(n4847), .ZN(n3826) );
  NOR2_X1 U3915 ( .A1(n6344), .A2(n4719), .ZN(n3102) );
  OR2_X1 U3916 ( .A1(n3743), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n3103)
         );
  OR2_X1 U3917 ( .A1(n3246), .A2(n3606), .ZN(n3104) );
  AND2_X1 U3918 ( .A1(n5613), .A2(n4430), .ZN(n6203) );
  AND4_X1 U3919 ( .A1(n3134), .A2(n3133), .A3(n3132), .A4(n3131), .ZN(n3105)
         );
  INV_X1 U3920 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6114) );
  INV_X1 U3921 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6757) );
  INV_X1 U3922 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n5335) );
  INV_X1 U3923 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n4723) );
  OR2_X1 U3924 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4257) );
  NAND2_X1 U3925 ( .A1(n4343), .A2(n5541), .ZN(n3217) );
  OR2_X1 U3926 ( .A1(n3283), .A2(n3282), .ZN(n3285) );
  INV_X1 U3927 ( .A(n4269), .ZN(n3267) );
  INV_X1 U3928 ( .A(n3404), .ZN(n3344) );
  AOI22_X1 U3929 ( .A1(n3037), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3150) );
  OR2_X1 U3930 ( .A1(n3471), .A2(n3470), .ZN(n3488) );
  AND2_X1 U3931 ( .A1(n4528), .A2(n3246), .ZN(n3416) );
  INV_X1 U3932 ( .A(n3402), .ZN(n3392) );
  OR2_X1 U3933 ( .A1(n3540), .A2(n3539), .ZN(n3568) );
  INV_X1 U3934 ( .A(n3702), .ZN(n3696) );
  OR2_X1 U3935 ( .A1(n6446), .A2(n6479), .ZN(n4260) );
  OR2_X1 U3936 ( .A1(n6053), .A2(n4257), .ZN(n4019) );
  INV_X1 U3937 ( .A(n5002), .ZN(n3841) );
  AND3_X1 U3938 ( .A1(n3347), .A2(n3346), .A3(n3345), .ZN(n3399) );
  NOR2_X1 U3939 ( .A1(n6185), .A2(n5385), .ZN(n5457) );
  OR2_X1 U3940 ( .A1(n5303), .A2(n3971), .ZN(n3972) );
  AND2_X1 U3941 ( .A1(n3638), .A2(n3637), .ZN(n4653) );
  AND2_X1 U3942 ( .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n4076), .ZN(n4077)
         );
  INV_X1 U3943 ( .A(n5601), .ZN(n4021) );
  NAND2_X1 U3944 ( .A1(n5700), .A2(n5683), .ZN(n5684) );
  OAI211_X1 U3945 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n5335), .A(n5334), .B(n5333), .ZN(n5364) );
  NAND2_X1 U3946 ( .A1(n3360), .A2(n3359), .ZN(n5066) );
  AND2_X1 U3947 ( .A1(n5520), .A2(n5463), .ZN(n5500) );
  NOR2_X1 U3948 ( .A1(n3884), .A2(n3885), .ZN(n3899) );
  AND2_X1 U3949 ( .A1(n3833), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3852)
         );
  OR2_X1 U3950 ( .A1(n5384), .A2(n5335), .ZN(n5180) );
  NAND2_X1 U3951 ( .A1(n3994), .A2(n3993), .ZN(n5315) );
  XNOR2_X1 U3952 ( .A(n4275), .B(n4274), .ZN(n5132) );
  AND2_X1 U3953 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n3828), .ZN(n3833)
         );
  OR2_X1 U3954 ( .A1(n6481), .A2(n6486), .ZN(n4289) );
  OR2_X1 U3955 ( .A1(n4269), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U3956 ( .A1(n3423), .A2(n3615), .ZN(n4408) );
  OR3_X1 U3957 ( .A1(n4773), .A2(n5860), .A3(n4772), .ZN(n5881) );
  NOR2_X1 U3958 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4494), .ZN(n4961) );
  INV_X1 U3959 ( .A(n6407), .ZN(n4891) );
  OR2_X1 U3960 ( .A1(n4852), .A2(n5856), .ZN(n4939) );
  INV_X1 U3961 ( .A(n5860), .ZN(n4758) );
  NOR2_X1 U3962 ( .A1(n4289), .A2(n4288), .ZN(n4308) );
  NOR2_X1 U3963 ( .A1(n6535), .A2(n6058), .ZN(n5960) );
  NAND2_X1 U3964 ( .A1(n3772), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3936)
         );
  NOR2_X1 U3965 ( .A1(n6586), .A2(n5123), .ZN(n5384) );
  INV_X1 U3966 ( .A(n6115), .ZN(n6178) );
  OR2_X1 U3967 ( .A1(n5464), .A2(n5143), .ZN(n6172) );
  INV_X1 U3968 ( .A(n6195), .ZN(n5559) );
  AND2_X1 U3969 ( .A1(n5613), .A2(n5612), .ZN(n5614) );
  AND2_X1 U3970 ( .A1(n5613), .A2(n4431), .ZN(n5375) );
  NOR2_X1 U3971 ( .A1(n6209), .A2(n6588), .ZN(n6238) );
  OR2_X1 U3972 ( .A1(n4310), .A2(n4535), .ZN(n4428) );
  INV_X1 U3973 ( .A(n4289), .ZN(n4385) );
  INV_X1 U3974 ( .A(n5660), .ZN(n5664) );
  NOR2_X1 U3975 ( .A1(n5983), .A2(n3740), .ZN(n5841) );
  INV_X1 U3976 ( .A(n6308), .ZN(n6284) );
  AND2_X1 U3977 ( .A1(n3722), .A2(n3707), .ZN(n6333) );
  INV_X1 U3978 ( .A(n4961), .ZN(n4856) );
  NOR2_X1 U3979 ( .A1(n4696), .A2(n4810), .ZN(n4716) );
  OAI21_X1 U3980 ( .B1(n5013), .B2(n5014), .A(n5334), .ZN(n5039) );
  INV_X1 U3981 ( .A(n4771), .ZN(n5043) );
  INV_X1 U3982 ( .A(n5881), .ZN(n5914) );
  AND2_X1 U3983 ( .A1(n4811), .A2(n4810), .ZN(n6392) );
  AND2_X1 U3984 ( .A1(n4805), .A2(n4675), .ZN(n6407) );
  INV_X1 U3985 ( .A(n4959), .ZN(n4893) );
  NOR2_X2 U3986 ( .A1(n4939), .A2(n3815), .ZN(n5368) );
  INV_X1 U3987 ( .A(n5115), .ZN(n6438) );
  OR2_X1 U3988 ( .A1(n5070), .A2(n5069), .ZN(n5105) );
  NAND2_X1 U3989 ( .A1(n4773), .A2(n4758), .ZN(n4852) );
  AND2_X1 U3990 ( .A1(n4635), .A2(n3815), .ZN(n5110) );
  INV_X1 U3991 ( .A(n3815), .ZN(n4810) );
  AND2_X1 U3992 ( .A1(n4489), .A2(n5860), .ZN(n4996) );
  AND2_X1 U3993 ( .A1(n6474), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3598) );
  INV_X1 U3994 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6474) );
  OR2_X1 U3995 ( .A1(n4308), .A2(n4302), .ZN(n6586) );
  OR2_X1 U3996 ( .A1(n5384), .A2(n6567), .ZN(n6115) );
  INV_X1 U3997 ( .A(n6158), .ZN(n6175) );
  OR2_X1 U3998 ( .A1(n5384), .A2(n5125), .ZN(n6151) );
  OR2_X1 U3999 ( .A1(n5384), .A2(n5133), .ZN(n6161) );
  NAND2_X1 U4000 ( .A1(n6195), .A2(n5612), .ZN(n5608) );
  INV_X1 U4001 ( .A(n6100), .ZN(n5294) );
  INV_X1 U4002 ( .A(n5375), .ZN(n4757) );
  INV_X1 U4003 ( .A(n6209), .ZN(n6241) );
  AOI21_X1 U4004 ( .B1(n6276), .B2(n5482), .A(n4285), .ZN(n4286) );
  NAND2_X1 U4005 ( .A1(n6297), .A2(n4270), .ZN(n6282) );
  AND2_X1 U4006 ( .A1(n3744), .A2(n3103), .ZN(n3745) );
  INV_X1 U4007 ( .A(n6331), .ZN(n6010) );
  INV_X1 U4008 ( .A(n4716), .ZN(n4754) );
  NAND2_X1 U4009 ( .A1(n4689), .A2(n4810), .ZN(n5046) );
  NAND2_X1 U4010 ( .A1(n4805), .A2(n4674), .ZN(n6415) );
  AOI21_X1 U4011 ( .B1(n4859), .B2(n4858), .A(n4857), .ZN(n4896) );
  NAND2_X1 U4012 ( .A1(n4853), .A2(n3815), .ZN(n4959) );
  OR2_X1 U4013 ( .A1(n4852), .A2(n4770), .ZN(n6444) );
  OR2_X1 U4014 ( .A1(n4852), .A2(n4772), .ZN(n5115) );
  NAND2_X1 U4015 ( .A1(n4635), .A2(n4810), .ZN(n4999) );
  INV_X1 U4016 ( .A(n4751), .ZN(n4668) );
  INV_X1 U4017 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6567) );
  OAI211_X1 U4018 ( .C1(n5759), .C2(n6297), .A(n3043), .B(n4286), .ZN(U2957)
         );
  OAI21_X1 U4019 ( .B1(n5442), .B2(n6307), .A(n3745), .ZN(U2991) );
  AND2_X4 U4020 ( .A1(n4578), .A2(n4351), .ZN(n4239) );
  NOR2_X4 U4021 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4352) );
  AOI22_X1 U4022 ( .A1(n4239), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3112) );
  AOI22_X1 U4023 ( .A1(n4222), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3203), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3111) );
  AOI22_X1 U4024 ( .A1(n3035), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3110) );
  INV_X1 U4025 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3108) );
  AND2_X2 U4026 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n3108), .ZN(n3114)
         );
  AOI22_X1 U4027 ( .A1(n3292), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3109) );
  AND2_X4 U4028 ( .A1(n3114), .A2(n4352), .ZN(n4140) );
  AOI22_X1 U4029 ( .A1(n4245), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3118) );
  AND2_X4 U4030 ( .A1(n3114), .A2(n3113), .ZN(n3311) );
  AND2_X2 U4031 ( .A1(n4357), .A2(n4573), .ZN(n3310) );
  AOI22_X1 U4032 ( .A1(n3310), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3116) );
  AOI22_X1 U4033 ( .A1(n4183), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U4034 ( .A1(n4239), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3029), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3124) );
  AOI22_X1 U4035 ( .A1(n3025), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3123) );
  AOI22_X1 U4036 ( .A1(n4245), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3122) );
  AOI22_X1 U4037 ( .A1(n3034), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3121) );
  AOI22_X1 U4038 ( .A1(n3310), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3128) );
  AOI22_X1 U4039 ( .A1(n3313), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3127) );
  AOI22_X1 U4040 ( .A1(n3331), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3126) );
  AOI22_X1 U4041 ( .A1(n4239), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3134) );
  AOI22_X1 U4042 ( .A1(n3025), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3310), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3133) );
  AOI22_X1 U4043 ( .A1(n4245), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3132) );
  AOI22_X1 U4044 ( .A1(n3277), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3131) );
  AOI22_X1 U4045 ( .A1(n3311), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3138) );
  AOI22_X1 U4046 ( .A1(n3035), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3028), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3137) );
  AOI22_X1 U4047 ( .A1(n4222), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3136) );
  AOI22_X1 U4048 ( .A1(n3203), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3135) );
  AND3_X2 U4049 ( .A1(n3105), .A2(n3138), .A3(n3042), .ZN(n4514) );
  AOI22_X1 U4050 ( .A1(n3310), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3203), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3142) );
  AOI22_X1 U4051 ( .A1(n3311), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3141) );
  AOI22_X1 U4052 ( .A1(n3025), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3140) );
  AOI22_X1 U4053 ( .A1(n4245), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3139) );
  NAND4_X1 U4054 ( .A1(n3142), .A2(n3141), .A3(n3140), .A4(n3139), .ZN(n3148)
         );
  AOI22_X1 U4055 ( .A1(n3034), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3145) );
  AOI22_X1 U4056 ( .A1(n4222), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3144) );
  AOI22_X1 U4057 ( .A1(n3028), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3143) );
  NAND4_X1 U4058 ( .A1(n3146), .A2(n3145), .A3(n3144), .A4(n3143), .ZN(n3147)
         );
  OR2_X2 U4059 ( .A1(n3148), .A2(n3147), .ZN(n5445) );
  AOI21_X1 U4060 ( .B1(n4376), .B2(n4514), .A(n5612), .ZN(n3159) );
  AOI22_X1 U4061 ( .A1(n3311), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3152) );
  AOI22_X1 U4062 ( .A1(n3310), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3203), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U4063 ( .A1(n3025), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3149) );
  AOI22_X1 U4064 ( .A1(n3032), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3156) );
  AOI22_X1 U4065 ( .A1(n3034), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3155) );
  NAND2_X1 U4066 ( .A1(n3045), .A2(n3816), .ZN(n3247) );
  NAND2_X1 U4067 ( .A1(n3247), .A2(n3708), .ZN(n3181) );
  NAND2_X1 U4068 ( .A1(n3034), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3163) );
  NAND2_X1 U4069 ( .A1(n3367), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3162)
         );
  NAND2_X1 U4070 ( .A1(n4183), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3161) );
  NAND2_X1 U4071 ( .A1(n3277), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3160)
         );
  NAND2_X1 U4072 ( .A1(n3310), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3167) );
  NAND2_X1 U4073 ( .A1(n3203), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3166) );
  NAND2_X1 U4074 ( .A1(n3311), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3165) );
  NAND2_X1 U4075 ( .A1(n3292), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3164) );
  NAND2_X1 U4076 ( .A1(n3026), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3173)
         );
  NAND2_X1 U4077 ( .A1(n4245), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3172)
         );
  NAND2_X1 U4078 ( .A1(n3331), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3171) );
  NAND2_X1 U4079 ( .A1(n4140), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3170) );
  NAND2_X1 U4080 ( .A1(n4239), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3177)
         );
  NAND2_X1 U4081 ( .A1(n3275), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3176) );
  NAND2_X1 U4082 ( .A1(n4222), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3175)
         );
  NAND2_X1 U4083 ( .A1(n2996), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3174) );
  NAND3_X1 U4084 ( .A1(n3249), .A2(n3181), .A3(n4535), .ZN(n3202) );
  NAND2_X1 U4085 ( .A1(n3035), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3185) );
  NAND2_X1 U4086 ( .A1(n3203), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3184) );
  NAND2_X1 U4087 ( .A1(n3275), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3183) );
  NAND2_X1 U4088 ( .A1(n4183), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3182) );
  NAND2_X1 U4089 ( .A1(n3292), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3189) );
  NAND2_X1 U4090 ( .A1(n3310), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3188) );
  NAND2_X1 U4091 ( .A1(n3026), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3187)
         );
  NAND2_X1 U4092 ( .A1(n3311), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3186) );
  NAND2_X1 U4093 ( .A1(n4245), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3192)
         );
  NAND2_X1 U4094 ( .A1(n3331), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3191) );
  NAND2_X1 U4095 ( .A1(n4239), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3197)
         );
  NAND2_X1 U4096 ( .A1(n3277), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3196)
         );
  NAND2_X1 U4097 ( .A1(n2996), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3195) );
  NAND2_X1 U4098 ( .A1(n3367), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3194)
         );
  NAND4_X4 U4099 ( .A1(n3201), .A2(n3200), .A3(n3199), .A4(n3198), .ZN(n3606)
         );
  NAND2_X1 U4100 ( .A1(n3202), .A2(n4528), .ZN(n3215) );
  AOI22_X1 U4101 ( .A1(n3310), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3203), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3207) );
  AOI22_X1 U4102 ( .A1(n3311), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3206) );
  AOI22_X1 U4103 ( .A1(n3025), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3205) );
  AOI22_X1 U4104 ( .A1(n4245), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3204) );
  NAND4_X1 U4105 ( .A1(n3207), .A2(n3206), .A3(n3205), .A4(n3204), .ZN(n3213)
         );
  AOI22_X1 U4106 ( .A1(n3028), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3211) );
  AOI22_X1 U4107 ( .A1(n4239), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3275), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U4108 ( .A1(n4222), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3209) );
  AOI22_X1 U4109 ( .A1(n3035), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3208) );
  NAND4_X1 U4110 ( .A1(n3211), .A2(n3210), .A3(n3209), .A4(n3208), .ZN(n3212)
         );
  NAND2_X1 U4111 ( .A1(n3416), .A2(n4429), .ZN(n3214) );
  NAND2_X1 U4112 ( .A1(n3215), .A2(n3214), .ZN(n3240) );
  NAND2_X1 U4113 ( .A1(n3045), .A2(n5445), .ZN(n3593) );
  NAND2_X1 U4114 ( .A1(n3593), .A2(n5139), .ZN(n3218) );
  AND2_X4 U4115 ( .A1(n3600), .A2(n3246), .ZN(n5541) );
  AND2_X1 U4116 ( .A1(n4376), .A2(n5445), .ZN(n3220) );
  NOR2_X1 U4117 ( .A1(n4344), .A2(n3710), .ZN(n3589) );
  XNOR2_X1 U4118 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n3522) );
  NAND2_X1 U4119 ( .A1(n4535), .A2(n3522), .ZN(n3245) );
  NAND2_X1 U4120 ( .A1(n3245), .A2(n3222), .ZN(n3223) );
  NAND3_X1 U4121 ( .A1(n3230), .A2(n3589), .A3(n3223), .ZN(n3224) );
  NAND2_X1 U4122 ( .A1(n3226), .A2(n3225), .ZN(n3262) );
  NAND2_X1 U4123 ( .A1(n3262), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3229) );
  INV_X1 U4124 ( .A(n3598), .ZN(n3266) );
  NAND2_X1 U4125 ( .A1(n6474), .A2(n6567), .ZN(n6575) );
  MUX2_X1 U4126 ( .A(n3266), .B(n3267), .S(n4930), .Z(n3227) );
  INV_X1 U4127 ( .A(n3227), .ZN(n3228) );
  NAND2_X1 U4128 ( .A1(n3229), .A2(n3228), .ZN(n3291) );
  OR2_X1 U4129 ( .A1(n6575), .A2(n6479), .ZN(n6487) );
  INV_X1 U4130 ( .A(n6487), .ZN(n3232) );
  NAND2_X1 U4131 ( .A1(n3710), .A2(n3606), .ZN(n3231) );
  OAI211_X1 U4132 ( .C1(n4429), .C2(n6591), .A(n3232), .B(n3231), .ZN(n3233)
         );
  INV_X1 U4133 ( .A(n3233), .ZN(n3239) );
  NAND2_X1 U4134 ( .A1(n4521), .A2(n4514), .ZN(n3250) );
  NOR2_X1 U4135 ( .A1(n3250), .A2(n3606), .ZN(n3235) );
  NAND2_X1 U4136 ( .A1(n3234), .A2(n3235), .ZN(n4579) );
  NAND2_X1 U4137 ( .A1(n4429), .A2(n3219), .ZN(n3236) );
  NAND2_X1 U4138 ( .A1(n3236), .A2(n3246), .ZN(n3237) );
  OAI21_X1 U4139 ( .B1(n4344), .B2(n3237), .A(n3600), .ZN(n3238) );
  NAND2_X1 U4140 ( .A1(n4343), .A2(n3600), .ZN(n3715) );
  NAND2_X1 U4141 ( .A1(n3240), .A2(n3715), .ZN(n3713) );
  NAND2_X1 U4142 ( .A1(n3291), .A2(n3289), .ZN(n3330) );
  INV_X1 U4143 ( .A(n3330), .ZN(n3261) );
  NAND2_X1 U4144 ( .A1(n3262), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3254) );
  INV_X1 U4145 ( .A(n3593), .ZN(n3244) );
  INV_X1 U4146 ( .A(n3245), .ZN(n3252) );
  NAND2_X1 U4147 ( .A1(n3249), .A2(n3248), .ZN(n3594) );
  INV_X1 U4148 ( .A(n3250), .ZN(n4378) );
  NOR2_X1 U4149 ( .A1(n3600), .A2(n3606), .ZN(n3543) );
  NAND3_X1 U4150 ( .A1(n4378), .A2(n3543), .A3(n3222), .ZN(n4346) );
  NAND2_X1 U4151 ( .A1(n5445), .A2(n3251), .ZN(n3776) );
  OAI211_X1 U4152 ( .C1(n4288), .C2(n3252), .A(n3602), .B(n3706), .ZN(n3253)
         );
  NAND2_X1 U4153 ( .A1(n3253), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3256) );
  XNOR2_X1 U4154 ( .A(n6453), .B(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6344)
         );
  AOI22_X1 U4155 ( .A1(n3267), .A2(n6344), .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n3266), .ZN(n3255) );
  INV_X1 U4156 ( .A(n3255), .ZN(n3258) );
  INV_X1 U4157 ( .A(n3256), .ZN(n3257) );
  OAI21_X1 U4158 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n3258), .A(n3257), 
        .ZN(n3259) );
  OAI21_X2 U4159 ( .B1(n3261), .B2(n3329), .A(n3260), .ZN(n3353) );
  NAND2_X1 U4160 ( .A1(n3262), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3269) );
  AND2_X1 U4161 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3263) );
  NAND2_X1 U4162 ( .A1(n3263), .A2(n6458), .ZN(n4762) );
  INV_X1 U4163 ( .A(n3263), .ZN(n3264) );
  NAND2_X1 U4164 ( .A1(n3264), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3265) );
  NAND2_X1 U4165 ( .A1(n4762), .A2(n3265), .ZN(n4724) );
  AOI22_X1 U4166 ( .A1(n3267), .A2(n4724), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3266), .ZN(n3268) );
  XNOR2_X1 U4167 ( .A(n3353), .B(n3354), .ZN(n4491) );
  AOI22_X1 U4168 ( .A1(n4236), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4169 ( .A1(n3312), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3273) );
  AOI22_X1 U4170 ( .A1(n3038), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3272) );
  AOI22_X1 U4171 ( .A1(n4245), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3271) );
  NAND4_X1 U4172 ( .A1(n3274), .A2(n3273), .A3(n3272), .A4(n3271), .ZN(n3283)
         );
  INV_X1 U4173 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6631) );
  AOI22_X1 U4174 ( .A1(n4239), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3281) );
  BUF_X1 U4175 ( .A(n3277), .Z(n4238) );
  AOI22_X1 U4176 ( .A1(n3035), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3280) );
  AOI22_X1 U4177 ( .A1(n3030), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3279) );
  BUF_X1 U4178 ( .A(n3367), .Z(n3332) );
  AOI22_X1 U4179 ( .A1(n3028), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3278) );
  NAND4_X1 U4180 ( .A1(n3281), .A2(n3280), .A3(n3279), .A4(n3278), .ZN(n3282)
         );
  NOR2_X1 U4181 ( .A1(n3362), .A2(n3394), .ZN(n3284) );
  AOI21_X1 U4182 ( .B1(n4491), .B2(n6479), .A(n3284), .ZN(n3288) );
  INV_X1 U4183 ( .A(n3361), .ZN(n3286) );
  AOI22_X1 U4184 ( .A1(n3566), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3286), 
        .B2(n3285), .ZN(n3287) );
  XNOR2_X1 U4185 ( .A(n3291), .B(n3290), .ZN(n3818) );
  AOI22_X1 U4186 ( .A1(n4239), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3296) );
  AOI22_X1 U4187 ( .A1(n4236), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3203), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3295) );
  AOI22_X1 U4188 ( .A1(n3292), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3294) );
  AOI22_X1 U4189 ( .A1(n3034), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3293) );
  NAND4_X1 U4190 ( .A1(n3296), .A2(n3295), .A3(n3294), .A4(n3293), .ZN(n3302)
         );
  AOI22_X1 U4191 ( .A1(n3038), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3312), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4192 ( .A1(n3305), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4193 ( .A1(n3030), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3298) );
  AOI22_X1 U4194 ( .A1(n4183), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3297) );
  NAND4_X1 U4195 ( .A1(n3300), .A2(n3299), .A3(n3298), .A4(n3297), .ZN(n3301)
         );
  NAND2_X1 U4196 ( .A1(n3270), .A2(n3500), .ZN(n3327) );
  INV_X1 U4197 ( .A(n3500), .ZN(n3303) );
  NAND2_X1 U4198 ( .A1(n3303), .A2(n3270), .ZN(n3320) );
  AOI22_X1 U4199 ( .A1(n4247), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3292), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4200 ( .A1(n3038), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3308) );
  AOI22_X1 U4201 ( .A1(n4245), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4202 ( .A1(n4183), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3306) );
  NAND4_X1 U4203 ( .A1(n3309), .A2(n3308), .A3(n3307), .A4(n3306), .ZN(n3319)
         );
  AOI22_X1 U4204 ( .A1(n4222), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3203), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4205 ( .A1(n4236), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3312), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4206 ( .A1(n3035), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3315) );
  AOI22_X1 U4207 ( .A1(n4239), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3314) );
  NAND4_X1 U4208 ( .A1(n3317), .A2(n3316), .A3(n3315), .A4(n3314), .ZN(n3318)
         );
  MUX2_X1 U4209 ( .A(n3327), .B(n3320), .S(n3417), .Z(n3321) );
  INV_X1 U4210 ( .A(n3321), .ZN(n3322) );
  NAND2_X1 U4211 ( .A1(n3322), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3411) );
  NAND2_X1 U4212 ( .A1(n3409), .A2(n3411), .ZN(n3326) );
  NAND2_X1 U4213 ( .A1(n3566), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3325) );
  AOI21_X1 U4214 ( .B1(n4528), .B2(n3417), .A(n6479), .ZN(n3323) );
  AND2_X1 U4215 ( .A1(n3323), .A2(n3327), .ZN(n3324) );
  NAND2_X1 U4216 ( .A1(n3325), .A2(n3324), .ZN(n3412) );
  NAND2_X1 U4217 ( .A1(n3326), .A2(n3412), .ZN(n3328) );
  XNOR2_X1 U4218 ( .A(n3330), .B(n3329), .ZN(n4341) );
  AOI22_X1 U4219 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n4246), .B1(n4244), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4220 ( .A1(n4127), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4221 ( .A1(n3312), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4222 ( .A1(n4236), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3333) );
  NAND4_X1 U4223 ( .A1(n3336), .A2(n3335), .A3(n3334), .A4(n3333), .ZN(n3342)
         );
  AOI22_X1 U4224 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n4239), .B1(n4222), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4225 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n3038), .B1(n4199), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4226 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n4237), .B1(n3028), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4227 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4247), .B1(n4238), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3337) );
  NAND4_X1 U4228 ( .A1(n3340), .A2(n3339), .A3(n3338), .A4(n3337), .ZN(n3341)
         );
  OAI21_X1 U4229 ( .B1(n4341), .B2(STATE2_REG_0__SCAN_IN), .A(n3343), .ZN(
        n3349) );
  NAND2_X1 U4230 ( .A1(n3350), .A2(n3349), .ZN(n3348) );
  NAND2_X1 U4231 ( .A1(n3566), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3347) );
  OR2_X1 U4232 ( .A1(n3362), .A2(n3500), .ZN(n3346) );
  OR2_X1 U4233 ( .A1(n3361), .A2(n3344), .ZN(n3345) );
  NAND2_X1 U4234 ( .A1(n3348), .A2(n3399), .ZN(n3352) );
  INV_X1 U4235 ( .A(n3349), .ZN(n3398) );
  INV_X1 U4236 ( .A(n3350), .ZN(n3400) );
  NOR2_X2 U4237 ( .A1(n3393), .A2(n3402), .ZN(n3425) );
  INV_X1 U4238 ( .A(n3353), .ZN(n3355) );
  NAND2_X1 U4239 ( .A1(n3262), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3360) );
  NAND3_X1 U4240 ( .A1(n6357), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6343) );
  INV_X1 U4241 ( .A(n6343), .ZN(n3356) );
  NAND2_X1 U4242 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3356), .ZN(n4540) );
  NAND2_X1 U4243 ( .A1(n6357), .A2(n4540), .ZN(n3357) );
  NAND3_X1 U4244 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4960) );
  INV_X1 U4245 ( .A(n4960), .ZN(n4493) );
  NAND2_X1 U4246 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4493), .ZN(n4663) );
  NAND2_X1 U4247 ( .A1(n3357), .A2(n4663), .ZN(n4855) );
  OAI22_X1 U4248 ( .A1(n4269), .A2(n4855), .B1(n3598), .B2(n6357), .ZN(n3358)
         );
  INV_X1 U4249 ( .A(n3358), .ZN(n3359) );
  XNOR2_X2 U4250 ( .A(n4589), .B(n5066), .ZN(n4490) );
  AOI22_X1 U4251 ( .A1(n4236), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4252 ( .A1(n3312), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4253 ( .A1(n3038), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4254 ( .A1(n4245), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3363) );
  NAND4_X1 U4255 ( .A1(n3366), .A2(n3365), .A3(n3364), .A4(n3363), .ZN(n3373)
         );
  AOI22_X1 U4256 ( .A1(n3032), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4257 ( .A1(n4127), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4258 ( .A1(n4222), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4259 ( .A1(n4183), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3368) );
  NAND4_X1 U4260 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n3372)
         );
  AOI22_X1 U4261 ( .A1(n3572), .A2(n3429), .B1(n3566), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3374) );
  AOI21_X2 U4262 ( .B1(n4490), .B2(n6479), .A(n3375), .ZN(n4601) );
  INV_X1 U4263 ( .A(n4601), .ZN(n4488) );
  AOI22_X1 U4264 ( .A1(n4127), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3379) );
  AOI22_X1 U4265 ( .A1(n4236), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3378) );
  AOI22_X1 U4266 ( .A1(n3038), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3377) );
  AOI22_X1 U4267 ( .A1(n4183), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3376) );
  NAND4_X1 U4268 ( .A1(n3379), .A2(n3378), .A3(n3377), .A4(n3376), .ZN(n3385)
         );
  AOI22_X1 U4269 ( .A1(n4246), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3312), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4270 ( .A1(n4245), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4271 ( .A1(n4222), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4272 ( .A1(n4247), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3380) );
  NAND4_X1 U4273 ( .A1(n3383), .A2(n3382), .A3(n3381), .A4(n3380), .ZN(n3384)
         );
  NAND2_X1 U4274 ( .A1(n3572), .A2(n3452), .ZN(n3387) );
  NAND2_X1 U4275 ( .A1(n3566), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3386) );
  NAND2_X1 U4276 ( .A1(n3794), .A2(n3792), .ZN(n3389) );
  NAND2_X1 U4277 ( .A1(n3417), .A2(n3404), .ZN(n3403) );
  NAND2_X1 U4278 ( .A1(n3403), .A2(n3394), .ZN(n3428) );
  NAND2_X1 U4279 ( .A1(n3428), .A2(n3429), .ZN(n3454) );
  XNOR2_X1 U4280 ( .A(n3454), .B(n3452), .ZN(n3390) );
  NAND2_X1 U4281 ( .A1(n3390), .A2(n5139), .ZN(n3391) );
  INV_X1 U4282 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3622) );
  XNOR2_X1 U4283 ( .A(n3435), .B(n3622), .ZN(n4607) );
  NAND2_X1 U4284 ( .A1(n3805), .A2(n3548), .ZN(n3397) );
  OAI21_X1 U4285 ( .B1(n3394), .B2(n3403), .A(n3428), .ZN(n3395) );
  AOI21_X1 U4286 ( .B1(n3395), .B2(n5139), .A(n3416), .ZN(n3396) );
  NAND2_X1 U4287 ( .A1(n3422), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4407)
         );
  NAND3_X1 U4288 ( .A1(n3400), .A2(n3398), .A3(n3399), .ZN(n3401) );
  OAI21_X1 U4289 ( .B1(n3417), .B2(n3404), .A(n3403), .ZN(n3406) );
  INV_X1 U4290 ( .A(n3710), .ZN(n3405) );
  OAI211_X1 U4291 ( .C1(n3406), .C2(n6591), .A(n3405), .B(n3242), .ZN(n3407)
         );
  INV_X1 U4292 ( .A(n3407), .ZN(n3408) );
  NAND2_X1 U4293 ( .A1(n3409), .A2(n3412), .ZN(n3410) );
  INV_X1 U4294 ( .A(n3411), .ZN(n3413) );
  NAND2_X1 U4295 ( .A1(n3413), .A2(n3412), .ZN(n3414) );
  INV_X1 U4296 ( .A(n3416), .ZN(n3714) );
  OAI21_X1 U4297 ( .B1(n6591), .B2(n3417), .A(n3714), .ZN(n3418) );
  INV_X1 U4298 ( .A(n3418), .ZN(n3419) );
  XNOR2_X1 U4299 ( .A(n4462), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4439)
         );
  NAND2_X1 U4300 ( .A1(n4440), .A2(n4439), .ZN(n4442) );
  INV_X1 U4301 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3607) );
  OR2_X1 U4302 ( .A1(n4462), .A2(n3607), .ZN(n3421) );
  NAND2_X1 U4303 ( .A1(n4407), .A2(n4410), .ZN(n3424) );
  INV_X1 U4304 ( .A(n3425), .ZN(n3426) );
  NAND2_X1 U4305 ( .A1(n3426), .A2(n4601), .ZN(n3427) );
  OAI211_X1 U4306 ( .C1(n3429), .C2(n3428), .A(n3454), .B(n5139), .ZN(n3430)
         );
  INV_X1 U4307 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3431) );
  XNOR2_X1 U4308 ( .A(n3432), .B(n3431), .ZN(n4447) );
  NAND2_X1 U4309 ( .A1(n4448), .A2(n4447), .ZN(n3434) );
  NAND2_X1 U4310 ( .A1(n3432), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3433)
         );
  NAND2_X1 U4311 ( .A1(n3434), .A2(n3433), .ZN(n4608) );
  NAND2_X1 U4312 ( .A1(n4607), .A2(n4608), .ZN(n3437) );
  NAND2_X1 U4313 ( .A1(n3435), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3436)
         );
  NAND2_X1 U4314 ( .A1(n3437), .A2(n3436), .ZN(n4906) );
  AOI22_X1 U4315 ( .A1(n4236), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3441) );
  AOI22_X1 U4316 ( .A1(n3312), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3440) );
  AOI22_X1 U4317 ( .A1(n3038), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4318 ( .A1(n4245), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3438) );
  NAND4_X1 U4319 ( .A1(n3441), .A2(n3440), .A3(n3439), .A4(n3438), .ZN(n3447)
         );
  AOI22_X1 U4320 ( .A1(n3032), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4321 ( .A1(n4127), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3444) );
  AOI22_X1 U4322 ( .A1(n4222), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3443) );
  INV_X1 U4323 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n6759) );
  AOI22_X1 U4324 ( .A1(n3028), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3442) );
  NAND4_X1 U4325 ( .A1(n3445), .A2(n3444), .A3(n3443), .A4(n3442), .ZN(n3446)
         );
  NAND2_X1 U4326 ( .A1(n3572), .A2(n3455), .ZN(n3449) );
  NAND2_X1 U4327 ( .A1(n3566), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3448) );
  NAND2_X1 U4328 ( .A1(n3450), .A2(n3048), .ZN(n3451) );
  NAND2_X1 U4329 ( .A1(n3791), .A2(n3451), .ZN(n3458) );
  INV_X1 U4330 ( .A(n3452), .ZN(n3453) );
  NOR2_X1 U4331 ( .A1(n3454), .A2(n3453), .ZN(n3456) );
  NAND2_X1 U4332 ( .A1(n3456), .A2(n3455), .ZN(n3487) );
  OAI211_X1 U4333 ( .C1(n3456), .C2(n3455), .A(n3487), .B(n5139), .ZN(n3457)
         );
  XNOR2_X1 U4334 ( .A(n3459), .B(n4909), .ZN(n4907) );
  NAND2_X1 U4335 ( .A1(n4906), .A2(n4907), .ZN(n3461) );
  NAND2_X1 U4336 ( .A1(n3459), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3460)
         );
  NAND2_X1 U4337 ( .A1(n3461), .A2(n3460), .ZN(n4897) );
  AOI22_X1 U4338 ( .A1(n3032), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U4339 ( .A1(n4236), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4340 ( .A1(n3305), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3463) );
  AOI22_X1 U4341 ( .A1(n4238), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3462) );
  NAND4_X1 U4342 ( .A1(n3465), .A2(n3464), .A3(n3463), .A4(n3462), .ZN(n3471)
         );
  AOI22_X1 U4343 ( .A1(n3030), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3312), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4344 ( .A1(n3038), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4345 ( .A1(n4127), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4346 ( .A1(n4247), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3466) );
  NAND4_X1 U4347 ( .A1(n3469), .A2(n3468), .A3(n3467), .A4(n3466), .ZN(n3470)
         );
  NAND2_X1 U4348 ( .A1(n3572), .A2(n3488), .ZN(n3473) );
  NAND2_X1 U4349 ( .A1(n3566), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3472) );
  INV_X1 U4350 ( .A(n3827), .ZN(n3479) );
  XNOR2_X1 U4351 ( .A(n3487), .B(n3488), .ZN(n3477) );
  NAND2_X1 U4352 ( .A1(n3477), .A2(n5139), .ZN(n3478) );
  INV_X1 U4353 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3634) );
  XNOR2_X1 U4354 ( .A(n3480), .B(n3634), .ZN(n4898) );
  NAND2_X1 U4355 ( .A1(n4897), .A2(n4898), .ZN(n3482) );
  NAND2_X1 U4356 ( .A1(n3480), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3481)
         );
  NAND2_X1 U4357 ( .A1(n3482), .A2(n3481), .ZN(n5151) );
  NAND2_X1 U4358 ( .A1(n3572), .A2(n3500), .ZN(n3484) );
  NAND2_X1 U4359 ( .A1(n3566), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3483) );
  NAND2_X1 U4360 ( .A1(n3484), .A2(n3483), .ZN(n3485) );
  INV_X1 U4361 ( .A(n3487), .ZN(n3489) );
  NAND2_X1 U4362 ( .A1(n3489), .A2(n3488), .ZN(n3499) );
  XNOR2_X1 U4363 ( .A(n3499), .B(n3500), .ZN(n3490) );
  NAND2_X1 U4364 ( .A1(n3490), .A2(n5139), .ZN(n3491) );
  NAND2_X1 U4365 ( .A1(n3492), .A2(n3491), .ZN(n3494) );
  INV_X1 U4366 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3493) );
  XNOR2_X1 U4367 ( .A(n3494), .B(n3493), .ZN(n5152) );
  NAND2_X1 U4368 ( .A1(n5151), .A2(n5152), .ZN(n3496) );
  NAND2_X1 U4369 ( .A1(n3494), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3495)
         );
  NAND2_X1 U4370 ( .A1(n3003), .A2(n3495), .ZN(n5163) );
  INV_X1 U4371 ( .A(n3499), .ZN(n3501) );
  NAND3_X1 U4372 ( .A1(n3501), .A2(n5139), .A3(n3500), .ZN(n3502) );
  NAND2_X1 U4373 ( .A1(n3508), .A2(n3502), .ZN(n3503) );
  INV_X1 U4374 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3641) );
  XNOR2_X1 U4375 ( .A(n3503), .B(n3641), .ZN(n5164) );
  NAND2_X1 U4376 ( .A1(n3503), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3504)
         );
  INV_X1 U4377 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6326) );
  NOR2_X1 U4378 ( .A1(n3007), .A2(n6326), .ZN(n3505) );
  INV_X4 U4379 ( .A(n3506), .ZN(n5727) );
  NAND2_X1 U4380 ( .A1(n3508), .A2(n6326), .ZN(n3507) );
  INV_X1 U4381 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6317) );
  AND2_X1 U4382 ( .A1(n3508), .A2(n6317), .ZN(n5210) );
  NAND2_X1 U4383 ( .A1(n3031), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5211) );
  INV_X1 U4384 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5261) );
  NAND2_X1 U4385 ( .A1(n3007), .A2(n5261), .ZN(n5255) );
  NAND2_X1 U4386 ( .A1(n3506), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5256) );
  INV_X1 U4387 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3654) );
  NOR2_X1 U4388 ( .A1(n5727), .A2(n3654), .ZN(n5271) );
  NAND2_X1 U4389 ( .A1(n5727), .A2(n3654), .ZN(n5269) );
  XNOR2_X1 U4390 ( .A(n5727), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5974)
         );
  INV_X1 U4391 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6004) );
  NAND2_X1 U4392 ( .A1(n5727), .A2(n6004), .ZN(n5393) );
  INV_X1 U4393 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6003) );
  NAND2_X1 U4394 ( .A1(n5727), .A2(n6003), .ZN(n3509) );
  NAND2_X1 U4395 ( .A1(n3506), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3510) );
  INV_X1 U4396 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6000) );
  INV_X1 U4397 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5992) );
  NAND2_X1 U4398 ( .A1(n5727), .A2(n5992), .ZN(n5736) );
  NAND2_X1 U4399 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3740) );
  NAND2_X1 U4400 ( .A1(n3506), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5737) );
  OAI21_X1 U4401 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n3506), .ZN(n3514) );
  INV_X1 U4402 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3516) );
  NOR2_X1 U4403 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5809) );
  INV_X1 U4404 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5803) );
  INV_X1 U4405 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3677) );
  INV_X1 U4406 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5792) );
  NAND4_X1 U4407 ( .A1(n5809), .A2(n5803), .A3(n3677), .A4(n5792), .ZN(n3519)
         );
  AND2_X1 U4408 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5790) );
  AND2_X1 U4409 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5810) );
  AND2_X1 U4410 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3727) );
  AND3_X1 U4411 ( .A1(n5790), .A2(n5810), .A3(n3727), .ZN(n3741) );
  NAND2_X1 U4412 ( .A1(n3517), .A2(n3741), .ZN(n3518) );
  XNOR2_X1 U4413 ( .A(n5727), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5674)
         );
  INV_X1 U4414 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5786) );
  NAND2_X1 U4415 ( .A1(n5727), .A2(n5786), .ZN(n3520) );
  NAND2_X1 U4416 ( .A1(n5727), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5661) );
  INV_X1 U4417 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5776) );
  NAND2_X1 U4418 ( .A1(n3506), .A2(n5776), .ZN(n5662) );
  NOR2_X1 U4419 ( .A1(n3747), .A2(n5652), .ZN(n3521) );
  INV_X1 U4420 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5647) );
  XNOR2_X1 U4421 ( .A(n3521), .B(n5647), .ZN(n5442) );
  INV_X1 U4422 ( .A(n3522), .ZN(n3523) );
  INV_X1 U4423 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U4424 ( .A1(n3523), .A2(n6506), .ZN(n6501) );
  XNOR2_X1 U4425 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3533) );
  NAND2_X1 U4426 ( .A1(n4930), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3545) );
  INV_X1 U4427 ( .A(n3545), .ZN(n3524) );
  NAND2_X1 U4428 ( .A1(n3533), .A2(n3524), .ZN(n3526) );
  NAND2_X1 U4429 ( .A1(n6453), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3525) );
  NAND2_X1 U4430 ( .A1(n3526), .A2(n3525), .ZN(n3534) );
  XNOR2_X1 U4431 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3535) );
  NAND2_X1 U4432 ( .A1(n3534), .A2(n3535), .ZN(n3528) );
  NAND2_X1 U4433 ( .A1(n6458), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3527) );
  NAND2_X1 U4434 ( .A1(n3528), .A2(n3527), .ZN(n3536) );
  XNOR2_X1 U4435 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3537) );
  NAND2_X1 U4436 ( .A1(n3536), .A2(n3537), .ZN(n3530) );
  NAND2_X1 U4437 ( .A1(n6357), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3529) );
  NAND2_X1 U4438 ( .A1(n3530), .A2(n3529), .ZN(n3540) );
  AND2_X1 U4439 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6738), .ZN(n3531)
         );
  INV_X1 U4440 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3779) );
  NAND2_X1 U4441 ( .A1(n3779), .A2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n3539) );
  XNOR2_X1 U4442 ( .A(n3533), .B(n3545), .ZN(n3549) );
  XOR2_X1 U4443 ( .A(n3535), .B(n3534), .Z(n3558) );
  XOR2_X1 U4444 ( .A(n3537), .B(n3536), .Z(n3567) );
  AND3_X1 U4445 ( .A1(n3549), .A2(n3558), .A3(n3567), .ZN(n3538) );
  OR2_X1 U4446 ( .A1(n3575), .A2(n3538), .ZN(n3541) );
  NAND2_X1 U4447 ( .A1(n3541), .A2(n3568), .ZN(n4294) );
  INV_X1 U4448 ( .A(n4294), .ZN(n4287) );
  NOR2_X1 U4449 ( .A1(n4287), .A2(READY_N), .ZN(n4365) );
  INV_X1 U4450 ( .A(n4365), .ZN(n3542) );
  AOI21_X1 U4451 ( .B1(n3600), .B2(n6501), .A(n3542), .ZN(n3585) );
  AOI21_X1 U4452 ( .B1(n3572), .B2(n3600), .A(n3222), .ZN(n3557) );
  NAND2_X1 U4453 ( .A1(n3549), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3556) );
  AND2_X1 U4454 ( .A1(n4535), .A2(n3242), .ZN(n3544) );
  NOR2_X1 U4455 ( .A1(n3543), .A2(n3544), .ZN(n3562) );
  OAI21_X1 U4456 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n4930), .A(n3545), 
        .ZN(n3550) );
  OAI21_X1 U4457 ( .B1(n4343), .B2(n3550), .A(n3546), .ZN(n3547) );
  AOI22_X1 U4458 ( .A1(n3557), .A2(n3556), .B1(n3562), .B2(n3547), .ZN(n3554)
         );
  NOR2_X1 U4459 ( .A1(n3577), .A2(n3549), .ZN(n3553) );
  INV_X1 U4460 ( .A(n3572), .ZN(n3551) );
  OAI21_X1 U4461 ( .B1(n3551), .B2(n3550), .A(n3577), .ZN(n3552) );
  OAI21_X1 U4462 ( .B1(n3554), .B2(n3553), .A(n3552), .ZN(n3555) );
  OAI21_X1 U4463 ( .B1(n3557), .B2(n3556), .A(n3555), .ZN(n3565) );
  INV_X1 U4464 ( .A(n3566), .ZN(n3559) );
  NAND2_X1 U4465 ( .A1(n3572), .A2(n3558), .ZN(n3561) );
  OAI211_X1 U4466 ( .C1(n3559), .C2(n3558), .A(n3562), .B(n3561), .ZN(n3564)
         );
  OAI22_X1 U4467 ( .A1(n3562), .A2(n3561), .B1(n3567), .B2(n3560), .ZN(n3563)
         );
  AOI21_X1 U4468 ( .B1(n3565), .B2(n3564), .A(n3563), .ZN(n3570) );
  AOI21_X1 U4469 ( .B1(n3567), .B2(n3568), .A(n3566), .ZN(n3569) );
  OAI22_X1 U4470 ( .A1(n3570), .A2(n3569), .B1(n3577), .B2(n3568), .ZN(n3571)
         );
  AOI21_X1 U4471 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6479), .A(n3571), 
        .ZN(n3574) );
  NAND2_X1 U4472 ( .A1(n3572), .A2(n3575), .ZN(n3573) );
  NAND2_X1 U4473 ( .A1(n3574), .A2(n3573), .ZN(n3579) );
  INV_X1 U4474 ( .A(n3575), .ZN(n3576) );
  NAND2_X1 U4475 ( .A1(n4535), .A2(n6501), .ZN(n5127) );
  INV_X1 U4476 ( .A(READY_N), .ZN(n4307) );
  NAND2_X1 U4477 ( .A1(n5127), .A2(n4307), .ZN(n3581) );
  OAI211_X1 U4478 ( .C1(n3580), .C2(n3581), .A(n3606), .B(n3776), .ZN(n3582)
         );
  INV_X1 U4479 ( .A(n3582), .ZN(n3583) );
  NOR2_X1 U4480 ( .A1(n6481), .A2(n3583), .ZN(n3584) );
  MUX2_X1 U4481 ( .A(n3585), .B(n3584), .S(n4514), .Z(n3586) );
  INV_X1 U4482 ( .A(n3586), .ZN(n3597) );
  NAND2_X1 U4483 ( .A1(n3234), .A2(n3242), .ZN(n6446) );
  NOR2_X1 U4484 ( .A1(n6446), .A2(n4535), .ZN(n3587) );
  NAND2_X1 U4485 ( .A1(n6481), .A2(n3587), .ZN(n4358) );
  NAND2_X1 U4486 ( .A1(n6446), .A2(n4528), .ZN(n3588) );
  AND2_X1 U4487 ( .A1(n3589), .A2(n3588), .ZN(n3603) );
  INV_X1 U4488 ( .A(n4429), .ZN(n3592) );
  NAND2_X1 U4489 ( .A1(n4429), .A2(n3606), .ZN(n3590) );
  NAND2_X1 U4490 ( .A1(n6591), .A2(n3590), .ZN(n3591) );
  OAI21_X1 U4491 ( .B1(n3593), .B2(n3592), .A(n3591), .ZN(n4347) );
  NAND2_X1 U4492 ( .A1(n3603), .A2(n4347), .ZN(n3595) );
  NAND2_X1 U4493 ( .A1(n3595), .A2(n3594), .ZN(n4362) );
  AND2_X1 U4494 ( .A1(n4358), .A2(n4362), .ZN(n3596) );
  NAND2_X1 U4495 ( .A1(n3597), .A2(n3596), .ZN(n3599) );
  NAND2_X1 U4496 ( .A1(n3598), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6486) );
  INV_X1 U4497 ( .A(n6486), .ZN(n4424) );
  AND2_X1 U4498 ( .A1(n3603), .A2(n4343), .ZN(n3770) );
  INV_X1 U4499 ( .A(n3770), .ZN(n6464) );
  OAI22_X1 U4500 ( .A1(n3580), .A2(n4379), .B1(n3270), .B2(n3706), .ZN(n3601)
         );
  INV_X1 U4501 ( .A(n3601), .ZN(n3604) );
  NAND2_X1 U4502 ( .A1(n3603), .A2(n3543), .ZN(n4565) );
  NAND4_X1 U4503 ( .A1(n6464), .A2(n3604), .A3(n2999), .A4(n4565), .ZN(n3605)
         );
  AND2_X4 U4504 ( .A1(n5541), .A2(n5134), .ZN(n3750) );
  INV_X1 U4505 ( .A(EBX_REG_1__SCAN_IN), .ZN(n5254) );
  NAND2_X1 U4506 ( .A1(n3750), .A2(n5254), .ZN(n3611) );
  NAND2_X2 U4507 ( .A1(n4521), .A2(n3606), .ZN(n3751) );
  NAND2_X1 U4508 ( .A1(n3751), .A2(n3607), .ZN(n3609) );
  NAND2_X1 U4509 ( .A1(n5134), .A2(n5254), .ZN(n3608) );
  NAND3_X1 U4510 ( .A1(n3609), .A2(n5596), .A3(n3608), .ZN(n3610) );
  NAND2_X1 U4511 ( .A1(n3751), .A2(EBX_REG_0__SCAN_IN), .ZN(n3612) );
  OAI21_X1 U4512 ( .B1(n5541), .B2(EBX_REG_0__SCAN_IN), .A(n3612), .ZN(n4373)
         );
  XNOR2_X1 U4513 ( .A(n3613), .B(n4373), .ZN(n5250) );
  INV_X1 U4514 ( .A(n3613), .ZN(n3614) );
  INV_X1 U4515 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3615) );
  NAND2_X1 U4516 ( .A1(n3751), .A2(n3615), .ZN(n3617) );
  INV_X1 U4517 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6707) );
  NAND2_X1 U4518 ( .A1(n5134), .A2(n6707), .ZN(n3616) );
  NAND3_X1 U4519 ( .A1(n3617), .A2(n5596), .A3(n3616), .ZN(n3618) );
  OAI21_X1 U4520 ( .B1(n3757), .B2(EBX_REG_2__SCAN_IN), .A(n3618), .ZN(n4412)
         );
  MUX2_X1 U4521 ( .A(n3702), .B(n5596), .S(EBX_REG_3__SCAN_IN), .Z(n3620) );
  NAND2_X1 U4522 ( .A1(n3756), .A2(n3431), .ZN(n3619) );
  NAND2_X1 U4523 ( .A1(n3620), .A2(n3619), .ZN(n4454) );
  INV_X1 U4524 ( .A(n4454), .ZN(n3621) );
  OAI21_X1 U4525 ( .B1(n5541), .B2(n3622), .A(n3751), .ZN(n3623) );
  OAI21_X1 U4526 ( .B1(EBX_REG_4__SCAN_IN), .B2(n4379), .A(n3623), .ZN(n3626)
         );
  INV_X1 U4527 ( .A(EBX_REG_4__SCAN_IN), .ZN(n3624) );
  NAND2_X1 U4528 ( .A1(n3750), .A2(n3624), .ZN(n3625) );
  INV_X1 U4529 ( .A(EBX_REG_5__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U4530 ( .A1(n3696), .A2(n6194), .ZN(n3631) );
  INV_X1 U4531 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4909) );
  NAND2_X1 U4532 ( .A1(n5134), .A2(n6194), .ZN(n3629) );
  OAI211_X1 U4533 ( .C1(n5541), .C2(n4909), .A(n3629), .B(n3751), .ZN(n3630)
         );
  NAND2_X1 U4534 ( .A1(n3631), .A2(n3630), .ZN(n4911) );
  INV_X1 U4535 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U4536 ( .A1(n3750), .A2(n6147), .ZN(n3638) );
  NAND2_X1 U4537 ( .A1(n3751), .A2(n3634), .ZN(n3636) );
  NAND2_X1 U4538 ( .A1(n5134), .A2(n6147), .ZN(n3635) );
  NAND3_X1 U4539 ( .A1(n3636), .A2(n5596), .A3(n3635), .ZN(n3637) );
  NOR2_X2 U4540 ( .A1(n4914), .A2(n4653), .ZN(n5005) );
  MUX2_X1 U4541 ( .A(n3702), .B(n5596), .S(EBX_REG_7__SCAN_IN), .Z(n3640) );
  NAND2_X1 U4542 ( .A1(n3493), .A2(n3756), .ZN(n3639) );
  NAND2_X1 U4543 ( .A1(n5005), .A2(n5004), .ZN(n5052) );
  INV_X1 U4544 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6126) );
  NAND2_X1 U4545 ( .A1(n3750), .A2(n6126), .ZN(n3645) );
  NAND2_X1 U4546 ( .A1(n3751), .A2(n3641), .ZN(n3643) );
  NAND2_X1 U4547 ( .A1(n5134), .A2(n6126), .ZN(n3642) );
  NAND3_X1 U4548 ( .A1(n3643), .A2(n5596), .A3(n3642), .ZN(n3644) );
  OR2_X2 U4549 ( .A1(n5052), .A2(n5051), .ZN(n5054) );
  NAND2_X1 U4550 ( .A1(n6326), .A2(n3756), .ZN(n3647) );
  MUX2_X1 U4551 ( .A(n3702), .B(n5596), .S(EBX_REG_9__SCAN_IN), .Z(n3646) );
  NAND2_X1 U4552 ( .A1(n3647), .A2(n3646), .ZN(n4924) );
  OAI21_X1 U4553 ( .B1(n5541), .B2(n6317), .A(n3751), .ZN(n3650) );
  INV_X1 U4554 ( .A(EBX_REG_10__SCAN_IN), .ZN(n3648) );
  NAND2_X1 U4555 ( .A1(n5134), .A2(n3648), .ZN(n3649) );
  NAND2_X1 U4556 ( .A1(n3650), .A2(n3649), .ZN(n3651) );
  OAI21_X1 U4557 ( .B1(EBX_REG_10__SCAN_IN), .B2(n3757), .A(n3651), .ZN(n5136)
         );
  AND2_X2 U4558 ( .A1(n5137), .A2(n5136), .ZN(n5195) );
  MUX2_X1 U4559 ( .A(n3702), .B(n5596), .S(EBX_REG_11__SCAN_IN), .Z(n3653) );
  NAND2_X1 U4560 ( .A1(n5261), .A2(n3756), .ZN(n3652) );
  INV_X1 U4561 ( .A(EBX_REG_12__SCAN_IN), .ZN(n3655) );
  NAND2_X1 U4562 ( .A1(n3750), .A2(n3655), .ZN(n3659) );
  NAND2_X1 U4563 ( .A1(n3751), .A2(n3654), .ZN(n3657) );
  NAND2_X1 U4564 ( .A1(n5134), .A2(n3655), .ZN(n3656) );
  NAND3_X1 U4565 ( .A1(n3657), .A2(n5596), .A3(n3656), .ZN(n3658) );
  AND2_X1 U4566 ( .A1(n3659), .A2(n3658), .ZN(n5223) );
  MUX2_X1 U4567 ( .A(n3702), .B(n5596), .S(EBX_REG_13__SCAN_IN), .Z(n3660) );
  OAI21_X1 U4568 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n4374), .A(n3660), 
        .ZN(n5292) );
  OAI21_X1 U4569 ( .B1(n5541), .B2(n6003), .A(n3751), .ZN(n3661) );
  OAI21_X1 U4570 ( .B1(EBX_REG_14__SCAN_IN), .B2(n4379), .A(n3661), .ZN(n3663)
         );
  INV_X1 U4571 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U4572 ( .A1(n3750), .A2(n5323), .ZN(n3662) );
  NAND2_X1 U4573 ( .A1(n4374), .A2(EBX_REG_15__SCAN_IN), .ZN(n3665) );
  NAND2_X1 U4574 ( .A1(n4379), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3664) );
  NAND2_X1 U4575 ( .A1(n3665), .A2(n3664), .ZN(n3666) );
  XNOR2_X1 U4576 ( .A(n3666), .B(n5596), .ZN(n5377) );
  OAI21_X1 U4577 ( .B1(n5541), .B2(n5992), .A(n3751), .ZN(n3667) );
  OAI21_X1 U4578 ( .B1(EBX_REG_16__SCAN_IN), .B2(n4379), .A(n3667), .ZN(n3669)
         );
  INV_X1 U4579 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5311) );
  NAND2_X1 U4580 ( .A1(n3750), .A2(n5311), .ZN(n3668) );
  AND2_X1 U4581 ( .A1(n3669), .A2(n3668), .ZN(n5308) );
  INV_X1 U4582 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6064) );
  NAND2_X1 U4583 ( .A1(n3696), .A2(n6064), .ZN(n3672) );
  INV_X1 U4584 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5850) );
  NAND2_X1 U4585 ( .A1(n5134), .A2(n6064), .ZN(n3670) );
  OAI211_X1 U4586 ( .C1(n5541), .C2(n5850), .A(n3670), .B(n3751), .ZN(n3671)
         );
  NAND2_X1 U4587 ( .A1(n3672), .A2(n3671), .ZN(n5300) );
  OAI21_X1 U4588 ( .B1(n5541), .B2(n3516), .A(n3751), .ZN(n3674) );
  INV_X1 U4589 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5600) );
  NAND2_X1 U4590 ( .A1(n5134), .A2(n5600), .ZN(n3673) );
  NAND2_X1 U4591 ( .A1(n3674), .A2(n3673), .ZN(n3675) );
  OAI21_X1 U4592 ( .B1(EBX_REG_19__SCAN_IN), .B2(n3757), .A(n3675), .ZN(n5544)
         );
  NOR2_X1 U4593 ( .A1(n4379), .A2(EBX_REG_20__SCAN_IN), .ZN(n3676) );
  AOI21_X1 U4594 ( .B1(n3756), .B2(n3677), .A(n3676), .ZN(n5597) );
  OR2_X1 U4595 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3678)
         );
  INV_X1 U4596 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U4597 ( .A1(n5134), .A2(n5609), .ZN(n5542) );
  NAND2_X1 U4598 ( .A1(n3678), .A2(n5542), .ZN(n5595) );
  NAND2_X1 U4599 ( .A1(n5541), .A2(EBX_REG_20__SCAN_IN), .ZN(n3680) );
  NAND2_X1 U4600 ( .A1(n5595), .A2(n5596), .ZN(n3679) );
  OAI211_X1 U4601 ( .C1(n5597), .C2(n5595), .A(n3680), .B(n3679), .ZN(n3681)
         );
  INV_X1 U4602 ( .A(n3681), .ZN(n3682) );
  MUX2_X1 U4603 ( .A(n3702), .B(n5596), .S(EBX_REG_21__SCAN_IN), .Z(n3683) );
  OAI21_X1 U4604 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n4374), .A(n3683), 
        .ZN(n5586) );
  INV_X1 U4605 ( .A(EBX_REG_23__SCAN_IN), .ZN(n3684) );
  MUX2_X1 U4606 ( .A(n5541), .B(n3696), .S(n3684), .Z(n3686) );
  NOR2_X1 U4607 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3685)
         );
  NOR2_X1 U4608 ( .A1(n3686), .A2(n3685), .ZN(n5575) );
  INV_X1 U4609 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5943) );
  NAND2_X1 U4610 ( .A1(n3750), .A2(n5943), .ZN(n3690) );
  INV_X1 U4611 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n6709) );
  NAND2_X1 U4612 ( .A1(n3751), .A2(n6709), .ZN(n3688) );
  NAND2_X1 U4613 ( .A1(n5134), .A2(n5943), .ZN(n3687) );
  NAND3_X1 U4614 ( .A1(n3688), .A2(n5596), .A3(n3687), .ZN(n3689) );
  NAND2_X1 U4615 ( .A1(n3690), .A2(n3689), .ZN(n5580) );
  NAND2_X1 U4616 ( .A1(n5575), .A2(n5580), .ZN(n3691) );
  NOR2_X2 U4617 ( .A1(n5588), .A2(n3691), .ZN(n5576) );
  NAND2_X1 U4618 ( .A1(n3751), .A2(n5792), .ZN(n3693) );
  INV_X1 U4619 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U4620 ( .A1(n5134), .A2(n5570), .ZN(n3692) );
  NAND3_X1 U4621 ( .A1(n3693), .A2(n5596), .A3(n3692), .ZN(n3694) );
  OAI21_X1 U4622 ( .B1(n3757), .B2(EBX_REG_24__SCAN_IN), .A(n3694), .ZN(n5567)
         );
  AND2_X2 U4623 ( .A1(n5576), .A2(n5567), .ZN(n5569) );
  INV_X1 U4624 ( .A(EBX_REG_25__SCAN_IN), .ZN(n3695) );
  MUX2_X1 U4625 ( .A(n5541), .B(n3696), .S(n3695), .Z(n3698) );
  NOR2_X1 U4626 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3697)
         );
  NOR2_X1 U4627 ( .A1(n3698), .A2(n3697), .ZN(n5529) );
  INV_X1 U4628 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5563) );
  NAND2_X1 U4629 ( .A1(n3750), .A2(n5563), .ZN(n3701) );
  NAND2_X1 U4630 ( .A1(n3751), .A2(n5776), .ZN(n3699) );
  OAI211_X1 U4631 ( .C1(EBX_REG_26__SCAN_IN), .C2(n4379), .A(n3699), .B(n5596), 
        .ZN(n3700) );
  AND2_X1 U4632 ( .A1(n3701), .A2(n3700), .ZN(n5514) );
  MUX2_X1 U4633 ( .A(n3702), .B(n5596), .S(EBX_REG_27__SCAN_IN), .Z(n3703) );
  OAI21_X1 U4634 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n4374), .A(n3703), 
        .ZN(n3704) );
  NAND2_X1 U4635 ( .A1(n5516), .A2(n3704), .ZN(n3705) );
  NAND2_X1 U4636 ( .A1(n5493), .A2(n3705), .ZN(n5561) );
  OR2_X1 U4637 ( .A1(n3580), .A2(n6591), .ZN(n6472) );
  OAI21_X1 U4638 ( .B1(n3706), .B2(n3219), .A(n6472), .ZN(n3707) );
  OAI21_X1 U4639 ( .B1(n3776), .B2(n3606), .A(n3708), .ZN(n3709) );
  NAND2_X1 U4640 ( .A1(n4528), .A2(n3600), .ZN(n5179) );
  OR2_X1 U4641 ( .A1(n5179), .A2(n3708), .ZN(n4363) );
  NAND3_X1 U4642 ( .A1(n3756), .A2(n3709), .A3(n4363), .ZN(n3711) );
  NAND2_X1 U4643 ( .A1(n3711), .A2(n3710), .ZN(n3712) );
  NAND2_X1 U4644 ( .A1(n3713), .A2(n3712), .ZN(n4350) );
  INV_X1 U4645 ( .A(n4350), .ZN(n3718) );
  OAI21_X1 U4646 ( .B1(n3715), .B2(n3714), .A(n4579), .ZN(n3716) );
  AOI21_X1 U4647 ( .B1(n5541), .B2(n4344), .A(n3716), .ZN(n3717) );
  NAND3_X1 U4648 ( .A1(n3718), .A2(n3717), .A3(n4347), .ZN(n3719) );
  NAND2_X1 U4649 ( .A1(n3722), .A2(n3719), .ZN(n3736) );
  INV_X1 U4650 ( .A(n3722), .ZN(n3720) );
  NAND2_X1 U4651 ( .A1(n3720), .A2(n6308), .ZN(n4467) );
  OAI21_X1 U4652 ( .B1(n3736), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4467), 
        .ZN(n4416) );
  INV_X1 U4653 ( .A(n4416), .ZN(n5154) );
  INV_X1 U4654 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6569) );
  OAI21_X1 U4655 ( .B1(n3607), .B2(n6569), .A(n3615), .ZN(n4899) );
  INV_X1 U4656 ( .A(n4899), .ZN(n4449) );
  NAND2_X1 U4657 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4910) );
  NOR2_X1 U4658 ( .A1(n4909), .A2(n4910), .ZN(n4902) );
  NAND2_X1 U4659 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4902), .ZN(n5150)
         );
  NOR2_X1 U4660 ( .A1(n4449), .A2(n5150), .ZN(n5156) );
  NAND2_X1 U4661 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U4662 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6314) );
  NOR2_X1 U4663 ( .A1(n6313), .A2(n6314), .ZN(n5260) );
  NAND2_X1 U4664 ( .A1(n5156), .A2(n5260), .ZN(n3735) );
  AND2_X1 U4665 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6009) );
  NAND2_X1 U4666 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6009), .ZN(n6016) );
  NOR2_X1 U4667 ( .A1(n6003), .A2(n6016), .ZN(n5987) );
  NAND3_X1 U4668 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5987), .ZN(n3734) );
  NOR2_X1 U4669 ( .A1(n6446), .A2(n4528), .ZN(n3721) );
  NAND2_X1 U4670 ( .A1(n3722), .A2(n4375), .ZN(n5155) );
  INV_X1 U4671 ( .A(n5155), .ZN(n5276) );
  OAI21_X1 U4672 ( .B1(n3735), .B2(n3734), .A(n5276), .ZN(n3724) );
  NAND2_X1 U4673 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4451) );
  NOR2_X1 U4674 ( .A1(n5150), .A2(n4451), .ZN(n5153) );
  NAND2_X1 U4675 ( .A1(n5260), .A2(n5153), .ZN(n3738) );
  NOR2_X1 U4676 ( .A1(n3594), .A2(n4535), .ZN(n6449) );
  NAND2_X1 U4677 ( .A1(n3722), .A2(n6449), .ZN(n4466) );
  NAND2_X1 U4678 ( .A1(n3736), .A2(n4466), .ZN(n5159) );
  OAI21_X1 U4679 ( .B1(n3734), .B2(n3738), .A(n5159), .ZN(n3723) );
  NAND3_X1 U4680 ( .A1(n5154), .A2(n3724), .A3(n3723), .ZN(n5979) );
  INV_X1 U4681 ( .A(n5979), .ZN(n5827) );
  INV_X1 U4682 ( .A(n5790), .ZN(n5831) );
  NAND2_X1 U4683 ( .A1(n5155), .A2(n3736), .ZN(n6331) );
  NAND2_X1 U4684 ( .A1(n6010), .A2(n4466), .ZN(n6329) );
  OAI21_X1 U4685 ( .B1(n5831), .B2(n3740), .A(n6329), .ZN(n3725) );
  AND2_X1 U4686 ( .A1(n5827), .A2(n3725), .ZN(n5817) );
  INV_X1 U4687 ( .A(n5810), .ZN(n5692) );
  NAND2_X1 U4688 ( .A1(n6329), .A2(n5692), .ZN(n3726) );
  AND2_X1 U4689 ( .A1(n5817), .A2(n3726), .ZN(n5799) );
  NAND2_X1 U4690 ( .A1(n4466), .A2(n6569), .ZN(n6328) );
  NAND2_X1 U4691 ( .A1(n5159), .A2(n6328), .ZN(n4450) );
  NAND2_X1 U4692 ( .A1(n4450), .A2(n5155), .ZN(n5825) );
  INV_X1 U4693 ( .A(n3727), .ZN(n3728) );
  NAND2_X1 U4694 ( .A1(n5825), .A2(n3728), .ZN(n3729) );
  AND2_X1 U4695 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3742) );
  INV_X1 U4696 ( .A(n3742), .ZN(n3762) );
  NAND2_X1 U4697 ( .A1(n6329), .A2(n3762), .ZN(n3730) );
  NAND2_X1 U4698 ( .A1(n5791), .A2(n3730), .ZN(n5764) );
  INV_X1 U4699 ( .A(n6308), .ZN(n6334) );
  NAND2_X1 U4700 ( .A1(n6334), .A2(REIP_REG_27__SCAN_IN), .ZN(n5436) );
  INV_X1 U4701 ( .A(n5436), .ZN(n3731) );
  AOI21_X1 U4702 ( .B1(n5764), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n3731), 
        .ZN(n3732) );
  OAI21_X1 U4703 ( .B1(n5561), .B2(n6309), .A(n3732), .ZN(n3733) );
  INV_X1 U4704 ( .A(n3733), .ZN(n3744) );
  INV_X1 U4705 ( .A(n3734), .ZN(n3739) );
  INV_X1 U4706 ( .A(n3735), .ZN(n3737) );
  NOR3_X1 U4707 ( .A1(n3736), .A2(n6569), .A3(n3738), .ZN(n5274) );
  AOI21_X1 U4708 ( .B1(n3737), .B2(n5276), .A(n5274), .ZN(n6005) );
  NOR2_X1 U4709 ( .A1(n4466), .A2(n3738), .ZN(n5275) );
  INV_X1 U4710 ( .A(n5275), .ZN(n6024) );
  NAND2_X1 U4711 ( .A1(n6005), .A2(n6024), .ZN(n6002) );
  NAND2_X1 U4712 ( .A1(n3739), .A2(n6002), .ZN(n5983) );
  INV_X1 U4713 ( .A(n5763), .ZN(n3743) );
  NAND2_X1 U4714 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5761) );
  INV_X1 U4715 ( .A(n5761), .ZN(n3746) );
  NOR2_X1 U4716 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5760) );
  NAND2_X1 U4717 ( .A1(n5652), .A2(n5760), .ZN(n5649) );
  INV_X1 U4718 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4356) );
  NAND2_X1 U4719 ( .A1(n3771), .A2(n6322), .ZN(n3769) );
  AND2_X1 U4720 ( .A1(n4379), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3748)
         );
  AOI21_X1 U4721 ( .B1(n4374), .B2(EBX_REG_30__SCAN_IN), .A(n3748), .ZN(n5417)
         );
  INV_X1 U4722 ( .A(EBX_REG_28__SCAN_IN), .ZN(n3749) );
  NAND2_X1 U4723 ( .A1(n3750), .A2(n3749), .ZN(n3754) );
  INV_X1 U4724 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5648) );
  NAND2_X1 U4725 ( .A1(n3751), .A2(n5648), .ZN(n3752) );
  OAI211_X1 U4726 ( .C1(EBX_REG_28__SCAN_IN), .C2(n4379), .A(n3752), .B(n5596), 
        .ZN(n3753) );
  AND2_X1 U4727 ( .A1(n3754), .A2(n3753), .ZN(n5492) );
  INV_X1 U4728 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5423) );
  NOR2_X1 U4729 ( .A1(n4379), .A2(EBX_REG_29__SCAN_IN), .ZN(n3755) );
  AOI21_X1 U4730 ( .B1(n3756), .B2(n5423), .A(n3755), .ZN(n5451) );
  OR2_X1 U4731 ( .A1(n5416), .A2(n5541), .ZN(n3759) );
  NOR2_X1 U4732 ( .A1(n3757), .A2(EBX_REG_29__SCAN_IN), .ZN(n5450) );
  NAND2_X1 U4733 ( .A1(n5495), .A2(n5450), .ZN(n3758) );
  NOR2_X1 U4734 ( .A1(n5418), .A2(n5541), .ZN(n5415) );
  AOI21_X1 U4735 ( .B1(n5417), .B2(n5449), .A(n5415), .ZN(n3761) );
  OAI22_X1 U4736 ( .A1(n4374), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4379), .ZN(n3760) );
  NAND2_X1 U4737 ( .A1(n5763), .A2(n3746), .ZN(n5755) );
  NAND2_X1 U4738 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3764) );
  NOR3_X1 U4739 ( .A1(n5755), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n3764), 
        .ZN(n3767) );
  OAI21_X1 U4740 ( .B1(n5761), .B2(n3762), .A(n6329), .ZN(n3763) );
  NAND2_X1 U4741 ( .A1(n5791), .A2(n3763), .ZN(n5752) );
  AOI21_X1 U4742 ( .B1(n6329), .B2(n3764), .A(n5752), .ZN(n3765) );
  NAND2_X1 U4743 ( .A1(n6334), .A2(REIP_REG_31__SCAN_IN), .ZN(n4277) );
  OAI21_X1 U4744 ( .B1(n3765), .B2(n4356), .A(n4277), .ZN(n3766) );
  AOI211_X1 U4745 ( .C1(n5553), .C2(n6333), .A(n3767), .B(n3766), .ZN(n3768)
         );
  NAND2_X1 U4746 ( .A1(n3769), .A2(n3768), .ZN(U2987) );
  NAND2_X1 U4747 ( .A1(n3771), .A2(n6289), .ZN(n4280) );
  NAND2_X1 U4748 ( .A1(n2997), .A2(EAX_REG_13__SCAN_IN), .ZN(n3774) );
  INV_X1 U4749 ( .A(n4257), .ZN(n4233) );
  OAI21_X1 U4750 ( .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n3772), .A(n3936), 
        .ZN(n6103) );
  NAND2_X1 U4751 ( .A1(n5335), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4122) );
  AOI22_X1 U4752 ( .A1(n4233), .A2(n6103), .B1(n4265), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3773) );
  NAND2_X1 U4753 ( .A1(n3774), .A2(n3773), .ZN(n3990) );
  NOR2_X2 U4754 ( .A1(n3251), .A2(n5335), .ZN(n3949) );
  INV_X1 U4755 ( .A(n3776), .ZN(n5444) );
  NAND2_X1 U4756 ( .A1(n5444), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3821) );
  NAND2_X1 U4757 ( .A1(n4723), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3778)
         );
  NAND2_X1 U4758 ( .A1(n2997), .A2(EAX_REG_4__SCAN_IN), .ZN(n3777) );
  OAI211_X1 U4759 ( .C1(n3821), .C2(n3779), .A(n3778), .B(n3777), .ZN(n3780)
         );
  NAND2_X1 U4760 ( .A1(n3780), .A2(n4257), .ZN(n3782) );
  OAI21_X1 U4761 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n3785), .A(n3797), 
        .ZN(n6179) );
  NAND2_X1 U4762 ( .A1(n4233), .A2(n6179), .ZN(n3781) );
  NAND2_X1 U4763 ( .A1(n3782), .A2(n3781), .ZN(n3783) );
  INV_X1 U4764 ( .A(n3807), .ZN(n3787) );
  INV_X1 U4765 ( .A(n3785), .ZN(n3786) );
  OAI21_X1 U4766 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3787), .A(n3786), 
        .ZN(n5234) );
  AOI22_X1 U4767 ( .A1(n4233), .A2(n5234), .B1(n4265), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3789) );
  NAND2_X1 U4768 ( .A1(n2997), .A2(EAX_REG_3__SCAN_IN), .ZN(n3788) );
  OAI211_X1 U4769 ( .C1(n3821), .C2(n3108), .A(n3789), .B(n3788), .ZN(n3790)
         );
  AOI21_X1 U4770 ( .B1(n4773), .B2(n3949), .A(n3790), .ZN(n4457) );
  INV_X1 U4771 ( .A(n3949), .ZN(n3939) );
  OR2_X1 U4772 ( .A1(n3792), .A2(n3939), .ZN(n3793) );
  OR2_X1 U4773 ( .A1(n3794), .A2(n3793), .ZN(n3796) );
  OR2_X1 U4774 ( .A1(n3939), .A2(n3048), .ZN(n3795) );
  NAND2_X1 U4775 ( .A1(n3796), .A2(n3795), .ZN(n3804) );
  INV_X1 U4776 ( .A(n3797), .ZN(n3799) );
  INV_X1 U4777 ( .A(n3828), .ZN(n3798) );
  OAI21_X1 U4778 ( .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n3799), .A(n3798), 
        .ZN(n6275) );
  NAND2_X1 U4779 ( .A1(n4233), .A2(n6275), .ZN(n3800) );
  OAI21_X1 U4780 ( .B1(n6283), .B2(n4122), .A(n3800), .ZN(n3801) );
  AOI21_X1 U4781 ( .B1(n2997), .B2(EAX_REG_5__SCAN_IN), .A(n3801), .ZN(n3802)
         );
  NAND2_X1 U4782 ( .A1(n3805), .A2(n3949), .ZN(n3806) );
  NAND2_X1 U4783 ( .A1(n3806), .A2(n4122), .ZN(n3824) );
  OAI21_X1 U4784 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3807), .ZN(n6293) );
  AOI22_X1 U4785 ( .A1(n4265), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n4233), 
        .B2(n6293), .ZN(n3809) );
  NAND2_X1 U4786 ( .A1(n2997), .A2(EAX_REG_2__SCAN_IN), .ZN(n3808) );
  OAI211_X1 U4787 ( .C1(n3821), .C2(n3107), .A(n3809), .B(n3808), .ZN(n3823)
         );
  NAND2_X1 U4788 ( .A1(n3824), .A2(n3823), .ZN(n3822) );
  AOI22_X1 U4789 ( .A1(n2997), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n4723), .ZN(n3812) );
  INV_X1 U4790 ( .A(n3821), .ZN(n3810) );
  NAND2_X1 U4791 ( .A1(n3810), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3811) );
  AND2_X1 U4792 ( .A1(n3812), .A2(n3811), .ZN(n3813) );
  NAND2_X1 U4793 ( .A1(n3814), .A2(n3813), .ZN(n4404) );
  INV_X1 U4794 ( .A(n3816), .ZN(n3817) );
  NAND2_X1 U4795 ( .A1(n3036), .A2(n3949), .ZN(n3820) );
  AOI22_X1 U4796 ( .A1(n2997), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n4723), .ZN(n3819) );
  OAI211_X1 U4797 ( .C1(n3821), .C2(n3076), .A(n3820), .B(n3819), .ZN(n4383)
         );
  MUX2_X1 U4798 ( .A(n4233), .B(n4384), .S(n4383), .Z(n4403) );
  NAND2_X1 U4799 ( .A1(n4404), .A2(n4403), .ZN(n4433) );
  NAND2_X1 U4800 ( .A1(n3822), .A2(n4433), .ZN(n3825) );
  NOR2_X1 U4801 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n3828), .ZN(n3829)
         );
  NOR2_X1 U4802 ( .A1(n3833), .A2(n3829), .ZN(n6149) );
  INV_X1 U4803 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n5059) );
  OAI22_X1 U4804 ( .A1(n6149), .A2(n4257), .B1(n4122), .B2(n5059), .ZN(n3830)
         );
  AOI21_X1 U4805 ( .B1(n2997), .B2(EAX_REG_6__SCAN_IN), .A(n3830), .ZN(n3831)
         );
  INV_X1 U4806 ( .A(EAX_REG_7__SCAN_IN), .ZN(n3838) );
  INV_X1 U4807 ( .A(n3852), .ZN(n3836) );
  INV_X1 U4808 ( .A(n3833), .ZN(n3834) );
  INV_X1 U4809 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6737) );
  NAND2_X1 U4810 ( .A1(n3834), .A2(n6737), .ZN(n3835) );
  NAND2_X1 U4811 ( .A1(n3836), .A2(n3835), .ZN(n6269) );
  AOI22_X1 U4812 ( .A1(n6269), .A2(n4233), .B1(n4265), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3837) );
  OAI21_X1 U4813 ( .B1(n3106), .B2(n3838), .A(n3837), .ZN(n3839) );
  AOI22_X1 U4814 ( .A1(n3038), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4815 ( .A1(n3037), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4816 ( .A1(n3032), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4817 ( .A1(n4183), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3842) );
  NAND4_X1 U4818 ( .A1(n3845), .A2(n3844), .A3(n3843), .A4(n3842), .ZN(n3851)
         );
  AOI22_X1 U4819 ( .A1(n4247), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3030), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4820 ( .A1(n4236), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4821 ( .A1(n3312), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4822 ( .A1(n4127), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3846) );
  NAND4_X1 U4823 ( .A1(n3849), .A2(n3848), .A3(n3847), .A4(n3846), .ZN(n3850)
         );
  OAI21_X1 U4824 ( .B1(n3851), .B2(n3850), .A(n3949), .ZN(n3855) );
  NAND2_X1 U4825 ( .A1(n2997), .A2(EAX_REG_8__SCAN_IN), .ZN(n3854) );
  XNOR2_X1 U4826 ( .A(n3852), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6128) );
  AOI22_X1 U4827 ( .A1(n6128), .A2(n4233), .B1(n4265), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3853) );
  NOR2_X2 U4828 ( .A1(n5000), .A2(n5047), .ZN(n5049) );
  XOR2_X1 U4829 ( .A(n6114), .B(n3856), .Z(n6118) );
  AOI22_X1 U4830 ( .A1(n2997), .A2(EAX_REG_9__SCAN_IN), .B1(n4265), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4831 ( .A1(n3032), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4832 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n3312), .B1(n4246), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4833 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n4245), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4834 ( .A1(n4127), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4835 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3866)
         );
  AOI22_X1 U4836 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n4236), .B1(n4244), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4837 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n3038), .B1(n3305), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4838 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n3030), .B1(n4199), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4839 ( .A1(n3028), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3861) );
  NAND4_X1 U4840 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), .ZN(n3865)
         );
  OAI21_X1 U4841 ( .B1(n3866), .B2(n3865), .A(n3949), .ZN(n3867) );
  OAI211_X1 U4842 ( .C1(n6118), .C2(n4257), .A(n3868), .B(n3867), .ZN(n4922)
         );
  NAND2_X1 U4843 ( .A1(n5049), .A2(n4922), .ZN(n4921) );
  XNOR2_X1 U4844 ( .A(n3869), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5216)
         );
  AOI22_X1 U4845 ( .A1(n4247), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4846 ( .A1(n3312), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3872) );
  AOI22_X1 U4847 ( .A1(n3305), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4848 ( .A1(n4238), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3870) );
  NAND4_X1 U4849 ( .A1(n3873), .A2(n3872), .A3(n3871), .A4(n3870), .ZN(n3879)
         );
  AOI22_X1 U4850 ( .A1(n4222), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4851 ( .A1(n3038), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3037), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3876) );
  AOI22_X1 U4852 ( .A1(n4127), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4853 ( .A1(n4239), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3874) );
  NAND4_X1 U4854 ( .A1(n3877), .A2(n3876), .A3(n3875), .A4(n3874), .ZN(n3878)
         );
  OAI21_X1 U4855 ( .B1(n3879), .B2(n3878), .A(n3949), .ZN(n3882) );
  NAND2_X1 U4856 ( .A1(n2997), .A2(EAX_REG_10__SCAN_IN), .ZN(n3881) );
  NAND2_X1 U4857 ( .A1(n4265), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3880)
         );
  NAND3_X1 U4858 ( .A1(n3882), .A2(n3881), .A3(n3880), .ZN(n3883) );
  AOI21_X1 U4859 ( .B1(n5216), .B2(n4233), .A(n3883), .ZN(n5119) );
  XOR2_X1 U4860 ( .A(n3885), .B(n3884), .Z(n6264) );
  AOI22_X1 U4861 ( .A1(n2997), .A2(EAX_REG_11__SCAN_IN), .B1(n4265), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4862 ( .A1(n3312), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4863 ( .A1(n3305), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4864 ( .A1(n3032), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4865 ( .A1(n4247), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3886) );
  NAND4_X1 U4866 ( .A1(n3889), .A2(n3888), .A3(n3887), .A4(n3886), .ZN(n3895)
         );
  AOI22_X1 U4867 ( .A1(n4127), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3030), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4868 ( .A1(n4236), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3892) );
  AOI22_X1 U4869 ( .A1(n3038), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3037), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3891) );
  AOI22_X1 U4870 ( .A1(n4183), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3890) );
  NAND4_X1 U4871 ( .A1(n3893), .A2(n3892), .A3(n3891), .A4(n3890), .ZN(n3894)
         );
  OAI21_X1 U4872 ( .B1(n3895), .B2(n3894), .A(n3949), .ZN(n3896) );
  OAI211_X1 U4873 ( .C1(n6264), .C2(n4257), .A(n3897), .B(n3896), .ZN(n3898)
         );
  INV_X1 U4874 ( .A(n3898), .ZN(n5190) );
  XNOR2_X1 U4875 ( .A(n3899), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5286)
         );
  INV_X1 U4876 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3900) );
  AOI21_X1 U4877 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n3900), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3902) );
  AND2_X1 U4878 ( .A1(n2997), .A2(EAX_REG_12__SCAN_IN), .ZN(n3901) );
  OAI22_X1 U4879 ( .A1(n5286), .A2(n4257), .B1(n3902), .B2(n3901), .ZN(n3914)
         );
  AOI22_X1 U4880 ( .A1(n3032), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4881 ( .A1(n3312), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4882 ( .A1(n3038), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4883 ( .A1(n4247), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3028), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3903) );
  NAND4_X1 U4884 ( .A1(n3906), .A2(n3905), .A3(n3904), .A4(n3903), .ZN(n3912)
         );
  AOI22_X1 U4885 ( .A1(n3030), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3910) );
  AOI22_X1 U4886 ( .A1(n3037), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4887 ( .A1(n4127), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4888 ( .A1(n2996), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3907) );
  NAND4_X1 U4889 ( .A1(n3910), .A2(n3909), .A3(n3908), .A4(n3907), .ZN(n3911)
         );
  OAI21_X1 U4890 ( .B1(n3912), .B2(n3911), .A(n3949), .ZN(n3913) );
  NAND2_X1 U4891 ( .A1(n3914), .A2(n3913), .ZN(n5220) );
  AND2_X2 U4892 ( .A1(n5191), .A2(n5220), .ZN(n3994) );
  AOI22_X1 U4893 ( .A1(n4127), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3918) );
  AOI22_X1 U4894 ( .A1(n4239), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4895 ( .A1(n3312), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4896 ( .A1(n3028), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3915) );
  NAND4_X1 U4897 ( .A1(n3918), .A2(n3917), .A3(n3916), .A4(n3915), .ZN(n3924)
         );
  AOI22_X1 U4898 ( .A1(n4222), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3922) );
  AOI22_X1 U4899 ( .A1(n3038), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4900 ( .A1(n3037), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4901 ( .A1(n4199), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3919) );
  NAND4_X1 U4902 ( .A1(n3922), .A2(n3921), .A3(n3920), .A4(n3919), .ZN(n3923)
         );
  OR2_X1 U4903 ( .A1(n3924), .A2(n3923), .ZN(n3925) );
  NAND2_X1 U4904 ( .A1(n3949), .A2(n3925), .ZN(n5266) );
  AOI22_X1 U4905 ( .A1(n4239), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4906 ( .A1(n4236), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3312), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4907 ( .A1(n3038), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3037), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4908 ( .A1(n4238), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3926) );
  NAND4_X1 U4909 ( .A1(n3929), .A2(n3928), .A3(n3927), .A4(n3926), .ZN(n3935)
         );
  AOI22_X1 U4910 ( .A1(n4246), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4911 ( .A1(n3331), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4912 ( .A1(n4222), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4913 ( .A1(n4127), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3028), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3930) );
  NAND4_X1 U4914 ( .A1(n3933), .A2(n3932), .A3(n3931), .A4(n3930), .ZN(n3934)
         );
  NOR2_X1 U4915 ( .A1(n3935), .A2(n3934), .ZN(n3940) );
  AOI21_X1 U4916 ( .B1(n6757), .B2(n3936), .A(n3956), .ZN(n6089) );
  OR2_X1 U4917 ( .A1(n6089), .A2(n4257), .ZN(n3938) );
  AOI22_X1 U4918 ( .A1(n2997), .A2(EAX_REG_14__SCAN_IN), .B1(n4265), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3937) );
  OAI211_X1 U4919 ( .C1(n3940), .C2(n3939), .A(n3938), .B(n3937), .ZN(n5317)
         );
  INV_X1 U4920 ( .A(n5317), .ZN(n3992) );
  OR2_X1 U4921 ( .A1(n5266), .A2(n3992), .ZN(n5314) );
  XNOR2_X1 U4922 ( .A(n3956), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n5748)
         );
  AOI22_X1 U4923 ( .A1(n3032), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3944) );
  AOI22_X1 U4924 ( .A1(n3312), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4925 ( .A1(n3038), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4926 ( .A1(n4246), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3941) );
  NAND4_X1 U4927 ( .A1(n3944), .A2(n3943), .A3(n3942), .A4(n3941), .ZN(n3951)
         );
  AOI22_X1 U4928 ( .A1(n4222), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4929 ( .A1(n3037), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4930 ( .A1(n3028), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3946) );
  AOI22_X1 U4931 ( .A1(n4127), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3945) );
  NAND4_X1 U4932 ( .A1(n3948), .A2(n3947), .A3(n3946), .A4(n3945), .ZN(n3950)
         );
  OAI21_X1 U4933 ( .B1(n3951), .B2(n3950), .A(n3949), .ZN(n3954) );
  NAND2_X1 U4934 ( .A1(n2997), .A2(EAX_REG_15__SCAN_IN), .ZN(n3953) );
  NAND2_X1 U4935 ( .A1(n4265), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3952)
         );
  NAND3_X1 U4936 ( .A1(n3954), .A2(n3953), .A3(n3952), .ZN(n3955) );
  AOI21_X1 U4937 ( .B1(n5748), .B2(n4233), .A(n3955), .ZN(n5374) );
  OR2_X1 U4938 ( .A1(n5314), .A2(n5374), .ZN(n5303) );
  XOR2_X1 U4939 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .B(n3973), .Z(n6076) );
  AOI22_X1 U4940 ( .A1(n3030), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4941 ( .A1(n3312), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4245), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4942 ( .A1(n4247), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3028), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3958) );
  AOI22_X1 U4943 ( .A1(n3032), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3957) );
  NAND4_X1 U4944 ( .A1(n3960), .A2(n3959), .A3(n3958), .A4(n3957), .ZN(n3966)
         );
  AOI22_X1 U4945 ( .A1(n3038), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4946 ( .A1(n3305), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4947 ( .A1(n4127), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4948 ( .A1(n4246), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3961) );
  NAND4_X1 U4949 ( .A1(n3964), .A2(n3963), .A3(n3962), .A4(n3961), .ZN(n3965)
         );
  NOR2_X1 U4950 ( .A1(n3966), .A2(n3965), .ZN(n3968) );
  AOI22_X1 U4951 ( .A1(n2997), .A2(EAX_REG_16__SCAN_IN), .B1(n4265), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3967) );
  OAI21_X1 U4952 ( .B1(n4260), .B2(n3968), .A(n3967), .ZN(n3969) );
  INV_X1 U4953 ( .A(n3969), .ZN(n3970) );
  OAI21_X1 U4954 ( .B1(n6076), .B2(n4257), .A(n3970), .ZN(n5307) );
  INV_X1 U4955 ( .A(n5307), .ZN(n3971) );
  NOR2_X2 U4956 ( .A1(n5265), .A2(n3972), .ZN(n5297) );
  XNOR2_X1 U4957 ( .A(n4013), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6066)
         );
  NAND2_X1 U4958 ( .A1(n6066), .A2(n4233), .ZN(n3989) );
  AOI22_X1 U4959 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n3038), .B1(n4222), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4960 ( .A1(n4236), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3037), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4961 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n4127), .B1(n4237), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4962 ( .A1(n4246), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3974) );
  NAND4_X1 U4963 ( .A1(n3977), .A2(n3976), .A3(n3975), .A4(n3974), .ZN(n3985)
         );
  NAND2_X1 U4964 ( .A1(n4247), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3979)
         );
  NAND2_X1 U4965 ( .A1(n3305), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3978)
         );
  AND3_X1 U4966 ( .A1(n3979), .A2(n3978), .A3(n4257), .ZN(n3983) );
  AOI22_X1 U4967 ( .A1(n4239), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3028), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4968 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n3312), .B1(n4199), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4969 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n4244), .B1(n3277), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3980) );
  NAND4_X1 U4970 ( .A1(n3983), .A2(n3982), .A3(n3981), .A4(n3980), .ZN(n3984)
         );
  NAND2_X1 U4971 ( .A1(n4260), .A2(n4257), .ZN(n4066) );
  OAI21_X1 U4972 ( .B1(n3985), .B2(n3984), .A(n4066), .ZN(n3987) );
  AOI22_X1 U4973 ( .A1(n2997), .A2(EAX_REG_17__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4723), .ZN(n3986) );
  NAND2_X1 U4974 ( .A1(n3987), .A2(n3986), .ZN(n3988) );
  NAND2_X1 U4975 ( .A1(n3989), .A2(n3988), .ZN(n5298) );
  INV_X1 U4976 ( .A(n5298), .ZN(n3995) );
  NAND2_X1 U4977 ( .A1(n5297), .A2(n3995), .ZN(n3998) );
  INV_X1 U4978 ( .A(n3990), .ZN(n3991) );
  NOR2_X1 U4979 ( .A1(n3992), .A2(n3991), .ZN(n3993) );
  NOR2_X2 U4980 ( .A1(n5315), .A2(n5374), .ZN(n5304) );
  AND2_X1 U4981 ( .A1(n5307), .A2(n3995), .ZN(n3996) );
  NAND2_X1 U4982 ( .A1(n5304), .A2(n3996), .ZN(n3997) );
  AOI22_X1 U4983 ( .A1(n3030), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4984 ( .A1(n3038), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4985 ( .A1(n3028), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4000) );
  AOI22_X1 U4986 ( .A1(n4127), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3999) );
  NAND4_X1 U4987 ( .A1(n4002), .A2(n4001), .A3(n4000), .A4(n3999), .ZN(n4008)
         );
  AOI22_X1 U4988 ( .A1(n3032), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4989 ( .A1(n4236), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U4990 ( .A1(n4245), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4991 ( .A1(n4246), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4003) );
  NAND4_X1 U4992 ( .A1(n4006), .A2(n4005), .A3(n4004), .A4(n4003), .ZN(n4007)
         );
  NOR2_X1 U4993 ( .A1(n4008), .A2(n4007), .ZN(n4012) );
  NAND2_X1 U4994 ( .A1(n4723), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4009)
         );
  NAND2_X1 U4995 ( .A1(n4257), .A2(n4009), .ZN(n4010) );
  AOI21_X1 U4996 ( .B1(n2997), .B2(EAX_REG_18__SCAN_IN), .A(n4010), .ZN(n4011)
         );
  OAI21_X1 U4997 ( .B1(n4260), .B2(n4012), .A(n4011), .ZN(n4020) );
  INV_X1 U4998 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6063) );
  INV_X1 U4999 ( .A(n4051), .ZN(n4018) );
  INV_X1 U5000 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4016) );
  INV_X1 U5001 ( .A(n4014), .ZN(n4015) );
  NAND2_X1 U5002 ( .A1(n4016), .A2(n4015), .ZN(n4017) );
  NAND2_X1 U5003 ( .A1(n4018), .A2(n4017), .ZN(n6053) );
  NAND2_X1 U5004 ( .A1(n4020), .A2(n4019), .ZN(n5601) );
  AOI22_X1 U5005 ( .A1(n3038), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U5006 ( .A1(n3032), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4024) );
  AOI22_X1 U5007 ( .A1(n3331), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U5008 ( .A1(n3311), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4022) );
  NAND4_X1 U5009 ( .A1(n4025), .A2(n4024), .A3(n4023), .A4(n4022), .ZN(n4033)
         );
  AOI22_X1 U5010 ( .A1(n4127), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U5011 ( .A1(n3030), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U5012 ( .A1(n4236), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4029) );
  NAND2_X1 U5013 ( .A1(n3037), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4027) );
  AOI21_X1 U5014 ( .B1(n3367), .B2(INSTQUEUE_REG_2__3__SCAN_IN), .A(n4233), 
        .ZN(n4026) );
  AND2_X1 U5015 ( .A1(n4027), .A2(n4026), .ZN(n4028) );
  NAND4_X1 U5016 ( .A1(n4031), .A2(n4030), .A3(n4029), .A4(n4028), .ZN(n4032)
         );
  OAI21_X1 U5017 ( .B1(n4033), .B2(n4032), .A(n4066), .ZN(n4035) );
  AOI22_X1 U5018 ( .A1(n2997), .A2(EAX_REG_19__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n4723), .ZN(n4034) );
  NAND2_X1 U5019 ( .A1(n4035), .A2(n4034), .ZN(n4037) );
  INV_X1 U5020 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5722) );
  XNOR2_X1 U5021 ( .A(n4051), .B(n5722), .ZN(n5720) );
  NAND2_X1 U5022 ( .A1(n5720), .A2(n4233), .ZN(n4036) );
  NAND2_X1 U5023 ( .A1(n4037), .A2(n4036), .ZN(n5545) );
  AOI22_X1 U5024 ( .A1(n3032), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4222), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U5025 ( .A1(n4236), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U5026 ( .A1(n3311), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3037), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U5027 ( .A1(n4127), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4038) );
  NAND4_X1 U5028 ( .A1(n4041), .A2(n4040), .A3(n4039), .A4(n4038), .ZN(n4047)
         );
  AOI22_X1 U5029 ( .A1(n3038), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U5030 ( .A1(n3305), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U5031 ( .A1(n4247), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U5032 ( .A1(n3028), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4042) );
  NAND4_X1 U5033 ( .A1(n4045), .A2(n4044), .A3(n4043), .A4(n4042), .ZN(n4046)
         );
  NOR2_X1 U5034 ( .A1(n4047), .A2(n4046), .ZN(n4048) );
  OR2_X1 U5035 ( .A1(n4260), .A2(n4048), .ZN(n4055) );
  NAND2_X1 U5036 ( .A1(n4723), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n4049)
         );
  NAND2_X1 U5037 ( .A1(n4257), .A2(n4049), .ZN(n4050) );
  AOI21_X1 U5038 ( .B1(n2997), .B2(EAX_REG_20__SCAN_IN), .A(n4050), .ZN(n4054)
         );
  OAI21_X1 U5039 ( .B1(n4052), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n4075), 
        .ZN(n5961) );
  NOR2_X1 U5040 ( .A1(n5961), .A2(n4257), .ZN(n4053) );
  AOI21_X1 U5041 ( .B1(n4055), .B2(n4054), .A(n4053), .ZN(n5590) );
  AOI22_X1 U5042 ( .A1(n4247), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U5043 ( .A1(n3038), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U5044 ( .A1(n4127), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U5045 ( .A1(n3030), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3028), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4056) );
  NAND4_X1 U5046 ( .A1(n4059), .A2(n4058), .A3(n4057), .A4(n4056), .ZN(n4068)
         );
  AOI22_X1 U5047 ( .A1(n4239), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4065) );
  AOI21_X1 U5048 ( .B1(n4238), .B2(INSTQUEUE_REG_15__5__SCAN_IN), .A(n4233), 
        .ZN(n4061) );
  NAND2_X1 U5049 ( .A1(n3037), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4060) );
  AND2_X1 U5050 ( .A1(n4061), .A2(n4060), .ZN(n4064) );
  AOI22_X1 U5051 ( .A1(n3311), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U5052 ( .A1(n4199), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4062) );
  NAND4_X1 U5053 ( .A1(n4065), .A2(n4064), .A3(n4063), .A4(n4062), .ZN(n4067)
         );
  OAI21_X1 U5054 ( .B1(n4068), .B2(n4067), .A(n4066), .ZN(n4070) );
  AOI22_X1 U5055 ( .A1(n2997), .A2(EAX_REG_21__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n4723), .ZN(n4069) );
  NAND2_X1 U5056 ( .A1(n4070), .A2(n4069), .ZN(n4072) );
  XNOR2_X1 U5057 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .B(n4075), .ZN(n5951)
         );
  NAND2_X1 U5058 ( .A1(n5951), .A2(n4233), .ZN(n4071) );
  NAND2_X1 U5059 ( .A1(n4072), .A2(n4071), .ZN(n5584) );
  NAND2_X1 U5060 ( .A1(n4074), .A2(n4073), .ZN(n5578) );
  OAI21_X1 U5061 ( .B1(n4077), .B2(PHYADDRPOINTER_REG_22__SCAN_IN), .A(n4119), 
        .ZN(n5937) );
  INV_X1 U5062 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5063 ( .A1(n4222), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4081) );
  AOI22_X1 U5064 ( .A1(n4236), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4080) );
  AOI22_X1 U5065 ( .A1(n4247), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4079) );
  AOI22_X1 U5066 ( .A1(n3035), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4183), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4078) );
  NAND4_X1 U5067 ( .A1(n4081), .A2(n4080), .A3(n4079), .A4(n4078), .ZN(n4088)
         );
  AOI22_X1 U5068 ( .A1(n3032), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U5069 ( .A1(n3038), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5070 ( .A1(n3037), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U5071 ( .A1(n3277), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4082) );
  NAND4_X1 U5072 ( .A1(n4085), .A2(n4084), .A3(n4083), .A4(n4082), .ZN(n4087)
         );
  INV_X1 U5073 ( .A(n4260), .ZN(n4086) );
  OAI21_X1 U5074 ( .B1(n4088), .B2(n4087), .A(n4086), .ZN(n4090) );
  AOI21_X1 U5075 ( .B1(PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n4723), .A(n4233), 
        .ZN(n4089) );
  OAI211_X1 U5076 ( .C1(n3106), .C2(n4091), .A(n4090), .B(n4089), .ZN(n4092)
         );
  OAI21_X1 U5077 ( .B1(n4257), .B2(n5937), .A(n4092), .ZN(n5579) );
  XNOR2_X1 U5078 ( .A(n4119), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5928)
         );
  INV_X1 U5079 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5936) );
  OAI21_X1 U5080 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5936), .A(n4257), .ZN(
        n4117) );
  AOI22_X1 U5081 ( .A1(n4236), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n4096) );
  INV_X1 U5082 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6772) );
  AOI22_X1 U5083 ( .A1(n3312), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n4095) );
  AOI22_X1 U5084 ( .A1(n3038), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4094) );
  AOI22_X1 U5085 ( .A1(n3037), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4093) );
  NAND4_X1 U5086 ( .A1(n4096), .A2(n4095), .A3(n4094), .A4(n4093), .ZN(n4102)
         );
  AOI22_X1 U5087 ( .A1(n3032), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U5088 ( .A1(n3035), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4099) );
  AOI22_X1 U5089 ( .A1(n3030), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4098) );
  AOI22_X1 U5090 ( .A1(n3028), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4097) );
  NAND4_X1 U5091 ( .A1(n4100), .A2(n4099), .A3(n4098), .A4(n4097), .ZN(n4101)
         );
  OR2_X1 U5092 ( .A1(n4102), .A2(n4101), .ZN(n4135) );
  INV_X1 U5093 ( .A(n4135), .ZN(n4114) );
  AOI22_X1 U5094 ( .A1(n4236), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4106) );
  AOI22_X1 U5095 ( .A1(n3312), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5096 ( .A1(n3038), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5097 ( .A1(n4245), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4103) );
  NAND4_X1 U5098 ( .A1(n4106), .A2(n4105), .A3(n4104), .A4(n4103), .ZN(n4112)
         );
  AOI22_X1 U5099 ( .A1(n3032), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U5100 ( .A1(n3034), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5101 ( .A1(n3030), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4108) );
  AOI22_X1 U5102 ( .A1(n4183), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4107) );
  NAND4_X1 U5103 ( .A1(n4110), .A2(n4109), .A3(n4108), .A4(n4107), .ZN(n4111)
         );
  OR2_X1 U5104 ( .A1(n4112), .A2(n4111), .ZN(n4134) );
  INV_X1 U5105 ( .A(n4134), .ZN(n4113) );
  XNOR2_X1 U5106 ( .A(n4114), .B(n4113), .ZN(n4115) );
  NOR2_X1 U5107 ( .A1(n4260), .A2(n4115), .ZN(n4116) );
  AOI211_X1 U5108 ( .C1(n2997), .C2(EAX_REG_23__SCAN_IN), .A(n4117), .B(n4116), 
        .ZN(n4118) );
  AOI21_X1 U5109 ( .B1(n4233), .B2(n5928), .A(n4118), .ZN(n5574) );
  INV_X1 U5110 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5687) );
  INV_X1 U5111 ( .A(n4120), .ZN(n4121) );
  AOI21_X1 U5112 ( .B1(n5687), .B2(n4121), .A(n4157), .ZN(n5919) );
  OAI22_X1 U5113 ( .A1(n5919), .A2(n4257), .B1(n4122), .B2(n5687), .ZN(n4138)
         );
  AOI22_X1 U5114 ( .A1(n4236), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4126) );
  AOI22_X1 U5115 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4244), .B1(n3312), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4125) );
  AOI22_X1 U5116 ( .A1(n3038), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4124) );
  AOI22_X1 U5117 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(n3037), .B1(n4237), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4123) );
  NAND4_X1 U5118 ( .A1(n4126), .A2(n4125), .A3(n4124), .A4(n4123), .ZN(n4133)
         );
  AOI22_X1 U5119 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n4239), .B1(n4247), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5120 ( .A1(n4127), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4130) );
  AOI22_X1 U5121 ( .A1(n4222), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4129) );
  AOI22_X1 U5122 ( .A1(n3028), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4128) );
  NAND4_X1 U5123 ( .A1(n4131), .A2(n4130), .A3(n4129), .A4(n4128), .ZN(n4132)
         );
  NOR2_X1 U5124 ( .A1(n4133), .A2(n4132), .ZN(n4152) );
  NAND2_X1 U5125 ( .A1(n4135), .A2(n4134), .ZN(n4151) );
  XNOR2_X1 U5126 ( .A(n4152), .B(n4151), .ZN(n4136) );
  NOR2_X1 U5127 ( .A1(n4260), .A2(n4136), .ZN(n4137) );
  INV_X1 U5128 ( .A(n4157), .ZN(n4139) );
  XNOR2_X1 U5129 ( .A(n4139), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5672)
         );
  INV_X1 U5130 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5670) );
  AOI21_X1 U5131 ( .B1(n5670), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4155) );
  AOI22_X1 U5132 ( .A1(n4236), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n4144) );
  AOI22_X1 U5133 ( .A1(n3312), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n4143) );
  AOI22_X1 U5134 ( .A1(n3038), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U5135 ( .A1(n3037), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4141) );
  NAND4_X1 U5136 ( .A1(n4144), .A2(n4143), .A3(n4142), .A4(n4141), .ZN(n4150)
         );
  AOI22_X1 U5137 ( .A1(n3032), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4148) );
  AOI22_X1 U5138 ( .A1(n3034), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4147) );
  AOI22_X1 U5139 ( .A1(n3030), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4146) );
  AOI22_X1 U5140 ( .A1(n4183), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4145) );
  NAND4_X1 U5141 ( .A1(n4148), .A2(n4147), .A3(n4146), .A4(n4145), .ZN(n4149)
         );
  OR2_X1 U5142 ( .A1(n4150), .A2(n4149), .ZN(n4171) );
  NOR2_X1 U5143 ( .A1(n4152), .A2(n4151), .ZN(n4172) );
  XNOR2_X1 U5144 ( .A(n4171), .B(n4172), .ZN(n4153) );
  NOR2_X1 U5145 ( .A1(n4260), .A2(n4153), .ZN(n4154) );
  AOI211_X1 U5146 ( .C1(n2997), .C2(EAX_REG_25__SCAN_IN), .A(n4155), .B(n4154), 
        .ZN(n4156) );
  AOI21_X1 U5147 ( .B1(n4233), .B2(n5672), .A(n4156), .ZN(n5527) );
  INV_X1 U5148 ( .A(n4158), .ZN(n4159) );
  INV_X1 U5149 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5513) );
  NAND2_X1 U5150 ( .A1(n4159), .A2(n5513), .ZN(n4160) );
  NAND2_X1 U5151 ( .A1(n4194), .A2(n4160), .ZN(n5666) );
  AOI22_X1 U5152 ( .A1(n4239), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4164) );
  AOI22_X1 U5153 ( .A1(n4236), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4163) );
  AOI22_X1 U5154 ( .A1(n3312), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3037), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4162) );
  AOI22_X1 U5155 ( .A1(n3028), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4161) );
  NAND4_X1 U5156 ( .A1(n4164), .A2(n4163), .A3(n4162), .A4(n4161), .ZN(n4170)
         );
  AOI22_X1 U5157 ( .A1(n3038), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3030), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4168) );
  AOI22_X1 U5158 ( .A1(n3305), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4167) );
  AOI22_X1 U5159 ( .A1(n4247), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4166) );
  AOI22_X1 U5160 ( .A1(n3035), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4165) );
  NAND4_X1 U5161 ( .A1(n4168), .A2(n4167), .A3(n4166), .A4(n4165), .ZN(n4169)
         );
  NOR2_X1 U5162 ( .A1(n4170), .A2(n4169), .ZN(n4178) );
  NAND2_X1 U5163 ( .A1(n4172), .A2(n4171), .ZN(n4177) );
  XNOR2_X1 U5164 ( .A(n4178), .B(n4177), .ZN(n4175) );
  AOI21_X1 U5165 ( .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n4723), .A(n4233), 
        .ZN(n4174) );
  NAND2_X1 U5166 ( .A1(n2997), .A2(EAX_REG_26__SCAN_IN), .ZN(n4173) );
  OAI211_X1 U5167 ( .C1(n4175), .C2(n4260), .A(n4174), .B(n4173), .ZN(n4176)
         );
  OAI21_X1 U5168 ( .B1(n4257), .B2(n5666), .A(n4176), .ZN(n5512) );
  XNOR2_X1 U5169 ( .A(n4194), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5504)
         );
  INV_X1 U5170 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5437) );
  OAI21_X1 U5171 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5437), .A(n4257), .ZN(
        n4192) );
  NOR2_X1 U5172 ( .A1(n4178), .A2(n4177), .ZN(n4211) );
  AOI22_X1 U5173 ( .A1(n4236), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4182) );
  AOI22_X1 U5174 ( .A1(n3311), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n4181) );
  AOI22_X1 U5175 ( .A1(n3038), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4180) );
  AOI22_X1 U5176 ( .A1(n4245), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4179) );
  NAND4_X1 U5177 ( .A1(n4182), .A2(n4181), .A3(n4180), .A4(n4179), .ZN(n4189)
         );
  AOI22_X1 U5178 ( .A1(n3032), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4187) );
  AOI22_X1 U5179 ( .A1(n3034), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4186) );
  AOI22_X1 U5180 ( .A1(n3030), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4185) );
  AOI22_X1 U5181 ( .A1(n4183), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3332), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4184) );
  NAND4_X1 U5182 ( .A1(n4187), .A2(n4186), .A3(n4185), .A4(n4184), .ZN(n4188)
         );
  OR2_X1 U5183 ( .A1(n4189), .A2(n4188), .ZN(n4210) );
  XNOR2_X1 U5184 ( .A(n4211), .B(n4210), .ZN(n4190) );
  NOR2_X1 U5185 ( .A1(n4190), .A2(n4260), .ZN(n4191) );
  AOI211_X1 U5186 ( .C1(n2997), .C2(EAX_REG_27__SCAN_IN), .A(n4192), .B(n4191), 
        .ZN(n4193) );
  AOI21_X1 U5187 ( .B1(n4233), .B2(n5504), .A(n4193), .ZN(n5439) );
  INV_X1 U5188 ( .A(n4194), .ZN(n4195) );
  INV_X1 U5189 ( .A(n4196), .ZN(n4197) );
  INV_X1 U5190 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U5191 ( .A1(n4197), .A2(n5496), .ZN(n4198) );
  NAND2_X1 U5192 ( .A1(n4262), .A2(n4198), .ZN(n5656) );
  AOI22_X1 U5193 ( .A1(n3034), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3032), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4203) );
  AOI22_X1 U5194 ( .A1(n4246), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4140), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4202) );
  AOI22_X1 U5195 ( .A1(n4222), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4199), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4201) );
  AOI22_X1 U5196 ( .A1(n4183), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4200) );
  NAND4_X1 U5197 ( .A1(n4203), .A2(n4202), .A3(n4201), .A4(n4200), .ZN(n4209)
         );
  AOI22_X1 U5198 ( .A1(n4236), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4207) );
  AOI22_X1 U5199 ( .A1(n3038), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3311), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4206) );
  AOI22_X1 U5200 ( .A1(n3037), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4205) );
  AOI22_X1 U5201 ( .A1(n4247), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4204) );
  NAND4_X1 U5202 ( .A1(n4207), .A2(n4206), .A3(n4205), .A4(n4204), .ZN(n4208)
         );
  NOR2_X1 U5203 ( .A1(n4209), .A2(n4208), .ZN(n4217) );
  NAND2_X1 U5204 ( .A1(n4211), .A2(n4210), .ZN(n4216) );
  XNOR2_X1 U5205 ( .A(n4217), .B(n4216), .ZN(n4214) );
  AOI21_X1 U5206 ( .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n4723), .A(n4233), 
        .ZN(n4213) );
  NAND2_X1 U5207 ( .A1(n2997), .A2(EAX_REG_28__SCAN_IN), .ZN(n4212) );
  OAI211_X1 U5208 ( .C1(n4214), .C2(n4260), .A(n4213), .B(n4212), .ZN(n4215)
         );
  OAI21_X1 U5209 ( .B1(n4257), .B2(n5656), .A(n4215), .ZN(n5491) );
  XNOR2_X1 U5210 ( .A(n4262), .B(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5482)
         );
  INV_X1 U5211 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5484) );
  AOI21_X1 U5212 ( .B1(n5484), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4231) );
  NOR2_X1 U5213 ( .A1(n4217), .A2(n4216), .ZN(n4235) );
  AOI22_X1 U5214 ( .A1(n4236), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4246), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4221) );
  AOI22_X1 U5215 ( .A1(n3311), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U5216 ( .A1(n3038), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3331), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4219) );
  AOI22_X1 U5217 ( .A1(n4245), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4218) );
  NAND4_X1 U5218 ( .A1(n4221), .A2(n4220), .A3(n4219), .A4(n4218), .ZN(n4228)
         );
  AOI22_X1 U5219 ( .A1(n3032), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4247), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4226) );
  AOI22_X1 U5220 ( .A1(n3035), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3277), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4225) );
  AOI22_X1 U5221 ( .A1(n3030), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4224) );
  AOI22_X1 U5222 ( .A1(n3028), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4223) );
  NAND4_X1 U5223 ( .A1(n4226), .A2(n4225), .A3(n4224), .A4(n4223), .ZN(n4227)
         );
  OR2_X1 U5224 ( .A1(n4228), .A2(n4227), .ZN(n4234) );
  XNOR2_X1 U5225 ( .A(n4235), .B(n4234), .ZN(n4229) );
  NOR2_X1 U5226 ( .A1(n4229), .A2(n4260), .ZN(n4230) );
  AOI211_X1 U5227 ( .C1(n2997), .C2(EAX_REG_29__SCAN_IN), .A(n4231), .B(n4230), 
        .ZN(n4232) );
  AOI21_X1 U5228 ( .B1(n4233), .B2(n5482), .A(n4232), .ZN(n4283) );
  NAND2_X1 U5229 ( .A1(n4235), .A2(n4234), .ZN(n4255) );
  AOI22_X1 U5230 ( .A1(n3029), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4236), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4243) );
  AOI22_X1 U5231 ( .A1(n3312), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4237), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4242) );
  AOI22_X1 U5232 ( .A1(n3034), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4241) );
  AOI22_X1 U5233 ( .A1(n4239), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4240) );
  NAND4_X1 U5234 ( .A1(n4243), .A2(n4242), .A3(n4241), .A4(n4240), .ZN(n4253)
         );
  AOI22_X1 U5235 ( .A1(n3038), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4244), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4251) );
  AOI22_X1 U5236 ( .A1(n3037), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4250) );
  AOI22_X1 U5237 ( .A1(n4246), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n2996), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4249) );
  AOI22_X1 U5238 ( .A1(n4247), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3367), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4248) );
  NAND4_X1 U5239 ( .A1(n4251), .A2(n4250), .A3(n4249), .A4(n4248), .ZN(n4252)
         );
  NOR2_X1 U5240 ( .A1(n4253), .A2(n4252), .ZN(n4254) );
  XNOR2_X1 U5241 ( .A(n4255), .B(n4254), .ZN(n4261) );
  NAND2_X1 U5242 ( .A1(n5335), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4256)
         );
  NAND2_X1 U5243 ( .A1(n4257), .A2(n4256), .ZN(n4258) );
  AOI21_X1 U5244 ( .B1(n2997), .B2(EAX_REG_30__SCAN_IN), .A(n4258), .ZN(n4259)
         );
  OAI21_X1 U5245 ( .B1(n4261), .B2(n4260), .A(n4259), .ZN(n4264) );
  XNOR2_X1 U5246 ( .A(n4273), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5474)
         );
  NAND2_X1 U5247 ( .A1(n5474), .A2(n4233), .ZN(n4263) );
  NAND2_X1 U5248 ( .A1(n4264), .A2(n4263), .ZN(n5429) );
  AOI22_X1 U5249 ( .A1(n2997), .A2(EAX_REG_31__SCAN_IN), .B1(n4265), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4266) );
  XNOR2_X1 U5250 ( .A(n4267), .B(n4266), .ZN(n5615) );
  NAND3_X1 U5251 ( .A1(n6479), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6493) );
  INV_X1 U5252 ( .A(n6493), .ZN(n4268) );
  NOR2_X2 U5253 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_3__SCAN_IN), .ZN(
        n6350) );
  INV_X1 U5254 ( .A(n6350), .ZN(n6347) );
  NAND2_X1 U5255 ( .A1(n6347), .A2(n4269), .ZN(n6587) );
  NAND2_X1 U5256 ( .A1(n6587), .A2(n6479), .ZN(n4270) );
  NAND2_X1 U5257 ( .A1(n6479), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4272) );
  INV_X1 U5258 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6760) );
  NAND2_X1 U5259 ( .A1(n6760), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4271) );
  NAND2_X1 U5260 ( .A1(n4272), .A2(n4271), .ZN(n6299) );
  INV_X1 U5261 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5432) );
  INV_X1 U5262 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4274) );
  NAND2_X1 U5263 ( .A1(n6300), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4276)
         );
  OAI211_X1 U5264 ( .C1(n6294), .C2(n5132), .A(n4277), .B(n4276), .ZN(n4278)
         );
  AOI21_X1 U5265 ( .B1(n5615), .B2(n6287), .A(n4278), .ZN(n4279) );
  NAND2_X1 U5266 ( .A1(n4280), .A2(n4279), .ZN(U2955) );
  INV_X1 U5267 ( .A(n5649), .ZN(n5413) );
  AOI21_X1 U5268 ( .B1(n3746), .B2(n3747), .A(n5413), .ZN(n4281) );
  XNOR2_X1 U5269 ( .A(n4281), .B(n5423), .ZN(n5759) );
  NAND2_X1 U5270 ( .A1(n6334), .A2(REIP_REG_29__SCAN_IN), .ZN(n5753) );
  OAI21_X1 U5271 ( .B1(n6282), .B2(n5484), .A(n5753), .ZN(n4285) );
  OR2_X1 U5272 ( .A1(n3594), .A2(n4287), .ZN(n4292) );
  NOR2_X1 U5273 ( .A1(n4292), .A2(n6486), .ZN(n4302) );
  INV_X1 U5274 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n4291) );
  INV_X1 U5275 ( .A(n4308), .ZN(n4290) );
  NAND2_X1 U5276 ( .A1(n6350), .A2(n6474), .ZN(n6033) );
  OAI211_X1 U5277 ( .C1(n4302), .C2(n4291), .A(n4290), .B(n6033), .ZN(U2788)
         );
  INV_X1 U5278 ( .A(n3543), .ZN(n4422) );
  AOI22_X1 U5279 ( .A1(n6481), .A2(n4422), .B1(n4288), .B2(n4292), .ZN(n6030)
         );
  INV_X1 U5280 ( .A(n5179), .ZN(n4293) );
  NOR2_X1 U5281 ( .A1(n4293), .A2(n5139), .ZN(n4304) );
  INV_X1 U5282 ( .A(n6501), .ZN(n4387) );
  OAI21_X1 U5283 ( .B1(n4304), .B2(n4387), .A(n4307), .ZN(n6589) );
  AND2_X1 U5284 ( .A1(n6030), .A2(n6589), .ZN(n6462) );
  NOR2_X1 U5285 ( .A1(n6462), .A2(n6486), .ZN(n6038) );
  INV_X1 U5286 ( .A(MORE_REG_SCAN_IN), .ZN(n4301) );
  NAND3_X1 U5287 ( .A1(n6464), .A2(n4565), .A3(n4288), .ZN(n4296) );
  NOR2_X1 U5288 ( .A1(n3594), .A2(n4294), .ZN(n4295) );
  AOI21_X1 U5289 ( .B1(n6481), .B2(n4296), .A(n4295), .ZN(n4298) );
  INV_X1 U5290 ( .A(n4375), .ZN(n4566) );
  OR2_X1 U5291 ( .A1(n6481), .A2(n4566), .ZN(n4297) );
  AND2_X1 U5292 ( .A1(n4298), .A2(n4297), .ZN(n6465) );
  INV_X1 U5293 ( .A(n6465), .ZN(n4299) );
  NAND2_X1 U5294 ( .A1(n6038), .A2(n4299), .ZN(n4300) );
  OAI21_X1 U5295 ( .B1(n6038), .B2(n4301), .A(n4300), .ZN(U3471) );
  INV_X1 U5296 ( .A(n6033), .ZN(n4303) );
  NOR2_X1 U5297 ( .A1(n4303), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4306) );
  NAND2_X1 U5298 ( .A1(n6586), .A2(n4304), .ZN(n4305) );
  OAI21_X1 U5299 ( .B1(n6586), .B2(n4306), .A(n4305), .ZN(U3474) );
  NAND2_X1 U5300 ( .A1(n4308), .A2(n4307), .ZN(n4310) );
  INV_X1 U5301 ( .A(n6472), .ZN(n4309) );
  NAND2_X1 U5302 ( .A1(n4385), .A2(n4309), .ZN(n6262) );
  AND2_X2 U5303 ( .A1(n4310), .A2(n6262), .ZN(n6259) );
  INV_X2 U5304 ( .A(n6262), .ZN(n6256) );
  AOI22_X1 U5305 ( .A1(n6259), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n6256), .ZN(n4311) );
  INV_X1 U5306 ( .A(DATAI_5_), .ZN(n4548) );
  OR2_X1 U5307 ( .A1(n4428), .A2(n4548), .ZN(n4312) );
  NAND2_X1 U5308 ( .A1(n4311), .A2(n4312), .ZN(U2944) );
  AOI22_X1 U5309 ( .A1(n6259), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n6256), .ZN(n4313) );
  NAND2_X1 U5310 ( .A1(n4313), .A2(n4312), .ZN(U2929) );
  AOI22_X1 U5311 ( .A1(n6259), .A2(UWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_16__SCAN_IN), .B2(n6256), .ZN(n4314) );
  NAND2_X1 U5312 ( .A1(n6260), .A2(DATAI_0_), .ZN(n4319) );
  NAND2_X1 U5313 ( .A1(n4314), .A2(n4319), .ZN(U2924) );
  AOI22_X1 U5314 ( .A1(n6259), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n6256), .ZN(n4315) );
  NAND2_X1 U5315 ( .A1(n6260), .A2(DATAI_4_), .ZN(n4337) );
  NAND2_X1 U5316 ( .A1(n4315), .A2(n4337), .ZN(U2943) );
  AOI22_X1 U5317 ( .A1(n6259), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n6256), .ZN(n4316) );
  NAND2_X1 U5318 ( .A1(n6260), .A2(DATAI_7_), .ZN(n4333) );
  NAND2_X1 U5319 ( .A1(n4316), .A2(n4333), .ZN(U2946) );
  AOI22_X1 U5320 ( .A1(n6259), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n6256), .ZN(n4317) );
  NAND2_X1 U5321 ( .A1(n6260), .A2(DATAI_12_), .ZN(n4321) );
  NAND2_X1 U5322 ( .A1(n4317), .A2(n4321), .ZN(U2951) );
  AOI22_X1 U5323 ( .A1(n6259), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n6256), .ZN(n4318) );
  NAND2_X1 U5324 ( .A1(n6260), .A2(DATAI_1_), .ZN(n4326) );
  NAND2_X1 U5325 ( .A1(n4318), .A2(n4326), .ZN(U2940) );
  AOI22_X1 U5326 ( .A1(n6259), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n6256), .ZN(n4320) );
  NAND2_X1 U5327 ( .A1(n4320), .A2(n4319), .ZN(U2939) );
  AOI22_X1 U5328 ( .A1(n6259), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n6256), .ZN(n4322) );
  NAND2_X1 U5329 ( .A1(n4322), .A2(n4321), .ZN(U2936) );
  AOI22_X1 U5330 ( .A1(n6259), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n6256), .ZN(n4323) );
  NAND2_X1 U5331 ( .A1(n6260), .A2(DATAI_6_), .ZN(n4328) );
  NAND2_X1 U5332 ( .A1(n4323), .A2(n4328), .ZN(U2945) );
  AOI22_X1 U5333 ( .A1(n6259), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n6256), .ZN(n4324) );
  NAND2_X1 U5334 ( .A1(n6260), .A2(DATAI_3_), .ZN(n4330) );
  NAND2_X1 U5335 ( .A1(n4324), .A2(n4330), .ZN(U2927) );
  AOI22_X1 U5336 ( .A1(n6259), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n6256), .ZN(n4325) );
  NAND2_X1 U5337 ( .A1(n6260), .A2(DATAI_2_), .ZN(n4339) );
  NAND2_X1 U5338 ( .A1(n4325), .A2(n4339), .ZN(U2926) );
  AOI22_X1 U5339 ( .A1(n6259), .A2(UWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_17__SCAN_IN), .B2(n6256), .ZN(n4327) );
  NAND2_X1 U5340 ( .A1(n4327), .A2(n4326), .ZN(U2925) );
  AOI22_X1 U5341 ( .A1(n6259), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n6256), .ZN(n4329) );
  NAND2_X1 U5342 ( .A1(n4329), .A2(n4328), .ZN(U2930) );
  AOI22_X1 U5343 ( .A1(n6259), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n6256), .ZN(n4331) );
  NAND2_X1 U5344 ( .A1(n4331), .A2(n4330), .ZN(U2942) );
  AOI22_X1 U5345 ( .A1(n6259), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n6256), .ZN(n4332) );
  NAND2_X1 U5346 ( .A1(n6260), .A2(DATAI_14_), .ZN(n4335) );
  NAND2_X1 U5347 ( .A1(n4332), .A2(n4335), .ZN(U2953) );
  AOI22_X1 U5348 ( .A1(n6259), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n6256), .ZN(n4334) );
  NAND2_X1 U5349 ( .A1(n4334), .A2(n4333), .ZN(U2931) );
  AOI22_X1 U5350 ( .A1(n6259), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n6256), .ZN(n4336) );
  NAND2_X1 U5351 ( .A1(n4336), .A2(n4335), .ZN(U2938) );
  AOI22_X1 U5352 ( .A1(n6259), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n6256), .ZN(n4338) );
  NAND2_X1 U5353 ( .A1(n4338), .A2(n4337), .ZN(U2928) );
  AOI22_X1 U5354 ( .A1(n6259), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n6256), .ZN(n4340) );
  NAND2_X1 U5355 ( .A1(n4340), .A2(n4339), .ZN(U2941) );
  OAI21_X1 U5356 ( .B1(n4344), .B2(n4343), .A(n5541), .ZN(n4345) );
  AND4_X1 U5357 ( .A1(n4347), .A2(n3580), .A3(n4346), .A4(n4345), .ZN(n4348)
         );
  NAND2_X1 U5358 ( .A1(n4348), .A2(n2999), .ZN(n4349) );
  NOR2_X1 U5359 ( .A1(n4350), .A2(n4349), .ZN(n4571) );
  NOR3_X1 U5360 ( .A1(n6446), .A2(n4351), .A3(n4352), .ZN(n4353) );
  AOI21_X1 U5361 ( .B1(n6449), .B2(n4354), .A(n4353), .ZN(n4355) );
  OAI21_X1 U5362 ( .B1(n4342), .B2(n4571), .A(n4355), .ZN(n6451) );
  INV_X1 U5363 ( .A(n6575), .ZN(n5407) );
  NOR2_X1 U5364 ( .A1(n6474), .A2(n6569), .ZN(n5401) );
  AOI22_X1 U5365 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4356), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3607), .ZN(n5402) );
  AOI222_X1 U5366 ( .A1(n6451), .A2(n5407), .B1(n5401), .B2(n5402), .C1(n4357), 
        .C2(n5400), .ZN(n4372) );
  INV_X1 U5367 ( .A(n4358), .ZN(n4370) );
  NOR2_X1 U5368 ( .A1(n5134), .A2(n4387), .ZN(n4360) );
  NAND2_X1 U5369 ( .A1(n6449), .A2(n4387), .ZN(n4359) );
  OAI21_X1 U5370 ( .B1(n4360), .B2(n3580), .A(n4359), .ZN(n4361) );
  NAND2_X1 U5371 ( .A1(n4361), .A2(n4307), .ZN(n4364) );
  OAI211_X1 U5372 ( .C1(n6481), .C2(n4364), .A(n4363), .B(n4362), .ZN(n4369)
         );
  OR2_X1 U5373 ( .A1(n6481), .A2(n4565), .ZN(n4368) );
  INV_X1 U5374 ( .A(n2999), .ZN(n4366) );
  NAND2_X1 U5375 ( .A1(n4366), .A2(n4365), .ZN(n4367) );
  NAND2_X1 U5376 ( .A1(n4368), .A2(n4367), .ZN(n4426) );
  NOR3_X1 U5377 ( .A1(n4370), .A2(n4369), .A3(n4426), .ZN(n4584) );
  INV_X1 U5378 ( .A(n4584), .ZN(n6450) );
  NAND2_X1 U5379 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4596) );
  NOR2_X1 U5380 ( .A1(n6479), .A2(n4596), .ZN(n4594) );
  AOI22_X1 U5381 ( .A1(n6450), .A2(n4424), .B1(FLUSH_REG_SCAN_IN), .B2(n4594), 
        .ZN(n6027) );
  NAND2_X1 U5382 ( .A1(n6479), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U5383 ( .A1(n6027), .A2(n6565), .ZN(n6573) );
  INV_X1 U5384 ( .A(n6573), .ZN(n5409) );
  INV_X1 U5385 ( .A(n5400), .ZN(n5865) );
  NOR2_X1 U5386 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n5865), .ZN(n6568)
         );
  OAI21_X1 U5387 ( .B1(n5409), .B2(n6568), .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), 
        .ZN(n4371) );
  OAI21_X1 U5388 ( .B1(n4372), .B2(n5409), .A(n4371), .ZN(U3460) );
  OAI21_X1 U5389 ( .B1(n4374), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4373), 
        .ZN(n5206) );
  NAND2_X1 U5390 ( .A1(n6481), .A2(n4375), .ZN(n4381) );
  INV_X1 U5391 ( .A(n4376), .ZN(n4377) );
  NAND4_X1 U5392 ( .A1(n4378), .A2(n4377), .A3(n3270), .A4(n5612), .ZN(n4423)
         );
  OR2_X1 U5393 ( .A1(n4423), .A2(n4379), .ZN(n4380) );
  NAND2_X1 U5394 ( .A1(n4381), .A2(n4380), .ZN(n4382) );
  INV_X1 U5395 ( .A(EBX_REG_0__SCAN_IN), .ZN(n5202) );
  AND2_X1 U5396 ( .A1(n6195), .A2(n5445), .ZN(n6192) );
  INV_X2 U5397 ( .A(n6192), .ZN(n5610) );
  XNOR2_X1 U5398 ( .A(n4384), .B(n4383), .ZN(n6304) );
  OAI222_X1 U5399 ( .A1(n5206), .A2(n5608), .B1(n5202), .B2(n6195), .C1(n5610), 
        .C2(n6304), .ZN(U2859) );
  INV_X1 U5400 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4390) );
  NAND2_X1 U5401 ( .A1(n4385), .A2(n6449), .ZN(n4386) );
  NAND2_X1 U5402 ( .A1(n6262), .A2(n4386), .ZN(n4388) );
  NAND2_X1 U5403 ( .A1(n6209), .A2(n3606), .ZN(n4484) );
  AOI22_X1 U5404 ( .A1(UWORD_REG_14__SCAN_IN), .A2(n6588), .B1(n6238), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4389) );
  OAI21_X1 U5405 ( .B1(n4390), .B2(n4484), .A(n4389), .ZN(U2893) );
  INV_X1 U5406 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4392) );
  AOI22_X1 U5407 ( .A1(UWORD_REG_10__SCAN_IN), .A2(n6588), .B1(n6238), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4391) );
  OAI21_X1 U5408 ( .B1(n4392), .B2(n4484), .A(n4391), .ZN(U2897) );
  INV_X1 U5409 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4394) );
  AOI22_X1 U5410 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n6588), .B1(n6238), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4393) );
  OAI21_X1 U5411 ( .B1(n4394), .B2(n4484), .A(n4393), .ZN(U2896) );
  INV_X1 U5412 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4396) );
  AOI22_X1 U5413 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n6588), .B1(n6238), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4395) );
  OAI21_X1 U5414 ( .B1(n4396), .B2(n4484), .A(n4395), .ZN(U2895) );
  INV_X1 U5415 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4398) );
  AOI22_X1 U5416 ( .A1(UWORD_REG_13__SCAN_IN), .A2(n6588), .B1(n6238), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4397) );
  OAI21_X1 U5417 ( .B1(n4398), .B2(n4484), .A(n4397), .ZN(U2894) );
  INV_X1 U5418 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4400) );
  AOI22_X1 U5419 ( .A1(UWORD_REG_8__SCAN_IN), .A2(n6588), .B1(n6238), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4399) );
  OAI21_X1 U5420 ( .B1(n4400), .B2(n4484), .A(n4399), .ZN(U2899) );
  INV_X1 U5421 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4402) );
  AOI22_X1 U5422 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n6588), .B1(n6238), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4401) );
  OAI21_X1 U5423 ( .B1(n4402), .B2(n4484), .A(n4401), .ZN(U2898) );
  OR2_X1 U5424 ( .A1(n4404), .A2(n4403), .ZN(n4405) );
  NAND2_X1 U5425 ( .A1(n4405), .A2(n4433), .ZN(n5246) );
  XNOR2_X1 U5426 ( .A(n5250), .B(n5134), .ZN(n6332) );
  AOI22_X1 U5427 ( .A1(n6191), .A2(n6332), .B1(EBX_REG_1__SCAN_IN), .B2(n5559), 
        .ZN(n4406) );
  OAI21_X1 U5428 ( .B1(n5610), .B2(n5246), .A(n4406), .ZN(U2858) );
  NAND2_X1 U5429 ( .A1(n4408), .A2(n4407), .ZN(n4409) );
  XNOR2_X1 U5430 ( .A(n4410), .B(n4409), .ZN(n6285) );
  NAND2_X1 U5431 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4411) );
  OAI21_X1 U5432 ( .B1(n4411), .B2(n3615), .A(n4899), .ZN(n4420) );
  NOR2_X1 U5433 ( .A1(n4413), .A2(n4412), .ZN(n4414) );
  OR2_X1 U5434 ( .A1(n4452), .A2(n4414), .ZN(n4437) );
  INV_X1 U5435 ( .A(REIP_REG_2__SCAN_IN), .ZN(n4415) );
  OAI22_X1 U5436 ( .A1(n6309), .A2(n4437), .B1(n6308), .B2(n4415), .ZN(n4419)
         );
  AOI21_X1 U5438 ( .B1(n5159), .B2(n4451), .A(n4416), .ZN(n4900) );
  OAI33_X1 U5439 ( .A1(1'b0), .A2(n4900), .A3(n3615), .B1(
        INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n3607), .B3(n4450), .ZN(n4418) );
  AOI211_X1 U5440 ( .C1(n5276), .C2(n4420), .A(n4419), .B(n4418), .ZN(n4421)
         );
  OAI21_X1 U5441 ( .B1(n6285), .B2(n6307), .A(n4421), .ZN(U3016) );
  NOR2_X1 U5442 ( .A1(n4423), .A2(n4422), .ZN(n4425) );
  OAI21_X1 U5443 ( .B1(n4426), .B2(n4425), .A(n4424), .ZN(n4427) );
  NAND2_X1 U5444 ( .A1(n4429), .A2(n5445), .ZN(n4430) );
  INV_X1 U5445 ( .A(n4430), .ZN(n4431) );
  INV_X1 U5446 ( .A(DATAI_1_), .ZN(n4536) );
  INV_X1 U5447 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6237) );
  OAI222_X1 U5448 ( .A1(n5246), .A2(n5626), .B1(n4757), .B2(n4536), .C1(n5613), 
        .C2(n6237), .ZN(U2890) );
  INV_X1 U5449 ( .A(n4432), .ZN(n4458) );
  INV_X1 U5450 ( .A(n4433), .ZN(n4434) );
  OR2_X1 U5451 ( .A1(n4435), .A2(n4434), .ZN(n4436) );
  NAND2_X1 U5452 ( .A1(n4458), .A2(n4436), .ZN(n6286) );
  INV_X1 U5453 ( .A(n4437), .ZN(n5184) );
  AOI22_X1 U5454 ( .A1(n6191), .A2(n5184), .B1(EBX_REG_2__SCAN_IN), .B2(n5559), 
        .ZN(n4438) );
  OAI21_X1 U5455 ( .B1(n6286), .B2(n5610), .A(n4438), .ZN(U2857) );
  INV_X2 U5456 ( .A(n6203), .ZN(n5626) );
  INV_X1 U5457 ( .A(DATAI_0_), .ZN(n4529) );
  INV_X1 U5458 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6242) );
  OAI222_X1 U5459 ( .A1(n5626), .A2(n6304), .B1(n4757), .B2(n4529), .C1(n5613), 
        .C2(n6242), .ZN(U2891) );
  INV_X1 U5460 ( .A(DATAI_2_), .ZN(n4515) );
  INV_X1 U5461 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6235) );
  OAI222_X1 U5462 ( .A1(n6286), .A2(n5626), .B1(n4757), .B2(n4515), .C1(n5613), 
        .C2(n6235), .ZN(U2889) );
  OR2_X1 U5463 ( .A1(n4440), .A2(n4439), .ZN(n4441) );
  NAND2_X1 U5464 ( .A1(n4442), .A2(n4441), .ZN(n6337) );
  INV_X1 U5465 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4445) );
  NOR2_X1 U5466 ( .A1(n5246), .A2(n6303), .ZN(n4444) );
  INV_X1 U5467 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5251) );
  OAI22_X1 U5468 ( .A1(n6282), .A2(n4445), .B1(n6308), .B2(n5251), .ZN(n4443)
         );
  AOI211_X1 U5469 ( .C1(n6276), .C2(n4445), .A(n4444), .B(n4443), .ZN(n4446)
         );
  OAI21_X1 U5470 ( .B1(n6297), .B2(n6337), .A(n4446), .ZN(U2985) );
  XNOR2_X1 U5471 ( .A(n4447), .B(n4448), .ZN(n4564) );
  OAI21_X1 U5472 ( .B1(n5155), .B2(n4899), .A(n4900), .ZN(n4613) );
  AOI221_X1 U5473 ( .B1(n4451), .B2(n5155), .C1(n4450), .C2(n5155), .A(n4449), 
        .ZN(n4908) );
  AOI22_X1 U5474 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4613), .B1(n4908), 
        .B2(n3431), .ZN(n4456) );
  INV_X1 U5475 ( .A(n4452), .ZN(n4453) );
  AOI21_X1 U5476 ( .B1(n4454), .B2(n4453), .A(n3628), .ZN(n4460) );
  INV_X1 U5477 ( .A(REIP_REG_3__SCAN_IN), .ZN(n5239) );
  NOR2_X1 U5478 ( .A1(n6308), .A2(n5239), .ZN(n4559) );
  AOI21_X1 U5479 ( .B1(n6333), .B2(n4460), .A(n4559), .ZN(n4455) );
  OAI211_X1 U5480 ( .C1(n4564), .C2(n6307), .A(n4456), .B(n4455), .ZN(U3015)
         );
  INV_X1 U5481 ( .A(n4457), .ZN(n4459) );
  OR2_X1 U5482 ( .A1(n4458), .A2(n4457), .ZN(n4618) );
  OAI21_X1 U5483 ( .B1(n4432), .B2(n4459), .A(n4618), .ZN(n5244) );
  INV_X1 U5484 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4461) );
  INV_X1 U5485 ( .A(n4460), .ZN(n5238) );
  OAI222_X1 U5486 ( .A1(n5244), .A2(n5610), .B1(n4461), .B2(n6195), .C1(n5238), 
        .C2(n5608), .ZN(U2856) );
  INV_X1 U5487 ( .A(DATAI_3_), .ZN(n4522) );
  INV_X1 U5488 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6233) );
  OAI222_X1 U5489 ( .A1(n5244), .A2(n5626), .B1(n4757), .B2(n4522), .C1(n5613), 
        .C2(n6233), .ZN(U2888) );
  INV_X1 U5490 ( .A(n5206), .ZN(n4465) );
  OAI21_X1 U5491 ( .B1(n4463), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4462), 
        .ZN(n6296) );
  NAND2_X1 U5492 ( .A1(n6334), .A2(REIP_REG_0__SCAN_IN), .ZN(n6295) );
  OAI21_X1 U5493 ( .B1(n6307), .B2(n6296), .A(n6295), .ZN(n4464) );
  AOI21_X1 U5494 ( .B1(n6333), .B2(n4465), .A(n4464), .ZN(n4469) );
  INV_X1 U5495 ( .A(n4466), .ZN(n6007) );
  INV_X1 U5496 ( .A(n4467), .ZN(n6330) );
  OAI21_X1 U5497 ( .B1(n6007), .B2(n6330), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4468) );
  OAI211_X1 U5498 ( .C1(INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n6010), .A(n4469), 
        .B(n4468), .ZN(U3018) );
  INV_X1 U5499 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4471) );
  AOI22_X1 U5500 ( .A1(UWORD_REG_2__SCAN_IN), .A2(n6239), .B1(n6229), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4470) );
  OAI21_X1 U5501 ( .B1(n4471), .B2(n4484), .A(n4470), .ZN(U2905) );
  INV_X1 U5502 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4473) );
  AOI22_X1 U5503 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6588), .B1(n6229), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4472) );
  OAI21_X1 U5504 ( .B1(n4473), .B2(n4484), .A(n4472), .ZN(U2902) );
  AOI22_X1 U5505 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n6588), .B1(n6229), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4474) );
  OAI21_X1 U5506 ( .B1(n4091), .B2(n4484), .A(n4474), .ZN(U2901) );
  INV_X1 U5507 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4476) );
  AOI22_X1 U5508 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n6588), .B1(n6229), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4475) );
  OAI21_X1 U5509 ( .B1(n4476), .B2(n4484), .A(n4475), .ZN(U2900) );
  INV_X1 U5510 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4478) );
  AOI22_X1 U5511 ( .A1(UWORD_REG_0__SCAN_IN), .A2(n6239), .B1(n6229), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4477) );
  OAI21_X1 U5512 ( .B1(n4478), .B2(n4484), .A(n4477), .ZN(U2907) );
  INV_X1 U5513 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4480) );
  AOI22_X1 U5514 ( .A1(UWORD_REG_1__SCAN_IN), .A2(n6239), .B1(n6229), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4479) );
  OAI21_X1 U5515 ( .B1(n4480), .B2(n4484), .A(n4479), .ZN(U2906) );
  INV_X1 U5516 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4482) );
  AOI22_X1 U5517 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6588), .B1(n6229), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4481) );
  OAI21_X1 U5518 ( .B1(n4482), .B2(n4484), .A(n4481), .ZN(U2903) );
  INV_X1 U5519 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4485) );
  AOI22_X1 U5520 ( .A1(UWORD_REG_3__SCAN_IN), .A2(n6588), .B1(n6229), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4483) );
  OAI21_X1 U5521 ( .B1(n4485), .B2(n4484), .A(n4483), .ZN(U2904) );
  NAND3_X1 U5522 ( .A1(n5860), .A2(n5856), .A3(n4488), .ZN(n4496) );
  INV_X1 U5523 ( .A(DATAI_23_), .ZN(n4486) );
  OR2_X1 U5524 ( .A1(n6303), .A2(n4486), .ZN(n6397) );
  INV_X1 U5525 ( .A(DATAI_31_), .ZN(n4487) );
  OR2_X1 U5526 ( .A1(n6303), .A2(n4487), .ZN(n6445) );
  INV_X1 U5527 ( .A(n6445), .ZN(n6393) );
  AND2_X1 U5528 ( .A1(n4674), .A2(n4488), .ZN(n4489) );
  NOR2_X1 U5529 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6592) );
  INV_X1 U5530 ( .A(n6592), .ZN(n5121) );
  NOR2_X1 U5531 ( .A1(n4549), .A2(n5612), .ZN(n6436) );
  INV_X1 U5532 ( .A(n6436), .ZN(n5085) );
  NAND2_X1 U5533 ( .A1(n4490), .A2(n3036), .ZN(n4928) );
  INV_X1 U5534 ( .A(n4342), .ZN(n5249) );
  NAND2_X1 U5535 ( .A1(n5183), .A2(n5249), .ZN(n4966) );
  OR2_X1 U5536 ( .A1(n4928), .A2(n4966), .ZN(n4492) );
  NAND2_X1 U5537 ( .A1(n4492), .A2(n4663), .ZN(n4498) );
  AOI22_X1 U5538 ( .A1(n4498), .A2(n6350), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4493), .ZN(n4662) );
  INV_X1 U5539 ( .A(DATAI_7_), .ZN(n6766) );
  NOR2_X1 U5540 ( .A1(n6766), .A2(n4856), .ZN(n6440) );
  INV_X1 U5541 ( .A(n6440), .ZN(n5355) );
  OAI22_X1 U5542 ( .A1(n5085), .A2(n4663), .B1(n4662), .B2(n5355), .ZN(n4495)
         );
  AOI21_X1 U5543 ( .B1(n6393), .B2(n4996), .A(n4495), .ZN(n4501) );
  NAND2_X1 U5544 ( .A1(n6350), .A2(n6760), .ZN(n5009) );
  INV_X1 U5545 ( .A(n5009), .ZN(n5874) );
  AOI21_X1 U5546 ( .B1(n4496), .B2(n6287), .A(n5874), .ZN(n4499) );
  OAI21_X1 U5547 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6567), .A(n4961), 
        .ZN(n4933) );
  AOI21_X1 U5548 ( .B1(n4960), .B2(n6347), .A(n4933), .ZN(n4497) );
  OAI21_X1 U5549 ( .B1(n4499), .B2(n4498), .A(n4497), .ZN(n4665) );
  NAND2_X1 U5550 ( .A1(n4665), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4500)
         );
  OAI211_X1 U5551 ( .C1(n4668), .C2(n6397), .A(n4501), .B(n4500), .ZN(U3147)
         );
  INV_X1 U5552 ( .A(DATAI_20_), .ZN(n4502) );
  OR2_X1 U5553 ( .A1(n6303), .A2(n4502), .ZN(n6381) );
  INV_X1 U5554 ( .A(DATAI_28_), .ZN(n4503) );
  OR2_X1 U5555 ( .A1(n6303), .A2(n4503), .ZN(n5084) );
  INV_X1 U5556 ( .A(n5084), .ZN(n6378) );
  NOR2_X1 U5557 ( .A1(n4549), .A2(n3270), .ZN(n6377) );
  INV_X1 U5558 ( .A(n6377), .ZN(n5079) );
  INV_X1 U5559 ( .A(DATAI_4_), .ZN(n4624) );
  NOR2_X1 U5560 ( .A1(n4624), .A2(n4856), .ZN(n6376) );
  INV_X1 U5561 ( .A(n6376), .ZN(n5351) );
  OAI22_X1 U5562 ( .A1(n5079), .A2(n4663), .B1(n4662), .B2(n5351), .ZN(n4504)
         );
  AOI21_X1 U5563 ( .B1(n6378), .B2(n4996), .A(n4504), .ZN(n4506) );
  NAND2_X1 U5564 ( .A1(n4665), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4505)
         );
  OAI211_X1 U5565 ( .C1(n4668), .C2(n6381), .A(n4506), .B(n4505), .ZN(U3144)
         );
  INV_X1 U5566 ( .A(DATAI_22_), .ZN(n4507) );
  OR2_X1 U5567 ( .A1(n6303), .A2(n4507), .ZN(n6389) );
  INV_X1 U5568 ( .A(DATAI_30_), .ZN(n4508) );
  OR2_X1 U5569 ( .A1(n6303), .A2(n4508), .ZN(n6416) );
  INV_X1 U5570 ( .A(n6416), .ZN(n6386) );
  INV_X1 U5571 ( .A(n6409), .ZN(n5089) );
  INV_X1 U5572 ( .A(DATAI_6_), .ZN(n4756) );
  NOR2_X1 U5573 ( .A1(n4756), .A2(n4856), .ZN(n6411) );
  INV_X1 U5574 ( .A(n6411), .ZN(n5347) );
  OAI22_X1 U5575 ( .A1(n5089), .A2(n4663), .B1(n4662), .B2(n5347), .ZN(n4509)
         );
  AOI21_X1 U5576 ( .B1(n6386), .B2(n4996), .A(n4509), .ZN(n4511) );
  NAND2_X1 U5577 ( .A1(n4665), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4510)
         );
  OAI211_X1 U5578 ( .C1(n4668), .C2(n6389), .A(n4511), .B(n4510), .ZN(U3146)
         );
  INV_X1 U5579 ( .A(DATAI_18_), .ZN(n4512) );
  OR2_X1 U5580 ( .A1(n6303), .A2(n4512), .ZN(n6371) );
  INV_X1 U5581 ( .A(DATAI_26_), .ZN(n4513) );
  OR2_X1 U5582 ( .A1(n6303), .A2(n4513), .ZN(n5114) );
  INV_X1 U5583 ( .A(n5114), .ZN(n6368) );
  NOR2_X1 U5584 ( .A1(n4549), .A2(n4514), .ZN(n6367) );
  INV_X1 U5585 ( .A(n6367), .ZN(n5108) );
  NOR2_X1 U5586 ( .A1(n4515), .A2(n4856), .ZN(n6366) );
  INV_X1 U5587 ( .A(n6366), .ZN(n5359) );
  OAI22_X1 U5588 ( .A1(n5108), .A2(n4663), .B1(n4662), .B2(n5359), .ZN(n4516)
         );
  AOI21_X1 U5589 ( .B1(n6368), .B2(n4996), .A(n4516), .ZN(n4518) );
  NAND2_X1 U5590 ( .A1(n4665), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4517)
         );
  OAI211_X1 U5591 ( .C1(n4668), .C2(n6371), .A(n4518), .B(n4517), .ZN(U3142)
         );
  INV_X1 U5592 ( .A(DATAI_19_), .ZN(n4519) );
  OR2_X1 U5593 ( .A1(n6303), .A2(n4519), .ZN(n6375) );
  INV_X1 U5594 ( .A(DATAI_27_), .ZN(n4520) );
  OR2_X1 U5595 ( .A1(n6303), .A2(n4520), .ZN(n6405) );
  INV_X1 U5596 ( .A(n6405), .ZN(n6372) );
  NOR2_X1 U5597 ( .A1(n4549), .A2(n4521), .ZN(n6401) );
  INV_X1 U5598 ( .A(n6401), .ZN(n5075) );
  NOR2_X1 U5599 ( .A1(n4522), .A2(n4856), .ZN(n6402) );
  INV_X1 U5600 ( .A(n6402), .ZN(n5343) );
  OAI22_X1 U5601 ( .A1(n5075), .A2(n4663), .B1(n4662), .B2(n5343), .ZN(n4523)
         );
  AOI21_X1 U5602 ( .B1(n6372), .B2(n4996), .A(n4523), .ZN(n4525) );
  NAND2_X1 U5603 ( .A1(n4665), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4524)
         );
  OAI211_X1 U5604 ( .C1(n4668), .C2(n6375), .A(n4525), .B(n4524), .ZN(U3143)
         );
  INV_X1 U5605 ( .A(DATAI_16_), .ZN(n4526) );
  OR2_X1 U5606 ( .A1(n6303), .A2(n4526), .ZN(n6361) );
  INV_X1 U5607 ( .A(DATAI_24_), .ZN(n4527) );
  OR2_X1 U5608 ( .A1(n6303), .A2(n4527), .ZN(n6422) );
  INV_X1 U5609 ( .A(n6422), .ZN(n6358) );
  NOR2_X1 U5610 ( .A1(n4549), .A2(n4528), .ZN(n6417) );
  INV_X1 U5611 ( .A(n6417), .ZN(n5097) );
  NOR2_X1 U5612 ( .A1(n4529), .A2(n4856), .ZN(n6419) );
  INV_X1 U5613 ( .A(n6419), .ZN(n5370) );
  OAI22_X1 U5614 ( .A1(n5097), .A2(n4663), .B1(n4662), .B2(n5370), .ZN(n4530)
         );
  AOI21_X1 U5615 ( .B1(n6358), .B2(n4996), .A(n4530), .ZN(n4532) );
  NAND2_X1 U5616 ( .A1(n4665), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4531)
         );
  OAI211_X1 U5617 ( .C1(n4668), .C2(n6361), .A(n4532), .B(n4531), .ZN(U3140)
         );
  INV_X1 U5618 ( .A(DATAI_17_), .ZN(n4533) );
  OR2_X1 U5619 ( .A1(n6303), .A2(n4533), .ZN(n6365) );
  INV_X1 U5620 ( .A(DATAI_25_), .ZN(n4534) );
  OR2_X1 U5621 ( .A1(n6303), .A2(n4534), .ZN(n6428) );
  INV_X1 U5622 ( .A(n6428), .ZN(n6362) );
  NOR2_X1 U5623 ( .A1(n4549), .A2(n4535), .ZN(n6423) );
  INV_X1 U5624 ( .A(n6423), .ZN(n5101) );
  NOR2_X1 U5625 ( .A1(n4536), .A2(n4856), .ZN(n6425) );
  INV_X1 U5626 ( .A(n6425), .ZN(n5339) );
  OAI22_X1 U5627 ( .A1(n5101), .A2(n4663), .B1(n4662), .B2(n5339), .ZN(n4537)
         );
  AOI21_X1 U5628 ( .B1(n6362), .B2(n4996), .A(n4537), .ZN(n4539) );
  NAND2_X1 U5629 ( .A1(n4665), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4538)
         );
  OAI211_X1 U5630 ( .C1(n4668), .C2(n6365), .A(n4539), .B(n4538), .ZN(U3141)
         );
  NOR2_X1 U5631 ( .A1(n4804), .A2(n6760), .ZN(n5859) );
  NAND2_X1 U5632 ( .A1(n4805), .A2(n5859), .ZN(n4603) );
  NAND2_X1 U5633 ( .A1(n6350), .A2(n4603), .ZN(n4544) );
  INV_X1 U5634 ( .A(n6349), .ZN(n4541) );
  INV_X1 U5635 ( .A(n4540), .ZN(n6408) );
  AOI21_X1 U5636 ( .B1(n4541), .B2(n3036), .A(n6408), .ZN(n4545) );
  INV_X1 U5637 ( .A(n4545), .ZN(n4543) );
  AOI21_X1 U5638 ( .B1(n6343), .B2(n6347), .A(n4933), .ZN(n4542) );
  OAI21_X1 U5639 ( .B1(n4544), .B2(n4543), .A(n4542), .ZN(n6412) );
  OAI22_X1 U5640 ( .A1(n4545), .A2(n4544), .B1(n5335), .B2(n6343), .ZN(n6410)
         );
  AOI22_X1 U5641 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6412), .B1(n6366), 
        .B2(n6410), .ZN(n4547) );
  NOR2_X1 U5642 ( .A1(n4804), .A2(n3815), .ZN(n4675) );
  INV_X1 U5643 ( .A(n6371), .ZN(n5111) );
  AOI22_X1 U5644 ( .A1(n6367), .A2(n6408), .B1(n6407), .B2(n5111), .ZN(n4546)
         );
  OAI211_X1 U5645 ( .C1(n5114), .C2(n6415), .A(n4547), .B(n4546), .ZN(U3078)
         );
  INV_X1 U5646 ( .A(DATAI_29_), .ZN(n6602) );
  OR2_X1 U5647 ( .A1(n6303), .A2(n6602), .ZN(n6434) );
  NOR2_X1 U5648 ( .A1(n4548), .A2(n4856), .ZN(n6431) );
  AOI22_X1 U5649 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6412), .B1(n6431), 
        .B2(n6410), .ZN(n4552) );
  NOR2_X1 U5650 ( .A1(n4549), .A2(n3222), .ZN(n6429) );
  INV_X1 U5651 ( .A(DATAI_21_), .ZN(n4550) );
  OR2_X1 U5652 ( .A1(n6303), .A2(n4550), .ZN(n6385) );
  INV_X1 U5653 ( .A(n6385), .ZN(n6430) );
  AOI22_X1 U5654 ( .A1(n6429), .A2(n6408), .B1(n6407), .B2(n6430), .ZN(n4551)
         );
  OAI211_X1 U5655 ( .C1(n6434), .C2(n6415), .A(n4552), .B(n4551), .ZN(U3081)
         );
  AOI22_X1 U5656 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6412), .B1(n6376), 
        .B2(n6410), .ZN(n4554) );
  INV_X1 U5657 ( .A(n6381), .ZN(n5081) );
  AOI22_X1 U5658 ( .A1(n6377), .A2(n6408), .B1(n6407), .B2(n5081), .ZN(n4553)
         );
  OAI211_X1 U5659 ( .C1(n5084), .C2(n6415), .A(n4554), .B(n4553), .ZN(U3080)
         );
  AOI22_X1 U5660 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6412), .B1(n6440), 
        .B2(n6410), .ZN(n4556) );
  INV_X1 U5661 ( .A(n6397), .ZN(n6437) );
  AOI22_X1 U5662 ( .A1(n6436), .A2(n6408), .B1(n6407), .B2(n6437), .ZN(n4555)
         );
  OAI211_X1 U5663 ( .C1(n6445), .C2(n6415), .A(n4556), .B(n4555), .ZN(U3083)
         );
  AOI22_X1 U5664 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6412), .B1(n6425), 
        .B2(n6410), .ZN(n4558) );
  INV_X1 U5665 ( .A(n6365), .ZN(n6424) );
  AOI22_X1 U5666 ( .A1(n6423), .A2(n6408), .B1(n6407), .B2(n6424), .ZN(n4557)
         );
  OAI211_X1 U5667 ( .C1(n6428), .C2(n6415), .A(n4558), .B(n4557), .ZN(U3077)
         );
  INV_X1 U5668 ( .A(n5244), .ZN(n4562) );
  AOI21_X1 U5669 ( .B1(n6300), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4559), 
        .ZN(n4560) );
  OAI21_X1 U5670 ( .B1(n5234), .B2(n6294), .A(n4560), .ZN(n4561) );
  AOI21_X1 U5671 ( .B1(n4562), .B2(n6287), .A(n4561), .ZN(n4563) );
  OAI21_X1 U5672 ( .B1(n4564), .B2(n6297), .A(n4563), .ZN(U2983) );
  INV_X1 U5673 ( .A(n5183), .ZN(n5862) );
  NAND2_X1 U5674 ( .A1(n4566), .A2(n4565), .ZN(n4572) );
  XNOR2_X1 U5675 ( .A(n4351), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4569)
         );
  INV_X1 U5676 ( .A(n6449), .ZN(n4581) );
  XNOR2_X1 U5677 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4567) );
  OAI22_X1 U5678 ( .A1(n4581), .A2(n4567), .B1(n4579), .B2(n4569), .ZN(n4568)
         );
  AOI21_X1 U5679 ( .B1(n4572), .B2(n4569), .A(n4568), .ZN(n4570) );
  OAI21_X1 U5680 ( .B1(n5862), .B2(n4571), .A(n4570), .ZN(n5408) );
  MUX2_X1 U5681 ( .A(n5408), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(n4584), 
        .Z(n6456) );
  NAND2_X1 U5682 ( .A1(n6456), .A2(n6474), .ZN(n4587) );
  INV_X1 U5683 ( .A(n4571), .ZN(n6448) );
  INV_X1 U5684 ( .A(n4572), .ZN(n4575) );
  MUX2_X1 U5685 ( .A(n4573), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4351), 
        .Z(n4574) );
  NOR3_X1 U5686 ( .A1(n4575), .A2(n4585), .A3(n4574), .ZN(n4583) );
  NAND2_X1 U5687 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4577) );
  INV_X1 U5688 ( .A(n4577), .ZN(n4576) );
  MUX2_X1 U5689 ( .A(n4577), .B(n4576), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4580) );
  INV_X1 U5690 ( .A(n4351), .ZN(n5404) );
  AOI211_X1 U5691 ( .C1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n5404), .A(n4578), .B(n3331), .ZN(n5866) );
  OAI22_X1 U5692 ( .A1(n4581), .A2(n4580), .B1(n5866), .B2(n4579), .ZN(n4582)
         );
  MUX2_X1 U5693 ( .A(n5867), .B(n3108), .S(n4584), .Z(n6459) );
  INV_X1 U5694 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6037) );
  NAND2_X1 U5695 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6037), .ZN(n4591) );
  INV_X1 U5696 ( .A(n4585), .ZN(n4586) );
  OAI22_X1 U5697 ( .A1(n4587), .A2(n6459), .B1(n4591), .B2(n4586), .ZN(n6467)
         );
  INV_X1 U5698 ( .A(n4352), .ZN(n4588) );
  NAND2_X1 U5699 ( .A1(n6467), .A2(n4588), .ZN(n4598) );
  INV_X1 U5700 ( .A(n5066), .ZN(n4801) );
  OR2_X1 U5701 ( .A1(n4589), .A2(n4801), .ZN(n4590) );
  XNOR2_X1 U5702 ( .A(n4590), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6171)
         );
  INV_X1 U5703 ( .A(n6171), .ZN(n6026) );
  OAI22_X1 U5704 ( .A1(n6450), .A2(n3779), .B1(n6026), .B2(n2999), .ZN(n4593)
         );
  INV_X1 U5705 ( .A(n4591), .ZN(n4592) );
  AOI22_X1 U5706 ( .A1(n4593), .A2(n6474), .B1(n4592), .B2(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6466) );
  AND3_X1 U5707 ( .A1(n4598), .A2(n6466), .A3(n6037), .ZN(n4595) );
  INV_X1 U5708 ( .A(n4594), .ZN(n6564) );
  OAI21_X1 U5709 ( .B1(n4595), .B2(n6564), .A(n4856), .ZN(n6342) );
  INV_X1 U5710 ( .A(n4596), .ZN(n4597) );
  AND3_X1 U5711 ( .A1(n4598), .A2(n6466), .A3(n4597), .ZN(n6476) );
  INV_X1 U5712 ( .A(n3036), .ZN(n5204) );
  AND2_X1 U5713 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6567), .ZN(n5861) );
  OAI22_X1 U5714 ( .A1(n3815), .A2(n6347), .B1(n5204), .B2(n5861), .ZN(n4599)
         );
  OAI21_X1 U5715 ( .B1(n6476), .B2(n4599), .A(n6342), .ZN(n4600) );
  OAI21_X1 U5716 ( .B1(n6342), .B2(n4930), .A(n4600), .ZN(U3465) );
  NOR2_X1 U5717 ( .A1(n5856), .A2(n4601), .ZN(n4602) );
  NAND2_X1 U5718 ( .A1(n4635), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4628) );
  AND2_X1 U5719 ( .A1(n4628), .A2(n4852), .ZN(n4759) );
  AOI21_X1 U5720 ( .B1(n4759), .B2(n4603), .A(n6347), .ZN(n4605) );
  OAI22_X1 U5721 ( .A1(n3001), .A2(n5009), .B1(n5877), .B2(n5861), .ZN(n4604)
         );
  OAI21_X1 U5722 ( .B1(n4605), .B2(n4604), .A(n6342), .ZN(n4606) );
  OAI21_X1 U5723 ( .B1(n6342), .B2(n6357), .A(n4606), .ZN(U3462) );
  XNOR2_X1 U5724 ( .A(n4608), .B(n4607), .ZN(n4623) );
  INV_X1 U5725 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6517) );
  NOR2_X1 U5726 ( .A1(n6308), .A2(n6517), .ZN(n4619) );
  NAND2_X1 U5727 ( .A1(n4610), .A2(n4609), .ZN(n4611) );
  NAND2_X1 U5728 ( .A1(n4912), .A2(n4611), .ZN(n6174) );
  NOR2_X1 U5729 ( .A1(n6309), .A2(n6174), .ZN(n4612) );
  AOI211_X1 U5730 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n4613), .A(n4619), 
        .B(n4612), .ZN(n4615) );
  OAI211_X1 U5731 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4908), .B(n4910), .ZN(n4614) );
  OAI211_X1 U5732 ( .C1(n6307), .C2(n4623), .A(n4615), .B(n4614), .ZN(U3014)
         );
  AND2_X1 U5733 ( .A1(n4432), .A2(n4617), .ZN(n4846) );
  AOI21_X1 U5734 ( .B1(n4616), .B2(n4618), .A(n4846), .ZN(n6183) );
  AOI21_X1 U5735 ( .B1(n6300), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n4619), 
        .ZN(n4620) );
  OAI21_X1 U5736 ( .B1(n6179), .B2(n6294), .A(n4620), .ZN(n4621) );
  AOI21_X1 U5737 ( .B1(n6183), .B2(n6287), .A(n4621), .ZN(n4622) );
  OAI21_X1 U5738 ( .B1(n6297), .B2(n4623), .A(n4622), .ZN(U2982) );
  INV_X1 U5739 ( .A(n6183), .ZN(n4755) );
  INV_X1 U5740 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6231) );
  OAI222_X1 U5741 ( .A1(n4755), .A2(n5626), .B1(n4757), .B2(n4624), .C1(n5613), 
        .C2(n6231), .ZN(U2887) );
  AND2_X1 U5742 ( .A1(n5183), .A2(n4342), .ZN(n5072) );
  INV_X1 U5743 ( .A(n5072), .ZN(n4625) );
  OR2_X1 U5744 ( .A1(n4625), .A2(n4928), .ZN(n4627) );
  NAND2_X1 U5745 ( .A1(n6453), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4632) );
  INV_X1 U5746 ( .A(n4632), .ZN(n4802) );
  NAND2_X1 U5747 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4802), .ZN(n5067) );
  NOR2_X1 U5748 ( .A1(n4930), .A2(n5067), .ZN(n4659) );
  INV_X1 U5749 ( .A(n4659), .ZN(n4626) );
  AND2_X1 U5750 ( .A1(n4627), .A2(n4626), .ZN(n4634) );
  INV_X1 U5751 ( .A(n4634), .ZN(n4630) );
  NAND2_X1 U5752 ( .A1(n6350), .A2(n4628), .ZN(n4633) );
  AOI21_X1 U5753 ( .B1(n6347), .B2(n5067), .A(n4933), .ZN(n4629) );
  OAI21_X1 U5754 ( .B1(n4630), .B2(n4633), .A(n4629), .ZN(n4658) );
  NAND2_X1 U5755 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4631) );
  OAI22_X1 U5756 ( .A1(n4634), .A2(n4633), .B1(n4632), .B2(n4631), .ZN(n4657)
         );
  AOI22_X1 U5757 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4658), .B1(n6411), 
        .B2(n4657), .ZN(n4637) );
  AOI22_X1 U5758 ( .A1(n6409), .A2(n4659), .B1(n5110), .B2(n6386), .ZN(n4636)
         );
  OAI211_X1 U5759 ( .C1(n6389), .C2(n4999), .A(n4637), .B(n4636), .ZN(U3130)
         );
  AOI22_X1 U5760 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4658), .B1(n6402), 
        .B2(n4657), .ZN(n4639) );
  AOI22_X1 U5761 ( .A1(n6401), .A2(n4659), .B1(n5110), .B2(n6372), .ZN(n4638)
         );
  OAI211_X1 U5762 ( .C1(n6375), .C2(n4999), .A(n4639), .B(n4638), .ZN(U3127)
         );
  AOI22_X1 U5763 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4658), .B1(n6419), 
        .B2(n4657), .ZN(n4641) );
  AOI22_X1 U5764 ( .A1(n6417), .A2(n4659), .B1(n5110), .B2(n6358), .ZN(n4640)
         );
  OAI211_X1 U5765 ( .C1(n6361), .C2(n4999), .A(n4641), .B(n4640), .ZN(U3124)
         );
  AOI22_X1 U5766 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4658), .B1(n6376), 
        .B2(n4657), .ZN(n4643) );
  AOI22_X1 U5767 ( .A1(n6377), .A2(n4659), .B1(n5110), .B2(n6378), .ZN(n4642)
         );
  OAI211_X1 U5768 ( .C1(n6381), .C2(n4999), .A(n4643), .B(n4642), .ZN(U3128)
         );
  AOI22_X1 U5769 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4658), .B1(n6440), 
        .B2(n4657), .ZN(n4645) );
  AOI22_X1 U5770 ( .A1(n6436), .A2(n4659), .B1(n5110), .B2(n6393), .ZN(n4644)
         );
  OAI211_X1 U5771 ( .C1(n6397), .C2(n4999), .A(n4645), .B(n4644), .ZN(U3131)
         );
  AOI22_X1 U5772 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4658), .B1(n6366), 
        .B2(n4657), .ZN(n4647) );
  AOI22_X1 U5773 ( .A1(n6367), .A2(n4659), .B1(n5110), .B2(n6368), .ZN(n4646)
         );
  OAI211_X1 U5774 ( .C1(n6371), .C2(n4999), .A(n4647), .B(n4646), .ZN(U3126)
         );
  AOI22_X1 U5775 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4658), .B1(n6425), 
        .B2(n4657), .ZN(n4649) );
  AOI22_X1 U5776 ( .A1(n6423), .A2(n4659), .B1(n5110), .B2(n6362), .ZN(n4648)
         );
  OAI211_X1 U5777 ( .C1(n6365), .C2(n4999), .A(n4649), .B(n4648), .ZN(U3125)
         );
  OAI21_X1 U5778 ( .B1(n4650), .B2(n4652), .A(n4651), .ZN(n6152) );
  AND2_X1 U5779 ( .A1(n4914), .A2(n4653), .ZN(n4654) );
  OR2_X1 U5780 ( .A1(n4654), .A2(n5005), .ZN(n6146) );
  INV_X1 U5781 ( .A(n6146), .ZN(n4655) );
  AOI22_X1 U5782 ( .A1(n6191), .A2(n4655), .B1(EBX_REG_6__SCAN_IN), .B2(n5559), 
        .ZN(n4656) );
  OAI21_X1 U5783 ( .B1(n6152), .B2(n5610), .A(n4656), .ZN(U2853) );
  AOI22_X1 U5784 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4658), .B1(n6431), 
        .B2(n4657), .ZN(n4661) );
  INV_X1 U5785 ( .A(n6434), .ZN(n6382) );
  AOI22_X1 U5786 ( .A1(n6429), .A2(n4659), .B1(n5110), .B2(n6382), .ZN(n4660)
         );
  OAI211_X1 U5787 ( .C1(n6385), .C2(n4999), .A(n4661), .B(n4660), .ZN(U3129)
         );
  INV_X1 U5788 ( .A(n6429), .ZN(n5093) );
  INV_X1 U5789 ( .A(n6431), .ZN(n5363) );
  OAI22_X1 U5790 ( .A1(n5093), .A2(n4663), .B1(n4662), .B2(n5363), .ZN(n4664)
         );
  AOI21_X1 U5791 ( .B1(n6382), .B2(n4996), .A(n4664), .ZN(n4667) );
  NAND2_X1 U5792 ( .A1(n4665), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4666)
         );
  OAI211_X1 U5793 ( .C1(n4668), .C2(n6385), .A(n4667), .B(n4666), .ZN(U3145)
         );
  INV_X1 U5794 ( .A(n5859), .ZN(n4669) );
  OAI21_X1 U5795 ( .B1(n4852), .B2(n4669), .A(n6350), .ZN(n4673) );
  NOR2_X1 U5796 ( .A1(n5183), .A2(n4342), .ZN(n4761) );
  NOR2_X1 U5797 ( .A1(n4762), .A2(n6357), .ZN(n6435) );
  AOI21_X1 U5798 ( .B1(n5329), .B2(n3036), .A(n6435), .ZN(n4670) );
  NAND3_X1 U5799 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6458), .ZN(n5328) );
  OAI22_X1 U5800 ( .A1(n4673), .A2(n4670), .B1(n5328), .B2(n5335), .ZN(n6439)
         );
  INV_X1 U5801 ( .A(n6439), .ZN(n4688) );
  INV_X1 U5802 ( .A(n4670), .ZN(n4672) );
  AOI21_X1 U5803 ( .B1(n5328), .B2(n6347), .A(n4933), .ZN(n4671) );
  OAI21_X1 U5804 ( .B1(n4673), .B2(n4672), .A(n4671), .ZN(n6441) );
  INV_X1 U5805 ( .A(n4674), .ZN(n4770) );
  INV_X1 U5806 ( .A(n4675), .ZN(n4772) );
  INV_X1 U5807 ( .A(n6375), .ZN(n6400) );
  AOI22_X1 U5808 ( .A1(n6438), .A2(n6400), .B1(n6401), .B2(n6435), .ZN(n4676)
         );
  OAI21_X1 U5809 ( .B1(n6405), .B2(n6444), .A(n4676), .ZN(n4677) );
  AOI21_X1 U5810 ( .B1(n6441), .B2(INSTQUEUE_REG_11__3__SCAN_IN), .A(n4677), 
        .ZN(n4678) );
  OAI21_X1 U5811 ( .B1(n4688), .B2(n5343), .A(n4678), .ZN(U3111) );
  AOI22_X1 U5812 ( .A1(n6438), .A2(n5081), .B1(n6377), .B2(n6435), .ZN(n4679)
         );
  OAI21_X1 U5813 ( .B1(n5084), .B2(n6444), .A(n4679), .ZN(n4680) );
  AOI21_X1 U5814 ( .B1(n6441), .B2(INSTQUEUE_REG_11__4__SCAN_IN), .A(n4680), 
        .ZN(n4681) );
  OAI21_X1 U5815 ( .B1(n4688), .B2(n5351), .A(n4681), .ZN(U3112) );
  AOI22_X1 U5816 ( .A1(n6438), .A2(n5111), .B1(n6367), .B2(n6435), .ZN(n4682)
         );
  OAI21_X1 U5817 ( .B1(n5114), .B2(n6444), .A(n4682), .ZN(n4683) );
  AOI21_X1 U5818 ( .B1(n6441), .B2(INSTQUEUE_REG_11__2__SCAN_IN), .A(n4683), 
        .ZN(n4684) );
  OAI21_X1 U5819 ( .B1(n4688), .B2(n5359), .A(n4684), .ZN(U3110) );
  INV_X1 U5820 ( .A(n6389), .ZN(n6406) );
  AOI22_X1 U5821 ( .A1(n6438), .A2(n6406), .B1(n6409), .B2(n6435), .ZN(n4685)
         );
  OAI21_X1 U5822 ( .B1(n6416), .B2(n6444), .A(n4685), .ZN(n4686) );
  AOI21_X1 U5823 ( .B1(n6441), .B2(INSTQUEUE_REG_11__6__SCAN_IN), .A(n4686), 
        .ZN(n4687) );
  OAI21_X1 U5824 ( .B1(n4688), .B2(n5347), .A(n4687), .ZN(U3114) );
  NAND3_X1 U5825 ( .A1(n3001), .A2(n4758), .A3(n4804), .ZN(n4696) );
  INV_X1 U5826 ( .A(n4696), .ZN(n4689) );
  OAI21_X1 U5827 ( .B1(n4696), .B2(n6760), .A(n6350), .ZN(n4695) );
  NOR2_X1 U5828 ( .A1(n5183), .A2(n5249), .ZN(n4927) );
  NAND2_X1 U5829 ( .A1(n5877), .A2(n4927), .ZN(n4722) );
  OR2_X1 U5830 ( .A1(n4722), .A2(n5204), .ZN(n4691) );
  NAND3_X1 U5831 ( .A1(n6357), .A2(n6458), .A3(n6453), .ZN(n4718) );
  NOR2_X1 U5832 ( .A1(n4930), .A2(n4718), .ZN(n4713) );
  INV_X1 U5833 ( .A(n4713), .ZN(n4690) );
  AND2_X1 U5834 ( .A1(n4691), .A2(n4690), .ZN(n4694) );
  INV_X1 U5835 ( .A(n4694), .ZN(n4693) );
  AOI21_X1 U5836 ( .B1(n6347), .B2(n4718), .A(n4933), .ZN(n4692) );
  OAI21_X1 U5837 ( .B1(n4695), .B2(n4693), .A(n4692), .ZN(n4712) );
  OAI22_X1 U5838 ( .A1(n4695), .A2(n4694), .B1(n5335), .B2(n4718), .ZN(n4711)
         );
  AOI22_X1 U5839 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4712), .B1(n6376), 
        .B2(n4711), .ZN(n4698) );
  AOI22_X1 U5840 ( .A1(n4716), .A2(n6378), .B1(n6377), .B2(n4713), .ZN(n4697)
         );
  OAI211_X1 U5841 ( .C1(n6381), .C2(n5046), .A(n4698), .B(n4697), .ZN(U3032)
         );
  AOI22_X1 U5842 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4712), .B1(n6402), 
        .B2(n4711), .ZN(n4700) );
  AOI22_X1 U5843 ( .A1(n4716), .A2(n6372), .B1(n6401), .B2(n4713), .ZN(n4699)
         );
  OAI211_X1 U5844 ( .C1(n6375), .C2(n5046), .A(n4700), .B(n4699), .ZN(U3031)
         );
  AOI22_X1 U5845 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4712), .B1(n6419), 
        .B2(n4711), .ZN(n4702) );
  AOI22_X1 U5846 ( .A1(n4716), .A2(n6358), .B1(n6417), .B2(n4713), .ZN(n4701)
         );
  OAI211_X1 U5847 ( .C1(n6361), .C2(n5046), .A(n4702), .B(n4701), .ZN(U3028)
         );
  AOI22_X1 U5848 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4712), .B1(n6431), 
        .B2(n4711), .ZN(n4704) );
  AOI22_X1 U5849 ( .A1(n4716), .A2(n6382), .B1(n6429), .B2(n4713), .ZN(n4703)
         );
  OAI211_X1 U5850 ( .C1(n6385), .C2(n5046), .A(n4704), .B(n4703), .ZN(U3033)
         );
  AOI22_X1 U5851 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4712), .B1(n6440), 
        .B2(n4711), .ZN(n4706) );
  AOI22_X1 U5852 ( .A1(n4716), .A2(n6393), .B1(n6436), .B2(n4713), .ZN(n4705)
         );
  OAI211_X1 U5853 ( .C1(n6397), .C2(n5046), .A(n4706), .B(n4705), .ZN(U3035)
         );
  AOI22_X1 U5854 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4712), .B1(n6425), 
        .B2(n4711), .ZN(n4708) );
  AOI22_X1 U5855 ( .A1(n4716), .A2(n6362), .B1(n6423), .B2(n4713), .ZN(n4707)
         );
  OAI211_X1 U5856 ( .C1(n6365), .C2(n5046), .A(n4708), .B(n4707), .ZN(U3029)
         );
  AOI22_X1 U5857 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4712), .B1(n6411), 
        .B2(n4711), .ZN(n4710) );
  AOI22_X1 U5858 ( .A1(n4716), .A2(n6386), .B1(n6409), .B2(n4713), .ZN(n4709)
         );
  OAI211_X1 U5859 ( .C1(n6389), .C2(n5046), .A(n4710), .B(n4709), .ZN(U3034)
         );
  AOI22_X1 U5860 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4712), .B1(n6366), 
        .B2(n4711), .ZN(n4715) );
  AOI22_X1 U5861 ( .A1(n4716), .A2(n6368), .B1(n6367), .B2(n4713), .ZN(n4714)
         );
  OAI211_X1 U5862 ( .C1(n6371), .C2(n5046), .A(n4715), .B(n4714), .ZN(U3030)
         );
  NOR3_X1 U5863 ( .A1(n4716), .A2(n4751), .A3(n6347), .ZN(n4717) );
  OAI21_X1 U5864 ( .B1(n4717), .B2(n5874), .A(n4722), .ZN(n4721) );
  OR2_X1 U5865 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4718), .ZN(n4749)
         );
  AND2_X1 U5866 ( .A1(n4724), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6345) );
  INV_X1 U5867 ( .A(n4855), .ZN(n4719) );
  OAI21_X1 U5868 ( .B1(n3102), .B2(n5335), .A(n4961), .ZN(n5870) );
  AOI211_X1 U5869 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4749), .A(n6345), .B(
        n5870), .ZN(n4720) );
  NAND2_X1 U5870 ( .A1(n4721), .A2(n4720), .ZN(n4747) );
  NAND2_X1 U5871 ( .A1(n4747), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4728) );
  INV_X1 U5872 ( .A(n4722), .ZN(n4725) );
  NOR2_X1 U5873 ( .A1(n4724), .A2(n4723), .ZN(n6353) );
  AOI22_X1 U5874 ( .A1(n4725), .A2(n6350), .B1(n6353), .B2(n3102), .ZN(n4748)
         );
  OAI22_X1 U5875 ( .A1(n5093), .A2(n4749), .B1(n4748), .B2(n5363), .ZN(n4726)
         );
  AOI21_X1 U5876 ( .B1(n6382), .B2(n4751), .A(n4726), .ZN(n4727) );
  OAI211_X1 U5877 ( .C1(n4754), .C2(n6385), .A(n4728), .B(n4727), .ZN(U3025)
         );
  NAND2_X1 U5878 ( .A1(n4747), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4731) );
  OAI22_X1 U5879 ( .A1(n5089), .A2(n4749), .B1(n4748), .B2(n5347), .ZN(n4729)
         );
  AOI21_X1 U5880 ( .B1(n6386), .B2(n4751), .A(n4729), .ZN(n4730) );
  OAI211_X1 U5881 ( .C1(n4754), .C2(n6389), .A(n4731), .B(n4730), .ZN(U3026)
         );
  NAND2_X1 U5882 ( .A1(n4747), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4734) );
  OAI22_X1 U5883 ( .A1(n5097), .A2(n4749), .B1(n4748), .B2(n5370), .ZN(n4732)
         );
  AOI21_X1 U5884 ( .B1(n6358), .B2(n4751), .A(n4732), .ZN(n4733) );
  OAI211_X1 U5885 ( .C1(n4754), .C2(n6361), .A(n4734), .B(n4733), .ZN(U3020)
         );
  NAND2_X1 U5886 ( .A1(n4747), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4737) );
  OAI22_X1 U5887 ( .A1(n5079), .A2(n4749), .B1(n4748), .B2(n5351), .ZN(n4735)
         );
  AOI21_X1 U5888 ( .B1(n6378), .B2(n4751), .A(n4735), .ZN(n4736) );
  OAI211_X1 U5889 ( .C1(n4754), .C2(n6381), .A(n4737), .B(n4736), .ZN(U3024)
         );
  NAND2_X1 U5890 ( .A1(n4747), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4740) );
  OAI22_X1 U5891 ( .A1(n5108), .A2(n4749), .B1(n4748), .B2(n5359), .ZN(n4738)
         );
  AOI21_X1 U5892 ( .B1(n6368), .B2(n4751), .A(n4738), .ZN(n4739) );
  OAI211_X1 U5893 ( .C1(n4754), .C2(n6371), .A(n4740), .B(n4739), .ZN(U3022)
         );
  NAND2_X1 U5894 ( .A1(n4747), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4743) );
  OAI22_X1 U5895 ( .A1(n5085), .A2(n4749), .B1(n4748), .B2(n5355), .ZN(n4741)
         );
  AOI21_X1 U5896 ( .B1(n6393), .B2(n4751), .A(n4741), .ZN(n4742) );
  OAI211_X1 U5897 ( .C1(n4754), .C2(n6397), .A(n4743), .B(n4742), .ZN(U3027)
         );
  NAND2_X1 U5898 ( .A1(n4747), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4746) );
  OAI22_X1 U5899 ( .A1(n5075), .A2(n4749), .B1(n4748), .B2(n5343), .ZN(n4744)
         );
  AOI21_X1 U5900 ( .B1(n6372), .B2(n4751), .A(n4744), .ZN(n4745) );
  OAI211_X1 U5901 ( .C1(n4754), .C2(n6375), .A(n4746), .B(n4745), .ZN(U3023)
         );
  NAND2_X1 U5902 ( .A1(n4747), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4753) );
  OAI22_X1 U5903 ( .A1(n5101), .A2(n4749), .B1(n4748), .B2(n5339), .ZN(n4750)
         );
  AOI21_X1 U5904 ( .B1(n6362), .B2(n4751), .A(n4750), .ZN(n4752) );
  OAI211_X1 U5905 ( .C1(n4754), .C2(n6365), .A(n4753), .B(n4752), .ZN(U3021)
         );
  OAI222_X1 U5906 ( .A1(n6174), .A2(n5608), .B1(n6195), .B2(n3624), .C1(n4755), 
        .C2(n5610), .ZN(U2855) );
  INV_X1 U5907 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6227) );
  OAI222_X1 U5908 ( .A1(n6152), .A2(n5626), .B1(n4757), .B2(n4756), .C1(n5613), 
        .C2(n6227), .ZN(U2885) );
  NAND3_X1 U5909 ( .A1(n4759), .A2(n5859), .A3(n4758), .ZN(n4760) );
  NAND2_X1 U5910 ( .A1(n4760), .A2(n6350), .ZN(n4768) );
  INV_X1 U5911 ( .A(n4768), .ZN(n4766) );
  NAND2_X1 U5912 ( .A1(n5877), .A2(n4761), .ZN(n5015) );
  OR2_X1 U5913 ( .A1(n5015), .A2(n5204), .ZN(n4764) );
  INV_X1 U5914 ( .A(n4762), .ZN(n4763) );
  NAND2_X1 U5915 ( .A1(n4763), .A2(n6357), .ZN(n4796) );
  NAND2_X1 U5916 ( .A1(n4764), .A2(n4796), .ZN(n4769) );
  NAND3_X1 U5917 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6357), .A3(n6458), .ZN(n5012) );
  INV_X1 U5918 ( .A(n5012), .ZN(n4765) );
  AOI22_X1 U5919 ( .A1(n4766), .A2(n4769), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4765), .ZN(n4800) );
  AOI21_X1 U5920 ( .B1(n5012), .B2(n6347), .A(n4933), .ZN(n4767) );
  OAI21_X1 U5921 ( .B1(n4769), .B2(n4768), .A(n4767), .ZN(n4795) );
  NAND2_X1 U5922 ( .A1(n4795), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4776) );
  OR3_X1 U5923 ( .A1(n4773), .A2(n5860), .A3(n4770), .ZN(n4771) );
  OAI22_X1 U5924 ( .A1(n5108), .A2(n4796), .B1(n6371), .B2(n5881), .ZN(n4774)
         );
  AOI21_X1 U5925 ( .B1(n6368), .B2(n5043), .A(n4774), .ZN(n4775) );
  OAI211_X1 U5926 ( .C1(n4800), .C2(n5359), .A(n4776), .B(n4775), .ZN(U3046)
         );
  NAND2_X1 U5927 ( .A1(n4795), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4779) );
  OAI22_X1 U5928 ( .A1(n5085), .A2(n4796), .B1(n6397), .B2(n5881), .ZN(n4777)
         );
  AOI21_X1 U5929 ( .B1(n6393), .B2(n5043), .A(n4777), .ZN(n4778) );
  OAI211_X1 U5930 ( .C1(n4800), .C2(n5355), .A(n4779), .B(n4778), .ZN(U3051)
         );
  NAND2_X1 U5931 ( .A1(n4795), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4782) );
  OAI22_X1 U5932 ( .A1(n5075), .A2(n4796), .B1(n6375), .B2(n5881), .ZN(n4780)
         );
  AOI21_X1 U5933 ( .B1(n6372), .B2(n5043), .A(n4780), .ZN(n4781) );
  OAI211_X1 U5934 ( .C1(n4800), .C2(n5343), .A(n4782), .B(n4781), .ZN(U3047)
         );
  NAND2_X1 U5935 ( .A1(n4795), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4785) );
  OAI22_X1 U5936 ( .A1(n5089), .A2(n4796), .B1(n6389), .B2(n5881), .ZN(n4783)
         );
  AOI21_X1 U5937 ( .B1(n6386), .B2(n5043), .A(n4783), .ZN(n4784) );
  OAI211_X1 U5938 ( .C1(n4800), .C2(n5347), .A(n4785), .B(n4784), .ZN(U3050)
         );
  NAND2_X1 U5939 ( .A1(n4795), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4788) );
  OAI22_X1 U5940 ( .A1(n5079), .A2(n4796), .B1(n6381), .B2(n5881), .ZN(n4786)
         );
  AOI21_X1 U5941 ( .B1(n6378), .B2(n5043), .A(n4786), .ZN(n4787) );
  OAI211_X1 U5942 ( .C1(n4800), .C2(n5351), .A(n4788), .B(n4787), .ZN(U3048)
         );
  NAND2_X1 U5943 ( .A1(n4795), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4791) );
  OAI22_X1 U5944 ( .A1(n5097), .A2(n4796), .B1(n6361), .B2(n5881), .ZN(n4789)
         );
  AOI21_X1 U5945 ( .B1(n6358), .B2(n5043), .A(n4789), .ZN(n4790) );
  OAI211_X1 U5946 ( .C1(n4800), .C2(n5370), .A(n4791), .B(n4790), .ZN(U3044)
         );
  NAND2_X1 U5947 ( .A1(n4795), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4794) );
  OAI22_X1 U5948 ( .A1(n5101), .A2(n4796), .B1(n6365), .B2(n5881), .ZN(n4792)
         );
  AOI21_X1 U5949 ( .B1(n6362), .B2(n5043), .A(n4792), .ZN(n4793) );
  OAI211_X1 U5950 ( .C1(n4800), .C2(n5339), .A(n4794), .B(n4793), .ZN(U3045)
         );
  NAND2_X1 U5951 ( .A1(n4795), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4799) );
  OAI22_X1 U5952 ( .A1(n5093), .A2(n4796), .B1(n6385), .B2(n5881), .ZN(n4797)
         );
  AOI21_X1 U5953 ( .B1(n6382), .B2(n5043), .A(n4797), .ZN(n4798) );
  OAI211_X1 U5954 ( .C1(n4800), .C2(n5363), .A(n4799), .B(n4798), .ZN(U3049)
         );
  NAND2_X1 U5955 ( .A1(n5072), .A2(n4801), .ZN(n5872) );
  INV_X1 U5956 ( .A(n5872), .ZN(n4803) );
  NAND2_X1 U5957 ( .A1(n4802), .A2(n6357), .ZN(n5869) );
  NOR2_X1 U5958 ( .A1(n4930), .A2(n5869), .ZN(n4839) );
  AOI21_X1 U5959 ( .B1(n4803), .B2(n3036), .A(n4839), .ZN(n4808) );
  AOI21_X1 U5960 ( .B1(n4811), .B2(STATEBS16_REG_SCAN_IN), .A(n6347), .ZN(
        n5873) );
  INV_X1 U5961 ( .A(n5869), .ZN(n4806) );
  NOR2_X1 U5962 ( .A1(n4806), .A2(n6350), .ZN(n4807) );
  AOI211_X2 U5963 ( .C1(n4808), .C2(n5873), .A(n4807), .B(n4933), .ZN(n4845)
         );
  INV_X1 U5964 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4815) );
  INV_X1 U5965 ( .A(n5873), .ZN(n4809) );
  OAI22_X1 U5966 ( .A1(n4809), .A2(n4808), .B1(n5869), .B2(n4723), .ZN(n4842)
         );
  NAND2_X1 U5967 ( .A1(n4811), .A2(n3815), .ZN(n5913) );
  INV_X1 U5968 ( .A(n6361), .ZN(n6418) );
  AOI22_X1 U5969 ( .A1(n6392), .A2(n6418), .B1(n6417), .B2(n4839), .ZN(n4812)
         );
  OAI21_X1 U5970 ( .B1(n6422), .B2(n5913), .A(n4812), .ZN(n4813) );
  AOI21_X1 U5971 ( .B1(n4842), .B2(n6419), .A(n4813), .ZN(n4814) );
  OAI21_X1 U5972 ( .B1(n4845), .B2(n4815), .A(n4814), .ZN(U3060) );
  AOI22_X1 U5973 ( .A1(n6392), .A2(n6424), .B1(n6423), .B2(n4839), .ZN(n4816)
         );
  OAI21_X1 U5974 ( .B1(n6428), .B2(n5913), .A(n4816), .ZN(n4817) );
  AOI21_X1 U5975 ( .B1(n4842), .B2(n6425), .A(n4817), .ZN(n4818) );
  OAI21_X1 U5976 ( .B1(n4845), .B2(n6720), .A(n4818), .ZN(U3061) );
  INV_X1 U5977 ( .A(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4822) );
  AOI22_X1 U5978 ( .A1(n6392), .A2(n6406), .B1(n6409), .B2(n4839), .ZN(n4819)
         );
  OAI21_X1 U5979 ( .B1(n6416), .B2(n5913), .A(n4819), .ZN(n4820) );
  AOI21_X1 U5980 ( .B1(n4842), .B2(n6411), .A(n4820), .ZN(n4821) );
  OAI21_X1 U5981 ( .B1(n4845), .B2(n4822), .A(n4821), .ZN(U3066) );
  INV_X1 U5982 ( .A(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4826) );
  AOI22_X1 U5983 ( .A1(n6392), .A2(n5081), .B1(n6377), .B2(n4839), .ZN(n4823)
         );
  OAI21_X1 U5984 ( .B1(n5084), .B2(n5913), .A(n4823), .ZN(n4824) );
  AOI21_X1 U5985 ( .B1(n4842), .B2(n6376), .A(n4824), .ZN(n4825) );
  OAI21_X1 U5986 ( .B1(n4845), .B2(n4826), .A(n4825), .ZN(U3064) );
  INV_X1 U5987 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4830) );
  AOI22_X1 U5988 ( .A1(n6392), .A2(n6400), .B1(n6401), .B2(n4839), .ZN(n4827)
         );
  OAI21_X1 U5989 ( .B1(n6405), .B2(n5913), .A(n4827), .ZN(n4828) );
  AOI21_X1 U5990 ( .B1(n4842), .B2(n6402), .A(n4828), .ZN(n4829) );
  OAI21_X1 U5991 ( .B1(n4845), .B2(n4830), .A(n4829), .ZN(U3063) );
  INV_X1 U5992 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4834) );
  AOI22_X1 U5993 ( .A1(n6392), .A2(n5111), .B1(n6367), .B2(n4839), .ZN(n4831)
         );
  OAI21_X1 U5994 ( .B1(n5114), .B2(n5913), .A(n4831), .ZN(n4832) );
  AOI21_X1 U5995 ( .B1(n4842), .B2(n6366), .A(n4832), .ZN(n4833) );
  OAI21_X1 U5996 ( .B1(n4845), .B2(n4834), .A(n4833), .ZN(U3062) );
  INV_X1 U5997 ( .A(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4838) );
  AOI22_X1 U5998 ( .A1(n6392), .A2(n6430), .B1(n6429), .B2(n4839), .ZN(n4835)
         );
  OAI21_X1 U5999 ( .B1(n6434), .B2(n5913), .A(n4835), .ZN(n4836) );
  AOI21_X1 U6000 ( .B1(n4842), .B2(n6431), .A(n4836), .ZN(n4837) );
  OAI21_X1 U6001 ( .B1(n4845), .B2(n4838), .A(n4837), .ZN(U3065) );
  INV_X1 U6002 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4844) );
  AOI22_X1 U6003 ( .A1(n6392), .A2(n6437), .B1(n6436), .B2(n4839), .ZN(n4840)
         );
  OAI21_X1 U6004 ( .B1(n6445), .B2(n5913), .A(n4840), .ZN(n4841) );
  AOI21_X1 U6005 ( .B1(n4842), .B2(n6440), .A(n4841), .ZN(n4843) );
  OAI21_X1 U6006 ( .B1(n4845), .B2(n4844), .A(n4843), .ZN(U3067) );
  INV_X1 U6007 ( .A(n4846), .ZN(n4848) );
  AND2_X1 U6008 ( .A1(n4848), .A2(n4847), .ZN(n4849) );
  NOR2_X1 U6009 ( .A1(n4650), .A2(n4849), .ZN(n6278) );
  INV_X1 U6010 ( .A(n6278), .ZN(n4851) );
  INV_X2 U6011 ( .A(n5613), .ZN(n6205) );
  AOI22_X1 U6012 ( .A1(n5375), .A2(DATAI_5_), .B1(n6205), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n4850) );
  OAI21_X1 U6013 ( .B1(n4851), .B2(n5626), .A(n4850), .ZN(U2886) );
  NAND2_X1 U6014 ( .A1(n4927), .A2(n4490), .ZN(n4859) );
  INV_X1 U6015 ( .A(n4939), .ZN(n4853) );
  NAND3_X1 U6016 ( .A1(n4959), .A2(n6350), .A3(n4891), .ZN(n4854) );
  NAND2_X1 U6017 ( .A1(n4854), .A2(n5009), .ZN(n4858) );
  NAND3_X1 U6018 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6458), .A3(n6453), .ZN(n4936) );
  NOR2_X1 U6019 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4936), .ZN(n4889)
         );
  INV_X1 U6020 ( .A(n6345), .ZN(n4967) );
  OR2_X1 U6021 ( .A1(n6344), .A2(n4855), .ZN(n5073) );
  AOI21_X1 U6022 ( .B1(n5073), .B2(STATE2_REG_2__SCAN_IN), .A(n4856), .ZN(
        n5068) );
  OAI211_X1 U6023 ( .C1(n6567), .C2(n4889), .A(n4967), .B(n5068), .ZN(n4857)
         );
  INV_X1 U6024 ( .A(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4863) );
  INV_X1 U6025 ( .A(n6353), .ZN(n5326) );
  OAI22_X1 U6026 ( .A1(n4859), .A2(n6347), .B1(n5326), .B2(n5073), .ZN(n4888)
         );
  AOI22_X1 U6027 ( .A1(n6423), .A2(n4889), .B1(n6425), .B2(n4888), .ZN(n4860)
         );
  OAI21_X1 U6028 ( .B1(n6428), .B2(n4891), .A(n4860), .ZN(n4861) );
  AOI21_X1 U6029 ( .B1(n4893), .B2(n6424), .A(n4861), .ZN(n4862) );
  OAI21_X1 U6030 ( .B1(n4896), .B2(n4863), .A(n4862), .ZN(U3085) );
  INV_X1 U6031 ( .A(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4867) );
  AOI22_X1 U6032 ( .A1(n6401), .A2(n4889), .B1(n6402), .B2(n4888), .ZN(n4864)
         );
  OAI21_X1 U6033 ( .B1(n6405), .B2(n4891), .A(n4864), .ZN(n4865) );
  AOI21_X1 U6034 ( .B1(n4893), .B2(n6400), .A(n4865), .ZN(n4866) );
  OAI21_X1 U6035 ( .B1(n4896), .B2(n4867), .A(n4866), .ZN(U3087) );
  INV_X1 U6036 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4871) );
  AOI22_X1 U6037 ( .A1(n6367), .A2(n4889), .B1(n6366), .B2(n4888), .ZN(n4868)
         );
  OAI21_X1 U6038 ( .B1(n5114), .B2(n4891), .A(n4868), .ZN(n4869) );
  AOI21_X1 U6039 ( .B1(n4893), .B2(n5111), .A(n4869), .ZN(n4870) );
  OAI21_X1 U6040 ( .B1(n4896), .B2(n4871), .A(n4870), .ZN(U3086) );
  INV_X1 U6041 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4875) );
  AOI22_X1 U6042 ( .A1(n6417), .A2(n4889), .B1(n6419), .B2(n4888), .ZN(n4872)
         );
  OAI21_X1 U6043 ( .B1(n6422), .B2(n4891), .A(n4872), .ZN(n4873) );
  AOI21_X1 U6044 ( .B1(n4893), .B2(n6418), .A(n4873), .ZN(n4874) );
  OAI21_X1 U6045 ( .B1(n4896), .B2(n4875), .A(n4874), .ZN(U3084) );
  INV_X1 U6046 ( .A(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4879) );
  AOI22_X1 U6047 ( .A1(n6409), .A2(n4889), .B1(n6411), .B2(n4888), .ZN(n4876)
         );
  OAI21_X1 U6048 ( .B1(n6416), .B2(n4891), .A(n4876), .ZN(n4877) );
  AOI21_X1 U6049 ( .B1(n4893), .B2(n6406), .A(n4877), .ZN(n4878) );
  OAI21_X1 U6050 ( .B1(n4896), .B2(n4879), .A(n4878), .ZN(U3090) );
  INV_X1 U6051 ( .A(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4883) );
  AOI22_X1 U6052 ( .A1(n6429), .A2(n4889), .B1(n6431), .B2(n4888), .ZN(n4880)
         );
  OAI21_X1 U6053 ( .B1(n6434), .B2(n4891), .A(n4880), .ZN(n4881) );
  AOI21_X1 U6054 ( .B1(n4893), .B2(n6430), .A(n4881), .ZN(n4882) );
  OAI21_X1 U6055 ( .B1(n4896), .B2(n4883), .A(n4882), .ZN(U3089) );
  INV_X1 U6056 ( .A(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4887) );
  AOI22_X1 U6057 ( .A1(n6436), .A2(n4889), .B1(n6440), .B2(n4888), .ZN(n4884)
         );
  OAI21_X1 U6058 ( .B1(n6445), .B2(n4891), .A(n4884), .ZN(n4885) );
  AOI21_X1 U6059 ( .B1(n4893), .B2(n6437), .A(n4885), .ZN(n4886) );
  OAI21_X1 U6060 ( .B1(n4896), .B2(n4887), .A(n4886), .ZN(U3091) );
  INV_X1 U6061 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4895) );
  AOI22_X1 U6062 ( .A1(n6377), .A2(n4889), .B1(n6376), .B2(n4888), .ZN(n4890)
         );
  OAI21_X1 U6063 ( .B1(n5084), .B2(n4891), .A(n4890), .ZN(n4892) );
  AOI21_X1 U6064 ( .B1(n4893), .B2(n5081), .A(n4892), .ZN(n4894) );
  OAI21_X1 U6065 ( .B1(n4896), .B2(n4895), .A(n4894), .ZN(U3088) );
  XNOR2_X1 U6066 ( .A(n4897), .B(n4898), .ZN(n5063) );
  INV_X1 U6067 ( .A(n6329), .ZN(n5985) );
  AND2_X1 U6068 ( .A1(n4902), .A2(n4899), .ZN(n4901) );
  OAI21_X1 U6069 ( .B1(n5985), .B2(n4901), .A(n4900), .ZN(n4917) );
  NAND3_X1 U6070 ( .A1(n4902), .A2(n4908), .A3(n3634), .ZN(n4903) );
  INV_X1 U6071 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6710) );
  OR2_X1 U6072 ( .A1(n6308), .A2(n6710), .ZN(n5058) );
  OAI211_X1 U6073 ( .C1(n6309), .C2(n6146), .A(n4903), .B(n5058), .ZN(n4904)
         );
  AOI21_X1 U6074 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n4917), .A(n4904), 
        .ZN(n4905) );
  OAI21_X1 U6075 ( .B1(n6307), .B2(n5063), .A(n4905), .ZN(U3012) );
  XOR2_X1 U6076 ( .A(n3024), .B(n4907), .Z(n6279) );
  INV_X1 U6077 ( .A(n6279), .ZN(n4920) );
  INV_X1 U6078 ( .A(n4908), .ZN(n5149) );
  OAI21_X1 U6079 ( .B1(n4910), .B2(n5149), .A(n4909), .ZN(n4918) );
  NAND2_X1 U6080 ( .A1(n4912), .A2(n4911), .ZN(n4913) );
  AND2_X1 U6081 ( .A1(n4914), .A2(n4913), .ZN(n6190) );
  INV_X1 U6082 ( .A(n6190), .ZN(n4915) );
  NAND2_X1 U6083 ( .A1(n6334), .A2(REIP_REG_5__SCAN_IN), .ZN(n6280) );
  OAI21_X1 U6084 ( .B1(n6309), .B2(n4915), .A(n6280), .ZN(n4916) );
  AOI21_X1 U6085 ( .B1(n4918), .B2(n4917), .A(n4916), .ZN(n4919) );
  OAI21_X1 U6086 ( .B1(n4920), .B2(n6307), .A(n4919), .ZN(U3013) );
  OR2_X1 U6087 ( .A1(n5049), .A2(n4922), .ZN(n4923) );
  NAND2_X1 U6088 ( .A1(n5118), .A2(n4923), .ZN(n6120) );
  AOI21_X1 U6089 ( .B1(n4924), .B2(n5054), .A(n5137), .ZN(n6320) );
  AOI22_X1 U6090 ( .A1(n6191), .A2(n6320), .B1(EBX_REG_9__SCAN_IN), .B2(n5559), 
        .ZN(n4925) );
  OAI21_X1 U6091 ( .B1(n6120), .B2(n5610), .A(n4925), .ZN(U2850) );
  AOI22_X1 U6092 ( .A1(n5375), .A2(DATAI_9_), .B1(n6205), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4926) );
  OAI21_X1 U6093 ( .B1(n6120), .B2(n5626), .A(n4926), .ZN(U2882) );
  OAI21_X1 U6094 ( .B1(n4939), .B2(n6760), .A(n6350), .ZN(n4937) );
  INV_X1 U6095 ( .A(n4927), .ZN(n4929) );
  OR2_X1 U6096 ( .A1(n4929), .A2(n4928), .ZN(n4932) );
  NOR2_X1 U6097 ( .A1(n4930), .A2(n4936), .ZN(n4956) );
  INV_X1 U6098 ( .A(n4956), .ZN(n4931) );
  AND2_X1 U6099 ( .A1(n4932), .A2(n4931), .ZN(n4938) );
  INV_X1 U6100 ( .A(n4938), .ZN(n4935) );
  AOI21_X1 U6101 ( .B1(n6347), .B2(n4936), .A(n4933), .ZN(n4934) );
  OAI21_X1 U6102 ( .B1(n4937), .B2(n4935), .A(n4934), .ZN(n4955) );
  OAI22_X1 U6103 ( .A1(n4938), .A2(n4937), .B1(n5335), .B2(n4936), .ZN(n4954)
         );
  AOI22_X1 U6104 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4955), .B1(n6376), 
        .B2(n4954), .ZN(n4941) );
  AOI22_X1 U6105 ( .A1(n5368), .A2(n5081), .B1(n4956), .B2(n6377), .ZN(n4940)
         );
  OAI211_X1 U6106 ( .C1(n4959), .C2(n5084), .A(n4941), .B(n4940), .ZN(U3096)
         );
  AOI22_X1 U6107 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4955), .B1(n6440), 
        .B2(n4954), .ZN(n4943) );
  AOI22_X1 U6108 ( .A1(n5368), .A2(n6437), .B1(n4956), .B2(n6436), .ZN(n4942)
         );
  OAI211_X1 U6109 ( .C1(n4959), .C2(n6445), .A(n4943), .B(n4942), .ZN(U3099)
         );
  AOI22_X1 U6110 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4955), .B1(n6411), 
        .B2(n4954), .ZN(n4945) );
  AOI22_X1 U6111 ( .A1(n5368), .A2(n6406), .B1(n4956), .B2(n6409), .ZN(n4944)
         );
  OAI211_X1 U6112 ( .C1(n4959), .C2(n6416), .A(n4945), .B(n4944), .ZN(U3098)
         );
  AOI22_X1 U6113 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4955), .B1(n6402), 
        .B2(n4954), .ZN(n4947) );
  AOI22_X1 U6114 ( .A1(n5368), .A2(n6400), .B1(n4956), .B2(n6401), .ZN(n4946)
         );
  OAI211_X1 U6115 ( .C1(n4959), .C2(n6405), .A(n4947), .B(n4946), .ZN(U3095)
         );
  AOI22_X1 U6116 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4955), .B1(n6366), 
        .B2(n4954), .ZN(n4949) );
  AOI22_X1 U6117 ( .A1(n5368), .A2(n5111), .B1(n4956), .B2(n6367), .ZN(n4948)
         );
  OAI211_X1 U6118 ( .C1(n4959), .C2(n5114), .A(n4949), .B(n4948), .ZN(U3094)
         );
  AOI22_X1 U6119 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4955), .B1(n6431), 
        .B2(n4954), .ZN(n4951) );
  AOI22_X1 U6120 ( .A1(n5368), .A2(n6430), .B1(n4956), .B2(n6429), .ZN(n4950)
         );
  OAI211_X1 U6121 ( .C1(n4959), .C2(n6434), .A(n4951), .B(n4950), .ZN(U3097)
         );
  AOI22_X1 U6122 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4955), .B1(n6419), 
        .B2(n4954), .ZN(n4953) );
  AOI22_X1 U6123 ( .A1(n5368), .A2(n6418), .B1(n6417), .B2(n4956), .ZN(n4952)
         );
  OAI211_X1 U6124 ( .C1(n4959), .C2(n6422), .A(n4953), .B(n4952), .ZN(U3092)
         );
  AOI22_X1 U6125 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4955), .B1(n6425), 
        .B2(n4954), .ZN(n4958) );
  AOI22_X1 U6126 ( .A1(n5368), .A2(n6424), .B1(n4956), .B2(n6423), .ZN(n4957)
         );
  OAI211_X1 U6127 ( .C1(n4959), .C2(n6428), .A(n4958), .B(n4957), .ZN(U3093)
         );
  NOR2_X1 U6128 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4960), .ZN(n4970)
         );
  OAI21_X1 U6129 ( .B1(n6344), .B2(n5335), .A(n4961), .ZN(n6352) );
  NOR3_X1 U6130 ( .A1(n6352), .A2(n6357), .A3(n6353), .ZN(n4965) );
  INV_X1 U6131 ( .A(n4999), .ZN(n4962) );
  OAI21_X1 U6132 ( .B1(n4962), .B2(n4996), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4963) );
  NAND3_X1 U6133 ( .A1(n4966), .A2(n6350), .A3(n4963), .ZN(n4964) );
  OAI211_X1 U6134 ( .C1(n4970), .C2(n6567), .A(n4965), .B(n4964), .ZN(n4992)
         );
  NAND2_X1 U6135 ( .A1(n4992), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4973)
         );
  INV_X1 U6136 ( .A(n6344), .ZN(n4968) );
  OAI33_X1 U6137 ( .A1(n4968), .A2(n6357), .A3(n4967), .B1(n4966), .B2(n6347), 
        .B3(n5877), .ZN(n4969) );
  INV_X1 U6138 ( .A(n4969), .ZN(n4994) );
  INV_X1 U6139 ( .A(n4970), .ZN(n4993) );
  OAI22_X1 U6140 ( .A1(n4994), .A2(n5359), .B1(n5108), .B2(n4993), .ZN(n4971)
         );
  AOI21_X1 U6141 ( .B1(n5111), .B2(n4996), .A(n4971), .ZN(n4972) );
  OAI211_X1 U6142 ( .C1(n4999), .C2(n5114), .A(n4973), .B(n4972), .ZN(U3134)
         );
  NAND2_X1 U6143 ( .A1(n4992), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4976)
         );
  OAI22_X1 U6144 ( .A1(n4994), .A2(n5347), .B1(n5089), .B2(n4993), .ZN(n4974)
         );
  AOI21_X1 U6145 ( .B1(n6406), .B2(n4996), .A(n4974), .ZN(n4975) );
  OAI211_X1 U6146 ( .C1(n4999), .C2(n6416), .A(n4976), .B(n4975), .ZN(U3138)
         );
  NAND2_X1 U6147 ( .A1(n4992), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4979)
         );
  OAI22_X1 U6148 ( .A1(n4994), .A2(n5351), .B1(n5079), .B2(n4993), .ZN(n4977)
         );
  AOI21_X1 U6149 ( .B1(n5081), .B2(n4996), .A(n4977), .ZN(n4978) );
  OAI211_X1 U6150 ( .C1(n4999), .C2(n5084), .A(n4979), .B(n4978), .ZN(U3136)
         );
  NAND2_X1 U6151 ( .A1(n4992), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4982)
         );
  OAI22_X1 U6152 ( .A1(n4994), .A2(n5363), .B1(n5093), .B2(n4993), .ZN(n4980)
         );
  AOI21_X1 U6153 ( .B1(n6430), .B2(n4996), .A(n4980), .ZN(n4981) );
  OAI211_X1 U6154 ( .C1(n4999), .C2(n6434), .A(n4982), .B(n4981), .ZN(U3137)
         );
  NAND2_X1 U6155 ( .A1(n4992), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4985)
         );
  OAI22_X1 U6156 ( .A1(n4994), .A2(n5355), .B1(n5085), .B2(n4993), .ZN(n4983)
         );
  AOI21_X1 U6157 ( .B1(n6437), .B2(n4996), .A(n4983), .ZN(n4984) );
  OAI211_X1 U6158 ( .C1(n4999), .C2(n6445), .A(n4985), .B(n4984), .ZN(U3139)
         );
  NAND2_X1 U6159 ( .A1(n4992), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4988)
         );
  OAI22_X1 U6160 ( .A1(n4994), .A2(n5343), .B1(n5075), .B2(n4993), .ZN(n4986)
         );
  AOI21_X1 U6161 ( .B1(n6400), .B2(n4996), .A(n4986), .ZN(n4987) );
  OAI211_X1 U6162 ( .C1(n4999), .C2(n6405), .A(n4988), .B(n4987), .ZN(U3135)
         );
  NAND2_X1 U6163 ( .A1(n4992), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4991)
         );
  OAI22_X1 U6164 ( .A1(n4994), .A2(n5370), .B1(n5097), .B2(n4993), .ZN(n4989)
         );
  AOI21_X1 U6165 ( .B1(n6418), .B2(n4996), .A(n4989), .ZN(n4990) );
  OAI211_X1 U6166 ( .C1(n4999), .C2(n6422), .A(n4991), .B(n4990), .ZN(U3132)
         );
  NAND2_X1 U6167 ( .A1(n4992), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4998)
         );
  OAI22_X1 U6168 ( .A1(n4994), .A2(n5339), .B1(n5101), .B2(n4993), .ZN(n4995)
         );
  AOI21_X1 U6169 ( .B1(n6424), .B2(n4996), .A(n4995), .ZN(n4997) );
  OAI211_X1 U6170 ( .C1(n4999), .C2(n6428), .A(n4998), .B(n4997), .ZN(U3133)
         );
  INV_X1 U6171 ( .A(n5000), .ZN(n5001) );
  AOI21_X1 U6172 ( .B1(n5002), .B2(n4651), .A(n5001), .ZN(n6271) );
  INV_X1 U6173 ( .A(n6271), .ZN(n5008) );
  AOI22_X1 U6174 ( .A1(n5375), .A2(DATAI_7_), .B1(n6205), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n5003) );
  OAI21_X1 U6175 ( .B1(n5008), .B2(n5626), .A(n5003), .ZN(U2884) );
  INV_X1 U6176 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5007) );
  OR2_X1 U6177 ( .A1(n5005), .A2(n5004), .ZN(n5006) );
  NAND2_X1 U6178 ( .A1(n5052), .A2(n5006), .ZN(n6140) );
  OAI222_X1 U6179 ( .A1(n5008), .A2(n5610), .B1(n5007), .B2(n6195), .C1(n5608), 
        .C2(n6140), .ZN(U2852) );
  INV_X1 U6180 ( .A(n5046), .ZN(n5010) );
  OAI21_X1 U6181 ( .B1(n5010), .B2(n5043), .A(n5009), .ZN(n5011) );
  AOI21_X1 U6182 ( .B1(n5011), .B2(n5015), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5013) );
  NOR2_X1 U6183 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5012), .ZN(n5014)
         );
  NOR2_X1 U6184 ( .A1(n6345), .A2(n6352), .ZN(n5334) );
  NAND2_X1 U6185 ( .A1(n5039), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n5020) );
  INV_X1 U6186 ( .A(n5014), .ZN(n5041) );
  INV_X1 U6187 ( .A(n5015), .ZN(n5017) );
  NOR2_X1 U6188 ( .A1(n5326), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5016)
         );
  AOI22_X1 U6189 ( .A1(n5017), .A2(n6350), .B1(n6344), .B2(n5016), .ZN(n5040)
         );
  OAI22_X1 U6190 ( .A1(n5097), .A2(n5041), .B1(n5040), .B2(n5370), .ZN(n5018)
         );
  AOI21_X1 U6191 ( .B1(n6418), .B2(n5043), .A(n5018), .ZN(n5019) );
  OAI211_X1 U6192 ( .C1(n5046), .C2(n6422), .A(n5020), .B(n5019), .ZN(U3036)
         );
  NAND2_X1 U6193 ( .A1(n5039), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n5023) );
  OAI22_X1 U6194 ( .A1(n5085), .A2(n5041), .B1(n5040), .B2(n5355), .ZN(n5021)
         );
  AOI21_X1 U6195 ( .B1(n6437), .B2(n5043), .A(n5021), .ZN(n5022) );
  OAI211_X1 U6196 ( .C1(n5046), .C2(n6445), .A(n5023), .B(n5022), .ZN(U3043)
         );
  NAND2_X1 U6197 ( .A1(n5039), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n5026) );
  OAI22_X1 U6198 ( .A1(n5089), .A2(n5041), .B1(n5040), .B2(n5347), .ZN(n5024)
         );
  AOI21_X1 U6199 ( .B1(n6406), .B2(n5043), .A(n5024), .ZN(n5025) );
  OAI211_X1 U6200 ( .C1(n5046), .C2(n6416), .A(n5026), .B(n5025), .ZN(U3042)
         );
  NAND2_X1 U6201 ( .A1(n5039), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n5029) );
  OAI22_X1 U6202 ( .A1(n5093), .A2(n5041), .B1(n5040), .B2(n5363), .ZN(n5027)
         );
  AOI21_X1 U6203 ( .B1(n6430), .B2(n5043), .A(n5027), .ZN(n5028) );
  OAI211_X1 U6204 ( .C1(n5046), .C2(n6434), .A(n5029), .B(n5028), .ZN(U3041)
         );
  NAND2_X1 U6205 ( .A1(n5039), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5032) );
  OAI22_X1 U6206 ( .A1(n5108), .A2(n5041), .B1(n5040), .B2(n5359), .ZN(n5030)
         );
  AOI21_X1 U6207 ( .B1(n5111), .B2(n5043), .A(n5030), .ZN(n5031) );
  OAI211_X1 U6208 ( .C1(n5046), .C2(n5114), .A(n5032), .B(n5031), .ZN(U3038)
         );
  NAND2_X1 U6209 ( .A1(n5039), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n5035) );
  OAI22_X1 U6210 ( .A1(n5101), .A2(n5041), .B1(n5040), .B2(n5339), .ZN(n5033)
         );
  AOI21_X1 U6211 ( .B1(n6424), .B2(n5043), .A(n5033), .ZN(n5034) );
  OAI211_X1 U6212 ( .C1(n5046), .C2(n6428), .A(n5035), .B(n5034), .ZN(U3037)
         );
  NAND2_X1 U6213 ( .A1(n5039), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n5038) );
  OAI22_X1 U6214 ( .A1(n5079), .A2(n5041), .B1(n5040), .B2(n5351), .ZN(n5036)
         );
  AOI21_X1 U6215 ( .B1(n5081), .B2(n5043), .A(n5036), .ZN(n5037) );
  OAI211_X1 U6216 ( .C1(n5046), .C2(n5084), .A(n5038), .B(n5037), .ZN(U3040)
         );
  NAND2_X1 U6217 ( .A1(n5039), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n5045) );
  OAI22_X1 U6218 ( .A1(n5075), .A2(n5041), .B1(n5040), .B2(n5343), .ZN(n5042)
         );
  AOI21_X1 U6219 ( .B1(n6400), .B2(n5043), .A(n5042), .ZN(n5044) );
  OAI211_X1 U6220 ( .C1(n5046), .C2(n6405), .A(n5045), .B(n5044), .ZN(U3039)
         );
  AND2_X1 U6221 ( .A1(n5000), .A2(n5047), .ZN(n5048) );
  NOR2_X1 U6222 ( .A1(n5049), .A2(n5048), .ZN(n6130) );
  INV_X1 U6223 ( .A(n6130), .ZN(n5057) );
  AOI22_X1 U6224 ( .A1(n5375), .A2(DATAI_8_), .B1(n6205), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n5050) );
  OAI21_X1 U6225 ( .B1(n5057), .B2(n5626), .A(n5050), .ZN(U2883) );
  NAND2_X1 U6226 ( .A1(n5052), .A2(n5051), .ZN(n5053) );
  NAND2_X1 U6227 ( .A1(n5054), .A2(n5053), .ZN(n6125) );
  INV_X1 U6228 ( .A(n6125), .ZN(n5055) );
  AOI22_X1 U6229 ( .A1(n6191), .A2(n5055), .B1(EBX_REG_8__SCAN_IN), .B2(n5559), 
        .ZN(n5056) );
  OAI21_X1 U6230 ( .B1(n5057), .B2(n5610), .A(n5056), .ZN(U2851) );
  OAI21_X1 U6231 ( .B1(n6282), .B2(n5059), .A(n5058), .ZN(n5061) );
  NOR2_X1 U6232 ( .A1(n6152), .A2(n6303), .ZN(n5060) );
  AOI211_X1 U6233 ( .C1(n6276), .C2(n6149), .A(n5061), .B(n5060), .ZN(n5062)
         );
  OAI21_X1 U6234 ( .B1(n6297), .B2(n5063), .A(n5062), .ZN(U2980) );
  INV_X1 U6235 ( .A(n5110), .ZN(n5064) );
  AOI21_X1 U6236 ( .B1(n5064), .B2(n5115), .A(n6760), .ZN(n5065) );
  AOI211_X1 U6237 ( .C1(n5072), .C2(n5066), .A(n6347), .B(n5065), .ZN(n5070)
         );
  NOR2_X1 U6238 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5067), .ZN(n5071)
         );
  OAI211_X1 U6239 ( .C1(n6567), .C2(n5071), .A(n5326), .B(n5068), .ZN(n5069)
         );
  NAND2_X1 U6240 ( .A1(n5105), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n5078)
         );
  INV_X1 U6241 ( .A(n5071), .ZN(n5107) );
  AND2_X1 U6242 ( .A1(n5072), .A2(n6350), .ZN(n5878) );
  INV_X1 U6243 ( .A(n5073), .ZN(n5074) );
  AOI22_X1 U6244 ( .A1(n5878), .A2(n4490), .B1(n6345), .B2(n5074), .ZN(n5106)
         );
  OAI22_X1 U6245 ( .A1(n5075), .A2(n5107), .B1(n5106), .B2(n5343), .ZN(n5076)
         );
  AOI21_X1 U6246 ( .B1(n6400), .B2(n5110), .A(n5076), .ZN(n5077) );
  OAI211_X1 U6247 ( .C1(n5115), .C2(n6405), .A(n5078), .B(n5077), .ZN(U3119)
         );
  NAND2_X1 U6248 ( .A1(n5105), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5083)
         );
  OAI22_X1 U6249 ( .A1(n5079), .A2(n5107), .B1(n5106), .B2(n5351), .ZN(n5080)
         );
  AOI21_X1 U6250 ( .B1(n5081), .B2(n5110), .A(n5080), .ZN(n5082) );
  OAI211_X1 U6251 ( .C1(n5115), .C2(n5084), .A(n5083), .B(n5082), .ZN(U3120)
         );
  NAND2_X1 U6252 ( .A1(n5105), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n5088)
         );
  OAI22_X1 U6253 ( .A1(n5085), .A2(n5107), .B1(n5106), .B2(n5355), .ZN(n5086)
         );
  AOI21_X1 U6254 ( .B1(n6437), .B2(n5110), .A(n5086), .ZN(n5087) );
  OAI211_X1 U6255 ( .C1(n5115), .C2(n6445), .A(n5088), .B(n5087), .ZN(U3123)
         );
  NAND2_X1 U6256 ( .A1(n5105), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n5092)
         );
  OAI22_X1 U6257 ( .A1(n5089), .A2(n5107), .B1(n5106), .B2(n5347), .ZN(n5090)
         );
  AOI21_X1 U6258 ( .B1(n6406), .B2(n5110), .A(n5090), .ZN(n5091) );
  OAI211_X1 U6259 ( .C1(n5115), .C2(n6416), .A(n5092), .B(n5091), .ZN(U3122)
         );
  NAND2_X1 U6260 ( .A1(n5105), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n5096)
         );
  OAI22_X1 U6261 ( .A1(n5093), .A2(n5107), .B1(n5106), .B2(n5363), .ZN(n5094)
         );
  AOI21_X1 U6262 ( .B1(n6430), .B2(n5110), .A(n5094), .ZN(n5095) );
  OAI211_X1 U6263 ( .C1(n5115), .C2(n6434), .A(n5096), .B(n5095), .ZN(U3121)
         );
  NAND2_X1 U6264 ( .A1(n5105), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n5100)
         );
  OAI22_X1 U6265 ( .A1(n5097), .A2(n5107), .B1(n5106), .B2(n5370), .ZN(n5098)
         );
  AOI21_X1 U6266 ( .B1(n6418), .B2(n5110), .A(n5098), .ZN(n5099) );
  OAI211_X1 U6267 ( .C1(n5115), .C2(n6422), .A(n5100), .B(n5099), .ZN(U3116)
         );
  NAND2_X1 U6268 ( .A1(n5105), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n5104)
         );
  OAI22_X1 U6269 ( .A1(n5101), .A2(n5107), .B1(n5106), .B2(n5339), .ZN(n5102)
         );
  AOI21_X1 U6270 ( .B1(n6424), .B2(n5110), .A(n5102), .ZN(n5103) );
  OAI211_X1 U6271 ( .C1(n5115), .C2(n6428), .A(n5104), .B(n5103), .ZN(U3117)
         );
  NAND2_X1 U6272 ( .A1(n5105), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n5113)
         );
  OAI22_X1 U6273 ( .A1(n5108), .A2(n5107), .B1(n5106), .B2(n5359), .ZN(n5109)
         );
  AOI21_X1 U6274 ( .B1(n5111), .B2(n5110), .A(n5109), .ZN(n5112) );
  OAI211_X1 U6275 ( .C1(n5115), .C2(n5114), .A(n5113), .B(n5112), .ZN(U3118)
         );
  INV_X1 U6276 ( .A(n5116), .ZN(n5117) );
  AOI21_X1 U6277 ( .B1(n5119), .B2(n5118), .A(n5117), .ZN(n5218) );
  INV_X1 U6278 ( .A(n5218), .ZN(n5168) );
  AOI22_X1 U6279 ( .A1(n5375), .A2(DATAI_10_), .B1(n6205), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n5120) );
  OAI21_X1 U6280 ( .B1(n5168), .B2(n5626), .A(n5120), .ZN(U2881) );
  NOR3_X1 U6281 ( .A1(n6479), .A2(n6567), .A3(n5121), .ZN(n6475) );
  NAND2_X1 U6282 ( .A1(n6479), .A2(n4723), .ZN(n6492) );
  NOR3_X1 U6283 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6492), .A3(n6474), .ZN(
        n6488) );
  OR2_X1 U6284 ( .A1(n6284), .A2(n6488), .ZN(n5122) );
  OR2_X1 U6285 ( .A1(n6475), .A2(n5122), .ZN(n5123) );
  INV_X1 U6286 ( .A(n5132), .ZN(n5124) );
  NAND2_X1 U6287 ( .A1(n5124), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5125) );
  NAND3_X1 U6288 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .A3(
        REIP_REG_7__SCAN_IN), .ZN(n6112) );
  INV_X1 U6289 ( .A(n6112), .ZN(n5130) );
  NAND3_X1 U6290 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6184) );
  NOR2_X1 U6291 ( .A1(n6517), .A2(n6184), .ZN(n6163) );
  NAND2_X1 U6292 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6163), .ZN(n5383) );
  NOR2_X1 U6293 ( .A1(n5384), .A2(n5383), .ZN(n6137) );
  NAND2_X1 U6294 ( .A1(n4307), .A2(n6760), .ZN(n5141) );
  INV_X1 U6295 ( .A(n5141), .ZN(n5126) );
  AND3_X1 U6296 ( .A1(n5127), .A2(n3606), .A3(n5126), .ZN(n5128) );
  INV_X1 U6297 ( .A(n5384), .ZN(n5129) );
  NAND2_X1 U6298 ( .A1(n6185), .A2(n5129), .ZN(n5547) );
  AOI21_X1 U6299 ( .B1(n5130), .B2(n6137), .A(n6138), .ZN(n6124) );
  INV_X1 U6300 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6722) );
  INV_X1 U6301 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6525) );
  OR2_X1 U6302 ( .A1(n6185), .A2(n5383), .ZN(n6135) );
  AOI211_X1 U6303 ( .C1(n6722), .C2(n6525), .A(n6112), .B(n6135), .ZN(n5131)
         );
  NAND2_X1 U6304 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .ZN(
        n5221) );
  AOI22_X1 U6305 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6124), .B1(n5131), .B2(
        n5221), .ZN(n5148) );
  NAND2_X1 U6306 ( .A1(n5132), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5133) );
  INV_X1 U6307 ( .A(n5216), .ZN(n5146) );
  NAND3_X1 U6308 ( .A1(n5134), .A2(EBX_REG_31__SCAN_IN), .A3(n5141), .ZN(n5135) );
  NOR2_X2 U6309 ( .A1(n5180), .A2(n5135), .ZN(n6158) );
  NOR2_X1 U6310 ( .A1(n5137), .A2(n5136), .ZN(n5138) );
  OR2_X1 U6311 ( .A1(n5195), .A2(n5138), .ZN(n6310) );
  OR2_X1 U6312 ( .A1(n6501), .A2(n5141), .ZN(n6471) );
  NAND2_X1 U6313 ( .A1(n5139), .A2(n6471), .ZN(n5140) );
  NOR2_X1 U6314 ( .A1(n5180), .A2(n5140), .ZN(n5464) );
  INV_X1 U6315 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5554) );
  NAND3_X1 U6316 ( .A1(n3606), .A2(n5141), .A3(n5554), .ZN(n5142) );
  NOR2_X1 U6317 ( .A1(n5180), .A2(n5142), .ZN(n5143) );
  AOI22_X1 U6318 ( .A1(EBX_REG_10__SCAN_IN), .A2(n6172), .B1(
        PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n6178), .ZN(n5144) );
  NOR2_X1 U6319 ( .A1(n6033), .A2(n5384), .ZN(n6177) );
  OAI211_X1 U6320 ( .C1(n6175), .C2(n6310), .A(n5144), .B(n6160), .ZN(n5145)
         );
  AOI21_X1 U6321 ( .B1(n6180), .B2(n5146), .A(n5145), .ZN(n5147) );
  OAI211_X1 U6322 ( .C1(n5168), .C2(n6151), .A(n5148), .B(n5147), .ZN(U2817)
         );
  XOR2_X1 U6323 ( .A(n5151), .B(n5152), .Z(n6272) );
  NAND2_X1 U6324 ( .A1(n6272), .A2(n6322), .ZN(n5162) );
  INV_X1 U6325 ( .A(n5153), .ZN(n5158) );
  OAI21_X1 U6326 ( .B1(n5156), .B2(n5155), .A(n5154), .ZN(n5157) );
  AOI21_X1 U6327 ( .B1(n5159), .B2(n5158), .A(n5157), .ZN(n5259) );
  INV_X1 U6328 ( .A(n5259), .ZN(n6305) );
  NAND2_X1 U6329 ( .A1(n6334), .A2(REIP_REG_7__SCAN_IN), .ZN(n6273) );
  OAI21_X1 U6330 ( .B1(n6309), .B2(n6140), .A(n6273), .ZN(n5160) );
  AOI21_X1 U6331 ( .B1(n6305), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n5160), 
        .ZN(n5161) );
  OAI211_X1 U6332 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n6312), .A(n5162), 
        .B(n5161), .ZN(U3011) );
  XNOR2_X1 U6333 ( .A(n5163), .B(n5164), .ZN(n5174) );
  NAND2_X1 U6334 ( .A1(n6334), .A2(REIP_REG_8__SCAN_IN), .ZN(n5169) );
  NAND2_X1 U6335 ( .A1(n6300), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5165)
         );
  OAI211_X1 U6336 ( .C1(n6294), .C2(n6128), .A(n5169), .B(n5165), .ZN(n5166)
         );
  AOI21_X1 U6337 ( .B1(n6130), .B2(n6287), .A(n5166), .ZN(n5167) );
  OAI21_X1 U6338 ( .B1(n5174), .B2(n6297), .A(n5167), .ZN(U2978) );
  OAI222_X1 U6339 ( .A1(n5168), .A2(n5610), .B1(n6195), .B2(n3648), .C1(n6310), 
        .C2(n5608), .ZN(U2849) );
  OAI21_X1 U6340 ( .B1(n6309), .B2(n6125), .A(n5169), .ZN(n5172) );
  OAI21_X1 U6341 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6313), .ZN(n5170) );
  NOR2_X1 U6342 ( .A1(n6312), .A2(n5170), .ZN(n5171) );
  AOI211_X1 U6343 ( .C1(INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n6305), .A(n5172), 
        .B(n5171), .ZN(n5173) );
  OAI21_X1 U6344 ( .B1(n6307), .B2(n5174), .A(n5173), .ZN(U3010) );
  NAND2_X1 U6345 ( .A1(n5175), .A2(n3543), .ZN(n5176) );
  OAI21_X1 U6346 ( .B1(n5384), .B2(n5251), .A(n5547), .ZN(n5177) );
  NAND2_X1 U6347 ( .A1(n5177), .A2(REIP_REG_2__SCAN_IN), .ZN(n5240) );
  OAI21_X1 U6348 ( .B1(n6185), .B2(n5251), .A(n4415), .ZN(n5178) );
  NAND2_X1 U6349 ( .A1(n5240), .A2(n5178), .ZN(n5188) );
  NOR2_X1 U6350 ( .A1(n5180), .A2(n5179), .ZN(n6170) );
  INV_X1 U6351 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5181) );
  OAI22_X1 U6352 ( .A1(n6293), .A2(n6161), .B1(n6115), .B2(n5181), .ZN(n5182)
         );
  AOI21_X1 U6353 ( .B1(n6170), .B2(n5183), .A(n5182), .ZN(n5187) );
  NAND2_X1 U6354 ( .A1(n6172), .A2(EBX_REG_2__SCAN_IN), .ZN(n5186) );
  NAND2_X1 U6355 ( .A1(n6158), .A2(n5184), .ZN(n5185) );
  AND4_X1 U6356 ( .A1(n5188), .A2(n5187), .A3(n5186), .A4(n5185), .ZN(n5189)
         );
  OAI21_X1 U6357 ( .B1(n6157), .B2(n6286), .A(n5189), .ZN(U2825) );
  AND2_X1 U6358 ( .A1(n5116), .A2(n5190), .ZN(n5192) );
  OR2_X1 U6359 ( .A1(n5192), .A2(n5191), .ZN(n6105) );
  AOI22_X1 U6360 ( .A1(n5375), .A2(DATAI_11_), .B1(n6205), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5193) );
  OAI21_X1 U6361 ( .B1(n6105), .B2(n5626), .A(n5193), .ZN(U2880) );
  INV_X1 U6362 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5196) );
  OAI21_X1 U6363 ( .B1(n5195), .B2(n5194), .A(n5224), .ZN(n5262) );
  OAI222_X1 U6364 ( .A1(n6105), .A2(n5610), .B1(n5196), .B2(n6195), .C1(n5608), 
        .C2(n5262), .ZN(U2848) );
  XNOR2_X1 U6365 ( .A(n5727), .B(n6326), .ZN(n5198) );
  XNOR2_X1 U6366 ( .A(n5197), .B(n5198), .ZN(n6323) );
  NAND2_X1 U6367 ( .A1(n6323), .A2(n6289), .ZN(n5201) );
  NAND2_X1 U6368 ( .A1(n6334), .A2(REIP_REG_9__SCAN_IN), .ZN(n6318) );
  OAI21_X1 U6369 ( .B1(n6282), .B2(n6114), .A(n6318), .ZN(n5199) );
  AOI21_X1 U6370 ( .B1(n6276), .B2(n6118), .A(n5199), .ZN(n5200) );
  OAI211_X1 U6371 ( .C1(n6303), .C2(n6120), .A(n5201), .B(n5200), .ZN(U2977)
         );
  INV_X1 U6372 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6582) );
  OAI22_X1 U6373 ( .A1(n6138), .A2(n6582), .B1(n6169), .B2(n5202), .ZN(n5209)
         );
  INV_X1 U6374 ( .A(n6170), .ZN(n5205) );
  OAI21_X1 U6375 ( .B1(n6178), .B2(n6180), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5203) );
  OAI21_X1 U6376 ( .B1(n5205), .B2(n5204), .A(n5203), .ZN(n5208) );
  OAI22_X1 U6377 ( .A1(n6175), .A2(n5206), .B1(n6157), .B2(n6304), .ZN(n5207)
         );
  OR3_X1 U6378 ( .A1(n5209), .A2(n5208), .A3(n5207), .ZN(U2827) );
  INV_X1 U6379 ( .A(n5210), .ZN(n5212) );
  NAND2_X1 U6380 ( .A1(n5212), .A2(n5211), .ZN(n5213) );
  XNOR2_X1 U6381 ( .A(n5214), .B(n5213), .ZN(n6306) );
  AOI22_X1 U6382 ( .A1(n6300), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6334), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5215) );
  OAI21_X1 U6383 ( .B1(n5216), .B2(n6294), .A(n5215), .ZN(n5217) );
  AOI21_X1 U6384 ( .B1(n5218), .B2(n6287), .A(n5217), .ZN(n5219) );
  OAI21_X1 U6385 ( .B1(n6297), .B2(n6306), .A(n5219), .ZN(U2976) );
  XOR2_X1 U6386 ( .A(n5220), .B(n5191), .Z(n5288) );
  NOR2_X1 U6387 ( .A1(n6112), .A2(n5221), .ZN(n6107) );
  NAND2_X1 U6388 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6107), .ZN(n5382) );
  INV_X1 U6389 ( .A(n5382), .ZN(n5222) );
  AOI21_X1 U6390 ( .B1(n5222), .B2(n6137), .A(n6138), .ZN(n6106) );
  OAI22_X1 U6391 ( .A1(n6169), .A2(n3655), .B1(n5286), .B2(n6161), .ZN(n5228)
         );
  NAND2_X1 U6392 ( .A1(n5224), .A2(n5223), .ZN(n5225) );
  NAND2_X1 U6393 ( .A1(n5291), .A2(n5225), .ZN(n5279) );
  NOR2_X1 U6394 ( .A1(n5382), .A2(n6135), .ZN(n6095) );
  INV_X1 U6395 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6528) );
  AOI22_X1 U6396 ( .A1(PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n6178), .B1(n6095), 
        .B2(n6528), .ZN(n5226) );
  OAI211_X1 U6397 ( .C1(n6175), .C2(n5279), .A(n5226), .B(n6160), .ZN(n5227)
         );
  AOI211_X1 U6398 ( .C1(n6106), .C2(REIP_REG_12__SCAN_IN), .A(n5228), .B(n5227), .ZN(n5229) );
  OAI21_X1 U6399 ( .B1(n5233), .B2(n6151), .A(n5229), .ZN(U2815) );
  INV_X1 U6400 ( .A(n5279), .ZN(n5230) );
  AOI22_X1 U6401 ( .A1(n5230), .A2(n6191), .B1(EBX_REG_12__SCAN_IN), .B2(n5559), .ZN(n5231) );
  OAI21_X1 U6402 ( .B1(n5233), .B2(n5610), .A(n5231), .ZN(U2847) );
  AOI22_X1 U6403 ( .A1(n5375), .A2(DATAI_12_), .B1(n6205), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n5232) );
  OAI21_X1 U6404 ( .B1(n5233), .B2(n5626), .A(n5232), .ZN(U2879) );
  OAI22_X1 U6405 ( .A1(n5235), .A2(n6115), .B1(n6161), .B2(n5234), .ZN(n5236)
         );
  AOI21_X1 U6406 ( .B1(n6170), .B2(n4490), .A(n5236), .ZN(n5237) );
  OAI21_X1 U6407 ( .B1(n6175), .B2(n5238), .A(n5237), .ZN(n5242) );
  OAI21_X1 U6408 ( .B1(n5384), .B2(n6184), .A(n5547), .ZN(n6173) );
  AOI21_X1 U6409 ( .B1(n5240), .B2(n5239), .A(n6173), .ZN(n5241) );
  AOI211_X1 U6410 ( .C1(EBX_REG_3__SCAN_IN), .C2(n6172), .A(n5242), .B(n5241), 
        .ZN(n5243) );
  OAI21_X1 U6411 ( .B1(n6157), .B2(n5244), .A(n5243), .ZN(U2824) );
  AOI22_X1 U6412 ( .A1(n6180), .A2(n4445), .B1(REIP_REG_1__SCAN_IN), .B2(n5384), .ZN(n5245) );
  OAI21_X1 U6413 ( .B1(n4445), .B2(n6115), .A(n5245), .ZN(n5248) );
  NOR2_X1 U6414 ( .A1(n6157), .A2(n5246), .ZN(n5247) );
  AOI211_X1 U6415 ( .C1(n6170), .C2(n5249), .A(n5248), .B(n5247), .ZN(n5253)
         );
  INV_X1 U6416 ( .A(n6185), .ZN(n6164) );
  AOI22_X1 U6417 ( .A1(n6164), .A2(n5251), .B1(n6158), .B2(n5250), .ZN(n5252)
         );
  OAI211_X1 U6418 ( .C1(n5254), .C2(n6169), .A(n5253), .B(n5252), .ZN(U2826)
         );
  NAND2_X1 U6419 ( .A1(n5256), .A2(n5255), .ZN(n5258) );
  XOR2_X1 U6420 ( .A(n5258), .B(n5257), .Z(n6268) );
  OAI21_X1 U6421 ( .B1(n5985), .B2(n5260), .A(n5259), .ZN(n6006) );
  AOI22_X1 U6422 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6006), .B1(n6002), .B2(n5261), .ZN(n5264) );
  INV_X1 U6423 ( .A(n5262), .ZN(n6104) );
  AOI22_X1 U6424 ( .A1(n6333), .A2(n6104), .B1(n6334), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n5263) );
  OAI211_X1 U6425 ( .C1(n6268), .C2(n6307), .A(n5264), .B(n5263), .ZN(U3007)
         );
  OR2_X1 U6426 ( .A1(n5265), .A2(n5266), .ZN(n5313) );
  NAND2_X1 U6427 ( .A1(n5265), .A2(n5266), .ZN(n5267) );
  AOI22_X1 U6428 ( .A1(n5375), .A2(DATAI_13_), .B1(n6205), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5268) );
  OAI21_X1 U6429 ( .B1(n5294), .B2(n5626), .A(n5268), .ZN(U2878) );
  INV_X1 U6430 ( .A(n5269), .ZN(n5270) );
  NOR2_X1 U6431 ( .A1(n5271), .A2(n5270), .ZN(n5272) );
  XNOR2_X1 U6432 ( .A(n3013), .B(n5272), .ZN(n5290) );
  NOR3_X1 U6433 ( .A1(n5276), .A2(n5275), .A3(n5274), .ZN(n5277) );
  INV_X1 U6434 ( .A(n6006), .ZN(n5984) );
  OAI21_X1 U6435 ( .B1(n6009), .B2(n5277), .A(n5984), .ZN(n5282) );
  AOI21_X1 U6436 ( .B1(n6002), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5278) );
  INV_X1 U6437 ( .A(n5278), .ZN(n5281) );
  NAND2_X1 U6438 ( .A1(n6334), .A2(REIP_REG_12__SCAN_IN), .ZN(n5285) );
  OAI21_X1 U6439 ( .B1(n6309), .B2(n5279), .A(n5285), .ZN(n5280) );
  AOI21_X1 U6440 ( .B1(n5282), .B2(n5281), .A(n5280), .ZN(n5283) );
  OAI21_X1 U6441 ( .B1(n5290), .B2(n6307), .A(n5283), .ZN(U3006) );
  NAND2_X1 U6442 ( .A1(n6300), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5284)
         );
  OAI211_X1 U6443 ( .C1(n6294), .C2(n5286), .A(n5285), .B(n5284), .ZN(n5287)
         );
  AOI21_X1 U6444 ( .B1(n5288), .B2(n6287), .A(n5287), .ZN(n5289) );
  OAI21_X1 U6445 ( .B1(n5290), .B2(n6297), .A(n5289), .ZN(U2974) );
  INV_X1 U6446 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5293) );
  OAI21_X1 U6447 ( .B1(n3062), .B2(n3061), .A(n5320), .ZN(n6098) );
  OAI222_X1 U6448 ( .A1(n5294), .A2(n5610), .B1(n5293), .B2(n6195), .C1(n5608), 
        .C2(n6098), .ZN(U2846) );
  AND2_X1 U6449 ( .A1(n5307), .A2(n5304), .ZN(n5296) );
  NOR2_X1 U6450 ( .A1(n5297), .A2(n5296), .ZN(n5306) );
  NAND2_X1 U6451 ( .A1(n5306), .A2(n5298), .ZN(n5299) );
  NAND2_X1 U6452 ( .A1(n5602), .A2(n5299), .ZN(n6067) );
  AND2_X1 U6453 ( .A1(n5310), .A2(n5300), .ZN(n5301) );
  NOR2_X1 U6454 ( .A1(n5607), .A2(n5301), .ZN(n6068) );
  AOI22_X1 U6455 ( .A1(n6068), .A2(n6191), .B1(EBX_REG_17__SCAN_IN), .B2(n5559), .ZN(n5302) );
  OAI21_X1 U6456 ( .B1(n6067), .B2(n5610), .A(n5302), .ZN(U2842) );
  NOR2_X1 U6457 ( .A1(n5265), .A2(n5303), .ZN(n5305) );
  OR2_X1 U6458 ( .A1(n5305), .A2(n5304), .ZN(n5372) );
  OAI21_X1 U6459 ( .B1(n5372), .B2(n5307), .A(n5306), .ZN(n5741) );
  NAND2_X1 U6460 ( .A1(n5379), .A2(n5308), .ZN(n5309) );
  NAND2_X1 U6461 ( .A1(n5310), .A2(n5309), .ZN(n6082) );
  OAI222_X1 U6462 ( .A1(n5741), .A2(n5610), .B1(n5311), .B2(n6195), .C1(n5608), 
        .C2(n6082), .ZN(U2843) );
  NAND2_X1 U6463 ( .A1(n5313), .A2(n5312), .ZN(n5318) );
  OR2_X1 U6464 ( .A1(n5265), .A2(n5314), .ZN(n5316) );
  AND2_X1 U6465 ( .A1(n5316), .A2(n5315), .ZN(n5373) );
  OAI21_X1 U6466 ( .B1(n5318), .B2(n5317), .A(n5373), .ZN(n6088) );
  AOI22_X1 U6467 ( .A1(n5375), .A2(DATAI_14_), .B1(n6205), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5319) );
  OAI21_X1 U6468 ( .B1(n6088), .B2(n5626), .A(n5319), .ZN(U2877) );
  AOI21_X1 U6469 ( .B1(n5321), .B2(n5320), .A(n5378), .ZN(n5322) );
  INV_X1 U6470 ( .A(n5322), .ZN(n6084) );
  OAI222_X1 U6471 ( .A1(n6088), .A2(n5610), .B1(n5323), .B2(n6195), .C1(n5608), 
        .C2(n6084), .ZN(U2845) );
  INV_X1 U6472 ( .A(n6444), .ZN(n5324) );
  OAI21_X1 U6473 ( .B1(n5368), .B2(n5324), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n5325) );
  NOR2_X1 U6474 ( .A1(n5326), .A2(n6357), .ZN(n5327) );
  NOR2_X1 U6475 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5328), .ZN(n5365)
         );
  INV_X1 U6476 ( .A(n5329), .ZN(n5331) );
  INV_X1 U6477 ( .A(n5365), .ZN(n5330) );
  AOI22_X1 U6478 ( .A1(n5332), .A2(n5331), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5330), .ZN(n5333) );
  AOI22_X1 U6479 ( .A1(n6423), .A2(n5365), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5364), .ZN(n5336) );
  OAI21_X1 U6480 ( .B1(n6365), .B2(n6444), .A(n5336), .ZN(n5337) );
  AOI21_X1 U6481 ( .B1(n5368), .B2(n6362), .A(n5337), .ZN(n5338) );
  OAI21_X1 U6482 ( .B1(n5371), .B2(n5339), .A(n5338), .ZN(U3101) );
  AOI22_X1 U6483 ( .A1(n6401), .A2(n5365), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5364), .ZN(n5340) );
  OAI21_X1 U6484 ( .B1(n6375), .B2(n6444), .A(n5340), .ZN(n5341) );
  AOI21_X1 U6485 ( .B1(n5368), .B2(n6372), .A(n5341), .ZN(n5342) );
  OAI21_X1 U6486 ( .B1(n5371), .B2(n5343), .A(n5342), .ZN(U3103) );
  AOI22_X1 U6487 ( .A1(n6409), .A2(n5365), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5364), .ZN(n5344) );
  OAI21_X1 U6488 ( .B1(n6389), .B2(n6444), .A(n5344), .ZN(n5345) );
  AOI21_X1 U6489 ( .B1(n5368), .B2(n6386), .A(n5345), .ZN(n5346) );
  OAI21_X1 U6490 ( .B1(n5371), .B2(n5347), .A(n5346), .ZN(U3106) );
  AOI22_X1 U6491 ( .A1(n6377), .A2(n5365), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5364), .ZN(n5348) );
  OAI21_X1 U6492 ( .B1(n6381), .B2(n6444), .A(n5348), .ZN(n5349) );
  AOI21_X1 U6493 ( .B1(n5368), .B2(n6378), .A(n5349), .ZN(n5350) );
  OAI21_X1 U6494 ( .B1(n5371), .B2(n5351), .A(n5350), .ZN(U3104) );
  AOI22_X1 U6495 ( .A1(n6436), .A2(n5365), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5364), .ZN(n5352) );
  OAI21_X1 U6496 ( .B1(n6397), .B2(n6444), .A(n5352), .ZN(n5353) );
  AOI21_X1 U6497 ( .B1(n5368), .B2(n6393), .A(n5353), .ZN(n5354) );
  OAI21_X1 U6498 ( .B1(n5371), .B2(n5355), .A(n5354), .ZN(U3107) );
  AOI22_X1 U6499 ( .A1(n6367), .A2(n5365), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5364), .ZN(n5356) );
  OAI21_X1 U6500 ( .B1(n6371), .B2(n6444), .A(n5356), .ZN(n5357) );
  AOI21_X1 U6501 ( .B1(n5368), .B2(n6368), .A(n5357), .ZN(n5358) );
  OAI21_X1 U6502 ( .B1(n5371), .B2(n5359), .A(n5358), .ZN(U3102) );
  AOI22_X1 U6503 ( .A1(n6429), .A2(n5365), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5364), .ZN(n5360) );
  OAI21_X1 U6504 ( .B1(n6385), .B2(n6444), .A(n5360), .ZN(n5361) );
  AOI21_X1 U6505 ( .B1(n5368), .B2(n6382), .A(n5361), .ZN(n5362) );
  OAI21_X1 U6506 ( .B1(n5371), .B2(n5363), .A(n5362), .ZN(U3105) );
  AOI22_X1 U6507 ( .A1(n6417), .A2(n5365), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5364), .ZN(n5366) );
  OAI21_X1 U6508 ( .B1(n6361), .B2(n6444), .A(n5366), .ZN(n5367) );
  AOI21_X1 U6509 ( .B1(n6358), .B2(n5368), .A(n5367), .ZN(n5369) );
  OAI21_X1 U6510 ( .B1(n5371), .B2(n5370), .A(n5369), .ZN(U3100) );
  AOI21_X1 U6511 ( .B1(n5374), .B2(n5373), .A(n5372), .ZN(n5750) );
  INV_X1 U6512 ( .A(n5750), .ZN(n5391) );
  AOI22_X1 U6513 ( .A1(n5375), .A2(DATAI_15_), .B1(n6205), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5376) );
  OAI21_X1 U6514 ( .B1(n5391), .B2(n5626), .A(n5376), .ZN(U2876) );
  OR2_X1 U6515 ( .A1(n5378), .A2(n5377), .ZN(n5380) );
  AND2_X1 U6516 ( .A1(n5380), .A2(n5379), .ZN(n5996) );
  AOI22_X1 U6517 ( .A1(n5996), .A2(n6191), .B1(EBX_REG_15__SCAN_IN), .B2(n5559), .ZN(n5381) );
  OAI21_X1 U6518 ( .B1(n5391), .B2(n5610), .A(n5381), .ZN(U2844) );
  INV_X1 U6519 ( .A(n5748), .ZN(n5389) );
  NAND2_X1 U6520 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n6094) );
  NOR3_X1 U6521 ( .A1(n5383), .A2(n5382), .A3(n6094), .ZN(n6086) );
  NAND2_X1 U6522 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6086), .ZN(n5385) );
  NOR2_X1 U6523 ( .A1(n5384), .A2(n5385), .ZN(n6074) );
  NOR2_X1 U6524 ( .A1(n6138), .A2(n6074), .ZN(n6083) );
  AOI22_X1 U6525 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6172), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6083), .ZN(n5387) );
  AOI22_X1 U6526 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n6178), .B1(n6158), 
        .B2(n5996), .ZN(n5386) );
  INV_X1 U6527 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6532) );
  NAND2_X1 U6528 ( .A1(n5457), .A2(n6532), .ZN(n6073) );
  NAND4_X1 U6529 ( .A1(n5387), .A2(n5386), .A3(n6160), .A4(n6073), .ZN(n5388)
         );
  AOI21_X1 U6530 ( .B1(n6180), .B2(n5389), .A(n5388), .ZN(n5390) );
  OAI21_X1 U6531 ( .B1(n5391), .B2(n6151), .A(n5390), .ZN(U2812) );
  NAND2_X1 U6532 ( .A1(n5392), .A2(n5393), .ZN(n5395) );
  XNOR2_X1 U6533 ( .A(n5727), .B(n6003), .ZN(n5394) );
  XNOR2_X1 U6534 ( .A(n5395), .B(n5394), .ZN(n6011) );
  INV_X1 U6535 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5396) );
  OAI22_X1 U6536 ( .A1(n6282), .A2(n6757), .B1(n6308), .B2(n5396), .ZN(n5397)
         );
  AOI21_X1 U6537 ( .B1(n6276), .B2(n6089), .A(n5397), .ZN(n5399) );
  OR2_X1 U6538 ( .A1(n6088), .A2(n6303), .ZN(n5398) );
  OAI211_X1 U6539 ( .C1(n6011), .C2(n6297), .A(n5399), .B(n5398), .ZN(U2972)
         );
  AOI21_X1 U6540 ( .B1(n5400), .B2(n5404), .A(n5409), .ZN(n5411) );
  INV_X1 U6541 ( .A(n5401), .ZN(n5403) );
  NOR2_X1 U6542 ( .A1(n5403), .A2(n5402), .ZN(n5406) );
  NOR3_X1 U6543 ( .A1(n5404), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5865), 
        .ZN(n5405) );
  AOI211_X1 U6544 ( .C1(n5408), .C2(n5407), .A(n5406), .B(n5405), .ZN(n5410)
         );
  OAI22_X1 U6545 ( .A1(n5411), .A2(n3107), .B1(n5410), .B2(n5409), .ZN(U3459)
         );
  XOR2_X1 U6546 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5414), .Z(n5435) );
  AOI211_X1 U6547 ( .C1(n5495), .C2(n5416), .A(n5417), .B(n5415), .ZN(n5421)
         );
  INV_X1 U6548 ( .A(n5495), .ZN(n5453) );
  INV_X1 U6549 ( .A(n5417), .ZN(n5419) );
  AOI211_X1 U6550 ( .C1(n5541), .C2(n5453), .A(n5419), .B(n5418), .ZN(n5420)
         );
  NOR2_X1 U6551 ( .A1(n5421), .A2(n5420), .ZN(n5556) );
  NOR3_X1 U6552 ( .A1(n5755), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5423), 
        .ZN(n5426) );
  NAND2_X1 U6553 ( .A1(n5791), .A2(n5985), .ZN(n5422) );
  OAI211_X1 U6554 ( .C1(n5752), .C2(n5423), .A(INSTADDRPOINTER_REG_30__SCAN_IN), .B(n5422), .ZN(n5424) );
  NAND2_X1 U6555 ( .A1(n6334), .A2(REIP_REG_30__SCAN_IN), .ZN(n5430) );
  NAND2_X1 U6556 ( .A1(n5424), .A2(n5430), .ZN(n5425) );
  AOI211_X1 U6557 ( .C1(n5556), .C2(n6333), .A(n5426), .B(n5425), .ZN(n5427)
         );
  OAI21_X1 U6558 ( .B1(n5435), .B2(n6307), .A(n5427), .ZN(U2988) );
  NAND2_X1 U6559 ( .A1(n6276), .A2(n5474), .ZN(n5431) );
  OAI211_X1 U6560 ( .C1(n5432), .C2(n6282), .A(n5431), .B(n5430), .ZN(n5433)
         );
  AOI21_X1 U6561 ( .B1(n5472), .B2(n6287), .A(n5433), .ZN(n5434) );
  OAI21_X1 U6562 ( .B1(n5435), .B2(n6297), .A(n5434), .ZN(U2956) );
  OAI21_X1 U6563 ( .B1(n6282), .B2(n5437), .A(n5436), .ZN(n5441) );
  INV_X1 U6564 ( .A(n5443), .ZN(n5480) );
  AOI22_X1 U6565 ( .A1(n6202), .A2(DATAI_29_), .B1(n6205), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5448) );
  AND2_X1 U6566 ( .A1(n3222), .A2(n5445), .ZN(n5446) );
  NAND2_X1 U6567 ( .A1(n6206), .A2(DATAI_13_), .ZN(n5447) );
  OAI211_X1 U6568 ( .C1(n5443), .C2(n5626), .A(n5448), .B(n5447), .ZN(U2862)
         );
  INV_X1 U6569 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5456) );
  INV_X1 U6570 ( .A(n5449), .ZN(n5455) );
  AOI21_X1 U6571 ( .B1(n5451), .B2(n5596), .A(n5450), .ZN(n5452) );
  NAND2_X1 U6572 ( .A1(n5453), .A2(n5452), .ZN(n5454) );
  NAND2_X1 U6573 ( .A1(n5455), .A2(n5454), .ZN(n5481) );
  OAI222_X1 U6574 ( .A1(n5610), .A2(n5443), .B1(n5456), .B2(n6195), .C1(n5481), 
        .C2(n5608), .ZN(U2830) );
  INV_X1 U6575 ( .A(n5615), .ZN(n5471) );
  INV_X1 U6576 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6535) );
  INV_X1 U6577 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6578 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5457), .ZN(n6078) );
  NOR2_X1 U6579 ( .A1(n5458), .A2(n6078), .ZN(n6062) );
  NAND2_X1 U6580 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6062), .ZN(n6058) );
  NAND3_X1 U6581 ( .A1(n5960), .A2(REIP_REG_20__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .ZN(n5959) );
  NAND2_X1 U6582 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5946) );
  NOR2_X1 U6583 ( .A1(n5959), .A2(n5946), .ZN(n5932) );
  NAND2_X1 U6584 ( .A1(n5932), .A2(REIP_REG_23__SCAN_IN), .ZN(n5927) );
  NAND3_X1 U6585 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .A3(
        REIP_REG_26__SCAN_IN), .ZN(n5460) );
  NOR2_X1 U6586 ( .A1(n5927), .A2(n5460), .ZN(n5509) );
  AND2_X1 U6587 ( .A1(REIP_REG_27__SCAN_IN), .A2(REIP_REG_28__SCAN_IN), .ZN(
        n5462) );
  NAND2_X1 U6588 ( .A1(n5509), .A2(n5462), .ZN(n5490) );
  INV_X1 U6589 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6557) );
  INV_X1 U6590 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6554) );
  NOR4_X1 U6591 ( .A1(n5490), .A2(REIP_REG_31__SCAN_IN), .A3(n6557), .A4(n6554), .ZN(n5469) );
  NAND2_X1 U6592 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n5459) );
  NAND4_X1 U6593 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .A4(n6074), .ZN(n5546) );
  NOR3_X1 U6594 ( .A1(n6535), .A2(n5459), .A3(n5546), .ZN(n5938) );
  NAND4_X1 U6595 ( .A1(n5938), .A2(REIP_REG_23__SCAN_IN), .A3(
        REIP_REG_22__SCAN_IN), .A4(REIP_REG_21__SCAN_IN), .ZN(n5534) );
  OR2_X1 U6596 ( .A1(n5534), .A2(n5460), .ZN(n5461) );
  NAND2_X1 U6597 ( .A1(n5461), .A2(n5547), .ZN(n5520) );
  OR2_X1 U6598 ( .A1(n6185), .A2(n5462), .ZN(n5463) );
  OAI21_X1 U6599 ( .B1(REIP_REG_29__SCAN_IN), .B2(n6185), .A(n5500), .ZN(n5473) );
  AOI21_X1 U6600 ( .B1(n6164), .B2(n6557), .A(n5473), .ZN(n5467) );
  INV_X1 U6601 ( .A(REIP_REG_31__SCAN_IN), .ZN(n5466) );
  AOI22_X1 U6602 ( .A1(n5464), .A2(EBX_REG_31__SCAN_IN), .B1(n6178), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5465) );
  OAI21_X1 U6603 ( .B1(n5467), .B2(n5466), .A(n5465), .ZN(n5468) );
  OAI21_X1 U6604 ( .B1(n5471), .B2(n6151), .A(n5470), .ZN(U2796) );
  NOR3_X1 U6605 ( .A1(n5490), .A2(REIP_REG_30__SCAN_IN), .A3(n6554), .ZN(n5478) );
  INV_X1 U6606 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5558) );
  NAND2_X1 U6607 ( .A1(n5473), .A2(REIP_REG_30__SCAN_IN), .ZN(n5476) );
  AOI22_X1 U6608 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n6178), .B1(n6180), 
        .B2(n5474), .ZN(n5475) );
  OAI211_X1 U6609 ( .C1(n6169), .C2(n5558), .A(n5476), .B(n5475), .ZN(n5477)
         );
  AOI211_X1 U6610 ( .C1(n5556), .C2(n6158), .A(n5478), .B(n5477), .ZN(n5479)
         );
  NAND2_X1 U6611 ( .A1(n5480), .A2(n6143), .ZN(n5489) );
  INV_X1 U6612 ( .A(n5481), .ZN(n5757) );
  INV_X1 U6613 ( .A(n5482), .ZN(n5483) );
  OAI22_X1 U6614 ( .A1(n5484), .A2(n6115), .B1(n6161), .B2(n5483), .ZN(n5485)
         );
  AOI21_X1 U6615 ( .B1(n6172), .B2(EBX_REG_29__SCAN_IN), .A(n5485), .ZN(n5486)
         );
  OAI21_X1 U6616 ( .B1(n5500), .B2(n6554), .A(n5486), .ZN(n5487) );
  AOI21_X1 U6617 ( .B1(n5757), .B2(n6158), .A(n5487), .ZN(n5488) );
  OAI211_X1 U6618 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5490), .A(n5489), .B(n5488), .ZN(U2798) );
  AOI21_X1 U6619 ( .B1(n5491), .B2(n5438), .A(n4282), .ZN(n5658) );
  INV_X1 U6620 ( .A(n5658), .ZN(n5623) );
  INV_X1 U6621 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6550) );
  NOR2_X1 U6622 ( .A1(n6550), .A2(REIP_REG_28__SCAN_IN), .ZN(n5502) );
  INV_X1 U6623 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6552) );
  AND2_X1 U6624 ( .A1(n5493), .A2(n5492), .ZN(n5494) );
  NOR2_X1 U6625 ( .A1(n5495), .A2(n5494), .ZN(n5769) );
  NAND2_X1 U6626 ( .A1(n5769), .A2(n6158), .ZN(n5499) );
  OAI22_X1 U6627 ( .A1(n5496), .A2(n6115), .B1(n6161), .B2(n5656), .ZN(n5497)
         );
  AOI21_X1 U6628 ( .B1(n6172), .B2(EBX_REG_28__SCAN_IN), .A(n5497), .ZN(n5498)
         );
  OAI211_X1 U6629 ( .C1(n5500), .C2(n6552), .A(n5499), .B(n5498), .ZN(n5501)
         );
  AOI21_X1 U6630 ( .B1(n5509), .B2(n5502), .A(n5501), .ZN(n5503) );
  OAI21_X1 U6631 ( .B1(n5623), .B2(n6151), .A(n5503), .ZN(U2799) );
  NOR2_X1 U6632 ( .A1(n5520), .A2(n6550), .ZN(n5508) );
  AOI22_X1 U6633 ( .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n6178), .B1(n6180), 
        .B2(n5504), .ZN(n5506) );
  NAND2_X1 U6634 ( .A1(n6172), .A2(EBX_REG_27__SCAN_IN), .ZN(n5505) );
  OAI211_X1 U6635 ( .C1(n5561), .C2(n6175), .A(n5506), .B(n5505), .ZN(n5507)
         );
  AOI211_X1 U6636 ( .C1(n5509), .C2(n6550), .A(n5508), .B(n5507), .ZN(n5510)
         );
  OAI21_X1 U6637 ( .B1(n5627), .B2(n6151), .A(n5510), .ZN(U2800) );
  AOI21_X1 U6638 ( .B1(n5512), .B2(n5526), .A(n5511), .ZN(n5668) );
  INV_X1 U6639 ( .A(n5668), .ZN(n5630) );
  OAI22_X1 U6640 ( .A1(n5513), .A2(n6115), .B1(n6161), .B2(n5666), .ZN(n5518)
         );
  NAND2_X1 U6641 ( .A1(n5531), .A2(n5514), .ZN(n5515) );
  NAND2_X1 U6642 ( .A1(n5516), .A2(n5515), .ZN(n5772) );
  NOR2_X1 U6643 ( .A1(n5772), .A2(n6175), .ZN(n5517) );
  AOI211_X1 U6644 ( .C1(EBX_REG_26__SCAN_IN), .C2(n6172), .A(n5518), .B(n5517), 
        .ZN(n5524) );
  INV_X1 U6645 ( .A(REIP_REG_25__SCAN_IN), .ZN(n5519) );
  NOR3_X1 U6646 ( .A1(n5927), .A2(n6599), .A3(n5519), .ZN(n5522) );
  INV_X1 U6647 ( .A(n5520), .ZN(n5521) );
  OAI21_X1 U6648 ( .B1(n5522), .B2(REIP_REG_26__SCAN_IN), .A(n5521), .ZN(n5523) );
  OAI211_X1 U6649 ( .C1(n5630), .C2(n6151), .A(n5524), .B(n5523), .ZN(U2801)
         );
  OAI21_X1 U6650 ( .B1(n5525), .B2(n5527), .A(n5526), .ZN(n5678) );
  INV_X1 U6651 ( .A(n5678), .ZN(n5539) );
  XNOR2_X1 U6652 ( .A(REIP_REG_24__SCAN_IN), .B(REIP_REG_25__SCAN_IN), .ZN(
        n5528) );
  NOR2_X1 U6653 ( .A1(n5927), .A2(n5528), .ZN(n5538) );
  OR2_X1 U6654 ( .A1(n5569), .A2(n5529), .ZN(n5530) );
  NAND2_X1 U6655 ( .A1(n5531), .A2(n5530), .ZN(n5783) );
  INV_X1 U6656 ( .A(n5672), .ZN(n5532) );
  OAI22_X1 U6657 ( .A1(n5670), .A2(n6115), .B1(n6161), .B2(n5532), .ZN(n5533)
         );
  AOI21_X1 U6658 ( .B1(n6172), .B2(EBX_REG_25__SCAN_IN), .A(n5533), .ZN(n5536)
         );
  AND2_X1 U6659 ( .A1(n5534), .A2(n5547), .ZN(n5933) );
  NAND2_X1 U6660 ( .A1(n5933), .A2(REIP_REG_25__SCAN_IN), .ZN(n5535) );
  OAI211_X1 U6661 ( .C1(n5783), .C2(n6175), .A(n5536), .B(n5535), .ZN(n5537)
         );
  AOI211_X1 U6662 ( .C1(n5539), .C2(n6143), .A(n5538), .B(n5537), .ZN(n5540)
         );
  INV_X1 U6663 ( .A(n5540), .ZN(U2802) );
  MUX2_X1 U6664 ( .A(n5595), .B(n5542), .S(n5541), .Z(n5543) );
  INV_X1 U6665 ( .A(n5543), .ZN(n5606) );
  NAND2_X1 U6666 ( .A1(n5607), .A2(n5606), .ZN(n5605) );
  XNOR2_X1 U6667 ( .A(n5605), .B(n3058), .ZN(n5839) );
  AOI21_X1 U6668 ( .B1(n5545), .B2(n5604), .A(n5591), .ZN(n5724) );
  NAND2_X1 U6669 ( .A1(n5724), .A2(n6143), .ZN(n5552) );
  INV_X1 U6670 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6538) );
  NAND2_X1 U6671 ( .A1(n5547), .A2(n5546), .ZN(n6071) );
  OAI21_X1 U6672 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6058), .A(n6071), .ZN(n5550) );
  AOI22_X1 U6673 ( .A1(EBX_REG_19__SCAN_IN), .A2(n6172), .B1(n5720), .B2(n6180), .ZN(n5548) );
  OAI211_X1 U6674 ( .C1(n6115), .C2(n5722), .A(n5548), .B(n6160), .ZN(n5549)
         );
  AOI221_X1 U6675 ( .B1(n5960), .B2(n6538), .C1(n5550), .C2(
        REIP_REG_19__SCAN_IN), .A(n5549), .ZN(n5551) );
  OAI211_X1 U6676 ( .C1(n5839), .C2(n6175), .A(n5552), .B(n5551), .ZN(U2808)
         );
  INV_X1 U6677 ( .A(n5553), .ZN(n5555) );
  OAI22_X1 U6678 ( .A1(n5555), .A2(n5608), .B1(n6195), .B2(n5554), .ZN(U2828)
         );
  INV_X1 U6679 ( .A(n5556), .ZN(n5557) );
  OAI222_X1 U6680 ( .A1(n5610), .A2(n5620), .B1(n5558), .B2(n6195), .C1(n5557), 
        .C2(n5608), .ZN(U2829) );
  AOI22_X1 U6681 ( .A1(n5769), .A2(n6191), .B1(EBX_REG_28__SCAN_IN), .B2(n5559), .ZN(n5560) );
  OAI21_X1 U6682 ( .B1(n5623), .B2(n5610), .A(n5560), .ZN(U2831) );
  INV_X1 U6683 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5562) );
  OAI222_X1 U6684 ( .A1(n5610), .A2(n5627), .B1(n5562), .B2(n6195), .C1(n5561), 
        .C2(n5608), .ZN(U2832) );
  OAI222_X1 U6685 ( .A1(n5610), .A2(n5630), .B1(n5563), .B2(n6195), .C1(n5772), 
        .C2(n5608), .ZN(U2833) );
  OAI222_X1 U6686 ( .A1(n5678), .A2(n5610), .B1(n6195), .B2(n3695), .C1(n5783), 
        .C2(n5608), .ZN(U2834) );
  AOI21_X1 U6687 ( .B1(n5565), .B2(n5564), .A(n5525), .ZN(n5566) );
  INV_X1 U6688 ( .A(n5566), .ZN(n5923) );
  NOR2_X1 U6689 ( .A1(n5576), .A2(n5567), .ZN(n5568) );
  OR2_X1 U6690 ( .A1(n5569), .A2(n5568), .ZN(n5922) );
  OAI22_X1 U6691 ( .A1(n5922), .A2(n5608), .B1(n5570), .B2(n6195), .ZN(n5571)
         );
  INV_X1 U6692 ( .A(n5571), .ZN(n5572) );
  OAI21_X1 U6693 ( .B1(n5923), .B2(n5610), .A(n5572), .ZN(U2835) );
  AOI21_X1 U6694 ( .B1(n3057), .B2(n5580), .A(n5575), .ZN(n5577) );
  OR2_X1 U6695 ( .A1(n5577), .A2(n5576), .ZN(n5929) );
  OAI222_X1 U6696 ( .A1(n5610), .A2(n5930), .B1(n6195), .B2(n3684), .C1(n5929), 
        .C2(n5608), .ZN(U2836) );
  AOI21_X1 U6697 ( .B1(n5579), .B2(n5578), .A(n5573), .ZN(n5945) );
  INV_X1 U6698 ( .A(n5945), .ZN(n5639) );
  INV_X1 U6699 ( .A(n5580), .ZN(n5581) );
  XNOR2_X1 U6700 ( .A(n5588), .B(n5581), .ZN(n5950) );
  OAI22_X1 U6701 ( .A1(n5950), .A2(n5608), .B1(n5943), .B2(n6195), .ZN(n5582)
         );
  INV_X1 U6702 ( .A(n5582), .ZN(n5583) );
  OAI21_X1 U6703 ( .B1(n5639), .B2(n5610), .A(n5583), .ZN(U2837) );
  NAND2_X1 U6704 ( .A1(n5593), .A2(n5584), .ZN(n5585) );
  NAND2_X1 U6705 ( .A1(n5578), .A2(n5585), .ZN(n5955) );
  INV_X1 U6706 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U6707 ( .A1(n3050), .A2(n5586), .ZN(n5587) );
  NAND2_X1 U6708 ( .A1(n5588), .A2(n5587), .ZN(n5954) );
  OAI222_X1 U6709 ( .A1(n5955), .A2(n5610), .B1(n5589), .B2(n6195), .C1(n5608), 
        .C2(n5954), .ZN(U2838) );
  OR2_X1 U6710 ( .A1(n5591), .A2(n5590), .ZN(n5592) );
  NAND2_X1 U6711 ( .A1(n5593), .A2(n5592), .ZN(n5965) );
  INV_X1 U6712 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5599) );
  MUX2_X1 U6713 ( .A(n5596), .B(n5595), .S(n5594), .Z(n5598) );
  XNOR2_X1 U6714 ( .A(n5598), .B(n5597), .ZN(n5830) );
  INV_X1 U6715 ( .A(n5830), .ZN(n5964) );
  OAI222_X1 U6716 ( .A1(n5965), .A2(n5610), .B1(n5599), .B2(n6195), .C1(n5608), 
        .C2(n5964), .ZN(U2839) );
  INV_X1 U6717 ( .A(n5724), .ZN(n5646) );
  OAI222_X1 U6718 ( .A1(n5646), .A2(n5610), .B1(n5600), .B2(n6195), .C1(n5608), 
        .C2(n5839), .ZN(U2840) );
  NAND2_X1 U6719 ( .A1(n5602), .A2(n5601), .ZN(n5603) );
  AND2_X1 U6720 ( .A1(n5604), .A2(n5603), .ZN(n6196) );
  INV_X1 U6721 ( .A(n6196), .ZN(n5611) );
  OAI21_X1 U6722 ( .B1(n5607), .B2(n5606), .A(n5605), .ZN(n6061) );
  OAI222_X1 U6723 ( .A1(n5611), .A2(n5610), .B1(n5609), .B2(n6195), .C1(n5608), 
        .C2(n6061), .ZN(U2841) );
  NAND2_X1 U6724 ( .A1(n5615), .A2(n5614), .ZN(n5617) );
  AOI22_X1 U6725 ( .A1(n6202), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6205), .ZN(n5616) );
  NAND2_X1 U6726 ( .A1(n5617), .A2(n5616), .ZN(U2860) );
  AOI22_X1 U6727 ( .A1(n6202), .A2(DATAI_30_), .B1(n6205), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U6728 ( .A1(n6206), .A2(DATAI_14_), .ZN(n5618) );
  OAI211_X1 U6729 ( .C1(n5620), .C2(n5626), .A(n5619), .B(n5618), .ZN(U2861)
         );
  AOI22_X1 U6730 ( .A1(n6202), .A2(DATAI_28_), .B1(n6205), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U6731 ( .A1(n6206), .A2(DATAI_12_), .ZN(n5621) );
  OAI211_X1 U6732 ( .C1(n5623), .C2(n5626), .A(n5622), .B(n5621), .ZN(U2863)
         );
  AOI22_X1 U6733 ( .A1(n6202), .A2(DATAI_27_), .B1(n6205), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U6734 ( .A1(n6206), .A2(DATAI_11_), .ZN(n5624) );
  OAI211_X1 U6735 ( .C1(n5627), .C2(n5626), .A(n5625), .B(n5624), .ZN(U2864)
         );
  AOI22_X1 U6736 ( .A1(n6202), .A2(DATAI_26_), .B1(n6205), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U6737 ( .A1(n6206), .A2(DATAI_10_), .ZN(n5628) );
  OAI211_X1 U6738 ( .C1(n5630), .C2(n5626), .A(n5629), .B(n5628), .ZN(U2865)
         );
  AOI22_X1 U6739 ( .A1(n6202), .A2(DATAI_25_), .B1(n6205), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5632) );
  NAND2_X1 U6740 ( .A1(n6206), .A2(DATAI_9_), .ZN(n5631) );
  OAI211_X1 U6741 ( .C1(n5678), .C2(n5626), .A(n5632), .B(n5631), .ZN(U2866)
         );
  AOI22_X1 U6742 ( .A1(n6202), .A2(DATAI_24_), .B1(n6205), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5634) );
  NAND2_X1 U6743 ( .A1(n6206), .A2(DATAI_8_), .ZN(n5633) );
  OAI211_X1 U6744 ( .C1(n5923), .C2(n5626), .A(n5634), .B(n5633), .ZN(U2867)
         );
  AOI22_X1 U6745 ( .A1(n6202), .A2(DATAI_23_), .B1(n6205), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5636) );
  NAND2_X1 U6746 ( .A1(n6206), .A2(DATAI_7_), .ZN(n5635) );
  OAI211_X1 U6747 ( .C1(n5930), .C2(n5626), .A(n5636), .B(n5635), .ZN(U2868)
         );
  AOI22_X1 U6748 ( .A1(n6202), .A2(DATAI_22_), .B1(n6205), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5638) );
  NAND2_X1 U6749 ( .A1(n6206), .A2(DATAI_6_), .ZN(n5637) );
  OAI211_X1 U6750 ( .C1(n5639), .C2(n5626), .A(n5638), .B(n5637), .ZN(U2869)
         );
  AOI22_X1 U6751 ( .A1(n6202), .A2(DATAI_21_), .B1(n6205), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5641) );
  NAND2_X1 U6752 ( .A1(n6206), .A2(DATAI_5_), .ZN(n5640) );
  OAI211_X1 U6753 ( .C1(n5955), .C2(n5626), .A(n5641), .B(n5640), .ZN(U2870)
         );
  AOI22_X1 U6754 ( .A1(n6202), .A2(DATAI_20_), .B1(n6205), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5643) );
  NAND2_X1 U6755 ( .A1(n6206), .A2(DATAI_4_), .ZN(n5642) );
  OAI211_X1 U6756 ( .C1(n5965), .C2(n5626), .A(n5643), .B(n5642), .ZN(U2871)
         );
  AOI22_X1 U6757 ( .A1(n6202), .A2(DATAI_19_), .B1(n6205), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5645) );
  NAND2_X1 U6758 ( .A1(n6206), .A2(DATAI_3_), .ZN(n5644) );
  OAI211_X1 U6759 ( .C1(n5646), .C2(n5626), .A(n5645), .B(n5644), .ZN(U2872)
         );
  INV_X1 U6760 ( .A(n3747), .ZN(n5654) );
  NAND2_X1 U6761 ( .A1(n5647), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5651) );
  NAND3_X1 U6762 ( .A1(n3747), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5648), .ZN(n5650) );
  OAI211_X1 U6763 ( .C1(n5652), .C2(n5651), .A(n5650), .B(n5649), .ZN(n5653)
         );
  AOI21_X1 U6764 ( .B1(n3746), .B2(n5654), .A(n5653), .ZN(n5771) );
  NAND2_X1 U6765 ( .A1(n6334), .A2(REIP_REG_28__SCAN_IN), .ZN(n5766) );
  NAND2_X1 U6766 ( .A1(n6300), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5655)
         );
  OAI211_X1 U6767 ( .C1(n6294), .C2(n5656), .A(n5766), .B(n5655), .ZN(n5657)
         );
  AOI21_X1 U6768 ( .B1(n5658), .B2(n6287), .A(n5657), .ZN(n5659) );
  OAI21_X1 U6769 ( .B1(n5771), .B2(n6297), .A(n5659), .ZN(U2958) );
  NAND2_X1 U6770 ( .A1(n5662), .A2(n5661), .ZN(n5663) );
  XNOR2_X1 U6771 ( .A(n5664), .B(n5663), .ZN(n5780) );
  NAND2_X1 U6772 ( .A1(n6334), .A2(REIP_REG_26__SCAN_IN), .ZN(n5773) );
  NAND2_X1 U6773 ( .A1(n6300), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5665)
         );
  OAI211_X1 U6774 ( .C1(n6294), .C2(n5666), .A(n5773), .B(n5665), .ZN(n5667)
         );
  AOI21_X1 U6775 ( .B1(n5668), .B2(n6287), .A(n5667), .ZN(n5669) );
  OAI21_X1 U6776 ( .B1(n5780), .B2(n6297), .A(n5669), .ZN(U2960) );
  NAND2_X1 U6777 ( .A1(n6334), .A2(REIP_REG_25__SCAN_IN), .ZN(n5782) );
  OAI21_X1 U6778 ( .B1(n6282), .B2(n5670), .A(n5782), .ZN(n5671) );
  AOI21_X1 U6779 ( .B1(n6276), .B2(n5672), .A(n5671), .ZN(n5677) );
  OAI21_X1 U6780 ( .B1(n5675), .B2(n5674), .A(n5673), .ZN(n5781) );
  NAND2_X1 U6781 ( .A1(n5781), .A2(n6289), .ZN(n5676) );
  OAI211_X1 U6782 ( .C1(n5678), .C2(n6303), .A(n5677), .B(n5676), .ZN(U2961)
         );
  BUF_X1 U6783 ( .A(n5679), .Z(n5691) );
  OAI21_X1 U6784 ( .B1(n5691), .B2(n3516), .A(n5727), .ZN(n5680) );
  AND2_X2 U6785 ( .A1(n5717), .A2(n5680), .ZN(n5711) );
  XNOR2_X1 U6786 ( .A(n5727), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5712)
         );
  XNOR2_X1 U6787 ( .A(n5727), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5705)
         );
  INV_X1 U6788 ( .A(n5700), .ZN(n5682) );
  NAND3_X1 U6789 ( .A1(n5727), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U6790 ( .A1(n5682), .A2(n5681), .ZN(n5685) );
  NAND3_X1 U6791 ( .A1(n3506), .A2(n5803), .A3(n6709), .ZN(n5683) );
  NAND2_X1 U6792 ( .A1(n5685), .A2(n5684), .ZN(n5686) );
  NAND2_X1 U6793 ( .A1(n5797), .A2(n6289), .ZN(n5690) );
  NAND2_X1 U6794 ( .A1(n6334), .A2(REIP_REG_24__SCAN_IN), .ZN(n5794) );
  OAI21_X1 U6795 ( .B1(n6282), .B2(n5687), .A(n5794), .ZN(n5688) );
  AOI21_X1 U6796 ( .B1(n6276), .B2(n5919), .A(n5688), .ZN(n5689) );
  OAI211_X1 U6797 ( .C1(n6303), .C2(n5923), .A(n5690), .B(n5689), .ZN(U2962)
         );
  NOR3_X1 U6798 ( .A1(n5691), .A2(n5831), .A3(n5692), .ZN(n5694) );
  NOR2_X1 U6799 ( .A1(n5704), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5693)
         );
  MUX2_X1 U6800 ( .A(n5694), .B(n5693), .S(n3506), .Z(n5695) );
  XNOR2_X1 U6801 ( .A(n5695), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5806)
         );
  NAND2_X1 U6802 ( .A1(n6334), .A2(REIP_REG_23__SCAN_IN), .ZN(n5800) );
  OAI21_X1 U6803 ( .B1(n6282), .B2(n5936), .A(n5800), .ZN(n5697) );
  NOR2_X1 U6804 ( .A1(n5930), .A2(n6303), .ZN(n5696) );
  AOI211_X1 U6805 ( .C1(n5928), .C2(n6276), .A(n5697), .B(n5696), .ZN(n5698)
         );
  OAI21_X1 U6806 ( .B1(n5806), .B2(n6297), .A(n5698), .ZN(U2963) );
  XNOR2_X1 U6807 ( .A(n5727), .B(n6709), .ZN(n5699) );
  XNOR2_X1 U6808 ( .A(n5700), .B(n5699), .ZN(n5815) );
  NAND2_X1 U6809 ( .A1(n6334), .A2(REIP_REG_22__SCAN_IN), .ZN(n5807) );
  NAND2_X1 U6810 ( .A1(n6300), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5701)
         );
  OAI211_X1 U6811 ( .C1(n6294), .C2(n5937), .A(n5807), .B(n5701), .ZN(n5702)
         );
  AOI21_X1 U6812 ( .B1(n5945), .B2(n6287), .A(n5702), .ZN(n5703) );
  OAI21_X1 U6813 ( .B1(n5815), .B2(n6297), .A(n5703), .ZN(U2964) );
  OAI21_X1 U6814 ( .B1(n5706), .B2(n5705), .A(n5704), .ZN(n5816) );
  NAND2_X1 U6815 ( .A1(n5816), .A2(n6289), .ZN(n5710) );
  INV_X1 U6816 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U6817 ( .A1(n6334), .A2(REIP_REG_21__SCAN_IN), .ZN(n5818) );
  OAI21_X1 U6818 ( .B1(n6282), .B2(n5707), .A(n5818), .ZN(n5708) );
  AOI21_X1 U6819 ( .B1(n6276), .B2(n5951), .A(n5708), .ZN(n5709) );
  OAI211_X1 U6820 ( .C1(n6303), .C2(n5955), .A(n5710), .B(n5709), .ZN(U2965)
         );
  XOR2_X1 U6821 ( .A(n5712), .B(n5711), .Z(n5824) );
  AND2_X1 U6822 ( .A1(n6334), .A2(REIP_REG_20__SCAN_IN), .ZN(n5829) );
  AOI21_X1 U6823 ( .B1(n6300), .B2(PHYADDRPOINTER_REG_20__SCAN_IN), .A(n5829), 
        .ZN(n5714) );
  OR2_X1 U6824 ( .A1(n6294), .A2(n5961), .ZN(n5713) );
  OAI211_X1 U6825 ( .C1(n5965), .C2(n6303), .A(n5714), .B(n5713), .ZN(n5715)
         );
  AOI21_X1 U6826 ( .B1(n5824), .B2(n6289), .A(n5715), .ZN(n5716) );
  INV_X1 U6827 ( .A(n5716), .ZN(U2966) );
  OAI21_X1 U6828 ( .B1(n5718), .B2(n3516), .A(n3000), .ZN(n5719) );
  XNOR2_X1 U6829 ( .A(n5719), .B(n5727), .ZN(n5843) );
  NAND2_X1 U6830 ( .A1(n6276), .A2(n5720), .ZN(n5721) );
  NAND2_X1 U6831 ( .A1(n6334), .A2(REIP_REG_19__SCAN_IN), .ZN(n5837) );
  OAI211_X1 U6832 ( .C1(n6282), .C2(n5722), .A(n5721), .B(n5837), .ZN(n5723)
         );
  AOI21_X1 U6833 ( .B1(n5724), .B2(n6287), .A(n5723), .ZN(n5725) );
  OAI21_X1 U6834 ( .B1(n5843), .B2(n6297), .A(n5725), .ZN(U2967) );
  NAND2_X1 U6835 ( .A1(n5727), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5845) );
  INV_X1 U6836 ( .A(n5726), .ZN(n5846) );
  NAND2_X1 U6837 ( .A1(n5846), .A2(n5737), .ZN(n5728) );
  OAI211_X1 U6838 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5727), .A(n5728), .B(n5845), .ZN(n5731) );
  NOR4_X1 U6839 ( .A1(n5727), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A4(INSTADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n5730) );
  NAND2_X1 U6840 ( .A1(n5729), .A2(n5730), .ZN(n5844) );
  OAI211_X1 U6841 ( .C1(n5726), .C2(n5845), .A(n5731), .B(n5844), .ZN(n5980)
         );
  NAND2_X1 U6842 ( .A1(n5980), .A2(n6289), .ZN(n5735) );
  INV_X1 U6843 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5732) );
  OAI22_X1 U6844 ( .A1(n6282), .A2(n6063), .B1(n6308), .B2(n5732), .ZN(n5733)
         );
  AOI21_X1 U6845 ( .B1(n6276), .B2(n6066), .A(n5733), .ZN(n5734) );
  OAI211_X1 U6846 ( .C1(n6303), .C2(n6067), .A(n5735), .B(n5734), .ZN(U2969)
         );
  INV_X1 U6847 ( .A(n5737), .ZN(n5740) );
  AND2_X1 U6848 ( .A1(n5737), .A2(n5736), .ZN(n5738) );
  OAI22_X1 U6849 ( .A1(n5846), .A2(n5740), .B1(n5739), .B2(n5738), .ZN(n5988)
         );
  INV_X1 U6850 ( .A(n5741), .ZN(n6204) );
  INV_X1 U6851 ( .A(n6076), .ZN(n5743) );
  AOI22_X1 U6852 ( .A1(n6300), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6334), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5742) );
  OAI21_X1 U6853 ( .B1(n5743), .B2(n6294), .A(n5742), .ZN(n5744) );
  AOI21_X1 U6854 ( .B1(n6204), .B2(n6287), .A(n5744), .ZN(n5745) );
  OAI21_X1 U6855 ( .B1(n5988), .B2(n6297), .A(n5745), .ZN(U2970) );
  XNOR2_X1 U6856 ( .A(n5727), .B(n6000), .ZN(n5746) );
  XNOR2_X1 U6857 ( .A(n5729), .B(n5746), .ZN(n5995) );
  AOI22_X1 U6858 ( .A1(n6300), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n6334), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5747) );
  OAI21_X1 U6859 ( .B1(n5748), .B2(n6294), .A(n5747), .ZN(n5749) );
  AOI21_X1 U6860 ( .B1(n5750), .B2(n6287), .A(n5749), .ZN(n5751) );
  OAI21_X1 U6861 ( .B1(n6297), .B2(n5995), .A(n5751), .ZN(U2971) );
  NAND2_X1 U6862 ( .A1(n5752), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5754) );
  OAI211_X1 U6863 ( .C1(n5755), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5754), .B(n5753), .ZN(n5756) );
  AOI21_X1 U6864 ( .B1(n5757), .B2(n6333), .A(n5756), .ZN(n5758) );
  OAI21_X1 U6865 ( .B1(n5759), .B2(n6307), .A(n5758), .ZN(U2989) );
  INV_X1 U6866 ( .A(n5760), .ZN(n5762) );
  NAND3_X1 U6867 ( .A1(n5763), .A2(n5762), .A3(n5761), .ZN(n5767) );
  NAND2_X1 U6868 ( .A1(n5764), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5765) );
  NAND3_X1 U6869 ( .A1(n5767), .A2(n5766), .A3(n5765), .ZN(n5768) );
  AOI21_X1 U6870 ( .B1(n5769), .B2(n6333), .A(n5768), .ZN(n5770) );
  OAI21_X1 U6871 ( .B1(n5771), .B2(n6307), .A(n5770), .ZN(U2990) );
  INV_X1 U6872 ( .A(n5772), .ZN(n5775) );
  OAI21_X1 U6873 ( .B1(n5791), .B2(n5776), .A(n5773), .ZN(n5774) );
  AOI21_X1 U6874 ( .B1(n5775), .B2(n6333), .A(n5774), .ZN(n5779) );
  XNOR2_X1 U6875 ( .A(n5776), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5777)
         );
  NAND2_X1 U6876 ( .A1(n5787), .A2(n5777), .ZN(n5778) );
  OAI211_X1 U6877 ( .C1(n5780), .C2(n6307), .A(n5779), .B(n5778), .ZN(U2992)
         );
  INV_X1 U6878 ( .A(n5781), .ZN(n5789) );
  NOR2_X1 U6879 ( .A1(n5791), .A2(n5786), .ZN(n5785) );
  OAI21_X1 U6880 ( .B1(n5783), .B2(n6309), .A(n5782), .ZN(n5784) );
  AOI211_X1 U6881 ( .C1(n5787), .C2(n5786), .A(n5785), .B(n5784), .ZN(n5788)
         );
  OAI21_X1 U6882 ( .B1(n5789), .B2(n6307), .A(n5788), .ZN(U2993) );
  AND2_X1 U6883 ( .A1(n5841), .A2(n5790), .ZN(n5808) );
  NAND3_X1 U6884 ( .A1(n5808), .A2(n5810), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5793) );
  AOI21_X1 U6885 ( .B1(n5793), .B2(n5792), .A(n5791), .ZN(n5796) );
  OAI21_X1 U6886 ( .B1(n5922), .B2(n6309), .A(n5794), .ZN(n5795) );
  INV_X1 U6887 ( .A(n5798), .ZN(U2994) );
  INV_X1 U6888 ( .A(n5799), .ZN(n5802) );
  OAI21_X1 U6889 ( .B1(n5929), .B2(n6309), .A(n5800), .ZN(n5801) );
  AOI21_X1 U6890 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5802), .A(n5801), 
        .ZN(n5805) );
  NAND3_X1 U6891 ( .A1(n5808), .A2(n5810), .A3(n5803), .ZN(n5804) );
  OAI211_X1 U6892 ( .C1(n5806), .C2(n6307), .A(n5805), .B(n5804), .ZN(U2995)
         );
  INV_X1 U6893 ( .A(n5950), .ZN(n5813) );
  OAI21_X1 U6894 ( .B1(n5817), .B2(n6709), .A(n5807), .ZN(n5812) );
  INV_X1 U6895 ( .A(n5808), .ZN(n5823) );
  NOR3_X1 U6896 ( .A1(n5823), .A2(n5810), .A3(n5809), .ZN(n5811) );
  AOI211_X1 U6897 ( .C1(n6333), .C2(n5813), .A(n5812), .B(n5811), .ZN(n5814)
         );
  OAI21_X1 U6898 ( .B1(n5815), .B2(n6307), .A(n5814), .ZN(U2996) );
  NAND2_X1 U6899 ( .A1(n5816), .A2(n6322), .ZN(n5822) );
  INV_X1 U6900 ( .A(n5817), .ZN(n5820) );
  OAI21_X1 U6901 ( .B1(n5954), .B2(n6309), .A(n5818), .ZN(n5819) );
  AOI21_X1 U6902 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5820), .A(n5819), 
        .ZN(n5821) );
  OAI211_X1 U6903 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5823), .A(n5822), .B(n5821), .ZN(U2997) );
  NAND2_X1 U6904 ( .A1(n5824), .A2(n6322), .ZN(n5835) );
  NAND2_X1 U6905 ( .A1(n5825), .A2(n5850), .ZN(n5826) );
  AND2_X1 U6906 ( .A1(n5827), .A2(n5826), .ZN(n5849) );
  INV_X1 U6907 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5847) );
  NAND2_X1 U6908 ( .A1(n6329), .A2(n5847), .ZN(n5828) );
  NAND2_X1 U6909 ( .A1(n5849), .A2(n5828), .ZN(n5836) );
  AOI21_X1 U6910 ( .B1(n5836), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5829), 
        .ZN(n5834) );
  NAND2_X1 U6911 ( .A1(n5830), .A2(n6333), .ZN(n5833) );
  OAI211_X1 U6912 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5841), .B(n5831), .ZN(n5832) );
  NAND4_X1 U6913 ( .A1(n5835), .A2(n5834), .A3(n5833), .A4(n5832), .ZN(U2998)
         );
  NAND2_X1 U6914 ( .A1(n5836), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5838) );
  OAI211_X1 U6915 ( .C1(n5839), .C2(n6309), .A(n5838), .B(n5837), .ZN(n5840)
         );
  AOI21_X1 U6916 ( .B1(n5841), .B2(n3516), .A(n5840), .ZN(n5842) );
  OAI21_X1 U6917 ( .B1(n5843), .B2(n6307), .A(n5842), .ZN(U2999) );
  OAI21_X1 U6918 ( .B1(n5846), .B2(n5845), .A(n5844), .ZN(n5848) );
  XNOR2_X1 U6919 ( .A(n5848), .B(n5847), .ZN(n5971) );
  INV_X1 U6920 ( .A(n5971), .ZN(n5855) );
  INV_X1 U6921 ( .A(n5849), .ZN(n5853) );
  OAI22_X1 U6922 ( .A1(n6061), .A2(n6309), .B1(n6535), .B2(n6308), .ZN(n5852)
         );
  NOR3_X1 U6923 ( .A1(n5983), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .A3(n5850), 
        .ZN(n5851) );
  AOI211_X1 U6924 ( .C1(INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n5853), .A(n5852), .B(n5851), .ZN(n5854) );
  OAI21_X1 U6925 ( .B1(n5855), .B2(n6307), .A(n5854), .ZN(U3000) );
  OAI21_X1 U6926 ( .B1(n5856), .B2(STATEBS16_REG_SCAN_IN), .A(n6350), .ZN(
        n5857) );
  OAI22_X1 U6927 ( .A1(n5857), .A2(n5859), .B1(n4342), .B2(n5861), .ZN(n5858)
         );
  MUX2_X1 U6928 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5858), .S(n6342), 
        .Z(U3464) );
  XNOR2_X1 U6929 ( .A(n5860), .B(n5859), .ZN(n5863) );
  OAI22_X1 U6930 ( .A1(n5863), .A2(n6347), .B1(n5862), .B2(n5861), .ZN(n5864)
         );
  MUX2_X1 U6931 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5864), .S(n6342), 
        .Z(U3463) );
  OAI22_X1 U6932 ( .A1(n5867), .A2(n6575), .B1(n5866), .B2(n5865), .ZN(n5868)
         );
  MUX2_X1 U6933 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n5868), .S(n6573), 
        .Z(U3456) );
  NOR2_X1 U6934 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5869), .ZN(n5912)
         );
  INV_X1 U6935 ( .A(n5912), .ZN(n5871) );
  AOI211_X1 U6936 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5871), .A(n6353), .B(
        n5870), .ZN(n5876) );
  OAI211_X1 U6937 ( .C1(n5874), .C2(n5881), .A(n5873), .B(n5872), .ZN(n5875)
         );
  NAND2_X1 U6938 ( .A1(n5876), .A2(n5875), .ZN(n5910) );
  NAND2_X1 U6939 ( .A1(n5910), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U6940 ( .A1(n5878), .A2(n5877), .ZN(n5880) );
  NAND2_X1 U6941 ( .A1(n3102), .A2(n6345), .ZN(n5879) );
  NAND2_X1 U6942 ( .A1(n5880), .A2(n5879), .ZN(n5911) );
  AOI22_X1 U6943 ( .A1(n6417), .A2(n5912), .B1(n6419), .B2(n5911), .ZN(n5884)
         );
  OR2_X1 U6944 ( .A1(n5913), .A2(n6361), .ZN(n5883) );
  NAND2_X1 U6945 ( .A1(n5914), .A2(n6358), .ZN(n5882) );
  NAND4_X1 U6946 ( .A1(n5885), .A2(n5884), .A3(n5883), .A4(n5882), .ZN(U3052)
         );
  NAND2_X1 U6947 ( .A1(n5910), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5889) );
  AOI22_X1 U6948 ( .A1(n6423), .A2(n5912), .B1(n6425), .B2(n5911), .ZN(n5888)
         );
  OR2_X1 U6949 ( .A1(n5913), .A2(n6365), .ZN(n5887) );
  NAND2_X1 U6950 ( .A1(n5914), .A2(n6362), .ZN(n5886) );
  NAND4_X1 U6951 ( .A1(n5889), .A2(n5888), .A3(n5887), .A4(n5886), .ZN(U3053)
         );
  NAND2_X1 U6952 ( .A1(n5910), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5893) );
  AOI22_X1 U6953 ( .A1(n6367), .A2(n5912), .B1(n6366), .B2(n5911), .ZN(n5892)
         );
  OR2_X1 U6954 ( .A1(n5913), .A2(n6371), .ZN(n5891) );
  NAND2_X1 U6955 ( .A1(n5914), .A2(n6368), .ZN(n5890) );
  NAND4_X1 U6956 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), .ZN(U3054)
         );
  NAND2_X1 U6957 ( .A1(n5910), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5897) );
  AOI22_X1 U6958 ( .A1(n6401), .A2(n5912), .B1(n6402), .B2(n5911), .ZN(n5896)
         );
  OR2_X1 U6959 ( .A1(n5913), .A2(n6375), .ZN(n5895) );
  NAND2_X1 U6960 ( .A1(n5914), .A2(n6372), .ZN(n5894) );
  NAND4_X1 U6961 ( .A1(n5897), .A2(n5896), .A3(n5895), .A4(n5894), .ZN(U3055)
         );
  NAND2_X1 U6962 ( .A1(n5910), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5901) );
  AOI22_X1 U6963 ( .A1(n6377), .A2(n5912), .B1(n6376), .B2(n5911), .ZN(n5900)
         );
  OR2_X1 U6964 ( .A1(n5913), .A2(n6381), .ZN(n5899) );
  NAND2_X1 U6965 ( .A1(n5914), .A2(n6378), .ZN(n5898) );
  NAND4_X1 U6966 ( .A1(n5901), .A2(n5900), .A3(n5899), .A4(n5898), .ZN(U3056)
         );
  NAND2_X1 U6967 ( .A1(n5910), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5905) );
  AOI22_X1 U6968 ( .A1(n6429), .A2(n5912), .B1(n6431), .B2(n5911), .ZN(n5904)
         );
  OR2_X1 U6969 ( .A1(n5913), .A2(n6385), .ZN(n5903) );
  NAND2_X1 U6970 ( .A1(n5914), .A2(n6382), .ZN(n5902) );
  NAND4_X1 U6971 ( .A1(n5905), .A2(n5904), .A3(n5903), .A4(n5902), .ZN(U3057)
         );
  NAND2_X1 U6972 ( .A1(n5910), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5909) );
  AOI22_X1 U6973 ( .A1(n6409), .A2(n5912), .B1(n6411), .B2(n5911), .ZN(n5908)
         );
  OR2_X1 U6974 ( .A1(n5913), .A2(n6389), .ZN(n5907) );
  NAND2_X1 U6975 ( .A1(n5914), .A2(n6386), .ZN(n5906) );
  NAND4_X1 U6976 ( .A1(n5909), .A2(n5908), .A3(n5907), .A4(n5906), .ZN(U3058)
         );
  NAND2_X1 U6977 ( .A1(n5910), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5918) );
  AOI22_X1 U6978 ( .A1(n6436), .A2(n5912), .B1(n6440), .B2(n5911), .ZN(n5917)
         );
  OR2_X1 U6979 ( .A1(n5913), .A2(n6397), .ZN(n5916) );
  NAND2_X1 U6980 ( .A1(n5914), .A2(n6393), .ZN(n5915) );
  NAND4_X1 U6981 ( .A1(n5918), .A2(n5917), .A3(n5916), .A4(n5915), .ZN(U3059)
         );
  AND2_X1 U6982 ( .A1(n6229), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6983 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n6178), .B1(n6180), 
        .B2(n5919), .ZN(n5921) );
  NAND2_X1 U6984 ( .A1(n6172), .A2(EBX_REG_24__SCAN_IN), .ZN(n5920) );
  OAI211_X1 U6985 ( .C1(n5922), .C2(n6175), .A(n5921), .B(n5920), .ZN(n5925)
         );
  NOR2_X1 U6986 ( .A1(n5923), .A2(n6151), .ZN(n5924) );
  OAI21_X1 U6987 ( .B1(REIP_REG_24__SCAN_IN), .B2(n5927), .A(n5926), .ZN(U2803) );
  AOI22_X1 U6988 ( .A1(EBX_REG_23__SCAN_IN), .A2(n6172), .B1(n5928), .B2(n6180), .ZN(n5935) );
  OAI22_X1 U6989 ( .A1(n5930), .A2(n6151), .B1(n5929), .B2(n6175), .ZN(n5931)
         );
  OAI211_X1 U6990 ( .C1(n5936), .C2(n6115), .A(n5935), .B(n5934), .ZN(U2804)
         );
  INV_X1 U6991 ( .A(n5937), .ZN(n5941) );
  INV_X1 U6992 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5939) );
  OR2_X1 U6993 ( .A1(n6138), .A2(n5938), .ZN(n5969) );
  INV_X1 U6994 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6541) );
  OAI22_X1 U6995 ( .A1(n6115), .A2(n5939), .B1(n5969), .B2(n6541), .ZN(n5940)
         );
  AOI21_X1 U6996 ( .B1(n5941), .B2(n6180), .A(n5940), .ZN(n5942) );
  OAI21_X1 U6997 ( .B1(n6169), .B2(n5943), .A(n5942), .ZN(n5944) );
  AOI21_X1 U6998 ( .B1(n5945), .B2(n6143), .A(n5944), .ZN(n5949) );
  INV_X1 U6999 ( .A(n5959), .ZN(n5947) );
  OAI211_X1 U7000 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5947), .B(n5946), .ZN(n5948) );
  OAI211_X1 U7001 ( .C1(n6175), .C2(n5950), .A(n5949), .B(n5948), .ZN(U2805)
         );
  INV_X1 U7002 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6540) );
  AOI22_X1 U7003 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6172), .B1(n5951), .B2(n6180), .ZN(n5952) );
  OAI21_X1 U7004 ( .B1(n6540), .B2(n5969), .A(n5952), .ZN(n5953) );
  AOI21_X1 U7005 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6178), .A(n5953), 
        .ZN(n5958) );
  OAI22_X1 U7006 ( .A1(n5955), .A2(n6151), .B1(n6175), .B2(n5954), .ZN(n5956)
         );
  INV_X1 U7007 ( .A(n5956), .ZN(n5957) );
  OAI211_X1 U7008 ( .C1(REIP_REG_21__SCAN_IN), .C2(n5959), .A(n5958), .B(n5957), .ZN(U2806) );
  AOI21_X1 U7009 ( .B1(n5960), .B2(REIP_REG_19__SCAN_IN), .A(
        REIP_REG_20__SCAN_IN), .ZN(n5970) );
  INV_X1 U7010 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5962) );
  OAI22_X1 U7011 ( .A1(n5962), .A2(n6115), .B1(n5961), .B2(n6161), .ZN(n5963)
         );
  AOI21_X1 U7012 ( .B1(EBX_REG_20__SCAN_IN), .B2(n6172), .A(n5963), .ZN(n5968)
         );
  OAI22_X1 U7013 ( .A1(n5965), .A2(n6151), .B1(n6175), .B2(n5964), .ZN(n5966)
         );
  INV_X1 U7014 ( .A(n5966), .ZN(n5967) );
  OAI211_X1 U7015 ( .C1(n5970), .C2(n5969), .A(n5968), .B(n5967), .ZN(U2807)
         );
  AOI22_X1 U7016 ( .A1(n6284), .A2(REIP_REG_18__SCAN_IN), .B1(n6300), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5973) );
  AOI22_X1 U7017 ( .A1(n5971), .A2(n6289), .B1(n6287), .B2(n6196), .ZN(n5972)
         );
  OAI211_X1 U7018 ( .C1(n6294), .C2(n6053), .A(n5973), .B(n5972), .ZN(U2968)
         );
  INV_X1 U7019 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5978) );
  OAI21_X1 U7020 ( .B1(n5975), .B2(n5974), .A(n5392), .ZN(n6017) );
  INV_X1 U7021 ( .A(n6103), .ZN(n5976) );
  AOI222_X1 U7022 ( .A1(n6017), .A2(n6289), .B1(n5976), .B2(n6276), .C1(n6287), 
        .C2(n6100), .ZN(n5977) );
  NAND2_X1 U7023 ( .A1(n6284), .A2(REIP_REG_13__SCAN_IN), .ZN(n6022) );
  OAI211_X1 U7024 ( .C1(n5978), .C2(n6282), .A(n5977), .B(n6022), .ZN(U2973)
         );
  AOI22_X1 U7025 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5979), .B1(n6284), .B2(REIP_REG_17__SCAN_IN), .ZN(n5982) );
  AOI22_X1 U7026 ( .A1(n5980), .A2(n6322), .B1(n6333), .B2(n6068), .ZN(n5981)
         );
  OAI211_X1 U7027 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5983), .A(n5982), .B(n5981), .ZN(U3001) );
  OAI21_X1 U7028 ( .B1(n5985), .B2(n5987), .A(n5984), .ZN(n5986) );
  INV_X1 U7029 ( .A(n5986), .ZN(n6001) );
  NAND2_X1 U7030 ( .A1(n5987), .A2(n6002), .ZN(n5993) );
  AOI221_X1 U7031 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n6000), .C2(n5992), .A(n5993), 
        .ZN(n5990) );
  OAI22_X1 U7032 ( .A1(n5988), .A2(n6307), .B1(n6309), .B2(n6082), .ZN(n5989)
         );
  AOI211_X1 U7033 ( .C1(REIP_REG_16__SCAN_IN), .C2(n6284), .A(n5990), .B(n5989), .ZN(n5991) );
  OAI21_X1 U7034 ( .B1(n6001), .B2(n5992), .A(n5991), .ZN(U3002) );
  OAI22_X1 U7035 ( .A1(n6532), .A2(n6308), .B1(n5993), .B2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5994) );
  INV_X1 U7036 ( .A(n5994), .ZN(n5999) );
  INV_X1 U7037 ( .A(n5995), .ZN(n5997) );
  AOI22_X1 U7038 ( .A1(n5997), .A2(n6322), .B1(n6333), .B2(n5996), .ZN(n5998)
         );
  OAI211_X1 U7039 ( .C1(n6001), .C2(n6000), .A(n5999), .B(n5998), .ZN(U3003)
         );
  NAND2_X1 U7040 ( .A1(n6003), .A2(n6002), .ZN(n6015) );
  NAND2_X1 U7041 ( .A1(n6009), .A2(n6004), .ZN(n6025) );
  NOR2_X1 U7042 ( .A1(n6005), .A2(n6025), .ZN(n6019) );
  AOI211_X1 U7043 ( .C1(n6007), .C2(n6016), .A(n6019), .B(n6006), .ZN(n6008)
         );
  OAI21_X1 U7044 ( .B1(n6010), .B2(n6009), .A(n6008), .ZN(n6021) );
  OAI22_X1 U7045 ( .A1(n6011), .A2(n6307), .B1(n6309), .B2(n6084), .ZN(n6012)
         );
  AOI21_X1 U7046 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n6021), .A(n6012), 
        .ZN(n6014) );
  NAND2_X1 U7047 ( .A1(n6284), .A2(REIP_REG_14__SCAN_IN), .ZN(n6013) );
  OAI211_X1 U7048 ( .C1(n6016), .C2(n6015), .A(n6014), .B(n6013), .ZN(U3004)
         );
  INV_X1 U7049 ( .A(n6017), .ZN(n6018) );
  OAI22_X1 U7050 ( .A1(n6018), .A2(n6307), .B1(n6309), .B2(n6098), .ZN(n6020)
         );
  AOI211_X1 U7051 ( .C1(n6021), .C2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n6020), .B(n6019), .ZN(n6023) );
  OAI211_X1 U7052 ( .C1(n6025), .C2(n6024), .A(n6023), .B(n6022), .ZN(U3005)
         );
  OR4_X1 U7053 ( .A1(n6027), .A2(n6026), .A3(n6575), .A4(n2999), .ZN(n6028) );
  OAI21_X1 U7054 ( .B1(n6573), .B2(n3779), .A(n6028), .ZN(U3455) );
  INV_X1 U7055 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6512) );
  AOI21_X1 U7056 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6512), .A(n6506), .ZN(n6035) );
  INV_X1 U7057 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6029) );
  INV_X1 U7058 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6502) );
  NOR2_X1 U7059 ( .A1(n6502), .A2(STATE_REG_0__SCAN_IN), .ZN(n6559) );
  AOI21_X1 U7060 ( .B1(n6035), .B2(n6029), .A(n6559), .ZN(U2789) );
  INV_X1 U7061 ( .A(n6030), .ZN(n6031) );
  OAI21_X1 U7062 ( .B1(n6031), .B2(n6486), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6032) );
  OAI21_X1 U7063 ( .B1(n6033), .B2(n6479), .A(n6032), .ZN(U2790) );
  NOR2_X1 U7064 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6036) );
  OAI21_X1 U7065 ( .B1(n6036), .B2(D_C_N_REG_SCAN_IN), .A(n6597), .ZN(n6034)
         );
  OAI21_X1 U7066 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6597), .A(n6034), .ZN(
        U2791) );
  NOR2_X1 U7067 ( .A1(n6559), .A2(n6035), .ZN(n6563) );
  OAI21_X1 U7068 ( .B1(n6036), .B2(BS16_N), .A(n6563), .ZN(n6561) );
  OAI21_X1 U7069 ( .B1(n6563), .B2(n6760), .A(n6561), .ZN(U2792) );
  OAI21_X1 U7070 ( .B1(n6038), .B2(n6037), .A(n6297), .ZN(U2793) );
  NOR4_X1 U7071 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(
        DATAWIDTH_REG_18__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n6042) );
  NOR4_X1 U7072 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_16__SCAN_IN), .ZN(n6041) );
  NOR4_X1 U7073 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6040) );
  NOR4_X1 U7074 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n6039) );
  NAND4_X1 U7075 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n6048)
         );
  NOR4_X1 U7076 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6046) );
  AOI211_X1 U7077 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_30__SCAN_IN), .B(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n6045) );
  NOR4_X1 U7078 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6044)
         );
  NOR4_X1 U7079 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n6043) );
  NAND4_X1 U7080 ( .A1(n6046), .A2(n6045), .A3(n6044), .A4(n6043), .ZN(n6047)
         );
  NOR2_X1 U7081 ( .A1(n6048), .A2(n6047), .ZN(n6580) );
  INV_X1 U7082 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n6050) );
  NOR3_X1 U7083 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6051) );
  OAI21_X1 U7084 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6051), .A(n6580), .ZN(n6049)
         );
  OAI21_X1 U7085 ( .B1(n6580), .B2(n6050), .A(n6049), .ZN(U2794) );
  INV_X1 U7086 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6562) );
  AOI21_X1 U7087 ( .B1(n5251), .B2(n6562), .A(n6051), .ZN(n6052) );
  INV_X1 U7088 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6558) );
  INV_X1 U7089 ( .A(n6580), .ZN(n6583) );
  AOI22_X1 U7090 ( .A1(n6580), .A2(n6052), .B1(n6558), .B2(n6583), .ZN(U2795)
         );
  INV_X1 U7091 ( .A(n6053), .ZN(n6056) );
  AOI22_X1 U7092 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6172), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6178), .ZN(n6054) );
  OAI211_X1 U7093 ( .C1(n6071), .C2(n6535), .A(n6054), .B(n6160), .ZN(n6055)
         );
  AOI21_X1 U7094 ( .B1(n6180), .B2(n6056), .A(n6055), .ZN(n6057) );
  OAI21_X1 U7095 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6058), .A(n6057), .ZN(n6059) );
  AOI21_X1 U7096 ( .B1(n6196), .B2(n6143), .A(n6059), .ZN(n6060) );
  OAI21_X1 U7097 ( .B1(n6175), .B2(n6061), .A(n6060), .ZN(U2809) );
  NOR2_X1 U7098 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6062), .ZN(n6072) );
  OAI22_X1 U7099 ( .A1(n6169), .A2(n6064), .B1(n6063), .B2(n6115), .ZN(n6065)
         );
  AOI211_X1 U7100 ( .C1(n6180), .C2(n6066), .A(n6177), .B(n6065), .ZN(n6070)
         );
  INV_X1 U7101 ( .A(n6067), .ZN(n6199) );
  AOI22_X1 U7102 ( .A1(n6199), .A2(n6143), .B1(n6158), .B2(n6068), .ZN(n6069)
         );
  OAI211_X1 U7103 ( .C1(n6072), .C2(n6071), .A(n6070), .B(n6069), .ZN(U2810)
         );
  OAI21_X1 U7104 ( .B1(n6138), .B2(n6074), .A(n6073), .ZN(n6075) );
  AOI22_X1 U7105 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6172), .B1(
        REIP_REG_16__SCAN_IN), .B2(n6075), .ZN(n6081) );
  AOI22_X1 U7106 ( .A1(PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n6178), .B1(n6076), 
        .B2(n6180), .ZN(n6077) );
  OAI211_X1 U7107 ( .C1(REIP_REG_16__SCAN_IN), .C2(n6078), .A(n6077), .B(n6160), .ZN(n6079) );
  AOI21_X1 U7108 ( .B1(n6204), .B2(n6143), .A(n6079), .ZN(n6080) );
  OAI211_X1 U7109 ( .C1(n6175), .C2(n6082), .A(n6081), .B(n6080), .ZN(U2811)
         );
  AOI22_X1 U7110 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6172), .B1(
        REIP_REG_14__SCAN_IN), .B2(n6083), .ZN(n6093) );
  NOR2_X1 U7111 ( .A1(n6185), .A2(REIP_REG_14__SCAN_IN), .ZN(n6087) );
  OAI22_X1 U7112 ( .A1(n6757), .A2(n6115), .B1(n6175), .B2(n6084), .ZN(n6085)
         );
  AOI21_X1 U7113 ( .B1(n6087), .B2(n6086), .A(n6085), .ZN(n6092) );
  INV_X1 U7114 ( .A(n6088), .ZN(n6090) );
  AOI22_X1 U7115 ( .A1(n6090), .A2(n6143), .B1(n6180), .B2(n6089), .ZN(n6091)
         );
  NAND4_X1 U7116 ( .A1(n6093), .A2(n6092), .A3(n6091), .A4(n6160), .ZN(U2813)
         );
  AOI22_X1 U7117 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6172), .B1(
        REIP_REG_13__SCAN_IN), .B2(n6106), .ZN(n6102) );
  OAI211_X1 U7118 ( .C1(REIP_REG_13__SCAN_IN), .C2(REIP_REG_12__SCAN_IN), .A(
        n6095), .B(n6094), .ZN(n6097) );
  AOI21_X1 U7119 ( .B1(n6178), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6177), 
        .ZN(n6096) );
  OAI211_X1 U7120 ( .C1(n6175), .C2(n6098), .A(n6097), .B(n6096), .ZN(n6099)
         );
  AOI21_X1 U7121 ( .B1(n6100), .B2(n6143), .A(n6099), .ZN(n6101) );
  OAI211_X1 U7122 ( .C1(n6103), .C2(n6161), .A(n6102), .B(n6101), .ZN(U2814)
         );
  AOI22_X1 U7123 ( .A1(EBX_REG_11__SCAN_IN), .A2(n6172), .B1(
        PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n6178), .ZN(n6111) );
  AOI21_X1 U7124 ( .B1(n6158), .B2(n6104), .A(n6177), .ZN(n6110) );
  INV_X1 U7125 ( .A(n6105), .ZN(n6265) );
  AOI22_X1 U7126 ( .A1(n6265), .A2(n6143), .B1(n6180), .B2(n6264), .ZN(n6109)
         );
  INV_X1 U7127 ( .A(n6135), .ZN(n6154) );
  OAI221_X1 U7128 ( .B1(REIP_REG_11__SCAN_IN), .B2(n6107), .C1(
        REIP_REG_11__SCAN_IN), .C2(n6154), .A(n6106), .ZN(n6108) );
  NAND4_X1 U7129 ( .A1(n6111), .A2(n6110), .A3(n6109), .A4(n6108), .ZN(U2816)
         );
  NOR2_X1 U7130 ( .A1(n6112), .A2(n6135), .ZN(n6117) );
  AOI22_X1 U7131 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6172), .B1(n6158), .B2(n6320), 
        .ZN(n6113) );
  OAI211_X1 U7132 ( .C1(n6115), .C2(n6114), .A(n6113), .B(n6160), .ZN(n6116)
         );
  AOI221_X1 U7133 ( .B1(n6117), .B2(n6722), .C1(n6124), .C2(
        REIP_REG_9__SCAN_IN), .A(n6116), .ZN(n6123) );
  INV_X1 U7134 ( .A(n6118), .ZN(n6119) );
  OAI22_X1 U7135 ( .A1(n6120), .A2(n6151), .B1(n6161), .B2(n6119), .ZN(n6121)
         );
  INV_X1 U7136 ( .A(n6121), .ZN(n6122) );
  NAND2_X1 U7137 ( .A1(n6123), .A2(n6122), .ZN(U2818) );
  INV_X1 U7138 ( .A(n6124), .ZN(n6134) );
  INV_X1 U7139 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6521) );
  NOR2_X1 U7140 ( .A1(n6710), .A2(n6521), .ZN(n6136) );
  AOI21_X1 U7141 ( .B1(n6136), .B2(n6154), .A(REIP_REG_8__SCAN_IN), .ZN(n6133)
         );
  OAI22_X1 U7142 ( .A1(n6169), .A2(n6126), .B1(n6175), .B2(n6125), .ZN(n6127)
         );
  AOI211_X1 U7143 ( .C1(n6178), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6177), 
        .B(n6127), .ZN(n6132) );
  NOR2_X1 U7144 ( .A1(n6161), .A2(n6128), .ZN(n6129) );
  AOI21_X1 U7145 ( .B1(n6130), .B2(n6143), .A(n6129), .ZN(n6131) );
  OAI211_X1 U7146 ( .C1(n6134), .C2(n6133), .A(n6132), .B(n6131), .ZN(U2819)
         );
  AOI211_X1 U7147 ( .C1(n6710), .C2(n6521), .A(n6136), .B(n6135), .ZN(n6142)
         );
  NOR2_X1 U7148 ( .A1(n6138), .A2(n6137), .ZN(n6165) );
  AOI22_X1 U7149 ( .A1(PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n6178), .B1(
        REIP_REG_7__SCAN_IN), .B2(n6165), .ZN(n6139) );
  OAI211_X1 U7150 ( .C1(n6175), .C2(n6140), .A(n6139), .B(n6160), .ZN(n6141)
         );
  AOI211_X1 U7151 ( .C1(EBX_REG_7__SCAN_IN), .C2(n6172), .A(n6142), .B(n6141), 
        .ZN(n6145) );
  NAND2_X1 U7152 ( .A1(n6271), .A2(n6143), .ZN(n6144) );
  OAI211_X1 U7153 ( .C1(n6161), .C2(n6269), .A(n6145), .B(n6144), .ZN(U2820)
         );
  OAI22_X1 U7154 ( .A1(n6169), .A2(n6147), .B1(n6175), .B2(n6146), .ZN(n6148)
         );
  AOI211_X1 U7155 ( .C1(n6178), .C2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6177), 
        .B(n6148), .ZN(n6156) );
  INV_X1 U7156 ( .A(n6149), .ZN(n6150) );
  OAI22_X1 U7157 ( .A1(n6152), .A2(n6151), .B1(n6150), .B2(n6161), .ZN(n6153)
         );
  AOI221_X1 U7158 ( .B1(n6165), .B2(REIP_REG_6__SCAN_IN), .C1(n6154), .C2(
        n6710), .A(n6153), .ZN(n6155) );
  NAND2_X1 U7159 ( .A1(n6156), .A2(n6155), .ZN(U2821) );
  INV_X1 U7160 ( .A(n6157), .ZN(n6182) );
  AOI22_X1 U7161 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n6178), .B1(n6158), 
        .B2(n6190), .ZN(n6159) );
  OAI211_X1 U7162 ( .C1(n6275), .C2(n6161), .A(n6160), .B(n6159), .ZN(n6162)
         );
  AOI21_X1 U7163 ( .B1(n6278), .B2(n6182), .A(n6162), .ZN(n6168) );
  AND2_X1 U7164 ( .A1(n6164), .A2(n6163), .ZN(n6166) );
  OAI21_X1 U7165 ( .B1(REIP_REG_5__SCAN_IN), .B2(n6166), .A(n6165), .ZN(n6167)
         );
  OAI211_X1 U7166 ( .C1(n6169), .C2(n6194), .A(n6168), .B(n6167), .ZN(U2822)
         );
  AOI22_X1 U7167 ( .A1(EBX_REG_4__SCAN_IN), .A2(n6172), .B1(n6171), .B2(n6170), 
        .ZN(n6189) );
  OAI22_X1 U7168 ( .A1(n6175), .A2(n6174), .B1(n6517), .B2(n6173), .ZN(n6176)
         );
  AOI211_X1 U7169 ( .C1(n6178), .C2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n6177), 
        .B(n6176), .ZN(n6188) );
  INV_X1 U7170 ( .A(n6179), .ZN(n6181) );
  AOI22_X1 U7171 ( .A1(n6183), .A2(n6182), .B1(n6181), .B2(n6180), .ZN(n6187)
         );
  OR3_X1 U7172 ( .A1(n6185), .A2(n6184), .A3(REIP_REG_4__SCAN_IN), .ZN(n6186)
         );
  NAND4_X1 U7173 ( .A1(n6189), .A2(n6188), .A3(n6187), .A4(n6186), .ZN(U2823)
         );
  AOI22_X1 U7174 ( .A1(n6278), .A2(n6192), .B1(n6191), .B2(n6190), .ZN(n6193)
         );
  OAI21_X1 U7175 ( .B1(n6195), .B2(n6194), .A(n6193), .ZN(U2854) );
  AOI22_X1 U7176 ( .A1(n6196), .A2(n6203), .B1(n6202), .B2(DATAI_18_), .ZN(
        n6198) );
  AOI22_X1 U7177 ( .A1(n6206), .A2(DATAI_2_), .B1(n6205), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U7178 ( .A1(n6198), .A2(n6197), .ZN(U2873) );
  AOI22_X1 U7179 ( .A1(n6199), .A2(n6203), .B1(n6202), .B2(DATAI_17_), .ZN(
        n6201) );
  AOI22_X1 U7180 ( .A1(n6206), .A2(DATAI_1_), .B1(n6205), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7181 ( .A1(n6201), .A2(n6200), .ZN(U2874) );
  AOI22_X1 U7182 ( .A1(n6204), .A2(n6203), .B1(n6202), .B2(DATAI_16_), .ZN(
        n6208) );
  AOI22_X1 U7183 ( .A1(n6206), .A2(DATAI_0_), .B1(n6205), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7184 ( .A1(n6208), .A2(n6207), .ZN(U2875) );
  INV_X1 U7185 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6263) );
  AOI22_X1 U7186 ( .A1(LWORD_REG_15__SCAN_IN), .A2(n6588), .B1(n6229), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6210) );
  OAI21_X1 U7187 ( .B1(n6263), .B2(n6241), .A(n6210), .ZN(U2908) );
  INV_X1 U7188 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6212) );
  AOI22_X1 U7189 ( .A1(LWORD_REG_14__SCAN_IN), .A2(n6588), .B1(n6229), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6211) );
  OAI21_X1 U7190 ( .B1(n6212), .B2(n6241), .A(n6211), .ZN(U2909) );
  INV_X1 U7191 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6214) );
  AOI22_X1 U7192 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6588), .B1(n6229), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6213) );
  OAI21_X1 U7193 ( .B1(n6214), .B2(n6241), .A(n6213), .ZN(U2910) );
  INV_X1 U7194 ( .A(EAX_REG_12__SCAN_IN), .ZN(n6216) );
  AOI22_X1 U7195 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n6588), .B1(n6229), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6215) );
  OAI21_X1 U7196 ( .B1(n6216), .B2(n6241), .A(n6215), .ZN(U2911) );
  INV_X1 U7197 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6218) );
  AOI22_X1 U7198 ( .A1(LWORD_REG_11__SCAN_IN), .A2(n6588), .B1(n6229), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6217) );
  OAI21_X1 U7199 ( .B1(n6218), .B2(n6241), .A(n6217), .ZN(U2912) );
  INV_X1 U7200 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6220) );
  AOI22_X1 U7201 ( .A1(LWORD_REG_10__SCAN_IN), .A2(n6588), .B1(n6229), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6219) );
  OAI21_X1 U7202 ( .B1(n6220), .B2(n6241), .A(n6219), .ZN(U2913) );
  INV_X1 U7203 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6222) );
  AOI22_X1 U7204 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n6588), .B1(n6229), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6221) );
  OAI21_X1 U7205 ( .B1(n6222), .B2(n6241), .A(n6221), .ZN(U2914) );
  INV_X1 U7206 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6224) );
  AOI22_X1 U7207 ( .A1(LWORD_REG_8__SCAN_IN), .A2(n6588), .B1(n6229), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6223) );
  OAI21_X1 U7208 ( .B1(n6224), .B2(n6241), .A(n6223), .ZN(U2915) );
  AOI22_X1 U7209 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6239), .B1(n6229), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6225) );
  OAI21_X1 U7210 ( .B1(n3838), .B2(n6241), .A(n6225), .ZN(U2916) );
  AOI22_X1 U7211 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6239), .B1(n6229), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6226) );
  OAI21_X1 U7212 ( .B1(n6227), .B2(n6241), .A(n6226), .ZN(U2917) );
  INV_X1 U7213 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6756) );
  AOI22_X1 U7214 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6239), .B1(n6229), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6228) );
  OAI21_X1 U7215 ( .B1(n6756), .B2(n6241), .A(n6228), .ZN(U2918) );
  AOI22_X1 U7216 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6239), .B1(n6229), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6230) );
  OAI21_X1 U7217 ( .B1(n6231), .B2(n6241), .A(n6230), .ZN(U2919) );
  AOI22_X1 U7218 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6239), .B1(n6238), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6232) );
  OAI21_X1 U7219 ( .B1(n6233), .B2(n6241), .A(n6232), .ZN(U2920) );
  AOI22_X1 U7220 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6239), .B1(n6238), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6234) );
  OAI21_X1 U7221 ( .B1(n6235), .B2(n6241), .A(n6234), .ZN(U2921) );
  AOI22_X1 U7222 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n6239), .B1(n6238), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6236) );
  OAI21_X1 U7223 ( .B1(n6237), .B2(n6241), .A(n6236), .ZN(U2922) );
  AOI22_X1 U7224 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n6239), .B1(n6238), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6240) );
  OAI21_X1 U7225 ( .B1(n6242), .B2(n6241), .A(n6240), .ZN(U2923) );
  AOI22_X1 U7226 ( .A1(EAX_REG_24__SCAN_IN), .A2(n6256), .B1(n6259), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n6243) );
  NAND2_X1 U7227 ( .A1(n6260), .A2(DATAI_8_), .ZN(n6248) );
  NAND2_X1 U7228 ( .A1(n6243), .A2(n6248), .ZN(U2932) );
  AOI22_X1 U7229 ( .A1(EAX_REG_25__SCAN_IN), .A2(n6256), .B1(n6259), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n6244) );
  NAND2_X1 U7230 ( .A1(n6260), .A2(DATAI_9_), .ZN(n6250) );
  NAND2_X1 U7231 ( .A1(n6244), .A2(n6250), .ZN(U2933) );
  AOI22_X1 U7232 ( .A1(EAX_REG_26__SCAN_IN), .A2(n6256), .B1(n6259), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6245) );
  NAND2_X1 U7233 ( .A1(n6260), .A2(DATAI_10_), .ZN(n6252) );
  NAND2_X1 U7234 ( .A1(n6245), .A2(n6252), .ZN(U2934) );
  AOI22_X1 U7235 ( .A1(EAX_REG_27__SCAN_IN), .A2(n6256), .B1(n6259), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n6246) );
  NAND2_X1 U7236 ( .A1(n6260), .A2(DATAI_11_), .ZN(n6254) );
  NAND2_X1 U7237 ( .A1(n6246), .A2(n6254), .ZN(U2935) );
  AOI22_X1 U7238 ( .A1(EAX_REG_29__SCAN_IN), .A2(n6256), .B1(n6259), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n6247) );
  NAND2_X1 U7239 ( .A1(n6260), .A2(DATAI_13_), .ZN(n6257) );
  NAND2_X1 U7240 ( .A1(n6247), .A2(n6257), .ZN(U2937) );
  AOI22_X1 U7241 ( .A1(EAX_REG_8__SCAN_IN), .A2(n6256), .B1(n6259), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n6249) );
  NAND2_X1 U7242 ( .A1(n6249), .A2(n6248), .ZN(U2947) );
  AOI22_X1 U7243 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6256), .B1(n6259), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U7244 ( .A1(n6251), .A2(n6250), .ZN(U2948) );
  AOI22_X1 U7245 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6256), .B1(n6259), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6253) );
  NAND2_X1 U7246 ( .A1(n6253), .A2(n6252), .ZN(U2949) );
  AOI22_X1 U7247 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6256), .B1(n6259), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7248 ( .A1(n6255), .A2(n6254), .ZN(U2950) );
  AOI22_X1 U7249 ( .A1(EAX_REG_13__SCAN_IN), .A2(n6256), .B1(n6259), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6258) );
  NAND2_X1 U7250 ( .A1(n6258), .A2(n6257), .ZN(U2952) );
  AOI22_X1 U7251 ( .A1(n6260), .A2(DATAI_15_), .B1(n6259), .B2(
        LWORD_REG_15__SCAN_IN), .ZN(n6261) );
  OAI21_X1 U7252 ( .B1(n6263), .B2(n6262), .A(n6261), .ZN(U2954) );
  AOI22_X1 U7253 ( .A1(n6284), .A2(REIP_REG_11__SCAN_IN), .B1(n6300), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6267) );
  AOI22_X1 U7254 ( .A1(n6265), .A2(n6287), .B1(n6276), .B2(n6264), .ZN(n6266)
         );
  OAI211_X1 U7255 ( .C1(n6268), .C2(n6297), .A(n6267), .B(n6266), .ZN(U2975)
         );
  INV_X1 U7256 ( .A(n6269), .ZN(n6270) );
  AOI222_X1 U7257 ( .A1(n6272), .A2(n6289), .B1(n6271), .B2(n6287), .C1(n6270), 
        .C2(n6276), .ZN(n6274) );
  OAI211_X1 U7258 ( .C1(n6737), .C2(n6282), .A(n6274), .B(n6273), .ZN(U2979)
         );
  INV_X1 U7259 ( .A(n6275), .ZN(n6277) );
  AOI222_X1 U7260 ( .A1(n6279), .A2(n6289), .B1(n6278), .B2(n6287), .C1(n6277), 
        .C2(n6276), .ZN(n6281) );
  OAI211_X1 U7261 ( .C1(n6283), .C2(n6282), .A(n6281), .B(n6280), .ZN(U2981)
         );
  AOI22_X1 U7262 ( .A1(n6284), .A2(REIP_REG_2__SCAN_IN), .B1(n6300), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6292) );
  INV_X1 U7263 ( .A(n6285), .ZN(n6290) );
  INV_X1 U7264 ( .A(n6286), .ZN(n6288) );
  AOI22_X1 U7265 ( .A1(n6290), .A2(n6289), .B1(n6288), .B2(n6287), .ZN(n6291)
         );
  OAI211_X1 U7266 ( .C1(n6294), .C2(n6293), .A(n6292), .B(n6291), .ZN(U2984)
         );
  OAI21_X1 U7267 ( .B1(n6297), .B2(n6296), .A(n6295), .ZN(n6298) );
  INV_X1 U7268 ( .A(n6298), .ZN(n6302) );
  OAI21_X1 U7269 ( .B1(n6300), .B2(n6299), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6301) );
  OAI211_X1 U7270 ( .C1(n6304), .C2(n6303), .A(n6302), .B(n6301), .ZN(U2986)
         );
  AOI21_X1 U7271 ( .B1(n6329), .B2(n6313), .A(n6305), .ZN(n6327) );
  OAI222_X1 U7272 ( .A1(n6310), .A2(n6309), .B1(n6308), .B2(n6525), .C1(n6307), 
        .C2(n6306), .ZN(n6311) );
  INV_X1 U7273 ( .A(n6311), .ZN(n6316) );
  NOR2_X1 U7274 ( .A1(n6313), .A2(n6312), .ZN(n6321) );
  OAI211_X1 U7275 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A(n6321), .B(n6314), .ZN(n6315) );
  OAI211_X1 U7276 ( .C1(n6327), .C2(n6317), .A(n6316), .B(n6315), .ZN(U3008)
         );
  INV_X1 U7277 ( .A(n6318), .ZN(n6319) );
  AOI21_X1 U7278 ( .B1(n6333), .B2(n6320), .A(n6319), .ZN(n6325) );
  AOI22_X1 U7279 ( .A1(n6323), .A2(n6322), .B1(n6321), .B2(n6326), .ZN(n6324)
         );
  OAI211_X1 U7280 ( .C1(n6327), .C2(n6326), .A(n6325), .B(n6324), .ZN(U3009)
         );
  NAND2_X1 U7281 ( .A1(n6329), .A2(n6328), .ZN(n6341) );
  AOI21_X1 U7282 ( .B1(n6331), .B2(n6569), .A(n6330), .ZN(n6340) );
  NAND2_X1 U7283 ( .A1(n6333), .A2(n6332), .ZN(n6336) );
  NAND2_X1 U7284 ( .A1(n6334), .A2(REIP_REG_1__SCAN_IN), .ZN(n6335) );
  OAI211_X1 U7285 ( .C1(n6337), .C2(n6307), .A(n6336), .B(n6335), .ZN(n6338)
         );
  INV_X1 U7286 ( .A(n6338), .ZN(n6339) );
  OAI221_X1 U7287 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n6341), .C1(n3607), .C2(n6340), .A(n6339), .ZN(U3017) );
  NOR2_X1 U7288 ( .A1(n6738), .A2(n6342), .ZN(U3019) );
  NOR2_X1 U7289 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6343), .ZN(n6391)
         );
  NAND3_X1 U7290 ( .A1(n6345), .A2(n6344), .A3(n6357), .ZN(n6346) );
  OAI21_X1 U7291 ( .B1(n6349), .B2(n6347), .A(n6346), .ZN(n6390) );
  AOI22_X1 U7292 ( .A1(n6417), .A2(n6391), .B1(n6419), .B2(n6390), .ZN(n6360)
         );
  INV_X1 U7293 ( .A(n6415), .ZN(n6348) );
  OAI21_X1 U7294 ( .B1(n6392), .B2(n6348), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6351) );
  NAND3_X1 U7295 ( .A1(n6351), .A2(n6350), .A3(n6349), .ZN(n6356) );
  INV_X1 U7296 ( .A(n6391), .ZN(n6354) );
  AOI211_X1 U7297 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6354), .A(n6353), .B(
        n6352), .ZN(n6355) );
  NAND3_X1 U7298 ( .A1(n6357), .A2(n6356), .A3(n6355), .ZN(n6394) );
  AOI22_X1 U7299 ( .A1(n6394), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6358), 
        .B2(n6392), .ZN(n6359) );
  OAI211_X1 U7300 ( .C1(n6361), .C2(n6415), .A(n6360), .B(n6359), .ZN(U3068)
         );
  AOI22_X1 U7301 ( .A1(n6423), .A2(n6391), .B1(n6425), .B2(n6390), .ZN(n6364)
         );
  AOI22_X1 U7302 ( .A1(n6394), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6362), 
        .B2(n6392), .ZN(n6363) );
  OAI211_X1 U7303 ( .C1(n6365), .C2(n6415), .A(n6364), .B(n6363), .ZN(U3069)
         );
  AOI22_X1 U7304 ( .A1(n6367), .A2(n6391), .B1(n6366), .B2(n6390), .ZN(n6370)
         );
  AOI22_X1 U7305 ( .A1(n6394), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6368), 
        .B2(n6392), .ZN(n6369) );
  OAI211_X1 U7306 ( .C1(n6371), .C2(n6415), .A(n6370), .B(n6369), .ZN(U3070)
         );
  AOI22_X1 U7307 ( .A1(n6401), .A2(n6391), .B1(n6402), .B2(n6390), .ZN(n6374)
         );
  AOI22_X1 U7308 ( .A1(n6394), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6372), 
        .B2(n6392), .ZN(n6373) );
  OAI211_X1 U7309 ( .C1(n6375), .C2(n6415), .A(n6374), .B(n6373), .ZN(U3071)
         );
  AOI22_X1 U7310 ( .A1(n6377), .A2(n6391), .B1(n6376), .B2(n6390), .ZN(n6380)
         );
  AOI22_X1 U7311 ( .A1(n6394), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6378), 
        .B2(n6392), .ZN(n6379) );
  OAI211_X1 U7312 ( .C1(n6381), .C2(n6415), .A(n6380), .B(n6379), .ZN(U3072)
         );
  AOI22_X1 U7313 ( .A1(n6429), .A2(n6391), .B1(n6431), .B2(n6390), .ZN(n6384)
         );
  AOI22_X1 U7314 ( .A1(n6394), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6382), 
        .B2(n6392), .ZN(n6383) );
  OAI211_X1 U7315 ( .C1(n6385), .C2(n6415), .A(n6384), .B(n6383), .ZN(U3073)
         );
  AOI22_X1 U7316 ( .A1(n6409), .A2(n6391), .B1(n6411), .B2(n6390), .ZN(n6388)
         );
  AOI22_X1 U7317 ( .A1(n6394), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6386), 
        .B2(n6392), .ZN(n6387) );
  OAI211_X1 U7318 ( .C1(n6389), .C2(n6415), .A(n6388), .B(n6387), .ZN(U3074)
         );
  AOI22_X1 U7319 ( .A1(n6436), .A2(n6391), .B1(n6440), .B2(n6390), .ZN(n6396)
         );
  AOI22_X1 U7320 ( .A1(n6394), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6393), 
        .B2(n6392), .ZN(n6395) );
  OAI211_X1 U7321 ( .C1(n6397), .C2(n6415), .A(n6396), .B(n6395), .ZN(U3075)
         );
  AOI22_X1 U7322 ( .A1(n6417), .A2(n6408), .B1(n6407), .B2(n6418), .ZN(n6399)
         );
  AOI22_X1 U7323 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6412), .B1(n6419), 
        .B2(n6410), .ZN(n6398) );
  OAI211_X1 U7324 ( .C1(n6422), .C2(n6415), .A(n6399), .B(n6398), .ZN(U3076)
         );
  AOI22_X1 U7325 ( .A1(n6401), .A2(n6408), .B1(n6407), .B2(n6400), .ZN(n6404)
         );
  AOI22_X1 U7326 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6412), .B1(n6402), 
        .B2(n6410), .ZN(n6403) );
  OAI211_X1 U7327 ( .C1(n6405), .C2(n6415), .A(n6404), .B(n6403), .ZN(U3079)
         );
  AOI22_X1 U7328 ( .A1(n6409), .A2(n6408), .B1(n6407), .B2(n6406), .ZN(n6414)
         );
  AOI22_X1 U7329 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6412), .B1(n6411), 
        .B2(n6410), .ZN(n6413) );
  OAI211_X1 U7330 ( .C1(n6416), .C2(n6415), .A(n6414), .B(n6413), .ZN(U3082)
         );
  AOI22_X1 U7331 ( .A1(n6438), .A2(n6418), .B1(n6417), .B2(n6435), .ZN(n6421)
         );
  AOI22_X1 U7332 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6441), .B1(n6419), 
        .B2(n6439), .ZN(n6420) );
  OAI211_X1 U7333 ( .C1(n6422), .C2(n6444), .A(n6421), .B(n6420), .ZN(U3108)
         );
  AOI22_X1 U7334 ( .A1(n6438), .A2(n6424), .B1(n6423), .B2(n6435), .ZN(n6427)
         );
  AOI22_X1 U7335 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6441), .B1(n6425), 
        .B2(n6439), .ZN(n6426) );
  OAI211_X1 U7336 ( .C1(n6428), .C2(n6444), .A(n6427), .B(n6426), .ZN(U3109)
         );
  AOI22_X1 U7337 ( .A1(n6438), .A2(n6430), .B1(n6429), .B2(n6435), .ZN(n6433)
         );
  AOI22_X1 U7338 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6441), .B1(n6431), 
        .B2(n6439), .ZN(n6432) );
  OAI211_X1 U7339 ( .C1(n6434), .C2(n6444), .A(n6433), .B(n6432), .ZN(U3113)
         );
  AOI22_X1 U7340 ( .A1(n6438), .A2(n6437), .B1(n6436), .B2(n6435), .ZN(n6443)
         );
  AOI22_X1 U7341 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6441), .B1(n6440), 
        .B2(n6439), .ZN(n6442) );
  OAI211_X1 U7342 ( .C1(n6445), .C2(n6444), .A(n6443), .B(n6442), .ZN(U3115)
         );
  AOI21_X1 U7343 ( .B1(n6459), .B2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6470) );
  INV_X1 U7344 ( .A(n6446), .ZN(n6447) );
  AOI22_X1 U7345 ( .A1(n3036), .A2(n6448), .B1(n6447), .B2(n3076), .ZN(n6571)
         );
  NAND2_X1 U7346 ( .A1(n6449), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6576) );
  NAND3_X1 U7347 ( .A1(n6571), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6576), .ZN(n6452) );
  OAI211_X1 U7348 ( .C1(n6453), .C2(n6452), .A(n6451), .B(n6450), .ZN(n6455)
         );
  NAND2_X1 U7349 ( .A1(n6453), .A2(n6452), .ZN(n6454) );
  NAND2_X1 U7350 ( .A1(n6455), .A2(n6454), .ZN(n6457) );
  AOI21_X1 U7351 ( .B1(n6457), .B2(n6458), .A(n6456), .ZN(n6461) );
  NOR2_X1 U7352 ( .A1(n6458), .A2(n6457), .ZN(n6460) );
  OAI22_X1 U7353 ( .A1(n6461), .A2(n6460), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n6459), .ZN(n6469) );
  OAI21_X1 U7354 ( .B1(MORE_REG_SCAN_IN), .B2(FLUSH_REG_SCAN_IN), .A(n6462), 
        .ZN(n6463) );
  NAND4_X1 U7355 ( .A1(n6466), .A2(n6465), .A3(n6464), .A4(n6463), .ZN(n6468)
         );
  AOI211_X1 U7356 ( .C1(n6470), .C2(n6469), .A(n6468), .B(n6467), .ZN(n6484)
         );
  OAI21_X1 U7357 ( .B1(n6472), .B2(n6471), .A(STATE2_REG_2__SCAN_IN), .ZN(
        n6473) );
  AOI221_X1 U7358 ( .B1(n6474), .B2(n6479), .C1(n4307), .C2(n6479), .A(n6473), 
        .ZN(n6477) );
  OAI221_X1 U7359 ( .B1(n6479), .B2(n6484), .C1(n6479), .C2(n6474), .A(n6477), 
        .ZN(n6566) );
  OAI21_X1 U7360 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4307), .A(n6566), .ZN(
        n6485) );
  AOI221_X1 U7361 ( .B1(n6476), .B2(STATE2_REG_0__SCAN_IN), .C1(n6485), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6475), .ZN(n6483) );
  NAND2_X1 U7362 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n6592), .ZN(n6480) );
  INV_X1 U7363 ( .A(n6477), .ZN(n6478) );
  OAI211_X1 U7364 ( .C1(n6481), .C2(n6480), .A(n6479), .B(n6478), .ZN(n6482)
         );
  OAI211_X1 U7365 ( .C1(n6484), .C2(n6486), .A(n6483), .B(n6482), .ZN(U3148)
         );
  NAND3_X1 U7366 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6492), .A3(n6485), .ZN(
        n6491) );
  OAI21_X1 U7367 ( .B1(READY_N), .B2(n6487), .A(n6486), .ZN(n6489) );
  AOI21_X1 U7368 ( .B1(n6489), .B2(n6566), .A(n6488), .ZN(n6490) );
  NAND2_X1 U7369 ( .A1(n6491), .A2(n6490), .ZN(U3149) );
  OAI211_X1 U7370 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n4307), .A(n6564), .B(
        n6492), .ZN(n6494) );
  OAI21_X1 U7371 ( .B1(n6592), .B2(n6494), .A(n6493), .ZN(U3150) );
  INV_X1 U7372 ( .A(n6563), .ZN(n6495) );
  AND2_X1 U7373 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6495), .ZN(U3151) );
  INV_X1 U7374 ( .A(DATAWIDTH_REG_30__SCAN_IN), .ZN(n6613) );
  NOR2_X1 U7375 ( .A1(n6563), .A2(n6613), .ZN(U3152) );
  AND2_X1 U7376 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6495), .ZN(U3153) );
  AND2_X1 U7377 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6495), .ZN(U3154) );
  AND2_X1 U7378 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6495), .ZN(U3155) );
  AND2_X1 U7379 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6495), .ZN(U3156) );
  INV_X1 U7380 ( .A(DATAWIDTH_REG_25__SCAN_IN), .ZN(n6629) );
  NOR2_X1 U7381 ( .A1(n6563), .A2(n6629), .ZN(U3157) );
  AND2_X1 U7382 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6495), .ZN(U3158) );
  AND2_X1 U7383 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6495), .ZN(U3159) );
  AND2_X1 U7384 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6495), .ZN(U3160) );
  AND2_X1 U7385 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6495), .ZN(U3161) );
  INV_X1 U7386 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6735) );
  NOR2_X1 U7387 ( .A1(n6563), .A2(n6735), .ZN(U3162) );
  AND2_X1 U7388 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6495), .ZN(U3163) );
  AND2_X1 U7389 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6495), .ZN(U3164) );
  AND2_X1 U7390 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6495), .ZN(U3165) );
  AND2_X1 U7391 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6495), .ZN(U3166) );
  AND2_X1 U7392 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6495), .ZN(U3167) );
  AND2_X1 U7393 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6495), .ZN(U3168) );
  AND2_X1 U7394 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6495), .ZN(U3169) );
  AND2_X1 U7395 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6495), .ZN(U3170) );
  AND2_X1 U7396 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6495), .ZN(U3171) );
  AND2_X1 U7397 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6495), .ZN(U3172) );
  AND2_X1 U7398 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6495), .ZN(U3173) );
  AND2_X1 U7399 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6495), .ZN(U3174) );
  INV_X1 U7400 ( .A(DATAWIDTH_REG_7__SCAN_IN), .ZN(n6751) );
  NOR2_X1 U7401 ( .A1(n6563), .A2(n6751), .ZN(U3175) );
  AND2_X1 U7402 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6495), .ZN(U3176) );
  AND2_X1 U7403 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6495), .ZN(U3177) );
  AND2_X1 U7404 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6495), .ZN(U3178) );
  AND2_X1 U7405 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6495), .ZN(U3179) );
  AND2_X1 U7406 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6495), .ZN(U3180) );
  NOR2_X1 U7407 ( .A1(n6502), .A2(n6512), .ZN(n6503) );
  AOI22_X1 U7408 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6511) );
  AND2_X1 U7409 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6499) );
  INV_X1 U7410 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6497) );
  INV_X1 U7411 ( .A(NA_N), .ZN(n6504) );
  AOI221_X1 U7412 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6504), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6508) );
  AOI221_X1 U7413 ( .B1(n6499), .B2(n6597), .C1(n6497), .C2(n6597), .A(n6508), 
        .ZN(n6496) );
  OAI21_X1 U7414 ( .B1(n6503), .B2(n6511), .A(n6496), .ZN(U3181) );
  NOR2_X1 U7415 ( .A1(n6506), .A2(n6497), .ZN(n6505) );
  NAND2_X1 U7416 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6498) );
  OAI21_X1 U7417 ( .B1(n6505), .B2(n6499), .A(n6498), .ZN(n6500) );
  OAI211_X1 U7418 ( .C1(n6502), .C2(n4307), .A(n6501), .B(n6500), .ZN(U3182)
         );
  AOI21_X1 U7419 ( .B1(n6505), .B2(n6504), .A(n6503), .ZN(n6510) );
  AOI221_X1 U7420 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n4307), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6507) );
  AOI221_X1 U7421 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6507), .C2(HOLD), .A(n6506), .ZN(n6509) );
  OAI22_X1 U7422 ( .A1(n6511), .A2(n6510), .B1(n6509), .B2(n6508), .ZN(U3183)
         );
  NAND2_X1 U7423 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6559), .ZN(n6556) );
  NAND2_X1 U7424 ( .A1(n6512), .A2(n6559), .ZN(n6546) );
  INV_X1 U7425 ( .A(n6546), .ZN(n6785) );
  AOI22_X1 U7426 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6597), .ZN(n6513) );
  OAI21_X1 U7427 ( .B1(n5251), .B2(n6556), .A(n6513), .ZN(U3184) );
  AOI22_X1 U7428 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6597), .ZN(n6514) );
  OAI21_X1 U7429 ( .B1(n4415), .B2(n6556), .A(n6514), .ZN(U3185) );
  INV_X1 U7430 ( .A(n6556), .ZN(n6786) );
  AOI22_X1 U7431 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6786), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6597), .ZN(n6515) );
  OAI21_X1 U7432 ( .B1(n6517), .B2(n6546), .A(n6515), .ZN(U3186) );
  AOI22_X1 U7433 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6597), .ZN(n6516) );
  OAI21_X1 U7434 ( .B1(n6517), .B2(n6556), .A(n6516), .ZN(U3187) );
  INV_X1 U7435 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6744) );
  AOI22_X1 U7436 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6597), .ZN(n6518) );
  OAI21_X1 U7437 ( .B1(n6744), .B2(n6556), .A(n6518), .ZN(U3188) );
  AOI22_X1 U7438 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6786), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6597), .ZN(n6519) );
  OAI21_X1 U7439 ( .B1(n6521), .B2(n6546), .A(n6519), .ZN(U3189) );
  INV_X1 U7440 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6610) );
  INV_X1 U7441 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6520) );
  OAI222_X1 U7442 ( .A1(n6556), .A2(n6521), .B1(n6610), .B2(n6559), .C1(n6520), 
        .C2(n6546), .ZN(U3190) );
  AOI22_X1 U7443 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6786), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6597), .ZN(n6522) );
  OAI21_X1 U7444 ( .B1(n6722), .B2(n6546), .A(n6522), .ZN(U3191) );
  AOI22_X1 U7445 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6786), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6597), .ZN(n6523) );
  OAI21_X1 U7446 ( .B1(n6525), .B2(n6546), .A(n6523), .ZN(U3192) );
  AOI22_X1 U7447 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6597), .ZN(n6524) );
  OAI21_X1 U7448 ( .B1(n6525), .B2(n6556), .A(n6524), .ZN(U3193) );
  AOI22_X1 U7449 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6786), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6597), .ZN(n6526) );
  OAI21_X1 U7450 ( .B1(n6528), .B2(n6546), .A(n6526), .ZN(U3194) );
  AOI22_X1 U7451 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6597), .ZN(n6527) );
  OAI21_X1 U7452 ( .B1(n6528), .B2(n6556), .A(n6527), .ZN(U3195) );
  AOI22_X1 U7453 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6786), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6597), .ZN(n6529) );
  OAI21_X1 U7454 ( .B1(n5396), .B2(n6546), .A(n6529), .ZN(U3196) );
  AOI22_X1 U7455 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6597), .ZN(n6530) );
  OAI21_X1 U7456 ( .B1(n5396), .B2(n6556), .A(n6530), .ZN(U3197) );
  AOI22_X1 U7457 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6597), .ZN(n6531) );
  OAI21_X1 U7458 ( .B1(n6532), .B2(n6556), .A(n6531), .ZN(U3198) );
  AOI22_X1 U7459 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6786), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6597), .ZN(n6533) );
  OAI21_X1 U7460 ( .B1(n5732), .B2(n6546), .A(n6533), .ZN(U3199) );
  AOI22_X1 U7461 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6786), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6597), .ZN(n6534) );
  OAI21_X1 U7462 ( .B1(n6535), .B2(n6546), .A(n6534), .ZN(U3200) );
  AOI222_X1 U7463 ( .A1(n6785), .A2(REIP_REG_19__SCAN_IN), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6597), .C1(REIP_REG_18__SCAN_IN), .C2(
        n6786), .ZN(n6536) );
  INV_X1 U7464 ( .A(n6536), .ZN(U3201) );
  AOI22_X1 U7465 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6597), .ZN(n6537) );
  OAI21_X1 U7466 ( .B1(n6538), .B2(n6556), .A(n6537), .ZN(U3202) );
  AOI22_X1 U7467 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6597), .ZN(n6539) );
  OAI21_X1 U7468 ( .B1(n6540), .B2(n6556), .A(n6539), .ZN(U3204) );
  INV_X1 U7469 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6741) );
  INV_X1 U7470 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6543) );
  OAI222_X1 U7471 ( .A1(n6556), .A2(n6541), .B1(n6741), .B2(n6559), .C1(n6543), 
        .C2(n6546), .ZN(U3205) );
  AOI22_X1 U7472 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6597), .ZN(n6542) );
  OAI21_X1 U7473 ( .B1(n6543), .B2(n6556), .A(n6542), .ZN(U3206) );
  INV_X1 U7474 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6599) );
  AOI22_X1 U7475 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6597), .ZN(n6544) );
  OAI21_X1 U7476 ( .B1(n6599), .B2(n6556), .A(n6544), .ZN(U3207) );
  INV_X1 U7477 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6548) );
  AOI22_X1 U7478 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6786), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6597), .ZN(n6545) );
  OAI21_X1 U7479 ( .B1(n6548), .B2(n6546), .A(n6545), .ZN(U3208) );
  AOI22_X1 U7480 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6597), .ZN(n6547) );
  OAI21_X1 U7481 ( .B1(n6548), .B2(n6556), .A(n6547), .ZN(U3209) );
  AOI22_X1 U7482 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6597), .ZN(n6549) );
  OAI21_X1 U7483 ( .B1(n6550), .B2(n6556), .A(n6549), .ZN(U3210) );
  AOI22_X1 U7484 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6597), .ZN(n6551) );
  OAI21_X1 U7485 ( .B1(n6552), .B2(n6556), .A(n6551), .ZN(U3211) );
  AOI22_X1 U7486 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6597), .ZN(n6553) );
  OAI21_X1 U7487 ( .B1(n6554), .B2(n6556), .A(n6553), .ZN(U3212) );
  AOI22_X1 U7488 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6785), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6597), .ZN(n6555) );
  OAI21_X1 U7489 ( .B1(n6557), .B2(n6556), .A(n6555), .ZN(U3213) );
  INV_X1 U7490 ( .A(BE_N_REG_3__SCAN_IN), .ZN(n6621) );
  AOI22_X1 U7491 ( .A1(n6559), .A2(n6558), .B1(n6621), .B2(n6597), .ZN(U3445)
         );
  MUX2_X1 U7492 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6597), .Z(U3446) );
  MUX2_X1 U7493 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6597), .Z(U3447) );
  MUX2_X1 U7494 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6597), .Z(U3448) );
  OAI21_X1 U7495 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6563), .A(n6561), .ZN(
        n6560) );
  INV_X1 U7496 ( .A(n6560), .ZN(U3451) );
  OAI21_X1 U7497 ( .B1(n6563), .B2(n6562), .A(n6561), .ZN(U3452) );
  OAI211_X1 U7498 ( .C1(n6567), .C2(n6566), .A(n6565), .B(n6564), .ZN(U3453)
         );
  AOI21_X1 U7499 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n6569), .A(n6568), .ZN(
        n6570) );
  OAI211_X1 U7500 ( .C1(n6571), .C2(n6575), .A(n6573), .B(n6570), .ZN(n6572)
         );
  OAI21_X1 U7501 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6573), .A(n6572), 
        .ZN(n6574) );
  OAI21_X1 U7502 ( .B1(n6576), .B2(n6575), .A(n6574), .ZN(U3461) );
  AOI21_X1 U7503 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6577) );
  AOI22_X1 U7504 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6577), .B2(n5251), .ZN(n6579) );
  INV_X1 U7505 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6578) );
  AOI22_X1 U7506 ( .A1(n6580), .A2(n6579), .B1(n6578), .B2(n6583), .ZN(U3468)
         );
  INV_X1 U7507 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6584) );
  NOR2_X1 U7508 ( .A1(n6583), .A2(REIP_REG_1__SCAN_IN), .ZN(n6581) );
  AOI22_X1 U7509 ( .A1(n6584), .A2(n6583), .B1(n6582), .B2(n6581), .ZN(U3469)
         );
  NAND2_X1 U7510 ( .A1(n6597), .A2(W_R_N_REG_SCAN_IN), .ZN(n6585) );
  OAI21_X1 U7511 ( .B1(n6597), .B2(READREQUEST_REG_SCAN_IN), .A(n6585), .ZN(
        U3470) );
  AOI211_X1 U7512 ( .C1(n6588), .C2(n4307), .A(n6587), .B(n6586), .ZN(n6596)
         );
  INV_X1 U7513 ( .A(n6589), .ZN(n6590) );
  OAI211_X1 U7514 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6591), .A(n6590), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6593) );
  AOI21_X1 U7515 ( .B1(n6593), .B2(STATE2_REG_0__SCAN_IN), .A(n6592), .ZN(
        n6595) );
  NAND2_X1 U7516 ( .A1(n6596), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6594) );
  OAI21_X1 U7517 ( .B1(n6596), .B2(n6595), .A(n6594), .ZN(U3472) );
  MUX2_X1 U7518 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6597), .Z(U3473) );
  AOI22_X1 U7519 ( .A1(n6772), .A2(keyinput78), .B1(keyinput113), .B2(n6599), 
        .ZN(n6598) );
  OAI221_X1 U7520 ( .B1(n6772), .B2(keyinput78), .C1(n6599), .C2(keyinput113), 
        .A(n6598), .ZN(n6607) );
  AOI22_X1 U7521 ( .A1(n6709), .A2(keyinput84), .B1(n6759), .B2(keyinput114), 
        .ZN(n6600) );
  OAI221_X1 U7522 ( .B1(n6709), .B2(keyinput84), .C1(n6759), .C2(keyinput114), 
        .A(n6600), .ZN(n6606) );
  AOI22_X1 U7523 ( .A1(n6602), .A2(keyinput65), .B1(n6760), .B2(keyinput117), 
        .ZN(n6601) );
  OAI221_X1 U7524 ( .B1(n6602), .B2(keyinput65), .C1(n6760), .C2(keyinput117), 
        .A(n6601), .ZN(n6605) );
  AOI22_X1 U7525 ( .A1(n5732), .A2(keyinput115), .B1(n6707), .B2(keyinput87), 
        .ZN(n6603) );
  OAI221_X1 U7526 ( .B1(n5732), .B2(keyinput115), .C1(n6707), .C2(keyinput87), 
        .A(n6603), .ZN(n6604) );
  NOR4_X1 U7527 ( .A1(n6607), .A2(n6606), .A3(n6605), .A4(n6604), .ZN(n6641)
         );
  AOI22_X1 U7528 ( .A1(n6751), .A2(keyinput74), .B1(n6757), .B2(keyinput68), 
        .ZN(n6608) );
  OAI221_X1 U7529 ( .B1(n6751), .B2(keyinput74), .C1(n6757), .C2(keyinput68), 
        .A(n6608), .ZN(n6617) );
  AOI22_X1 U7530 ( .A1(n6610), .A2(keyinput106), .B1(n5513), .B2(keyinput69), 
        .ZN(n6609) );
  OAI221_X1 U7531 ( .B1(n6610), .B2(keyinput106), .C1(n5513), .C2(keyinput69), 
        .A(n6609), .ZN(n6616) );
  AOI22_X1 U7532 ( .A1(n6722), .A2(keyinput76), .B1(n6710), .B2(keyinput96), 
        .ZN(n6611) );
  OAI221_X1 U7533 ( .B1(n6722), .B2(keyinput76), .C1(n6710), .C2(keyinput96), 
        .A(n6611), .ZN(n6615) );
  AOI22_X1 U7534 ( .A1(n6613), .A2(keyinput111), .B1(n6738), .B2(keyinput116), 
        .ZN(n6612) );
  OAI221_X1 U7535 ( .B1(n6613), .B2(keyinput111), .C1(n6738), .C2(keyinput116), 
        .A(n6612), .ZN(n6614) );
  NOR4_X1 U7536 ( .A1(n6617), .A2(n6616), .A3(n6615), .A4(n6614), .ZN(n6640)
         );
  INV_X1 U7537 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n6619) );
  AOI22_X1 U7538 ( .A1(n6619), .A2(keyinput121), .B1(n6756), .B2(keyinput103), 
        .ZN(n6618) );
  OAI221_X1 U7539 ( .B1(n6619), .B2(keyinput121), .C1(n6756), .C2(keyinput103), 
        .A(n6618), .ZN(n6627) );
  AOI22_X1 U7540 ( .A1(n5396), .A2(keyinput67), .B1(keyinput81), .B2(n6621), 
        .ZN(n6620) );
  OAI221_X1 U7541 ( .B1(n5396), .B2(keyinput67), .C1(n6621), .C2(keyinput81), 
        .A(n6620), .ZN(n6626) );
  INV_X1 U7542 ( .A(DATAI_14_), .ZN(n6765) );
  INV_X1 U7543 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n6770) );
  AOI22_X1 U7544 ( .A1(n6765), .A2(keyinput102), .B1(keyinput123), .B2(n6770), 
        .ZN(n6622) );
  OAI221_X1 U7545 ( .B1(n6765), .B2(keyinput102), .C1(n6770), .C2(keyinput123), 
        .A(n6622), .ZN(n6625) );
  INV_X1 U7546 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n6740) );
  AOI22_X1 U7547 ( .A1(n6740), .A2(keyinput95), .B1(keyinput97), .B2(n4091), 
        .ZN(n6623) );
  OAI221_X1 U7548 ( .B1(n6740), .B2(keyinput95), .C1(n4091), .C2(keyinput97), 
        .A(n6623), .ZN(n6624) );
  NOR4_X1 U7549 ( .A1(n6627), .A2(n6626), .A3(n6625), .A4(n6624), .ZN(n6639)
         );
  INV_X1 U7550 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n6726) );
  AOI22_X1 U7551 ( .A1(n6726), .A2(keyinput92), .B1(keyinput107), .B2(n6629), 
        .ZN(n6628) );
  OAI221_X1 U7552 ( .B1(n6726), .B2(keyinput92), .C1(n6629), .C2(keyinput107), 
        .A(n6628), .ZN(n6637) );
  AOI22_X1 U7553 ( .A1(n4507), .A2(keyinput99), .B1(n6631), .B2(keyinput119), 
        .ZN(n6630) );
  OAI221_X1 U7554 ( .B1(n4507), .B2(keyinput99), .C1(n6631), .C2(keyinput119), 
        .A(n6630), .ZN(n6636) );
  INV_X1 U7555 ( .A(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n6723) );
  INV_X1 U7556 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n6706) );
  AOI22_X1 U7557 ( .A1(n6723), .A2(keyinput109), .B1(n6706), .B2(keyinput105), 
        .ZN(n6632) );
  OAI221_X1 U7558 ( .B1(n6723), .B2(keyinput109), .C1(n6706), .C2(keyinput105), 
        .A(n6632), .ZN(n6635) );
  AOI22_X1 U7559 ( .A1(n6766), .A2(keyinput66), .B1(keyinput88), .B2(n6735), 
        .ZN(n6633) );
  OAI221_X1 U7560 ( .B1(n6766), .B2(keyinput66), .C1(n6735), .C2(keyinput88), 
        .A(n6633), .ZN(n6634) );
  NOR4_X1 U7561 ( .A1(n6637), .A2(n6636), .A3(n6635), .A4(n6634), .ZN(n6638)
         );
  AND4_X1 U7562 ( .A1(n6641), .A2(n6640), .A3(n6639), .A4(n6638), .ZN(n6784)
         );
  OAI22_X1 U7563 ( .A1(INSTQUEUE_REG_12__3__SCAN_IN), .A2(keyinput75), .B1(
        keyinput73), .B2(STATE_REG_2__SCAN_IN), .ZN(n6642) );
  AOI221_X1 U7564 ( .B1(INSTQUEUE_REG_12__3__SCAN_IN), .B2(keyinput75), .C1(
        STATE_REG_2__SCAN_IN), .C2(keyinput73), .A(n6642), .ZN(n6649) );
  OAI22_X1 U7565 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(keyinput98), .B1(
        keyinput89), .B2(DATAI_18_), .ZN(n6643) );
  AOI221_X1 U7566 ( .B1(INSTQUEUE_REG_12__6__SCAN_IN), .B2(keyinput98), .C1(
        DATAI_18_), .C2(keyinput89), .A(n6643), .ZN(n6648) );
  OAI22_X1 U7567 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(keyinput71), .B1(
        EBX_REG_31__SCAN_IN), .B2(keyinput90), .ZN(n6644) );
  AOI221_X1 U7568 ( .B1(INSTQUEUE_REG_5__4__SCAN_IN), .B2(keyinput71), .C1(
        keyinput90), .C2(EBX_REG_31__SCAN_IN), .A(n6644), .ZN(n6647) );
  OAI22_X1 U7569 ( .A1(EBX_REG_15__SCAN_IN), .A2(keyinput100), .B1(keyinput94), 
        .B2(DATAO_REG_31__SCAN_IN), .ZN(n6645) );
  AOI221_X1 U7570 ( .B1(EBX_REG_15__SCAN_IN), .B2(keyinput100), .C1(
        DATAO_REG_31__SCAN_IN), .C2(keyinput94), .A(n6645), .ZN(n6646) );
  NAND4_X1 U7571 ( .A1(n6649), .A2(n6648), .A3(n6647), .A4(n6646), .ZN(n6678)
         );
  OAI22_X1 U7572 ( .A1(INSTQUEUE_REG_2__2__SCAN_IN), .A2(keyinput118), .B1(
        keyinput64), .B2(HOLD), .ZN(n6650) );
  AOI221_X1 U7573 ( .B1(INSTQUEUE_REG_2__2__SCAN_IN), .B2(keyinput118), .C1(
        HOLD), .C2(keyinput64), .A(n6650), .ZN(n6657) );
  OAI22_X1 U7574 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(keyinput77), .B1(
        DATAO_REG_8__SCAN_IN), .B2(keyinput85), .ZN(n6651) );
  AOI221_X1 U7575 ( .B1(INSTQUEUE_REG_5__1__SCAN_IN), .B2(keyinput77), .C1(
        keyinput85), .C2(DATAO_REG_8__SCAN_IN), .A(n6651), .ZN(n6656) );
  OAI22_X1 U7576 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(keyinput122), .B1(
        REIP_REG_5__SCAN_IN), .B2(keyinput112), .ZN(n6652) );
  AOI221_X1 U7577 ( .B1(INSTQUEUE_REG_6__7__SCAN_IN), .B2(keyinput122), .C1(
        keyinput112), .C2(REIP_REG_5__SCAN_IN), .A(n6652), .ZN(n6655) );
  OAI22_X1 U7578 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(keyinput93), .B1(
        keyinput124), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6653) );
  AOI221_X1 U7579 ( .B1(INSTQUEUE_REG_9__4__SCAN_IN), .B2(keyinput93), .C1(
        PHYADDRPOINTER_REG_7__SCAN_IN), .C2(keyinput124), .A(n6653), .ZN(n6654) );
  NAND4_X1 U7580 ( .A1(n6657), .A2(n6656), .A3(n6655), .A4(n6654), .ZN(n6677)
         );
  OAI22_X1 U7581 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(keyinput86), .B1(
        DATAO_REG_7__SCAN_IN), .B2(keyinput70), .ZN(n6658) );
  AOI221_X1 U7582 ( .B1(INSTQUEUE_REG_4__4__SCAN_IN), .B2(keyinput86), .C1(
        keyinput70), .C2(DATAO_REG_7__SCAN_IN), .A(n6658), .ZN(n6666) );
  OAI22_X1 U7583 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(keyinput104), 
        .B1(keyinput83), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6659) );
  AOI221_X1 U7584 ( .B1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(keyinput104), 
        .C1(INSTADDRPOINTER_REG_27__SCAN_IN), .C2(keyinput83), .A(n6659), .ZN(
        n6665) );
  INV_X1 U7585 ( .A(DATAI_12_), .ZN(n6661) );
  OAI22_X1 U7586 ( .A1(n6661), .A2(keyinput80), .B1(keyinput120), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n6660) );
  AOI221_X1 U7587 ( .B1(n6661), .B2(keyinput80), .C1(UWORD_REG_11__SCAN_IN), 
        .C2(keyinput120), .A(n6660), .ZN(n6664) );
  OAI22_X1 U7588 ( .A1(n6741), .A2(keyinput72), .B1(LWORD_REG_7__SCAN_IN), 
        .B2(keyinput101), .ZN(n6662) );
  AOI221_X1 U7589 ( .B1(n6741), .B2(keyinput72), .C1(keyinput101), .C2(
        LWORD_REG_7__SCAN_IN), .A(n6662), .ZN(n6663) );
  NAND4_X1 U7590 ( .A1(n6666), .A2(n6665), .A3(n6664), .A4(n6663), .ZN(n6676)
         );
  OAI22_X1 U7591 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(keyinput127), 
        .B1(keyinput110), .B2(LWORD_REG_10__SCAN_IN), .ZN(n6667) );
  AOI221_X1 U7592 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(keyinput127), 
        .C1(LWORD_REG_10__SCAN_IN), .C2(keyinput110), .A(n6667), .ZN(n6674) );
  OAI22_X1 U7593 ( .A1(INSTQUEUE_REG_8__2__SCAN_IN), .A2(keyinput125), .B1(
        keyinput82), .B2(DATAO_REG_24__SCAN_IN), .ZN(n6668) );
  AOI221_X1 U7594 ( .B1(INSTQUEUE_REG_8__2__SCAN_IN), .B2(keyinput125), .C1(
        DATAO_REG_24__SCAN_IN), .C2(keyinput82), .A(n6668), .ZN(n6673) );
  OAI22_X1 U7595 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(keyinput91), .B1(
        DATAO_REG_20__SCAN_IN), .B2(keyinput126), .ZN(n6669) );
  AOI221_X1 U7596 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(keyinput91), 
        .C1(keyinput126), .C2(DATAO_REG_20__SCAN_IN), .A(n6669), .ZN(n6672) );
  OAI22_X1 U7597 ( .A1(DATAI_17_), .A2(keyinput79), .B1(keyinput108), .B2(
        ADDRESS_REG_17__SCAN_IN), .ZN(n6670) );
  AOI221_X1 U7598 ( .B1(DATAI_17_), .B2(keyinput79), .C1(
        ADDRESS_REG_17__SCAN_IN), .C2(keyinput108), .A(n6670), .ZN(n6671) );
  NAND4_X1 U7599 ( .A1(n6674), .A2(n6673), .A3(n6672), .A4(n6671), .ZN(n6675)
         );
  NOR4_X1 U7600 ( .A1(n6678), .A2(n6677), .A3(n6676), .A4(n6675), .ZN(n6783)
         );
  AOI22_X1 U7601 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(keyinput47), .B1(
        DATAI_17_), .B2(keyinput15), .ZN(n6679) );
  OAI221_X1 U7602 ( .B1(DATAWIDTH_REG_30__SCAN_IN), .B2(keyinput47), .C1(
        DATAI_17_), .C2(keyinput15), .A(n6679), .ZN(n6686) );
  AOI22_X1 U7603 ( .A1(LWORD_REG_10__SCAN_IN), .A2(keyinput46), .B1(
        STATE_REG_2__SCAN_IN), .B2(keyinput9), .ZN(n6680) );
  OAI221_X1 U7604 ( .B1(LWORD_REG_10__SCAN_IN), .B2(keyinput46), .C1(
        STATE_REG_2__SCAN_IN), .C2(keyinput9), .A(n6680), .ZN(n6685) );
  AOI22_X1 U7605 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(keyinput63), .B1(
        INSTQUEUE_REG_5__4__SCAN_IN), .B2(keyinput7), .ZN(n6681) );
  OAI221_X1 U7606 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(keyinput63), 
        .C1(INSTQUEUE_REG_5__4__SCAN_IN), .C2(keyinput7), .A(n6681), .ZN(n6684) );
  AOI22_X1 U7607 ( .A1(REIP_REG_24__SCAN_IN), .A2(keyinput49), .B1(
        INSTADDRPOINTER_REG_27__SCAN_IN), .B2(keyinput19), .ZN(n6682) );
  OAI221_X1 U7608 ( .B1(REIP_REG_24__SCAN_IN), .B2(keyinput49), .C1(
        INSTADDRPOINTER_REG_27__SCAN_IN), .C2(keyinput19), .A(n6682), .ZN(
        n6683) );
  NOR4_X1 U7609 ( .A1(n6686), .A2(n6685), .A3(n6684), .A4(n6683), .ZN(n6718)
         );
  AOI22_X1 U7610 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(keyinput27), .B1(
        INSTQUEUE_REG_2__2__SCAN_IN), .B2(keyinput54), .ZN(n6687) );
  OAI221_X1 U7611 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(keyinput27), 
        .C1(INSTQUEUE_REG_2__2__SCAN_IN), .C2(keyinput54), .A(n6687), .ZN(
        n6694) );
  AOI22_X1 U7612 ( .A1(DATAO_REG_24__SCAN_IN), .A2(keyinput18), .B1(DATAI_12_), 
        .B2(keyinput16), .ZN(n6688) );
  OAI221_X1 U7613 ( .B1(DATAO_REG_24__SCAN_IN), .B2(keyinput18), .C1(DATAI_12_), .C2(keyinput16), .A(n6688), .ZN(n6693) );
  AOI22_X1 U7614 ( .A1(EBX_REG_31__SCAN_IN), .A2(keyinput26), .B1(
        INSTQUEUE_REG_6__7__SCAN_IN), .B2(keyinput58), .ZN(n6689) );
  OAI221_X1 U7615 ( .B1(EBX_REG_31__SCAN_IN), .B2(keyinput26), .C1(
        INSTQUEUE_REG_6__7__SCAN_IN), .C2(keyinput58), .A(n6689), .ZN(n6692)
         );
  AOI22_X1 U7616 ( .A1(ADDRESS_REG_6__SCAN_IN), .A2(keyinput42), .B1(
        INSTQUEUE_REG_12__2__SCAN_IN), .B2(keyinput55), .ZN(n6690) );
  OAI221_X1 U7617 ( .B1(ADDRESS_REG_6__SCAN_IN), .B2(keyinput42), .C1(
        INSTQUEUE_REG_12__2__SCAN_IN), .C2(keyinput55), .A(n6690), .ZN(n6691)
         );
  NOR4_X1 U7618 ( .A1(n6694), .A2(n6693), .A3(n6692), .A4(n6691), .ZN(n6717)
         );
  AOI22_X1 U7619 ( .A1(DATAI_29_), .A2(keyinput1), .B1(
        INSTQUEUE_REG_12__3__SCAN_IN), .B2(keyinput11), .ZN(n6695) );
  OAI221_X1 U7620 ( .B1(DATAI_29_), .B2(keyinput1), .C1(
        INSTQUEUE_REG_12__3__SCAN_IN), .C2(keyinput11), .A(n6695), .ZN(n6702)
         );
  AOI22_X1 U7621 ( .A1(HOLD), .A2(keyinput0), .B1(EAX_REG_22__SCAN_IN), .B2(
        keyinput33), .ZN(n6696) );
  OAI221_X1 U7622 ( .B1(HOLD), .B2(keyinput0), .C1(EAX_REG_22__SCAN_IN), .C2(
        keyinput33), .A(n6696), .ZN(n6701) );
  AOI22_X1 U7623 ( .A1(ADDRESS_REG_17__SCAN_IN), .A2(keyinput44), .B1(
        DATAO_REG_20__SCAN_IN), .B2(keyinput62), .ZN(n6697) );
  OAI221_X1 U7624 ( .B1(ADDRESS_REG_17__SCAN_IN), .B2(keyinput44), .C1(
        DATAO_REG_20__SCAN_IN), .C2(keyinput62), .A(n6697), .ZN(n6700) );
  AOI22_X1 U7625 ( .A1(BE_N_REG_3__SCAN_IN), .A2(keyinput17), .B1(
        DATAO_REG_25__SCAN_IN), .B2(keyinput57), .ZN(n6698) );
  OAI221_X1 U7626 ( .B1(BE_N_REG_3__SCAN_IN), .B2(keyinput17), .C1(
        DATAO_REG_25__SCAN_IN), .C2(keyinput57), .A(n6698), .ZN(n6699) );
  NOR4_X1 U7627 ( .A1(n6702), .A2(n6701), .A3(n6700), .A4(n6699), .ZN(n6716)
         );
  AOI22_X1 U7628 ( .A1(DATAO_REG_7__SCAN_IN), .A2(keyinput6), .B1(
        INSTQUEUE_REG_4__4__SCAN_IN), .B2(keyinput22), .ZN(n6703) );
  OAI221_X1 U7629 ( .B1(DATAO_REG_7__SCAN_IN), .B2(keyinput6), .C1(
        INSTQUEUE_REG_4__4__SCAN_IN), .C2(keyinput22), .A(n6703), .ZN(n6714)
         );
  AOI22_X1 U7630 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(keyinput43), .B1(
        INSTQUEUE_REG_9__4__SCAN_IN), .B2(keyinput29), .ZN(n6704) );
  OAI221_X1 U7631 ( .B1(DATAWIDTH_REG_25__SCAN_IN), .B2(keyinput43), .C1(
        INSTQUEUE_REG_9__4__SCAN_IN), .C2(keyinput29), .A(n6704), .ZN(n6713)
         );
  AOI22_X1 U7632 ( .A1(n6707), .A2(keyinput23), .B1(n6706), .B2(keyinput41), 
        .ZN(n6705) );
  OAI221_X1 U7633 ( .B1(n6707), .B2(keyinput23), .C1(n6706), .C2(keyinput41), 
        .A(n6705), .ZN(n6712) );
  AOI22_X1 U7634 ( .A1(n6710), .A2(keyinput32), .B1(n6709), .B2(keyinput20), 
        .ZN(n6708) );
  OAI221_X1 U7635 ( .B1(n6710), .B2(keyinput32), .C1(n6709), .C2(keyinput20), 
        .A(n6708), .ZN(n6711) );
  NOR4_X1 U7636 ( .A1(n6714), .A2(n6713), .A3(n6712), .A4(n6711), .ZN(n6715)
         );
  NAND4_X1 U7637 ( .A1(n6718), .A2(n6717), .A3(n6716), .A4(n6715), .ZN(n6782)
         );
  INV_X1 U7638 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6720) );
  AOI22_X1 U7639 ( .A1(n6720), .A2(keyinput13), .B1(keyinput51), .B2(n5732), 
        .ZN(n6719) );
  OAI221_X1 U7640 ( .B1(n6720), .B2(keyinput13), .C1(n5732), .C2(keyinput51), 
        .A(n6719), .ZN(n6732) );
  AOI22_X1 U7641 ( .A1(n6723), .A2(keyinput45), .B1(keyinput12), .B2(n6722), 
        .ZN(n6721) );
  OAI221_X1 U7642 ( .B1(n6723), .B2(keyinput45), .C1(n6722), .C2(keyinput12), 
        .A(n6721), .ZN(n6731) );
  INV_X1 U7643 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n6725) );
  AOI22_X1 U7644 ( .A1(n6725), .A2(keyinput37), .B1(n5513), .B2(keyinput5), 
        .ZN(n6724) );
  OAI221_X1 U7645 ( .B1(n6725), .B2(keyinput37), .C1(n5513), .C2(keyinput5), 
        .A(n6724), .ZN(n6730) );
  XOR2_X1 U7646 ( .A(n6726), .B(keyinput28), .Z(n6728) );
  XNOR2_X1 U7647 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(keyinput40), .ZN(
        n6727) );
  NAND2_X1 U7648 ( .A1(n6728), .A2(n6727), .ZN(n6729) );
  NOR4_X1 U7649 ( .A1(n6732), .A2(n6731), .A3(n6730), .A4(n6729), .ZN(n6780)
         );
  INV_X1 U7650 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n6734) );
  AOI22_X1 U7651 ( .A1(n6735), .A2(keyinput24), .B1(n6734), .B2(keyinput30), 
        .ZN(n6733) );
  OAI221_X1 U7652 ( .B1(n6735), .B2(keyinput24), .C1(n6734), .C2(keyinput30), 
        .A(n6733), .ZN(n6748) );
  AOI22_X1 U7653 ( .A1(n6738), .A2(keyinput52), .B1(keyinput60), .B2(n6737), 
        .ZN(n6736) );
  OAI221_X1 U7654 ( .B1(n6738), .B2(keyinput52), .C1(n6737), .C2(keyinput60), 
        .A(n6736), .ZN(n6747) );
  AOI22_X1 U7655 ( .A1(n6741), .A2(keyinput8), .B1(n6740), .B2(keyinput31), 
        .ZN(n6739) );
  OAI221_X1 U7656 ( .B1(n6741), .B2(keyinput8), .C1(n6740), .C2(keyinput31), 
        .A(n6739), .ZN(n6746) );
  INV_X1 U7657 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n6743) );
  AOI22_X1 U7658 ( .A1(n6744), .A2(keyinput48), .B1(keyinput56), .B2(n6743), 
        .ZN(n6742) );
  OAI221_X1 U7659 ( .B1(n6744), .B2(keyinput48), .C1(n6743), .C2(keyinput56), 
        .A(n6742), .ZN(n6745) );
  NOR4_X1 U7660 ( .A1(n6748), .A2(n6747), .A3(n6746), .A4(n6745), .ZN(n6779)
         );
  INV_X1 U7661 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n6750) );
  AOI22_X1 U7662 ( .A1(n6750), .A2(keyinput21), .B1(n4871), .B2(keyinput61), 
        .ZN(n6749) );
  OAI221_X1 U7663 ( .B1(n6750), .B2(keyinput21), .C1(n4871), .C2(keyinput61), 
        .A(n6749), .ZN(n6754) );
  XOR2_X1 U7664 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .B(keyinput34), .Z(n6753)
         );
  XNOR2_X1 U7665 ( .A(n6751), .B(keyinput10), .ZN(n6752) );
  OR3_X1 U7666 ( .A1(n6754), .A2(n6753), .A3(n6752), .ZN(n6763) );
  AOI22_X1 U7667 ( .A1(n6757), .A2(keyinput4), .B1(keyinput39), .B2(n6756), 
        .ZN(n6755) );
  OAI221_X1 U7668 ( .B1(n6757), .B2(keyinput4), .C1(n6756), .C2(keyinput39), 
        .A(n6755), .ZN(n6762) );
  AOI22_X1 U7669 ( .A1(n6760), .A2(keyinput53), .B1(n6759), .B2(keyinput50), 
        .ZN(n6758) );
  OAI221_X1 U7670 ( .B1(n6760), .B2(keyinput53), .C1(n6759), .C2(keyinput50), 
        .A(n6758), .ZN(n6761) );
  NOR3_X1 U7671 ( .A1(n6763), .A2(n6762), .A3(n6761), .ZN(n6778) );
  AOI22_X1 U7672 ( .A1(n6766), .A2(keyinput2), .B1(n6765), .B2(keyinput38), 
        .ZN(n6764) );
  OAI221_X1 U7673 ( .B1(n6766), .B2(keyinput2), .C1(n6765), .C2(keyinput38), 
        .A(n6764), .ZN(n6776) );
  INV_X1 U7674 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6768) );
  AOI22_X1 U7675 ( .A1(n5396), .A2(keyinput3), .B1(n6768), .B2(keyinput36), 
        .ZN(n6767) );
  OAI221_X1 U7676 ( .B1(n5396), .B2(keyinput3), .C1(n6768), .C2(keyinput36), 
        .A(n6767), .ZN(n6775) );
  AOI22_X1 U7677 ( .A1(n6770), .A2(keyinput59), .B1(n4512), .B2(keyinput25), 
        .ZN(n6769) );
  OAI221_X1 U7678 ( .B1(n6770), .B2(keyinput59), .C1(n4512), .C2(keyinput25), 
        .A(n6769), .ZN(n6774) );
  AOI22_X1 U7679 ( .A1(n4507), .A2(keyinput35), .B1(n6772), .B2(keyinput14), 
        .ZN(n6771) );
  OAI221_X1 U7680 ( .B1(n4507), .B2(keyinput35), .C1(n6772), .C2(keyinput14), 
        .A(n6771), .ZN(n6773) );
  NOR4_X1 U7681 ( .A1(n6776), .A2(n6775), .A3(n6774), .A4(n6773), .ZN(n6777)
         );
  NAND4_X1 U7682 ( .A1(n6780), .A2(n6779), .A3(n6778), .A4(n6777), .ZN(n6781)
         );
  AOI211_X1 U7683 ( .C1(n6784), .C2(n6783), .A(n6782), .B(n6781), .ZN(n6788)
         );
  AOI222_X1 U7684 ( .A1(n6597), .A2(ADDRESS_REG_19__SCAN_IN), .B1(
        REIP_REG_20__SCAN_IN), .B2(n6786), .C1(REIP_REG_21__SCAN_IN), .C2(
        n6785), .ZN(n6787) );
  XNOR2_X1 U7685 ( .A(n6788), .B(n6787), .ZN(U3203) );
  CLKBUF_X1 U3449 ( .A(n2996), .Z(n4199) );
  BUF_X1 U3454 ( .A(n3304), .Z(n3026) );
  CLKBUF_X1 U34590 ( .A(n3331), .Z(n3305) );
  CLKBUF_X1 U34640 ( .A(n3221), .Z(n4429) );
  CLKBUF_X1 U34710 ( .A(n3818), .Z(n3036) );
  CLKBUF_X1 U3488 ( .A(n3216), .Z(n4535) );
  CLKBUF_X1 U3499 ( .A(n6239), .Z(n6588) );
endmodule

