

module b15_C_AntiSAT_k_128_5 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696,
         n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706,
         n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726,
         n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736,
         n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
         n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766,
         n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776,
         n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786,
         n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796,
         n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806,
         n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816,
         n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826,
         n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836,
         n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846,
         n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856,
         n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
         n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
         n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
         n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
         n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
         n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
         n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
         n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
         n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
         n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
         n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
         n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
         n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
         n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
         n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006,
         n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016,
         n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026,
         n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036,
         n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046,
         n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056,
         n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066,
         n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076,
         n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086,
         n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096,
         n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106,
         n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116,
         n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126,
         n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136,
         n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146,
         n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156,
         n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166,
         n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176,
         n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
         n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196,
         n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216,
         n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226,
         n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236,
         n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
         n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
         n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266,
         n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276,
         n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286,
         n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296,
         n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
         n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
         n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
         n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
         n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346,
         n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356,
         n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366,
         n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376,
         n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
         n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416,
         n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426,
         n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436,
         n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446,
         n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456,
         n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466,
         n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476,
         n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486,
         n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496,
         n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506,
         n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516,
         n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526,
         n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536,
         n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546,
         n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566,
         n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576,
         n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586,
         n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596,
         n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606,
         n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616,
         n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626,
         n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636,
         n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
         n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
         n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
         n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
         n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
         n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
         n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
         n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
         n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
         n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
         n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756,
         n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766,
         n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776,
         n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786,
         n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796,
         n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
         n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816,
         n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846,
         n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
         n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
         n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
         n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
         n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
         n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
         n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
         n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
         n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
         n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
         n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
         n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966,
         n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976,
         n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986,
         n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996,
         n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006,
         n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016,
         n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026,
         n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036,
         n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046,
         n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056,
         n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066,
         n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076,
         n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086,
         n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096,
         n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106,
         n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
         n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
         n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
         n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
         n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156,
         n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166,
         n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176,
         n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186,
         n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236,
         n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246,
         n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256,
         n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266,
         n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276,
         n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286,
         n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296,
         n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306,
         n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316,
         n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326,
         n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336,
         n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
         n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
         n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
         n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
         n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386,
         n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396,
         n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406,
         n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416,
         n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426,
         n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436,
         n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
         n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
         n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
         n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476,
         n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486,
         n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496,
         n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506,
         n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
         n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526,
         n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536,
         n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546,
         n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556,
         n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566,
         n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576,
         n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
         n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596,
         n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606,
         n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616,
         n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626,
         n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
         n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656,
         n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666,
         n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676,
         n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686,
         n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696,
         n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706,
         n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
         n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
         n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
         n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746,
         n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756,
         n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776,
         n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786,
         n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796,
         n6797, n6798, n6799, n6800, n6801, n6802, n6803;

  NAND2_X1 U34740 ( .A1(n5516), .A2(n5296), .ZN(n5069) );
  NOR2_X1 U3475 ( .A1(n5008), .A2(n5009), .ZN(n5006) );
  NOR2_X1 U3476 ( .A1(n4676), .A2(n4607), .ZN(n4608) );
  OAI211_X1 U3477 ( .C1(n3236), .C2(n3231), .A(n3234), .B(n3233), .ZN(n3321)
         );
  CLKBUF_X2 U3478 ( .A(n3156), .Z(n5148) );
  CLKBUF_X2 U3479 ( .A(n3248), .Z(n5138) );
  CLKBUF_X2 U3480 ( .A(n3243), .Z(n5145) );
  CLKBUF_X2 U3481 ( .A(n3265), .Z(n5147) );
  CLKBUF_X2 U3482 ( .A(n3270), .Z(n5137) );
  CLKBUF_X2 U3483 ( .A(n3272), .Z(n5146) );
  CLKBUF_X2 U3484 ( .A(n3303), .Z(n5149) );
  CLKBUF_X2 U3485 ( .A(n3288), .Z(n5139) );
  CLKBUF_X2 U3486 ( .A(n3967), .Z(n4968) );
  AND4_X1 U3487 ( .A1(n3155), .A2(n3154), .A3(n3153), .A4(n3152), .ZN(n3162)
         );
  AND4_X1 U3488 ( .A1(n3116), .A2(n3115), .A3(n3114), .A4(n3113), .ZN(n3042)
         );
  AND4_X1 U3489 ( .A1(n3112), .A2(n3111), .A3(n3110), .A4(n3109), .ZN(n3117)
         );
  BUF_X2 U3490 ( .A(n3134), .Z(n3250) );
  AND2_X2 U3491 ( .A1(n3065), .A2(n4418), .ZN(n3287) );
  AND2_X2 U3492 ( .A1(n3064), .A2(n4219), .ZN(n5124) );
  AND2_X2 U3493 ( .A1(n3060), .A2(n4220), .ZN(n3308) );
  AND2_X2 U3494 ( .A1(n3065), .A2(n4416), .ZN(n3265) );
  INV_X1 U3495 ( .A(n6199), .ZN(n6183) );
  OR2_X1 U3496 ( .A1(n3967), .A2(n3944), .ZN(n3208) );
  NAND2_X1 U3497 ( .A1(n3400), .A2(n3302), .ZN(n3385) );
  NOR2_X1 U3498 ( .A1(n3280), .A2(n3337), .ZN(n3477) );
  AND4_X1 U3499 ( .A1(n3084), .A2(n3083), .A3(n3082), .A4(n3081), .ZN(n3085)
         );
  NAND2_X2 U3500 ( .A1(n4303), .A2(n4065), .ZN(n4056) );
  INV_X1 U3501 ( .A(n4065), .ZN(n5381) );
  BUF_X1 U3503 ( .A(n3982), .Z(n4303) );
  AND2_X2 U3504 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4219) );
  INV_X1 U3505 ( .A(n3379), .ZN(n4384) );
  AND2_X2 U3506 ( .A1(n4402), .A2(n3030), .ZN(n4958) );
  INV_X1 U3507 ( .A(n6039), .ZN(n6012) );
  AND2_X1 U3508 ( .A1(n6026), .A2(n4954), .ZN(n6053) );
  XNOR2_X1 U3509 ( .A(n6193), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4276)
         );
  NAND2_X1 U3510 ( .A1(n6189), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6193)
         );
  INV_X2 U3513 ( .A(n6053), .ZN(n6070) );
  OR3_X1 U3514 ( .A1(n4232), .A2(n6461), .A3(n3556), .ZN(n6190) );
  NAND2_X2 U3515 ( .A1(n3350), .A2(n4542), .ZN(n3433) );
  XNOR2_X2 U3516 ( .A(n3413), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4316)
         );
  XNOR2_X1 U3517 ( .A(n5279), .B(n5278), .ZN(n5299) );
  NAND2_X1 U3518 ( .A1(n5331), .A2(n5290), .ZN(n5789) );
  OAI22_X1 U3519 ( .A1(n5594), .A2(n3504), .B1(n4119), .B2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3505) );
  XNOR2_X1 U3520 ( .A(n4121), .B(n4120), .ZN(n5227) );
  OR2_X1 U3521 ( .A1(n5845), .A2(n5844), .ZN(n5882) );
  OR2_X1 U3522 ( .A1(n5561), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5066)
         );
  INV_X1 U3523 ( .A(n3503), .ZN(n4135) );
  NAND2_X1 U3524 ( .A1(n5173), .A2(n5343), .ZN(n5344) );
  NOR2_X1 U3525 ( .A1(n4133), .A2(n4132), .ZN(n3503) );
  OR2_X1 U3526 ( .A1(n5603), .A2(n4117), .ZN(n4118) );
  NAND2_X1 U3527 ( .A1(n4122), .A2(n3896), .ZN(n3920) );
  CLKBUF_X1 U3528 ( .A(n5402), .Z(n5421) );
  NAND2_X1 U3529 ( .A1(n3727), .A2(n3726), .ZN(n5422) );
  CLKBUF_X1 U3530 ( .A(n5013), .Z(n5256) );
  CLKBUF_X1 U3531 ( .A(n4939), .Z(n4992) );
  CLKBUF_X1 U3532 ( .A(n4920), .Z(n4941) );
  NAND3_X1 U3534 ( .A1(n4270), .A2(n3590), .A3(n4269), .ZN(n4351) );
  OAI21_X1 U3535 ( .B1(n3601), .B2(n3950), .A(n3443), .ZN(n3444) );
  NAND2_X1 U3536 ( .A1(n3412), .A2(n6176), .ZN(n4315) );
  XNOR2_X1 U3537 ( .A(n3480), .B(n3467), .ZN(n3617) );
  OR2_X1 U3538 ( .A1(n3589), .A2(n3588), .ZN(n4269) );
  NOR2_X1 U3539 ( .A1(n5197), .A2(n5572), .ZN(n5200) );
  OR2_X1 U3540 ( .A1(n3433), .A2(n3432), .ZN(n3462) );
  INV_X1 U3541 ( .A(n3557), .ZN(n3376) );
  NAND2_X1 U3542 ( .A1(n3372), .A2(n3371), .ZN(n3373) );
  AND2_X1 U3543 ( .A1(n3349), .A2(n3348), .ZN(n4506) );
  NAND2_X1 U3545 ( .A1(n3258), .A2(n3257), .ZN(n3261) );
  NAND2_X1 U3546 ( .A1(n3328), .A2(n3330), .ZN(n4445) );
  OAI21_X1 U3547 ( .B1(n4212), .B2(STATE2_REG_0__SCAN_IN), .A(n3325), .ZN(
        n3386) );
  NAND2_X1 U3548 ( .A1(n4003), .A2(n3041), .ZN(n4766) );
  CLKBUF_X1 U3549 ( .A(n4212), .Z(n5731) );
  NAND2_X1 U3550 ( .A1(n3335), .A2(n3334), .ZN(n6295) );
  AND2_X2 U3551 ( .A1(n3551), .A2(n3550), .ZN(n4232) );
  XNOR2_X1 U3552 ( .A(n3324), .B(n3323), .ZN(n4212) );
  NAND2_X1 U3553 ( .A1(n3235), .A2(n3321), .ZN(n3329) );
  OAI21_X1 U3554 ( .B1(n3236), .B2(n3237), .A(n3242), .ZN(n3328) );
  NAND2_X1 U3555 ( .A1(n3337), .A2(n3336), .ZN(n3548) );
  NAND2_X1 U3556 ( .A1(n3299), .A2(n4968), .ZN(n4076) );
  CLKBUF_X1 U3557 ( .A(n3206), .Z(n3207) );
  OR2_X1 U3558 ( .A1(n3279), .A2(n3278), .ZN(n3476) );
  BUF_X2 U3559 ( .A(n3189), .Z(n3026) );
  AND4_X1 U3560 ( .A1(n3168), .A2(n3167), .A3(n3166), .A4(n3165), .ZN(n3184)
         );
  AND4_X1 U3561 ( .A1(n3072), .A2(n3071), .A3(n3070), .A4(n3069), .ZN(n3088)
         );
  AND4_X1 U3562 ( .A1(n3104), .A2(n3103), .A3(n3102), .A4(n3101), .ZN(n3105)
         );
  AND4_X1 U3563 ( .A1(n3100), .A2(n3099), .A3(n3098), .A4(n3097), .ZN(n3106)
         );
  AND4_X1 U3564 ( .A1(n3096), .A2(n3095), .A3(n3094), .A4(n3093), .ZN(n3107)
         );
  AND4_X1 U3565 ( .A1(n3092), .A2(n3091), .A3(n3090), .A4(n3089), .ZN(n3108)
         );
  AND4_X1 U3566 ( .A1(n3138), .A2(n3137), .A3(n3136), .A4(n3135), .ZN(n3048)
         );
  AND3_X1 U3567 ( .A1(n3063), .A2(n3062), .A3(n3061), .ZN(n3067) );
  AND4_X1 U3568 ( .A1(n3080), .A2(n3079), .A3(n3078), .A4(n3077), .ZN(n3086)
         );
  AND4_X1 U3569 ( .A1(n3076), .A2(n3075), .A3(n3074), .A4(n3073), .ZN(n3087)
         );
  BUF_X2 U3570 ( .A(n3287), .Z(n5144) );
  BUF_X2 U3571 ( .A(n3249), .Z(n3027) );
  AND2_X2 U3572 ( .A1(n3054), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4226)
         );
  CLKBUF_X1 U3573 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n6575) );
  AND2_X2 U3574 ( .A1(n3060), .A2(n3065), .ZN(n3243) );
  NAND2_X1 U3576 ( .A1(n4301), .A2(n4303), .ZN(n4302) );
  XNOR2_X1 U3577 ( .A(n3981), .B(n4196), .ZN(n4301) );
  XNOR2_X1 U3578 ( .A(n3329), .B(n3328), .ZN(n4375) );
  OAI22_X2 U3579 ( .A1(n4316), .A2(n4315), .B1(n3414), .B2(n5055), .ZN(n5050)
         );
  AND2_X2 U3580 ( .A1(n4084), .A2(n3205), .ZN(n3227) );
  AND2_X1 U3582 ( .A1(n3064), .A2(n4219), .ZN(n3028) );
  AND2_X2 U3583 ( .A1(n5265), .A2(n5264), .ZN(n5367) );
  NOR2_X2 U3584 ( .A1(n5380), .A2(n4041), .ZN(n5265) );
  BUF_X2 U3585 ( .A(n3151), .Z(n3290) );
  NAND4_X1 U3586 ( .A1(n3164), .A2(n3163), .A3(n3162), .A4(n3161), .ZN(n3029)
         );
  NAND4_X1 U3587 ( .A1(n3164), .A2(n3163), .A3(n3162), .A4(n3161), .ZN(n3030)
         );
  NAND4_X4 U3588 ( .A1(n3184), .A2(n3183), .A3(n3182), .A4(n3181), .ZN(n3967)
         );
  OAI21_X2 U3589 ( .B1(n6152), .B2(n6153), .A(n6154), .ZN(n5017) );
  AOI21_X2 U3590 ( .B1(n4978), .B2(n4979), .A(n4981), .ZN(n6152) );
  AND2_X1 U3591 ( .A1(n5576), .A2(n3935), .ZN(n5560) );
  NAND2_X1 U3592 ( .A1(n3400), .A2(n3399), .ZN(n3569) );
  MUX2_X2 U3593 ( .A(n5070), .B(n5381), .S(n5069), .Z(n5073) );
  AOI21_X2 U3594 ( .B1(n4532), .B2(n4531), .A(n3034), .ZN(n4934) );
  NAND4_X1 U3595 ( .A1(n3164), .A2(n3163), .A3(n3162), .A4(n3161), .ZN(n3033)
         );
  AOI21_X2 U3596 ( .B1(n4909), .B2(n4910), .A(n3485), .ZN(n4997) );
  OAI21_X2 U3597 ( .B1(n4934), .B2(n4933), .A(n3475), .ZN(n4909) );
  NOR2_X2 U3598 ( .A1(n5348), .A2(n5347), .ZN(n5522) );
  OR2_X2 U3599 ( .A1(n5228), .A2(n5217), .ZN(n5348) );
  NOR2_X2 U3600 ( .A1(n4344), .A2(n4345), .ZN(n4364) );
  NOR2_X1 U3601 ( .A1(n3226), .A2(n3225), .ZN(n3229) );
  CLKBUF_X1 U3602 ( .A(n3227), .Z(n3228) );
  NAND2_X1 U3603 ( .A1(n4431), .A2(n3219), .ZN(n3226) );
  OR2_X1 U3604 ( .A1(n4072), .A2(n6780), .ZN(n3337) );
  NAND3_X1 U3605 ( .A1(n4072), .A2(n3030), .A3(STATE2_REG_0__SCAN_IN), .ZN(
        n3536) );
  NAND2_X1 U3606 ( .A1(n3264), .A2(n3262), .ZN(n3322) );
  XNOR2_X1 U3607 ( .A(n4445), .B(n6295), .ZN(n4374) );
  CLKBUF_X1 U3608 ( .A(n3308), .Z(n5136) );
  OR2_X1 U3609 ( .A1(n3256), .A2(n3255), .ZN(n3365) );
  NOR2_X1 U3610 ( .A1(n4075), .A2(n3210), .ZN(n3211) );
  AOI22_X1 U3611 ( .A1(n3248), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3063) );
  NAND2_X1 U3613 ( .A1(n3459), .A2(n3460), .ZN(n3480) );
  AND2_X2 U3614 ( .A1(n4226), .A2(n4418), .ZN(n3146) );
  AND2_X2 U3615 ( .A1(n4226), .A2(n4416), .ZN(n3272) );
  AND2_X2 U3616 ( .A1(n3060), .A2(n4226), .ZN(n3270) );
  NOR2_X2 U3617 ( .A1(n5344), .A2(n5518), .ZN(n5508) );
  NOR2_X2 U3618 ( .A1(n3920), .A2(n3919), .ZN(n5173) );
  AND2_X1 U3619 ( .A1(n5402), .A2(n5403), .ZN(n4122) );
  NOR2_X1 U3620 ( .A1(n5422), .A2(n5423), .ZN(n5402) );
  NAND2_X1 U3621 ( .A1(n3462), .A2(n3461), .ZN(n3614) );
  NAND2_X1 U3622 ( .A1(n3433), .A2(n3430), .ZN(n3364) );
  INV_X1 U3623 ( .A(n3724), .ZN(n3739) );
  NAND2_X1 U3624 ( .A1(n5890), .A2(n3491), .ZN(n3492) );
  INV_X1 U3625 ( .A(n4415), .ZN(n4200) );
  NOR2_X2 U3626 ( .A1(n5331), .A2(n5332), .ZN(n5330) );
  NAND2_X1 U3627 ( .A1(n5895), .A2(n5894), .ZN(n5897) );
  CLKBUF_X1 U3628 ( .A(n4122), .Z(n5895) );
  NOR2_X1 U3629 ( .A1(n3484), .A2(n4005), .ZN(n3485) );
  AND2_X1 U3630 ( .A1(n4608), .A2(n4787), .ZN(n4922) );
  NOR2_X1 U3631 ( .A1(n3602), .A2(n6175), .ZN(n3609) );
  NAND2_X1 U3632 ( .A1(n3609), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3618)
         );
  NAND2_X1 U3633 ( .A1(n3616), .A2(n3615), .ZN(n4676) );
  INV_X1 U3634 ( .A(n4679), .ZN(n3615) );
  INV_X1 U3635 ( .A(n4678), .ZN(n3616) );
  NAND2_X1 U3636 ( .A1(n3595), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3602)
         );
  INV_X1 U3637 ( .A(n4198), .ZN(n4069) );
  NAND2_X1 U3638 ( .A1(n3500), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3498) );
  OR2_X1 U3639 ( .A1(n6583), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3926) );
  INV_X1 U3640 ( .A(n5025), .ZN(n6236) );
  CLKBUF_X1 U3641 ( .A(n3941), .Z(n3942) );
  NAND2_X1 U3642 ( .A1(n3044), .A2(n3186), .ZN(n4073) );
  OR2_X1 U3643 ( .A1(n5733), .A2(n4542), .ZN(n5737) );
  INV_X1 U3644 ( .A(n3549), .ZN(n3550) );
  AOI21_X1 U3645 ( .B1(n3548), .B2(n3958), .A(n3547), .ZN(n3549) );
  OR2_X1 U3646 ( .A1(n5737), .A2(n5744), .ZN(n6260) );
  OR2_X1 U3647 ( .A1(n5737), .A2(n4614), .ZN(n6288) );
  NOR2_X1 U3648 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4383), .ZN(n4582) );
  AND2_X1 U3649 ( .A1(n6765), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3555) );
  INV_X1 U3650 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6486) );
  AND2_X1 U3651 ( .A1(n5293), .A2(n3186), .ZN(n6610) );
  INV_X1 U3652 ( .A(n5293), .ZN(n6608) );
  AND2_X1 U3653 ( .A1(n5293), .A2(n4299), .ZN(n5557) );
  INV_X1 U3654 ( .A(n6174), .ZN(n6196) );
  NAND2_X1 U3655 ( .A1(n4119), .A2(n4118), .ZN(n4121) );
  INV_X1 U3656 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6256) );
  AND2_X1 U3657 ( .A1(n3218), .A2(n6485), .ZN(n3219) );
  NOR2_X1 U3658 ( .A1(n3518), .A2(n3517), .ZN(n3516) );
  OAI211_X1 U3659 ( .C1(n3026), .C2(n3192), .A(n3191), .B(n3194), .ZN(n3193)
         );
  NAND2_X1 U3660 ( .A1(n3026), .A2(n3190), .ZN(n3191) );
  AND2_X2 U3661 ( .A1(n3053), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3065)
         );
  CLKBUF_X1 U3662 ( .A(n5124), .Z(n3734) );
  OR2_X1 U3663 ( .A1(n3427), .A2(n3426), .ZN(n3441) );
  NAND2_X1 U3664 ( .A1(n3196), .A2(n4072), .ZN(n3222) );
  AND2_X2 U3665 ( .A1(n3059), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3064)
         );
  INV_X1 U3666 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3059) );
  OR2_X1 U3668 ( .A1(n3315), .A2(n3314), .ZN(n3390) );
  AOI22_X1 U3669 ( .A1(n3544), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3259), 
        .B2(n3365), .ZN(n3260) );
  OR2_X1 U3670 ( .A1(n3033), .A2(n6780), .ZN(n3336) );
  AOI21_X1 U3671 ( .B1(n6575), .B2(n6458), .A(n3516), .ZN(n3514) );
  NOR2_X1 U3672 ( .A1(n6460), .A2(n3974), .ZN(n4086) );
  NAND2_X1 U3673 ( .A1(n3194), .A2(n3379), .ZN(n4077) );
  AND2_X2 U3674 ( .A1(n4219), .A2(n4416), .ZN(n3134) );
  AND2_X2 U3675 ( .A1(n3060), .A2(n4219), .ZN(n3156) );
  INV_X1 U3676 ( .A(n3536), .ZN(n3544) );
  OR2_X1 U3677 ( .A1(n3347), .A2(n3346), .ZN(n3369) );
  AND2_X2 U3678 ( .A1(n4418), .A2(n4219), .ZN(n3151) );
  AND2_X1 U3679 ( .A1(n3895), .A2(n4123), .ZN(n3896) );
  NAND2_X1 U3680 ( .A1(n3697), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3710)
         );
  NAND2_X1 U3681 ( .A1(n3665), .A2(n3664), .ZN(n4939) );
  INV_X1 U3682 ( .A(n4920), .ZN(n3665) );
  INV_X1 U3683 ( .A(n6575), .ZN(n3585) );
  NAND2_X1 U3684 ( .A1(n3560), .A2(n3912), .ZN(n3589) );
  OR2_X1 U3685 ( .A1(n4371), .A2(n3724), .ZN(n3560) );
  BUF_X1 U3686 ( .A(n3190), .Z(n3187) );
  OR2_X1 U3687 ( .A1(n3983), .A2(EBX_REG_1__SCAN_IN), .ZN(n3977) );
  INV_X1 U3688 ( .A(n4077), .ZN(n3391) );
  INV_X1 U3689 ( .A(n4072), .ZN(n3298) );
  AND2_X2 U3690 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4416) );
  INV_X1 U3691 ( .A(n3204), .ZN(n3954) );
  INV_X1 U3692 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6445) );
  INV_X1 U3693 ( .A(n4965), .ZN(n3299) );
  CLKBUF_X1 U3694 ( .A(n4144), .Z(n4145) );
  AND3_X1 U3695 ( .A1(n3744), .A2(n3743), .A3(n3742), .ZN(n5423) );
  INV_X1 U3696 ( .A(n5510), .ZN(n5191) );
  AND2_X1 U3697 ( .A1(n5172), .A2(n5171), .ZN(n5343) );
  OR2_X1 U3698 ( .A1(n5881), .A2(n5211), .ZN(n5171) );
  NAND2_X1 U3699 ( .A1(n3786), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3910)
         );
  NOR2_X1 U3700 ( .A1(n3910), .A2(n6636), .ZN(n5169) );
  NOR2_X1 U3701 ( .A1(n3835), .A2(n5606), .ZN(n3802) );
  NAND2_X1 U3702 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n3851), .ZN(n3835)
         );
  NOR2_X1 U3703 ( .A1(n3870), .A2(n6758), .ZN(n3851) );
  AND2_X1 U3704 ( .A1(n3784), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3871)
         );
  NAND2_X1 U3705 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n3871), .ZN(n3870)
         );
  NOR2_X1 U3706 ( .A1(n3729), .A2(n6771), .ZN(n3784) );
  NOR2_X1 U3707 ( .A1(n3710), .A2(n5982), .ZN(n3728) );
  INV_X1 U3708 ( .A(n5257), .ZN(n3726) );
  INV_X1 U3709 ( .A(n5013), .ZN(n3727) );
  NOR2_X1 U3710 ( .A1(n3681), .A2(n5996), .ZN(n3697) );
  CLKBUF_X1 U3711 ( .A(n5006), .Z(n5007) );
  NAND2_X1 U3712 ( .A1(n3666), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3681)
         );
  NOR2_X1 U3713 ( .A1(n3500), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6153)
         );
  NAND2_X1 U3714 ( .A1(n3680), .A2(n3679), .ZN(n5008) );
  INV_X1 U3715 ( .A(n4939), .ZN(n3680) );
  NOR2_X1 U3716 ( .A1(n3649), .A2(n6006), .ZN(n3666) );
  NAND2_X1 U3717 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n3636), .ZN(n3649)
         );
  AOI21_X1 U3718 ( .B1(n3617), .B2(n3739), .A(n3622), .ZN(n4607) );
  CLKBUF_X1 U3719 ( .A(n4608), .Z(n4609) );
  AOI21_X1 U3720 ( .B1(n3614), .B2(n3739), .A(n3613), .ZN(n4679) );
  NAND2_X1 U3721 ( .A1(n3608), .A2(n3607), .ZN(n4347) );
  OR2_X1 U3722 ( .A1(n3601), .A2(n3724), .ZN(n3608) );
  AOI21_X1 U3723 ( .B1(n3600), .B2(n3739), .A(n3599), .ZN(n4343) );
  NOR2_X2 U3724 ( .A1(n4351), .A2(n4343), .ZN(n4348) );
  NOR2_X1 U3725 ( .A1(n3581), .A2(n4359), .ZN(n3595) );
  AND2_X1 U3726 ( .A1(n5513), .A2(n5514), .ZN(n5516) );
  AND2_X1 U3727 ( .A1(n5522), .A2(n5521), .ZN(n5513) );
  NOR2_X1 U3728 ( .A1(n5698), .A2(n3933), .ZN(n3934) );
  OR2_X1 U3729 ( .A1(n5369), .A2(n5230), .ZN(n5228) );
  NAND2_X1 U3730 ( .A1(n5367), .A2(n5366), .ZN(n5369) );
  AND2_X1 U3731 ( .A1(n5890), .A2(n5705), .ZN(n3497) );
  XOR2_X1 U3733 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .B(n5890), .Z(n5629) );
  CLKBUF_X1 U3734 ( .A(n5613), .Z(n5614) );
  NOR2_X1 U3735 ( .A1(n4101), .A2(n4415), .ZN(n5025) );
  AND2_X1 U3736 ( .A1(n5890), .A2(n6234), .ZN(n3486) );
  AND2_X1 U3737 ( .A1(n4011), .A2(n4010), .ZN(n4925) );
  NAND2_X1 U3738 ( .A1(n4926), .A2(n4925), .ZN(n4988) );
  NOR2_X2 U3739 ( .A1(n4766), .A2(n4765), .ZN(n4913) );
  INV_X1 U3740 ( .A(n6213), .ZN(n5720) );
  AND2_X1 U3741 ( .A1(n3994), .A2(n3993), .ZN(n4345) );
  NAND2_X1 U3742 ( .A1(n3990), .A2(n3989), .ZN(n4344) );
  INV_X1 U3743 ( .A(n4321), .ZN(n3990) );
  NOR2_X1 U3744 ( .A1(n4319), .A2(n4320), .ZN(n3989) );
  AND2_X1 U3745 ( .A1(n4048), .A2(n3031), .ZN(n4198) );
  BUF_X1 U3746 ( .A(n3557), .Z(n4371) );
  CLKBUF_X1 U3747 ( .A(n4375), .Z(n5491) );
  INV_X1 U3748 ( .A(n3507), .ZN(n6438) );
  CLKBUF_X1 U3749 ( .A(n3571), .Z(n6441) );
  INV_X1 U3750 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6765) );
  NAND2_X1 U3751 ( .A1(n3199), .A2(n3954), .ZN(n4216) );
  NOR2_X1 U3752 ( .A1(n4147), .A2(n6460), .ZN(n3199) );
  AND2_X1 U3753 ( .A1(n4211), .A2(n4210), .ZN(n6448) );
  CLKBUF_X1 U3754 ( .A(n4374), .Z(n5747) );
  OR2_X1 U3755 ( .A1(n6260), .A2(n6487), .ZN(n4543) );
  NOR2_X1 U3756 ( .A1(n5742), .A2(n3376), .ZN(n6371) );
  INV_X1 U3757 ( .A(n6263), .ZN(n6380) );
  CLKBUF_X1 U3758 ( .A(n3299), .Z(n4409) );
  CLKBUF_X1 U3759 ( .A(n3558), .Z(n3559) );
  OR2_X1 U3760 ( .A1(n6567), .A2(n4383), .ZN(n4583) );
  INV_X1 U3761 ( .A(n6064), .ZN(n6048) );
  AND2_X1 U3762 ( .A1(n6094), .A2(n5286), .ZN(n6081) );
  CLKBUF_X1 U3763 ( .A(n5533), .Z(n6085) );
  INV_X1 U3764 ( .A(n6081), .ZN(n6090) );
  INV_X1 U3765 ( .A(n5882), .ZN(n5870) );
  NAND2_X1 U3766 ( .A1(n4297), .A2(n4296), .ZN(n5293) );
  INV_X1 U3767 ( .A(n5557), .ZN(n5010) );
  INV_X1 U3768 ( .A(n6133), .ZN(n6103) );
  OR2_X1 U3769 ( .A1(n5202), .A2(n5323), .ZN(n4949) );
  XOR2_X1 U3770 ( .A(n5274), .B(n5330), .Z(n5319) );
  AND2_X1 U3771 ( .A1(n5897), .A2(n5896), .ZN(n6612) );
  INV_X1 U3772 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6175) );
  INV_X1 U3773 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n4359) );
  NAND2_X1 U3774 ( .A1(n6190), .A2(n3923), .ZN(n6174) );
  XNOR2_X1 U3775 ( .A(n3940), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5285)
         );
  NOR2_X1 U3776 ( .A1(n5682), .A2(n4112), .ZN(n5906) );
  NAND2_X1 U3777 ( .A1(n4133), .A2(n4132), .ZN(n4134) );
  NOR2_X1 U3778 ( .A1(n5247), .A2(n5024), .ZN(n6201) );
  INV_X1 U3779 ( .A(n6203), .ZN(n6247) );
  AND2_X1 U3780 ( .A1(n4093), .A2(n4074), .ZN(n6240) );
  CLKBUF_X1 U3781 ( .A(n4371), .Z(n5733) );
  INV_X1 U3782 ( .A(n5747), .ZN(n5740) );
  CLKBUF_X1 U3783 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n3507) );
  INV_X1 U3784 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3054) );
  NOR2_X1 U3785 ( .A1(n6569), .A2(n4232), .ZN(n5038) );
  OR2_X1 U3786 ( .A1(n6260), .A2(n6287), .ZN(n6266) );
  OR3_X1 U3787 ( .A1(n6302), .A2(n6301), .A3(n6300), .ZN(n6334) );
  OAI211_X1 U3788 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6486), .A(n5755), .B(n5754), .ZN(n5777) );
  OR2_X1 U3789 ( .A1(n4465), .A2(n6287), .ZN(n4807) );
  INV_X1 U3790 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6569) );
  INV_X1 U3791 ( .A(n6492), .ZN(n6568) );
  INV_X1 U3792 ( .A(n4129), .ZN(n4130) );
  OAI21_X1 U3793 ( .B1(n5823), .B2(n6199), .A(n4128), .ZN(n4129) );
  NAND2_X1 U3794 ( .A1(n3480), .A2(n3479), .ZN(n3488) );
  AND2_X1 U3795 ( .A1(n3465), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3034)
         );
  NOR2_X2 U3796 ( .A1(n6767), .A2(n6605), .ZN(n6556) );
  CLKBUF_X3 U3797 ( .A(n3271), .Z(n5100) );
  AND2_X2 U3798 ( .A1(n4220), .A2(n4416), .ZN(n3303) );
  AND2_X1 U3799 ( .A1(n3996), .A2(n3995), .ZN(n3035) );
  OR2_X1 U3800 ( .A1(n3500), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3036)
         );
  AND2_X1 U3801 ( .A1(n3500), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3037)
         );
  AND2_X1 U3802 ( .A1(n5890), .A2(n4094), .ZN(n3038) );
  AND2_X1 U3803 ( .A1(n5890), .A2(n5721), .ZN(n3039) );
  OR2_X1 U3804 ( .A1(n3500), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3040)
         );
  NAND2_X1 U3805 ( .A1(n4002), .A2(n4001), .ZN(n3041) );
  INV_X1 U3806 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3367) );
  AND3_X1 U3807 ( .A1(n3144), .A2(n3143), .A3(n3142), .ZN(n3043) );
  AND3_X1 U3808 ( .A1(n3969), .A2(n3185), .A3(n4384), .ZN(n3044) );
  INV_X1 U3809 ( .A(n3946), .ZN(n3186) );
  NAND2_X1 U3810 ( .A1(n3558), .A2(n5291), .ZN(n3215) );
  AND4_X1 U3811 ( .A1(n3133), .A2(n3132), .A3(n3131), .A4(n3130), .ZN(n3045)
         );
  AND2_X1 U3812 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3046) );
  INV_X1 U3813 ( .A(n4534), .ZN(n4003) );
  NOR2_X2 U3814 ( .A1(n6288), .A2(n3032), .ZN(n3047) );
  INV_X1 U3815 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3237) );
  OR2_X1 U3816 ( .A1(n3366), .A2(n6599), .ZN(n3049) );
  AND2_X1 U3817 ( .A1(n3362), .A2(n3361), .ZN(n3430) );
  BUF_X1 U3818 ( .A(n3983), .Z(n4065) );
  INV_X1 U3819 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3231) );
  OR2_X1 U3820 ( .A1(n3463), .A2(n6599), .ZN(n3050) );
  AND2_X1 U3821 ( .A1(n3188), .A2(n5291), .ZN(n3051) );
  INV_X1 U3822 ( .A(n3430), .ZN(n3431) );
  NAND2_X1 U3823 ( .A1(n3434), .A2(n3431), .ZN(n3432) );
  OR2_X1 U3824 ( .A1(n3360), .A2(n3359), .ZN(n3438) );
  NAND2_X1 U3825 ( .A1(n3051), .A2(n3298), .ZN(n3951) );
  INV_X1 U3826 ( .A(n4420), .ZN(n5129) );
  AOI21_X1 U3827 ( .B1(n3535), .B2(n3512), .A(n3511), .ZN(n3518) );
  INV_X1 U3828 ( .A(n4942), .ZN(n3664) );
  OR2_X1 U3829 ( .A1(n4188), .A2(n4576), .ZN(n3216) );
  INV_X1 U3830 ( .A(n3462), .ZN(n3459) );
  NAND2_X1 U3831 ( .A1(n3376), .A2(n3375), .ZN(n3382) );
  NAND2_X1 U3832 ( .A1(n3379), .A2(n3967), .ZN(n3974) );
  AND2_X1 U3833 ( .A1(n3220), .A2(n5291), .ZN(n3197) );
  INV_X1 U3834 ( .A(n3891), .ZN(n3785) );
  INV_X1 U3835 ( .A(n3888), .ZN(n3916) );
  OR2_X1 U3836 ( .A1(n6437), .A2(n6780), .ZN(n5208) );
  INV_X1 U3837 ( .A(n3916), .ZN(n5276) );
  NAND4_X2 U3838 ( .A1(n3088), .A2(n3087), .A3(n3086), .A4(n3085), .ZN(n3190)
         );
  INV_X1 U3839 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3491) );
  OR2_X1 U3840 ( .A1(n3297), .A2(n3296), .ZN(n3403) );
  INV_X1 U3841 ( .A(n3329), .ZN(n3330) );
  NAND2_X1 U3842 ( .A1(n4374), .A2(n6780), .ZN(n3349) );
  AND2_X1 U3843 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n3785), .ZN(n3786)
         );
  CLKBUF_X1 U3844 ( .A(n3969), .Z(n4948) );
  OR2_X1 U3845 ( .A1(n4092), .A2(n4090), .ZN(n4415) );
  NAND2_X1 U3846 ( .A1(n5124), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3145)
         );
  OR2_X1 U3847 ( .A1(n5179), .A2(n5590), .ZN(n5187) );
  OR2_X1 U3848 ( .A1(n5897), .A2(n5390), .ZN(n5843) );
  INV_X1 U3849 ( .A(n6177), .ZN(n6178) );
  NOR2_X1 U3850 ( .A1(n3536), .A2(n3950), .ZN(n3533) );
  INV_X1 U3851 ( .A(n3488), .ZN(n3500) );
  INV_X1 U3852 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3410) );
  NAND2_X1 U3854 ( .A1(n3571), .A2(n6780), .ZN(n3400) );
  NOR2_X1 U3855 ( .A1(n6167), .A2(n3618), .ZN(n3636) );
  INV_X1 U3856 ( .A(n6034), .ZN(n6069) );
  NAND2_X1 U3857 ( .A1(n4971), .A2(n4970), .ZN(n6046) );
  INV_X1 U3858 ( .A(n5071), .ZN(n5072) );
  AND2_X1 U3859 ( .A1(n4136), .A2(n3894), .ZN(n4123) );
  NAND2_X1 U3860 ( .A1(n4922), .A2(n4921), .ZN(n4920) );
  AND2_X1 U3861 ( .A1(n3043), .A2(n3145), .ZN(n3164) );
  OR2_X1 U3862 ( .A1(n5187), .A2(n5580), .ZN(n5197) );
  OR2_X1 U3863 ( .A1(n5377), .A2(n4139), .ZN(n4140) );
  NOR2_X1 U3864 ( .A1(n5890), .A2(n6224), .ZN(n4981) );
  OR2_X1 U3865 ( .A1(n5875), .A2(n3937), .ZN(n3938) );
  NOR2_X1 U3866 ( .A1(n5617), .A2(n5712), .ZN(n5686) );
  NAND2_X1 U3867 ( .A1(n4135), .A2(n3502), .ZN(n5594) );
  AND2_X1 U3868 ( .A1(n5890), .A2(n3494), .ZN(n3495) );
  NOR2_X2 U3869 ( .A1(n5425), .A2(n5424), .ZN(n5427) );
  XNOR2_X1 U3870 ( .A(n5890), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5638)
         );
  INV_X1 U3871 ( .A(n6240), .ZN(n6229) );
  INV_X1 U3872 ( .A(n4287), .ZN(n5241) );
  OR2_X1 U3874 ( .A1(n4541), .A2(n3032), .ZN(n4769) );
  INV_X1 U3875 ( .A(n5744), .ZN(n4614) );
  INV_X1 U3876 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6452) );
  INV_X1 U3877 ( .A(n6430), .ZN(n5780) );
  AOI21_X1 U3878 ( .B1(n6493), .B2(n4453), .A(n5038), .ZN(n4383) );
  OR2_X1 U3879 ( .A1(n4465), .A2(n3032), .ZN(n4806) );
  INV_X1 U3880 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6458) );
  NAND2_X1 U3881 ( .A1(n4229), .A2(n4163), .ZN(n6594) );
  AND2_X1 U3882 ( .A1(n6026), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6034) );
  NAND2_X1 U3883 ( .A1(n3802), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3891)
         );
  AND2_X1 U3884 ( .A1(n4964), .A2(n4963), .ZN(n6064) );
  OR2_X1 U3885 ( .A1(n6594), .A2(n4947), .ZN(n6026) );
  AND2_X1 U3886 ( .A1(n6026), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4971) );
  AND2_X1 U3887 ( .A1(n4971), .A2(n4961), .ZN(n6051) );
  AND2_X1 U3888 ( .A1(n4138), .A2(n4137), .ZN(n5377) );
  OR2_X1 U3889 ( .A1(n4988), .A2(n4987), .ZN(n5993) );
  AND2_X1 U3890 ( .A1(n5293), .A2(n5292), .ZN(n6609) );
  NAND2_X1 U3891 ( .A1(n5169), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5179)
         );
  AND2_X1 U3892 ( .A1(n5360), .A2(n4140), .ZN(n5864) );
  NAND2_X1 U3893 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3581) );
  INV_X1 U3894 ( .A(n6188), .ZN(n6168) );
  NAND2_X1 U3895 ( .A1(n3939), .A2(n3938), .ZN(n3940) );
  INV_X1 U3896 ( .A(n5576), .ZN(n5589) );
  AND2_X1 U3897 ( .A1(n5686), .A2(n4095), .ZN(n5900) );
  OR2_X1 U3898 ( .A1(n5271), .A2(n5677), .ZN(n5682) );
  NOR2_X1 U3899 ( .A1(n5698), .A2(n5697), .ZN(n5696) );
  CLKBUF_X1 U3900 ( .A(n5017), .Z(n5019) );
  NAND2_X1 U3901 ( .A1(n5241), .A2(n4285), .ZN(n6213) );
  AND2_X1 U3902 ( .A1(n3966), .A2(n6484), .ZN(n4093) );
  AND2_X1 U3903 ( .A1(n4483), .A2(n3032), .ZN(n4704) );
  NOR2_X1 U3904 ( .A1(n4699), .A2(n3032), .ZN(n4782) );
  INV_X1 U3905 ( .A(n4769), .ZN(n4592) );
  INV_X1 U3906 ( .A(n6266), .ZN(n6282) );
  INV_X1 U3907 ( .A(n6294), .ZN(n6333) );
  INV_X1 U3908 ( .A(n6342), .ZN(n6364) );
  AND2_X1 U3909 ( .A1(n6371), .A2(n5745), .ZN(n6430) );
  AND2_X1 U3910 ( .A1(n6371), .A2(n4505), .ZN(n6429) );
  INV_X1 U3911 ( .A(n3032), .ZN(n6287) );
  INV_X1 U3912 ( .A(n4807), .ZN(n4670) );
  INV_X1 U3913 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6767) );
  OR3_X1 U3914 ( .A1(n4232), .A2(n6482), .A3(n4145), .ZN(n4229) );
  INV_X1 U3915 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6780) );
  NAND2_X1 U3916 ( .A1(n6026), .A2(n4950), .ZN(n6039) );
  INV_X1 U3917 ( .A(n6051), .ZN(n6078) );
  XNOR2_X1 U3918 ( .A(n5069), .B(n5335), .ZN(n5643) );
  OR2_X1 U3919 ( .A1(n5377), .A2(n5376), .ZN(n5607) );
  INV_X1 U3920 ( .A(n5319), .ZN(n5543) );
  OAI21_X1 U3921 ( .B1(n5520), .B2(n5519), .A(n5509), .ZN(n5806) );
  NAND2_X1 U3922 ( .A1(n5293), .A2(n4298), .ZN(n5857) );
  NOR2_X1 U3923 ( .A1(n6597), .A2(n6103), .ZN(n6120) );
  OR3_X1 U3924 ( .A1(n4232), .A2(n4168), .A3(n4167), .ZN(n6133) );
  AND2_X1 U3925 ( .A1(n3930), .A2(n3929), .ZN(n3931) );
  INV_X1 U3926 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6167) );
  NAND2_X1 U3927 ( .A1(n6174), .A2(n6195), .ZN(n6188) );
  XNOR2_X1 U3928 ( .A(n5068), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5216)
         );
  NAND2_X1 U3929 ( .A1(n4093), .A2(n3973), .ZN(n6203) );
  AND2_X1 U3930 ( .A1(n4378), .A2(n4377), .ZN(n4606) );
  INV_X1 U3931 ( .A(n4782), .ZN(n4844) );
  OR2_X1 U3932 ( .A1(n6288), .A2(n6287), .ZN(n6342) );
  NAND2_X1 U3933 ( .A1(n4612), .A2(n3032), .ZN(n4891) );
  INV_X1 U3934 ( .A(n6429), .ZN(n4831) );
  NOR2_X1 U3935 ( .A1(n4642), .A2(n4641), .ZN(n4675) );
  AND2_X1 U3936 ( .A1(n6477), .A2(n6476), .ZN(n6492) );
  INV_X1 U3937 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3052) );
  AND2_X2 U3938 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n3052), .ZN(n3060)
         );
  INV_X1 U3939 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3053) );
  NOR2_X4 U3940 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4220) );
  NOR2_X4 U3942 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4418) );
  AOI22_X1 U3944 ( .A1(n3265), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3057) );
  AOI22_X1 U3945 ( .A1(n3303), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3056) );
  AOI22_X1 U3946 ( .A1(n3272), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3055) );
  AND2_X2 U3948 ( .A1(n3064), .A2(n3065), .ZN(n3248) );
  AND2_X2 U3949 ( .A1(n3064), .A2(n4220), .ZN(n3249) );
  AOI22_X1 U3950 ( .A1(n3249), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3062) );
  AND2_X2 U3951 ( .A1(n3064), .A2(n4226), .ZN(n3288) );
  AOI22_X1 U3952 ( .A1(n3288), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3146), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3061) );
  AOI22_X1 U3953 ( .A1(n5124), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3066) );
  NAND3_X2 U3954 ( .A1(n3068), .A2(n3067), .A3(n3066), .ZN(n3189) );
  INV_X2 U3955 ( .A(n3189), .ZN(n3558) );
  NAND2_X1 U3956 ( .A1(n3287), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3072) );
  NAND2_X1 U3957 ( .A1(n3308), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3071) );
  NAND2_X1 U3958 ( .A1(n3288), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3070) );
  NAND2_X1 U3959 ( .A1(n3146), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3069) );
  NAND2_X1 U3960 ( .A1(n3248), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3076)
         );
  NAND2_X1 U3961 ( .A1(n3270), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3075) );
  NAND2_X1 U3962 ( .A1(n3249), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3074) );
  NAND2_X1 U3963 ( .A1(n3156), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3073) );
  NAND2_X1 U3964 ( .A1(n3265), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3080)
         );
  NAND2_X1 U3965 ( .A1(n3272), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3079)
         );
  NAND2_X1 U3966 ( .A1(n3151), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3078) );
  NAND2_X1 U3967 ( .A1(n3134), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3077)
         );
  NAND2_X1 U3968 ( .A1(n5124), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3084)
         );
  NAND2_X1 U3969 ( .A1(n3243), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3083) );
  NAND2_X1 U3970 ( .A1(n3303), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3082)
         );
  NAND2_X1 U3971 ( .A1(n3309), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3081) );
  NAND2_X2 U3972 ( .A1(n3558), .A2(n3190), .ZN(n3196) );
  NAND2_X1 U3973 ( .A1(n3248), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3092)
         );
  NAND2_X1 U3974 ( .A1(n3270), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3091) );
  NAND2_X1 U3975 ( .A1(n3249), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3090) );
  NAND2_X1 U3976 ( .A1(n3156), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3089) );
  NAND2_X1 U3977 ( .A1(n3288), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3096) );
  NAND2_X1 U3978 ( .A1(n3146), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3095) );
  NAND2_X1 U3979 ( .A1(n3265), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3094)
         );
  NAND2_X1 U3980 ( .A1(n3309), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3093) );
  NAND2_X1 U3981 ( .A1(n5124), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3100)
         );
  NAND2_X1 U3982 ( .A1(n3308), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3099) );
  NAND2_X1 U3983 ( .A1(n3243), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3098) );
  NAND2_X1 U3984 ( .A1(n3287), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3097) );
  NAND2_X1 U3985 ( .A1(n3272), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3104)
         );
  NAND2_X1 U3986 ( .A1(n3151), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3103) );
  NAND2_X1 U3987 ( .A1(n3303), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3102)
         );
  NAND2_X1 U3988 ( .A1(n3134), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3101)
         );
  AND4_X2 U3989 ( .A1(n3108), .A2(n3107), .A3(n3106), .A4(n3105), .ZN(n4576)
         );
  INV_X1 U3990 ( .A(n4576), .ZN(n4072) );
  AOI22_X1 U3991 ( .A1(n3243), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3028), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3112) );
  AOI22_X1 U3992 ( .A1(n3248), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3270), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3111) );
  AOI22_X1 U3993 ( .A1(n3146), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3110) );
  AOI22_X1 U3994 ( .A1(n3272), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3109) );
  AOI22_X1 U3995 ( .A1(n3308), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3116) );
  AOI22_X1 U3996 ( .A1(n3288), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U3997 ( .A1(n3249), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3114) );
  AOI22_X1 U3998 ( .A1(n3303), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3113) );
  NAND2_X2 U3999 ( .A1(n3117), .A2(n3042), .ZN(n4188) );
  BUF_X1 U4000 ( .A(n3308), .Z(n3281) );
  AOI22_X1 U4001 ( .A1(n5124), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3121) );
  AOI22_X1 U4002 ( .A1(n3243), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3120) );
  AOI22_X1 U4003 ( .A1(n3270), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3249), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3119) );
  AOI22_X1 U4004 ( .A1(n3265), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3118) );
  NAND4_X1 U4005 ( .A1(n3121), .A2(n3120), .A3(n3119), .A4(n3118), .ZN(n3127)
         );
  AOI22_X1 U4006 ( .A1(n3288), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3146), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3125) );
  AOI22_X1 U4007 ( .A1(n3248), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3124) );
  AOI22_X1 U4008 ( .A1(n3309), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3290), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3123) );
  AOI22_X1 U4009 ( .A1(n3272), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3303), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3122) );
  NAND4_X1 U4010 ( .A1(n3125), .A2(n3124), .A3(n3123), .A4(n3122), .ZN(n3126)
         );
  OR2_X2 U4011 ( .A1(n3127), .A2(n3126), .ZN(n3379) );
  NOR2_X1 U4012 ( .A1(n4077), .A2(n4187), .ZN(n3128) );
  AND2_X1 U4013 ( .A1(n3128), .A2(n3222), .ZN(n3141) );
  INV_X1 U4014 ( .A(n3196), .ZN(n3129) );
  NAND2_X1 U4015 ( .A1(n3129), .A2(n4576), .ZN(n3139) );
  INV_X1 U4016 ( .A(n3190), .ZN(n3206) );
  NAND2_X1 U4017 ( .A1(n3206), .A2(n3189), .ZN(n3188) );
  AOI22_X1 U4018 ( .A1(n5124), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3133) );
  AOI22_X1 U4019 ( .A1(n3288), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3265), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3132) );
  AOI22_X1 U4020 ( .A1(n3249), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3131) );
  AOI22_X1 U4021 ( .A1(n3270), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3151), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3130) );
  AOI22_X1 U4022 ( .A1(n3243), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3138) );
  AOI22_X1 U4023 ( .A1(n3146), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3309), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3137) );
  AOI22_X1 U4024 ( .A1(n3248), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3134), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3136) );
  AOI22_X1 U4025 ( .A1(n3272), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3303), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3135) );
  NAND2_X2 U4026 ( .A1(n3045), .A2(n3048), .ZN(n5291) );
  NAND2_X2 U4027 ( .A1(n3139), .A2(n3051), .ZN(n4075) );
  INV_X1 U4028 ( .A(n4075), .ZN(n3140) );
  NAND2_X1 U4030 ( .A1(n3287), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3144) );
  NAND2_X1 U4031 ( .A1(n3265), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3143)
         );
  NAND2_X1 U4032 ( .A1(n3288), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3142) );
  NAND2_X1 U4033 ( .A1(n3243), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3150) );
  NAND2_X1 U4034 ( .A1(n3308), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U4035 ( .A1(n3271), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3148) );
  NAND2_X1 U4036 ( .A1(n3309), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3147) );
  AND4_X2 U4037 ( .A1(n3150), .A2(n3149), .A3(n3148), .A4(n3147), .ZN(n3163)
         );
  NAND2_X1 U4038 ( .A1(n3270), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3155) );
  NAND2_X1 U4039 ( .A1(n3272), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3154)
         );
  NAND2_X1 U4040 ( .A1(n3290), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3153) );
  NAND2_X1 U4041 ( .A1(n3303), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3152)
         );
  NAND2_X1 U4042 ( .A1(n3248), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3160)
         );
  NAND2_X1 U4043 ( .A1(n3249), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3159) );
  NAND2_X1 U4044 ( .A1(n3156), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3158) );
  NAND2_X1 U4045 ( .A1(n3250), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3157)
         );
  AND4_X2 U4046 ( .A1(n3160), .A2(n3159), .A3(n3158), .A4(n3157), .ZN(n3161)
         );
  NAND4_X4 U4047 ( .A1(n3164), .A2(n3163), .A3(n3162), .A4(n3161), .ZN(n4965)
         );
  NAND2_X1 U4048 ( .A1(n3941), .A2(n4965), .ZN(n4144) );
  NAND2_X1 U4049 ( .A1(n3028), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3168)
         );
  NAND2_X1 U4050 ( .A1(n3308), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3167) );
  NAND2_X1 U4051 ( .A1(n3243), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3166) );
  NAND2_X1 U4052 ( .A1(n3287), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3165) );
  NAND2_X1 U4053 ( .A1(n3248), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3172)
         );
  NAND2_X1 U4054 ( .A1(n3270), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3171) );
  NAND2_X1 U4055 ( .A1(n3249), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3170) );
  NAND2_X1 U4056 ( .A1(n3156), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3169) );
  NAND2_X1 U4058 ( .A1(n3288), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3176) );
  NAND2_X1 U4059 ( .A1(n3271), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3175) );
  NAND2_X1 U4060 ( .A1(n3265), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3174)
         );
  NAND2_X1 U4061 ( .A1(n3309), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3173) );
  AND4_X2 U4062 ( .A1(n3176), .A2(n3175), .A3(n3174), .A4(n3173), .ZN(n3182)
         );
  NAND2_X1 U4063 ( .A1(n3272), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3180)
         );
  NAND2_X1 U4064 ( .A1(n3290), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3179) );
  NAND2_X1 U4065 ( .A1(n3303), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3178)
         );
  NAND2_X1 U4066 ( .A1(n3250), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3177)
         );
  AND4_X2 U4067 ( .A1(n3180), .A2(n3179), .A3(n3178), .A4(n3177), .ZN(n3181)
         );
  INV_X1 U4068 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6504) );
  NOR2_X1 U4069 ( .A1(n6504), .A2(n6767), .ZN(n6505) );
  AOI21_X1 U4070 ( .B1(n6767), .B2(n6504), .A(n6505), .ZN(n3944) );
  INV_X1 U4071 ( .A(n3208), .ZN(n3200) );
  NOR2_X2 U4072 ( .A1(n4965), .A2(n3967), .ZN(n3969) );
  NOR2_X1 U4073 ( .A1(n4187), .A2(n4188), .ZN(n3185) );
  NAND2_X1 U4074 ( .A1(n5291), .A2(n3026), .ZN(n3946) );
  INV_X1 U4075 ( .A(n3969), .ZN(n4147) );
  NAND2_X2 U4076 ( .A1(n4576), .A2(n3187), .ZN(n6460) );
  NAND3_X1 U4077 ( .A1(n3215), .A2(n3188), .A3(n4576), .ZN(n3195) );
  INV_X2 U4078 ( .A(n4188), .ZN(n3194) );
  INV_X1 U4079 ( .A(n4576), .ZN(n3192) );
  OAI21_X1 U4080 ( .B1(n3195), .B2(n3194), .A(n3193), .ZN(n3198) );
  NAND2_X1 U4081 ( .A1(n3196), .A2(n3379), .ZN(n3220) );
  NAND2_X1 U4082 ( .A1(n3198), .A2(n3197), .ZN(n3204) );
  OAI211_X1 U4083 ( .C1(n4144), .C2(n3200), .A(n4073), .B(n4216), .ZN(n3201)
         );
  NAND2_X1 U4084 ( .A1(n3201), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3233) );
  INV_X1 U4085 ( .A(n3233), .ZN(n3203) );
  NAND2_X1 U4086 ( .A1(n6569), .A2(n6765), .ZN(n6583) );
  XNOR2_X1 U4087 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n5749) );
  OAI22_X1 U4088 ( .A1(n3926), .A2(n5749), .B1(n3555), .B2(n6445), .ZN(n3232)
         );
  OR2_X1 U4089 ( .A1(n3232), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3202)
         );
  NAND2_X1 U4090 ( .A1(n3203), .A2(n3202), .ZN(n3320) );
  NAND2_X1 U4091 ( .A1(n3204), .A2(n3969), .ZN(n4084) );
  INV_X2 U4092 ( .A(n3967), .ZN(n4402) );
  AOI21_X1 U4093 ( .B1(n3951), .B2(n4958), .A(n4086), .ZN(n3205) );
  NAND2_X1 U4094 ( .A1(n3208), .A2(n3207), .ZN(n3209) );
  NAND4_X1 U4095 ( .A1(n3209), .A2(n3222), .A3(n3391), .A4(n4076), .ZN(n3210)
         );
  NAND2_X1 U4096 ( .A1(n3227), .A2(n3211), .ZN(n3212) );
  NAND2_X1 U4097 ( .A1(n3212), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3230) );
  INV_X1 U4098 ( .A(n3555), .ZN(n4186) );
  INV_X1 U4099 ( .A(n3926), .ZN(n3241) );
  MUX2_X1 U4100 ( .A(n4186), .B(n3241), .S(n6256), .Z(n3213) );
  INV_X1 U4101 ( .A(n3213), .ZN(n3214) );
  OAI21_X2 U4102 ( .B1(n3230), .B2(n6438), .A(n3214), .ZN(n3264) );
  NOR2_X1 U4103 ( .A1(n3215), .A2(n3216), .ZN(n3552) );
  NOR2_X1 U4104 ( .A1(n3379), .A2(n4965), .ZN(n3217) );
  NAND2_X1 U4105 ( .A1(n3552), .A2(n3217), .ZN(n4431) );
  NAND2_X1 U4106 ( .A1(n4188), .A2(n3033), .ZN(n3218) );
  NOR2_X1 U4107 ( .A1(n6583), .A2(n6780), .ZN(n6485) );
  NAND2_X1 U4108 ( .A1(n3220), .A2(n4958), .ZN(n3221) );
  NAND2_X1 U4109 ( .A1(n3222), .A2(n3379), .ZN(n3223) );
  OAI21_X1 U4110 ( .B1(n4075), .B2(n3223), .A(n4968), .ZN(n3224) );
  INV_X1 U4111 ( .A(n4076), .ZN(n4952) );
  NAND2_X1 U4112 ( .A1(n4952), .A2(n6460), .ZN(n4081) );
  NAND3_X1 U4113 ( .A1(n3221), .A2(n3224), .A3(n4081), .ZN(n3225) );
  NAND2_X1 U4114 ( .A1(n3229), .A2(n3228), .ZN(n3262) );
  NAND2_X1 U4115 ( .A1(n3320), .A2(n3322), .ZN(n3235) );
  BUF_X2 U4116 ( .A(n3230), .Z(n3236) );
  INV_X1 U4117 ( .A(n3232), .ZN(n3234) );
  AND2_X1 U4118 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3238) );
  NAND2_X1 U4119 ( .A1(n3238), .A2(n6452), .ZN(n4728) );
  INV_X1 U4120 ( .A(n3238), .ZN(n3239) );
  NAND2_X1 U4121 ( .A1(n3239), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U4122 ( .A1(n4728), .A2(n3240), .ZN(n4380) );
  AOI22_X1 U4123 ( .A1(n3241), .A2(n4380), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n4186), .ZN(n3242) );
  NAND2_X1 U4124 ( .A1(n4375), .A2(n6780), .ZN(n3258) );
  INV_X1 U4125 ( .A(n3337), .ZN(n4192) );
  AOI22_X1 U4127 ( .A1(n5124), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3247) );
  AOI22_X1 U4128 ( .A1(n5145), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3246) );
  AOI22_X1 U4129 ( .A1(n5139), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3245) );
  BUF_X1 U4130 ( .A(n3309), .Z(n3289) );
  AOI22_X1 U4131 ( .A1(n5147), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3244) );
  NAND4_X1 U4132 ( .A1(n3247), .A2(n3246), .A3(n3245), .A4(n3244), .ZN(n3256)
         );
  AOI22_X1 U4133 ( .A1(n5138), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U4134 ( .A1(n3027), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3253) );
  AOI22_X1 U4136 ( .A1(n5146), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3291), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3252) );
  INV_X1 U4137 ( .A(n3250), .ZN(n4420) );
  AOI22_X1 U4138 ( .A1(n5149), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3251) );
  NAND4_X1 U4139 ( .A1(n3254), .A2(n3253), .A3(n3252), .A4(n3251), .ZN(n3255)
         );
  NAND2_X1 U4140 ( .A1(n4192), .A2(n3365), .ZN(n3257) );
  INV_X1 U4141 ( .A(n3336), .ZN(n3259) );
  INV_X1 U4143 ( .A(n3262), .ZN(n3263) );
  XNOR2_X1 U4144 ( .A(n3264), .B(n3263), .ZN(n3571) );
  AOI22_X1 U4145 ( .A1(n5145), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3028), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3269) );
  AOI22_X1 U4146 ( .A1(n5139), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5147), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3268) );
  AOI22_X1 U4147 ( .A1(n3248), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3267) );
  AOI22_X1 U4148 ( .A1(n5149), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3266) );
  NAND4_X1 U4149 ( .A1(n3269), .A2(n3268), .A3(n3267), .A4(n3266), .ZN(n3279)
         );
  AOI22_X1 U4150 ( .A1(n3281), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3277) );
  AOI22_X1 U4151 ( .A1(n5137), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3276) );
  AOI22_X1 U4152 ( .A1(n5100), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3275) );
  AOI22_X1 U4153 ( .A1(n5146), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3274) );
  NAND4_X1 U4154 ( .A1(n3277), .A2(n3276), .A3(n3275), .A4(n3274), .ZN(n3278)
         );
  INV_X1 U4155 ( .A(n3476), .ZN(n3280) );
  NOR2_X1 U4156 ( .A1(n3337), .A2(n3476), .ZN(n3316) );
  AOI22_X1 U4157 ( .A1(n5124), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3281), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4158 ( .A1(n5145), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4159 ( .A1(n3027), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3156), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4160 ( .A1(n5146), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5149), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3283) );
  NAND4_X1 U4161 ( .A1(n3286), .A2(n3285), .A3(n3284), .A4(n3283), .ZN(n3297)
         );
  AOI22_X1 U4162 ( .A1(n5138), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3295) );
  AOI22_X1 U4163 ( .A1(n3288), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3294) );
  AOI22_X1 U4164 ( .A1(n5147), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3293) );
  BUF_X1 U4165 ( .A(n3290), .Z(n3291) );
  AOI22_X1 U4166 ( .A1(n3291), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3292) );
  NAND4_X1 U4167 ( .A1(n3295), .A2(n3294), .A3(n3293), .A4(n3292), .ZN(n3296)
         );
  MUX2_X1 U4168 ( .A(n3477), .B(n3316), .S(n3403), .Z(n3398) );
  INV_X1 U4169 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4413) );
  AOI21_X1 U4170 ( .B1(n3298), .B2(n3476), .A(n6780), .ZN(n3301) );
  NAND2_X1 U4171 ( .A1(n4409), .A2(n3403), .ZN(n3300) );
  OAI211_X1 U4172 ( .C1(n3536), .C2(n4413), .A(n3301), .B(n3300), .ZN(n3396)
         );
  AOI21_X1 U4173 ( .B1(n3398), .B2(n3396), .A(n3477), .ZN(n3302) );
  AOI22_X1 U4174 ( .A1(n5145), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n5124), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3307) );
  AOI22_X1 U4175 ( .A1(n5138), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3306) );
  AOI22_X1 U4176 ( .A1(n5139), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5147), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3305) );
  AOI22_X1 U4177 ( .A1(n3291), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n5149), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3304) );
  NAND4_X1 U4178 ( .A1(n3307), .A2(n3306), .A3(n3305), .A4(n3304), .ZN(n3315)
         );
  AOI22_X1 U4179 ( .A1(n5136), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3313) );
  AOI22_X1 U4180 ( .A1(n3027), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3312) );
  BUF_X1 U4181 ( .A(n3309), .Z(n5083) );
  AOI22_X1 U4182 ( .A1(n5100), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4183 ( .A1(n5146), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3310) );
  NAND4_X1 U4184 ( .A1(n3313), .A2(n3312), .A3(n3311), .A4(n3310), .ZN(n3314)
         );
  INV_X1 U4185 ( .A(n3390), .ZN(n3319) );
  INV_X1 U4186 ( .A(n3316), .ZN(n3318) );
  NAND2_X1 U4187 ( .A1(n3544), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3317) );
  OAI211_X1 U4188 ( .C1(n3319), .C2(n3336), .A(n3318), .B(n3317), .ZN(n3383)
         );
  NAND2_X1 U4189 ( .A1(n3321), .A2(n3320), .ZN(n3324) );
  NAND2_X1 U4190 ( .A1(n4192), .A2(n3390), .ZN(n3325) );
  OAI21_X1 U4191 ( .B1(n3385), .B2(n3383), .A(n3386), .ZN(n3327) );
  NAND2_X1 U4192 ( .A1(n3385), .A2(n3383), .ZN(n3326) );
  NAND2_X1 U4193 ( .A1(n3327), .A2(n3326), .ZN(n3371) );
  INV_X1 U4194 ( .A(n3373), .ZN(n3350) );
  INV_X1 U4195 ( .A(n3236), .ZN(n3331) );
  NAND2_X1 U4196 ( .A1(n3331), .A2(n6575), .ZN(n3335) );
  NOR3_X1 U4197 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6452), .A3(n6445), 
        .ZN(n6341) );
  NAND2_X1 U4198 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6341), .ZN(n6338) );
  NAND2_X1 U4199 ( .A1(n6458), .A2(n6338), .ZN(n3332) );
  NAND3_X1 U4200 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n4638) );
  INV_X1 U4201 ( .A(n4638), .ZN(n4463) );
  NAND2_X1 U4202 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4463), .ZN(n4804) );
  NAND2_X1 U4203 ( .A1(n3332), .A2(n4804), .ZN(n4369) );
  OAI22_X1 U4204 ( .A1(n3926), .A2(n4369), .B1(n3555), .B2(n6458), .ZN(n3333)
         );
  INV_X1 U4205 ( .A(n3333), .ZN(n3334) );
  AOI22_X1 U4206 ( .A1(n5124), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3341) );
  AOI22_X1 U4207 ( .A1(n5145), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4208 ( .A1(n5139), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4209 ( .A1(n5147), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3338) );
  NAND4_X1 U4210 ( .A1(n3341), .A2(n3340), .A3(n3339), .A4(n3338), .ZN(n3347)
         );
  AOI22_X1 U4211 ( .A1(n5138), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3345) );
  AOI22_X1 U4212 ( .A1(n3027), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3344) );
  AOI22_X1 U4213 ( .A1(n5146), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3291), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3343) );
  AOI22_X1 U4214 ( .A1(n5149), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3342) );
  NAND4_X1 U4215 ( .A1(n3345), .A2(n3344), .A3(n3343), .A4(n3342), .ZN(n3346)
         );
  AOI22_X1 U4216 ( .A1(n3548), .A2(n3369), .B1(n3544), .B2(
        INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3348) );
  INV_X1 U4217 ( .A(n4506), .ZN(n4542) );
  INV_X1 U4218 ( .A(n3433), .ZN(n3363) );
  AOI22_X1 U4219 ( .A1(n5105), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3354) );
  AOI22_X1 U4220 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n5138), .B1(n5148), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4221 ( .A1(n5139), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3291), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4222 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n5146), .B1(n5149), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3351) );
  NAND4_X1 U4223 ( .A1(n3354), .A2(n3353), .A3(n3352), .A4(n3351), .ZN(n3360)
         );
  AOI22_X1 U4224 ( .A1(n5145), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3028), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4225 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n5137), .B1(n3027), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4226 ( .A1(n5144), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3356) );
  AOI22_X1 U4227 ( .A1(n5147), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3355) );
  NAND4_X1 U4228 ( .A1(n3358), .A2(n3357), .A3(n3356), .A4(n3355), .ZN(n3359)
         );
  NAND2_X1 U4229 ( .A1(n3548), .A2(n3438), .ZN(n3362) );
  NAND2_X1 U4230 ( .A1(n3544), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3361) );
  NAND2_X1 U4231 ( .A1(n3363), .A2(n3431), .ZN(n3436) );
  NAND2_X1 U4232 ( .A1(n3436), .A2(n3364), .ZN(n3591) );
  NAND2_X1 U4233 ( .A1(n4968), .A2(n4187), .ZN(n3950) );
  NAND2_X1 U4234 ( .A1(n3390), .A2(n3403), .ZN(n3389) );
  INV_X1 U4235 ( .A(n3365), .ZN(n3378) );
  NAND2_X1 U4236 ( .A1(n3389), .A2(n3378), .ZN(n3377) );
  NAND2_X1 U4237 ( .A1(n3377), .A2(n3369), .ZN(n3440) );
  XOR2_X1 U4238 ( .A(n3438), .B(n3440), .Z(n3366) );
  INV_X1 U4239 ( .A(n4958), .ZN(n6599) );
  OAI21_X1 U4240 ( .B1(n3591), .B2(n3950), .A(n3049), .ZN(n3415) );
  XNOR2_X1 U4241 ( .A(n3415), .B(n3367), .ZN(n5049) );
  NAND2_X1 U4242 ( .A1(n3373), .A2(n4506), .ZN(n3368) );
  NAND2_X1 U4243 ( .A1(n3433), .A2(n3368), .ZN(n3580) );
  OAI211_X1 U4244 ( .C1(n3369), .C2(n3377), .A(n3440), .B(n4958), .ZN(n3370)
         );
  OAI21_X2 U4245 ( .B1(n3580), .B2(n3950), .A(n3370), .ZN(n3413) );
  NAND2_X1 U4246 ( .A1(n3374), .A2(n3373), .ZN(n3557) );
  INV_X1 U4247 ( .A(n3950), .ZN(n3375) );
  OAI21_X1 U4248 ( .B1(n3378), .B2(n3389), .A(n3377), .ZN(n3380) );
  AND2_X1 U4249 ( .A1(n4409), .A2(n3379), .ZN(n3401) );
  AOI21_X1 U4250 ( .B1(n3380), .B2(n4958), .A(n3401), .ZN(n3381) );
  NAND2_X1 U4251 ( .A1(n3382), .A2(n3381), .ZN(n3409) );
  NAND2_X1 U4252 ( .A1(n3409), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6177)
         );
  INV_X1 U4253 ( .A(n3383), .ZN(n3384) );
  XNOR2_X1 U4254 ( .A(n3385), .B(n3384), .ZN(n3388) );
  INV_X1 U4255 ( .A(n3386), .ZN(n3387) );
  XNOR2_X1 U4256 ( .A(n3388), .B(n3387), .ZN(n3563) );
  NAND2_X1 U4257 ( .A1(n3563), .A2(n3375), .ZN(n3395) );
  OAI21_X1 U4258 ( .B1(n3403), .B2(n3390), .A(n3389), .ZN(n3392) );
  OAI211_X1 U4259 ( .C1(n3392), .C2(n6599), .A(n3391), .B(n4187), .ZN(n3393)
         );
  INV_X1 U4260 ( .A(n3393), .ZN(n3394) );
  NAND2_X1 U4261 ( .A1(n3395), .A2(n3394), .ZN(n4277) );
  INV_X1 U4262 ( .A(n3396), .ZN(n3397) );
  XNOR2_X1 U4263 ( .A(n3398), .B(n3397), .ZN(n3399) );
  OR2_X1 U4264 ( .A1(n3569), .A2(n3950), .ZN(n3406) );
  INV_X1 U4265 ( .A(n3401), .ZN(n3402) );
  OAI21_X1 U4266 ( .B1(n6599), .B2(n3403), .A(n3402), .ZN(n3404) );
  INV_X1 U4267 ( .A(n3404), .ZN(n3405) );
  NAND2_X1 U4268 ( .A1(n3406), .A2(n3405), .ZN(n6189) );
  NAND2_X1 U4269 ( .A1(n4277), .A2(n4276), .ZN(n4275) );
  INV_X1 U4270 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6246) );
  OR2_X1 U4271 ( .A1(n6193), .A2(n6246), .ZN(n3407) );
  NAND2_X1 U4272 ( .A1(n4275), .A2(n3407), .ZN(n6181) );
  INV_X1 U4273 ( .A(n6181), .ZN(n3408) );
  NAND2_X1 U4274 ( .A1(n6177), .A2(n3408), .ZN(n3412) );
  INV_X1 U4275 ( .A(n3409), .ZN(n3411) );
  NAND2_X1 U4276 ( .A1(n3411), .A2(n3410), .ZN(n6176) );
  INV_X1 U4277 ( .A(n3413), .ZN(n3414) );
  NAND2_X1 U4278 ( .A1(n5049), .A2(n5050), .ZN(n3417) );
  NAND2_X1 U4279 ( .A1(n3415), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3416)
         );
  AND2_X2 U4280 ( .A1(n3417), .A2(n3416), .ZN(n4688) );
  AOI22_X1 U4281 ( .A1(n5124), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3421) );
  AOI22_X1 U4282 ( .A1(n5145), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3420) );
  AOI22_X1 U4283 ( .A1(n5139), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3419) );
  AOI22_X1 U4284 ( .A1(n5147), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3418) );
  NAND4_X1 U4285 ( .A1(n3421), .A2(n3420), .A3(n3419), .A4(n3418), .ZN(n3427)
         );
  AOI22_X1 U4286 ( .A1(n5138), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4287 ( .A1(n3027), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3424) );
  AOI22_X1 U4288 ( .A1(n5146), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3291), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3423) );
  AOI22_X1 U4289 ( .A1(n5149), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3422) );
  NAND4_X1 U4290 ( .A1(n3425), .A2(n3424), .A3(n3423), .A4(n3422), .ZN(n3426)
         );
  NAND2_X1 U4291 ( .A1(n3548), .A2(n3441), .ZN(n3429) );
  NAND2_X1 U4292 ( .A1(n3544), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3428) );
  NAND2_X1 U4293 ( .A1(n3429), .A2(n3428), .ZN(n3434) );
  INV_X1 U4294 ( .A(n3434), .ZN(n3435) );
  NAND2_X1 U4295 ( .A1(n3436), .A2(n3435), .ZN(n3437) );
  NAND2_X1 U4296 ( .A1(n3462), .A2(n3437), .ZN(n3601) );
  INV_X1 U4297 ( .A(n3438), .ZN(n3439) );
  NOR2_X1 U4298 ( .A1(n3440), .A2(n3439), .ZN(n3442) );
  NAND2_X1 U4299 ( .A1(n3442), .A2(n3441), .ZN(n3468) );
  OAI211_X1 U4300 ( .C1(n3442), .C2(n3441), .A(n3468), .B(n4958), .ZN(n3443)
         );
  XNOR2_X1 U4301 ( .A(n3444), .B(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4689)
         );
  INV_X1 U4302 ( .A(n3444), .ZN(n3446) );
  INV_X1 U4303 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3445) );
  OAI22_X2 U4304 ( .A1(n4688), .A2(n4689), .B1(n3446), .B2(n3445), .ZN(n4532)
         );
  AOI22_X1 U4305 ( .A1(n3028), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4306 ( .A1(n5138), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4307 ( .A1(n5139), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3448) );
  AOI22_X1 U4308 ( .A1(n5137), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3291), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3447) );
  NAND4_X1 U4309 ( .A1(n3450), .A2(n3449), .A3(n3448), .A4(n3447), .ZN(n3456)
         );
  AOI22_X1 U4310 ( .A1(n5145), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4311 ( .A1(n5144), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5147), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3453) );
  AOI22_X1 U4312 ( .A1(n5146), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5149), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3452) );
  AOI22_X1 U4313 ( .A1(n3027), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3451) );
  NAND4_X1 U4314 ( .A1(n3454), .A2(n3453), .A3(n3452), .A4(n3451), .ZN(n3455)
         );
  OR2_X1 U4315 ( .A1(n3456), .A2(n3455), .ZN(n3469) );
  NAND2_X1 U4316 ( .A1(n3548), .A2(n3469), .ZN(n3458) );
  NAND2_X1 U4317 ( .A1(n3544), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3457) );
  NAND2_X1 U4318 ( .A1(n3458), .A2(n3457), .ZN(n3460) );
  INV_X1 U4319 ( .A(n3460), .ZN(n3461) );
  NAND3_X1 U4320 ( .A1(n3480), .A2(n3614), .A3(n3375), .ZN(n3464) );
  XOR2_X1 U4321 ( .A(n3469), .B(n3468), .Z(n3463) );
  NAND2_X1 U4322 ( .A1(n3464), .A2(n3050), .ZN(n3465) );
  XOR2_X1 U4323 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .B(n3465), .Z(n4531) );
  INV_X1 U4324 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4399) );
  NAND2_X1 U4325 ( .A1(n3548), .A2(n3476), .ZN(n3466) );
  OAI21_X1 U4326 ( .B1(n4399), .B2(n3536), .A(n3466), .ZN(n3467) );
  NAND2_X1 U4327 ( .A1(n3617), .A2(n3375), .ZN(n3473) );
  INV_X1 U4328 ( .A(n3468), .ZN(n3470) );
  NAND2_X1 U4329 ( .A1(n3470), .A2(n3469), .ZN(n3482) );
  XNOR2_X1 U4330 ( .A(n3482), .B(n3476), .ZN(n3471) );
  NAND2_X1 U4331 ( .A1(n3471), .A2(n4958), .ZN(n3472) );
  NAND2_X1 U4332 ( .A1(n3473), .A2(n3472), .ZN(n3474) );
  XNOR2_X1 U4333 ( .A(n3474), .B(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4933)
         );
  NAND2_X1 U4334 ( .A1(n3474), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3475)
         );
  NAND2_X1 U4335 ( .A1(n4958), .A2(n3476), .ZN(n3481) );
  INV_X1 U4336 ( .A(n3477), .ZN(n3478) );
  NOR2_X1 U4337 ( .A1(n3478), .A2(n3950), .ZN(n3479) );
  OAI21_X1 U4338 ( .B1(n3482), .B2(n3481), .A(n3488), .ZN(n3483) );
  XOR2_X1 U4339 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .B(n3483), .Z(n4910) );
  INV_X1 U4340 ( .A(n3483), .ZN(n3484) );
  NAND2_X1 U4341 ( .A1(n3500), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3487)
         );
  INV_X1 U4342 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6234) );
  AOI21_X2 U4343 ( .B1(n4997), .B2(n3487), .A(n3486), .ZN(n4978) );
  INV_X1 U4344 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U4345 ( .A1(n5890), .A2(n6224), .ZN(n4979) );
  NAND2_X1 U4346 ( .A1(n3500), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6154) );
  INV_X1 U4347 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5240) );
  NAND2_X1 U4348 ( .A1(n5890), .A2(n5240), .ZN(n3489) );
  AOI21_X1 U4349 ( .B1(n5017), .B2(n3489), .A(n3037), .ZN(n5635) );
  NAND2_X1 U4350 ( .A1(n5635), .A2(n5638), .ZN(n5636) );
  NAND2_X1 U4351 ( .A1(n5636), .A2(n3036), .ZN(n5238) );
  NAND2_X1 U4352 ( .A1(n3500), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3490) );
  INV_X1 U4353 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5721) );
  AOI21_X2 U4354 ( .B1(n5238), .B2(n3490), .A(n3039), .ZN(n5613) );
  OAI21_X2 U4355 ( .B1(n5613), .B2(n5629), .A(n3492), .ZN(n5612) );
  INV_X1 U4356 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5617) );
  INV_X1 U4357 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5913) );
  NAND2_X1 U4358 ( .A1(n5617), .A2(n5913), .ZN(n3493) );
  OAI21_X1 U4359 ( .B1(INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n3493), .A(n3500), 
        .ZN(n3496) );
  NAND3_X1 U4360 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .A3(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n3494) );
  AOI21_X2 U4361 ( .B1(n5612), .B2(n3496), .A(n3495), .ZN(n5698) );
  INV_X1 U4362 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5705) );
  XNOR2_X1 U4363 ( .A(n5890), .B(n5705), .ZN(n5697) );
  NOR2_X1 U4364 ( .A1(n5696), .A2(n3497), .ZN(n5605) );
  NAND2_X1 U4365 ( .A1(n5605), .A2(n3040), .ZN(n3499) );
  NAND2_X1 U4366 ( .A1(n3499), .A2(n3498), .ZN(n4133) );
  XNOR2_X1 U4367 ( .A(n3500), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4132)
         );
  INV_X1 U4368 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3501) );
  NAND2_X1 U4369 ( .A1(n5890), .A2(n3501), .ZN(n3502) );
  NAND3_X1 U4370 ( .A1(n5890), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3504) );
  NOR2_X1 U4371 ( .A1(n5890), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5595)
         );
  NAND2_X1 U4372 ( .A1(n3503), .A2(n5595), .ZN(n4119) );
  XNOR2_X1 U4373 ( .A(n3505), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5226)
         );
  NAND2_X1 U4374 ( .A1(n6445), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3508) );
  NAND2_X1 U4375 ( .A1(n3231), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3506) );
  NAND2_X1 U4376 ( .A1(n3508), .A2(n3506), .ZN(n3520) );
  NAND2_X1 U4377 ( .A1(n3507), .A2(n6256), .ZN(n3519) );
  OAI21_X1 U4378 ( .B1(n3520), .B2(n3519), .A(n3508), .ZN(n3535) );
  NAND2_X1 U4379 ( .A1(n6452), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3510) );
  NAND2_X1 U4380 ( .A1(n3237), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3509) );
  NAND2_X1 U4381 ( .A1(n3510), .A2(n3509), .ZN(n3534) );
  INV_X1 U4382 ( .A(n3534), .ZN(n3512) );
  INV_X1 U4383 ( .A(n3510), .ZN(n3511) );
  XNOR2_X1 U4384 ( .A(n3585), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3517)
         );
  INV_X1 U4385 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5946) );
  INV_X1 U4386 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6456) );
  NOR2_X1 U4387 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n6456), .ZN(n3513)
         );
  AOI221_X1 U4388 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n3514), .C1(
        n5946), .C2(n3514), .A(n3513), .ZN(n3958) );
  NAND2_X1 U4389 ( .A1(n3958), .A2(n3533), .ZN(n3551) );
  AND3_X1 U4390 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3514), .A3(n5946), 
        .ZN(n3515) );
  AOI211_X1 U4391 ( .C1(n3518), .C2(n3517), .A(n3516), .B(n3515), .ZN(n3543)
         );
  INV_X1 U4392 ( .A(n3543), .ZN(n3961) );
  AOI22_X1 U4393 ( .A1(n3533), .A2(n3961), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6780), .ZN(n3546) );
  INV_X1 U4394 ( .A(n3519), .ZN(n3521) );
  XNOR2_X1 U4395 ( .A(n3520), .B(n3521), .ZN(n3956) );
  AOI21_X1 U4396 ( .B1(n3207), .B2(n4965), .A(n4968), .ZN(n3538) );
  AOI21_X1 U4397 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6438), .A(n3521), 
        .ZN(n3526) );
  AOI21_X1 U4398 ( .B1(n3526), .B2(n6460), .A(n4409), .ZN(n3523) );
  AND2_X1 U4399 ( .A1(n3956), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3525) );
  NAND2_X1 U4400 ( .A1(n3548), .A2(n4968), .ZN(n3522) );
  NAND2_X1 U4401 ( .A1(n3522), .A2(n4187), .ZN(n3524) );
  OAI22_X1 U4402 ( .A1(n3538), .A2(n3523), .B1(n3525), .B2(n3524), .ZN(n3527)
         );
  NAND2_X1 U4403 ( .A1(n3956), .A2(n3527), .ZN(n3532) );
  INV_X1 U4404 ( .A(n3524), .ZN(n3530) );
  INV_X1 U4405 ( .A(n3525), .ZN(n3529) );
  NAND2_X1 U4406 ( .A1(n3526), .A2(n3548), .ZN(n3528) );
  OAI22_X1 U4407 ( .A1(n3530), .A2(n3529), .B1(n3528), .B2(n3527), .ZN(n3531)
         );
  AOI21_X1 U4408 ( .B1(n3533), .B2(n3532), .A(n3531), .ZN(n3541) );
  XNOR2_X1 U4409 ( .A(n3535), .B(n3534), .ZN(n3957) );
  NOR2_X1 U4410 ( .A1(n3536), .A2(n3957), .ZN(n3537) );
  AOI211_X1 U4411 ( .C1(n3548), .C2(n3957), .A(n3537), .B(n3538), .ZN(n3540)
         );
  NAND3_X1 U4412 ( .A1(n3538), .A2(n3548), .A3(n3957), .ZN(n3539) );
  OAI21_X1 U4413 ( .B1(n3541), .B2(n3540), .A(n3539), .ZN(n3542) );
  OAI21_X1 U4414 ( .B1(n3544), .B2(n3543), .A(n3542), .ZN(n3545) );
  NAND2_X1 U4415 ( .A1(n3546), .A2(n3545), .ZN(n3547) );
  NOR2_X1 U4416 ( .A1(n4075), .A2(n4384), .ZN(n3554) );
  NAND2_X1 U4417 ( .A1(n3552), .A2(n4187), .ZN(n6437) );
  NAND2_X1 U4418 ( .A1(n3194), .A2(n3033), .ZN(n4087) );
  NAND2_X1 U4419 ( .A1(n6437), .A2(n4087), .ZN(n3553) );
  NAND2_X1 U4420 ( .A1(n3554), .A2(n3553), .ZN(n6461) );
  AND2_X1 U4421 ( .A1(n3555), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6484) );
  INV_X1 U4422 ( .A(n6484), .ZN(n6482) );
  OR2_X1 U4423 ( .A1(n6460), .A2(n6482), .ZN(n3556) );
  NAND2_X1 U4424 ( .A1(n3559), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3724) );
  NAND2_X1 U4425 ( .A1(n6486), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3912) );
  NAND2_X1 U4426 ( .A1(n3186), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3593) );
  OAI21_X1 U4427 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3581), .ZN(n6187) );
  NOR2_X2 U4428 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n5205) );
  INV_X1 U4429 ( .A(n3912), .ZN(n5275) );
  AOI22_X1 U4430 ( .A1(n6187), .A2(n5205), .B1(n5275), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3562) );
  NOR2_X2 U4431 ( .A1(n5291), .A2(n6486), .ZN(n3888) );
  NAND2_X1 U4432 ( .A1(n5276), .A2(EAX_REG_2__SCAN_IN), .ZN(n3561) );
  OAI211_X1 U4433 ( .C1(n3593), .C2(n3237), .A(n3562), .B(n3561), .ZN(n3588)
         );
  NAND2_X1 U4434 ( .A1(n3589), .A2(n3588), .ZN(n3579) );
  NAND2_X1 U4435 ( .A1(n5744), .A2(n3739), .ZN(n3568) );
  NAND2_X1 U4436 ( .A1(n3888), .A2(EAX_REG_1__SCAN_IN), .ZN(n3565) );
  NAND2_X1 U4437 ( .A1(n6486), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3564)
         );
  OAI211_X1 U4438 ( .C1(n3593), .C2(n3231), .A(n3565), .B(n3564), .ZN(n3566)
         );
  INV_X1 U4439 ( .A(n3566), .ZN(n3567) );
  NAND2_X1 U4440 ( .A1(n3568), .A2(n3567), .ZN(n4280) );
  INV_X1 U4441 ( .A(n3215), .ZN(n3570) );
  NAND2_X1 U4442 ( .A1(n3032), .A2(n3570), .ZN(n4182) );
  NAND2_X1 U4443 ( .A1(n6441), .A2(n3739), .ZN(n3576) );
  NAND2_X1 U4444 ( .A1(n6486), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3573)
         );
  NAND2_X1 U4445 ( .A1(n3888), .A2(EAX_REG_0__SCAN_IN), .ZN(n3572) );
  OAI211_X1 U4446 ( .C1(n3593), .C2(n6438), .A(n3573), .B(n3572), .ZN(n3574)
         );
  INV_X1 U4447 ( .A(n3574), .ZN(n3575) );
  NAND2_X1 U4448 ( .A1(n3576), .A2(n3575), .ZN(n4184) );
  AND2_X1 U4449 ( .A1(n4184), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3577) );
  NAND2_X1 U4450 ( .A1(n4182), .A2(n3577), .ZN(n4183) );
  INV_X1 U4451 ( .A(n5205), .ZN(n5211) );
  OR2_X1 U4452 ( .A1(n4184), .A2(n5211), .ZN(n3578) );
  NAND2_X1 U4453 ( .A1(n4183), .A2(n3578), .ZN(n4279) );
  NAND2_X1 U4454 ( .A1(n4280), .A2(n4279), .ZN(n4278) );
  NAND2_X1 U4455 ( .A1(n3579), .A2(n4278), .ZN(n4270) );
  INV_X1 U4456 ( .A(n5742), .ZN(n3587) );
  AOI21_X1 U4457 ( .B1(n3581), .B2(n4359), .A(n3595), .ZN(n5478) );
  OAI22_X1 U4458 ( .A1(n5478), .A2(n5211), .B1(n3912), .B2(n4359), .ZN(n3582)
         );
  INV_X1 U4459 ( .A(n3582), .ZN(n3584) );
  NAND2_X1 U4460 ( .A1(n3888), .A2(EAX_REG_3__SCAN_IN), .ZN(n3583) );
  OAI211_X1 U4461 ( .C1(n3593), .C2(n3585), .A(n3584), .B(n3583), .ZN(n3586)
         );
  AOI21_X1 U4462 ( .B1(n3587), .B2(n3739), .A(n3586), .ZN(n4354) );
  INV_X1 U4463 ( .A(n4354), .ZN(n3590) );
  INV_X1 U4464 ( .A(n3591), .ZN(n3600) );
  INV_X1 U4465 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6068) );
  AOI21_X1 U4466 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n6068), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3592) );
  AOI21_X1 U4467 ( .B1(n3888), .B2(EAX_REG_4__SCAN_IN), .A(n3592), .ZN(n3598)
         );
  INV_X1 U4468 ( .A(n3593), .ZN(n3594) );
  NAND2_X1 U4469 ( .A1(n3594), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3597) );
  OAI21_X1 U4470 ( .B1(n3595), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3602), 
        .ZN(n6071) );
  NOR2_X1 U4471 ( .A1(n6071), .A2(n5211), .ZN(n3596) );
  AOI21_X1 U4472 ( .B1(n3598), .B2(n3597), .A(n3596), .ZN(n3599) );
  NAND2_X1 U4473 ( .A1(n3602), .A2(n6175), .ZN(n3604) );
  INV_X1 U4474 ( .A(n3609), .ZN(n3603) );
  NAND2_X1 U4475 ( .A1(n3604), .A2(n3603), .ZN(n6052) );
  NAND2_X1 U4476 ( .A1(n6052), .A2(n5205), .ZN(n3605) );
  OAI21_X1 U4477 ( .B1(n6175), .B2(n3912), .A(n3605), .ZN(n3606) );
  AOI21_X1 U4478 ( .B1(n3888), .B2(EAX_REG_5__SCAN_IN), .A(n3606), .ZN(n3607)
         );
  NAND2_X1 U4479 ( .A1(n4348), .A2(n4347), .ZN(n4678) );
  NAND2_X1 U4480 ( .A1(n3888), .A2(EAX_REG_6__SCAN_IN), .ZN(n3612) );
  INV_X1 U4481 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6487) );
  OAI21_X1 U4482 ( .B1(n6487), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6486), 
        .ZN(n3611) );
  OAI21_X1 U4483 ( .B1(n3609), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n3618), 
        .ZN(n6038) );
  INV_X1 U4484 ( .A(n6038), .ZN(n3610) );
  AOI22_X1 U4485 ( .A1(n3612), .A2(n3611), .B1(n3610), .B2(n5205), .ZN(n3613)
         );
  AOI21_X1 U4486 ( .B1(n6167), .B2(n3618), .A(n3636), .ZN(n3619) );
  INV_X1 U4487 ( .A(n3619), .ZN(n6161) );
  NAND2_X1 U4488 ( .A1(n6161), .A2(n5205), .ZN(n3621) );
  AOI22_X1 U4489 ( .A1(n5276), .A2(EAX_REG_7__SCAN_IN), .B1(n5275), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3620) );
  NAND2_X1 U4490 ( .A1(n3621), .A2(n3620), .ZN(n3622) );
  AOI22_X1 U4491 ( .A1(n3734), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3626) );
  AOI22_X1 U4492 ( .A1(n5138), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3625) );
  AOI22_X1 U4493 ( .A1(n5147), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3624) );
  AOI22_X1 U4494 ( .A1(n5137), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3623) );
  NAND4_X1 U4495 ( .A1(n3626), .A2(n3625), .A3(n3624), .A4(n3623), .ZN(n3632)
         );
  AOI22_X1 U4496 ( .A1(n5145), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4497 ( .A1(n5139), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4498 ( .A1(n5146), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3291), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3628) );
  AOI22_X1 U4499 ( .A1(n5148), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5149), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3627) );
  NAND4_X1 U4500 ( .A1(n3630), .A2(n3629), .A3(n3628), .A4(n3627), .ZN(n3631)
         );
  NOR2_X1 U4501 ( .A1(n3632), .A2(n3631), .ZN(n3635) );
  XNOR2_X1 U4502 ( .A(n3636), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n5467) );
  NAND2_X1 U4503 ( .A1(n5467), .A2(n5205), .ZN(n3634) );
  AOI22_X1 U4504 ( .A1(n5276), .A2(EAX_REG_8__SCAN_IN), .B1(n5275), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3633) );
  OAI211_X1 U4505 ( .C1(n3635), .C2(n3724), .A(n3634), .B(n3633), .ZN(n4787)
         );
  INV_X1 U4506 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6006) );
  XOR2_X1 U4507 ( .A(n6006), .B(n3649), .Z(n6011) );
  AOI22_X1 U4508 ( .A1(n5276), .A2(EAX_REG_9__SCAN_IN), .B1(n5275), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4509 ( .A1(n5145), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4510 ( .A1(n3027), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4511 ( .A1(n5100), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3638) );
  AOI22_X1 U4512 ( .A1(n5146), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3291), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3637) );
  NAND4_X1 U4513 ( .A1(n3640), .A2(n3639), .A3(n3638), .A4(n3637), .ZN(n3646)
         );
  AOI22_X1 U4514 ( .A1(n3734), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3644) );
  AOI22_X1 U4515 ( .A1(n5138), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3643) );
  AOI22_X1 U4516 ( .A1(n5139), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5147), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3642) );
  AOI22_X1 U4517 ( .A1(n5149), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3641) );
  NAND4_X1 U4518 ( .A1(n3644), .A2(n3643), .A3(n3642), .A4(n3641), .ZN(n3645)
         );
  OAI21_X1 U4519 ( .B1(n3646), .B2(n3645), .A(n3739), .ZN(n3647) );
  OAI211_X1 U4520 ( .C1(n6011), .C2(n5211), .A(n3648), .B(n3647), .ZN(n4921)
         );
  XNOR2_X1 U4521 ( .A(n3666), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5456)
         );
  AOI22_X1 U4522 ( .A1(n3734), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3653) );
  AOI22_X1 U4523 ( .A1(n5139), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3652) );
  AOI22_X1 U4524 ( .A1(n5147), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n5146), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3651) );
  AOI22_X1 U4525 ( .A1(n5137), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3650) );
  NAND4_X1 U4526 ( .A1(n3653), .A2(n3652), .A3(n3651), .A4(n3650), .ZN(n3659)
         );
  AOI22_X1 U4527 ( .A1(n5145), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3657) );
  AOI22_X1 U4528 ( .A1(n5138), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4529 ( .A1(n5083), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3291), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3655) );
  AOI22_X1 U4530 ( .A1(n5149), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3654) );
  NAND4_X1 U4531 ( .A1(n3657), .A2(n3656), .A3(n3655), .A4(n3654), .ZN(n3658)
         );
  NOR2_X1 U4532 ( .A1(n3659), .A2(n3658), .ZN(n3662) );
  NAND2_X1 U4533 ( .A1(n5276), .A2(EAX_REG_10__SCAN_IN), .ZN(n3661) );
  NAND2_X1 U4534 ( .A1(n5275), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3660)
         );
  OAI211_X1 U4535 ( .C1(n3724), .C2(n3662), .A(n3661), .B(n3660), .ZN(n3663)
         );
  AOI21_X1 U4536 ( .B1(n5456), .B2(n5205), .A(n3663), .ZN(n4942) );
  INV_X1 U4537 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n5996) );
  XOR2_X1 U4538 ( .A(n5996), .B(n3681), .Z(n6157) );
  AOI22_X1 U4539 ( .A1(n5276), .A2(EAX_REG_11__SCAN_IN), .B1(n5275), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3678) );
  AOI22_X1 U4540 ( .A1(n5145), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4541 ( .A1(n5138), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3669) );
  AOI22_X1 U4542 ( .A1(n5144), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4543 ( .A1(n5146), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3667) );
  NAND4_X1 U4544 ( .A1(n3670), .A2(n3669), .A3(n3668), .A4(n3667), .ZN(n3676)
         );
  AOI22_X1 U4545 ( .A1(n3734), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3674) );
  AOI22_X1 U4546 ( .A1(n5139), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n5147), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3673) );
  AOI22_X1 U4547 ( .A1(n5137), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4548 ( .A1(n3291), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5149), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3671) );
  NAND4_X1 U4549 ( .A1(n3674), .A2(n3673), .A3(n3672), .A4(n3671), .ZN(n3675)
         );
  OAI21_X1 U4550 ( .B1(n3676), .B2(n3675), .A(n3739), .ZN(n3677) );
  OAI211_X1 U4551 ( .C1(n6157), .C2(n5211), .A(n3678), .B(n3677), .ZN(n3679)
         );
  INV_X1 U4552 ( .A(n3679), .ZN(n4991) );
  XNOR2_X1 U4553 ( .A(n3697), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5445)
         );
  INV_X1 U4554 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5012) );
  INV_X1 U4555 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3682) );
  OAI22_X1 U4556 ( .A1(n3916), .A2(n5012), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3682), .ZN(n3683) );
  NAND2_X1 U4557 ( .A1(n3683), .A2(n5211), .ZN(n3695) );
  AOI22_X1 U4558 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n5139), .B1(n3734), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4559 ( .A1(n5147), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4560 ( .A1(n5146), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4561 ( .A1(n5138), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5149), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3684) );
  NAND4_X1 U4562 ( .A1(n3687), .A2(n3686), .A3(n3685), .A4(n3684), .ZN(n3693)
         );
  AOI22_X1 U4563 ( .A1(n5145), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4564 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n5144), .B1(n5100), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4565 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5148), .B1(n3027), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4566 ( .A1(n5137), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3688) );
  NAND4_X1 U4567 ( .A1(n3691), .A2(n3690), .A3(n3689), .A4(n3688), .ZN(n3692)
         );
  OAI21_X1 U4568 ( .B1(n3693), .B2(n3692), .A(n3739), .ZN(n3694) );
  NAND2_X1 U4569 ( .A1(n3695), .A2(n3694), .ZN(n3696) );
  AOI21_X1 U4570 ( .B1(n5445), .B2(n5205), .A(n3696), .ZN(n5009) );
  INV_X1 U4571 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5982) );
  XOR2_X1 U4572 ( .A(n5982), .B(n3710), .Z(n5984) );
  AOI22_X1 U4573 ( .A1(n5276), .A2(EAX_REG_13__SCAN_IN), .B1(n5275), .B2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3709) );
  AOI22_X1 U4574 ( .A1(n5139), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4575 ( .A1(n5138), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5146), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4576 ( .A1(n3027), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4577 ( .A1(n5083), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3698) );
  NAND4_X1 U4578 ( .A1(n3701), .A2(n3700), .A3(n3699), .A4(n3698), .ZN(n3707)
         );
  AOI22_X1 U4579 ( .A1(n3734), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4580 ( .A1(n5145), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4581 ( .A1(n5147), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n5149), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4582 ( .A1(n5137), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3702) );
  NAND4_X1 U4583 ( .A1(n3705), .A2(n3704), .A3(n3703), .A4(n3702), .ZN(n3706)
         );
  OAI21_X1 U4584 ( .B1(n3707), .B2(n3706), .A(n3739), .ZN(n3708) );
  OAI211_X1 U4585 ( .C1(n5984), .C2(n5211), .A(n3709), .B(n3708), .ZN(n5014)
         );
  NAND2_X1 U4586 ( .A1(n5006), .A2(n5014), .ZN(n5013) );
  XNOR2_X1 U4587 ( .A(n3728), .B(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5435)
         );
  AOI22_X1 U4588 ( .A1(n5145), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3734), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4589 ( .A1(n5137), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n5146), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3713) );
  AOI22_X1 U4590 ( .A1(n5138), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3712) );
  AOI22_X1 U4591 ( .A1(n5147), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3711) );
  NAND4_X1 U4592 ( .A1(n3714), .A2(n3713), .A3(n3712), .A4(n3711), .ZN(n3720)
         );
  AOI22_X1 U4593 ( .A1(n5105), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4594 ( .A1(n5139), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4595 ( .A1(n3289), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5149), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4596 ( .A1(n3027), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3715) );
  NAND4_X1 U4597 ( .A1(n3718), .A2(n3717), .A3(n3716), .A4(n3715), .ZN(n3719)
         );
  NOR2_X1 U4598 ( .A1(n3720), .A2(n3719), .ZN(n3723) );
  NAND2_X1 U4599 ( .A1(n5276), .A2(EAX_REG_14__SCAN_IN), .ZN(n3722) );
  NAND2_X1 U4600 ( .A1(n5275), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3721)
         );
  OAI211_X1 U4601 ( .C1(n3724), .C2(n3723), .A(n3722), .B(n3721), .ZN(n3725)
         );
  AOI21_X1 U4602 ( .B1(n5435), .B2(n5205), .A(n3725), .ZN(n5257) );
  NAND2_X1 U4603 ( .A1(n3728), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3729)
         );
  INV_X1 U4604 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6771) );
  AOI21_X1 U4605 ( .B1(n3729), .B2(n6771), .A(n3784), .ZN(n5631) );
  OR2_X1 U4606 ( .A1(n5631), .A2(n5211), .ZN(n3744) );
  AOI22_X1 U4607 ( .A1(n5276), .A2(EAX_REG_15__SCAN_IN), .B1(n5275), .B2(
        PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3743) );
  AOI22_X1 U4608 ( .A1(n5145), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4609 ( .A1(n5139), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n5147), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3732) );
  AOI22_X1 U4610 ( .A1(n5137), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5146), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4611 ( .A1(n3027), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3730) );
  NAND4_X1 U4612 ( .A1(n3733), .A2(n3732), .A3(n3731), .A4(n3730), .ZN(n3741)
         );
  AOI22_X1 U4613 ( .A1(n3734), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4614 ( .A1(n5144), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4615 ( .A1(n3291), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n5149), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4616 ( .A1(n5138), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3735) );
  NAND4_X1 U4617 ( .A1(n3738), .A2(n3737), .A3(n3736), .A4(n3735), .ZN(n3740)
         );
  OAI21_X1 U4618 ( .B1(n3741), .B2(n3740), .A(n3739), .ZN(n3742) );
  XNOR2_X1 U4619 ( .A(n3784), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5625)
         );
  NAND2_X1 U4620 ( .A1(n5625), .A2(n5205), .ZN(n3759) );
  AOI22_X1 U4621 ( .A1(n3734), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3748) );
  AOI22_X1 U4622 ( .A1(n5145), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3747) );
  AOI22_X1 U4623 ( .A1(n5147), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3746) );
  AOI22_X1 U4624 ( .A1(n5148), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5149), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3745) );
  NAND4_X1 U4625 ( .A1(n3748), .A2(n3747), .A3(n3746), .A4(n3745), .ZN(n3754)
         );
  AOI22_X1 U4626 ( .A1(n5139), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4627 ( .A1(n5138), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4628 ( .A1(n5146), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4629 ( .A1(n5137), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3749) );
  NAND4_X1 U4630 ( .A1(n3752), .A2(n3751), .A3(n3750), .A4(n3749), .ZN(n3753)
         );
  NOR2_X1 U4631 ( .A1(n3754), .A2(n3753), .ZN(n3756) );
  AOI22_X1 U4632 ( .A1(n5276), .A2(EAX_REG_16__SCAN_IN), .B1(n5275), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3755) );
  OAI21_X1 U4633 ( .B1(n5208), .B2(n3756), .A(n3755), .ZN(n3757) );
  INV_X1 U4634 ( .A(n3757), .ZN(n3758) );
  NAND2_X1 U4635 ( .A1(n3759), .A2(n3758), .ZN(n5403) );
  AOI22_X1 U4636 ( .A1(n5105), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3763) );
  AOI22_X1 U4637 ( .A1(n5138), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3762) );
  AOI22_X1 U4638 ( .A1(n5146), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3761) );
  AOI22_X1 U4639 ( .A1(n5137), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3760) );
  NAND4_X1 U4640 ( .A1(n3763), .A2(n3762), .A3(n3761), .A4(n3760), .ZN(n3769)
         );
  AOI22_X1 U4641 ( .A1(n5145), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3734), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3767) );
  AOI22_X1 U4642 ( .A1(n5139), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3766) );
  AOI22_X1 U4643 ( .A1(n5147), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3765) );
  AOI22_X1 U4644 ( .A1(n5148), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5149), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3764) );
  NAND4_X1 U4645 ( .A1(n3767), .A2(n3766), .A3(n3765), .A4(n3764), .ZN(n3768)
         );
  NOR2_X1 U4646 ( .A1(n3769), .A2(n3768), .ZN(n3897) );
  AOI22_X1 U4647 ( .A1(n5145), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4648 ( .A1(n5138), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3772) );
  AOI22_X1 U4649 ( .A1(n5147), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5149), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3771) );
  AOI22_X1 U4650 ( .A1(n5137), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3770) );
  NAND4_X1 U4651 ( .A1(n3773), .A2(n3772), .A3(n3771), .A4(n3770), .ZN(n3779)
         );
  AOI22_X1 U4652 ( .A1(n3734), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3777) );
  AOI22_X1 U4653 ( .A1(n5139), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3776) );
  AOI22_X1 U4654 ( .A1(n5146), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4655 ( .A1(n3289), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3774) );
  NAND4_X1 U4656 ( .A1(n3777), .A2(n3776), .A3(n3775), .A4(n3774), .ZN(n3778)
         );
  NOR2_X1 U4657 ( .A1(n3779), .A2(n3778), .ZN(n3898) );
  XNOR2_X1 U4658 ( .A(n3897), .B(n3898), .ZN(n3783) );
  NAND2_X1 U4659 ( .A1(n6486), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3780)
         );
  NAND2_X1 U4660 ( .A1(n5211), .A2(n3780), .ZN(n3781) );
  AOI21_X1 U4661 ( .B1(n3888), .B2(EAX_REG_23__SCAN_IN), .A(n3781), .ZN(n3782)
         );
  OAI21_X1 U4662 ( .B1(n5208), .B2(n3783), .A(n3782), .ZN(n3788) );
  INV_X1 U4663 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6758) );
  INV_X1 U4664 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5606) );
  OAI21_X1 U4665 ( .B1(n3786), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n3910), 
        .ZN(n5821) );
  OR2_X1 U4666 ( .A1(n5821), .A2(n5211), .ZN(n3787) );
  NAND2_X1 U4667 ( .A1(n3788), .A2(n3787), .ZN(n4124) );
  INV_X1 U4668 ( .A(n4124), .ZN(n3895) );
  AOI22_X1 U4669 ( .A1(n3734), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5146), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3792) );
  AOI22_X1 U4670 ( .A1(n5138), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3791) );
  AOI22_X1 U4671 ( .A1(n3027), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3790) );
  AOI22_X1 U4672 ( .A1(n5149), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3789) );
  NAND4_X1 U4673 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(n3798)
         );
  AOI22_X1 U4674 ( .A1(n5145), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4675 ( .A1(n5144), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3795) );
  AOI22_X1 U4676 ( .A1(n5139), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3794) );
  AOI22_X1 U4677 ( .A1(n5147), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3291), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3793) );
  NAND4_X1 U4678 ( .A1(n3796), .A2(n3795), .A3(n3794), .A4(n3793), .ZN(n3797)
         );
  NOR2_X1 U4679 ( .A1(n3798), .A2(n3797), .ZN(n3799) );
  OR2_X1 U4680 ( .A1(n5208), .A2(n3799), .ZN(n3805) );
  NAND2_X1 U4681 ( .A1(n6486), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3800)
         );
  NAND2_X1 U4682 ( .A1(n5211), .A2(n3800), .ZN(n3801) );
  AOI21_X1 U4683 ( .B1(n3888), .B2(EAX_REG_21__SCAN_IN), .A(n3801), .ZN(n3804)
         );
  OAI21_X1 U4684 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n3802), .A(n3891), 
        .ZN(n5836) );
  NOR2_X1 U4685 ( .A1(n5836), .A2(n5211), .ZN(n3803) );
  AOI21_X1 U4686 ( .B1(n3805), .B2(n3804), .A(n3803), .ZN(n4139) );
  AOI22_X1 U4687 ( .A1(n3734), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3809) );
  AOI22_X1 U4688 ( .A1(n5145), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3808) );
  AOI22_X1 U4689 ( .A1(n5139), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3807) );
  AOI22_X1 U4690 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5147), .B1(n5083), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3806) );
  NAND4_X1 U4691 ( .A1(n3809), .A2(n3808), .A3(n3807), .A4(n3806), .ZN(n3815)
         );
  AOI22_X1 U4692 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n5138), .B1(n5137), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4693 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n3027), .B1(n5148), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4694 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n5146), .B1(n3291), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3811) );
  AOI22_X1 U4695 ( .A1(n5149), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3810) );
  NAND4_X1 U4696 ( .A1(n3813), .A2(n3812), .A3(n3811), .A4(n3810), .ZN(n3814)
         );
  NOR2_X1 U4697 ( .A1(n3815), .A2(n3814), .ZN(n3818) );
  AOI21_X1 U4698 ( .B1(n5606), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3816) );
  AOI21_X1 U4699 ( .B1(n3888), .B2(EAX_REG_20__SCAN_IN), .A(n3816), .ZN(n3817)
         );
  OAI21_X1 U4700 ( .B1(n5208), .B2(n3818), .A(n3817), .ZN(n3820) );
  XNOR2_X1 U4701 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n3835), .ZN(n5610)
         );
  NAND2_X1 U4702 ( .A1(n5205), .A2(n5610), .ZN(n3819) );
  AND2_X1 U4703 ( .A1(n3820), .A2(n3819), .ZN(n5375) );
  INV_X1 U4704 ( .A(n5375), .ZN(n3856) );
  AOI22_X1 U4705 ( .A1(n5145), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3734), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3824) );
  AOI22_X1 U4706 ( .A1(n5144), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3823) );
  AOI22_X1 U4707 ( .A1(n5138), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3822) );
  AOI22_X1 U4708 ( .A1(n5147), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3821) );
  NAND4_X1 U4709 ( .A1(n3824), .A2(n3823), .A3(n3822), .A4(n3821), .ZN(n3830)
         );
  AOI22_X1 U4710 ( .A1(n5139), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4711 ( .A1(n5137), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4712 ( .A1(n5146), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4713 ( .A1(n5149), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3825) );
  NAND4_X1 U4714 ( .A1(n3828), .A2(n3827), .A3(n3826), .A4(n3825), .ZN(n3829)
         );
  NOR2_X1 U4715 ( .A1(n3830), .A2(n3829), .ZN(n3834) );
  OAI21_X1 U4716 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6487), .A(n6486), 
        .ZN(n3831) );
  INV_X1 U4717 ( .A(n3831), .ZN(n3832) );
  AOI21_X1 U4718 ( .B1(n3888), .B2(EAX_REG_19__SCAN_IN), .A(n3832), .ZN(n3833)
         );
  OAI21_X1 U4719 ( .B1(n5208), .B2(n3834), .A(n3833), .ZN(n3837) );
  OAI21_X1 U4720 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n3851), .A(n3835), 
        .ZN(n5884) );
  OR2_X1 U4721 ( .A1(n5211), .A2(n5884), .ZN(n3836) );
  NAND2_X1 U4722 ( .A1(n3837), .A2(n3836), .ZN(n5842) );
  AOI22_X1 U4723 ( .A1(n3734), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4724 ( .A1(n5100), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5147), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4725 ( .A1(n5137), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3839) );
  AOI22_X1 U4726 ( .A1(n5146), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n5149), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3838) );
  NAND4_X1 U4727 ( .A1(n3841), .A2(n3840), .A3(n3839), .A4(n3838), .ZN(n3847)
         );
  AOI22_X1 U4728 ( .A1(n5145), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4729 ( .A1(n5138), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4730 ( .A1(n5139), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3843) );
  AOI22_X1 U4731 ( .A1(n3273), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3842) );
  NAND4_X1 U4732 ( .A1(n3845), .A2(n3844), .A3(n3843), .A4(n3842), .ZN(n3846)
         );
  NOR2_X1 U4733 ( .A1(n3847), .A2(n3846), .ZN(n3850) );
  OAI21_X1 U4734 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6758), .A(n5211), .ZN(
        n3848) );
  AOI21_X1 U4735 ( .B1(n5276), .B2(EAX_REG_18__SCAN_IN), .A(n3848), .ZN(n3849)
         );
  OAI21_X1 U4736 ( .B1(n5208), .B2(n3850), .A(n3849), .ZN(n3855) );
  INV_X1 U4737 ( .A(n3870), .ZN(n3853) );
  INV_X1 U4738 ( .A(n3851), .ZN(n3852) );
  OAI21_X1 U4739 ( .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n3853), .A(n3852), 
        .ZN(n5620) );
  OR2_X1 U4740 ( .A1(n5211), .A2(n5620), .ZN(n3854) );
  NAND2_X1 U4741 ( .A1(n3855), .A2(n3854), .ZN(n5390) );
  OR2_X1 U4742 ( .A1(n5842), .A2(n5390), .ZN(n5374) );
  NOR2_X1 U4743 ( .A1(n3856), .A2(n5374), .ZN(n4137) );
  AND2_X1 U4744 ( .A1(n4139), .A2(n4137), .ZN(n3875) );
  AOI22_X1 U4745 ( .A1(n5144), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4746 ( .A1(n5138), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4747 ( .A1(n5147), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n5146), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3858) );
  AOI22_X1 U4748 ( .A1(n5149), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3857) );
  NAND4_X1 U4749 ( .A1(n3860), .A2(n3859), .A3(n3858), .A4(n3857), .ZN(n3866)
         );
  AOI22_X1 U4750 ( .A1(n3734), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4751 ( .A1(n5145), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n5139), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4752 ( .A1(n3027), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4753 ( .A1(n5083), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3861) );
  NAND4_X1 U4754 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), .ZN(n3865)
         );
  NOR2_X1 U4755 ( .A1(n3866), .A2(n3865), .ZN(n3867) );
  OR2_X1 U4756 ( .A1(n5208), .A2(n3867), .ZN(n3874) );
  NAND2_X1 U4757 ( .A1(n6486), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3868)
         );
  NAND2_X1 U4758 ( .A1(n5211), .A2(n3868), .ZN(n3869) );
  AOI21_X1 U4759 ( .B1(n3888), .B2(EAX_REG_17__SCAN_IN), .A(n3869), .ZN(n3873)
         );
  OAI21_X1 U4760 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3871), .A(n3870), 
        .ZN(n5977) );
  NOR2_X1 U4761 ( .A1(n5977), .A2(n5211), .ZN(n3872) );
  AOI21_X1 U4762 ( .B1(n3874), .B2(n3873), .A(n3872), .ZN(n5894) );
  AND2_X1 U4763 ( .A1(n3875), .A2(n5894), .ZN(n4136) );
  AOI22_X1 U4764 ( .A1(n3734), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4765 ( .A1(n5145), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3878) );
  AOI22_X1 U4766 ( .A1(n5138), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3877) );
  AOI22_X1 U4767 ( .A1(n5100), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3876) );
  NAND4_X1 U4768 ( .A1(n3879), .A2(n3878), .A3(n3877), .A4(n3876), .ZN(n3885)
         );
  AOI22_X1 U4769 ( .A1(n5139), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5147), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4770 ( .A1(n5137), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3027), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4771 ( .A1(n5146), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4772 ( .A1(n5149), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3880) );
  NAND4_X1 U4773 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3884)
         );
  NOR2_X1 U4774 ( .A1(n3885), .A2(n3884), .ZN(n3890) );
  NAND2_X1 U4775 ( .A1(n6486), .A2(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n3886)
         );
  NAND2_X1 U4776 ( .A1(n5211), .A2(n3886), .ZN(n3887) );
  AOI21_X1 U4777 ( .B1(n3888), .B2(EAX_REG_22__SCAN_IN), .A(n3887), .ZN(n3889)
         );
  OAI21_X1 U4778 ( .B1(n5208), .B2(n3890), .A(n3889), .ZN(n3893) );
  XNOR2_X1 U4779 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .B(n3891), .ZN(n5601)
         );
  NAND2_X1 U4780 ( .A1(n5205), .A2(n5601), .ZN(n3892) );
  NAND2_X1 U4781 ( .A1(n3893), .A2(n3892), .ZN(n5359) );
  INV_X1 U4782 ( .A(n5359), .ZN(n3894) );
  NOR2_X1 U4783 ( .A1(n3898), .A2(n3897), .ZN(n5113) );
  AOI22_X1 U4784 ( .A1(n3734), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4785 ( .A1(n5145), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4786 ( .A1(n5139), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3900) );
  AOI22_X1 U4787 ( .A1(n5147), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3899) );
  NAND4_X1 U4788 ( .A1(n3902), .A2(n3901), .A3(n3900), .A4(n3899), .ZN(n3908)
         );
  AOI22_X1 U4789 ( .A1(n5138), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3906) );
  AOI22_X1 U4790 ( .A1(n3027), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3905) );
  AOI22_X1 U4791 ( .A1(n5146), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3904) );
  AOI22_X1 U4792 ( .A1(n5149), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3903) );
  NAND4_X1 U4793 ( .A1(n3906), .A2(n3905), .A3(n3904), .A4(n3903), .ZN(n3907)
         );
  OR2_X1 U4794 ( .A1(n3908), .A2(n3907), .ZN(n5112) );
  INV_X1 U4795 ( .A(n5112), .ZN(n3909) );
  XNOR2_X1 U4796 ( .A(n5113), .B(n3909), .ZN(n3918) );
  INV_X1 U4797 ( .A(n5208), .ZN(n5158) );
  INV_X1 U4798 ( .A(EAX_REG_24__SCAN_IN), .ZN(n3915) );
  INV_X1 U4799 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6636) );
  AND2_X1 U4800 ( .A1(n3910), .A2(n6636), .ZN(n3911) );
  NOR2_X1 U4801 ( .A1(n5169), .A2(n3911), .ZN(n5812) );
  OAI22_X1 U4802 ( .A1(n5812), .A2(n5211), .B1(n6636), .B2(n3912), .ZN(n3913)
         );
  INV_X1 U4803 ( .A(n3913), .ZN(n3914) );
  OAI21_X1 U4804 ( .B1(n3916), .B2(n3915), .A(n3914), .ZN(n3917) );
  AOI21_X1 U4805 ( .B1(n3918), .B2(n5158), .A(n3917), .ZN(n3919) );
  AND2_X1 U4806 ( .A1(n3920), .A2(n3919), .ZN(n3921) );
  OR2_X1 U4807 ( .A1(n3921), .A2(n5173), .ZN(n5815) );
  INV_X1 U4808 ( .A(n5815), .ZN(n3922) );
  AND2_X1 U4809 ( .A1(n6780), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4944) );
  NAND2_X1 U4810 ( .A1(n4944), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6494) );
  NOR2_X2 U4811 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6343) );
  INV_X1 U4812 ( .A(n6343), .ZN(n6382) );
  OR2_X2 U4813 ( .A1(n6494), .A2(n6382), .ZN(n6199) );
  NAND2_X1 U4814 ( .A1(n3922), .A2(n6183), .ZN(n3930) );
  NAND2_X1 U4815 ( .A1(n6382), .A2(n3926), .ZN(n6595) );
  NAND2_X1 U4816 ( .A1(n6595), .A2(n6780), .ZN(n3923) );
  NAND2_X1 U4817 ( .A1(n6780), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3925) );
  NAND2_X1 U4818 ( .A1(n6487), .A2(STATE2_REG_1__SCAN_IN), .ZN(n3924) );
  NAND2_X1 U4819 ( .A1(n3925), .A2(n3924), .ZN(n6195) );
  OR2_X1 U4820 ( .A1(n3926), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6242) );
  INV_X2 U4821 ( .A(n6242), .ZN(n6218) );
  AND2_X1 U4822 ( .A1(n6218), .A2(REIP_REG_24__SCAN_IN), .ZN(n5223) );
  INV_X1 U4823 ( .A(n5223), .ZN(n3927) );
  OAI21_X1 U4824 ( .B1(n6174), .B2(n6636), .A(n3927), .ZN(n3928) );
  AOI21_X1 U4825 ( .B1(n6168), .B2(n5812), .A(n3928), .ZN(n3929) );
  OAI21_X1 U4826 ( .B1(n5226), .B2(n6190), .A(n3931), .ZN(U2962) );
  INV_X1 U4827 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6744) );
  NOR2_X1 U4828 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5687) );
  NOR4_X1 U4829 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .A3(INSTADDRPOINTER_REG_22__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3932) );
  AOI21_X1 U4830 ( .B1(n5687), .B2(n3932), .A(n5890), .ZN(n3933) );
  AND2_X1 U4831 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5688) );
  AND2_X1 U4832 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5231) );
  AND2_X1 U4833 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4110) );
  NAND3_X1 U4834 ( .A1(n5688), .A2(n5231), .A3(n4110), .ZN(n4094) );
  NOR2_X2 U4835 ( .A1(n3934), .A2(n3038), .ZN(n5874) );
  XOR2_X1 U4836 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .B(n5890), .Z(n5873) );
  NOR2_X2 U4837 ( .A1(n5874), .A2(n5873), .ZN(n3936) );
  AOI21_X2 U4838 ( .B1(n5890), .B2(n6744), .A(n3936), .ZN(n5576) );
  INV_X1 U4839 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5668) );
  NOR2_X1 U4840 ( .A1(n3500), .A2(n5668), .ZN(n5587) );
  NAND2_X1 U4841 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5644) );
  INV_X1 U4842 ( .A(n5644), .ZN(n4096) );
  AND2_X1 U4843 ( .A1(n5587), .A2(n4096), .ZN(n3935) );
  NAND2_X1 U4844 ( .A1(n5560), .A2(n3046), .ZN(n3939) );
  INV_X1 U4845 ( .A(n3936), .ZN(n5875) );
  NAND2_X1 U4846 ( .A1(n3500), .A2(n5668), .ZN(n5585) );
  NOR3_X1 U4847 ( .A1(n5585), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5065) );
  INV_X1 U4848 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n6735) );
  INV_X1 U4849 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5648) );
  NAND3_X1 U4850 ( .A1(n5065), .A2(n6735), .A3(n5648), .ZN(n3937) );
  INV_X1 U4851 ( .A(READY_N), .ZN(n6596) );
  NAND2_X1 U4852 ( .A1(n3942), .A2(n6596), .ZN(n3943) );
  NAND2_X1 U4853 ( .A1(n3943), .A2(n3030), .ZN(n3945) );
  INV_X1 U4854 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6508) );
  NAND2_X1 U4855 ( .A1(n3944), .A2(n6508), .ZN(n6503) );
  INV_X1 U4856 ( .A(n6503), .ZN(n4967) );
  OAI22_X1 U4857 ( .A1(n4232), .A2(n3945), .B1(n4967), .B2(n6599), .ZN(n3947)
         );
  NAND2_X1 U4858 ( .A1(n3947), .A2(n3946), .ZN(n3949) );
  OAI22_X1 U4859 ( .A1(n4232), .A2(n4188), .B1(n4402), .B2(n6437), .ZN(n3948)
         );
  NAND2_X1 U4860 ( .A1(n3949), .A2(n3948), .ZN(n3965) );
  OR2_X1 U4861 ( .A1(n3950), .A2(n3026), .ZN(n4090) );
  OAI211_X1 U4862 ( .C1(n3951), .C2(n3129), .A(n4965), .B(n4090), .ZN(n4082)
         );
  INV_X1 U4863 ( .A(n4082), .ZN(n3952) );
  OR2_X1 U4864 ( .A1(n3952), .A2(n6461), .ZN(n3955) );
  NOR2_X1 U4865 ( .A1(n6460), .A2(n4965), .ZN(n3953) );
  NAND2_X1 U4866 ( .A1(n3954), .A2(n3953), .ZN(n4153) );
  NAND2_X1 U4867 ( .A1(n3955), .A2(n4153), .ZN(n4205) );
  NAND2_X1 U4868 ( .A1(n4968), .A2(n6503), .ZN(n3962) );
  NAND2_X1 U4869 ( .A1(n3957), .A2(n3956), .ZN(n3960) );
  INV_X1 U4870 ( .A(n3958), .ZN(n3959) );
  OAI21_X1 U4871 ( .B1(n3961), .B2(n3960), .A(n3959), .ZN(n4154) );
  NOR2_X1 U4872 ( .A1(READY_N), .A2(n4154), .ZN(n4207) );
  NAND3_X1 U4873 ( .A1(n3962), .A2(n4207), .A3(n4188), .ZN(n3963) );
  AND2_X1 U4874 ( .A1(n4205), .A2(n3963), .ZN(n3964) );
  NAND2_X1 U4875 ( .A1(n3965), .A2(n3964), .ZN(n3966) );
  AND2_X1 U4876 ( .A1(n3029), .A2(n3967), .ZN(n3982) );
  INV_X1 U4877 ( .A(n4073), .ZN(n3968) );
  AOI22_X1 U4878 ( .A1(n3942), .A2(n4303), .B1(n3968), .B2(n4072), .ZN(n3972)
         );
  INV_X1 U4879 ( .A(n6460), .ZN(n3970) );
  NOR2_X1 U4880 ( .A1(n3970), .A2(n4948), .ZN(n3971) );
  OR2_X1 U4881 ( .A1(n6461), .A2(n3971), .ZN(n4152) );
  NAND3_X1 U4882 ( .A1(n3972), .A2(n4152), .A3(n4216), .ZN(n3973) );
  NAND2_X1 U4883 ( .A1(n4384), .A2(n3033), .ZN(n3986) );
  INV_X1 U4884 ( .A(n3986), .ZN(n4024) );
  NAND2_X1 U4885 ( .A1(n3986), .A2(n6246), .ZN(n3976) );
  BUF_X2 U4886 ( .A(n3974), .Z(n3983) );
  INV_X1 U4887 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4973) );
  NAND2_X1 U4888 ( .A1(n3982), .A2(n4973), .ZN(n3975) );
  NAND3_X1 U4889 ( .A1(n3976), .A2(n3983), .A3(n3975), .ZN(n3978) );
  NAND2_X1 U4890 ( .A1(n3978), .A2(n3977), .ZN(n3981) );
  NAND2_X1 U4891 ( .A1(n3986), .A2(EBX_REG_0__SCAN_IN), .ZN(n3980) );
  INV_X1 U4892 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4199) );
  NAND2_X1 U4893 ( .A1(n3983), .A2(n4199), .ZN(n3979) );
  NAND2_X1 U4894 ( .A1(n3980), .A2(n3979), .ZN(n4196) );
  NAND2_X1 U4895 ( .A1(n4302), .A2(n3981), .ZN(n4321) );
  INV_X2 U4896 ( .A(n3982), .ZN(n4962) );
  NAND2_X1 U4897 ( .A1(n3983), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3984)
         );
  OAI211_X1 U4898 ( .C1(n4962), .C2(EBX_REG_3__SCAN_IN), .A(n4048), .B(n3984), 
        .ZN(n3985) );
  OAI21_X1 U4899 ( .B1(n4056), .B2(EBX_REG_3__SCAN_IN), .A(n3985), .ZN(n4319)
         );
  MUX2_X1 U4900 ( .A(n3983), .B(n3986), .S(EBX_REG_2__SCAN_IN), .Z(n3988) );
  NAND2_X1 U4901 ( .A1(n4962), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3987)
         );
  NAND2_X1 U4902 ( .A1(n3988), .A2(n3987), .ZN(n4273) );
  INV_X1 U4903 ( .A(n4273), .ZN(n4320) );
  NAND2_X1 U4904 ( .A1(n4048), .A2(n3367), .ZN(n3992) );
  INV_X1 U4905 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U4906 ( .A1(n4303), .A2(n6079), .ZN(n3991) );
  NAND3_X1 U4907 ( .A1(n3992), .A2(n3031), .A3(n3991), .ZN(n3994) );
  NAND2_X1 U4908 ( .A1(n5381), .A2(n6079), .ZN(n3993) );
  MUX2_X1 U4909 ( .A(n4056), .B(n3031), .S(EBX_REG_5__SCAN_IN), .Z(n3996) );
  NAND2_X1 U4910 ( .A1(n4198), .A2(n3445), .ZN(n3995) );
  NAND2_X1 U4911 ( .A1(n4364), .A2(n3035), .ZN(n4534) );
  INV_X1 U4912 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3997) );
  NAND2_X1 U4913 ( .A1(n4048), .A2(n3997), .ZN(n3999) );
  INV_X1 U4914 ( .A(EBX_REG_6__SCAN_IN), .ZN(n4000) );
  NAND2_X1 U4915 ( .A1(n4303), .A2(n4000), .ZN(n3998) );
  NAND3_X1 U4916 ( .A1(n3999), .A2(n3031), .A3(n3998), .ZN(n4002) );
  NAND2_X1 U4917 ( .A1(n5381), .A2(n4000), .ZN(n4001) );
  MUX2_X1 U4918 ( .A(n4056), .B(n3031), .S(EBX_REG_7__SCAN_IN), .Z(n4004) );
  OAI21_X1 U4919 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n4069), .A(n4004), 
        .ZN(n4765) );
  INV_X1 U4920 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4005) );
  NAND2_X1 U4921 ( .A1(n4048), .A2(n4005), .ZN(n4007) );
  INV_X1 U4922 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U4923 ( .A1(n4303), .A2(n5470), .ZN(n4006) );
  NAND3_X1 U4924 ( .A1(n4007), .A2(n3031), .A3(n4006), .ZN(n4009) );
  NAND2_X1 U4925 ( .A1(n5381), .A2(n5470), .ZN(n4008) );
  NAND2_X1 U4926 ( .A1(n4009), .A2(n4008), .ZN(n4912) );
  AND2_X2 U4927 ( .A1(n4913), .A2(n4912), .ZN(n4926) );
  MUX2_X1 U4928 ( .A(n4056), .B(n3031), .S(EBX_REG_9__SCAN_IN), .Z(n4011) );
  OR2_X1 U4929 ( .A1(n4069), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4010)
         );
  MUX2_X1 U4930 ( .A(n3031), .B(n4048), .S(EBX_REG_10__SCAN_IN), .Z(n4013) );
  NAND2_X1 U4931 ( .A1(n4962), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4012) );
  AND2_X1 U4932 ( .A1(n4013), .A2(n4012), .ZN(n4987) );
  NAND2_X1 U4933 ( .A1(n3031), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4014) );
  OAI211_X1 U4934 ( .C1(n4962), .C2(EBX_REG_11__SCAN_IN), .A(n4048), .B(n4014), 
        .ZN(n4015) );
  OAI21_X1 U4935 ( .B1(n4056), .B2(EBX_REG_11__SCAN_IN), .A(n4015), .ZN(n5992)
         );
  NOR2_X2 U4936 ( .A1(n5993), .A2(n5992), .ZN(n5994) );
  MUX2_X1 U4937 ( .A(n3031), .B(n4048), .S(EBX_REG_12__SCAN_IN), .Z(n4017) );
  NAND2_X1 U4938 ( .A1(n4962), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4016) );
  NAND2_X1 U4939 ( .A1(n4017), .A2(n4016), .ZN(n5028) );
  NAND2_X1 U4940 ( .A1(n5994), .A2(n5028), .ZN(n5927) );
  NAND2_X1 U4941 ( .A1(n3031), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4018) );
  OAI211_X1 U4942 ( .C1(n4962), .C2(EBX_REG_13__SCAN_IN), .A(n4048), .B(n4018), 
        .ZN(n4019) );
  OAI21_X1 U4943 ( .B1(n4056), .B2(EBX_REG_13__SCAN_IN), .A(n4019), .ZN(n5926)
         );
  OR2_X2 U4944 ( .A1(n5927), .A2(n5926), .ZN(n5929) );
  MUX2_X1 U4945 ( .A(n4065), .B(n4048), .S(EBX_REG_14__SCAN_IN), .Z(n4021) );
  NAND2_X1 U4946 ( .A1(n4962), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4020) );
  AND2_X1 U4947 ( .A1(n4021), .A2(n4020), .ZN(n5248) );
  OR2_X2 U4948 ( .A1(n5929), .A2(n5248), .ZN(n5425) );
  NAND2_X1 U4949 ( .A1(n3031), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4022) );
  OAI211_X1 U4950 ( .C1(n4962), .C2(EBX_REG_15__SCAN_IN), .A(n4048), .B(n4022), 
        .ZN(n4023) );
  OAI21_X1 U4951 ( .B1(n4056), .B2(EBX_REG_15__SCAN_IN), .A(n4023), .ZN(n5424)
         );
  INV_X1 U4952 ( .A(n4024), .ZN(n4048) );
  MUX2_X1 U4953 ( .A(n4065), .B(n4048), .S(EBX_REG_16__SCAN_IN), .Z(n4026) );
  NAND2_X1 U4954 ( .A1(n4962), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4025) );
  NAND2_X1 U4955 ( .A1(n4026), .A2(n4025), .ZN(n5405) );
  AND2_X2 U4956 ( .A1(n5427), .A2(n5405), .ZN(n5908) );
  INV_X1 U4957 ( .A(n4056), .ZN(n4027) );
  INV_X1 U4958 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6083) );
  NAND2_X1 U4959 ( .A1(n4027), .A2(n6083), .ZN(n4030) );
  NAND2_X1 U4960 ( .A1(n4065), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4028) );
  OAI211_X1 U4961 ( .C1(n4962), .C2(EBX_REG_17__SCAN_IN), .A(n4048), .B(n4028), 
        .ZN(n4029) );
  AND2_X1 U4962 ( .A1(n4030), .A2(n4029), .ZN(n5907) );
  NAND2_X1 U4963 ( .A1(n5908), .A2(n5907), .ZN(n5391) );
  NAND2_X1 U4964 ( .A1(n4048), .A2(n5705), .ZN(n4032) );
  INV_X1 U4965 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5856) );
  NAND2_X1 U4966 ( .A1(n4303), .A2(n5856), .ZN(n4031) );
  NAND3_X1 U4967 ( .A1(n4032), .A2(n4065), .A3(n4031), .ZN(n4034) );
  NAND2_X1 U4968 ( .A1(n5381), .A2(n5856), .ZN(n4033) );
  AND2_X1 U4969 ( .A1(n4034), .A2(n4033), .ZN(n5701) );
  OR2_X2 U4970 ( .A1(n5391), .A2(n5701), .ZN(n5380) );
  NAND2_X1 U4971 ( .A1(n4069), .A2(EBX_REG_18__SCAN_IN), .ZN(n4036) );
  NAND2_X1 U4972 ( .A1(n4962), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4035) );
  NAND2_X1 U4973 ( .A1(n4036), .A2(n4035), .ZN(n5382) );
  OR2_X1 U4974 ( .A1(n5382), .A2(n3031), .ZN(n5393) );
  AND2_X1 U4975 ( .A1(n4962), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4037)
         );
  AOI21_X1 U4976 ( .B1(n4069), .B2(EBX_REG_20__SCAN_IN), .A(n4037), .ZN(n5383)
         );
  NAND2_X1 U4977 ( .A1(n5393), .A2(n5383), .ZN(n4040) );
  NAND2_X1 U4978 ( .A1(n5382), .A2(n4065), .ZN(n5392) );
  INV_X1 U4979 ( .A(n5383), .ZN(n4038) );
  NAND2_X1 U4980 ( .A1(n5392), .A2(n4038), .ZN(n4039) );
  NAND2_X1 U4981 ( .A1(n4040), .A2(n4039), .ZN(n4041) );
  MUX2_X1 U4982 ( .A(n4056), .B(n4065), .S(EBX_REG_21__SCAN_IN), .Z(n4043) );
  OR2_X1 U4983 ( .A1(n4069), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4042)
         );
  AND2_X1 U4984 ( .A1(n4043), .A2(n4042), .ZN(n5264) );
  MUX2_X1 U4985 ( .A(n3031), .B(n4048), .S(EBX_REG_22__SCAN_IN), .Z(n4045) );
  NAND2_X1 U4986 ( .A1(n4962), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4044) );
  NAND2_X1 U4987 ( .A1(n4045), .A2(n4044), .ZN(n5366) );
  NAND2_X1 U4988 ( .A1(n3031), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4046) );
  OAI211_X1 U4989 ( .C1(n4962), .C2(EBX_REG_23__SCAN_IN), .A(n4048), .B(n4046), 
        .ZN(n4047) );
  OAI21_X1 U4990 ( .B1(n4056), .B2(EBX_REG_23__SCAN_IN), .A(n4047), .ZN(n5230)
         );
  MUX2_X1 U4991 ( .A(n4065), .B(n4048), .S(EBX_REG_24__SCAN_IN), .Z(n4050) );
  NAND2_X1 U4992 ( .A1(n4962), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4049) );
  AND2_X1 U4993 ( .A1(n4050), .A2(n4049), .ZN(n5217) );
  MUX2_X1 U4994 ( .A(n4056), .B(n4065), .S(EBX_REG_25__SCAN_IN), .Z(n4051) );
  OAI21_X1 U4995 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n4069), .A(n4051), 
        .ZN(n5347) );
  NAND2_X1 U4996 ( .A1(n4048), .A2(n5668), .ZN(n4053) );
  INV_X1 U4997 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6738) );
  NAND2_X1 U4998 ( .A1(n4303), .A2(n6738), .ZN(n4052) );
  NAND3_X1 U4999 ( .A1(n4053), .A2(n3031), .A3(n4052), .ZN(n4055) );
  NAND2_X1 U5000 ( .A1(n5381), .A2(n6738), .ZN(n4054) );
  NAND2_X1 U5001 ( .A1(n4055), .A2(n4054), .ZN(n5521) );
  MUX2_X1 U5002 ( .A(n4056), .B(n4065), .S(EBX_REG_27__SCAN_IN), .Z(n4058) );
  OR2_X1 U5003 ( .A1(n4069), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4057)
         );
  AND2_X1 U5004 ( .A1(n4058), .A2(n4057), .ZN(n5514) );
  MUX2_X1 U5005 ( .A(n4065), .B(n4048), .S(EBX_REG_28__SCAN_IN), .Z(n4060) );
  NAND2_X1 U5006 ( .A1(n4962), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4059) );
  NAND2_X1 U5007 ( .A1(n4060), .A2(n4059), .ZN(n5296) );
  NAND2_X1 U5008 ( .A1(n4069), .A2(EBX_REG_29__SCAN_IN), .ZN(n4062) );
  NAND2_X1 U5009 ( .A1(n4962), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4061) );
  NAND2_X1 U5010 ( .A1(n4062), .A2(n4061), .ZN(n5070) );
  OAI21_X1 U5011 ( .B1(n5069), .B2(n5070), .A(n5381), .ZN(n4068) );
  INV_X1 U5012 ( .A(n5069), .ZN(n4066) );
  NAND2_X1 U5013 ( .A1(n4069), .A2(EBX_REG_30__SCAN_IN), .ZN(n4064) );
  NAND2_X1 U5014 ( .A1(n4962), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4063) );
  NAND2_X1 U5015 ( .A1(n4064), .A2(n4063), .ZN(n5071) );
  XNOR2_X1 U5016 ( .A(n5070), .B(n4065), .ZN(n5334) );
  NAND3_X1 U5017 ( .A1(n4066), .A2(n5071), .A3(n5334), .ZN(n4067) );
  NAND2_X1 U5018 ( .A1(n4068), .A2(n4067), .ZN(n4071) );
  OAI22_X1 U5019 ( .A1(n4069), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4962), .ZN(n4070) );
  XNOR2_X1 U5020 ( .A(n4071), .B(n4070), .ZN(n5502) );
  NAND2_X1 U5021 ( .A1(n3942), .A2(n4958), .ZN(n4231) );
  OAI21_X1 U5022 ( .B1(n4073), .B2(n4072), .A(n4231), .ZN(n4074) );
  NAND2_X1 U5023 ( .A1(n6218), .A2(REIP_REG_31__SCAN_IN), .ZN(n5281) );
  INV_X1 U5024 ( .A(n5281), .ZN(n4099) );
  INV_X1 U5025 ( .A(n4093), .ZN(n4101) );
  NAND2_X1 U5026 ( .A1(n4075), .A2(n5381), .ZN(n4080) );
  OR2_X1 U5027 ( .A1(n4076), .A2(n4188), .ZN(n4204) );
  NAND2_X1 U5028 ( .A1(n4198), .A2(n4204), .ZN(n4078) );
  NAND2_X1 U5029 ( .A1(n4078), .A2(n4077), .ZN(n4079) );
  AND4_X1 U5030 ( .A1(n4082), .A2(n4081), .A3(n4080), .A4(n4079), .ZN(n4083)
         );
  AND2_X1 U5031 ( .A1(n4084), .A2(n4083), .ZN(n4218) );
  AOI21_X1 U5032 ( .B1(n3186), .B2(n4409), .A(n3194), .ZN(n4085) );
  OR2_X1 U5033 ( .A1(n4086), .A2(n4085), .ZN(n4213) );
  NAND2_X1 U5034 ( .A1(n4213), .A2(n4087), .ZN(n4088) );
  AND2_X1 U5035 ( .A1(n4088), .A2(n4431), .ZN(n4089) );
  NAND2_X1 U5036 ( .A1(n4218), .A2(n4089), .ZN(n4092) );
  NAND2_X1 U5037 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4690) );
  INV_X1 U5038 ( .A(n4690), .ZN(n5054) );
  NAND2_X1 U5039 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n5054), .ZN(n4533)
         );
  OR2_X1 U5040 ( .A1(n3997), .A2(n4533), .ZN(n4911) );
  AOI21_X1 U5041 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4691) );
  NOR2_X1 U5042 ( .A1(n4911), .A2(n4691), .ZN(n4104) );
  INV_X1 U5043 ( .A(n4104), .ZN(n4091) );
  NAND2_X1 U5044 ( .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6212) );
  INV_X1 U5045 ( .A(n6212), .ZN(n6216) );
  NAND3_X1 U5046 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n6216), .ZN(n4105) );
  NOR3_X1 U5047 ( .A1(n6236), .A2(n4091), .A3(n4105), .ZN(n5247) );
  NAND2_X1 U5048 ( .A1(n4093), .A2(n4092), .ZN(n5244) );
  NOR2_X1 U5049 ( .A1(n4153), .A2(n4402), .ZN(n6442) );
  NAND2_X1 U5050 ( .A1(n4093), .A2(n6442), .ZN(n4285) );
  NAND2_X1 U5051 ( .A1(n5244), .A2(n4285), .ZN(n4318) );
  INV_X1 U5052 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6577) );
  NAND2_X1 U5053 ( .A1(n6577), .A2(n4285), .ZN(n4306) );
  NAND2_X1 U5054 ( .A1(n4318), .A2(n4306), .ZN(n6245) );
  NAND2_X1 U5055 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6237) );
  OR2_X1 U5056 ( .A1(n4911), .A2(n6237), .ZN(n4102) );
  NOR2_X1 U5057 ( .A1(n4102), .A2(n4105), .ZN(n5935) );
  INV_X1 U5058 ( .A(n5935), .ZN(n5243) );
  NOR2_X1 U5059 ( .A1(n6245), .A2(n5243), .ZN(n5024) );
  NAND3_X1 U5060 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .A3(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5722) );
  NOR2_X1 U5061 ( .A1(n5721), .A2(n5722), .ZN(n5719) );
  NAND3_X1 U5062 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5719), .ZN(n4100) );
  NOR2_X1 U5063 ( .A1(n6201), .A2(n4100), .ZN(n5914) );
  NAND2_X1 U5064 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5914), .ZN(n5712) );
  INV_X1 U5065 ( .A(n4094), .ZN(n4095) );
  AND2_X1 U5066 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5666) );
  NAND2_X1 U5067 ( .A1(n5900), .A2(n5666), .ZN(n5659) );
  NAND2_X1 U5068 ( .A1(n4096), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4097) );
  OR2_X1 U5069 ( .A1(n5659), .A2(n4097), .ZN(n5075) );
  NOR3_X1 U5070 ( .A1(n5075), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n6735), 
        .ZN(n4098) );
  AOI211_X1 U5071 ( .C1(n5502), .C2(n6240), .A(n4099), .B(n4098), .ZN(n4115)
         );
  NAND2_X1 U5072 ( .A1(n5244), .A2(n6236), .ZN(n4287) );
  INV_X1 U5073 ( .A(n4100), .ZN(n4106) );
  NAND2_X1 U5074 ( .A1(n4101), .A2(n6242), .ZN(n4308) );
  OAI21_X1 U5075 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n5244), .A(n4308), 
        .ZN(n4317) );
  AOI21_X1 U5076 ( .B1(n4318), .B2(n4102), .A(n4317), .ZN(n4103) );
  OAI21_X1 U5077 ( .B1(n4104), .B2(n6236), .A(n4103), .ZN(n6211) );
  AOI21_X1 U5078 ( .B1(n6213), .B2(n4105), .A(n6211), .ZN(n6210) );
  OAI21_X1 U5079 ( .B1(n5720), .B2(n4106), .A(n6210), .ZN(n5912) );
  NAND2_X1 U5080 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5710) );
  AND2_X1 U5081 ( .A1(n6213), .A2(n5710), .ZN(n4107) );
  NOR2_X1 U5082 ( .A1(n5912), .A2(n4107), .ZN(n5704) );
  INV_X1 U5083 ( .A(n5688), .ZN(n4108) );
  NAND2_X1 U5084 ( .A1(n6213), .A2(n4108), .ZN(n4109) );
  NAND2_X1 U5085 ( .A1(n5704), .A2(n4109), .ZN(n5271) );
  NAND2_X1 U5086 ( .A1(n5686), .A2(n5688), .ZN(n5268) );
  NOR2_X1 U5087 ( .A1(n5268), .A2(n5231), .ZN(n5677) );
  NAND2_X1 U5088 ( .A1(n6236), .A2(n6245), .ZN(n5709) );
  INV_X1 U5089 ( .A(n4110), .ZN(n4111) );
  AND2_X1 U5090 ( .A1(n5709), .A2(n4111), .ZN(n4112) );
  OAI21_X1 U5091 ( .B1(n5720), .B2(n5666), .A(n5906), .ZN(n5663) );
  AOI21_X1 U5092 ( .B1(n5644), .B2(n6213), .A(n5663), .ZN(n5649) );
  OAI21_X1 U5093 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5720), .A(n5649), 
        .ZN(n5077) );
  NOR2_X1 U5094 ( .A1(n5720), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4113)
         );
  OAI21_X1 U5095 ( .B1(n5077), .B2(n4113), .A(INSTADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n4114) );
  AND2_X1 U5096 ( .A1(n4115), .A2(n4114), .ZN(n4116) );
  OAI21_X1 U5097 ( .B1(n5285), .B2(n6203), .A(n4116), .ZN(U2987) );
  XNOR2_X1 U5098 ( .A(n5890), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5604)
         );
  NAND2_X1 U5099 ( .A1(n5605), .A2(n5604), .ZN(n5603) );
  NAND2_X1 U5100 ( .A1(n5688), .A2(n5231), .ZN(n4117) );
  INV_X1 U5101 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4120) );
  INV_X1 U5102 ( .A(n6190), .ZN(n6182) );
  NAND2_X1 U5103 ( .A1(n5227), .A2(n6182), .ZN(n4131) );
  NAND2_X1 U5104 ( .A1(n5895), .A2(n4123), .ZN(n5362) );
  NAND2_X1 U5105 ( .A1(n5362), .A2(n4124), .ZN(n4125) );
  NAND2_X1 U5106 ( .A1(n3920), .A2(n4125), .ZN(n5823) );
  INV_X1 U5107 ( .A(REIP_REG_23__SCAN_IN), .ZN(n4126) );
  NOR2_X1 U5108 ( .A1(n6242), .A2(n4126), .ZN(n5234) );
  NOR2_X1 U5109 ( .A1(n6188), .A2(n5821), .ZN(n4127) );
  AOI211_X1 U5110 ( .C1(n6196), .C2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n5234), 
        .B(n4127), .ZN(n4128) );
  NAND2_X1 U5111 ( .A1(n4131), .A2(n4130), .ZN(U2963) );
  NAND2_X1 U5112 ( .A1(n4135), .A2(n4134), .ZN(n5263) );
  INV_X1 U5113 ( .A(n5836), .ZN(n4141) );
  NAND2_X1 U5114 ( .A1(n5895), .A2(n4136), .ZN(n5360) );
  AND2_X1 U5115 ( .A1(n5895), .A2(n5894), .ZN(n4138) );
  AOI222_X1 U5116 ( .A1(n5263), .A2(n6182), .B1(n4141), .B2(n6168), .C1(n6183), 
        .C2(n5864), .ZN(n4143) );
  NAND2_X1 U5117 ( .A1(n6218), .A2(REIP_REG_21__SCAN_IN), .ZN(n5267) );
  INV_X1 U5118 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5829) );
  OR2_X1 U5119 ( .A1(n6174), .A2(n5829), .ZN(n4142) );
  NAND3_X1 U5120 ( .A1(n4143), .A2(n5267), .A3(n4142), .ZN(U2965) );
  NOR2_X1 U5121 ( .A1(n4154), .A2(n4153), .ZN(n4149) );
  NAND2_X1 U5122 ( .A1(n4149), .A2(n6484), .ZN(n4163) );
  INV_X1 U5123 ( .A(n4163), .ZN(n4146) );
  INV_X1 U5124 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n6606) );
  NAND2_X1 U5125 ( .A1(n6343), .A2(n6765), .ZN(n5950) );
  OAI211_X1 U5126 ( .C1(n4146), .C2(n6606), .A(n4229), .B(n5950), .ZN(U2788)
         );
  NAND2_X1 U5127 ( .A1(n4232), .A2(n4147), .ZN(n4151) );
  INV_X1 U5128 ( .A(n4145), .ZN(n4148) );
  OR2_X1 U5129 ( .A1(n4149), .A2(n4148), .ZN(n4150) );
  NAND2_X1 U5130 ( .A1(n4151), .A2(n4150), .ZN(n5948) );
  OR2_X1 U5131 ( .A1(n4958), .A2(n4952), .ZN(n4165) );
  AOI21_X1 U5132 ( .B1(n4165), .B2(n6503), .A(READY_N), .ZN(n6598) );
  OR2_X1 U5133 ( .A1(n5948), .A2(n6598), .ZN(n6465) );
  AND2_X1 U5134 ( .A1(n6465), .A2(n6484), .ZN(n5955) );
  INV_X1 U5135 ( .A(MORE_REG_SCAN_IN), .ZN(n4162) );
  NAND2_X1 U5136 ( .A1(n4152), .A2(n4145), .ZN(n4156) );
  INV_X1 U5137 ( .A(n4153), .ZN(n4155) );
  AOI22_X1 U5138 ( .A1(n4232), .A2(n4156), .B1(n4155), .B2(n4154), .ZN(n4159)
         );
  INV_X1 U5139 ( .A(n4232), .ZN(n4157) );
  NAND2_X1 U5140 ( .A1(n4157), .A2(n4200), .ZN(n4158) );
  AND2_X1 U5141 ( .A1(n4159), .A2(n4158), .ZN(n6463) );
  INV_X1 U5142 ( .A(n6463), .ZN(n4160) );
  NAND2_X1 U5143 ( .A1(n5955), .A2(n4160), .ZN(n4161) );
  OAI21_X1 U5144 ( .B1(n5955), .B2(n4162), .A(n4161), .ZN(U3471) );
  INV_X1 U5145 ( .A(n6594), .ZN(n4166) );
  INV_X1 U5146 ( .A(n5950), .ZN(n5394) );
  OAI21_X1 U5147 ( .B1(n5394), .B2(READREQUEST_REG_SCAN_IN), .A(n4166), .ZN(
        n4164) );
  OAI21_X1 U5148 ( .B1(n4166), .B2(n4165), .A(n4164), .ZN(U3474) );
  INV_X1 U5149 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4170) );
  INV_X1 U5150 ( .A(n4231), .ZN(n6475) );
  NOR2_X1 U5151 ( .A1(n6442), .A2(n6475), .ZN(n4168) );
  NAND2_X1 U5152 ( .A1(n4967), .A2(n6484), .ZN(n4167) );
  NAND2_X1 U5153 ( .A1(n6103), .A2(n4965), .ZN(n4341) );
  NAND2_X1 U5154 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4453) );
  OR2_X1 U5155 ( .A1(n4453), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6105) );
  INV_X2 U5156 ( .A(n6105), .ZN(n6597) );
  AOI22_X1 U5157 ( .A1(DATAO_REG_19__SCAN_IN), .A2(n6120), .B1(n6597), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n4169) );
  OAI21_X1 U5158 ( .B1(n4170), .B2(n4341), .A(n4169), .ZN(U2904) );
  INV_X1 U5159 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4172) );
  AOI22_X1 U5160 ( .A1(DATAO_REG_20__SCAN_IN), .A2(n6120), .B1(n6597), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n4171) );
  OAI21_X1 U5161 ( .B1(n4172), .B2(n4341), .A(n4171), .ZN(U2903) );
  AOI22_X1 U5162 ( .A1(n6597), .A2(UWORD_REG_8__SCAN_IN), .B1(n6120), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4173) );
  OAI21_X1 U5163 ( .B1(n3915), .B2(n4341), .A(n4173), .ZN(U2899) );
  INV_X1 U5164 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U5165 ( .A1(n6597), .A2(UWORD_REG_12__SCAN_IN), .B1(n6120), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4174) );
  OAI21_X1 U5166 ( .B1(n4175), .B2(n4341), .A(n4174), .ZN(U2895) );
  INV_X1 U5167 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4177) );
  AOI22_X1 U5168 ( .A1(n6597), .A2(UWORD_REG_9__SCAN_IN), .B1(n6120), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4176) );
  OAI21_X1 U5169 ( .B1(n4177), .B2(n4341), .A(n4176), .ZN(U2898) );
  INV_X1 U5170 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4179) );
  AOI22_X1 U5171 ( .A1(n6597), .A2(UWORD_REG_10__SCAN_IN), .B1(n6120), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4178) );
  OAI21_X1 U5172 ( .B1(n4179), .B2(n4341), .A(n4178), .ZN(U2897) );
  INV_X1 U5173 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4181) );
  AOI22_X1 U5174 ( .A1(n6597), .A2(UWORD_REG_14__SCAN_IN), .B1(n6120), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4180) );
  OAI21_X1 U5175 ( .B1(n4181), .B2(n4341), .A(n4180), .ZN(U2893) );
  AND2_X1 U5176 ( .A1(n4182), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4185) );
  OAI21_X1 U5177 ( .B1(n4185), .B2(n4184), .A(n4183), .ZN(n6200) );
  NAND3_X1 U5178 ( .A1(n4200), .A2(n6484), .A3(n4232), .ZN(n4195) );
  AND2_X1 U5179 ( .A1(n3026), .A2(n4384), .ZN(n4191) );
  NOR2_X1 U5180 ( .A1(n4187), .A2(n4186), .ZN(n4190) );
  NOR2_X1 U5181 ( .A1(n5291), .A2(n4188), .ZN(n4189) );
  NAND4_X1 U5182 ( .A1(n4192), .A2(n4191), .A3(n4190), .A4(n4189), .ZN(n4293)
         );
  INV_X1 U5183 ( .A(n4293), .ZN(n4193) );
  NAND2_X1 U5184 ( .A1(n4193), .A2(n4303), .ZN(n4194) );
  NAND2_X2 U5185 ( .A1(n4195), .A2(n4194), .ZN(n6094) );
  NAND2_X1 U5186 ( .A1(n6094), .A2(n5291), .ZN(n5533) );
  INV_X1 U5187 ( .A(n4196), .ZN(n4197) );
  AOI21_X1 U5188 ( .B1(n4198), .B2(n6577), .A(n4197), .ZN(n4289) );
  INV_X1 U5189 ( .A(n4289), .ZN(n5002) );
  INV_X1 U5190 ( .A(n5291), .ZN(n5286) );
  OAI222_X1 U5191 ( .A1(n6200), .A2(n5533), .B1(n6094), .B2(n4199), .C1(n5002), 
        .C2(n6090), .ZN(U2859) );
  NAND2_X1 U5192 ( .A1(n4200), .A2(n4232), .ZN(n4206) );
  NAND2_X1 U5193 ( .A1(n4962), .A2(n6503), .ZN(n4201) );
  AOI22_X1 U5194 ( .A1(n6442), .A2(n4967), .B1(n3942), .B2(n4201), .ZN(n4202)
         );
  OR3_X1 U5195 ( .A1(n4232), .A2(READY_N), .A3(n4202), .ZN(n4203) );
  AND4_X1 U5196 ( .A1(n4206), .A2(n4205), .A3(n4204), .A4(n4203), .ZN(n4211)
         );
  OR2_X1 U5197 ( .A1(n6461), .A2(n4147), .ZN(n4414) );
  OR2_X1 U5198 ( .A1(n4232), .A2(n4414), .ZN(n4209) );
  INV_X1 U5199 ( .A(n4216), .ZN(n5944) );
  NAND2_X1 U5200 ( .A1(n5944), .A2(n4207), .ZN(n4208) );
  NAND2_X1 U5201 ( .A1(n4209), .A2(n4208), .ZN(n4295) );
  INV_X1 U5202 ( .A(n4295), .ZN(n4210) );
  OR2_X1 U5203 ( .A1(n6780), .A2(n4453), .ZN(n6566) );
  INV_X1 U5204 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5954) );
  OAI22_X1 U5205 ( .A1(n6448), .A2(n6482), .B1(n6566), .B2(n5954), .ZN(n5942)
         );
  NOR2_X1 U5206 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6569), .ZN(n4382) );
  NOR2_X1 U5207 ( .A1(n5942), .A2(n4382), .ZN(n5941) );
  NOR2_X1 U5208 ( .A1(n4213), .A2(n3044), .ZN(n4215) );
  INV_X1 U5209 ( .A(n3942), .ZN(n4214) );
  AND3_X1 U5210 ( .A1(n4216), .A2(n4215), .A3(n4214), .ZN(n4217) );
  NAND2_X1 U5211 ( .A1(n4218), .A2(n4217), .ZN(n6440) );
  INV_X1 U5212 ( .A(n6440), .ZN(n4224) );
  CLKBUF_X1 U5213 ( .A(n4219), .Z(n5046) );
  CLKBUF_X1 U5214 ( .A(n4220), .Z(n4221) );
  NOR3_X1 U5215 ( .A1(n6437), .A2(n5046), .A3(n4221), .ZN(n4222) );
  AOI21_X1 U5216 ( .B1(n6442), .B2(n3231), .A(n4222), .ZN(n4223) );
  OAI21_X1 U5217 ( .B1(n5731), .B2(n4224), .A(n4223), .ZN(n6443) );
  INV_X1 U5218 ( .A(n6583), .ZN(n5943) );
  INV_X1 U5219 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4225) );
  AOI22_X1 U5220 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4225), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n6246), .ZN(n5040) );
  NOR2_X1 U5221 ( .A1(n6765), .A2(n6577), .ZN(n5039) );
  AOI222_X1 U5222 ( .A1(n6443), .A2(n5943), .B1(n5040), .B2(n5039), .C1(n4226), 
        .C2(n5038), .ZN(n4228) );
  INV_X1 U5223 ( .A(n5038), .ZN(n6571) );
  NOR2_X1 U5224 ( .A1(n3507), .A2(n6571), .ZN(n6576) );
  OAI21_X1 U5225 ( .B1(n5941), .B2(n6576), .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), 
        .ZN(n4227) );
  OAI21_X1 U5226 ( .B1(n5941), .B2(n4228), .A(n4227), .ZN(U3460) );
  NOR2_X1 U5227 ( .A1(n4229), .A2(READY_N), .ZN(n4234) );
  NAND2_X1 U5228 ( .A1(n4234), .A2(n4968), .ZN(n4297) );
  INV_X1 U5229 ( .A(DATAI_7_), .ZN(n4230) );
  OR2_X1 U5230 ( .A1(n4297), .A2(n4230), .ZN(n4260) );
  OR3_X1 U5231 ( .A1(n4232), .A2(n6482), .A3(n4231), .ZN(n4233) );
  INV_X2 U5232 ( .A(n4233), .ZN(n6148) );
  OR2_X1 U5233 ( .A1(n4234), .A2(n6148), .ZN(n6151) );
  AOI22_X1 U5234 ( .A1(n6148), .A2(EAX_REG_7__SCAN_IN), .B1(n6145), .B2(
        LWORD_REG_7__SCAN_IN), .ZN(n4235) );
  NAND2_X1 U5235 ( .A1(n4260), .A2(n4235), .ZN(U2946) );
  INV_X1 U5236 ( .A(n4297), .ZN(n6149) );
  NAND2_X1 U5237 ( .A1(n6149), .A2(DATAI_8_), .ZN(n4266) );
  AOI22_X1 U5238 ( .A1(n6148), .A2(EAX_REG_8__SCAN_IN), .B1(n6145), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n4236) );
  NAND2_X1 U5239 ( .A1(n4266), .A2(n4236), .ZN(U2947) );
  NAND2_X1 U5240 ( .A1(n6149), .A2(DATAI_3_), .ZN(n4250) );
  AOI22_X1 U5241 ( .A1(n6148), .A2(EAX_REG_3__SCAN_IN), .B1(n6145), .B2(
        LWORD_REG_3__SCAN_IN), .ZN(n4237) );
  NAND2_X1 U5242 ( .A1(n4250), .A2(n4237), .ZN(U2942) );
  INV_X1 U5243 ( .A(DATAI_6_), .ZN(n4698) );
  OR2_X1 U5244 ( .A1(n4297), .A2(n4698), .ZN(n4252) );
  AOI22_X1 U5245 ( .A1(n6148), .A2(EAX_REG_6__SCAN_IN), .B1(n6145), .B2(
        LWORD_REG_6__SCAN_IN), .ZN(n4238) );
  NAND2_X1 U5246 ( .A1(n4252), .A2(n4238), .ZN(U2945) );
  INV_X1 U5247 ( .A(DATAI_9_), .ZN(n4924) );
  OR2_X1 U5248 ( .A1(n4297), .A2(n4924), .ZN(n4254) );
  AOI22_X1 U5249 ( .A1(n6148), .A2(EAX_REG_9__SCAN_IN), .B1(n6145), .B2(
        LWORD_REG_9__SCAN_IN), .ZN(n4239) );
  NAND2_X1 U5250 ( .A1(n4254), .A2(n4239), .ZN(U2948) );
  NAND2_X1 U5251 ( .A1(n6149), .A2(DATAI_11_), .ZN(n4248) );
  AOI22_X1 U5252 ( .A1(n6148), .A2(EAX_REG_11__SCAN_IN), .B1(n6145), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n4240) );
  NAND2_X1 U5253 ( .A1(n4248), .A2(n4240), .ZN(U2950) );
  INV_X1 U5254 ( .A(DATAI_1_), .ZN(n4300) );
  OR2_X1 U5255 ( .A1(n4297), .A2(n4300), .ZN(n4264) );
  AOI22_X1 U5256 ( .A1(n6148), .A2(EAX_REG_1__SCAN_IN), .B1(n6145), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n4241) );
  NAND2_X1 U5257 ( .A1(n4264), .A2(n4241), .ZN(U2940) );
  INV_X1 U5258 ( .A(DATAI_5_), .ZN(n4242) );
  OR2_X1 U5259 ( .A1(n4297), .A2(n4242), .ZN(n4268) );
  AOI22_X1 U5260 ( .A1(n6148), .A2(EAX_REG_5__SCAN_IN), .B1(n6145), .B2(
        LWORD_REG_5__SCAN_IN), .ZN(n4243) );
  NAND2_X1 U5261 ( .A1(n4268), .A2(n4243), .ZN(U2944) );
  INV_X1 U5262 ( .A(DATAI_4_), .ZN(n4367) );
  OR2_X1 U5263 ( .A1(n4297), .A2(n4367), .ZN(n4258) );
  AOI22_X1 U5264 ( .A1(n6148), .A2(EAX_REG_4__SCAN_IN), .B1(n6145), .B2(
        LWORD_REG_4__SCAN_IN), .ZN(n4244) );
  NAND2_X1 U5265 ( .A1(n4258), .A2(n4244), .ZN(U2943) );
  INV_X1 U5266 ( .A(DATAI_2_), .ZN(n4482) );
  OR2_X1 U5267 ( .A1(n4297), .A2(n4482), .ZN(n4262) );
  AOI22_X1 U5268 ( .A1(n6148), .A2(EAX_REG_2__SCAN_IN), .B1(n6145), .B2(
        LWORD_REG_2__SCAN_IN), .ZN(n4245) );
  NAND2_X1 U5269 ( .A1(n4262), .A2(n4245), .ZN(U2941) );
  INV_X1 U5270 ( .A(DATAI_0_), .ZN(n4481) );
  OR2_X1 U5271 ( .A1(n4297), .A2(n4481), .ZN(n4256) );
  INV_X2 U5272 ( .A(n6151), .ZN(n6145) );
  AOI22_X1 U5273 ( .A1(n6148), .A2(EAX_REG_0__SCAN_IN), .B1(n6145), .B2(
        LWORD_REG_0__SCAN_IN), .ZN(n4246) );
  NAND2_X1 U5274 ( .A1(n4256), .A2(n4246), .ZN(U2939) );
  AOI22_X1 U5275 ( .A1(n6148), .A2(EAX_REG_27__SCAN_IN), .B1(n6145), .B2(
        UWORD_REG_11__SCAN_IN), .ZN(n4247) );
  NAND2_X1 U5276 ( .A1(n4248), .A2(n4247), .ZN(U2935) );
  AOI22_X1 U5277 ( .A1(n6148), .A2(EAX_REG_19__SCAN_IN), .B1(n6145), .B2(
        UWORD_REG_3__SCAN_IN), .ZN(n4249) );
  NAND2_X1 U5278 ( .A1(n4250), .A2(n4249), .ZN(U2927) );
  AOI22_X1 U5279 ( .A1(n6148), .A2(EAX_REG_22__SCAN_IN), .B1(n6145), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n4251) );
  NAND2_X1 U5280 ( .A1(n4252), .A2(n4251), .ZN(U2930) );
  AOI22_X1 U5281 ( .A1(n6148), .A2(EAX_REG_25__SCAN_IN), .B1(n6145), .B2(
        UWORD_REG_9__SCAN_IN), .ZN(n4253) );
  NAND2_X1 U5282 ( .A1(n4254), .A2(n4253), .ZN(U2933) );
  AOI22_X1 U5283 ( .A1(n6148), .A2(EAX_REG_16__SCAN_IN), .B1(n6145), .B2(
        UWORD_REG_0__SCAN_IN), .ZN(n4255) );
  NAND2_X1 U5284 ( .A1(n4256), .A2(n4255), .ZN(U2924) );
  AOI22_X1 U5285 ( .A1(n6148), .A2(EAX_REG_20__SCAN_IN), .B1(n6145), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n4257) );
  NAND2_X1 U5286 ( .A1(n4258), .A2(n4257), .ZN(U2928) );
  AOI22_X1 U5287 ( .A1(n6148), .A2(EAX_REG_23__SCAN_IN), .B1(n6145), .B2(
        UWORD_REG_7__SCAN_IN), .ZN(n4259) );
  NAND2_X1 U5288 ( .A1(n4260), .A2(n4259), .ZN(U2931) );
  AOI22_X1 U5289 ( .A1(n6148), .A2(EAX_REG_18__SCAN_IN), .B1(n6145), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n4261) );
  NAND2_X1 U5290 ( .A1(n4262), .A2(n4261), .ZN(U2926) );
  AOI22_X1 U5291 ( .A1(n6148), .A2(EAX_REG_17__SCAN_IN), .B1(n6145), .B2(
        UWORD_REG_1__SCAN_IN), .ZN(n4263) );
  NAND2_X1 U5292 ( .A1(n4264), .A2(n4263), .ZN(U2925) );
  AOI22_X1 U5293 ( .A1(n6148), .A2(EAX_REG_24__SCAN_IN), .B1(n6145), .B2(
        UWORD_REG_8__SCAN_IN), .ZN(n4265) );
  NAND2_X1 U5294 ( .A1(n4266), .A2(n4265), .ZN(U2932) );
  AOI22_X1 U5295 ( .A1(n6148), .A2(EAX_REG_21__SCAN_IN), .B1(n6145), .B2(
        UWORD_REG_5__SCAN_IN), .ZN(n4267) );
  NAND2_X1 U5296 ( .A1(n4268), .A2(n4267), .ZN(U2929) );
  INV_X1 U5297 ( .A(n4269), .ZN(n4272) );
  NAND2_X1 U5298 ( .A1(n4270), .A2(n4269), .ZN(n4353) );
  INV_X1 U5299 ( .A(n4353), .ZN(n4271) );
  AOI21_X1 U5300 ( .B1(n4272), .B2(n4278), .A(n4271), .ZN(n6184) );
  INV_X1 U5301 ( .A(n6184), .ZN(n5501) );
  XNOR2_X1 U5302 ( .A(n4321), .B(n4273), .ZN(n6239) );
  INV_X1 U5303 ( .A(n6094), .ZN(n5505) );
  AOI22_X1 U5304 ( .A1(n6081), .A2(n6239), .B1(n5505), .B2(EBX_REG_2__SCAN_IN), 
        .ZN(n4274) );
  OAI21_X1 U5305 ( .B1(n5501), .B2(n5533), .A(n4274), .ZN(U2857) );
  OAI21_X1 U5306 ( .B1(n4277), .B2(n4276), .A(n4275), .ZN(n4314) );
  OAI21_X1 U5307 ( .B1(n4280), .B2(n4279), .A(n4278), .ZN(n4305) );
  INV_X1 U5308 ( .A(n4305), .ZN(n4976) );
  NAND2_X1 U5309 ( .A1(n4976), .A2(n6183), .ZN(n4284) );
  INV_X1 U5310 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4282) );
  AND2_X1 U5311 ( .A1(n6218), .A2(REIP_REG_1__SCAN_IN), .ZN(n4309) );
  AND2_X1 U5312 ( .A1(n6196), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4281)
         );
  AOI211_X1 U5313 ( .C1(n6168), .C2(n4282), .A(n4309), .B(n4281), .ZN(n4283)
         );
  OAI211_X1 U5314 ( .C1(n4314), .C2(n6190), .A(n4284), .B(n4283), .ZN(U2985)
         );
  INV_X1 U5315 ( .A(n4308), .ZN(n4286) );
  INV_X1 U5316 ( .A(n4285), .ZN(n5936) );
  AOI211_X1 U5317 ( .C1(n6193), .C2(n6247), .A(n4286), .B(n5936), .ZN(n4292)
         );
  INV_X1 U5318 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6586) );
  NOR2_X1 U5319 ( .A1(n6242), .A2(n6586), .ZN(n6192) );
  NAND2_X1 U5320 ( .A1(n6577), .A2(n4287), .ZN(n4307) );
  INV_X1 U5321 ( .A(n4307), .ZN(n4288) );
  AOI211_X1 U5322 ( .C1(n6240), .C2(n4289), .A(n6192), .B(n4288), .ZN(n4291)
         );
  NAND3_X1 U5323 ( .A1(n6193), .A2(n6247), .A3(n6189), .ZN(n4290) );
  OAI211_X1 U5324 ( .C1(n4292), .C2(n6577), .A(n4291), .B(n4290), .ZN(U3018)
         );
  NOR2_X1 U5325 ( .A1(n4293), .A2(n4147), .ZN(n4294) );
  AOI21_X1 U5326 ( .B1(n4295), .B2(n6484), .A(n4294), .ZN(n4296) );
  NAND2_X1 U5327 ( .A1(n3196), .A2(n5291), .ZN(n4298) );
  INV_X1 U5328 ( .A(n4298), .ZN(n4299) );
  INV_X1 U5329 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6130) );
  OAI222_X1 U5330 ( .A1(n4305), .A2(n5857), .B1(n5010), .B2(n4300), .C1(n5293), 
        .C2(n6130), .ZN(U2890) );
  OAI21_X1 U5331 ( .B1(n4301), .B2(n4303), .A(n4302), .ZN(n4311) );
  AOI22_X1 U5332 ( .A1(n6081), .A2(n4311), .B1(n5505), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n4304) );
  OAI21_X1 U5333 ( .B1(n4305), .B2(n6085), .A(n4304), .ZN(U2858) );
  NAND3_X1 U5334 ( .A1(n6213), .A2(n4306), .A3(n6246), .ZN(n4313) );
  AOI21_X1 U5335 ( .B1(n4308), .B2(n4307), .A(n6246), .ZN(n4310) );
  AOI211_X1 U5336 ( .C1(n6240), .C2(n4311), .A(n4310), .B(n4309), .ZN(n4312)
         );
  OAI211_X1 U5337 ( .C1(n6203), .C2(n4314), .A(n4313), .B(n4312), .ZN(U3017)
         );
  XNOR2_X1 U5338 ( .A(n4315), .B(n4316), .ZN(n4362) );
  INV_X1 U5339 ( .A(n4691), .ZN(n6238) );
  AOI21_X1 U5340 ( .B1(n4318), .B2(n6237), .A(n4317), .ZN(n6253) );
  OAI21_X1 U5341 ( .B1(n6236), .B2(n6238), .A(n6253), .ZN(n5051) );
  OAI21_X1 U5342 ( .B1(n4321), .B2(n4320), .A(n4319), .ZN(n4322) );
  NAND2_X1 U5343 ( .A1(n4322), .A2(n4344), .ZN(n4355) );
  NAND2_X1 U5344 ( .A1(n6218), .A2(REIP_REG_3__SCAN_IN), .ZN(n4357) );
  OAI21_X1 U5345 ( .B1(n6229), .B2(n4355), .A(n4357), .ZN(n4324) );
  OAI21_X1 U5346 ( .B1(n6237), .B2(n6245), .A(n6236), .ZN(n4535) );
  NAND2_X1 U5347 ( .A1(n6238), .A2(n4535), .ZN(n5053) );
  NOR2_X1 U5348 ( .A1(n5053), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4323)
         );
  AOI211_X1 U5349 ( .C1(n5051), .C2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n4324), 
        .B(n4323), .ZN(n4325) );
  OAI21_X1 U5350 ( .B1(n4362), .B2(n6203), .A(n4325), .ZN(U3015) );
  INV_X1 U5351 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4327) );
  AOI22_X1 U5352 ( .A1(n6597), .A2(UWORD_REG_0__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4326) );
  OAI21_X1 U5353 ( .B1(n4327), .B2(n4341), .A(n4326), .ZN(U2907) );
  INV_X1 U5354 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4329) );
  AOI22_X1 U5355 ( .A1(n6597), .A2(UWORD_REG_5__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4328) );
  OAI21_X1 U5356 ( .B1(n4329), .B2(n4341), .A(n4328), .ZN(U2902) );
  INV_X1 U5357 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4331) );
  AOI22_X1 U5358 ( .A1(n6597), .A2(UWORD_REG_6__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4330) );
  OAI21_X1 U5359 ( .B1(n4331), .B2(n4341), .A(n4330), .ZN(U2901) );
  INV_X1 U5360 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4333) );
  AOI22_X1 U5361 ( .A1(n6597), .A2(UWORD_REG_11__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4332) );
  OAI21_X1 U5362 ( .B1(n4333), .B2(n4341), .A(n4332), .ZN(U2896) );
  INV_X1 U5363 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4335) );
  AOI22_X1 U5364 ( .A1(n6597), .A2(UWORD_REG_1__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4334) );
  OAI21_X1 U5365 ( .B1(n4335), .B2(n4341), .A(n4334), .ZN(U2906) );
  INV_X1 U5366 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4337) );
  AOI22_X1 U5367 ( .A1(n6597), .A2(UWORD_REG_2__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4336) );
  OAI21_X1 U5368 ( .B1(n4337), .B2(n4341), .A(n4336), .ZN(U2905) );
  INV_X1 U5369 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4339) );
  AOI22_X1 U5370 ( .A1(n6597), .A2(UWORD_REG_7__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4338) );
  OAI21_X1 U5371 ( .B1(n4339), .B2(n4341), .A(n4338), .ZN(U2900) );
  INV_X1 U5372 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4342) );
  AOI22_X1 U5373 ( .A1(n6597), .A2(UWORD_REG_13__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4340) );
  OAI21_X1 U5374 ( .B1(n4342), .B2(n4341), .A(n4340), .ZN(U2894) );
  AOI21_X1 U5375 ( .B1(n4343), .B2(n4351), .A(n4348), .ZN(n5062) );
  INV_X1 U5376 ( .A(n5062), .ZN(n6073) );
  AOI21_X1 U5377 ( .B1(n4345), .B2(n4344), .A(n4364), .ZN(n6063) );
  AOI22_X1 U5378 ( .A1(n6081), .A2(n6063), .B1(n5505), .B2(EBX_REG_4__SCAN_IN), 
        .ZN(n4346) );
  OAI21_X1 U5379 ( .B1(n6073), .B2(n6085), .A(n4346), .ZN(U2855) );
  OR2_X1 U5380 ( .A1(n4348), .A2(n4347), .ZN(n4349) );
  AND2_X1 U5381 ( .A1(n4678), .A2(n4349), .ZN(n6170) );
  INV_X1 U5382 ( .A(n6170), .ZN(n4366) );
  AOI22_X1 U5383 ( .A1(n5557), .A2(DATAI_5_), .B1(n6608), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n4350) );
  OAI21_X1 U5384 ( .B1(n4366), .B2(n5857), .A(n4350), .ZN(U2886) );
  INV_X1 U5385 ( .A(n4351), .ZN(n4352) );
  AOI21_X1 U5386 ( .B1(n4354), .B2(n4353), .A(n4352), .ZN(n5476) );
  INV_X1 U5387 ( .A(n5476), .ZN(n4363) );
  INV_X1 U5388 ( .A(n4355), .ZN(n5477) );
  AOI22_X1 U5389 ( .A1(n6081), .A2(n5477), .B1(n5505), .B2(EBX_REG_3__SCAN_IN), 
        .ZN(n4356) );
  OAI21_X1 U5390 ( .B1(n4363), .B2(n5533), .A(n4356), .ZN(U2856) );
  NAND2_X1 U5391 ( .A1(n6168), .A2(n5478), .ZN(n4358) );
  OAI211_X1 U5392 ( .C1(n6174), .C2(n4359), .A(n4358), .B(n4357), .ZN(n4360)
         );
  AOI21_X1 U5393 ( .B1(n5476), .B2(n6183), .A(n4360), .ZN(n4361) );
  OAI21_X1 U5394 ( .B1(n4362), .B2(n6190), .A(n4361), .ZN(U2983) );
  INV_X1 U5395 ( .A(DATAI_3_), .ZN(n6742) );
  INV_X1 U5396 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6127) );
  OAI222_X1 U5397 ( .A1(n4363), .A2(n5857), .B1(n5010), .B2(n6742), .C1(n5293), 
        .C2(n6127), .ZN(U2888) );
  INV_X1 U5398 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4365) );
  OAI21_X1 U5399 ( .B1(n4364), .B2(n3035), .A(n4534), .ZN(n6047) );
  OAI222_X1 U5400 ( .A1(n4366), .A2(n5533), .B1(n6094), .B2(n4365), .C1(n6090), 
        .C2(n6047), .ZN(U2854) );
  INV_X1 U5401 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6759) );
  OAI222_X1 U5402 ( .A1(n5857), .A2(n6073), .B1(n5293), .B2(n6759), .C1(n5010), 
        .C2(n4367), .ZN(U2887) );
  NAND3_X1 U5403 ( .A1(n6458), .A2(n6452), .A3(n6445), .ZN(n4706) );
  NOR2_X1 U5404 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4706), .ZN(n4600)
         );
  INV_X1 U5405 ( .A(n4600), .ZN(n4370) );
  INV_X1 U5406 ( .A(n4380), .ZN(n4368) );
  NOR2_X1 U5407 ( .A1(n4368), .A2(n6486), .ZN(n6290) );
  INV_X1 U5408 ( .A(n4369), .ZN(n4507) );
  INV_X1 U5409 ( .A(n5749), .ZN(n6289) );
  NOR2_X1 U5410 ( .A1(n4507), .A2(n6289), .ZN(n4381) );
  NOR2_X1 U5411 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6600) );
  INV_X1 U5412 ( .A(n6600), .ZN(n6493) );
  OAI21_X1 U5413 ( .B1(n4381), .B2(n6486), .A(n4582), .ZN(n4545) );
  AOI211_X1 U5414 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4370), .A(n6290), .B(
        n4545), .ZN(n4378) );
  AND2_X1 U5415 ( .A1(n5733), .A2(n4614), .ZN(n4372) );
  AND2_X1 U5416 ( .A1(n4372), .A2(n5742), .ZN(n4483) );
  OR3_X1 U5417 ( .A1(n5733), .A2(n4506), .A3(n4614), .ZN(n4465) );
  INV_X1 U5418 ( .A(n4806), .ZN(n4373) );
  NOR3_X1 U5419 ( .A1(n4704), .A2(n4373), .A3(n6382), .ZN(n4376) );
  AND2_X1 U5420 ( .A1(n6343), .A2(n6487), .ZN(n4616) );
  INV_X1 U5421 ( .A(n5731), .ZN(n4457) );
  OR2_X1 U5422 ( .A1(n5491), .A2(n4457), .ZN(n4700) );
  OAI22_X1 U5423 ( .A1(n4376), .A2(n4616), .B1(n5747), .B2(n4700), .ZN(n4377)
         );
  INV_X1 U5424 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4388) );
  INV_X1 U5425 ( .A(DATAI_19_), .ZN(n4379) );
  NOR2_X1 U5426 ( .A1(n6199), .A2(n4379), .ZN(n6404) );
  NAND2_X1 U5427 ( .A1(n6183), .A2(DATAI_27_), .ZN(n4860) );
  NAND2_X1 U5428 ( .A1(DATAI_3_), .A2(n4582), .ZN(n6407) );
  INV_X1 U5429 ( .A(n6407), .ZN(n6314) );
  NAND2_X1 U5430 ( .A1(n5740), .A2(n6343), .ZN(n6292) );
  NOR2_X1 U5431 ( .A1(n4380), .A2(n6486), .ZN(n4639) );
  INV_X1 U5432 ( .A(n4639), .ZN(n6299) );
  INV_X1 U5433 ( .A(n4381), .ZN(n4547) );
  OAI22_X1 U5434 ( .A1(n6292), .A2(n4700), .B1(n6299), .B2(n4547), .ZN(n4601)
         );
  INV_X1 U5435 ( .A(n4382), .ZN(n6567) );
  NOR2_X1 U5436 ( .A1(n4583), .A2(n4384), .ZN(n6402) );
  AOI22_X1 U5437 ( .A1(n6314), .A2(n4601), .B1(n6402), .B2(n4600), .ZN(n4385)
         );
  OAI21_X1 U5438 ( .B1(n4860), .B2(n4806), .A(n4385), .ZN(n4386) );
  AOI21_X1 U5439 ( .B1(n6404), .B2(n4704), .A(n4386), .ZN(n4387) );
  OAI21_X1 U5440 ( .B1(n4606), .B2(n4388), .A(n4387), .ZN(U3023) );
  INV_X1 U5441 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4394) );
  INV_X1 U5442 ( .A(DATAI_18_), .ZN(n4389) );
  NOR2_X1 U5443 ( .A1(n6199), .A2(n4389), .ZN(n6398) );
  INV_X1 U5444 ( .A(DATAI_26_), .ZN(n4390) );
  NOR2_X1 U5445 ( .A1(n6199), .A2(n4390), .ZN(n6397) );
  INV_X1 U5446 ( .A(n6397), .ZN(n4890) );
  NAND2_X1 U5447 ( .A1(DATAI_2_), .A2(n4582), .ZN(n6401) );
  INV_X1 U5448 ( .A(n6401), .ZN(n6310) );
  NOR2_X1 U5449 ( .A1(n3194), .A2(n4583), .ZN(n6396) );
  AOI22_X1 U5450 ( .A1(n6310), .A2(n4601), .B1(n6396), .B2(n4600), .ZN(n4391)
         );
  OAI21_X1 U5451 ( .B1(n4890), .B2(n4806), .A(n4391), .ZN(n4392) );
  AOI21_X1 U5452 ( .B1(n6398), .B2(n4704), .A(n4392), .ZN(n4393) );
  OAI21_X1 U5453 ( .B1(n4606), .B2(n4394), .A(n4393), .ZN(U3022) );
  NAND2_X1 U5454 ( .A1(n6183), .A2(DATAI_23_), .ZN(n6337) );
  INV_X1 U5455 ( .A(n6337), .ZN(n6428) );
  INV_X1 U5456 ( .A(DATAI_31_), .ZN(n4395) );
  NOR2_X1 U5457 ( .A1(n6199), .A2(n4395), .ZN(n6431) );
  INV_X1 U5458 ( .A(n6431), .ZN(n4857) );
  NAND2_X1 U5459 ( .A1(DATAI_7_), .A2(n4582), .ZN(n6435) );
  INV_X1 U5460 ( .A(n6435), .ZN(n6332) );
  NOR2_X1 U5461 ( .A1(n4583), .A2(n5286), .ZN(n6427) );
  AOI22_X1 U5462 ( .A1(n6332), .A2(n4601), .B1(n6427), .B2(n4600), .ZN(n4396)
         );
  OAI21_X1 U5463 ( .B1(n4857), .B2(n4806), .A(n4396), .ZN(n4397) );
  AOI21_X1 U5464 ( .B1(n6428), .B2(n4704), .A(n4397), .ZN(n4398) );
  OAI21_X1 U5465 ( .B1(n4606), .B2(n4399), .A(n4398), .ZN(U3027) );
  INV_X1 U5466 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4406) );
  INV_X1 U5467 ( .A(DATAI_17_), .ZN(n4400) );
  NOR2_X1 U5468 ( .A1(n6199), .A2(n4400), .ZN(n6391) );
  INV_X1 U5469 ( .A(DATAI_25_), .ZN(n4401) );
  NOR2_X1 U5470 ( .A1(n6199), .A2(n4401), .ZN(n6392) );
  INV_X1 U5471 ( .A(n6392), .ZN(n4884) );
  NAND2_X1 U5472 ( .A1(DATAI_1_), .A2(n4582), .ZN(n6395) );
  INV_X1 U5473 ( .A(n6395), .ZN(n6306) );
  NOR2_X1 U5474 ( .A1(n4583), .A2(n4402), .ZN(n6390) );
  AOI22_X1 U5475 ( .A1(n6306), .A2(n4601), .B1(n6390), .B2(n4600), .ZN(n4403)
         );
  OAI21_X1 U5476 ( .B1(n4884), .B2(n4806), .A(n4403), .ZN(n4404) );
  AOI21_X1 U5477 ( .B1(n6391), .B2(n4704), .A(n4404), .ZN(n4405) );
  OAI21_X1 U5478 ( .B1(n4606), .B2(n4406), .A(n4405), .ZN(U3021) );
  INV_X1 U5479 ( .A(DATAI_16_), .ZN(n4407) );
  NOR2_X1 U5480 ( .A1(n6199), .A2(n4407), .ZN(n6377) );
  INV_X1 U5481 ( .A(DATAI_24_), .ZN(n4408) );
  NOR2_X1 U5482 ( .A1(n6199), .A2(n4408), .ZN(n6386) );
  INV_X1 U5483 ( .A(n6386), .ZN(n4873) );
  NAND2_X1 U5484 ( .A1(DATAI_0_), .A2(n4582), .ZN(n6389) );
  INV_X1 U5485 ( .A(n6389), .ZN(n6293) );
  NOR2_X1 U5486 ( .A1(n4583), .A2(n4409), .ZN(n6376) );
  AOI22_X1 U5487 ( .A1(n6293), .A2(n4601), .B1(n6376), .B2(n4600), .ZN(n4410)
         );
  OAI21_X1 U5488 ( .B1(n4873), .B2(n4806), .A(n4410), .ZN(n4411) );
  AOI21_X1 U5489 ( .B1(n6377), .B2(n4704), .A(n4411), .ZN(n4412) );
  OAI21_X1 U5490 ( .B1(n4606), .B2(n4413), .A(n4412), .ZN(U3020) );
  NAND2_X1 U5491 ( .A1(n5747), .A2(n6440), .ZN(n4428) );
  NAND2_X1 U5492 ( .A1(n4415), .A2(n4414), .ZN(n4429) );
  MUX2_X1 U5493 ( .A(n4418), .B(n6575), .S(n5046), .Z(n4417) );
  CLKBUF_X1 U5494 ( .A(n4416), .Z(n4442) );
  NOR2_X1 U5495 ( .A1(n4417), .A2(n4442), .ZN(n4426) );
  INV_X1 U5496 ( .A(n4418), .ZN(n4419) );
  OAI211_X1 U5497 ( .C1(n5046), .C2(n6575), .A(n4420), .B(n4419), .ZN(n6572)
         );
  AND2_X1 U5498 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4422) );
  INV_X1 U5499 ( .A(n4422), .ZN(n4421) );
  MUX2_X1 U5500 ( .A(n4422), .B(n4421), .S(n6575), .Z(n4423) );
  NAND2_X1 U5501 ( .A1(n6442), .A2(n4423), .ZN(n4424) );
  OAI21_X1 U5502 ( .B1(n4431), .B2(n6572), .A(n4424), .ZN(n4425) );
  AOI21_X1 U5503 ( .B1(n4429), .B2(n4426), .A(n4425), .ZN(n4427) );
  NAND2_X1 U5504 ( .A1(n4428), .A2(n4427), .ZN(n6570) );
  INV_X1 U5505 ( .A(n6448), .ZN(n4437) );
  MUX2_X1 U5506 ( .A(n6575), .B(n6570), .S(n4437), .Z(n6459) );
  XNOR2_X1 U5507 ( .A(n5046), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4430)
         );
  NAND2_X1 U5508 ( .A1(n4429), .A2(n4430), .ZN(n4435) );
  XNOR2_X1 U5509 ( .A(n3231), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4433)
         );
  NOR2_X1 U5510 ( .A1(n4431), .A2(n4430), .ZN(n4432) );
  AOI21_X1 U5511 ( .B1(n6442), .B2(n4433), .A(n4432), .ZN(n4434) );
  NAND2_X1 U5512 ( .A1(n4435), .A2(n4434), .ZN(n4436) );
  AOI21_X1 U5513 ( .B1(n5491), .B2(n6440), .A(n4436), .ZN(n5042) );
  NAND2_X1 U5514 ( .A1(n5042), .A2(n4437), .ZN(n4439) );
  NAND2_X1 U5515 ( .A1(n6448), .A2(n3237), .ZN(n4438) );
  NAND2_X1 U5516 ( .A1(n4439), .A2(n4438), .ZN(n6450) );
  INV_X1 U5517 ( .A(n6450), .ZN(n4440) );
  NAND3_X1 U5518 ( .A1(n6459), .A2(n4440), .A3(n6765), .ZN(n4444) );
  NAND2_X1 U5519 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5954), .ZN(n4449) );
  INV_X1 U5520 ( .A(n4449), .ZN(n4441) );
  NAND2_X1 U5521 ( .A1(n4442), .A2(n4441), .ZN(n4443) );
  AND2_X1 U5522 ( .A1(n4444), .A2(n4443), .ZN(n6469) );
  NOR2_X1 U5523 ( .A1(n6469), .A2(n4221), .ZN(n4454) );
  INV_X1 U5524 ( .A(n6295), .ZN(n4509) );
  OR2_X1 U5525 ( .A1(n4445), .A2(n4509), .ZN(n4446) );
  XNOR2_X1 U5526 ( .A(n4446), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6061)
         );
  NAND2_X1 U5527 ( .A1(n6061), .A2(n5944), .ZN(n4448) );
  NAND2_X1 U5528 ( .A1(n6448), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4447) );
  AOI21_X1 U5529 ( .B1(n4448), .B2(n4447), .A(STATE2_REG_1__SCAN_IN), .ZN(
        n4451) );
  NOR2_X1 U5530 ( .A1(n5946), .A2(n4449), .ZN(n4450) );
  OR2_X1 U5531 ( .A1(n4451), .A2(n4450), .ZN(n6467) );
  NOR3_X1 U5532 ( .A1(n4454), .A2(n6467), .A3(FLUSH_REG_SCAN_IN), .ZN(n4452)
         );
  INV_X1 U5533 ( .A(n4582), .ZN(n4511) );
  OAI21_X1 U5534 ( .B1(n4452), .B2(n6566), .A(n4511), .ZN(n6254) );
  NOR3_X1 U5535 ( .A1(n4454), .A2(n4453), .A3(n6467), .ZN(n6479) );
  INV_X1 U5536 ( .A(n6441), .ZN(n6373) );
  AND2_X1 U5537 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6569), .ZN(n5741) );
  OAI22_X1 U5538 ( .A1(n3032), .A2(n6382), .B1(n6373), .B2(n5741), .ZN(n4455)
         );
  OAI21_X1 U5539 ( .B1(n6479), .B2(n4455), .A(n6254), .ZN(n4456) );
  OAI21_X1 U5540 ( .B1(n6254), .B2(n6256), .A(n4456), .ZN(U3465) );
  AOI21_X1 U5541 ( .B1(n6256), .B2(STATE2_REG_3__SCAN_IN), .A(n4511), .ZN(
        n6263) );
  AND2_X1 U5542 ( .A1(n5747), .A2(n6441), .ZN(n4863) );
  AND2_X1 U5543 ( .A1(n5491), .A2(n4457), .ZN(n4644) );
  INV_X1 U5544 ( .A(n4804), .ZN(n4458) );
  AOI21_X1 U5545 ( .B1(n4863), .B2(n4644), .A(n4458), .ZN(n4462) );
  INV_X1 U5546 ( .A(n4465), .ZN(n4459) );
  INV_X1 U5547 ( .A(n4616), .ZN(n6297) );
  OAI21_X1 U5548 ( .B1(n4459), .B2(n6199), .A(n6297), .ZN(n4460) );
  AOI22_X1 U5549 ( .A1(n4462), .A2(n4460), .B1(n4638), .B2(n6382), .ZN(n4461)
         );
  NAND2_X1 U5550 ( .A1(n6263), .A2(n4461), .ZN(n4810) );
  INV_X1 U5551 ( .A(n4462), .ZN(n4464) );
  AOI22_X1 U5552 ( .A1(n4464), .A2(n6343), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4463), .ZN(n4805) );
  INV_X1 U5553 ( .A(n6396), .ZN(n4752) );
  OAI22_X1 U5554 ( .A1(n6401), .A2(n4805), .B1(n4804), .B2(n4752), .ZN(n4467)
         );
  INV_X1 U5555 ( .A(n6398), .ZN(n6313) );
  OAI22_X1 U5556 ( .A1(n4890), .A2(n4807), .B1(n4806), .B2(n6313), .ZN(n4466)
         );
  AOI211_X1 U5557 ( .C1(n4810), .C2(INSTQUEUE_REG_15__2__SCAN_IN), .A(n4467), 
        .B(n4466), .ZN(n4468) );
  INV_X1 U5558 ( .A(n4468), .ZN(U3142) );
  INV_X1 U5559 ( .A(n6427), .ZN(n4731) );
  OAI22_X1 U5560 ( .A1(n6435), .A2(n4805), .B1(n4804), .B2(n4731), .ZN(n4470)
         );
  OAI22_X1 U5561 ( .A1(n4857), .A2(n4807), .B1(n4806), .B2(n6337), .ZN(n4469)
         );
  AOI211_X1 U5562 ( .C1(n4810), .C2(INSTQUEUE_REG_15__7__SCAN_IN), .A(n4470), 
        .B(n4469), .ZN(n4471) );
  INV_X1 U5563 ( .A(n4471), .ZN(U3147) );
  INV_X1 U5564 ( .A(n6390), .ZN(n4744) );
  OAI22_X1 U5565 ( .A1(n6395), .A2(n4805), .B1(n4804), .B2(n4744), .ZN(n4473)
         );
  INV_X1 U5566 ( .A(n6391), .ZN(n6309) );
  OAI22_X1 U5567 ( .A1(n4884), .A2(n4807), .B1(n4806), .B2(n6309), .ZN(n4472)
         );
  AOI211_X1 U5568 ( .C1(n4810), .C2(INSTQUEUE_REG_15__1__SCAN_IN), .A(n4473), 
        .B(n4472), .ZN(n4474) );
  INV_X1 U5569 ( .A(n4474), .ZN(U3141) );
  INV_X1 U5570 ( .A(n6402), .ZN(n4748) );
  OAI22_X1 U5571 ( .A1(n6407), .A2(n4805), .B1(n4804), .B2(n4748), .ZN(n4476)
         );
  INV_X1 U5572 ( .A(n6404), .ZN(n6317) );
  OAI22_X1 U5573 ( .A1(n4860), .A2(n4807), .B1(n4806), .B2(n6317), .ZN(n4475)
         );
  AOI211_X1 U5574 ( .C1(n4810), .C2(INSTQUEUE_REG_15__3__SCAN_IN), .A(n4476), 
        .B(n4475), .ZN(n4477) );
  INV_X1 U5575 ( .A(n4477), .ZN(U3143) );
  INV_X1 U5576 ( .A(n6376), .ZN(n4740) );
  OAI22_X1 U5577 ( .A1(n6389), .A2(n4805), .B1(n4804), .B2(n4740), .ZN(n4479)
         );
  INV_X1 U5578 ( .A(n6377), .ZN(n6305) );
  OAI22_X1 U5579 ( .A1(n4873), .A2(n4807), .B1(n4806), .B2(n6305), .ZN(n4478)
         );
  AOI211_X1 U5580 ( .C1(n4810), .C2(INSTQUEUE_REG_15__0__SCAN_IN), .A(n4479), 
        .B(n4478), .ZN(n4480) );
  INV_X1 U5581 ( .A(n4480), .ZN(U3140) );
  INV_X1 U5582 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6134) );
  OAI222_X1 U5583 ( .A1(n6200), .A2(n5857), .B1(n5010), .B2(n4481), .C1(n5293), 
        .C2(n6134), .ZN(U2891) );
  INV_X1 U5584 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6773) );
  OAI222_X1 U5585 ( .A1(n5501), .A2(n5857), .B1(n5010), .B2(n4482), .C1(n5293), 
        .C2(n6773), .ZN(U2889) );
  INV_X1 U5586 ( .A(n4483), .ZN(n4699) );
  AND2_X1 U5587 ( .A1(n5733), .A2(n5744), .ZN(n4484) );
  NAND2_X1 U5588 ( .A1(n4484), .A2(n5742), .ZN(n4541) );
  NOR2_X2 U5589 ( .A1(n4541), .A2(n6287), .ZN(n4841) );
  OAI21_X1 U5590 ( .B1(n4782), .B2(n4841), .A(n6297), .ZN(n4485) );
  NOR2_X1 U5591 ( .A1(n5491), .A2(n5731), .ZN(n5748) );
  NAND2_X1 U5592 ( .A1(n5740), .A2(n5748), .ZN(n4727) );
  AOI21_X1 U5593 ( .B1(n4485), .B2(n4727), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4486) );
  NAND3_X1 U5594 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6458), .A3(n6452), .ZN(n4734) );
  NOR2_X1 U5595 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4734), .ZN(n4489)
         );
  OAI21_X1 U5596 ( .B1(n6289), .B2(n6486), .A(n4582), .ZN(n6301) );
  NOR2_X1 U5597 ( .A1(n6290), .A2(n6301), .ZN(n5755) );
  OAI21_X1 U5598 ( .B1(n4486), .B2(n4489), .A(n5755), .ZN(n4836) );
  NAND2_X1 U5599 ( .A1(n4836), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4492) );
  INV_X1 U5600 ( .A(n4727), .ZN(n4488) );
  NOR3_X1 U5601 ( .A1(n6299), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n5749), 
        .ZN(n4487) );
  AOI21_X1 U5602 ( .B1(n4488), .B2(n6343), .A(n4487), .ZN(n4839) );
  INV_X1 U5603 ( .A(n4489), .ZN(n4837) );
  OAI22_X1 U5604 ( .A1(n6435), .A2(n4839), .B1(n4731), .B2(n4837), .ZN(n4490)
         );
  AOI21_X1 U5605 ( .B1(n6428), .B2(n4841), .A(n4490), .ZN(n4491) );
  OAI211_X1 U5606 ( .C1(n4844), .C2(n4857), .A(n4492), .B(n4491), .ZN(U3043)
         );
  NAND2_X1 U5607 ( .A1(n4836), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4495) );
  OAI22_X1 U5608 ( .A1(n6395), .A2(n4839), .B1(n4744), .B2(n4837), .ZN(n4493)
         );
  AOI21_X1 U5609 ( .B1(n6391), .B2(n4841), .A(n4493), .ZN(n4494) );
  OAI211_X1 U5610 ( .C1(n4844), .C2(n4884), .A(n4495), .B(n4494), .ZN(U3037)
         );
  NAND2_X1 U5611 ( .A1(n4836), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4498) );
  OAI22_X1 U5612 ( .A1(n6401), .A2(n4839), .B1(n4752), .B2(n4837), .ZN(n4496)
         );
  AOI21_X1 U5613 ( .B1(n6398), .B2(n4841), .A(n4496), .ZN(n4497) );
  OAI211_X1 U5614 ( .C1(n4844), .C2(n4890), .A(n4498), .B(n4497), .ZN(U3038)
         );
  NAND2_X1 U5615 ( .A1(n4836), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4501) );
  OAI22_X1 U5616 ( .A1(n6407), .A2(n4839), .B1(n4748), .B2(n4837), .ZN(n4499)
         );
  AOI21_X1 U5617 ( .B1(n6404), .B2(n4841), .A(n4499), .ZN(n4500) );
  OAI211_X1 U5618 ( .C1(n4844), .C2(n4860), .A(n4501), .B(n4500), .ZN(U3039)
         );
  NAND2_X1 U5619 ( .A1(n4836), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4504) );
  OAI22_X1 U5620 ( .A1(n6389), .A2(n4839), .B1(n4740), .B2(n4837), .ZN(n4502)
         );
  AOI21_X1 U5621 ( .B1(n6377), .B2(n4841), .A(n4502), .ZN(n4503) );
  OAI211_X1 U5622 ( .C1(n4844), .C2(n4873), .A(n4504), .B(n4503), .ZN(U3036)
         );
  AND2_X1 U5623 ( .A1(n5744), .A2(n6287), .ZN(n4505) );
  OR3_X1 U5624 ( .A1(n5733), .A2(n4506), .A3(n5744), .ZN(n4636) );
  NOR2_X2 U5625 ( .A1(n4636), .A2(n6287), .ZN(n4904) );
  NOR2_X1 U5626 ( .A1(n5740), .A2(n6382), .ZN(n4643) );
  AND2_X1 U5627 ( .A1(n5491), .A2(n5731), .ZN(n4862) );
  NAND2_X1 U5628 ( .A1(n4507), .A2(n5749), .ZN(n4512) );
  INV_X1 U5629 ( .A(n4512), .ZN(n4620) );
  AOI22_X1 U5630 ( .A1(n4643), .A2(n4862), .B1(n4620), .B2(n6290), .ZN(n4826)
         );
  NAND3_X1 U5631 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6445), .ZN(n4866) );
  NOR2_X1 U5632 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4866), .ZN(n4516)
         );
  INV_X1 U5633 ( .A(n4516), .ZN(n4825) );
  OAI22_X1 U5634 ( .A1(n6395), .A2(n4826), .B1(n4744), .B2(n4825), .ZN(n4508)
         );
  AOI21_X1 U5635 ( .B1(n6391), .B2(n4904), .A(n4508), .ZN(n4518) );
  NOR3_X1 U5636 ( .A1(n6429), .A2(n4904), .A3(n6382), .ZN(n4510) );
  INV_X1 U5637 ( .A(n4862), .ZN(n4549) );
  OAI22_X1 U5638 ( .A1(n4510), .A2(n4616), .B1(n4509), .B2(n4549), .ZN(n4515)
         );
  AOI21_X1 U5639 ( .B1(n4512), .B2(STATE2_REG_2__SCAN_IN), .A(n4511), .ZN(
        n4513) );
  INV_X1 U5640 ( .A(n4513), .ZN(n4613) );
  NOR2_X1 U5641 ( .A1(n4639), .A2(n4613), .ZN(n4514) );
  OAI211_X1 U5642 ( .C1(n4516), .C2(n6569), .A(n4515), .B(n4514), .ZN(n4828)
         );
  NAND2_X1 U5643 ( .A1(n4828), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4517)
         );
  OAI211_X1 U5644 ( .C1(n4831), .C2(n4884), .A(n4518), .B(n4517), .ZN(U3117)
         );
  OAI22_X1 U5645 ( .A1(n6407), .A2(n4826), .B1(n4748), .B2(n4825), .ZN(n4519)
         );
  AOI21_X1 U5646 ( .B1(n6404), .B2(n4904), .A(n4519), .ZN(n4521) );
  NAND2_X1 U5647 ( .A1(n4828), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4520)
         );
  OAI211_X1 U5648 ( .C1(n4831), .C2(n4860), .A(n4521), .B(n4520), .ZN(U3119)
         );
  OAI22_X1 U5649 ( .A1(n6435), .A2(n4826), .B1(n4731), .B2(n4825), .ZN(n4522)
         );
  AOI21_X1 U5650 ( .B1(n6428), .B2(n4904), .A(n4522), .ZN(n4524) );
  NAND2_X1 U5651 ( .A1(n4828), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4523)
         );
  OAI211_X1 U5652 ( .C1(n4831), .C2(n4857), .A(n4524), .B(n4523), .ZN(U3123)
         );
  OAI22_X1 U5653 ( .A1(n6389), .A2(n4826), .B1(n4740), .B2(n4825), .ZN(n4525)
         );
  AOI21_X1 U5654 ( .B1(n6377), .B2(n4904), .A(n4525), .ZN(n4527) );
  NAND2_X1 U5655 ( .A1(n4828), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4526)
         );
  OAI211_X1 U5656 ( .C1(n4831), .C2(n4873), .A(n4527), .B(n4526), .ZN(U3116)
         );
  OAI22_X1 U5657 ( .A1(n6401), .A2(n4826), .B1(n4752), .B2(n4825), .ZN(n4528)
         );
  AOI21_X1 U5658 ( .B1(n6398), .B2(n4904), .A(n4528), .ZN(n4530) );
  NAND2_X1 U5659 ( .A1(n4828), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4529)
         );
  OAI211_X1 U5660 ( .C1(n4831), .C2(n4890), .A(n4530), .B(n4529), .ZN(U3118)
         );
  XNOR2_X1 U5661 ( .A(n4532), .B(n4531), .ZN(n4684) );
  NOR2_X1 U5662 ( .A1(n4691), .A2(n4533), .ZN(n4536) );
  OAI21_X1 U5663 ( .B1(n5720), .B2(n4536), .A(n6253), .ZN(n4692) );
  OAI21_X1 U5664 ( .B1(n4003), .B2(n3041), .A(n4766), .ZN(n6037) );
  NAND3_X1 U5665 ( .A1(n4536), .A2(n3997), .A3(n4535), .ZN(n4538) );
  INV_X1 U5666 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6521) );
  NOR2_X1 U5667 ( .A1(n6242), .A2(n6521), .ZN(n4680) );
  INV_X1 U5668 ( .A(n4680), .ZN(n4537) );
  OAI211_X1 U5669 ( .C1(n6229), .C2(n6037), .A(n4538), .B(n4537), .ZN(n4539)
         );
  AOI21_X1 U5670 ( .B1(n4692), .B2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n4539), 
        .ZN(n4540) );
  OAI21_X1 U5671 ( .B1(n4684), .B2(n6203), .A(n4540), .ZN(U3012) );
  NOR2_X1 U5672 ( .A1(n4549), .A2(n6295), .ZN(n6257) );
  NAND2_X1 U5673 ( .A1(n4543), .A2(n6343), .ZN(n6255) );
  AOI211_X1 U5674 ( .C1(n4592), .C2(n6297), .A(n6257), .B(n6255), .ZN(n4546)
         );
  NAND3_X1 U5675 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6458), .A3(n6445), .ZN(n6258) );
  NOR2_X1 U5676 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6258), .ZN(n4588)
         );
  NOR2_X1 U5677 ( .A1(n6569), .A2(n4588), .ZN(n4544) );
  NOR4_X2 U5678 ( .A1(n4546), .A2(n4639), .A3(n4545), .A4(n4544), .ZN(n4595)
         );
  INV_X1 U5679 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4553) );
  INV_X1 U5680 ( .A(n4860), .ZN(n6403) );
  INV_X1 U5681 ( .A(n6290), .ZN(n4548) );
  OAI22_X1 U5682 ( .A1(n6292), .A2(n4549), .B1(n4548), .B2(n4547), .ZN(n4589)
         );
  AOI22_X1 U5683 ( .A1(n6314), .A2(n4589), .B1(n6402), .B2(n4588), .ZN(n4550)
         );
  OAI21_X1 U5684 ( .B1(n6317), .B2(n6266), .A(n4550), .ZN(n4551) );
  AOI21_X1 U5685 ( .B1(n6403), .B2(n4592), .A(n4551), .ZN(n4552) );
  OAI21_X1 U5686 ( .B1(n4595), .B2(n4553), .A(n4552), .ZN(U3055) );
  INV_X1 U5687 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4557) );
  AOI22_X1 U5688 ( .A1(n6310), .A2(n4589), .B1(n6396), .B2(n4588), .ZN(n4554)
         );
  OAI21_X1 U5689 ( .B1(n6313), .B2(n6266), .A(n4554), .ZN(n4555) );
  AOI21_X1 U5690 ( .B1(n6397), .B2(n4592), .A(n4555), .ZN(n4556) );
  OAI21_X1 U5691 ( .B1(n4595), .B2(n4557), .A(n4556), .ZN(U3054) );
  INV_X1 U5692 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4561) );
  AOI22_X1 U5693 ( .A1(n6332), .A2(n4589), .B1(n6427), .B2(n4588), .ZN(n4558)
         );
  OAI21_X1 U5694 ( .B1(n6337), .B2(n6266), .A(n4558), .ZN(n4559) );
  AOI21_X1 U5695 ( .B1(n6431), .B2(n4592), .A(n4559), .ZN(n4560) );
  OAI21_X1 U5696 ( .B1(n4595), .B2(n4561), .A(n4560), .ZN(U3059) );
  INV_X1 U5697 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4565) );
  AOI22_X1 U5698 ( .A1(n6293), .A2(n4589), .B1(n6376), .B2(n4588), .ZN(n4562)
         );
  OAI21_X1 U5699 ( .B1(n6305), .B2(n6266), .A(n4562), .ZN(n4563) );
  AOI21_X1 U5700 ( .B1(n6386), .B2(n4592), .A(n4563), .ZN(n4564) );
  OAI21_X1 U5701 ( .B1(n4595), .B2(n4565), .A(n4564), .ZN(U3052) );
  INV_X1 U5702 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4569) );
  AOI22_X1 U5703 ( .A1(n6306), .A2(n4589), .B1(n6390), .B2(n4588), .ZN(n4566)
         );
  OAI21_X1 U5704 ( .B1(n6309), .B2(n6266), .A(n4566), .ZN(n4567) );
  AOI21_X1 U5705 ( .B1(n6392), .B2(n4592), .A(n4567), .ZN(n4568) );
  OAI21_X1 U5706 ( .B1(n4595), .B2(n4569), .A(n4568), .ZN(U3053) );
  INV_X1 U5707 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4574) );
  NAND2_X1 U5708 ( .A1(n6183), .A2(DATAI_30_), .ZN(n4876) );
  INV_X1 U5709 ( .A(n4876), .ZN(n6421) );
  INV_X1 U5710 ( .A(DATAI_22_), .ZN(n4570) );
  NOR2_X1 U5711 ( .A1(n6199), .A2(n4570), .ZN(n6422) );
  INV_X1 U5712 ( .A(n6422), .ZN(n6329) );
  NAND2_X1 U5713 ( .A1(DATAI_6_), .A2(n4582), .ZN(n6425) );
  INV_X1 U5714 ( .A(n6425), .ZN(n6326) );
  NOR2_X1 U5715 ( .A1(n4583), .A2(n3559), .ZN(n6420) );
  AOI22_X1 U5716 ( .A1(n6326), .A2(n4589), .B1(n6420), .B2(n4588), .ZN(n4571)
         );
  OAI21_X1 U5717 ( .B1(n6329), .B2(n6266), .A(n4571), .ZN(n4572) );
  AOI21_X1 U5718 ( .B1(n6421), .B2(n4592), .A(n4572), .ZN(n4573) );
  OAI21_X1 U5719 ( .B1(n4595), .B2(n4574), .A(n4573), .ZN(U3058) );
  INV_X1 U5720 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4580) );
  NAND2_X1 U5721 ( .A1(n6183), .A2(DATAI_28_), .ZN(n4854) );
  INV_X1 U5722 ( .A(n4854), .ZN(n6409) );
  INV_X1 U5723 ( .A(DATAI_20_), .ZN(n4575) );
  NOR2_X1 U5724 ( .A1(n6199), .A2(n4575), .ZN(n6410) );
  INV_X1 U5725 ( .A(n6410), .ZN(n6321) );
  NAND2_X1 U5726 ( .A1(DATAI_4_), .A2(n4582), .ZN(n6413) );
  INV_X1 U5727 ( .A(n6413), .ZN(n6318) );
  NOR2_X1 U5728 ( .A1(n4583), .A2(n4576), .ZN(n6408) );
  AOI22_X1 U5729 ( .A1(n6318), .A2(n4589), .B1(n6408), .B2(n4588), .ZN(n4577)
         );
  OAI21_X1 U5730 ( .B1(n6321), .B2(n6266), .A(n4577), .ZN(n4578) );
  AOI21_X1 U5731 ( .B1(n6409), .B2(n4592), .A(n4578), .ZN(n4579) );
  OAI21_X1 U5732 ( .B1(n4595), .B2(n4580), .A(n4579), .ZN(U3056) );
  INV_X1 U5733 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4587) );
  NAND2_X1 U5734 ( .A1(n6183), .A2(DATAI_21_), .ZN(n6325) );
  INV_X1 U5735 ( .A(n6325), .ZN(n6415) );
  INV_X1 U5736 ( .A(DATAI_29_), .ZN(n4581) );
  NOR2_X1 U5737 ( .A1(n6199), .A2(n4581), .ZN(n6416) );
  INV_X1 U5738 ( .A(n6416), .ZN(n4881) );
  NAND2_X1 U5739 ( .A1(DATAI_5_), .A2(n4582), .ZN(n6419) );
  INV_X1 U5740 ( .A(n6419), .ZN(n6322) );
  NOR2_X1 U5741 ( .A1(n4583), .A2(n3207), .ZN(n6414) );
  AOI22_X1 U5742 ( .A1(n6322), .A2(n4601), .B1(n6414), .B2(n4600), .ZN(n4584)
         );
  OAI21_X1 U5743 ( .B1(n4881), .B2(n4806), .A(n4584), .ZN(n4585) );
  AOI21_X1 U5744 ( .B1(n6415), .B2(n4704), .A(n4585), .ZN(n4586) );
  OAI21_X1 U5745 ( .B1(n4606), .B2(n4587), .A(n4586), .ZN(U3025) );
  INV_X1 U5746 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4594) );
  AOI22_X1 U5747 ( .A1(n6322), .A2(n4589), .B1(n6414), .B2(n4588), .ZN(n4590)
         );
  OAI21_X1 U5748 ( .B1(n6325), .B2(n6266), .A(n4590), .ZN(n4591) );
  AOI21_X1 U5749 ( .B1(n6416), .B2(n4592), .A(n4591), .ZN(n4593) );
  OAI21_X1 U5750 ( .B1(n4595), .B2(n4594), .A(n4593), .ZN(U3057) );
  INV_X1 U5751 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4599) );
  AOI22_X1 U5752 ( .A1(n6318), .A2(n4601), .B1(n6408), .B2(n4600), .ZN(n4596)
         );
  OAI21_X1 U5753 ( .B1(n4854), .B2(n4806), .A(n4596), .ZN(n4597) );
  AOI21_X1 U5754 ( .B1(n6410), .B2(n4704), .A(n4597), .ZN(n4598) );
  OAI21_X1 U5755 ( .B1(n4606), .B2(n4599), .A(n4598), .ZN(U3024) );
  INV_X1 U5756 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4605) );
  AOI22_X1 U5757 ( .A1(n6326), .A2(n4601), .B1(n6420), .B2(n4600), .ZN(n4602)
         );
  OAI21_X1 U5758 ( .B1(n4876), .B2(n4806), .A(n4602), .ZN(n4603) );
  AOI21_X1 U5759 ( .B1(n6422), .B2(n4704), .A(n4603), .ZN(n4604) );
  OAI21_X1 U5760 ( .B1(n4606), .B2(n4605), .A(n4604), .ZN(U3026) );
  AND2_X1 U5761 ( .A1(n4676), .A2(n4607), .ZN(n4610) );
  OR2_X1 U5762 ( .A1(n4610), .A2(n4609), .ZN(n6162) );
  AOI22_X1 U5763 ( .A1(n5557), .A2(DATAI_7_), .B1(n6608), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4611) );
  OAI21_X1 U5764 ( .B1(n6162), .B2(n5857), .A(n4611), .ZN(U2884) );
  NAND2_X1 U5765 ( .A1(n6371), .A2(n4614), .ZN(n4851) );
  INV_X1 U5766 ( .A(n4851), .ZN(n4612) );
  NAND3_X1 U5767 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6452), .A3(n6445), .ZN(n4848) );
  OR2_X1 U5768 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4848), .ZN(n4816)
         );
  AOI211_X1 U5769 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4816), .A(n6290), .B(
        n4613), .ZN(n4619) );
  INV_X1 U5770 ( .A(n4891), .ZN(n4615) );
  NOR3_X1 U5771 ( .A1(n4615), .A2(n3047), .A3(n6382), .ZN(n4617) );
  OAI22_X1 U5772 ( .A1(n4617), .A2(n4616), .B1(n5740), .B2(n4700), .ZN(n4618)
         );
  NAND2_X1 U5773 ( .A1(n4619), .A2(n4618), .ZN(n4815) );
  NAND2_X1 U5774 ( .A1(n4815), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4623) );
  INV_X1 U5775 ( .A(n4700), .ZN(n4845) );
  AOI22_X1 U5776 ( .A1(n4643), .A2(n4845), .B1(n4639), .B2(n4620), .ZN(n4818)
         );
  OAI22_X1 U5777 ( .A1(n6401), .A2(n4818), .B1(n4752), .B2(n4816), .ZN(n4621)
         );
  AOI21_X1 U5778 ( .B1(n6397), .B2(n3047), .A(n4621), .ZN(n4622) );
  OAI211_X1 U5779 ( .C1(n6313), .C2(n4891), .A(n4623), .B(n4622), .ZN(U3086)
         );
  NAND2_X1 U5780 ( .A1(n4815), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4626) );
  OAI22_X1 U5781 ( .A1(n6395), .A2(n4818), .B1(n4744), .B2(n4816), .ZN(n4624)
         );
  AOI21_X1 U5782 ( .B1(n6392), .B2(n3047), .A(n4624), .ZN(n4625) );
  OAI211_X1 U5783 ( .C1(n6309), .C2(n4891), .A(n4626), .B(n4625), .ZN(U3085)
         );
  NAND2_X1 U5784 ( .A1(n4815), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4629) );
  OAI22_X1 U5785 ( .A1(n6435), .A2(n4818), .B1(n4731), .B2(n4816), .ZN(n4627)
         );
  AOI21_X1 U5786 ( .B1(n6431), .B2(n3047), .A(n4627), .ZN(n4628) );
  OAI211_X1 U5787 ( .C1(n6337), .C2(n4891), .A(n4629), .B(n4628), .ZN(U3091)
         );
  NAND2_X1 U5788 ( .A1(n4815), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4632) );
  OAI22_X1 U5789 ( .A1(n6389), .A2(n4818), .B1(n4740), .B2(n4816), .ZN(n4630)
         );
  AOI21_X1 U5790 ( .B1(n6386), .B2(n3047), .A(n4630), .ZN(n4631) );
  OAI211_X1 U5791 ( .C1(n6305), .C2(n4891), .A(n4632), .B(n4631), .ZN(U3084)
         );
  NAND2_X1 U5792 ( .A1(n4815), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4635) );
  OAI22_X1 U5793 ( .A1(n6407), .A2(n4818), .B1(n4748), .B2(n4816), .ZN(n4633)
         );
  AOI21_X1 U5794 ( .B1(n6403), .B2(n3047), .A(n4633), .ZN(n4634) );
  OAI211_X1 U5795 ( .C1(n6317), .C2(n4891), .A(n4635), .B(n4634), .ZN(U3087)
         );
  INV_X1 U5796 ( .A(n4636), .ZN(n4724) );
  NAND2_X1 U5797 ( .A1(n4724), .A2(n6287), .ZN(n4908) );
  AOI21_X1 U5798 ( .B1(n4908), .B2(n4807), .A(n6487), .ZN(n4637) );
  NOR3_X1 U5799 ( .A1(n4637), .A2(n4644), .A3(n6382), .ZN(n4642) );
  NOR2_X1 U5800 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4638), .ZN(n4668)
         );
  NOR3_X1 U5801 ( .A1(n6301), .A2(n6458), .A3(n4639), .ZN(n4640) );
  OAI21_X1 U5802 ( .B1(n6569), .B2(n4668), .A(n4640), .ZN(n4641) );
  INV_X1 U5803 ( .A(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4649) );
  INV_X1 U5804 ( .A(n4643), .ZN(n4646) );
  INV_X1 U5805 ( .A(n4644), .ZN(n6296) );
  NAND3_X1 U5806 ( .A1(n6290), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6289), .ZN(n4645) );
  OAI21_X1 U5807 ( .B1(n4646), .B2(n6296), .A(n4645), .ZN(n4669) );
  AOI22_X1 U5808 ( .A1(n6310), .A2(n4669), .B1(n6396), .B2(n4668), .ZN(n4648)
         );
  INV_X1 U5809 ( .A(n4908), .ZN(n4671) );
  AOI22_X1 U5810 ( .A1(n4671), .A2(n6397), .B1(n4670), .B2(n6398), .ZN(n4647)
         );
  OAI211_X1 U5811 ( .C1(n4675), .C2(n4649), .A(n4648), .B(n4647), .ZN(U3134)
         );
  INV_X1 U5812 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4652) );
  AOI22_X1 U5813 ( .A1(n6306), .A2(n4669), .B1(n6390), .B2(n4668), .ZN(n4651)
         );
  AOI22_X1 U5814 ( .A1(n4671), .A2(n6392), .B1(n4670), .B2(n6391), .ZN(n4650)
         );
  OAI211_X1 U5815 ( .C1(n4675), .C2(n4652), .A(n4651), .B(n4650), .ZN(U3133)
         );
  INV_X1 U5816 ( .A(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4655) );
  AOI22_X1 U5817 ( .A1(n6293), .A2(n4669), .B1(n6376), .B2(n4668), .ZN(n4654)
         );
  AOI22_X1 U5818 ( .A1(n4671), .A2(n6386), .B1(n4670), .B2(n6377), .ZN(n4653)
         );
  OAI211_X1 U5819 ( .C1(n4675), .C2(n4655), .A(n4654), .B(n4653), .ZN(U3132)
         );
  INV_X1 U5820 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4658) );
  AOI22_X1 U5821 ( .A1(n6318), .A2(n4669), .B1(n6408), .B2(n4668), .ZN(n4657)
         );
  AOI22_X1 U5822 ( .A1(n4671), .A2(n6409), .B1(n4670), .B2(n6410), .ZN(n4656)
         );
  OAI211_X1 U5823 ( .C1(n4675), .C2(n4658), .A(n4657), .B(n4656), .ZN(U3136)
         );
  INV_X1 U5824 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4661) );
  AOI22_X1 U5825 ( .A1(n6332), .A2(n4669), .B1(n6427), .B2(n4668), .ZN(n4660)
         );
  AOI22_X1 U5826 ( .A1(n4671), .A2(n6431), .B1(n4670), .B2(n6428), .ZN(n4659)
         );
  OAI211_X1 U5827 ( .C1(n4675), .C2(n4661), .A(n4660), .B(n4659), .ZN(U3139)
         );
  INV_X1 U5828 ( .A(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4664) );
  AOI22_X1 U5829 ( .A1(n6326), .A2(n4669), .B1(n6420), .B2(n4668), .ZN(n4663)
         );
  AOI22_X1 U5830 ( .A1(n4671), .A2(n6421), .B1(n4670), .B2(n6422), .ZN(n4662)
         );
  OAI211_X1 U5831 ( .C1(n4675), .C2(n4664), .A(n4663), .B(n4662), .ZN(U3138)
         );
  INV_X1 U5832 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4667) );
  AOI22_X1 U5833 ( .A1(n6322), .A2(n4669), .B1(n6414), .B2(n4668), .ZN(n4666)
         );
  AOI22_X1 U5834 ( .A1(n4671), .A2(n6416), .B1(n4670), .B2(n6415), .ZN(n4665)
         );
  OAI211_X1 U5835 ( .C1(n4675), .C2(n4667), .A(n4666), .B(n4665), .ZN(U3137)
         );
  INV_X1 U5836 ( .A(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4674) );
  AOI22_X1 U5837 ( .A1(n6314), .A2(n4669), .B1(n6402), .B2(n4668), .ZN(n4673)
         );
  AOI22_X1 U5838 ( .A1(n4671), .A2(n6403), .B1(n4670), .B2(n6404), .ZN(n4672)
         );
  OAI211_X1 U5839 ( .C1(n4675), .C2(n4674), .A(n4673), .B(n4672), .ZN(U3135)
         );
  INV_X1 U5840 ( .A(n4676), .ZN(n4677) );
  AOI21_X1 U5841 ( .B1(n4679), .B2(n4678), .A(n4677), .ZN(n4685) );
  AOI21_X1 U5842 ( .B1(n6196), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n4680), 
        .ZN(n4681) );
  OAI21_X1 U5843 ( .B1(n6038), .B2(n6188), .A(n4681), .ZN(n4682) );
  AOI21_X1 U5844 ( .B1(n4685), .B2(n6183), .A(n4682), .ZN(n4683) );
  OAI21_X1 U5845 ( .B1(n4684), .B2(n6190), .A(n4683), .ZN(U2980) );
  INV_X1 U5846 ( .A(n4685), .ZN(n6040) );
  INV_X1 U5847 ( .A(n6037), .ZN(n4686) );
  AOI22_X1 U5848 ( .A1(n4686), .A2(n6081), .B1(n5505), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n4687) );
  OAI21_X1 U5849 ( .B1(n6040), .B2(n6085), .A(n4687), .ZN(U2853) );
  XOR2_X1 U5850 ( .A(n4688), .B(n4689), .Z(n6171) );
  NOR4_X1 U5851 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4690), .A3(n6237), 
        .A4(n6245), .ZN(n4696) );
  NOR3_X1 U5852 ( .A1(n4691), .A2(n6236), .A3(n4690), .ZN(n4693) );
  OAI21_X1 U5853 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n4693), .A(n4692), 
        .ZN(n4694) );
  NAND2_X1 U5854 ( .A1(n6218), .A2(REIP_REG_5__SCAN_IN), .ZN(n6172) );
  OAI211_X1 U5855 ( .C1(n6229), .C2(n6047), .A(n4694), .B(n6172), .ZN(n4695)
         );
  AOI211_X1 U5856 ( .C1(n6171), .C2(n6247), .A(n4696), .B(n4695), .ZN(n4697)
         );
  INV_X1 U5857 ( .A(n4697), .ZN(U3013) );
  INV_X1 U5858 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6122) );
  OAI222_X1 U5859 ( .A1(n6040), .A2(n5857), .B1(n5010), .B2(n4698), .C1(n6122), 
        .C2(n5293), .ZN(U2885) );
  OAI21_X1 U5860 ( .B1(n4699), .B2(n6487), .A(n6343), .ZN(n4709) );
  INV_X1 U5861 ( .A(n4709), .ZN(n4703) );
  OR3_X1 U5862 ( .A1(n4700), .A2(n5747), .A3(n6373), .ZN(n4701) );
  OR2_X1 U5863 ( .A1(n6256), .A2(n4706), .ZN(n4780) );
  NAND2_X1 U5864 ( .A1(n4701), .A2(n4780), .ZN(n4708) );
  INV_X1 U5865 ( .A(n4706), .ZN(n4702) );
  AOI22_X1 U5866 ( .A1(n4703), .A2(n4708), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4702), .ZN(n4786) );
  INV_X1 U5867 ( .A(n4704), .ZN(n4779) );
  OAI22_X1 U5868 ( .A1(n4744), .A2(n4780), .B1(n4779), .B2(n4884), .ZN(n4705)
         );
  AOI21_X1 U5869 ( .B1(n6391), .B2(n4782), .A(n4705), .ZN(n4711) );
  AOI21_X1 U5870 ( .B1(n6382), .B2(n4706), .A(n6380), .ZN(n4707) );
  OAI21_X1 U5871 ( .B1(n4709), .B2(n4708), .A(n4707), .ZN(n4783) );
  NAND2_X1 U5872 ( .A1(n4783), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4710) );
  OAI211_X1 U5873 ( .C1(n4786), .C2(n6395), .A(n4711), .B(n4710), .ZN(U3029)
         );
  OAI22_X1 U5874 ( .A1(n4740), .A2(n4780), .B1(n4779), .B2(n4873), .ZN(n4712)
         );
  AOI21_X1 U5875 ( .B1(n6377), .B2(n4782), .A(n4712), .ZN(n4714) );
  NAND2_X1 U5876 ( .A1(n4783), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4713) );
  OAI211_X1 U5877 ( .C1(n4786), .C2(n6389), .A(n4714), .B(n4713), .ZN(U3028)
         );
  OAI22_X1 U5878 ( .A1(n4748), .A2(n4780), .B1(n4779), .B2(n4860), .ZN(n4715)
         );
  AOI21_X1 U5879 ( .B1(n6404), .B2(n4782), .A(n4715), .ZN(n4717) );
  NAND2_X1 U5880 ( .A1(n4783), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4716) );
  OAI211_X1 U5881 ( .C1(n4786), .C2(n6407), .A(n4717), .B(n4716), .ZN(U3031)
         );
  OAI22_X1 U5882 ( .A1(n4731), .A2(n4780), .B1(n4779), .B2(n4857), .ZN(n4718)
         );
  AOI21_X1 U5883 ( .B1(n6428), .B2(n4782), .A(n4718), .ZN(n4720) );
  NAND2_X1 U5884 ( .A1(n4783), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4719) );
  OAI211_X1 U5885 ( .C1(n4786), .C2(n6435), .A(n4720), .B(n4719), .ZN(U3035)
         );
  OAI22_X1 U5886 ( .A1(n4752), .A2(n4780), .B1(n4779), .B2(n4890), .ZN(n4721)
         );
  AOI21_X1 U5887 ( .B1(n6398), .B2(n4782), .A(n4721), .ZN(n4723) );
  NAND2_X1 U5888 ( .A1(n4783), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4722) );
  OAI211_X1 U5889 ( .C1(n4786), .C2(n6401), .A(n4723), .B(n4722), .ZN(U3030)
         );
  INV_X1 U5890 ( .A(n6371), .ZN(n4725) );
  NAND2_X1 U5891 ( .A1(n4724), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4861) );
  NAND2_X1 U5892 ( .A1(n4725), .A2(n4861), .ZN(n5738) );
  NAND2_X1 U5893 ( .A1(n5744), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6369) );
  NOR3_X1 U5894 ( .A1(n5738), .A2(n3376), .A3(n6369), .ZN(n4726) );
  NOR2_X1 U5895 ( .A1(n4726), .A2(n6382), .ZN(n4733) );
  OR2_X1 U5896 ( .A1(n4727), .A2(n6373), .ZN(n4729) );
  INV_X1 U5897 ( .A(n4728), .ZN(n6372) );
  NAND2_X1 U5898 ( .A1(n6372), .A2(n6458), .ZN(n4770) );
  NAND2_X1 U5899 ( .A1(n4729), .A2(n4770), .ZN(n4736) );
  INV_X1 U5900 ( .A(n4734), .ZN(n4730) );
  AOI22_X1 U5901 ( .A1(n4733), .A2(n4736), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4730), .ZN(n4775) );
  OAI22_X1 U5902 ( .A1(n4731), .A2(n4770), .B1(n6337), .B2(n4769), .ZN(n4732)
         );
  AOI21_X1 U5903 ( .B1(n6431), .B2(n4841), .A(n4732), .ZN(n4739) );
  INV_X1 U5904 ( .A(n4733), .ZN(n4737) );
  AOI21_X1 U5905 ( .B1(n6382), .B2(n4734), .A(n6380), .ZN(n4735) );
  OAI21_X1 U5906 ( .B1(n4737), .B2(n4736), .A(n4735), .ZN(n4772) );
  NAND2_X1 U5907 ( .A1(n4772), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4738) );
  OAI211_X1 U5908 ( .C1(n4775), .C2(n6435), .A(n4739), .B(n4738), .ZN(U3051)
         );
  OAI22_X1 U5909 ( .A1(n4740), .A2(n4770), .B1(n6305), .B2(n4769), .ZN(n4741)
         );
  AOI21_X1 U5910 ( .B1(n6386), .B2(n4841), .A(n4741), .ZN(n4743) );
  NAND2_X1 U5911 ( .A1(n4772), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4742) );
  OAI211_X1 U5912 ( .C1(n4775), .C2(n6389), .A(n4743), .B(n4742), .ZN(U3044)
         );
  OAI22_X1 U5913 ( .A1(n4744), .A2(n4770), .B1(n6309), .B2(n4769), .ZN(n4745)
         );
  AOI21_X1 U5914 ( .B1(n6392), .B2(n4841), .A(n4745), .ZN(n4747) );
  NAND2_X1 U5915 ( .A1(n4772), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4746) );
  OAI211_X1 U5916 ( .C1(n4775), .C2(n6395), .A(n4747), .B(n4746), .ZN(U3045)
         );
  OAI22_X1 U5917 ( .A1(n4748), .A2(n4770), .B1(n6317), .B2(n4769), .ZN(n4749)
         );
  AOI21_X1 U5918 ( .B1(n6403), .B2(n4841), .A(n4749), .ZN(n4751) );
  NAND2_X1 U5919 ( .A1(n4772), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4750) );
  OAI211_X1 U5920 ( .C1(n4775), .C2(n6407), .A(n4751), .B(n4750), .ZN(U3047)
         );
  OAI22_X1 U5921 ( .A1(n4752), .A2(n4770), .B1(n6313), .B2(n4769), .ZN(n4753)
         );
  AOI21_X1 U5922 ( .B1(n6397), .B2(n4841), .A(n4753), .ZN(n4755) );
  NAND2_X1 U5923 ( .A1(n4772), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4754) );
  OAI211_X1 U5924 ( .C1(n4775), .C2(n6401), .A(n4755), .B(n4754), .ZN(U3046)
         );
  INV_X1 U5925 ( .A(n6420), .ZN(n4832) );
  OAI22_X1 U5926 ( .A1(n4832), .A2(n4770), .B1(n6329), .B2(n4769), .ZN(n4756)
         );
  AOI21_X1 U5927 ( .B1(n6421), .B2(n4841), .A(n4756), .ZN(n4758) );
  NAND2_X1 U5928 ( .A1(n4772), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4757) );
  OAI211_X1 U5929 ( .C1(n4775), .C2(n6425), .A(n4758), .B(n4757), .ZN(U3050)
         );
  INV_X1 U5930 ( .A(n6408), .ZN(n4838) );
  OAI22_X1 U5931 ( .A1(n4838), .A2(n4770), .B1(n6321), .B2(n4769), .ZN(n4759)
         );
  AOI21_X1 U5932 ( .B1(n6409), .B2(n4841), .A(n4759), .ZN(n4761) );
  NAND2_X1 U5933 ( .A1(n4772), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4760) );
  OAI211_X1 U5934 ( .C1(n4775), .C2(n6413), .A(n4761), .B(n4760), .ZN(U3048)
         );
  INV_X1 U5935 ( .A(n6414), .ZN(n4817) );
  OAI22_X1 U5936 ( .A1(n4817), .A2(n4780), .B1(n4779), .B2(n4881), .ZN(n4762)
         );
  AOI21_X1 U5937 ( .B1(n6415), .B2(n4782), .A(n4762), .ZN(n4764) );
  NAND2_X1 U5938 ( .A1(n4783), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4763) );
  OAI211_X1 U5939 ( .C1(n4786), .C2(n6419), .A(n4764), .B(n4763), .ZN(U3033)
         );
  AND2_X1 U5940 ( .A1(n4766), .A2(n4765), .ZN(n4767) );
  OR2_X1 U5941 ( .A1(n4767), .A2(n4913), .ZN(n6019) );
  INV_X1 U5942 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4768) );
  OAI222_X1 U5943 ( .A1(n6019), .A2(n6090), .B1(n4768), .B2(n6094), .C1(n6162), 
        .C2(n6085), .ZN(U2852) );
  OAI22_X1 U5944 ( .A1(n4817), .A2(n4770), .B1(n6325), .B2(n4769), .ZN(n4771)
         );
  AOI21_X1 U5945 ( .B1(n6416), .B2(n4841), .A(n4771), .ZN(n4774) );
  NAND2_X1 U5946 ( .A1(n4772), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4773) );
  OAI211_X1 U5947 ( .C1(n4775), .C2(n6419), .A(n4774), .B(n4773), .ZN(U3049)
         );
  OAI22_X1 U5948 ( .A1(n4838), .A2(n4780), .B1(n4779), .B2(n4854), .ZN(n4776)
         );
  AOI21_X1 U5949 ( .B1(n6410), .B2(n4782), .A(n4776), .ZN(n4778) );
  NAND2_X1 U5950 ( .A1(n4783), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4777) );
  OAI211_X1 U5951 ( .C1(n4786), .C2(n6413), .A(n4778), .B(n4777), .ZN(U3032)
         );
  OAI22_X1 U5952 ( .A1(n4832), .A2(n4780), .B1(n4779), .B2(n4876), .ZN(n4781)
         );
  AOI21_X1 U5953 ( .B1(n6422), .B2(n4782), .A(n4781), .ZN(n4785) );
  NAND2_X1 U5954 ( .A1(n4783), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4784) );
  OAI211_X1 U5955 ( .C1(n4786), .C2(n6425), .A(n4785), .B(n4784), .ZN(U3034)
         );
  NOR2_X1 U5956 ( .A1(n4609), .A2(n4787), .ZN(n4788) );
  OR2_X1 U5957 ( .A1(n4922), .A2(n4788), .ZN(n5475) );
  INV_X1 U5958 ( .A(DATAI_8_), .ZN(n6781) );
  INV_X1 U5959 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6117) );
  OAI222_X1 U5960 ( .A1(n5475), .A2(n5857), .B1(n5010), .B2(n6781), .C1(n5293), 
        .C2(n6117), .ZN(U2883) );
  NAND2_X1 U5961 ( .A1(n4815), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4791) );
  OAI22_X1 U5962 ( .A1(n6413), .A2(n4818), .B1(n4838), .B2(n4816), .ZN(n4789)
         );
  AOI21_X1 U5963 ( .B1(n6409), .B2(n3047), .A(n4789), .ZN(n4790) );
  OAI211_X1 U5964 ( .C1(n6321), .C2(n4891), .A(n4791), .B(n4790), .ZN(U3088)
         );
  NAND2_X1 U5965 ( .A1(n4815), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4794) );
  OAI22_X1 U5966 ( .A1(n6425), .A2(n4818), .B1(n4832), .B2(n4816), .ZN(n4792)
         );
  AOI21_X1 U5967 ( .B1(n6421), .B2(n3047), .A(n4792), .ZN(n4793) );
  OAI211_X1 U5968 ( .C1(n6329), .C2(n4891), .A(n4794), .B(n4793), .ZN(U3090)
         );
  OAI22_X1 U5969 ( .A1(n6419), .A2(n4826), .B1(n4817), .B2(n4825), .ZN(n4795)
         );
  AOI21_X1 U5970 ( .B1(n6415), .B2(n4904), .A(n4795), .ZN(n4797) );
  NAND2_X1 U5971 ( .A1(n4828), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4796)
         );
  OAI211_X1 U5972 ( .C1(n4831), .C2(n4881), .A(n4797), .B(n4796), .ZN(U3121)
         );
  OAI22_X1 U5973 ( .A1(n6413), .A2(n4805), .B1(n4804), .B2(n4838), .ZN(n4799)
         );
  OAI22_X1 U5974 ( .A1(n4854), .A2(n4807), .B1(n4806), .B2(n6321), .ZN(n4798)
         );
  AOI211_X1 U5975 ( .C1(n4810), .C2(INSTQUEUE_REG_15__4__SCAN_IN), .A(n4799), 
        .B(n4798), .ZN(n4800) );
  INV_X1 U5976 ( .A(n4800), .ZN(U3144) );
  OAI22_X1 U5977 ( .A1(n6425), .A2(n4805), .B1(n4804), .B2(n4832), .ZN(n4802)
         );
  OAI22_X1 U5978 ( .A1(n4876), .A2(n4807), .B1(n4806), .B2(n6329), .ZN(n4801)
         );
  AOI211_X1 U5979 ( .C1(n4810), .C2(INSTQUEUE_REG_15__6__SCAN_IN), .A(n4802), 
        .B(n4801), .ZN(n4803) );
  INV_X1 U5980 ( .A(n4803), .ZN(U3146) );
  OAI22_X1 U5981 ( .A1(n6419), .A2(n4805), .B1(n4804), .B2(n4817), .ZN(n4809)
         );
  OAI22_X1 U5982 ( .A1(n4881), .A2(n4807), .B1(n4806), .B2(n6325), .ZN(n4808)
         );
  AOI211_X1 U5983 ( .C1(n4810), .C2(INSTQUEUE_REG_15__5__SCAN_IN), .A(n4809), 
        .B(n4808), .ZN(n4811) );
  INV_X1 U5984 ( .A(n4811), .ZN(U3145) );
  NAND2_X1 U5985 ( .A1(n4836), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4814) );
  OAI22_X1 U5986 ( .A1(n6419), .A2(n4839), .B1(n4817), .B2(n4837), .ZN(n4812)
         );
  AOI21_X1 U5987 ( .B1(n6415), .B2(n4841), .A(n4812), .ZN(n4813) );
  OAI211_X1 U5988 ( .C1(n4844), .C2(n4881), .A(n4814), .B(n4813), .ZN(U3041)
         );
  NAND2_X1 U5989 ( .A1(n4815), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4821) );
  OAI22_X1 U5990 ( .A1(n6419), .A2(n4818), .B1(n4817), .B2(n4816), .ZN(n4819)
         );
  AOI21_X1 U5991 ( .B1(n6416), .B2(n3047), .A(n4819), .ZN(n4820) );
  OAI211_X1 U5992 ( .C1(n6325), .C2(n4891), .A(n4821), .B(n4820), .ZN(U3089)
         );
  OAI22_X1 U5993 ( .A1(n6413), .A2(n4826), .B1(n4838), .B2(n4825), .ZN(n4822)
         );
  AOI21_X1 U5994 ( .B1(n6410), .B2(n4904), .A(n4822), .ZN(n4824) );
  NAND2_X1 U5995 ( .A1(n4828), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4823)
         );
  OAI211_X1 U5996 ( .C1(n4831), .C2(n4854), .A(n4824), .B(n4823), .ZN(U3120)
         );
  OAI22_X1 U5997 ( .A1(n6425), .A2(n4826), .B1(n4832), .B2(n4825), .ZN(n4827)
         );
  AOI21_X1 U5998 ( .B1(n6422), .B2(n4904), .A(n4827), .ZN(n4830) );
  NAND2_X1 U5999 ( .A1(n4828), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4829)
         );
  OAI211_X1 U6000 ( .C1(n4831), .C2(n4876), .A(n4830), .B(n4829), .ZN(U3122)
         );
  NAND2_X1 U6001 ( .A1(n4836), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4835) );
  OAI22_X1 U6002 ( .A1(n6425), .A2(n4839), .B1(n4832), .B2(n4837), .ZN(n4833)
         );
  AOI21_X1 U6003 ( .B1(n6422), .B2(n4841), .A(n4833), .ZN(n4834) );
  OAI211_X1 U6004 ( .C1(n4844), .C2(n4876), .A(n4835), .B(n4834), .ZN(U3042)
         );
  NAND2_X1 U6005 ( .A1(n4836), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4843) );
  OAI22_X1 U6006 ( .A1(n6413), .A2(n4839), .B1(n4838), .B2(n4837), .ZN(n4840)
         );
  AOI21_X1 U6007 ( .B1(n6410), .B2(n4841), .A(n4840), .ZN(n4842) );
  OAI211_X1 U6008 ( .C1(n4844), .C2(n4854), .A(n4843), .B(n4842), .ZN(U3040)
         );
  OAI21_X1 U6009 ( .B1(n4851), .B2(n6487), .A(n6343), .ZN(n4850) );
  NOR2_X1 U6010 ( .A1(n6256), .A2(n4848), .ZN(n4887) );
  AOI21_X1 U6011 ( .B1(n4863), .B2(n4845), .A(n4887), .ZN(n4849) );
  INV_X1 U6012 ( .A(n4849), .ZN(n4847) );
  AOI21_X1 U6013 ( .B1(n6382), .B2(n4848), .A(n6380), .ZN(n4846) );
  OAI21_X1 U6014 ( .B1(n4850), .B2(n4847), .A(n4846), .ZN(n4886) );
  OAI22_X1 U6015 ( .A1(n4850), .A2(n4849), .B1(n6486), .B2(n4848), .ZN(n4885)
         );
  AOI22_X1 U6016 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4886), .B1(n6318), 
        .B2(n4885), .ZN(n4853) );
  NOR2_X2 U6017 ( .A1(n4851), .A2(n3032), .ZN(n5782) );
  AOI22_X1 U6018 ( .A1(n5782), .A2(n6410), .B1(n4887), .B2(n6408), .ZN(n4852)
         );
  OAI211_X1 U6019 ( .C1(n4891), .C2(n4854), .A(n4853), .B(n4852), .ZN(U3096)
         );
  AOI22_X1 U6020 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4886), .B1(n6332), 
        .B2(n4885), .ZN(n4856) );
  AOI22_X1 U6021 ( .A1(n5782), .A2(n6428), .B1(n4887), .B2(n6427), .ZN(n4855)
         );
  OAI211_X1 U6022 ( .C1(n4891), .C2(n4857), .A(n4856), .B(n4855), .ZN(U3099)
         );
  AOI22_X1 U6023 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4886), .B1(n6314), 
        .B2(n4885), .ZN(n4859) );
  AOI22_X1 U6024 ( .A1(n5782), .A2(n6404), .B1(n4887), .B2(n6402), .ZN(n4858)
         );
  OAI211_X1 U6025 ( .C1(n4891), .C2(n4860), .A(n4859), .B(n4858), .ZN(U3095)
         );
  NAND2_X1 U6026 ( .A1(n6343), .A2(n4861), .ZN(n4867) );
  NOR2_X1 U6027 ( .A1(n6256), .A2(n4866), .ZN(n4905) );
  AOI21_X1 U6028 ( .B1(n4863), .B2(n4862), .A(n4905), .ZN(n4868) );
  INV_X1 U6029 ( .A(n4868), .ZN(n4865) );
  AOI21_X1 U6030 ( .B1(n6382), .B2(n4866), .A(n6380), .ZN(n4864) );
  OAI21_X1 U6031 ( .B1(n4867), .B2(n4865), .A(n4864), .ZN(n4903) );
  OAI22_X1 U6032 ( .A1(n4868), .A2(n4867), .B1(n6486), .B2(n4866), .ZN(n4902)
         );
  AOI22_X1 U6033 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4903), .B1(n6293), 
        .B2(n4902), .ZN(n4870) );
  AOI22_X1 U6034 ( .A1(n6376), .A2(n4905), .B1(n6386), .B2(n4904), .ZN(n4869)
         );
  OAI211_X1 U6035 ( .C1(n6305), .C2(n4908), .A(n4870), .B(n4869), .ZN(U3124)
         );
  AOI22_X1 U6036 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4886), .B1(n6293), 
        .B2(n4885), .ZN(n4872) );
  AOI22_X1 U6037 ( .A1(n5782), .A2(n6377), .B1(n6376), .B2(n4887), .ZN(n4871)
         );
  OAI211_X1 U6038 ( .C1(n4891), .C2(n4873), .A(n4872), .B(n4871), .ZN(U3092)
         );
  AOI22_X1 U6039 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4886), .B1(n6326), 
        .B2(n4885), .ZN(n4875) );
  AOI22_X1 U6040 ( .A1(n5782), .A2(n6422), .B1(n4887), .B2(n6420), .ZN(n4874)
         );
  OAI211_X1 U6041 ( .C1(n4891), .C2(n4876), .A(n4875), .B(n4874), .ZN(U3098)
         );
  AOI22_X1 U6042 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4903), .B1(n6332), 
        .B2(n4902), .ZN(n4878) );
  AOI22_X1 U6043 ( .A1(n6427), .A2(n4905), .B1(n6431), .B2(n4904), .ZN(n4877)
         );
  OAI211_X1 U6044 ( .C1(n6337), .C2(n4908), .A(n4878), .B(n4877), .ZN(U3131)
         );
  AOI22_X1 U6045 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4886), .B1(n6322), 
        .B2(n4885), .ZN(n4880) );
  AOI22_X1 U6046 ( .A1(n5782), .A2(n6415), .B1(n4887), .B2(n6414), .ZN(n4879)
         );
  OAI211_X1 U6047 ( .C1(n4891), .C2(n4881), .A(n4880), .B(n4879), .ZN(U3097)
         );
  AOI22_X1 U6048 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4886), .B1(n6306), 
        .B2(n4885), .ZN(n4883) );
  AOI22_X1 U6049 ( .A1(n5782), .A2(n6391), .B1(n4887), .B2(n6390), .ZN(n4882)
         );
  OAI211_X1 U6050 ( .C1(n4891), .C2(n4884), .A(n4883), .B(n4882), .ZN(U3093)
         );
  AOI22_X1 U6051 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4886), .B1(n6310), 
        .B2(n4885), .ZN(n4889) );
  AOI22_X1 U6052 ( .A1(n5782), .A2(n6398), .B1(n4887), .B2(n6396), .ZN(n4888)
         );
  OAI211_X1 U6053 ( .C1(n4891), .C2(n4890), .A(n4889), .B(n4888), .ZN(U3094)
         );
  AOI22_X1 U6054 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4903), .B1(n6326), 
        .B2(n4902), .ZN(n4893) );
  AOI22_X1 U6055 ( .A1(n6420), .A2(n4905), .B1(n6421), .B2(n4904), .ZN(n4892)
         );
  OAI211_X1 U6056 ( .C1(n6329), .C2(n4908), .A(n4893), .B(n4892), .ZN(U3130)
         );
  AOI22_X1 U6057 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4903), .B1(n6322), 
        .B2(n4902), .ZN(n4895) );
  AOI22_X1 U6058 ( .A1(n6414), .A2(n4905), .B1(n6416), .B2(n4904), .ZN(n4894)
         );
  OAI211_X1 U6059 ( .C1(n6325), .C2(n4908), .A(n4895), .B(n4894), .ZN(U3129)
         );
  AOI22_X1 U6060 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4903), .B1(n6310), 
        .B2(n4902), .ZN(n4897) );
  AOI22_X1 U6061 ( .A1(n6396), .A2(n4905), .B1(n6397), .B2(n4904), .ZN(n4896)
         );
  OAI211_X1 U6062 ( .C1(n6313), .C2(n4908), .A(n4897), .B(n4896), .ZN(U3126)
         );
  AOI22_X1 U6063 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4903), .B1(n6314), 
        .B2(n4902), .ZN(n4899) );
  AOI22_X1 U6064 ( .A1(n6402), .A2(n4905), .B1(n6403), .B2(n4904), .ZN(n4898)
         );
  OAI211_X1 U6065 ( .C1(n6317), .C2(n4908), .A(n4899), .B(n4898), .ZN(U3127)
         );
  AOI22_X1 U6066 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4903), .B1(n6318), 
        .B2(n4902), .ZN(n4901) );
  AOI22_X1 U6067 ( .A1(n6408), .A2(n4905), .B1(n6409), .B2(n4904), .ZN(n4900)
         );
  OAI211_X1 U6068 ( .C1(n6321), .C2(n4908), .A(n4901), .B(n4900), .ZN(U3128)
         );
  AOI22_X1 U6069 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4903), .B1(n6306), 
        .B2(n4902), .ZN(n4907) );
  AOI22_X1 U6070 ( .A1(n6390), .A2(n4905), .B1(n6392), .B2(n4904), .ZN(n4906)
         );
  OAI211_X1 U6071 ( .C1(n6309), .C2(n4908), .A(n4907), .B(n4906), .ZN(U3125)
         );
  XNOR2_X1 U6072 ( .A(n4909), .B(n4910), .ZN(n4932) );
  NOR2_X1 U6073 ( .A1(n4911), .A2(n5053), .ZN(n6215) );
  OAI211_X1 U6074 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n6215), .B(n6212), .ZN(n4917) );
  NOR2_X1 U6075 ( .A1(n4913), .A2(n4912), .ZN(n4914) );
  OR2_X1 U6076 ( .A1(n4926), .A2(n4914), .ZN(n5466) );
  INV_X1 U6077 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6524) );
  OAI22_X1 U6078 ( .A1(n6229), .A2(n5466), .B1(n6524), .B2(n6242), .ZN(n4915)
         );
  AOI21_X1 U6079 ( .B1(n6211), .B2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n4915), 
        .ZN(n4916) );
  OAI211_X1 U6080 ( .C1(n4932), .C2(n6203), .A(n4917), .B(n4916), .ZN(U3010)
         );
  INV_X1 U6081 ( .A(n5475), .ZN(n4930) );
  INV_X1 U6082 ( .A(n5533), .ZN(n6092) );
  OAI22_X1 U6083 ( .A1(n5466), .A2(n6090), .B1(n5470), .B2(n6094), .ZN(n4918)
         );
  AOI21_X1 U6084 ( .B1(n4930), .B2(n6092), .A(n4918), .ZN(n4919) );
  INV_X1 U6085 ( .A(n4919), .ZN(U2851) );
  OR2_X1 U6086 ( .A1(n4922), .A2(n4921), .ZN(n4923) );
  NAND2_X1 U6087 ( .A1(n4941), .A2(n4923), .ZN(n6010) );
  INV_X1 U6088 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6789) );
  OAI222_X1 U6089 ( .A1(n6010), .A2(n5857), .B1(n5010), .B2(n4924), .C1(n5293), 
        .C2(n6789), .ZN(U2882) );
  OAI21_X1 U6090 ( .B1(n4926), .B2(n4925), .A(n4988), .ZN(n6228) );
  INV_X1 U6091 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4927) );
  OAI222_X1 U6092 ( .A1(n6228), .A2(n6090), .B1(n4927), .B2(n6094), .C1(n6010), 
        .C2(n6085), .ZN(U2850) );
  AOI22_X1 U6093 ( .A1(n6196), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n6218), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n4928) );
  OAI21_X1 U6094 ( .B1(n5467), .B2(n6188), .A(n4928), .ZN(n4929) );
  AOI21_X1 U6095 ( .B1(n4930), .B2(n6183), .A(n4929), .ZN(n4931) );
  OAI21_X1 U6096 ( .B1(n4932), .B2(n6190), .A(n4931), .ZN(U2978) );
  INV_X1 U6097 ( .A(n6215), .ZN(n4938) );
  XOR2_X1 U6098 ( .A(n4934), .B(n4933), .Z(n6164) );
  NAND2_X1 U6099 ( .A1(n6164), .A2(n6247), .ZN(n4937) );
  NAND2_X1 U6100 ( .A1(n6218), .A2(REIP_REG_7__SCAN_IN), .ZN(n6165) );
  OAI21_X1 U6101 ( .B1(n6229), .B2(n6019), .A(n6165), .ZN(n4935) );
  AOI21_X1 U6102 ( .B1(n6211), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n4935), 
        .ZN(n4936) );
  OAI211_X1 U6103 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n4938), .A(n4937), 
        .B(n4936), .ZN(U3011) );
  INV_X1 U6104 ( .A(n4992), .ZN(n4940) );
  AOI21_X1 U6105 ( .B1(n4942), .B2(n4941), .A(n4940), .ZN(n4985) );
  INV_X1 U6106 ( .A(n4985), .ZN(n5465) );
  AOI22_X1 U6107 ( .A1(n5557), .A2(DATAI_10_), .B1(n6608), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4943) );
  OAI21_X1 U6108 ( .B1(n5465), .B2(n5857), .A(n4943), .ZN(U2881) );
  NOR3_X1 U6109 ( .A1(n6780), .A2(n6569), .A3(n6493), .ZN(n6478) );
  AND2_X1 U6110 ( .A1(n4944), .A2(n5205), .ZN(n4945) );
  OR2_X1 U6111 ( .A1(n6218), .A2(n4945), .ZN(n4946) );
  OR2_X1 U6112 ( .A1(n6478), .A2(n4946), .ZN(n4947) );
  NAND2_X1 U6113 ( .A1(n4971), .A2(n4948), .ZN(n4951) );
  INV_X1 U6114 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5590) );
  INV_X1 U6115 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5580) );
  INV_X1 U6116 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U6117 ( .A1(n5200), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5202)
         );
  INV_X1 U6118 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5323) );
  INV_X1 U6119 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5303) );
  XNOR2_X1 U6120 ( .A(n4949), .B(n5303), .ZN(n5282) );
  NOR2_X1 U6121 ( .A1(n5282), .A2(n6765), .ZN(n4950) );
  NAND2_X1 U6122 ( .A1(n4951), .A2(n6039), .ZN(n6054) );
  NAND2_X1 U6123 ( .A1(n4971), .A2(n4952), .ZN(n6059) );
  INV_X1 U6124 ( .A(n6026), .ZN(n4953) );
  AOI22_X1 U6125 ( .A1(n6034), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n4953), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4956) );
  AND2_X1 U6126 ( .A1(n5282), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4954) );
  NAND2_X1 U6127 ( .A1(n6053), .A2(n4282), .ZN(n4955) );
  OAI211_X1 U6128 ( .C1(n6059), .C2(n5731), .A(n4956), .B(n4955), .ZN(n4975)
         );
  NOR2_X1 U6129 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4966) );
  INV_X1 U6130 ( .A(n4966), .ZN(n4957) );
  OR2_X1 U6131 ( .A1(n6503), .A2(n4957), .ZN(n6473) );
  NAND2_X1 U6132 ( .A1(n4958), .A2(n6473), .ZN(n5301) );
  NOR2_X1 U6133 ( .A1(n4966), .A2(EBX_REG_31__SCAN_IN), .ZN(n4959) );
  NAND2_X1 U6134 ( .A1(n4965), .A2(n4959), .ZN(n4960) );
  NAND2_X1 U6135 ( .A1(n5301), .A2(n4960), .ZN(n4961) );
  NAND2_X1 U6136 ( .A1(n4971), .A2(EBX_REG_31__SCAN_IN), .ZN(n5302) );
  INV_X1 U6137 ( .A(n5302), .ZN(n4964) );
  NOR2_X1 U6138 ( .A1(n4962), .A2(n4966), .ZN(n4963) );
  NAND2_X1 U6139 ( .A1(n6064), .A2(n4301), .ZN(n4972) );
  OAI211_X1 U6140 ( .C1(n4968), .C2(n4967), .A(n4966), .B(n4965), .ZN(n4969)
         );
  INV_X1 U6141 ( .A(n4969), .ZN(n4970) );
  INV_X1 U6142 ( .A(n6046), .ZN(n5460) );
  INV_X1 U6143 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U6144 ( .A1(n5460), .A2(n5490), .ZN(n5483) );
  OAI211_X1 U6145 ( .C1(n4973), .C2(n6078), .A(n4972), .B(n5483), .ZN(n4974)
         );
  AOI211_X1 U6146 ( .C1(n4976), .C2(n6054), .A(n4975), .B(n4974), .ZN(n4977)
         );
  INV_X1 U6147 ( .A(n4977), .ZN(U2826) );
  INV_X1 U6148 ( .A(n4979), .ZN(n4980) );
  NOR2_X1 U6149 ( .A1(n4981), .A2(n4980), .ZN(n4982) );
  XNOR2_X1 U6150 ( .A(n4978), .B(n4982), .ZN(n6214) );
  AOI22_X1 U6151 ( .A1(n6196), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6218), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n4983) );
  OAI21_X1 U6152 ( .B1(n5456), .B2(n6188), .A(n4983), .ZN(n4984) );
  AOI21_X1 U6153 ( .B1(n4985), .B2(n6183), .A(n4984), .ZN(n4986) );
  OAI21_X1 U6154 ( .B1(n6214), .B2(n6190), .A(n4986), .ZN(U2976) );
  NAND2_X1 U6155 ( .A1(n4988), .A2(n4987), .ZN(n4989) );
  NAND2_X1 U6156 ( .A1(n5993), .A2(n4989), .ZN(n6220) );
  INV_X1 U6157 ( .A(EBX_REG_10__SCAN_IN), .ZN(n4990) );
  OAI222_X1 U6158 ( .A1(n6220), .A2(n6090), .B1(n6094), .B2(n4990), .C1(n6085), 
        .C2(n5465), .ZN(U2849) );
  NAND2_X1 U6159 ( .A1(n4992), .A2(n4991), .ZN(n4993) );
  AND2_X1 U6160 ( .A1(n5008), .A2(n4993), .ZN(n6158) );
  INV_X1 U6161 ( .A(n6158), .ZN(n4995) );
  AOI22_X1 U6162 ( .A1(n5557), .A2(DATAI_11_), .B1(n6608), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n4994) );
  OAI21_X1 U6163 ( .B1(n4995), .B2(n5857), .A(n4994), .ZN(U2880) );
  XNOR2_X1 U6164 ( .A(n5890), .B(n6234), .ZN(n4996) );
  XNOR2_X1 U6165 ( .A(n4997), .B(n4996), .ZN(n6225) );
  NAND2_X1 U6166 ( .A1(n6218), .A2(REIP_REG_9__SCAN_IN), .ZN(n6227) );
  OAI21_X1 U6167 ( .B1(n6174), .B2(n6006), .A(n6227), .ZN(n4999) );
  NOR2_X1 U6168 ( .A1(n6010), .A2(n6199), .ZN(n4998) );
  AOI211_X1 U6169 ( .C1(n6168), .C2(n6011), .A(n4999), .B(n4998), .ZN(n5000)
         );
  OAI21_X1 U6170 ( .B1(n6225), .B2(n6190), .A(n5000), .ZN(U2977) );
  INV_X1 U6171 ( .A(n6054), .ZN(n6072) );
  OAI21_X1 U6172 ( .B1(n6034), .B2(n6053), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5001) );
  OAI21_X1 U6173 ( .B1(n6059), .B2(n6373), .A(n5001), .ZN(n5004) );
  NAND2_X1 U6174 ( .A1(n6046), .A2(n6026), .ZN(n6028) );
  INV_X1 U6175 ( .A(n6028), .ZN(n5321) );
  OAI22_X1 U6176 ( .A1(n6048), .A2(n5002), .B1(n5321), .B2(n6586), .ZN(n5003)
         );
  AOI211_X1 U6177 ( .C1(n6051), .C2(EBX_REG_0__SCAN_IN), .A(n5004), .B(n5003), 
        .ZN(n5005) );
  OAI21_X1 U6178 ( .B1(n6072), .B2(n6200), .A(n5005), .ZN(U2827) );
  AOI21_X1 U6179 ( .B1(n5009), .B2(n5008), .A(n5007), .ZN(n5022) );
  INV_X1 U6180 ( .A(n5022), .ZN(n5452) );
  INV_X1 U6181 ( .A(DATAI_12_), .ZN(n5011) );
  OAI222_X1 U6182 ( .A1(n5452), .A2(n5857), .B1(n5293), .B2(n5012), .C1(n5011), 
        .C2(n5010), .ZN(U2879) );
  OR2_X1 U6183 ( .A1(n5007), .A2(n5014), .ZN(n5015) );
  NAND2_X1 U6184 ( .A1(n5256), .A2(n5015), .ZN(n6086) );
  AOI22_X1 U6185 ( .A1(n5557), .A2(DATAI_13_), .B1(n6608), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5016) );
  OAI21_X1 U6186 ( .B1(n6086), .B2(n5857), .A(n5016), .ZN(U2878) );
  XNOR2_X1 U6187 ( .A(n5890), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5018)
         );
  XNOR2_X1 U6188 ( .A(n5019), .B(n5018), .ZN(n5035) );
  NAND2_X1 U6189 ( .A1(n6218), .A2(REIP_REG_12__SCAN_IN), .ZN(n5027) );
  NAND2_X1 U6190 ( .A1(n6196), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5020)
         );
  OAI211_X1 U6191 ( .C1(n6188), .C2(n5445), .A(n5027), .B(n5020), .ZN(n5021)
         );
  AOI21_X1 U6192 ( .B1(n5022), .B2(n6183), .A(n5021), .ZN(n5023) );
  OAI21_X1 U6193 ( .B1(n5035), .B2(n6190), .A(n5023), .ZN(U2974) );
  INV_X1 U6194 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6209) );
  OAI21_X1 U6195 ( .B1(n5025), .B2(n5024), .A(n6209), .ZN(n5026) );
  AOI21_X1 U6196 ( .B1(n6210), .B2(n5026), .A(n5240), .ZN(n5033) );
  INV_X1 U6197 ( .A(n5027), .ZN(n5032) );
  OR2_X1 U6198 ( .A1(n5994), .A2(n5028), .ZN(n5029) );
  NAND2_X1 U6199 ( .A1(n5927), .A2(n5029), .ZN(n5444) );
  NOR2_X1 U6200 ( .A1(n5444), .A2(n6229), .ZN(n5031) );
  NOR3_X1 U6201 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n6201), .A3(n6209), 
        .ZN(n5030) );
  NOR4_X1 U6202 ( .A1(n5033), .A2(n5032), .A3(n5031), .A4(n5030), .ZN(n5034)
         );
  OAI21_X1 U6203 ( .B1(n5035), .B2(n6203), .A(n5034), .ZN(U3006) );
  INV_X1 U6204 ( .A(EBX_REG_12__SCAN_IN), .ZN(n5036) );
  OAI222_X1 U6205 ( .A1(n5444), .A2(n6090), .B1(n6094), .B2(n5036), .C1(n5533), 
        .C2(n5452), .ZN(U2847) );
  INV_X1 U6206 ( .A(n5046), .ZN(n5037) );
  AOI21_X1 U6207 ( .B1(n5038), .B2(n5037), .A(n5941), .ZN(n5048) );
  NOR2_X1 U6208 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n6571), .ZN(n5045)
         );
  INV_X1 U6209 ( .A(n5039), .ZN(n5041) );
  NOR2_X1 U6210 ( .A1(n5041), .A2(n5040), .ZN(n5044) );
  NOR2_X1 U6211 ( .A1(n5042), .A2(n6583), .ZN(n5043) );
  AOI211_X1 U6212 ( .C1(n5046), .C2(n5045), .A(n5044), .B(n5043), .ZN(n5047)
         );
  OAI22_X1 U6213 ( .A1(n5048), .A2(n3237), .B1(n5941), .B2(n5047), .ZN(U3459)
         );
  XNOR2_X1 U6214 ( .A(n5049), .B(n5050), .ZN(n5064) );
  NAND2_X1 U6215 ( .A1(n6218), .A2(REIP_REG_4__SCAN_IN), .ZN(n5059) );
  NAND2_X1 U6216 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n5051), .ZN(n5052)
         );
  NAND2_X1 U6217 ( .A1(n5059), .A2(n5052), .ZN(n5057) );
  INV_X1 U6218 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n5055) );
  AOI211_X1 U6219 ( .C1(n5055), .C2(n3367), .A(n5054), .B(n5053), .ZN(n5056)
         );
  AOI211_X1 U6220 ( .C1(n6240), .C2(n6063), .A(n5057), .B(n5056), .ZN(n5058)
         );
  OAI21_X1 U6221 ( .B1(n6203), .B2(n5064), .A(n5058), .ZN(U3014) );
  NAND2_X1 U6222 ( .A1(n6196), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n5060)
         );
  OAI211_X1 U6223 ( .C1(n6188), .C2(n6071), .A(n5060), .B(n5059), .ZN(n5061)
         );
  AOI21_X1 U6224 ( .B1(n5062), .B2(n6183), .A(n5061), .ZN(n5063) );
  OAI21_X1 U6225 ( .B1(n5064), .B2(n6190), .A(n5063), .ZN(U2982) );
  NAND2_X1 U6226 ( .A1(n5560), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5067) );
  NAND2_X1 U6227 ( .A1(n5589), .A2(n5065), .ZN(n5561) );
  NAND2_X1 U6228 ( .A1(n5067), .A2(n5066), .ZN(n5068) );
  XNOR2_X2 U6229 ( .A(n5073), .B(n5072), .ZN(n5506) );
  NAND2_X1 U6230 ( .A1(n5506), .A2(n6240), .ZN(n5074) );
  NAND2_X1 U6231 ( .A1(n6218), .A2(REIP_REG_30__SCAN_IN), .ZN(n5212) );
  OAI211_X1 U6232 ( .C1(INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n5075), .A(n5074), .B(n5212), .ZN(n5076) );
  AOI21_X1 U6233 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5077), .A(n5076), 
        .ZN(n5078) );
  OAI21_X1 U6234 ( .B1(n5216), .B2(n6203), .A(n5078), .ZN(U2988) );
  AOI22_X1 U6235 ( .A1(n5145), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n5082) );
  AOI22_X1 U6236 ( .A1(n5147), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n5081) );
  AOI22_X1 U6237 ( .A1(n5146), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n5149), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n5080) );
  AOI22_X1 U6238 ( .A1(n5138), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n5079) );
  NAND4_X1 U6239 ( .A1(n5082), .A2(n5081), .A3(n5080), .A4(n5079), .ZN(n5089)
         );
  AOI22_X1 U6240 ( .A1(n3734), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n5087) );
  AOI22_X1 U6241 ( .A1(n5139), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n5086) );
  AOI22_X1 U6242 ( .A1(n3027), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n5085) );
  AOI22_X1 U6243 ( .A1(n5137), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5084) );
  NAND4_X1 U6244 ( .A1(n5087), .A2(n5086), .A3(n5085), .A4(n5084), .ZN(n5088)
         );
  NOR2_X1 U6245 ( .A1(n5089), .A2(n5088), .ZN(n5204) );
  AOI22_X1 U6246 ( .A1(n3734), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n5093) );
  AOI22_X1 U6247 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n5147), .B1(n5083), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5092) );
  AOI22_X1 U6248 ( .A1(n5146), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n5149), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n5091) );
  AOI22_X1 U6249 ( .A1(n5138), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n5090) );
  NAND4_X1 U6250 ( .A1(n5093), .A2(n5092), .A3(n5091), .A4(n5090), .ZN(n5099)
         );
  AOI22_X1 U6251 ( .A1(n5145), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n5097) );
  AOI22_X1 U6252 ( .A1(n5139), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n5096) );
  AOI22_X1 U6253 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n5148), .B1(n3027), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n5095) );
  AOI22_X1 U6254 ( .A1(n5137), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3273), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n5094) );
  NAND4_X1 U6255 ( .A1(n5097), .A2(n5096), .A3(n5095), .A4(n5094), .ZN(n5098)
         );
  NOR2_X1 U6256 ( .A1(n5099), .A2(n5098), .ZN(n5183) );
  AOI22_X1 U6257 ( .A1(n3734), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n5104) );
  AOI22_X1 U6258 ( .A1(n3027), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n5103) );
  AOI22_X1 U6259 ( .A1(n5100), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n5083), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5102) );
  AOI22_X1 U6260 ( .A1(n3273), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n5101) );
  NAND4_X1 U6261 ( .A1(n5104), .A2(n5103), .A3(n5102), .A4(n5101), .ZN(n5111)
         );
  AOI22_X1 U6262 ( .A1(n5145), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n5105), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n5109) );
  AOI22_X1 U6263 ( .A1(n5138), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n5108) );
  AOI22_X1 U6264 ( .A1(n5139), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n5147), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n5107) );
  AOI22_X1 U6265 ( .A1(n5146), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n5149), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n5106) );
  NAND4_X1 U6266 ( .A1(n5109), .A2(n5108), .A3(n5107), .A4(n5106), .ZN(n5110)
         );
  NOR2_X1 U6267 ( .A1(n5111), .A2(n5110), .ZN(n5165) );
  NAND2_X1 U6268 ( .A1(n5113), .A2(n5112), .ZN(n5164) );
  NOR2_X1 U6269 ( .A1(n5165), .A2(n5164), .ZN(n5175) );
  AOI22_X1 U6270 ( .A1(n3734), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n5117) );
  AOI22_X1 U6271 ( .A1(n5145), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n5116) );
  AOI22_X1 U6272 ( .A1(n5139), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n5115) );
  AOI22_X1 U6273 ( .A1(n5147), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5114) );
  NAND4_X1 U6274 ( .A1(n5117), .A2(n5116), .A3(n5115), .A4(n5114), .ZN(n5123)
         );
  AOI22_X1 U6275 ( .A1(n5138), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n5121) );
  AOI22_X1 U6276 ( .A1(n3027), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n5120) );
  AOI22_X1 U6277 ( .A1(n5146), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3291), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n5119) );
  AOI22_X1 U6278 ( .A1(n5149), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n5118) );
  NAND4_X1 U6279 ( .A1(n5121), .A2(n5120), .A3(n5119), .A4(n5118), .ZN(n5122)
         );
  OR2_X1 U6280 ( .A1(n5123), .A2(n5122), .ZN(n5174) );
  NAND2_X1 U6281 ( .A1(n5175), .A2(n5174), .ZN(n5182) );
  NOR2_X1 U6282 ( .A1(n5183), .A2(n5182), .ZN(n5193) );
  AOI22_X1 U6283 ( .A1(n3734), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n5128) );
  AOI22_X1 U6284 ( .A1(n5145), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n5127) );
  AOI22_X1 U6285 ( .A1(n5139), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n5126) );
  AOI22_X1 U6286 ( .A1(n5147), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3289), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5125) );
  NAND4_X1 U6287 ( .A1(n5128), .A2(n5127), .A3(n5126), .A4(n5125), .ZN(n5135)
         );
  AOI22_X1 U6288 ( .A1(n5138), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n5133) );
  AOI22_X1 U6289 ( .A1(n3027), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n5132) );
  AOI22_X1 U6290 ( .A1(n5146), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3291), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n5131) );
  AOI22_X1 U6291 ( .A1(n5149), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n5129), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n5130) );
  NAND4_X1 U6292 ( .A1(n5133), .A2(n5132), .A3(n5131), .A4(n5130), .ZN(n5134)
         );
  OR2_X1 U6293 ( .A1(n5135), .A2(n5134), .ZN(n5192) );
  NAND2_X1 U6294 ( .A1(n5193), .A2(n5192), .ZN(n5203) );
  NOR2_X1 U6295 ( .A1(n5204), .A2(n5203), .ZN(n5157) );
  AOI22_X1 U6296 ( .A1(n3734), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n5136), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n5143) );
  AOI22_X1 U6297 ( .A1(n5138), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n5137), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n5142) );
  AOI22_X1 U6298 ( .A1(n5139), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n5100), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n5141) );
  AOI22_X1 U6299 ( .A1(n5083), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3291), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n5140) );
  NAND4_X1 U6300 ( .A1(n5143), .A2(n5142), .A3(n5141), .A4(n5140), .ZN(n5155)
         );
  AOI22_X1 U6301 ( .A1(n5145), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n5144), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n5153) );
  AOI22_X1 U6302 ( .A1(n5147), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n5146), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n5152) );
  AOI22_X1 U6303 ( .A1(n3027), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n5148), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n5151) );
  AOI22_X1 U6304 ( .A1(n5149), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3250), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n5150) );
  NAND4_X1 U6305 ( .A1(n5153), .A2(n5152), .A3(n5151), .A4(n5150), .ZN(n5154)
         );
  NOR2_X1 U6306 ( .A1(n5155), .A2(n5154), .ZN(n5156) );
  XNOR2_X1 U6307 ( .A(n5157), .B(n5156), .ZN(n5159) );
  NAND2_X1 U6308 ( .A1(n5159), .A2(n5158), .ZN(n5163) );
  AOI21_X1 U6309 ( .B1(n5323), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n5160) );
  AOI21_X1 U6310 ( .B1(n3888), .B2(EAX_REG_30__SCAN_IN), .A(n5160), .ZN(n5162)
         );
  XNOR2_X1 U6311 ( .A(n5202), .B(n5323), .ZN(n5322) );
  INV_X1 U6312 ( .A(n5322), .ZN(n5161) );
  AOI22_X1 U6313 ( .A1(n5163), .A2(n5162), .B1(n5205), .B2(n5161), .ZN(n5274)
         );
  XNOR2_X1 U6314 ( .A(n5165), .B(n5164), .ZN(n5168) );
  INV_X1 U6315 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5351) );
  AOI21_X1 U6316 ( .B1(n5351), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n5166) );
  AOI21_X1 U6317 ( .B1(n3888), .B2(EAX_REG_25__SCAN_IN), .A(n5166), .ZN(n5167)
         );
  OAI21_X1 U6318 ( .B1(n5168), .B2(n5208), .A(n5167), .ZN(n5172) );
  OR2_X1 U6319 ( .A1(n5169), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5170)
         );
  NAND2_X1 U6320 ( .A1(n5179), .A2(n5170), .ZN(n5881) );
  XNOR2_X1 U6321 ( .A(n5175), .B(n5174), .ZN(n5178) );
  OAI21_X1 U6322 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5590), .A(n5211), .ZN(
        n5176) );
  AOI21_X1 U6323 ( .B1(n3888), .B2(EAX_REG_26__SCAN_IN), .A(n5176), .ZN(n5177)
         );
  OAI21_X1 U6324 ( .B1(n5178), .B2(n5208), .A(n5177), .ZN(n5181) );
  XNOR2_X1 U6325 ( .A(n5179), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5803)
         );
  NAND2_X1 U6326 ( .A1(n5803), .A2(n5205), .ZN(n5180) );
  NAND2_X1 U6327 ( .A1(n5181), .A2(n5180), .ZN(n5518) );
  XNOR2_X1 U6328 ( .A(n5183), .B(n5182), .ZN(n5186) );
  OAI21_X1 U6329 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5580), .A(n5211), .ZN(
        n5184) );
  AOI21_X1 U6330 ( .B1(n3888), .B2(EAX_REG_27__SCAN_IN), .A(n5184), .ZN(n5185)
         );
  OAI21_X1 U6331 ( .B1(n5186), .B2(n5208), .A(n5185), .ZN(n5190) );
  NAND2_X1 U6332 ( .A1(n5187), .A2(n5580), .ZN(n5188) );
  NAND2_X1 U6333 ( .A1(n5197), .A2(n5188), .ZN(n5795) );
  INV_X1 U6334 ( .A(n5795), .ZN(n5583) );
  NAND2_X1 U6335 ( .A1(n5583), .A2(n5205), .ZN(n5189) );
  NAND2_X1 U6336 ( .A1(n5190), .A2(n5189), .ZN(n5510) );
  AND2_X2 U6337 ( .A1(n5508), .A2(n5191), .ZN(n5511) );
  XNOR2_X1 U6338 ( .A(n5193), .B(n5192), .ZN(n5196) );
  OAI21_X1 U6339 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5572), .A(n5211), .ZN(
        n5194) );
  AOI21_X1 U6340 ( .B1(n3888), .B2(EAX_REG_28__SCAN_IN), .A(n5194), .ZN(n5195)
         );
  OAI21_X1 U6341 ( .B1(n5196), .B2(n5208), .A(n5195), .ZN(n5199) );
  XNOR2_X1 U6342 ( .A(n5197), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5785)
         );
  NAND2_X1 U6343 ( .A1(n5785), .A2(n5205), .ZN(n5198) );
  AND2_X1 U6344 ( .A1(n5199), .A2(n5198), .ZN(n5289) );
  OR2_X1 U6346 ( .A1(n5200), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5201)
         );
  NAND2_X1 U6347 ( .A1(n5202), .A2(n5201), .ZN(n5566) );
  XNOR2_X1 U6348 ( .A(n5204), .B(n5203), .ZN(n5209) );
  AOI21_X1 U6349 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6486), .A(n5205), 
        .ZN(n5207) );
  NAND2_X1 U6350 ( .A1(n5276), .A2(EAX_REG_29__SCAN_IN), .ZN(n5206) );
  OAI211_X1 U6351 ( .C1(n5209), .C2(n5208), .A(n5207), .B(n5206), .ZN(n5210)
         );
  OAI21_X1 U6352 ( .B1(n5211), .B2(n5566), .A(n5210), .ZN(n5332) );
  NOR2_X1 U6353 ( .A1(n6188), .A2(n5322), .ZN(n5214) );
  OAI21_X1 U6354 ( .B1(n6174), .B2(n5323), .A(n5212), .ZN(n5213) );
  AOI211_X1 U6355 ( .C1(n5319), .C2(n6183), .A(n5214), .B(n5213), .ZN(n5215)
         );
  OAI21_X1 U6356 ( .B1(n5216), .B2(n6190), .A(n5215), .ZN(U2956) );
  NAND2_X1 U6357 ( .A1(n5228), .A2(n5217), .ZN(n5218) );
  NAND2_X1 U6358 ( .A1(n5348), .A2(n5218), .ZN(n5814) );
  INV_X1 U6359 ( .A(n5814), .ZN(n5224) );
  INV_X1 U6360 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5221) );
  INV_X1 U6361 ( .A(n5268), .ZN(n5219) );
  NAND3_X1 U6362 ( .A1(n5219), .A2(n5231), .A3(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5220) );
  AOI21_X1 U6363 ( .B1(n5221), .B2(n5220), .A(n5906), .ZN(n5222) );
  AOI211_X1 U6364 ( .C1(n6240), .C2(n5224), .A(n5223), .B(n5222), .ZN(n5225)
         );
  OAI21_X1 U6365 ( .B1(n5226), .B2(n6203), .A(n5225), .ZN(U2994) );
  INV_X1 U6366 ( .A(n5227), .ZN(n5237) );
  INV_X1 U6367 ( .A(n5228), .ZN(n5229) );
  AOI21_X1 U6368 ( .B1(n5230), .B2(n5369), .A(n5229), .ZN(n5848) );
  INV_X1 U6369 ( .A(n5231), .ZN(n5232) );
  NOR3_X1 U6370 ( .A1(n5268), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n5232), 
        .ZN(n5233) );
  AOI211_X1 U6371 ( .C1(n6240), .C2(n5848), .A(n5234), .B(n5233), .ZN(n5236)
         );
  NAND2_X1 U6372 ( .A1(n5682), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5235) );
  OAI211_X1 U6373 ( .C1(n5237), .C2(n6203), .A(n5236), .B(n5235), .ZN(U2995)
         );
  XNOR2_X1 U6374 ( .A(n5890), .B(n5721), .ZN(n5239) );
  XNOR2_X1 U6375 ( .A(n5238), .B(n5239), .ZN(n5262) );
  NOR2_X1 U6376 ( .A1(n6209), .A2(n5240), .ZN(n5245) );
  OAI21_X1 U6377 ( .B1(n5241), .B2(n5245), .A(n6210), .ZN(n5242) );
  AOI21_X1 U6378 ( .B1(n5936), .B2(n5722), .A(n5242), .ZN(n5931) );
  NOR3_X1 U6379 ( .A1(n6577), .A2(n5244), .A3(n5243), .ZN(n5246) );
  INV_X1 U6380 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5930) );
  AND2_X1 U6381 ( .A1(n5930), .A2(n5245), .ZN(n5934) );
  OAI21_X1 U6382 ( .B1(n5247), .B2(n5246), .A(n5934), .ZN(n5939) );
  AOI21_X1 U6383 ( .B1(n5931), .B2(n5939), .A(n5721), .ZN(n5253) );
  NAND2_X1 U6384 ( .A1(n6218), .A2(REIP_REG_14__SCAN_IN), .ZN(n5259) );
  INV_X1 U6385 ( .A(n5259), .ZN(n5252) );
  NAND2_X1 U6386 ( .A1(n5929), .A2(n5248), .ZN(n5249) );
  NAND2_X1 U6387 ( .A1(n5425), .A2(n5249), .ZN(n5540) );
  NOR2_X1 U6388 ( .A1(n5540), .A2(n6229), .ZN(n5251) );
  NOR3_X1 U6389 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6201), .A3(n5722), 
        .ZN(n5250) );
  NOR4_X1 U6390 ( .A1(n5253), .A2(n5252), .A3(n5251), .A4(n5250), .ZN(n5254)
         );
  OAI21_X1 U6391 ( .B1(n5262), .B2(n6203), .A(n5254), .ZN(U3004) );
  INV_X1 U6392 ( .A(n5422), .ZN(n5255) );
  AOI21_X1 U6393 ( .B1(n5257), .B2(n5256), .A(n5255), .ZN(n5434) );
  NAND2_X1 U6394 ( .A1(n6196), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5258)
         );
  OAI211_X1 U6395 ( .C1(n6188), .C2(n5435), .A(n5259), .B(n5258), .ZN(n5260)
         );
  AOI21_X1 U6396 ( .B1(n5434), .B2(n6183), .A(n5260), .ZN(n5261) );
  OAI21_X1 U6397 ( .B1(n5262), .B2(n6190), .A(n5261), .ZN(U2972) );
  INV_X1 U6398 ( .A(n5263), .ZN(n5273) );
  NOR2_X1 U6399 ( .A1(n5265), .A2(n5264), .ZN(n5266) );
  OR2_X1 U6400 ( .A1(n5367), .A2(n5266), .ZN(n5850) );
  OAI21_X1 U6401 ( .B1(n5850), .B2(n6229), .A(n5267), .ZN(n5270) );
  NOR2_X1 U6402 ( .A1(n5268), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5269)
         );
  AOI211_X1 U6403 ( .C1(INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n5271), .A(n5270), .B(n5269), .ZN(n5272) );
  OAI21_X1 U6404 ( .B1(n5273), .B2(n6203), .A(n5272), .ZN(U2997) );
  NAND2_X1 U6405 ( .A1(n5330), .A2(n5274), .ZN(n5279) );
  AOI22_X1 U6406 ( .A1(n5276), .A2(EAX_REG_31__SCAN_IN), .B1(n5275), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5277) );
  INV_X1 U6407 ( .A(n5277), .ZN(n5278) );
  NAND2_X1 U6408 ( .A1(n6196), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5280)
         );
  OAI211_X1 U6409 ( .C1(n6188), .C2(n5282), .A(n5281), .B(n5280), .ZN(n5283)
         );
  AOI21_X1 U6410 ( .B1(n5299), .B2(n6183), .A(n5283), .ZN(n5284) );
  OAI21_X1 U6411 ( .B1(n5285), .B2(n6190), .A(n5284), .ZN(U2955) );
  NAND3_X1 U6412 ( .A1(n5299), .A2(n5286), .A3(n5293), .ZN(n5288) );
  AOI22_X1 U6413 ( .A1(n6610), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6608), .ZN(n5287) );
  NAND2_X1 U6414 ( .A1(n5288), .A2(n5287), .ZN(U2860) );
  OR2_X1 U6415 ( .A1(n5511), .A2(n5289), .ZN(n5290) );
  AND2_X1 U6416 ( .A1(n3207), .A2(n5291), .ZN(n5292) );
  AOI22_X1 U6417 ( .A1(n6609), .A2(DATAI_12_), .B1(n6608), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5295) );
  NAND2_X1 U6418 ( .A1(n6610), .A2(DATAI_28_), .ZN(n5294) );
  OAI211_X1 U6419 ( .C1(n5789), .C2(n5857), .A(n5295), .B(n5294), .ZN(U2863)
         );
  INV_X1 U6420 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5298) );
  OR2_X1 U6421 ( .A1(n5516), .A2(n5296), .ZN(n5297) );
  NAND2_X1 U6422 ( .A1(n5069), .A2(n5297), .ZN(n5788) );
  OAI222_X1 U6423 ( .A1(n6085), .A2(n5789), .B1(n6094), .B2(n5298), .C1(n5788), 
        .C2(n6090), .ZN(U2831) );
  INV_X1 U6424 ( .A(n5299), .ZN(n5318) );
  INV_X1 U6425 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5300) );
  INV_X1 U6426 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6529) );
  INV_X1 U6427 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6527) );
  NAND3_X1 U6428 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6045) );
  INV_X1 U6429 ( .A(n6045), .ZN(n5484) );
  NAND3_X1 U6430 ( .A1(n5484), .A2(REIP_REG_5__SCAN_IN), .A3(
        REIP_REG_4__SCAN_IN), .ZN(n6024) );
  NAND3_X1 U6431 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_6__SCAN_IN), .ZN(n5461) );
  NOR2_X1 U6432 ( .A1(n6024), .A2(n5461), .ZN(n5462) );
  NAND2_X1 U6433 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5462), .ZN(n5453) );
  NOR3_X1 U6434 ( .A1(n6529), .A2(n6527), .A3(n5453), .ZN(n5446) );
  NAND4_X1 U6435 ( .A1(REIP_REG_14__SCAN_IN), .A2(n5446), .A3(
        REIP_REG_13__SCAN_IN), .A4(REIP_REG_12__SCAN_IN), .ZN(n5410) );
  NOR2_X1 U6436 ( .A1(n5300), .A2(n5410), .ZN(n5413) );
  NAND2_X1 U6437 ( .A1(REIP_REG_16__SCAN_IN), .A2(n5413), .ZN(n5306) );
  NOR2_X1 U6438 ( .A1(n6046), .A2(n5306), .ZN(n5970) );
  NAND2_X1 U6439 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5970), .ZN(n5839) );
  INV_X1 U6440 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6542) );
  INV_X1 U6441 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6540) );
  NOR2_X1 U6442 ( .A1(n6542), .A2(n6540), .ZN(n5309) );
  INV_X1 U6443 ( .A(n5309), .ZN(n5837) );
  NOR2_X1 U6444 ( .A1(n5839), .A2(n5837), .ZN(n5379) );
  NAND2_X1 U6445 ( .A1(REIP_REG_20__SCAN_IN), .A2(n5379), .ZN(n5828) );
  NAND2_X1 U6446 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5363) );
  NOR2_X1 U6447 ( .A1(n5828), .A2(n5363), .ZN(n5820) );
  NAND2_X1 U6448 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5820), .ZN(n5819) );
  NAND3_X1 U6449 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5312) );
  NOR2_X1 U6450 ( .A1(n5819), .A2(n5312), .ZN(n5797) );
  NAND3_X1 U6451 ( .A1(n5797), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_27__SCAN_IN), .ZN(n5338) );
  INV_X1 U6452 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6562) );
  INV_X1 U6453 ( .A(REIP_REG_29__SCAN_IN), .ZN(n5564) );
  NOR4_X1 U6454 ( .A1(n5338), .A2(REIP_REG_31__SCAN_IN), .A3(n6562), .A4(n5564), .ZN(n5305) );
  OAI22_X1 U6455 ( .A1(n5303), .A2(n6069), .B1(n5302), .B2(n5301), .ZN(n5304)
         );
  AOI211_X1 U6456 ( .C1(n5502), .C2(n6064), .A(n5305), .B(n5304), .ZN(n5317)
         );
  INV_X1 U6457 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6538) );
  NOR2_X1 U6458 ( .A1(n6538), .A2(n5306), .ZN(n5307) );
  NAND2_X1 U6459 ( .A1(n6026), .A2(n5307), .ZN(n5308) );
  NAND2_X1 U6460 ( .A1(n6028), .A2(n5308), .ZN(n5973) );
  NAND2_X1 U6461 ( .A1(n5309), .A2(REIP_REG_20__SCAN_IN), .ZN(n5310) );
  NAND2_X1 U6462 ( .A1(n5460), .A2(n5310), .ZN(n5311) );
  NAND2_X1 U6463 ( .A1(n5973), .A2(n5311), .ZN(n5831) );
  AOI221_X1 U6464 ( .B1(n4126), .B2(n6028), .C1(n5363), .C2(n6028), .A(n5831), 
        .ZN(n5827) );
  NAND2_X1 U6465 ( .A1(n6028), .A2(n5312), .ZN(n5313) );
  NAND2_X1 U6466 ( .A1(n5827), .A2(n5313), .ZN(n5809) );
  AND2_X1 U6467 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5314) );
  NOR2_X1 U6468 ( .A1(n6046), .A2(n5314), .ZN(n5315) );
  NOR2_X1 U6469 ( .A1(n5809), .A2(n5315), .ZN(n5787) );
  AND2_X1 U6470 ( .A1(n5787), .A2(REIP_REG_29__SCAN_IN), .ZN(n5320) );
  INV_X1 U6471 ( .A(n5320), .ZN(n5339) );
  OAI211_X1 U6472 ( .C1(n5339), .C2(n6562), .A(REIP_REG_31__SCAN_IN), .B(n6028), .ZN(n5316) );
  OAI211_X1 U6473 ( .C1(n5318), .C2(n6039), .A(n5317), .B(n5316), .ZN(U2796)
         );
  NOR3_X1 U6474 ( .A1(n5338), .A2(REIP_REG_30__SCAN_IN), .A3(n5564), .ZN(n5328) );
  NOR3_X1 U6475 ( .A1(n5321), .A2(n5320), .A3(n6562), .ZN(n5325) );
  OAI22_X1 U6476 ( .A1(n5323), .A2(n6069), .B1(n5322), .B2(n6070), .ZN(n5324)
         );
  AOI211_X1 U6477 ( .C1(n6051), .C2(EBX_REG_30__SCAN_IN), .A(n5325), .B(n5324), 
        .ZN(n5326) );
  INV_X1 U6478 ( .A(n5326), .ZN(n5327) );
  AOI211_X1 U6479 ( .C1(n5506), .C2(n6064), .A(n5328), .B(n5327), .ZN(n5329)
         );
  OAI21_X1 U6480 ( .B1(n5543), .B2(n6039), .A(n5329), .ZN(U2797) );
  AOI21_X1 U6481 ( .B1(n5332), .B2(n5331), .A(n5330), .ZN(n5568) );
  INV_X1 U6482 ( .A(n5568), .ZN(n5546) );
  INV_X1 U6483 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5333) );
  OAI22_X1 U6484 ( .A1(n5333), .A2(n6069), .B1(n6070), .B2(n5566), .ZN(n5337)
         );
  INV_X1 U6485 ( .A(n5334), .ZN(n5335) );
  NOR2_X1 U6486 ( .A1(n5643), .A2(n6048), .ZN(n5336) );
  AOI211_X1 U6487 ( .C1(n6051), .C2(EBX_REG_29__SCAN_IN), .A(n5337), .B(n5336), 
        .ZN(n5342) );
  INV_X1 U6488 ( .A(n5338), .ZN(n5340) );
  OAI21_X1 U6489 ( .B1(REIP_REG_29__SCAN_IN), .B2(n5340), .A(n5339), .ZN(n5341) );
  OAI211_X1 U6490 ( .C1(n5546), .C2(n6039), .A(n5342), .B(n5341), .ZN(U2798)
         );
  INV_X1 U6491 ( .A(n5343), .ZN(n5346) );
  INV_X1 U6492 ( .A(n5173), .ZN(n5345) );
  INV_X1 U6493 ( .A(n5344), .ZN(n5520) );
  AOI21_X1 U6494 ( .B1(n5346), .B2(n5345), .A(n5520), .ZN(n5878) );
  INV_X1 U6495 ( .A(n5878), .ZN(n5553) );
  INV_X1 U6496 ( .A(n5522), .ZN(n5350) );
  NAND2_X1 U6497 ( .A1(n5348), .A2(n5347), .ZN(n5349) );
  NAND2_X1 U6498 ( .A1(n5350), .A2(n5349), .ZN(n5901) );
  OAI21_X1 U6499 ( .B1(REIP_REG_24__SCAN_IN), .B2(n5819), .A(n5827), .ZN(n5353) );
  OAI22_X1 U6500 ( .A1(n5351), .A2(n6069), .B1(n5881), .B2(n6070), .ZN(n5352)
         );
  AOI21_X1 U6501 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5353), .A(n5352), .ZN(n5355) );
  NAND2_X1 U6502 ( .A1(n6051), .A2(EBX_REG_25__SCAN_IN), .ZN(n5354) );
  OAI211_X1 U6503 ( .C1(n5901), .C2(n6048), .A(n5355), .B(n5354), .ZN(n5357)
         );
  INV_X1 U6504 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6783) );
  NOR3_X1 U6505 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6783), .A3(n5819), .ZN(n5356) );
  NOR2_X1 U6506 ( .A1(n5357), .A2(n5356), .ZN(n5358) );
  OAI21_X1 U6507 ( .B1(n5553), .B2(n6039), .A(n5358), .ZN(U2802) );
  NAND2_X1 U6508 ( .A1(n5360), .A2(n5359), .ZN(n5361) );
  NAND2_X1 U6509 ( .A1(n5362), .A2(n5361), .ZN(n5598) );
  INV_X1 U6510 ( .A(n5598), .ZN(n5861) );
  OAI21_X1 U6511 ( .B1(REIP_REG_22__SCAN_IN), .B2(REIP_REG_21__SCAN_IN), .A(
        n5363), .ZN(n5365) );
  AOI22_X1 U6512 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n6034), .B1(
        REIP_REG_22__SCAN_IN), .B2(n5831), .ZN(n5364) );
  OAI21_X1 U6513 ( .B1(n5828), .B2(n5365), .A(n5364), .ZN(n5372) );
  OR2_X1 U6514 ( .A1(n5367), .A2(n5366), .ZN(n5368) );
  NAND2_X1 U6515 ( .A1(n5369), .A2(n5368), .ZN(n5680) );
  AOI22_X1 U6516 ( .A1(n6051), .A2(EBX_REG_22__SCAN_IN), .B1(n6053), .B2(n5601), .ZN(n5370) );
  OAI21_X1 U6517 ( .B1(n5680), .B2(n6048), .A(n5370), .ZN(n5371) );
  AOI211_X1 U6518 ( .C1(n5861), .C2(n6012), .A(n5372), .B(n5371), .ZN(n5373)
         );
  INV_X1 U6519 ( .A(n5373), .ZN(U2805) );
  NOR2_X1 U6520 ( .A1(n5897), .A2(n5374), .ZN(n5844) );
  NOR2_X1 U6521 ( .A1(n5844), .A2(n5375), .ZN(n5376) );
  INV_X1 U6522 ( .A(n5607), .ZN(n5867) );
  NAND2_X1 U6523 ( .A1(n5867), .A2(n6012), .ZN(n5388) );
  INV_X1 U6524 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5529) );
  OAI22_X1 U6525 ( .A1(n5529), .A2(n6078), .B1(n5606), .B2(n6069), .ZN(n5378)
         );
  AOI21_X1 U6526 ( .B1(n6053), .B2(n5610), .A(n5378), .ZN(n5387) );
  OAI21_X1 U6527 ( .B1(n5379), .B2(REIP_REG_20__SCAN_IN), .A(n5831), .ZN(n5386) );
  MUX2_X1 U6528 ( .A(n5382), .B(n5381), .S(n5380), .Z(n5384) );
  XNOR2_X1 U6529 ( .A(n5384), .B(n5383), .ZN(n5691) );
  NAND2_X1 U6530 ( .A1(n5691), .A2(n6064), .ZN(n5385) );
  NAND4_X1 U6531 ( .A1(n5388), .A2(n5387), .A3(n5386), .A4(n5385), .ZN(U2807)
         );
  INV_X1 U6532 ( .A(n5843), .ZN(n5389) );
  AOI21_X1 U6533 ( .B1(n5390), .B2(n5897), .A(n5389), .ZN(n6096) );
  INV_X1 U6534 ( .A(n6096), .ZN(n5532) );
  NAND2_X1 U6535 ( .A1(n5393), .A2(n5392), .ZN(n5699) );
  XNOR2_X1 U6536 ( .A(n5391), .B(n5699), .ZN(n5715) );
  INV_X1 U6537 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5398) );
  INV_X1 U6538 ( .A(n5620), .ZN(n5396) );
  NAND2_X1 U6539 ( .A1(n6026), .A2(n5394), .ZN(n6066) );
  OAI21_X1 U6540 ( .B1(n6069), .B2(n6758), .A(n6066), .ZN(n5395) );
  AOI21_X1 U6541 ( .B1(n6053), .B2(n5396), .A(n5395), .ZN(n5397) );
  OAI21_X1 U6542 ( .B1(n6078), .B2(n5398), .A(n5397), .ZN(n5400) );
  AOI22_X1 U6543 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5973), .B1(n5839), .B2(
        n6540), .ZN(n5399) );
  AOI211_X1 U6544 ( .C1(n6064), .C2(n5715), .A(n5400), .B(n5399), .ZN(n5401)
         );
  OAI21_X1 U6545 ( .B1(n5532), .B2(n6039), .A(n5401), .ZN(U2809) );
  NOR2_X1 U6546 ( .A1(n5421), .A2(n5403), .ZN(n5404) );
  OR2_X1 U6547 ( .A1(n5895), .A2(n5404), .ZN(n6099) );
  NOR2_X1 U6548 ( .A1(n5427), .A2(n5405), .ZN(n5406) );
  OR2_X1 U6549 ( .A1(n5908), .A2(n5406), .ZN(n5726) );
  INV_X1 U6550 ( .A(n5726), .ZN(n5419) );
  NAND2_X1 U6551 ( .A1(n6034), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5409)
         );
  INV_X1 U6552 ( .A(n5625), .ZN(n5407) );
  NAND2_X1 U6553 ( .A1(n6053), .A2(n5407), .ZN(n5408) );
  NAND3_X1 U6554 ( .A1(n5409), .A2(n5408), .A3(n6066), .ZN(n5418) );
  INV_X1 U6555 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5534) );
  INV_X1 U6556 ( .A(n5410), .ZN(n5411) );
  OAI21_X1 U6557 ( .B1(n6046), .B2(n5411), .A(n6026), .ZN(n5441) );
  NAND2_X1 U6558 ( .A1(n5300), .A2(n5411), .ZN(n5412) );
  NOR2_X1 U6559 ( .A1(n6046), .A2(n5412), .ZN(n5428) );
  OAI21_X1 U6560 ( .B1(n5441), .B2(n5428), .A(REIP_REG_16__SCAN_IN), .ZN(n5416) );
  INV_X1 U6561 ( .A(REIP_REG_16__SCAN_IN), .ZN(n5414) );
  NAND3_X1 U6562 ( .A1(n5460), .A2(n5414), .A3(n5413), .ZN(n5415) );
  OAI211_X1 U6563 ( .C1(n6078), .C2(n5534), .A(n5416), .B(n5415), .ZN(n5417)
         );
  AOI211_X1 U6564 ( .C1(n5419), .C2(n6064), .A(n5418), .B(n5417), .ZN(n5420)
         );
  OAI21_X1 U6565 ( .B1(n6099), .B2(n6039), .A(n5420), .ZN(U2811) );
  AOI21_X1 U6566 ( .B1(n5423), .B2(n5422), .A(n5421), .ZN(n5535) );
  INV_X1 U6567 ( .A(n5535), .ZN(n5634) );
  AND2_X1 U6568 ( .A1(n5425), .A2(n5424), .ZN(n5426) );
  NOR2_X1 U6569 ( .A1(n5427), .A2(n5426), .ZN(n5920) );
  AOI21_X1 U6570 ( .B1(n5631), .B2(n6053), .A(n5428), .ZN(n5429) );
  INV_X1 U6571 ( .A(n5429), .ZN(n5432) );
  AOI22_X1 U6572 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6051), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5441), .ZN(n5430) );
  OAI211_X1 U6573 ( .C1(n6069), .C2(n6771), .A(n5430), .B(n6066), .ZN(n5431)
         );
  AOI211_X1 U6574 ( .C1(n5920), .C2(n6064), .A(n5432), .B(n5431), .ZN(n5433)
         );
  OAI21_X1 U6575 ( .B1(n5634), .B2(n6039), .A(n5433), .ZN(U2812) );
  INV_X1 U6576 ( .A(n5434), .ZN(n5559) );
  NAND2_X1 U6577 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n5979) );
  NAND2_X1 U6578 ( .A1(n5460), .A2(n5446), .ZN(n5981) );
  INV_X1 U6579 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6534) );
  OAI21_X1 U6580 ( .B1(n5979), .B2(n5981), .A(n6534), .ZN(n5442) );
  NOR2_X1 U6581 ( .A1(n6070), .A2(n5435), .ZN(n5438) );
  INV_X1 U6582 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5436) );
  OAI21_X1 U6583 ( .B1(n6069), .B2(n5436), .A(n6066), .ZN(n5437) );
  AOI211_X1 U6584 ( .C1(n6051), .C2(EBX_REG_14__SCAN_IN), .A(n5438), .B(n5437), 
        .ZN(n5439) );
  OAI21_X1 U6585 ( .B1(n5540), .B2(n6048), .A(n5439), .ZN(n5440) );
  AOI21_X1 U6586 ( .B1(n5442), .B2(n5441), .A(n5440), .ZN(n5443) );
  OAI21_X1 U6587 ( .B1(n5559), .B2(n6039), .A(n5443), .ZN(U2813) );
  INV_X1 U6588 ( .A(n5444), .ZN(n5450) );
  OAI22_X1 U6589 ( .A1(n5981), .A2(REIP_REG_12__SCAN_IN), .B1(n5445), .B2(
        n6070), .ZN(n5449) );
  OAI21_X1 U6590 ( .B1(n6046), .B2(n5446), .A(n6026), .ZN(n5991) );
  AOI22_X1 U6591 ( .A1(EBX_REG_12__SCAN_IN), .A2(n6051), .B1(
        REIP_REG_12__SCAN_IN), .B2(n5991), .ZN(n5447) );
  OAI211_X1 U6592 ( .C1(n6069), .C2(n3682), .A(n5447), .B(n6066), .ZN(n5448)
         );
  AOI211_X1 U6593 ( .C1(n5450), .C2(n6064), .A(n5449), .B(n5448), .ZN(n5451)
         );
  OAI21_X1 U6594 ( .B1(n5452), .B2(n6039), .A(n5451), .ZN(U2815) );
  NOR2_X1 U6595 ( .A1(n6046), .A2(n5453), .ZN(n5990) );
  INV_X1 U6596 ( .A(n6066), .ZN(n6050) );
  AOI21_X1 U6597 ( .B1(n6034), .B2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6050), 
        .ZN(n5455) );
  NAND2_X1 U6598 ( .A1(n6051), .A2(EBX_REG_10__SCAN_IN), .ZN(n5454) );
  OAI211_X1 U6599 ( .C1(n6070), .C2(n5456), .A(n5455), .B(n5454), .ZN(n5458)
         );
  NOR2_X1 U6600 ( .A1(n6048), .A2(n6220), .ZN(n5457) );
  AOI211_X1 U6601 ( .C1(n6527), .C2(n5990), .A(n5458), .B(n5457), .ZN(n5464)
         );
  AND3_X1 U6602 ( .A1(REIP_REG_5__SCAN_IN), .A2(REIP_REG_4__SCAN_IN), .A3(
        n5484), .ZN(n5459) );
  NAND2_X1 U6603 ( .A1(n5460), .A2(n5459), .ZN(n6044) );
  NOR3_X1 U6604 ( .A1(REIP_REG_9__SCAN_IN), .A2(n5461), .A3(n6044), .ZN(n6008)
         );
  OAI21_X1 U6605 ( .B1(n6046), .B2(n5462), .A(n6026), .ZN(n6009) );
  OAI21_X1 U6606 ( .B1(n6008), .B2(n6009), .A(REIP_REG_10__SCAN_IN), .ZN(n5463) );
  OAI211_X1 U6607 ( .C1(n5465), .C2(n6039), .A(n5464), .B(n5463), .ZN(U2817)
         );
  NAND2_X1 U6608 ( .A1(REIP_REG_7__SCAN_IN), .A2(REIP_REG_6__SCAN_IN), .ZN(
        n6016) );
  OAI21_X1 U6609 ( .B1(n6016), .B2(n6044), .A(n6524), .ZN(n5473) );
  NOR2_X1 U6610 ( .A1(n6048), .A2(n5466), .ZN(n5472) );
  NOR2_X1 U6611 ( .A1(n6070), .A2(n5467), .ZN(n5468) );
  AOI211_X1 U6612 ( .C1(n6034), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6050), 
        .B(n5468), .ZN(n5469) );
  OAI21_X1 U6613 ( .B1(n5470), .B2(n6078), .A(n5469), .ZN(n5471) );
  AOI211_X1 U6614 ( .C1(n5473), .C2(n6009), .A(n5472), .B(n5471), .ZN(n5474)
         );
  OAI21_X1 U6615 ( .B1(n5475), .B2(n6039), .A(n5474), .ZN(U2819) );
  NAND2_X1 U6616 ( .A1(n5476), .A2(n6054), .ZN(n5488) );
  OAI21_X1 U6617 ( .B1(n6046), .B2(n5484), .A(n6026), .ZN(n6065) );
  INV_X1 U6618 ( .A(EBX_REG_3__SCAN_IN), .ZN(n5481) );
  NAND2_X1 U6619 ( .A1(n6064), .A2(n5477), .ZN(n5480) );
  AOI22_X1 U6620 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n6034), .B1(n6053), 
        .B2(n5478), .ZN(n5479) );
  OAI211_X1 U6621 ( .C1(n5481), .C2(n6078), .A(n5480), .B(n5479), .ZN(n5486)
         );
  AND2_X1 U6622 ( .A1(n6026), .A2(REIP_REG_2__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U6623 ( .A1(n5483), .A2(n5482), .ZN(n5499) );
  NOR3_X1 U6624 ( .A1(n5499), .A2(n6046), .A3(n5484), .ZN(n5485) );
  AOI211_X1 U6625 ( .C1(REIP_REG_3__SCAN_IN), .C2(n6065), .A(n5486), .B(n5485), 
        .ZN(n5487) );
  OAI211_X1 U6626 ( .C1(n5740), .C2(n6059), .A(n5488), .B(n5487), .ZN(U2824)
         );
  INV_X1 U6627 ( .A(REIP_REG_2__SCAN_IN), .ZN(n5489) );
  OAI21_X1 U6628 ( .B1(n6046), .B2(n5490), .A(n5489), .ZN(n5498) );
  INV_X1 U6629 ( .A(n5491), .ZN(n5734) );
  NOR2_X1 U6630 ( .A1(n5734), .A2(n6059), .ZN(n5497) );
  NAND2_X1 U6631 ( .A1(n6064), .A2(n6239), .ZN(n5495) );
  INV_X1 U6632 ( .A(n6187), .ZN(n5492) );
  AOI22_X1 U6633 ( .A1(n6034), .A2(PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n6053), 
        .B2(n5492), .ZN(n5494) );
  NAND2_X1 U6634 ( .A1(n6051), .A2(EBX_REG_2__SCAN_IN), .ZN(n5493) );
  NAND3_X1 U6635 ( .A1(n5495), .A2(n5494), .A3(n5493), .ZN(n5496) );
  AOI211_X1 U6636 ( .C1(n5499), .C2(n5498), .A(n5497), .B(n5496), .ZN(n5500)
         );
  OAI21_X1 U6637 ( .B1(n5501), .B2(n6072), .A(n5500), .ZN(U2825) );
  INV_X1 U6638 ( .A(n5502), .ZN(n5504) );
  INV_X1 U6639 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5503) );
  OAI22_X1 U6640 ( .A1(n5504), .A2(n6090), .B1(n6094), .B2(n5503), .ZN(U2828)
         );
  AOI22_X1 U6641 ( .A1(n5506), .A2(n6081), .B1(EBX_REG_30__SCAN_IN), .B2(n5505), .ZN(n5507) );
  OAI21_X1 U6642 ( .B1(n5543), .B2(n5533), .A(n5507), .ZN(U2829) );
  INV_X1 U6643 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6648) );
  OAI222_X1 U6644 ( .A1(n5546), .A2(n5533), .B1(n6090), .B2(n5643), .C1(n6094), 
        .C2(n6648), .ZN(U2830) );
  INV_X1 U6645 ( .A(n5508), .ZN(n5509) );
  AND2_X1 U6646 ( .A1(n5509), .A2(n5510), .ZN(n5512) );
  OR2_X1 U6647 ( .A1(n5512), .A2(n5511), .ZN(n5799) );
  INV_X1 U6648 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5517) );
  NOR2_X1 U6649 ( .A1(n5513), .A2(n5514), .ZN(n5515) );
  OR2_X1 U6650 ( .A1(n5516), .A2(n5515), .ZN(n5798) );
  OAI222_X1 U6651 ( .A1(n5533), .A2(n5799), .B1(n6094), .B2(n5517), .C1(n5798), 
        .C2(n6090), .ZN(U2832) );
  INV_X1 U6652 ( .A(n5518), .ZN(n5519) );
  NOR2_X1 U6653 ( .A1(n5522), .A2(n5521), .ZN(n5523) );
  OR2_X1 U6654 ( .A1(n5513), .A2(n5523), .ZN(n5805) );
  OAI22_X1 U6655 ( .A1(n5805), .A2(n6090), .B1(n6738), .B2(n6094), .ZN(n5524)
         );
  INV_X1 U6656 ( .A(n5524), .ZN(n5525) );
  OAI21_X1 U6657 ( .B1(n5806), .B2(n5533), .A(n5525), .ZN(U2833) );
  INV_X1 U6658 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5526) );
  OAI222_X1 U6659 ( .A1(n5901), .A2(n6090), .B1(n5526), .B2(n6094), .C1(n5553), 
        .C2(n5533), .ZN(U2834) );
  INV_X1 U6660 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5527) );
  OAI222_X1 U6661 ( .A1(n5533), .A2(n5815), .B1(n6094), .B2(n5527), .C1(n5814), 
        .C2(n6090), .ZN(U2835) );
  INV_X1 U6662 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5528) );
  OAI222_X1 U6663 ( .A1(n6090), .A2(n5680), .B1(n6094), .B2(n5528), .C1(n5598), 
        .C2(n5533), .ZN(U2837) );
  INV_X1 U6664 ( .A(n5691), .ZN(n5530) );
  OAI222_X1 U6665 ( .A1(n5530), .A2(n6090), .B1(n6094), .B2(n5529), .C1(n5533), 
        .C2(n5607), .ZN(U2839) );
  INV_X1 U6666 ( .A(n5715), .ZN(n5531) );
  OAI222_X1 U6667 ( .A1(n5532), .A2(n5533), .B1(n6090), .B2(n5531), .C1(n6094), 
        .C2(n5398), .ZN(U2841) );
  OAI222_X1 U6668 ( .A1(n5726), .A2(n6090), .B1(n6094), .B2(n5534), .C1(n5533), 
        .C2(n6099), .ZN(U2843) );
  INV_X1 U6669 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U6670 ( .A1(n5535), .A2(n6092), .ZN(n5537) );
  NAND2_X1 U6671 ( .A1(n5920), .A2(n6081), .ZN(n5536) );
  OAI211_X1 U6672 ( .C1(n5538), .C2(n6094), .A(n5537), .B(n5536), .ZN(U2844)
         );
  INV_X1 U6673 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5539) );
  OAI222_X1 U6674 ( .A1(n5540), .A2(n6090), .B1(n6094), .B2(n5539), .C1(n6085), 
        .C2(n5559), .ZN(U2845) );
  AOI22_X1 U6675 ( .A1(n6610), .A2(DATAI_30_), .B1(n6608), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5542) );
  NAND2_X1 U6676 ( .A1(n6609), .A2(DATAI_14_), .ZN(n5541) );
  OAI211_X1 U6677 ( .C1(n5543), .C2(n5857), .A(n5542), .B(n5541), .ZN(U2861)
         );
  AOI22_X1 U6678 ( .A1(n6610), .A2(DATAI_29_), .B1(n6608), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5545) );
  NAND2_X1 U6679 ( .A1(n6609), .A2(DATAI_13_), .ZN(n5544) );
  OAI211_X1 U6680 ( .C1(n5546), .C2(n5857), .A(n5545), .B(n5544), .ZN(U2862)
         );
  AOI22_X1 U6681 ( .A1(n6609), .A2(DATAI_11_), .B1(n6608), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5548) );
  NAND2_X1 U6682 ( .A1(n6610), .A2(DATAI_27_), .ZN(n5547) );
  OAI211_X1 U6683 ( .C1(n5799), .C2(n5857), .A(n5548), .B(n5547), .ZN(U2864)
         );
  AOI22_X1 U6684 ( .A1(n6609), .A2(DATAI_10_), .B1(n6608), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U6685 ( .A1(n6610), .A2(DATAI_26_), .ZN(n5549) );
  OAI211_X1 U6686 ( .C1(n5806), .C2(n5857), .A(n5550), .B(n5549), .ZN(U2865)
         );
  AOI22_X1 U6687 ( .A1(n6610), .A2(DATAI_25_), .B1(n6608), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U6688 ( .A1(n6609), .A2(DATAI_9_), .ZN(n5551) );
  OAI211_X1 U6689 ( .C1(n5553), .C2(n5857), .A(n5552), .B(n5551), .ZN(U2866)
         );
  AOI22_X1 U6690 ( .A1(n6609), .A2(DATAI_8_), .B1(n6608), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5555) );
  NAND2_X1 U6691 ( .A1(n6610), .A2(DATAI_24_), .ZN(n5554) );
  OAI211_X1 U6692 ( .C1(n5815), .C2(n5857), .A(n5555), .B(n5554), .ZN(U2867)
         );
  AOI22_X1 U6693 ( .A1(n5557), .A2(DATAI_15_), .B1(n6608), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5556) );
  OAI21_X1 U6694 ( .B1(n5634), .B2(n5857), .A(n5556), .ZN(U2876) );
  AOI22_X1 U6695 ( .A1(n5557), .A2(DATAI_14_), .B1(n6608), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5558) );
  OAI21_X1 U6696 ( .B1(n5559), .B2(n5857), .A(n5558), .ZN(U2877) );
  INV_X1 U6697 ( .A(n5560), .ZN(n5562) );
  NAND2_X1 U6698 ( .A1(n5562), .A2(n5561), .ZN(n5563) );
  XNOR2_X1 U6699 ( .A(n5563), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5652)
         );
  NOR2_X1 U6700 ( .A1(n6242), .A2(n5564), .ZN(n5646) );
  AOI21_X1 U6701 ( .B1(n6196), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5646), 
        .ZN(n5565) );
  OAI21_X1 U6702 ( .B1(n5566), .B2(n6188), .A(n5565), .ZN(n5567) );
  AOI21_X1 U6703 ( .B1(n5568), .B2(n6183), .A(n5567), .ZN(n5569) );
  OAI21_X1 U6704 ( .B1(n5652), .B2(n6190), .A(n5569), .ZN(U2957) );
  NAND3_X1 U6705 ( .A1(n5576), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(n5890), .ZN(n5570) );
  OR3_X1 U6706 ( .A1(n5874), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .A3(n5585), 
        .ZN(n5577) );
  AOI22_X1 U6707 ( .A1(n5570), .A2(n5577), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5668), .ZN(n5571) );
  XNOR2_X1 U6708 ( .A(n5571), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5658)
         );
  NAND2_X1 U6709 ( .A1(n6218), .A2(REIP_REG_28__SCAN_IN), .ZN(n5654) );
  OAI21_X1 U6710 ( .B1(n6174), .B2(n5572), .A(n5654), .ZN(n5574) );
  NOR2_X1 U6711 ( .A1(n5789), .A2(n6199), .ZN(n5573) );
  AOI211_X1 U6712 ( .C1(n6168), .C2(n5785), .A(n5574), .B(n5573), .ZN(n5575)
         );
  OAI21_X1 U6713 ( .B1(n5658), .B2(n6190), .A(n5575), .ZN(U2958) );
  NAND2_X1 U6714 ( .A1(n5576), .A2(n5587), .ZN(n5578) );
  NAND2_X1 U6715 ( .A1(n5578), .A2(n5577), .ZN(n5579) );
  XNOR2_X1 U6716 ( .A(n5579), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5665)
         );
  NAND2_X1 U6717 ( .A1(n6218), .A2(REIP_REG_27__SCAN_IN), .ZN(n5660) );
  OAI21_X1 U6718 ( .B1(n6174), .B2(n5580), .A(n5660), .ZN(n5582) );
  NOR2_X1 U6719 ( .A1(n5799), .A2(n6199), .ZN(n5581) );
  AOI211_X1 U6720 ( .C1(n6168), .C2(n5583), .A(n5582), .B(n5581), .ZN(n5584)
         );
  OAI21_X1 U6721 ( .B1(n5665), .B2(n6190), .A(n5584), .ZN(U2959) );
  INV_X1 U6722 ( .A(n5585), .ZN(n5586) );
  NOR2_X1 U6723 ( .A1(n5587), .A2(n5586), .ZN(n5588) );
  XNOR2_X1 U6724 ( .A(n5589), .B(n5588), .ZN(n5676) );
  NAND2_X1 U6725 ( .A1(n6218), .A2(REIP_REG_26__SCAN_IN), .ZN(n5672) );
  OAI21_X1 U6726 ( .B1(n6174), .B2(n5590), .A(n5672), .ZN(n5592) );
  NOR2_X1 U6727 ( .A1(n5806), .A2(n6199), .ZN(n5591) );
  AOI211_X1 U6728 ( .C1(n6168), .C2(n5803), .A(n5592), .B(n5591), .ZN(n5593)
         );
  OAI21_X1 U6729 ( .B1(n5676), .B2(n6190), .A(n5593), .ZN(U2960) );
  AOI21_X1 U6730 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5890), .A(n5595), 
        .ZN(n5596) );
  XNOR2_X1 U6731 ( .A(n5594), .B(n5596), .ZN(n5684) );
  INV_X1 U6732 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5597) );
  NAND2_X1 U6733 ( .A1(n6218), .A2(REIP_REG_22__SCAN_IN), .ZN(n5678) );
  OAI21_X1 U6734 ( .B1(n6174), .B2(n5597), .A(n5678), .ZN(n5600) );
  NOR2_X1 U6735 ( .A1(n5598), .A2(n6199), .ZN(n5599) );
  AOI211_X1 U6736 ( .C1(n6168), .C2(n5601), .A(n5600), .B(n5599), .ZN(n5602)
         );
  OAI21_X1 U6737 ( .B1(n5684), .B2(n6190), .A(n5602), .ZN(U2964) );
  OAI21_X1 U6738 ( .B1(n5605), .B2(n5604), .A(n5603), .ZN(n5695) );
  NAND2_X1 U6739 ( .A1(n6218), .A2(REIP_REG_20__SCAN_IN), .ZN(n5685) );
  OAI21_X1 U6740 ( .B1(n6174), .B2(n5606), .A(n5685), .ZN(n5609) );
  NOR2_X1 U6741 ( .A1(n5607), .A2(n6199), .ZN(n5608) );
  AOI211_X1 U6742 ( .C1(n6168), .C2(n5610), .A(n5609), .B(n5608), .ZN(n5611)
         );
  OAI21_X1 U6743 ( .B1(n5695), .B2(n6190), .A(n5611), .ZN(U2966) );
  INV_X1 U6744 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5889) );
  NOR2_X1 U6745 ( .A1(n5624), .A2(n5889), .ZN(n5892) );
  NOR2_X1 U6746 ( .A1(n3500), .A2(n5913), .ZN(n5616) );
  NOR3_X1 U6747 ( .A1(n5614), .A2(n5890), .A3(n5629), .ZN(n5891) );
  NOR2_X1 U6748 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5615) );
  AOI22_X1 U6749 ( .A1(n5892), .A2(n5616), .B1(n5891), .B2(n5615), .ZN(n5618)
         );
  XNOR2_X1 U6750 ( .A(n5618), .B(n5617), .ZN(n5717) );
  NOR2_X1 U6751 ( .A1(n6242), .A2(n6540), .ZN(n5714) );
  AOI21_X1 U6752 ( .B1(n6196), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5714), 
        .ZN(n5619) );
  OAI21_X1 U6753 ( .B1(n5620), .B2(n6188), .A(n5619), .ZN(n5621) );
  AOI21_X1 U6754 ( .B1(n6096), .B2(n6183), .A(n5621), .ZN(n5622) );
  OAI21_X1 U6755 ( .B1(n5717), .B2(n6190), .A(n5622), .ZN(U2968) );
  XNOR2_X1 U6756 ( .A(n5890), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5623)
         );
  XNOR2_X1 U6757 ( .A(n5624), .B(n5623), .ZN(n5718) );
  NAND2_X1 U6758 ( .A1(n5718), .A2(n6182), .ZN(n5628) );
  NOR2_X1 U6759 ( .A1(n6242), .A2(n5414), .ZN(n5723) );
  NOR2_X1 U6760 ( .A1(n6188), .A2(n5625), .ZN(n5626) );
  AOI211_X1 U6761 ( .C1(n6196), .C2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5723), 
        .B(n5626), .ZN(n5627) );
  OAI211_X1 U6762 ( .C1(n6199), .C2(n6099), .A(n5628), .B(n5627), .ZN(U2970)
         );
  XNOR2_X1 U6763 ( .A(n5614), .B(n5629), .ZN(n5922) );
  NAND2_X1 U6764 ( .A1(n5922), .A2(n6182), .ZN(n5633) );
  NAND2_X1 U6765 ( .A1(n6218), .A2(REIP_REG_15__SCAN_IN), .ZN(n5918) );
  OAI21_X1 U6766 ( .B1(n6174), .B2(n6771), .A(n5918), .ZN(n5630) );
  AOI21_X1 U6767 ( .B1(n6168), .B2(n5631), .A(n5630), .ZN(n5632) );
  OAI211_X1 U6768 ( .C1(n6199), .C2(n5634), .A(n5633), .B(n5632), .ZN(U2971)
         );
  CLKBUF_X1 U6769 ( .A(n5636), .Z(n5637) );
  OAI21_X1 U6770 ( .B1(n5635), .B2(n5638), .A(n5637), .ZN(n5933) );
  AOI22_X1 U6771 ( .A1(n6196), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .B1(n6218), 
        .B2(REIP_REG_13__SCAN_IN), .ZN(n5640) );
  NAND2_X1 U6772 ( .A1(n6168), .A2(n5984), .ZN(n5639) );
  OAI211_X1 U6773 ( .C1(n6086), .C2(n6199), .A(n5640), .B(n5639), .ZN(n5641)
         );
  AOI21_X1 U6774 ( .B1(n5933), .B2(n6182), .A(n5641), .ZN(n5642) );
  INV_X1 U6775 ( .A(n5642), .ZN(U2973) );
  INV_X1 U6776 ( .A(n5643), .ZN(n5647) );
  NOR3_X1 U6777 ( .A1(n5659), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5644), 
        .ZN(n5645) );
  AOI211_X1 U6778 ( .C1(n5647), .C2(n6240), .A(n5646), .B(n5645), .ZN(n5651)
         );
  OR2_X1 U6779 ( .A1(n5649), .A2(n5648), .ZN(n5650) );
  OAI211_X1 U6780 ( .C1(n5652), .C2(n6203), .A(n5651), .B(n5650), .ZN(U2989)
         );
  XNOR2_X1 U6781 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .B(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5653) );
  NOR2_X1 U6782 ( .A1(n5659), .A2(n5653), .ZN(n5656) );
  OAI21_X1 U6783 ( .B1(n5788), .B2(n6229), .A(n5654), .ZN(n5655) );
  AOI211_X1 U6784 ( .C1(n5663), .C2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5656), .B(n5655), .ZN(n5657) );
  OAI21_X1 U6785 ( .B1(n5658), .B2(n6203), .A(n5657), .ZN(U2990) );
  NOR2_X1 U6786 ( .A1(n5659), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5662)
         );
  OAI21_X1 U6787 ( .B1(n5798), .B2(n6229), .A(n5660), .ZN(n5661) );
  AOI211_X1 U6788 ( .C1(n5663), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5662), .B(n5661), .ZN(n5664) );
  OAI21_X1 U6789 ( .B1(n5665), .B2(n6203), .A(n5664), .ZN(U2991) );
  INV_X1 U6790 ( .A(n5906), .ZN(n5674) );
  INV_X1 U6791 ( .A(n5666), .ZN(n5670) );
  INV_X1 U6792 ( .A(n5900), .ZN(n5667) );
  AOI21_X1 U6793 ( .B1(n5668), .B2(n6744), .A(n5667), .ZN(n5669) );
  NAND2_X1 U6794 ( .A1(n5670), .A2(n5669), .ZN(n5671) );
  OAI211_X1 U6795 ( .C1(n5805), .C2(n6229), .A(n5672), .B(n5671), .ZN(n5673)
         );
  AOI21_X1 U6796 ( .B1(n5674), .B2(INSTADDRPOINTER_REG_26__SCAN_IN), .A(n5673), 
        .ZN(n5675) );
  OAI21_X1 U6797 ( .B1(n5676), .B2(n6203), .A(n5675), .ZN(U2992) );
  NAND2_X1 U6798 ( .A1(n5677), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5679) );
  OAI211_X1 U6799 ( .C1(n6229), .C2(n5680), .A(n5679), .B(n5678), .ZN(n5681)
         );
  AOI21_X1 U6800 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5682), .A(n5681), 
        .ZN(n5683) );
  OAI21_X1 U6801 ( .B1(n5684), .B2(n6203), .A(n5683), .ZN(U2996) );
  INV_X1 U6802 ( .A(n5685), .ZN(n5690) );
  INV_X1 U6803 ( .A(n5686), .ZN(n5706) );
  NOR3_X1 U6804 ( .A1(n5688), .A2(n5687), .A3(n5706), .ZN(n5689) );
  AOI211_X1 U6805 ( .C1(n5691), .C2(n6240), .A(n5690), .B(n5689), .ZN(n5694)
         );
  INV_X1 U6806 ( .A(n5704), .ZN(n5692) );
  NAND2_X1 U6807 ( .A1(n5692), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5693) );
  OAI211_X1 U6808 ( .C1(n5695), .C2(n6203), .A(n5694), .B(n5693), .ZN(U2998)
         );
  AOI21_X1 U6809 ( .B1(n5698), .B2(n5697), .A(n5696), .ZN(n5883) );
  INV_X1 U6810 ( .A(n5699), .ZN(n5700) );
  OR2_X1 U6811 ( .A1(n5391), .A2(n5700), .ZN(n5703) );
  INV_X1 U6812 ( .A(n5701), .ZN(n5702) );
  XNOR2_X1 U6813 ( .A(n5703), .B(n5702), .ZN(n5854) );
  NAND2_X1 U6814 ( .A1(n6218), .A2(REIP_REG_19__SCAN_IN), .ZN(n5886) );
  OAI221_X1 U6815 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5706), .C1(
        n5705), .C2(n5704), .A(n5886), .ZN(n5707) );
  AOI21_X1 U6816 ( .B1(n6240), .B2(n5854), .A(n5707), .ZN(n5708) );
  OAI21_X1 U6817 ( .B1(n5883), .B2(n6203), .A(n5708), .ZN(U2999) );
  AOI21_X1 U6818 ( .B1(n5710), .B2(n5709), .A(n5912), .ZN(n5711) );
  AOI21_X1 U6819 ( .B1(n5617), .B2(n5712), .A(n5711), .ZN(n5713) );
  AOI211_X1 U6820 ( .C1(n6240), .C2(n5715), .A(n5714), .B(n5713), .ZN(n5716)
         );
  OAI21_X1 U6821 ( .B1(n5717), .B2(n6203), .A(n5716), .ZN(U3000) );
  INV_X1 U6822 ( .A(n5718), .ZN(n5729) );
  OAI21_X1 U6823 ( .B1(n5720), .B2(n5719), .A(n6210), .ZN(n5917) );
  NOR3_X1 U6824 ( .A1(n6201), .A2(n5722), .A3(n5721), .ZN(n5921) );
  AOI22_X1 U6825 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .B1(n5889), .B2(n3491), .ZN(n5724)
         );
  AOI21_X1 U6826 ( .B1(n5921), .B2(n5724), .A(n5723), .ZN(n5725) );
  OAI21_X1 U6827 ( .B1(n5726), .B2(n6229), .A(n5725), .ZN(n5727) );
  AOI21_X1 U6828 ( .B1(n5917), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5727), 
        .ZN(n5728) );
  OAI21_X1 U6829 ( .B1(n5729), .B2(n6203), .A(n5728), .ZN(U3002) );
  OAI211_X1 U6830 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5744), .A(n6369), .B(
        n6343), .ZN(n5730) );
  OAI21_X1 U6831 ( .B1(n5741), .B2(n5731), .A(n5730), .ZN(n5732) );
  MUX2_X1 U6832 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5732), .S(n6254), 
        .Z(U3464) );
  XNOR2_X1 U6833 ( .A(n5733), .B(n6369), .ZN(n5735) );
  OAI22_X1 U6834 ( .A1(n5735), .A2(n6382), .B1(n5734), .B2(n5741), .ZN(n5736)
         );
  MUX2_X1 U6835 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5736), .S(n6254), 
        .Z(U3463) );
  NOR2_X1 U6836 ( .A1(n5737), .A2(n6369), .ZN(n6348) );
  NOR2_X1 U6837 ( .A1(n5738), .A2(n6348), .ZN(n5739) );
  OAI222_X1 U6838 ( .A1(n5742), .A2(n6297), .B1(n5741), .B2(n5740), .C1(n6382), 
        .C2(n5739), .ZN(n5743) );
  MUX2_X1 U6839 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5743), .S(n6254), 
        .Z(U3462) );
  AND2_X1 U6840 ( .A1(n5744), .A2(n3032), .ZN(n5745) );
  NAND2_X1 U6841 ( .A1(n5780), .A2(n6343), .ZN(n5746) );
  OAI21_X1 U6842 ( .B1(n5746), .B2(n5782), .A(n6297), .ZN(n5752) );
  AND2_X1 U6843 ( .A1(n5748), .A2(n5747), .ZN(n5751) );
  NOR3_X1 U6844 ( .A1(n6299), .A2(n6458), .A3(n5749), .ZN(n5750) );
  AOI21_X1 U6845 ( .B1(n5752), .B2(n5751), .A(n5750), .ZN(n5784) );
  NOR3_X1 U6846 ( .A1(n6458), .A2(n6445), .A3(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), 
        .ZN(n6379) );
  NAND2_X1 U6847 ( .A1(n6256), .A2(n6379), .ZN(n5753) );
  INV_X1 U6848 ( .A(n5753), .ZN(n5778) );
  INV_X1 U6849 ( .A(n5751), .ZN(n6374) );
  AOI22_X1 U6850 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5753), .B1(n5752), .B2(
        n6374), .ZN(n5754) );
  AOI22_X1 U6851 ( .A1(n6376), .A2(n5778), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5777), .ZN(n5756) );
  OAI21_X1 U6852 ( .B1(n5780), .B2(n6305), .A(n5756), .ZN(n5757) );
  AOI21_X1 U6853 ( .B1(n6386), .B2(n5782), .A(n5757), .ZN(n5758) );
  OAI21_X1 U6854 ( .B1(n5784), .B2(n6389), .A(n5758), .ZN(U3100) );
  AOI22_X1 U6855 ( .A1(n6390), .A2(n5778), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5777), .ZN(n5759) );
  OAI21_X1 U6856 ( .B1(n5780), .B2(n6309), .A(n5759), .ZN(n5760) );
  AOI21_X1 U6857 ( .B1(n5782), .B2(n6392), .A(n5760), .ZN(n5761) );
  OAI21_X1 U6858 ( .B1(n5784), .B2(n6395), .A(n5761), .ZN(U3101) );
  AOI22_X1 U6859 ( .A1(n6396), .A2(n5778), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5777), .ZN(n5762) );
  OAI21_X1 U6860 ( .B1(n5780), .B2(n6313), .A(n5762), .ZN(n5763) );
  AOI21_X1 U6861 ( .B1(n5782), .B2(n6397), .A(n5763), .ZN(n5764) );
  OAI21_X1 U6862 ( .B1(n5784), .B2(n6401), .A(n5764), .ZN(U3102) );
  AOI22_X1 U6863 ( .A1(n6402), .A2(n5778), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5777), .ZN(n5765) );
  OAI21_X1 U6864 ( .B1(n5780), .B2(n6317), .A(n5765), .ZN(n5766) );
  AOI21_X1 U6865 ( .B1(n5782), .B2(n6403), .A(n5766), .ZN(n5767) );
  OAI21_X1 U6866 ( .B1(n5784), .B2(n6407), .A(n5767), .ZN(U3103) );
  AOI22_X1 U6867 ( .A1(n6408), .A2(n5778), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5777), .ZN(n5768) );
  OAI21_X1 U6868 ( .B1(n5780), .B2(n6321), .A(n5768), .ZN(n5769) );
  AOI21_X1 U6869 ( .B1(n5782), .B2(n6409), .A(n5769), .ZN(n5770) );
  OAI21_X1 U6870 ( .B1(n5784), .B2(n6413), .A(n5770), .ZN(U3104) );
  AOI22_X1 U6871 ( .A1(n6414), .A2(n5778), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5777), .ZN(n5771) );
  OAI21_X1 U6872 ( .B1(n5780), .B2(n6325), .A(n5771), .ZN(n5772) );
  AOI21_X1 U6873 ( .B1(n5782), .B2(n6416), .A(n5772), .ZN(n5773) );
  OAI21_X1 U6874 ( .B1(n5784), .B2(n6419), .A(n5773), .ZN(U3105) );
  AOI22_X1 U6875 ( .A1(n6420), .A2(n5778), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5777), .ZN(n5774) );
  OAI21_X1 U6876 ( .B1(n5780), .B2(n6329), .A(n5774), .ZN(n5775) );
  AOI21_X1 U6877 ( .B1(n5782), .B2(n6421), .A(n5775), .ZN(n5776) );
  OAI21_X1 U6878 ( .B1(n5784), .B2(n6425), .A(n5776), .ZN(U3106) );
  AOI22_X1 U6879 ( .A1(n6427), .A2(n5778), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5777), .ZN(n5779) );
  OAI21_X1 U6880 ( .B1(n5780), .B2(n6337), .A(n5779), .ZN(n5781) );
  AOI21_X1 U6881 ( .B1(n5782), .B2(n6431), .A(n5781), .ZN(n5783) );
  OAI21_X1 U6882 ( .B1(n5784), .B2(n6435), .A(n5783), .ZN(U3107) );
  AND2_X1 U6883 ( .A1(n6120), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  NAND2_X1 U6884 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5797), .ZN(n5793) );
  INV_X1 U6885 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6555) );
  AOI22_X1 U6886 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n6034), .B1(n5785), 
        .B2(n6053), .ZN(n5786) );
  OAI21_X1 U6887 ( .B1(n5787), .B2(n6555), .A(n5786), .ZN(n5791) );
  OAI22_X1 U6888 ( .A1(n5789), .A2(n6039), .B1(n5788), .B2(n6048), .ZN(n5790)
         );
  AOI211_X1 U6889 ( .C1(EBX_REG_28__SCAN_IN), .C2(n6051), .A(n5791), .B(n5790), 
        .ZN(n5792) );
  OAI21_X1 U6890 ( .B1(REIP_REG_28__SCAN_IN), .B2(n5793), .A(n5792), .ZN(U2799) );
  INV_X1 U6891 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6552) );
  AOI22_X1 U6892 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6051), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6034), .ZN(n5794) );
  OAI21_X1 U6893 ( .B1(n5795), .B2(n6070), .A(n5794), .ZN(n5796) );
  AOI221_X1 U6894 ( .B1(n5797), .B2(n6552), .C1(n5809), .C2(
        REIP_REG_27__SCAN_IN), .A(n5796), .ZN(n5802) );
  OAI22_X1 U6895 ( .A1(n5799), .A2(n6039), .B1(n5798), .B2(n6048), .ZN(n5800)
         );
  INV_X1 U6896 ( .A(n5800), .ZN(n5801) );
  NAND2_X1 U6897 ( .A1(n5802), .A2(n5801), .ZN(U2800) );
  AOI22_X1 U6898 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6034), .B1(n5803), 
        .B2(n6053), .ZN(n5811) );
  NAND2_X1 U6899 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_25__SCAN_IN), .ZN(
        n5804) );
  INV_X1 U6900 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6550) );
  OAI21_X1 U6901 ( .B1(n5819), .B2(n5804), .A(n6550), .ZN(n5808) );
  OAI22_X1 U6902 ( .A1(n5806), .A2(n6039), .B1(n5805), .B2(n6048), .ZN(n5807)
         );
  AOI21_X1 U6903 ( .B1(n5809), .B2(n5808), .A(n5807), .ZN(n5810) );
  OAI211_X1 U6904 ( .C1(n6738), .C2(n6078), .A(n5811), .B(n5810), .ZN(U2801)
         );
  AOI22_X1 U6905 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n6034), .B1(n5812), 
        .B2(n6053), .ZN(n5813) );
  OAI21_X1 U6906 ( .B1(n5827), .B2(n6783), .A(n5813), .ZN(n5817) );
  OAI22_X1 U6907 ( .A1(n5815), .A2(n6039), .B1(n5814), .B2(n6048), .ZN(n5816)
         );
  AOI211_X1 U6908 ( .C1(EBX_REG_24__SCAN_IN), .C2(n6051), .A(n5817), .B(n5816), 
        .ZN(n5818) );
  OAI21_X1 U6909 ( .B1(REIP_REG_24__SCAN_IN), .B2(n5819), .A(n5818), .ZN(U2803) );
  NOR2_X1 U6910 ( .A1(REIP_REG_23__SCAN_IN), .A2(n5820), .ZN(n5826) );
  INV_X1 U6911 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n6638) );
  OAI22_X1 U6912 ( .A1(n6638), .A2(n6069), .B1(n5821), .B2(n6070), .ZN(n5822)
         );
  AOI21_X1 U6913 ( .B1(EBX_REG_23__SCAN_IN), .B2(n6051), .A(n5822), .ZN(n5825)
         );
  INV_X1 U6914 ( .A(n5823), .ZN(n5858) );
  AOI22_X1 U6915 ( .A1(n5858), .A2(n6012), .B1(n5848), .B2(n6064), .ZN(n5824)
         );
  OAI211_X1 U6916 ( .C1(n5827), .C2(n5826), .A(n5825), .B(n5824), .ZN(U2804)
         );
  INV_X1 U6917 ( .A(n5828), .ZN(n5832) );
  INV_X1 U6918 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6545) );
  INV_X1 U6919 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5853) );
  OAI22_X1 U6920 ( .A1(n5853), .A2(n6078), .B1(n5829), .B2(n6069), .ZN(n5830)
         );
  AOI221_X1 U6921 ( .B1(n5832), .B2(n6545), .C1(n5831), .C2(
        REIP_REG_21__SCAN_IN), .A(n5830), .ZN(n5835) );
  NOR2_X1 U6922 ( .A1(n5850), .A2(n6048), .ZN(n5833) );
  AOI21_X1 U6923 ( .B1(n5864), .B2(n6012), .A(n5833), .ZN(n5834) );
  OAI211_X1 U6924 ( .C1(n5836), .C2(n6070), .A(n5835), .B(n5834), .ZN(U2806)
         );
  INV_X1 U6925 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5888) );
  OAI21_X1 U6926 ( .B1(n6069), .B2(n5888), .A(n6066), .ZN(n5841) );
  OAI21_X1 U6927 ( .B1(REIP_REG_19__SCAN_IN), .B2(REIP_REG_18__SCAN_IN), .A(
        n5837), .ZN(n5838) );
  OAI22_X1 U6928 ( .A1(n5973), .A2(n6542), .B1(n5839), .B2(n5838), .ZN(n5840)
         );
  AOI211_X1 U6929 ( .C1(EBX_REG_19__SCAN_IN), .C2(n6051), .A(n5841), .B(n5840), 
        .ZN(n5847) );
  AND2_X1 U6930 ( .A1(n5843), .A2(n5842), .ZN(n5845) );
  AOI22_X1 U6931 ( .A1(n5870), .A2(n6012), .B1(n6064), .B2(n5854), .ZN(n5846)
         );
  OAI211_X1 U6932 ( .C1(n5884), .C2(n6070), .A(n5847), .B(n5846), .ZN(U2808)
         );
  INV_X1 U6933 ( .A(EBX_REG_23__SCAN_IN), .ZN(n6642) );
  AOI22_X1 U6934 ( .A1(n5858), .A2(n6092), .B1(n5848), .B2(n6081), .ZN(n5849)
         );
  OAI21_X1 U6935 ( .B1(n6642), .B2(n6094), .A(n5849), .ZN(U2836) );
  NOR2_X1 U6936 ( .A1(n5850), .A2(n6090), .ZN(n5851) );
  AOI21_X1 U6937 ( .B1(n5864), .B2(n6092), .A(n5851), .ZN(n5852) );
  OAI21_X1 U6938 ( .B1(n5853), .B2(n6094), .A(n5852), .ZN(U2838) );
  AOI22_X1 U6939 ( .A1(n5870), .A2(n6092), .B1(n6081), .B2(n5854), .ZN(n5855)
         );
  OAI21_X1 U6940 ( .B1(n5856), .B2(n6094), .A(n5855), .ZN(U2840) );
  INV_X1 U6941 ( .A(n5857), .ZN(n6611) );
  AOI22_X1 U6942 ( .A1(n5858), .A2(n6611), .B1(n6610), .B2(DATAI_23_), .ZN(
        n5860) );
  AOI22_X1 U6943 ( .A1(n6609), .A2(DATAI_7_), .B1(n6608), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5859) );
  NAND2_X1 U6944 ( .A1(n5860), .A2(n5859), .ZN(U2868) );
  AOI22_X1 U6945 ( .A1(n5861), .A2(n6611), .B1(n6610), .B2(DATAI_22_), .ZN(
        n5863) );
  AOI22_X1 U6946 ( .A1(n6609), .A2(DATAI_6_), .B1(n6608), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U6947 ( .A1(n5863), .A2(n5862), .ZN(U2869) );
  AOI22_X1 U6948 ( .A1(n5864), .A2(n6611), .B1(n6610), .B2(DATAI_21_), .ZN(
        n5866) );
  AOI22_X1 U6949 ( .A1(n6609), .A2(DATAI_5_), .B1(n6608), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U6950 ( .A1(n5866), .A2(n5865), .ZN(U2870) );
  AOI22_X1 U6951 ( .A1(n5867), .A2(n6611), .B1(n6610), .B2(DATAI_20_), .ZN(
        n5869) );
  AOI22_X1 U6952 ( .A1(n6609), .A2(DATAI_4_), .B1(n6608), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5868) );
  NAND2_X1 U6953 ( .A1(n5869), .A2(n5868), .ZN(U2871) );
  AOI22_X1 U6954 ( .A1(n5870), .A2(n6611), .B1(n6610), .B2(DATAI_19_), .ZN(
        n5872) );
  AOI22_X1 U6955 ( .A1(n6609), .A2(DATAI_3_), .B1(n6608), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U6956 ( .A1(n5872), .A2(n5871), .ZN(U2872) );
  AOI22_X1 U6957 ( .A1(n6218), .A2(REIP_REG_25__SCAN_IN), .B1(n6196), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5880) );
  INV_X1 U6958 ( .A(n5873), .ZN(n5877) );
  INV_X1 U6959 ( .A(n5874), .ZN(n5876) );
  OAI21_X1 U6960 ( .B1(n5877), .B2(n5876), .A(n5875), .ZN(n5903) );
  AOI22_X1 U6961 ( .A1(n5903), .A2(n6182), .B1(n6183), .B2(n5878), .ZN(n5879)
         );
  OAI211_X1 U6962 ( .C1(n6188), .C2(n5881), .A(n5880), .B(n5879), .ZN(U2961)
         );
  OAI222_X1 U6963 ( .A1(n6188), .A2(n5884), .B1(n6190), .B2(n5883), .C1(n6199), 
        .C2(n5882), .ZN(n5885) );
  INV_X1 U6964 ( .A(n5885), .ZN(n5887) );
  OAI211_X1 U6965 ( .C1(n5888), .C2(n6174), .A(n5887), .B(n5886), .ZN(U2967)
         );
  AOI22_X1 U6966 ( .A1(n6218), .A2(REIP_REG_17__SCAN_IN), .B1(n6196), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5899) );
  OAI22_X1 U6967 ( .A1(n5892), .A2(n5891), .B1(n5890), .B2(n5889), .ZN(n5893)
         );
  XNOR2_X1 U6968 ( .A(n5893), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5910)
         );
  OR2_X1 U6969 ( .A1(n5895), .A2(n5894), .ZN(n5896) );
  AOI22_X1 U6970 ( .A1(n5910), .A2(n6182), .B1(n6183), .B2(n6612), .ZN(n5898)
         );
  OAI211_X1 U6971 ( .C1(n6188), .C2(n5977), .A(n5899), .B(n5898), .ZN(U2969)
         );
  AOI22_X1 U6972 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6218), .B1(n5900), .B2(
        n6744), .ZN(n5905) );
  INV_X1 U6973 ( .A(n5901), .ZN(n5902) );
  AOI22_X1 U6974 ( .A1(n5903), .A2(n6247), .B1(n6240), .B2(n5902), .ZN(n5904)
         );
  OAI211_X1 U6975 ( .C1(n5906), .C2(n6744), .A(n5905), .B(n5904), .ZN(U2993)
         );
  OR2_X1 U6976 ( .A1(n5908), .A2(n5907), .ZN(n5909) );
  AND2_X1 U6977 ( .A1(n5391), .A2(n5909), .ZN(n6080) );
  AOI22_X1 U6978 ( .A1(n5910), .A2(n6247), .B1(n6240), .B2(n6080), .ZN(n5916)
         );
  NOR2_X1 U6979 ( .A1(n6242), .A2(n6538), .ZN(n5911) );
  AOI221_X1 U6980 ( .B1(n5914), .B2(n5913), .C1(n5912), .C2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5911), .ZN(n5915) );
  NAND2_X1 U6981 ( .A1(n5916), .A2(n5915), .ZN(U3001) );
  INV_X1 U6982 ( .A(n5917), .ZN(n5925) );
  INV_X1 U6983 ( .A(n5918), .ZN(n5919) );
  AOI21_X1 U6984 ( .B1(n5920), .B2(n6240), .A(n5919), .ZN(n5924) );
  AOI22_X1 U6985 ( .A1(n5922), .A2(n6247), .B1(n5921), .B2(n3491), .ZN(n5923)
         );
  OAI211_X1 U6986 ( .C1(n5925), .C2(n3491), .A(n5924), .B(n5923), .ZN(U3003)
         );
  NAND2_X1 U6987 ( .A1(n5927), .A2(n5926), .ZN(n5928) );
  NAND2_X1 U6988 ( .A1(n5929), .A2(n5928), .ZN(n6084) );
  OAI22_X1 U6989 ( .A1(n5931), .A2(n5930), .B1(n6229), .B2(n6084), .ZN(n5932)
         );
  AOI21_X1 U6990 ( .B1(n5933), .B2(n6247), .A(n5932), .ZN(n5940) );
  NAND2_X1 U6991 ( .A1(n6218), .A2(REIP_REG_13__SCAN_IN), .ZN(n5938) );
  NAND3_X1 U6992 ( .A1(n5936), .A2(n5935), .A3(n5934), .ZN(n5937) );
  NAND4_X1 U6993 ( .A1(n5940), .A2(n5939), .A3(n5938), .A4(n5937), .ZN(U3005)
         );
  INV_X1 U6994 ( .A(n5941), .ZN(n6581) );
  NAND4_X1 U6995 ( .A1(n6061), .A2(n5944), .A3(n5943), .A4(n5942), .ZN(n5945)
         );
  OAI21_X1 U6996 ( .B1(n6581), .B2(n5946), .A(n5945), .ZN(U3455) );
  AOI21_X1 U6997 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6767), .A(n6508), .ZN(n5952) );
  INV_X1 U6998 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5947) );
  AND2_X1 U6999 ( .A1(n6508), .A2(STATE_REG_1__SCAN_IN), .ZN(n6607) );
  AOI21_X1 U7000 ( .B1(n5952), .B2(n5947), .A(n6607), .ZN(U2789) );
  OAI21_X1 U7001 ( .B1(n5948), .B2(n6482), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5949) );
  OAI21_X1 U7002 ( .B1(n5950), .B2(n6780), .A(n5949), .ZN(U2790) );
  INV_X2 U7003 ( .A(n6607), .ZN(n6605) );
  NOR2_X1 U7004 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5953) );
  OAI21_X1 U7005 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5953), .A(n6605), .ZN(n5951)
         );
  OAI21_X1 U7006 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6605), .A(n5951), .ZN(
        U2791) );
  NOR2_X1 U7007 ( .A1(n6607), .A2(n5952), .ZN(n6565) );
  OAI21_X1 U7008 ( .B1(n5953), .B2(BS16_N), .A(n6565), .ZN(n6564) );
  OAI21_X1 U7009 ( .B1(n6565), .B2(n6487), .A(n6564), .ZN(U2792) );
  OAI21_X1 U7010 ( .B1(n5955), .B2(n5954), .A(n6190), .ZN(U2793) );
  NOR4_X1 U7011 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n5959) );
  NOR4_X1 U7012 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n5958) );
  NOR4_X1 U7013 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5957) );
  NOR4_X1 U7014 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_24__SCAN_IN), .A4(
        DATAWIDTH_REG_25__SCAN_IN), .ZN(n5956) );
  NAND4_X1 U7015 ( .A1(n5959), .A2(n5958), .A3(n5957), .A4(n5956), .ZN(n5965)
         );
  NOR4_X1 U7016 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(DATAWIDTH_REG_2__SCAN_IN), .A3(DATAWIDTH_REG_3__SCAN_IN), .A4(DATAWIDTH_REG_4__SCAN_IN), .ZN(n5963) );
  AOI211_X1 U7017 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_13__SCAN_IN), .B(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5962) );
  NOR4_X1 U7018 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n5961)
         );
  NOR4_X1 U7019 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(DATAWIDTH_REG_6__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n5960) );
  NAND4_X1 U7020 ( .A1(n5963), .A2(n5962), .A3(n5961), .A4(n5960), .ZN(n5964)
         );
  NOR2_X1 U7021 ( .A1(n5965), .A2(n5964), .ZN(n6590) );
  INV_X1 U7022 ( .A(n6590), .ZN(n5968) );
  NAND2_X1 U7023 ( .A1(n6590), .A2(n6586), .ZN(n6587) );
  NOR3_X1 U7024 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(n6587), .ZN(n5967) );
  AOI21_X1 U7025 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(n5968), .A(n5967), .ZN(
        n5966) );
  OAI21_X1 U7026 ( .B1(n5490), .B2(n5968), .A(n5966), .ZN(U2794) );
  NAND2_X1 U7027 ( .A1(n6590), .A2(n5490), .ZN(n6591) );
  AOI21_X1 U7028 ( .B1(BYTEENABLE_REG_3__SCAN_IN), .B2(n5968), .A(n5967), .ZN(
        n5969) );
  OAI21_X1 U7029 ( .B1(DATAWIDTH_REG_1__SCAN_IN), .B2(n6591), .A(n5969), .ZN(
        U2795) );
  NOR2_X1 U7030 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5970), .ZN(n5972) );
  INV_X1 U7031 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5971) );
  OAI22_X1 U7032 ( .A1(n5973), .A2(n5972), .B1(n5971), .B2(n6069), .ZN(n5974)
         );
  AOI211_X1 U7033 ( .C1(n6051), .C2(EBX_REG_17__SCAN_IN), .A(n6050), .B(n5974), 
        .ZN(n5976) );
  AOI22_X1 U7034 ( .A1(n6612), .A2(n6012), .B1(n6064), .B2(n6080), .ZN(n5975)
         );
  OAI211_X1 U7035 ( .C1(n5977), .C2(n6070), .A(n5976), .B(n5975), .ZN(U2810)
         );
  INV_X1 U7036 ( .A(n6084), .ZN(n5978) );
  AOI22_X1 U7037 ( .A1(n5978), .A2(n6064), .B1(REIP_REG_13__SCAN_IN), .B2(
        n5991), .ZN(n5989) );
  OAI21_X1 U7038 ( .B1(REIP_REG_13__SCAN_IN), .B2(REIP_REG_12__SCAN_IN), .A(
        n5979), .ZN(n5980) );
  OAI22_X1 U7039 ( .A1(n5982), .A2(n6069), .B1(n5981), .B2(n5980), .ZN(n5983)
         );
  AOI211_X1 U7040 ( .C1(n6051), .C2(EBX_REG_13__SCAN_IN), .A(n6050), .B(n5983), 
        .ZN(n5988) );
  INV_X1 U7041 ( .A(n5984), .ZN(n5985) );
  OAI22_X1 U7042 ( .A1(n6086), .A2(n6039), .B1(n6070), .B2(n5985), .ZN(n5986)
         );
  INV_X1 U7043 ( .A(n5986), .ZN(n5987) );
  NAND3_X1 U7044 ( .A1(n5989), .A2(n5988), .A3(n5987), .ZN(U2814) );
  AOI21_X1 U7045 ( .B1(REIP_REG_10__SCAN_IN), .B2(n5990), .A(
        REIP_REG_11__SCAN_IN), .ZN(n6003) );
  INV_X1 U7046 ( .A(n5991), .ZN(n6002) );
  AND2_X1 U7047 ( .A1(n5993), .A2(n5992), .ZN(n5995) );
  OR2_X1 U7048 ( .A1(n5995), .A2(n5994), .ZN(n6202) );
  INV_X1 U7049 ( .A(n6202), .ZN(n5999) );
  INV_X1 U7050 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6095) );
  NOR2_X1 U7051 ( .A1(n6078), .A2(n6095), .ZN(n5998) );
  OAI21_X1 U7052 ( .B1(n6069), .B2(n5996), .A(n6066), .ZN(n5997) );
  AOI211_X1 U7053 ( .C1(n5999), .C2(n6064), .A(n5998), .B(n5997), .ZN(n6001)
         );
  AOI22_X1 U7054 ( .A1(n6158), .A2(n6012), .B1(n6053), .B2(n6157), .ZN(n6000)
         );
  OAI211_X1 U7055 ( .C1(n6003), .C2(n6002), .A(n6001), .B(n6000), .ZN(U2816)
         );
  INV_X1 U7056 ( .A(n6228), .ZN(n6004) );
  AOI22_X1 U7057 ( .A1(n6004), .A2(n6064), .B1(n6051), .B2(EBX_REG_9__SCAN_IN), 
        .ZN(n6005) );
  OAI211_X1 U7058 ( .C1(n6069), .C2(n6006), .A(n6005), .B(n6066), .ZN(n6007)
         );
  AOI211_X1 U7059 ( .C1(n6009), .C2(REIP_REG_9__SCAN_IN), .A(n6008), .B(n6007), 
        .ZN(n6015) );
  INV_X1 U7060 ( .A(n6010), .ZN(n6013) );
  AOI22_X1 U7061 ( .A1(n6013), .A2(n6012), .B1(n6053), .B2(n6011), .ZN(n6014)
         );
  NAND2_X1 U7062 ( .A1(n6015), .A2(n6014), .ZN(U2818) );
  OAI21_X1 U7063 ( .B1(REIP_REG_7__SCAN_IN), .B2(REIP_REG_6__SCAN_IN), .A(
        n6016), .ZN(n6023) );
  NAND2_X1 U7064 ( .A1(n6034), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6017)
         );
  NAND2_X1 U7065 ( .A1(n6017), .A2(n6066), .ZN(n6018) );
  AOI21_X1 U7066 ( .B1(n6051), .B2(EBX_REG_7__SCAN_IN), .A(n6018), .ZN(n6022)
         );
  INV_X1 U7067 ( .A(n6019), .ZN(n6020) );
  NAND2_X1 U7068 ( .A1(n6064), .A2(n6020), .ZN(n6021) );
  OAI211_X1 U7069 ( .C1(n6044), .C2(n6023), .A(n6022), .B(n6021), .ZN(n6030)
         );
  INV_X1 U7070 ( .A(n6024), .ZN(n6025) );
  NAND2_X1 U7071 ( .A1(n6026), .A2(n6025), .ZN(n6027) );
  NAND2_X1 U7072 ( .A1(n6028), .A2(n6027), .ZN(n6057) );
  INV_X1 U7073 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6522) );
  NOR2_X1 U7074 ( .A1(n6057), .A2(n6522), .ZN(n6029) );
  NOR2_X1 U7075 ( .A1(n6030), .A2(n6029), .ZN(n6031) );
  OAI21_X1 U7076 ( .B1(n6162), .B2(n6039), .A(n6031), .ZN(n6032) );
  INV_X1 U7077 ( .A(n6032), .ZN(n6033) );
  OAI21_X1 U7078 ( .B1(n6161), .B2(n6070), .A(n6033), .ZN(U2820) );
  AOI21_X1 U7079 ( .B1(n6034), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n6050), 
        .ZN(n6036) );
  NAND2_X1 U7080 ( .A1(n6051), .A2(EBX_REG_6__SCAN_IN), .ZN(n6035) );
  OAI211_X1 U7081 ( .C1(n6048), .C2(n6037), .A(n6036), .B(n6035), .ZN(n6042)
         );
  OAI22_X1 U7082 ( .A1(n6040), .A2(n6039), .B1(n6038), .B2(n6070), .ZN(n6041)
         );
  NOR2_X1 U7083 ( .A1(n6042), .A2(n6041), .ZN(n6043) );
  OAI221_X1 U7084 ( .B1(REIP_REG_6__SCAN_IN), .B2(n6044), .C1(n6521), .C2(
        n6057), .A(n6043), .ZN(U2821) );
  NOR2_X1 U7085 ( .A1(n6046), .A2(n6045), .ZN(n6060) );
  AOI21_X1 U7086 ( .B1(REIP_REG_4__SCAN_IN), .B2(n6060), .A(
        REIP_REG_5__SCAN_IN), .ZN(n6058) );
  OAI22_X1 U7087 ( .A1(n6048), .A2(n6047), .B1(n6175), .B2(n6069), .ZN(n6049)
         );
  AOI211_X1 U7088 ( .C1(n6051), .C2(EBX_REG_5__SCAN_IN), .A(n6050), .B(n6049), 
        .ZN(n6056) );
  INV_X1 U7089 ( .A(n6052), .ZN(n6169) );
  AOI22_X1 U7090 ( .A1(n6170), .A2(n6054), .B1(n6169), .B2(n6053), .ZN(n6055)
         );
  OAI211_X1 U7091 ( .C1(n6058), .C2(n6057), .A(n6056), .B(n6055), .ZN(U2822)
         );
  INV_X1 U7092 ( .A(n6059), .ZN(n6062) );
  INV_X1 U7093 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6518) );
  AOI22_X1 U7094 ( .A1(n6062), .A2(n6061), .B1(n6060), .B2(n6518), .ZN(n6077)
         );
  AOI22_X1 U7095 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6065), .B1(n6064), .B2(n6063), .ZN(n6067) );
  OAI211_X1 U7096 ( .C1(n6069), .C2(n6068), .A(n6067), .B(n6066), .ZN(n6075)
         );
  OAI22_X1 U7097 ( .A1(n6073), .A2(n6072), .B1(n6071), .B2(n6070), .ZN(n6074)
         );
  NOR2_X1 U7098 ( .A1(n6075), .A2(n6074), .ZN(n6076) );
  OAI211_X1 U7099 ( .C1(n6079), .C2(n6078), .A(n6077), .B(n6076), .ZN(U2823)
         );
  AOI22_X1 U7100 ( .A1(n6612), .A2(n6092), .B1(n6081), .B2(n6080), .ZN(n6082)
         );
  OAI21_X1 U7101 ( .B1(n6083), .B2(n6094), .A(n6082), .ZN(U2842) );
  INV_X1 U7102 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6089) );
  OAI22_X1 U7103 ( .A1(n6086), .A2(n6085), .B1(n6090), .B2(n6084), .ZN(n6087)
         );
  INV_X1 U7104 ( .A(n6087), .ZN(n6088) );
  OAI21_X1 U7105 ( .B1(n6089), .B2(n6094), .A(n6088), .ZN(U2846) );
  NOR2_X1 U7106 ( .A1(n6202), .A2(n6090), .ZN(n6091) );
  AOI21_X1 U7107 ( .B1(n6158), .B2(n6092), .A(n6091), .ZN(n6093) );
  OAI21_X1 U7108 ( .B1(n6095), .B2(n6094), .A(n6093), .ZN(U2848) );
  AOI22_X1 U7109 ( .A1(n6096), .A2(n6611), .B1(n6610), .B2(DATAI_18_), .ZN(
        n6098) );
  AOI22_X1 U7110 ( .A1(n6609), .A2(DATAI_2_), .B1(n6608), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7111 ( .A1(n6098), .A2(n6097), .ZN(U2873) );
  INV_X1 U7112 ( .A(n6099), .ZN(n6100) );
  AOI22_X1 U7113 ( .A1(n6100), .A2(n6611), .B1(n6610), .B2(DATAI_16_), .ZN(
        n6102) );
  AOI22_X1 U7114 ( .A1(n6609), .A2(DATAI_0_), .B1(n6608), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6101) );
  NAND2_X1 U7115 ( .A1(n6102), .A2(n6101), .ZN(U2875) );
  INV_X1 U7116 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n6754) );
  AOI22_X1 U7117 ( .A1(EAX_REG_15__SCAN_IN), .A2(n6103), .B1(n6131), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6104) );
  OAI21_X1 U7118 ( .B1(n6754), .B2(n6105), .A(n6104), .ZN(U2908) );
  INV_X1 U7119 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6107) );
  AOI22_X1 U7120 ( .A1(n6597), .A2(LWORD_REG_14__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6106) );
  OAI21_X1 U7121 ( .B1(n6107), .B2(n6133), .A(n6106), .ZN(U2909) );
  INV_X1 U7122 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6109) );
  AOI22_X1 U7123 ( .A1(DATAO_REG_13__SCAN_IN), .A2(n6131), .B1(n6597), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6108) );
  OAI21_X1 U7124 ( .B1(n6109), .B2(n6133), .A(n6108), .ZN(U2910) );
  AOI22_X1 U7125 ( .A1(n6597), .A2(LWORD_REG_12__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6110) );
  OAI21_X1 U7126 ( .B1(n5012), .B2(n6133), .A(n6110), .ZN(U2911) );
  INV_X1 U7127 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6112) );
  AOI22_X1 U7128 ( .A1(n6597), .A2(LWORD_REG_11__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6111) );
  OAI21_X1 U7129 ( .B1(n6112), .B2(n6133), .A(n6111), .ZN(U2912) );
  INV_X1 U7130 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6114) );
  AOI22_X1 U7131 ( .A1(n6597), .A2(LWORD_REG_10__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6113) );
  OAI21_X1 U7132 ( .B1(n6114), .B2(n6133), .A(n6113), .ZN(U2913) );
  AOI22_X1 U7133 ( .A1(n6597), .A2(LWORD_REG_9__SCAN_IN), .B1(n6120), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6115) );
  OAI21_X1 U7134 ( .B1(n6789), .B2(n6133), .A(n6115), .ZN(U2914) );
  AOI22_X1 U7135 ( .A1(n6597), .A2(LWORD_REG_8__SCAN_IN), .B1(n6120), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6116) );
  OAI21_X1 U7136 ( .B1(n6117), .B2(n6133), .A(n6116), .ZN(U2915) );
  INV_X1 U7137 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6119) );
  AOI22_X1 U7138 ( .A1(n6597), .A2(LWORD_REG_7__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6118) );
  OAI21_X1 U7139 ( .B1(n6119), .B2(n6133), .A(n6118), .ZN(U2916) );
  AOI22_X1 U7140 ( .A1(n6597), .A2(LWORD_REG_6__SCAN_IN), .B1(n6120), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6121) );
  OAI21_X1 U7141 ( .B1(n6122), .B2(n6133), .A(n6121), .ZN(U2917) );
  INV_X1 U7142 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6124) );
  AOI22_X1 U7143 ( .A1(n6597), .A2(LWORD_REG_5__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6123) );
  OAI21_X1 U7144 ( .B1(n6124), .B2(n6133), .A(n6123), .ZN(U2918) );
  AOI22_X1 U7145 ( .A1(n6597), .A2(LWORD_REG_4__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6125) );
  OAI21_X1 U7146 ( .B1(n6759), .B2(n6133), .A(n6125), .ZN(U2919) );
  AOI22_X1 U7147 ( .A1(n6597), .A2(LWORD_REG_3__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6126) );
  OAI21_X1 U7148 ( .B1(n6127), .B2(n6133), .A(n6126), .ZN(U2920) );
  AOI22_X1 U7149 ( .A1(n6597), .A2(LWORD_REG_2__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6128) );
  OAI21_X1 U7150 ( .B1(n6773), .B2(n6133), .A(n6128), .ZN(U2921) );
  AOI22_X1 U7151 ( .A1(DATAO_REG_1__SCAN_IN), .A2(n6131), .B1(n6597), .B2(
        LWORD_REG_1__SCAN_IN), .ZN(n6129) );
  OAI21_X1 U7152 ( .B1(n6130), .B2(n6133), .A(n6129), .ZN(U2922) );
  AOI22_X1 U7153 ( .A1(n6597), .A2(LWORD_REG_0__SCAN_IN), .B1(n6131), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6132) );
  OAI21_X1 U7154 ( .B1(n6134), .B2(n6133), .A(n6132), .ZN(U2923) );
  AOI22_X1 U7155 ( .A1(EAX_REG_26__SCAN_IN), .A2(n6148), .B1(n6145), .B2(
        UWORD_REG_10__SCAN_IN), .ZN(n6135) );
  NAND2_X1 U7156 ( .A1(n6149), .A2(DATAI_10_), .ZN(n6139) );
  NAND2_X1 U7157 ( .A1(n6135), .A2(n6139), .ZN(U2934) );
  AOI22_X1 U7158 ( .A1(EAX_REG_28__SCAN_IN), .A2(n6148), .B1(n6145), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7159 ( .A1(n6149), .A2(DATAI_12_), .ZN(n6141) );
  NAND2_X1 U7160 ( .A1(n6136), .A2(n6141), .ZN(U2936) );
  AOI22_X1 U7161 ( .A1(EAX_REG_29__SCAN_IN), .A2(n6148), .B1(n6145), .B2(
        UWORD_REG_13__SCAN_IN), .ZN(n6137) );
  NAND2_X1 U7162 ( .A1(n6149), .A2(DATAI_13_), .ZN(n6143) );
  NAND2_X1 U7163 ( .A1(n6137), .A2(n6143), .ZN(U2937) );
  AOI22_X1 U7164 ( .A1(EAX_REG_30__SCAN_IN), .A2(n6148), .B1(n6145), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7165 ( .A1(n6149), .A2(DATAI_14_), .ZN(n6146) );
  NAND2_X1 U7166 ( .A1(n6138), .A2(n6146), .ZN(U2938) );
  AOI22_X1 U7167 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6148), .B1(n6145), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7168 ( .A1(n6140), .A2(n6139), .ZN(U2949) );
  AOI22_X1 U7169 ( .A1(EAX_REG_12__SCAN_IN), .A2(n6148), .B1(n6145), .B2(
        LWORD_REG_12__SCAN_IN), .ZN(n6142) );
  NAND2_X1 U7170 ( .A1(n6142), .A2(n6141), .ZN(U2951) );
  AOI22_X1 U7171 ( .A1(EAX_REG_13__SCAN_IN), .A2(n6148), .B1(n6145), .B2(
        LWORD_REG_13__SCAN_IN), .ZN(n6144) );
  NAND2_X1 U7172 ( .A1(n6144), .A2(n6143), .ZN(U2952) );
  AOI22_X1 U7173 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6148), .B1(n6145), .B2(
        LWORD_REG_14__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U7174 ( .A1(n6147), .A2(n6146), .ZN(U2953) );
  AOI22_X1 U7175 ( .A1(n6149), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6148), .ZN(n6150) );
  OAI21_X1 U7176 ( .B1(n6754), .B2(n6151), .A(n6150), .ZN(U2954) );
  INV_X1 U7177 ( .A(n6153), .ZN(n6155) );
  NAND2_X1 U7178 ( .A1(n6155), .A2(n6154), .ZN(n6156) );
  XNOR2_X1 U7179 ( .A(n6152), .B(n6156), .ZN(n6204) );
  AOI22_X1 U7180 ( .A1(n6218), .A2(REIP_REG_11__SCAN_IN), .B1(n6196), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6160) );
  AOI22_X1 U7181 ( .A1(n6158), .A2(n6183), .B1(n6168), .B2(n6157), .ZN(n6159)
         );
  OAI211_X1 U7182 ( .C1(n6204), .C2(n6190), .A(n6160), .B(n6159), .ZN(U2975)
         );
  OAI22_X1 U7183 ( .A1(n6162), .A2(n6199), .B1(n6161), .B2(n6188), .ZN(n6163)
         );
  AOI21_X1 U7184 ( .B1(n6164), .B2(n6182), .A(n6163), .ZN(n6166) );
  OAI211_X1 U7185 ( .C1(n6167), .C2(n6174), .A(n6166), .B(n6165), .ZN(U2979)
         );
  AOI222_X1 U7186 ( .A1(n6171), .A2(n6182), .B1(n6183), .B2(n6170), .C1(n6169), 
        .C2(n6168), .ZN(n6173) );
  OAI211_X1 U7187 ( .C1(n6175), .C2(n6174), .A(n6173), .B(n6172), .ZN(U2981)
         );
  AOI22_X1 U7188 ( .A1(n6218), .A2(REIP_REG_2__SCAN_IN), .B1(n6196), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6186) );
  INV_X1 U7189 ( .A(n6176), .ZN(n6179) );
  OR2_X1 U7190 ( .A1(n6179), .A2(n6178), .ZN(n6180) );
  XNOR2_X1 U7191 ( .A(n6181), .B(n6180), .ZN(n6248) );
  AOI22_X1 U7192 ( .A1(n6184), .A2(n6183), .B1(n6182), .B2(n6248), .ZN(n6185)
         );
  OAI211_X1 U7193 ( .C1(n6188), .C2(n6187), .A(n6186), .B(n6185), .ZN(U2984)
         );
  INV_X1 U7194 ( .A(n6189), .ZN(n6191) );
  AOI21_X1 U7195 ( .B1(n6191), .B2(n6577), .A(n6190), .ZN(n6194) );
  AOI21_X1 U7196 ( .B1(n6194), .B2(n6193), .A(n6192), .ZN(n6198) );
  OAI21_X1 U7197 ( .B1(n6196), .B2(n6195), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6197) );
  OAI211_X1 U7198 ( .C1(n6200), .C2(n6199), .A(n6198), .B(n6197), .ZN(U2986)
         );
  INV_X1 U7199 ( .A(n6201), .ZN(n6207) );
  OAI22_X1 U7200 ( .A1(n6202), .A2(n6229), .B1(n6529), .B2(n6242), .ZN(n6206)
         );
  NOR2_X1 U7201 ( .A1(n6204), .A2(n6203), .ZN(n6205) );
  AOI211_X1 U7202 ( .C1(n6209), .C2(n6207), .A(n6206), .B(n6205), .ZN(n6208)
         );
  OAI21_X1 U7203 ( .B1(n6210), .B2(n6209), .A(n6208), .ZN(U3007) );
  AOI21_X1 U7204 ( .B1(n6213), .B2(n6212), .A(n6211), .ZN(n6235) );
  INV_X1 U7205 ( .A(n6214), .ZN(n6222) );
  NAND2_X1 U7206 ( .A1(n6216), .A2(n6215), .ZN(n6226) );
  AOI221_X1 U7207 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n6234), .C2(n6224), .A(n6226), 
        .ZN(n6217) );
  AOI21_X1 U7208 ( .B1(n6218), .B2(REIP_REG_10__SCAN_IN), .A(n6217), .ZN(n6219) );
  OAI21_X1 U7209 ( .B1(n6220), .B2(n6229), .A(n6219), .ZN(n6221) );
  AOI21_X1 U7210 ( .B1(n6222), .B2(n6247), .A(n6221), .ZN(n6223) );
  OAI21_X1 U7211 ( .B1(n6235), .B2(n6224), .A(n6223), .ZN(U3008) );
  INV_X1 U7212 ( .A(n6225), .ZN(n6232) );
  NOR2_X1 U7213 ( .A1(n6226), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6231)
         );
  OAI21_X1 U7214 ( .B1(n6229), .B2(n6228), .A(n6227), .ZN(n6230) );
  AOI211_X1 U7215 ( .C1(n6232), .C2(n6247), .A(n6231), .B(n6230), .ZN(n6233)
         );
  OAI21_X1 U7216 ( .B1(n6235), .B2(n6234), .A(n6233), .ZN(U3009) );
  AOI221_X1 U7217 ( .B1(n6577), .B2(n6238), .C1(n6237), .C2(n6238), .A(n6236), 
        .ZN(n6244) );
  NAND2_X1 U7218 ( .A1(n6240), .A2(n6239), .ZN(n6241) );
  OAI21_X1 U7219 ( .B1(n5489), .B2(n6242), .A(n6241), .ZN(n6243) );
  NOR2_X1 U7220 ( .A1(n6244), .A2(n6243), .ZN(n6252) );
  NOR3_X1 U7221 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n6246), .A3(n6245), 
        .ZN(n6250) );
  AND2_X1 U7222 ( .A1(n6248), .A2(n6247), .ZN(n6249) );
  NOR2_X1 U7223 ( .A1(n6250), .A2(n6249), .ZN(n6251) );
  OAI211_X1 U7224 ( .C1(n6253), .C2(n3410), .A(n6252), .B(n6251), .ZN(U3016)
         );
  NOR2_X1 U7225 ( .A1(n6456), .A2(n6254), .ZN(U3019) );
  INV_X1 U7226 ( .A(n6255), .ZN(n6262) );
  NOR2_X1 U7227 ( .A1(n6256), .A2(n6258), .ZN(n6281) );
  AOI21_X1 U7228 ( .B1(n6257), .B2(n6441), .A(n6281), .ZN(n6261) );
  INV_X1 U7229 ( .A(n6261), .ZN(n6259) );
  INV_X1 U7230 ( .A(n6258), .ZN(n6265) );
  AOI22_X1 U7231 ( .A1(n6262), .A2(n6259), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6265), .ZN(n6286) );
  OR2_X1 U7232 ( .A1(n6260), .A2(n3032), .ZN(n6294) );
  AOI22_X1 U7233 ( .A1(n6377), .A2(n6333), .B1(n6376), .B2(n6281), .ZN(n6268)
         );
  NAND2_X1 U7234 ( .A1(n6262), .A2(n6261), .ZN(n6264) );
  OAI211_X1 U7235 ( .C1(n6343), .C2(n6265), .A(n6264), .B(n6263), .ZN(n6283)
         );
  AOI22_X1 U7236 ( .A1(n6283), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n6386), 
        .B2(n6282), .ZN(n6267) );
  OAI211_X1 U7237 ( .C1(n6286), .C2(n6389), .A(n6268), .B(n6267), .ZN(U3060)
         );
  AOI22_X1 U7238 ( .A1(n6391), .A2(n6333), .B1(n6390), .B2(n6281), .ZN(n6270)
         );
  AOI22_X1 U7239 ( .A1(n6283), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n6392), 
        .B2(n6282), .ZN(n6269) );
  OAI211_X1 U7240 ( .C1(n6286), .C2(n6395), .A(n6270), .B(n6269), .ZN(U3061)
         );
  AOI22_X1 U7241 ( .A1(n6398), .A2(n6333), .B1(n6396), .B2(n6281), .ZN(n6272)
         );
  AOI22_X1 U7242 ( .A1(n6283), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n6397), 
        .B2(n6282), .ZN(n6271) );
  OAI211_X1 U7243 ( .C1(n6286), .C2(n6401), .A(n6272), .B(n6271), .ZN(U3062)
         );
  AOI22_X1 U7244 ( .A1(n6404), .A2(n6333), .B1(n6402), .B2(n6281), .ZN(n6274)
         );
  AOI22_X1 U7245 ( .A1(n6283), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n6403), 
        .B2(n6282), .ZN(n6273) );
  OAI211_X1 U7246 ( .C1(n6286), .C2(n6407), .A(n6274), .B(n6273), .ZN(U3063)
         );
  AOI22_X1 U7247 ( .A1(n6410), .A2(n6333), .B1(n6408), .B2(n6281), .ZN(n6276)
         );
  AOI22_X1 U7248 ( .A1(n6283), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n6409), 
        .B2(n6282), .ZN(n6275) );
  OAI211_X1 U7249 ( .C1(n6286), .C2(n6413), .A(n6276), .B(n6275), .ZN(U3064)
         );
  AOI22_X1 U7250 ( .A1(n6415), .A2(n6333), .B1(n6414), .B2(n6281), .ZN(n6278)
         );
  AOI22_X1 U7251 ( .A1(n6283), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n6416), 
        .B2(n6282), .ZN(n6277) );
  OAI211_X1 U7252 ( .C1(n6286), .C2(n6419), .A(n6278), .B(n6277), .ZN(U3065)
         );
  AOI22_X1 U7253 ( .A1(n6422), .A2(n6333), .B1(n6420), .B2(n6281), .ZN(n6280)
         );
  AOI22_X1 U7254 ( .A1(n6283), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n6421), 
        .B2(n6282), .ZN(n6279) );
  OAI211_X1 U7255 ( .C1(n6286), .C2(n6425), .A(n6280), .B(n6279), .ZN(U3066)
         );
  AOI22_X1 U7256 ( .A1(n6428), .A2(n6333), .B1(n6427), .B2(n6281), .ZN(n6285)
         );
  AOI22_X1 U7257 ( .A1(n6283), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n6431), 
        .B2(n6282), .ZN(n6284) );
  OAI211_X1 U7258 ( .C1(n6286), .C2(n6435), .A(n6285), .B(n6284), .ZN(U3067)
         );
  NAND3_X1 U7259 ( .A1(n6290), .A2(n6289), .A3(n6458), .ZN(n6291) );
  OAI21_X1 U7260 ( .B1(n6292), .B2(n6296), .A(n6291), .ZN(n6331) );
  INV_X1 U7261 ( .A(n6341), .ZN(n6345) );
  NOR2_X1 U7262 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6345), .ZN(n6330)
         );
  AOI22_X1 U7263 ( .A1(n6293), .A2(n6331), .B1(n6376), .B2(n6330), .ZN(n6304)
         );
  NAND3_X1 U7264 ( .A1(n6342), .A2(n6294), .A3(n6343), .ZN(n6298) );
  NOR2_X1 U7265 ( .A1(n6296), .A2(n6295), .ZN(n6339) );
  AOI21_X1 U7266 ( .B1(n6298), .B2(n6297), .A(n6339), .ZN(n6302) );
  OAI211_X1 U7267 ( .C1(n6330), .C2(n6569), .A(n6299), .B(n6458), .ZN(n6300)
         );
  AOI22_X1 U7268 ( .A1(n6334), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6386), 
        .B2(n6333), .ZN(n6303) );
  OAI211_X1 U7269 ( .C1(n6305), .C2(n6342), .A(n6304), .B(n6303), .ZN(U3068)
         );
  AOI22_X1 U7270 ( .A1(n6306), .A2(n6331), .B1(n6390), .B2(n6330), .ZN(n6308)
         );
  AOI22_X1 U7271 ( .A1(n6334), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6392), 
        .B2(n6333), .ZN(n6307) );
  OAI211_X1 U7272 ( .C1(n6309), .C2(n6342), .A(n6308), .B(n6307), .ZN(U3069)
         );
  AOI22_X1 U7273 ( .A1(n6310), .A2(n6331), .B1(n6396), .B2(n6330), .ZN(n6312)
         );
  AOI22_X1 U7274 ( .A1(n6334), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6397), 
        .B2(n6333), .ZN(n6311) );
  OAI211_X1 U7275 ( .C1(n6313), .C2(n6342), .A(n6312), .B(n6311), .ZN(U3070)
         );
  AOI22_X1 U7276 ( .A1(n6314), .A2(n6331), .B1(n6402), .B2(n6330), .ZN(n6316)
         );
  AOI22_X1 U7277 ( .A1(n6334), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6403), 
        .B2(n6333), .ZN(n6315) );
  OAI211_X1 U7278 ( .C1(n6317), .C2(n6342), .A(n6316), .B(n6315), .ZN(U3071)
         );
  AOI22_X1 U7279 ( .A1(n6318), .A2(n6331), .B1(n6408), .B2(n6330), .ZN(n6320)
         );
  AOI22_X1 U7280 ( .A1(n6334), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6409), 
        .B2(n6333), .ZN(n6319) );
  OAI211_X1 U7281 ( .C1(n6321), .C2(n6342), .A(n6320), .B(n6319), .ZN(U3072)
         );
  AOI22_X1 U7282 ( .A1(n6322), .A2(n6331), .B1(n6414), .B2(n6330), .ZN(n6324)
         );
  AOI22_X1 U7283 ( .A1(n6334), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6416), 
        .B2(n6333), .ZN(n6323) );
  OAI211_X1 U7284 ( .C1(n6325), .C2(n6342), .A(n6324), .B(n6323), .ZN(U3073)
         );
  AOI22_X1 U7285 ( .A1(n6326), .A2(n6331), .B1(n6420), .B2(n6330), .ZN(n6328)
         );
  AOI22_X1 U7286 ( .A1(n6334), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6421), 
        .B2(n6333), .ZN(n6327) );
  OAI211_X1 U7287 ( .C1(n6329), .C2(n6342), .A(n6328), .B(n6327), .ZN(U3074)
         );
  AOI22_X1 U7288 ( .A1(n6332), .A2(n6331), .B1(n6427), .B2(n6330), .ZN(n6336)
         );
  AOI22_X1 U7289 ( .A1(n6334), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6431), 
        .B2(n6333), .ZN(n6335) );
  OAI211_X1 U7290 ( .C1(n6337), .C2(n6342), .A(n6336), .B(n6335), .ZN(U3075)
         );
  INV_X1 U7291 ( .A(n6338), .ZN(n6363) );
  AOI21_X1 U7292 ( .B1(n6339), .B2(n6441), .A(n6363), .ZN(n6344) );
  NOR2_X1 U7293 ( .A1(n6344), .A2(n6382), .ZN(n6340) );
  AOI21_X1 U7294 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6341), .A(n6340), .ZN(
        n6368) );
  AOI22_X1 U7295 ( .A1(n6386), .A2(n6364), .B1(n6376), .B2(n6363), .ZN(n6350)
         );
  NAND2_X1 U7296 ( .A1(n6344), .A2(n6343), .ZN(n6347) );
  AOI21_X1 U7297 ( .B1(n6382), .B2(n6345), .A(n6380), .ZN(n6346) );
  OAI21_X1 U7298 ( .B1(n6348), .B2(n6347), .A(n6346), .ZN(n6365) );
  AOI22_X1 U7299 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6365), .B1(n6377), 
        .B2(n3047), .ZN(n6349) );
  OAI211_X1 U7300 ( .C1(n6368), .C2(n6389), .A(n6350), .B(n6349), .ZN(U3076)
         );
  AOI22_X1 U7301 ( .A1(n6392), .A2(n6364), .B1(n6390), .B2(n6363), .ZN(n6352)
         );
  AOI22_X1 U7302 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6365), .B1(n6391), 
        .B2(n3047), .ZN(n6351) );
  OAI211_X1 U7303 ( .C1(n6368), .C2(n6395), .A(n6352), .B(n6351), .ZN(U3077)
         );
  AOI22_X1 U7304 ( .A1(n6398), .A2(n3047), .B1(n6396), .B2(n6363), .ZN(n6354)
         );
  AOI22_X1 U7305 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6365), .B1(n6397), 
        .B2(n6364), .ZN(n6353) );
  OAI211_X1 U7306 ( .C1(n6368), .C2(n6401), .A(n6354), .B(n6353), .ZN(U3078)
         );
  AOI22_X1 U7307 ( .A1(n6403), .A2(n6364), .B1(n6402), .B2(n6363), .ZN(n6356)
         );
  AOI22_X1 U7308 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6365), .B1(n6404), 
        .B2(n3047), .ZN(n6355) );
  OAI211_X1 U7309 ( .C1(n6368), .C2(n6407), .A(n6356), .B(n6355), .ZN(U3079)
         );
  AOI22_X1 U7310 ( .A1(n6409), .A2(n6364), .B1(n6408), .B2(n6363), .ZN(n6358)
         );
  AOI22_X1 U7311 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6365), .B1(n6410), 
        .B2(n3047), .ZN(n6357) );
  OAI211_X1 U7312 ( .C1(n6368), .C2(n6413), .A(n6358), .B(n6357), .ZN(U3080)
         );
  AOI22_X1 U7313 ( .A1(n6415), .A2(n3047), .B1(n6414), .B2(n6363), .ZN(n6360)
         );
  AOI22_X1 U7314 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6365), .B1(n6416), 
        .B2(n6364), .ZN(n6359) );
  OAI211_X1 U7315 ( .C1(n6368), .C2(n6419), .A(n6360), .B(n6359), .ZN(U3081)
         );
  AOI22_X1 U7316 ( .A1(n6421), .A2(n6364), .B1(n6420), .B2(n6363), .ZN(n6362)
         );
  AOI22_X1 U7317 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6365), .B1(n6422), 
        .B2(n3047), .ZN(n6361) );
  OAI211_X1 U7318 ( .C1(n6368), .C2(n6425), .A(n6362), .B(n6361), .ZN(U3082)
         );
  AOI22_X1 U7319 ( .A1(n6428), .A2(n3047), .B1(n6427), .B2(n6363), .ZN(n6367)
         );
  AOI22_X1 U7320 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6365), .B1(n6431), 
        .B2(n6364), .ZN(n6366) );
  OAI211_X1 U7321 ( .C1(n6368), .C2(n6435), .A(n6367), .B(n6366), .ZN(U3083)
         );
  INV_X1 U7322 ( .A(n6369), .ZN(n6370) );
  AOI21_X1 U7323 ( .B1(n6371), .B2(n6370), .A(n6382), .ZN(n6378) );
  NAND2_X1 U7324 ( .A1(n6372), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6375) );
  OAI21_X1 U7325 ( .B1(n6374), .B2(n6373), .A(n6375), .ZN(n6384) );
  AOI22_X1 U7326 ( .A1(n6378), .A2(n6384), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n6379), .ZN(n6436) );
  INV_X1 U7327 ( .A(n6375), .ZN(n6426) );
  AOI22_X1 U7328 ( .A1(n6429), .A2(n6377), .B1(n6376), .B2(n6426), .ZN(n6388)
         );
  INV_X1 U7329 ( .A(n6378), .ZN(n6385) );
  INV_X1 U7330 ( .A(n6379), .ZN(n6381) );
  AOI21_X1 U7331 ( .B1(n6382), .B2(n6381), .A(n6380), .ZN(n6383) );
  OAI21_X1 U7332 ( .B1(n6385), .B2(n6384), .A(n6383), .ZN(n6432) );
  AOI22_X1 U7333 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6432), .B1(n6386), 
        .B2(n6430), .ZN(n6387) );
  OAI211_X1 U7334 ( .C1(n6436), .C2(n6389), .A(n6388), .B(n6387), .ZN(U3108)
         );
  AOI22_X1 U7335 ( .A1(n6429), .A2(n6391), .B1(n6390), .B2(n6426), .ZN(n6394)
         );
  AOI22_X1 U7336 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6432), .B1(n6392), 
        .B2(n6430), .ZN(n6393) );
  OAI211_X1 U7337 ( .C1(n6436), .C2(n6395), .A(n6394), .B(n6393), .ZN(U3109)
         );
  AOI22_X1 U7338 ( .A1(n6430), .A2(n6397), .B1(n6396), .B2(n6426), .ZN(n6400)
         );
  AOI22_X1 U7339 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6432), .B1(n6398), 
        .B2(n6429), .ZN(n6399) );
  OAI211_X1 U7340 ( .C1(n6436), .C2(n6401), .A(n6400), .B(n6399), .ZN(U3110)
         );
  AOI22_X1 U7341 ( .A1(n6430), .A2(n6403), .B1(n6402), .B2(n6426), .ZN(n6406)
         );
  AOI22_X1 U7342 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6432), .B1(n6404), 
        .B2(n6429), .ZN(n6405) );
  OAI211_X1 U7343 ( .C1(n6436), .C2(n6407), .A(n6406), .B(n6405), .ZN(U3111)
         );
  AOI22_X1 U7344 ( .A1(n6430), .A2(n6409), .B1(n6408), .B2(n6426), .ZN(n6412)
         );
  AOI22_X1 U7345 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6432), .B1(n6410), 
        .B2(n6429), .ZN(n6411) );
  OAI211_X1 U7346 ( .C1(n6436), .C2(n6413), .A(n6412), .B(n6411), .ZN(U3112)
         );
  AOI22_X1 U7347 ( .A1(n6429), .A2(n6415), .B1(n6414), .B2(n6426), .ZN(n6418)
         );
  AOI22_X1 U7348 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6432), .B1(n6416), 
        .B2(n6430), .ZN(n6417) );
  OAI211_X1 U7349 ( .C1(n6436), .C2(n6419), .A(n6418), .B(n6417), .ZN(U3113)
         );
  AOI22_X1 U7350 ( .A1(n6430), .A2(n6421), .B1(n6420), .B2(n6426), .ZN(n6424)
         );
  AOI22_X1 U7351 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6432), .B1(n6422), 
        .B2(n6429), .ZN(n6423) );
  OAI211_X1 U7352 ( .C1(n6436), .C2(n6425), .A(n6424), .B(n6423), .ZN(U3114)
         );
  AOI22_X1 U7353 ( .A1(n6429), .A2(n6428), .B1(n6427), .B2(n6426), .ZN(n6434)
         );
  AOI22_X1 U7354 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6432), .B1(n6431), 
        .B2(n6430), .ZN(n6433) );
  OAI211_X1 U7355 ( .C1(n6436), .C2(n6435), .A(n6434), .B(n6433), .ZN(U3115)
         );
  NAND2_X1 U7356 ( .A1(n6459), .A2(n6458), .ZN(n6455) );
  INV_X1 U7357 ( .A(n6437), .ZN(n6439) );
  AOI22_X1 U7358 ( .A1(n6441), .A2(n6440), .B1(n6439), .B2(n6438), .ZN(n6579)
         );
  NAND2_X1 U7359 ( .A1(n6442), .A2(n3507), .ZN(n6584) );
  NAND3_X1 U7360 ( .A1(n6579), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6584), .ZN(n6444) );
  OAI21_X1 U7361 ( .B1(n6445), .B2(n6444), .A(n6443), .ZN(n6447) );
  NAND2_X1 U7362 ( .A1(n6445), .A2(n6444), .ZN(n6446) );
  OAI21_X1 U7363 ( .B1(n6448), .B2(n6447), .A(n6446), .ZN(n6453) );
  NAND2_X1 U7364 ( .A1(n6452), .A2(n6453), .ZN(n6449) );
  NAND2_X1 U7365 ( .A1(n6450), .A2(n6449), .ZN(n6451) );
  OAI21_X1 U7366 ( .B1(n6453), .B2(n6452), .A(n6451), .ZN(n6454) );
  NAND2_X1 U7367 ( .A1(n6455), .A2(n6454), .ZN(n6457) );
  OAI211_X1 U7368 ( .C1(n6459), .C2(n6458), .A(n6457), .B(n6456), .ZN(n6470)
         );
  NOR2_X1 U7369 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6464) );
  OR2_X1 U7370 ( .A1(n6461), .A2(n6460), .ZN(n6462) );
  OAI211_X1 U7371 ( .C1(n6465), .C2(n6464), .A(n6463), .B(n6462), .ZN(n6466)
         );
  NOR2_X1 U7372 ( .A1(n6467), .A2(n6466), .ZN(n6468) );
  AND3_X1 U7373 ( .A1(n6470), .A2(n6469), .A3(n6468), .ZN(n6483) );
  NAND2_X1 U7374 ( .A1(n6483), .A2(n6484), .ZN(n6472) );
  NAND2_X1 U7375 ( .A1(READY_N), .A2(n6597), .ZN(n6471) );
  NAND2_X1 U7376 ( .A1(n6472), .A2(n6471), .ZN(n6477) );
  INV_X1 U7377 ( .A(n6473), .ZN(n6474) );
  NAND2_X1 U7378 ( .A1(n6475), .A2(n6474), .ZN(n6476) );
  OAI21_X1 U7379 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6596), .A(n6568), .ZN(
        n6489) );
  AOI221_X1 U7380 ( .B1(n6479), .B2(STATE2_REG_0__SCAN_IN), .C1(n6489), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6478), .ZN(n6481) );
  OAI211_X1 U7381 ( .C1(n6493), .C2(n6571), .A(n6780), .B(n6568), .ZN(n6480)
         );
  OAI211_X1 U7382 ( .C1(n6483), .C2(n6482), .A(n6481), .B(n6480), .ZN(U3148)
         );
  AOI21_X1 U7383 ( .B1(n6485), .B2(n6596), .A(n6484), .ZN(n6491) );
  NAND2_X1 U7384 ( .A1(n6780), .A2(n6486), .ZN(n6488) );
  INV_X1 U7385 ( .A(n6488), .ZN(n6496) );
  OAI221_X1 U7386 ( .B1(n6496), .B2(n6489), .C1(n6488), .C2(n6487), .A(
        STATE2_REG_1__SCAN_IN), .ZN(n6490) );
  OAI21_X1 U7387 ( .B1(n6492), .B2(n6491), .A(n6490), .ZN(U3149) );
  OAI211_X1 U7388 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6596), .A(n6566), .B(
        n6493), .ZN(n6495) );
  OAI21_X1 U7389 ( .B1(n6496), .B2(n6495), .A(n6494), .ZN(U3150) );
  INV_X1 U7390 ( .A(n6565), .ZN(n6497) );
  AND2_X1 U7391 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6497), .ZN(U3151) );
  AND2_X1 U7392 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6497), .ZN(U3152) );
  INV_X1 U7393 ( .A(DATAWIDTH_REG_29__SCAN_IN), .ZN(n6784) );
  NOR2_X1 U7394 ( .A1(n6565), .A2(n6784), .ZN(U3153) );
  AND2_X1 U7395 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6497), .ZN(U3154) );
  INV_X1 U7396 ( .A(DATAWIDTH_REG_27__SCAN_IN), .ZN(n6619) );
  NOR2_X1 U7397 ( .A1(n6565), .A2(n6619), .ZN(U3155) );
  AND2_X1 U7398 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6497), .ZN(U3156) );
  AND2_X1 U7399 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6497), .ZN(U3157) );
  AND2_X1 U7400 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6497), .ZN(U3158) );
  AND2_X1 U7401 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6497), .ZN(U3159) );
  AND2_X1 U7402 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6497), .ZN(U3160) );
  AND2_X1 U7403 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6497), .ZN(U3161) );
  AND2_X1 U7404 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6497), .ZN(U3162) );
  AND2_X1 U7405 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6497), .ZN(U3163) );
  AND2_X1 U7406 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6497), .ZN(U3164) );
  AND2_X1 U7407 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6497), .ZN(U3165) );
  AND2_X1 U7408 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6497), .ZN(U3166) );
  AND2_X1 U7409 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6497), .ZN(U3167) );
  AND2_X1 U7410 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6497), .ZN(U3168) );
  INV_X1 U7411 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6741) );
  NOR2_X1 U7412 ( .A1(n6565), .A2(n6741), .ZN(U3169) );
  AND2_X1 U7413 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6497), .ZN(U3170) );
  AND2_X1 U7414 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6497), .ZN(U3171) );
  AND2_X1 U7415 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6497), .ZN(U3172) );
  AND2_X1 U7416 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6497), .ZN(U3173) );
  AND2_X1 U7417 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6497), .ZN(U3174) );
  AND2_X1 U7418 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6497), .ZN(U3175) );
  AND2_X1 U7419 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6497), .ZN(U3176) );
  AND2_X1 U7420 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6497), .ZN(U3177) );
  AND2_X1 U7421 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6497), .ZN(U3178) );
  AND2_X1 U7422 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6497), .ZN(U3179) );
  AND2_X1 U7423 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6497), .ZN(U3180) );
  AOI22_X1 U7424 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6513) );
  AND2_X1 U7425 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6501) );
  INV_X1 U7426 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6499) );
  INV_X1 U7427 ( .A(NA_N), .ZN(n6506) );
  AOI221_X1 U7428 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6506), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6510) );
  AOI221_X1 U7429 ( .B1(n6501), .B2(n6605), .C1(n6499), .C2(n6605), .A(n6510), 
        .ZN(n6498) );
  OAI21_X1 U7430 ( .B1(n6505), .B2(n6513), .A(n6498), .ZN(U3181) );
  NOR2_X1 U7431 ( .A1(n6508), .A2(n6499), .ZN(n6507) );
  NAND2_X1 U7432 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6500) );
  OAI21_X1 U7433 ( .B1(n6507), .B2(n6501), .A(n6500), .ZN(n6502) );
  OAI211_X1 U7434 ( .C1(n6504), .C2(n6596), .A(n6503), .B(n6502), .ZN(U3182)
         );
  AOI21_X1 U7435 ( .B1(n6507), .B2(n6506), .A(n6505), .ZN(n6512) );
  AOI221_X1 U7436 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6596), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6509) );
  AOI221_X1 U7437 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6509), .C2(HOLD), .A(n6508), .ZN(n6511) );
  OAI22_X1 U7438 ( .A1(n6513), .A2(n6512), .B1(n6511), .B2(n6510), .ZN(U3183)
         );
  INV_X1 U7439 ( .A(n6556), .ZN(n6561) );
  NAND2_X1 U7440 ( .A1(n6767), .A2(n6607), .ZN(n6558) );
  INV_X1 U7441 ( .A(n6558), .ZN(n6559) );
  AOI22_X1 U7442 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6605), .ZN(n6514) );
  OAI21_X1 U7443 ( .B1(n5490), .B2(n6561), .A(n6514), .ZN(U3184) );
  AOI22_X1 U7444 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6605), .ZN(n6515) );
  OAI21_X1 U7445 ( .B1(n5489), .B2(n6561), .A(n6515), .ZN(U3185) );
  AOI22_X1 U7446 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6556), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6605), .ZN(n6516) );
  OAI21_X1 U7447 ( .B1(n6518), .B2(n6558), .A(n6516), .ZN(U3186) );
  AOI22_X1 U7448 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6605), .ZN(n6517) );
  OAI21_X1 U7449 ( .B1(n6518), .B2(n6561), .A(n6517), .ZN(U3187) );
  AOI22_X1 U7450 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6556), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6605), .ZN(n6519) );
  OAI21_X1 U7451 ( .B1(n6521), .B2(n6558), .A(n6519), .ZN(U3188) );
  AOI22_X1 U7452 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6605), .ZN(n6520) );
  OAI21_X1 U7453 ( .B1(n6521), .B2(n6561), .A(n6520), .ZN(U3189) );
  INV_X1 U7454 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6739) );
  OAI222_X1 U7455 ( .A1(n6561), .A2(n6522), .B1(n6739), .B2(n6607), .C1(n6524), 
        .C2(n6558), .ZN(U3190) );
  AOI22_X1 U7456 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6605), .ZN(n6523) );
  OAI21_X1 U7457 ( .B1(n6524), .B2(n6561), .A(n6523), .ZN(U3191) );
  AOI22_X1 U7458 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6556), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6605), .ZN(n6525) );
  OAI21_X1 U7459 ( .B1(n6527), .B2(n6558), .A(n6525), .ZN(U3192) );
  AOI22_X1 U7460 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6605), .ZN(n6526) );
  OAI21_X1 U7461 ( .B1(n6527), .B2(n6561), .A(n6526), .ZN(U3193) );
  AOI22_X1 U7462 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6605), .ZN(n6528) );
  OAI21_X1 U7463 ( .B1(n6529), .B2(n6561), .A(n6528), .ZN(U3194) );
  INV_X1 U7464 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6531) );
  AOI22_X1 U7465 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6605), .ZN(n6530) );
  OAI21_X1 U7466 ( .B1(n6531), .B2(n6561), .A(n6530), .ZN(U3195) );
  AOI22_X1 U7467 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6556), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6605), .ZN(n6532) );
  OAI21_X1 U7468 ( .B1(n6534), .B2(n6558), .A(n6532), .ZN(U3196) );
  AOI22_X1 U7469 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6605), .ZN(n6533) );
  OAI21_X1 U7470 ( .B1(n6534), .B2(n6561), .A(n6533), .ZN(U3197) );
  AOI222_X1 U7471 ( .A1(n6556), .A2(REIP_REG_15__SCAN_IN), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6605), .C1(REIP_REG_16__SCAN_IN), .C2(
        n6559), .ZN(n6535) );
  INV_X1 U7472 ( .A(n6535), .ZN(U3198) );
  AOI22_X1 U7473 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6556), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6605), .ZN(n6536) );
  OAI21_X1 U7474 ( .B1(n6538), .B2(n6558), .A(n6536), .ZN(U3199) );
  AOI22_X1 U7475 ( .A1(REIP_REG_18__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6605), .ZN(n6537) );
  OAI21_X1 U7476 ( .B1(n6538), .B2(n6561), .A(n6537), .ZN(U3200) );
  AOI22_X1 U7477 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6605), .ZN(n6539) );
  OAI21_X1 U7478 ( .B1(n6540), .B2(n6561), .A(n6539), .ZN(U3201) );
  AOI22_X1 U7479 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6605), .ZN(n6541) );
  OAI21_X1 U7480 ( .B1(n6542), .B2(n6561), .A(n6541), .ZN(U3202) );
  AOI22_X1 U7481 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6556), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6605), .ZN(n6543) );
  OAI21_X1 U7482 ( .B1(n6545), .B2(n6558), .A(n6543), .ZN(U3203) );
  AOI22_X1 U7483 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6605), .ZN(n6544) );
  OAI21_X1 U7484 ( .B1(n6545), .B2(n6561), .A(n6544), .ZN(U3204) );
  AOI222_X1 U7485 ( .A1(n6556), .A2(REIP_REG_22__SCAN_IN), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6605), .C1(REIP_REG_23__SCAN_IN), .C2(
        n6559), .ZN(n6546) );
  INV_X1 U7486 ( .A(n6546), .ZN(U3205) );
  AOI22_X1 U7487 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6556), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6605), .ZN(n6547) );
  OAI21_X1 U7488 ( .B1(n6783), .B2(n6558), .A(n6547), .ZN(U3206) );
  AOI22_X1 U7489 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6605), .ZN(n6548) );
  OAI21_X1 U7490 ( .B1(n6783), .B2(n6561), .A(n6548), .ZN(U3207) );
  AOI22_X1 U7491 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6556), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6605), .ZN(n6549) );
  OAI21_X1 U7492 ( .B1(n6550), .B2(n6558), .A(n6549), .ZN(U3208) );
  AOI22_X1 U7493 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6556), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6605), .ZN(n6551) );
  OAI21_X1 U7494 ( .B1(n6552), .B2(n6558), .A(n6551), .ZN(U3209) );
  AOI22_X1 U7495 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6556), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6605), .ZN(n6553) );
  OAI21_X1 U7496 ( .B1(n6555), .B2(n6558), .A(n6553), .ZN(U3210) );
  AOI22_X1 U7497 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6605), .ZN(n6554) );
  OAI21_X1 U7498 ( .B1(n6555), .B2(n6561), .A(n6554), .ZN(U3211) );
  AOI22_X1 U7499 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6556), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6605), .ZN(n6557) );
  OAI21_X1 U7500 ( .B1(n6562), .B2(n6558), .A(n6557), .ZN(U3212) );
  AOI22_X1 U7501 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6559), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6605), .ZN(n6560) );
  OAI21_X1 U7502 ( .B1(n6562), .B2(n6561), .A(n6560), .ZN(U3213) );
  MUX2_X1 U7503 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6605), .Z(U3445) );
  MUX2_X1 U7504 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6605), .Z(U3446) );
  MUX2_X1 U7505 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6605), .Z(U3447) );
  MUX2_X1 U7506 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6605), .Z(U3448) );
  OAI21_X1 U7507 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6565), .A(n6564), .ZN(
        n6563) );
  INV_X1 U7508 ( .A(n6563), .ZN(U3451) );
  INV_X1 U7509 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6585) );
  OAI21_X1 U7510 ( .B1(n6565), .B2(n6585), .A(n6564), .ZN(U3452) );
  OAI211_X1 U7511 ( .C1(n6569), .C2(n6568), .A(n6567), .B(n6566), .ZN(U3453)
         );
  INV_X1 U7512 ( .A(n6570), .ZN(n6573) );
  OAI22_X1 U7513 ( .A1(n6573), .A2(n6583), .B1(n6572), .B2(n6571), .ZN(n6574)
         );
  MUX2_X1 U7514 ( .A(n6575), .B(n6574), .S(n6581), .Z(U3456) );
  AOI21_X1 U7515 ( .B1(STATE2_REG_1__SCAN_IN), .B2(n6577), .A(n6576), .ZN(
        n6578) );
  OAI211_X1 U7516 ( .C1(n6579), .C2(n6583), .A(n6581), .B(n6578), .ZN(n6580)
         );
  OAI21_X1 U7517 ( .B1(n3507), .B2(n6581), .A(n6580), .ZN(n6582) );
  OAI21_X1 U7518 ( .B1(n6584), .B2(n6583), .A(n6582), .ZN(U3461) );
  INV_X1 U7519 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6752) );
  AOI22_X1 U7520 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(n6586), .B1(n6585), .B2(
        n6752), .ZN(n6589) );
  OAI211_X1 U7521 ( .C1(n6590), .C2(BYTEENABLE_REG_2__SCAN_IN), .A(n6587), .B(
        n6591), .ZN(n6588) );
  OAI21_X1 U7522 ( .B1(n6589), .B2(n6591), .A(n6588), .ZN(U3468) );
  OAI22_X1 U7523 ( .A1(n6591), .A2(REIP_REG_0__SCAN_IN), .B1(n6590), .B2(
        BYTEENABLE_REG_0__SCAN_IN), .ZN(n6592) );
  INV_X1 U7524 ( .A(n6592), .ZN(U3469) );
  NAND2_X1 U7525 ( .A1(n6605), .A2(W_R_N_REG_SCAN_IN), .ZN(n6593) );
  OAI21_X1 U7526 ( .B1(n6605), .B2(READREQUEST_REG_SCAN_IN), .A(n6593), .ZN(
        U3470) );
  AOI211_X1 U7527 ( .C1(n6597), .C2(n6596), .A(n6595), .B(n6594), .ZN(n6604)
         );
  OAI211_X1 U7528 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6599), .A(n6598), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6601) );
  AOI21_X1 U7529 ( .B1(n6601), .B2(STATE2_REG_0__SCAN_IN), .A(n6600), .ZN(
        n6603) );
  NAND2_X1 U7530 ( .A1(n6604), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6602) );
  OAI21_X1 U7531 ( .B1(n6604), .B2(n6603), .A(n6602), .ZN(U3472) );
  INV_X1 U7532 ( .A(M_IO_N_REG_SCAN_IN), .ZN(n6768) );
  AOI22_X1 U7533 ( .A1(n6607), .A2(n6606), .B1(n6768), .B2(n6605), .ZN(U3473)
         );
  AOI22_X1 U7534 ( .A1(n6609), .A2(DATAI_1_), .B1(n6608), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6614) );
  AOI22_X1 U7535 ( .A1(n6612), .A2(n6611), .B1(n6610), .B2(DATAI_17_), .ZN(
        n6613) );
  NAND2_X1 U7536 ( .A1(n6614), .A2(n6613), .ZN(n6803) );
  INV_X1 U7537 ( .A(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n6745) );
  INV_X1 U7538 ( .A(ADDRESS_REG_21__SCAN_IN), .ZN(n6616) );
  AOI22_X1 U7539 ( .A1(n6745), .A2(keyinput107), .B1(keyinput83), .B2(n6616), 
        .ZN(n6615) );
  OAI221_X1 U7540 ( .B1(n6745), .B2(keyinput107), .C1(n6616), .C2(keyinput83), 
        .A(n6615), .ZN(n6624) );
  INV_X1 U7541 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n6788) );
  AOI22_X1 U7542 ( .A1(n6788), .A2(keyinput106), .B1(keyinput111), .B2(n4553), 
        .ZN(n6617) );
  OAI221_X1 U7543 ( .B1(n6788), .B2(keyinput106), .C1(n4553), .C2(keyinput111), 
        .A(n6617), .ZN(n6623) );
  AOI22_X1 U7544 ( .A1(n4390), .A2(keyinput77), .B1(keyinput81), .B2(n6619), 
        .ZN(n6618) );
  OAI221_X1 U7545 ( .B1(n4390), .B2(keyinput77), .C1(n6619), .C2(keyinput81), 
        .A(n6618), .ZN(n6622) );
  INV_X1 U7546 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n6751) );
  AOI22_X1 U7547 ( .A1(n6751), .A2(keyinput97), .B1(n6781), .B2(keyinput99), 
        .ZN(n6620) );
  OAI221_X1 U7548 ( .B1(n6751), .B2(keyinput97), .C1(n6781), .C2(keyinput99), 
        .A(n6620), .ZN(n6621) );
  NOR4_X1 U7549 ( .A1(n6624), .A2(n6623), .A3(n6622), .A4(n6621), .ZN(n6661)
         );
  AOI22_X1 U7550 ( .A1(ADDRESS_REG_14__SCAN_IN), .A2(keyinput105), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput113), .ZN(n6625) );
  OAI221_X1 U7551 ( .B1(ADDRESS_REG_14__SCAN_IN), .B2(keyinput105), .C1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .C2(keyinput113), .A(n6625), .ZN(
        n6633) );
  AOI22_X1 U7552 ( .A1(EBX_REG_15__SCAN_IN), .A2(keyinput80), .B1(
        INSTQUEUE_REG_8__2__SCAN_IN), .B2(keyinput67), .ZN(n6626) );
  OAI221_X1 U7553 ( .B1(EBX_REG_15__SCAN_IN), .B2(keyinput80), .C1(
        INSTQUEUE_REG_8__2__SCAN_IN), .C2(keyinput67), .A(n6626), .ZN(n6632)
         );
  AOI22_X1 U7554 ( .A1(n6789), .A2(keyinput108), .B1(n6738), .B2(keyinput85), 
        .ZN(n6627) );
  OAI221_X1 U7555 ( .B1(n6789), .B2(keyinput108), .C1(n6738), .C2(keyinput85), 
        .A(n6627), .ZN(n6631) );
  INV_X1 U7556 ( .A(DATAI_11_), .ZN(n6629) );
  INV_X1 U7557 ( .A(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n6736) );
  AOI22_X1 U7558 ( .A1(n6629), .A2(keyinput119), .B1(n6736), .B2(keyinput115), 
        .ZN(n6628) );
  OAI221_X1 U7559 ( .B1(n6629), .B2(keyinput119), .C1(n6736), .C2(keyinput115), 
        .A(n6628), .ZN(n6630) );
  NOR4_X1 U7560 ( .A1(n6633), .A2(n6632), .A3(n6631), .A4(n6630), .ZN(n6660)
         );
  INV_X1 U7561 ( .A(DATAI_21_), .ZN(n6635) );
  AOI22_X1 U7562 ( .A1(n6636), .A2(keyinput65), .B1(keyinput87), .B2(n6635), 
        .ZN(n6634) );
  OAI221_X1 U7563 ( .B1(n6636), .B2(keyinput65), .C1(n6635), .C2(keyinput87), 
        .A(n6634), .ZN(n6646) );
  AOI22_X1 U7564 ( .A1(n4594), .A2(keyinput75), .B1(keyinput93), .B2(n6638), 
        .ZN(n6637) );
  OAI221_X1 U7565 ( .B1(n4594), .B2(keyinput75), .C1(n6638), .C2(keyinput93), 
        .A(n6637), .ZN(n6645) );
  INV_X1 U7566 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6770) );
  AOI22_X1 U7567 ( .A1(n6771), .A2(keyinput116), .B1(n6770), .B2(keyinput127), 
        .ZN(n6639) );
  OAI221_X1 U7568 ( .B1(n6771), .B2(keyinput116), .C1(n6770), .C2(keyinput127), 
        .A(n6639), .ZN(n6644) );
  INV_X1 U7569 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n6641) );
  AOI22_X1 U7570 ( .A1(n6642), .A2(keyinput88), .B1(n6641), .B2(keyinput82), 
        .ZN(n6640) );
  OAI221_X1 U7571 ( .B1(n6642), .B2(keyinput88), .C1(n6641), .C2(keyinput82), 
        .A(n6640), .ZN(n6643) );
  NOR4_X1 U7572 ( .A1(n6646), .A2(n6645), .A3(n6644), .A4(n6643), .ZN(n6659)
         );
  INV_X1 U7573 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6649) );
  AOI22_X1 U7574 ( .A1(n6649), .A2(keyinput125), .B1(keyinput94), .B2(n6648), 
        .ZN(n6647) );
  OAI221_X1 U7575 ( .B1(n6649), .B2(keyinput125), .C1(n6648), .C2(keyinput94), 
        .A(n6647), .ZN(n6657) );
  AOI22_X1 U7576 ( .A1(n6767), .A2(keyinput89), .B1(keyinput100), .B2(n6768), 
        .ZN(n6650) );
  OAI221_X1 U7577 ( .B1(n6767), .B2(keyinput89), .C1(n6768), .C2(keyinput100), 
        .A(n6650), .ZN(n6656) );
  INV_X1 U7578 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n6652) );
  AOI22_X1 U7579 ( .A1(n6652), .A2(keyinput68), .B1(keyinput110), .B2(n6741), 
        .ZN(n6651) );
  OAI221_X1 U7580 ( .B1(n6652), .B2(keyinput68), .C1(n6741), .C2(keyinput110), 
        .A(n6651), .ZN(n6655) );
  AOI22_X1 U7581 ( .A1(n6735), .A2(keyinput64), .B1(keyinput118), .B2(n6773), 
        .ZN(n6653) );
  OAI221_X1 U7582 ( .B1(n6735), .B2(keyinput64), .C1(n6773), .C2(keyinput118), 
        .A(n6653), .ZN(n6654) );
  NOR4_X1 U7583 ( .A1(n6657), .A2(n6656), .A3(n6655), .A4(n6654), .ZN(n6658)
         );
  NAND4_X1 U7584 ( .A1(n6661), .A2(n6660), .A3(n6659), .A4(n6658), .ZN(n6801)
         );
  AOI22_X1 U7585 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(keyinput84), .B1(
        INSTADDRPOINTER_REG_25__SCAN_IN), .B2(keyinput109), .ZN(n6662) );
  OAI221_X1 U7586 ( .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(keyinput84), 
        .C1(INSTADDRPOINTER_REG_25__SCAN_IN), .C2(keyinput109), .A(n6662), 
        .ZN(n6669) );
  AOI22_X1 U7587 ( .A1(DATAO_REG_20__SCAN_IN), .A2(keyinput73), .B1(
        EBX_REG_4__SCAN_IN), .B2(keyinput95), .ZN(n6663) );
  OAI221_X1 U7588 ( .B1(DATAO_REG_20__SCAN_IN), .B2(keyinput73), .C1(
        EBX_REG_4__SCAN_IN), .C2(keyinput95), .A(n6663), .ZN(n6668) );
  AOI22_X1 U7589 ( .A1(EAX_REG_4__SCAN_IN), .A2(keyinput121), .B1(
        INSTQUEUE_REG_7__7__SCAN_IN), .B2(keyinput112), .ZN(n6664) );
  OAI221_X1 U7590 ( .B1(EAX_REG_4__SCAN_IN), .B2(keyinput121), .C1(
        INSTQUEUE_REG_7__7__SCAN_IN), .C2(keyinput112), .A(n6664), .ZN(n6667)
         );
  AOI22_X1 U7591 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(keyinput70), .B1(
        INSTQUEUE_REG_13__5__SCAN_IN), .B2(keyinput69), .ZN(n6665) );
  OAI221_X1 U7592 ( .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .B2(keyinput70), .C1(
        INSTQUEUE_REG_13__5__SCAN_IN), .C2(keyinput69), .A(n6665), .ZN(n6666)
         );
  NOR4_X1 U7593 ( .A1(n6669), .A2(n6668), .A3(n6667), .A4(n6666), .ZN(n6697)
         );
  AOI22_X1 U7594 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(keyinput71), .B1(
        EBX_REG_20__SCAN_IN), .B2(keyinput79), .ZN(n6670) );
  OAI221_X1 U7595 ( .B1(INSTADDRPOINTER_REG_15__SCAN_IN), .B2(keyinput71), 
        .C1(EBX_REG_20__SCAN_IN), .C2(keyinput79), .A(n6670), .ZN(n6677) );
  AOI22_X1 U7596 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(keyinput103), .B1(
        STATE2_REG_0__SCAN_IN), .B2(keyinput101), .ZN(n6671) );
  OAI221_X1 U7597 ( .B1(INSTQUEUE_REG_0__7__SCAN_IN), .B2(keyinput103), .C1(
        STATE2_REG_0__SCAN_IN), .C2(keyinput101), .A(n6671), .ZN(n6676) );
  AOI22_X1 U7598 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(keyinput126), .B1(
        INSTQUEUE_REG_8__4__SCAN_IN), .B2(keyinput90), .ZN(n6672) );
  OAI221_X1 U7599 ( .B1(DATAWIDTH_REG_29__SCAN_IN), .B2(keyinput126), .C1(
        INSTQUEUE_REG_8__4__SCAN_IN), .C2(keyinput90), .A(n6672), .ZN(n6675)
         );
  AOI22_X1 U7600 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(keyinput76), .B1(
        MEMORYFETCH_REG_SCAN_IN), .B2(keyinput72), .ZN(n6673) );
  OAI221_X1 U7601 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(keyinput76), .C1(
        MEMORYFETCH_REG_SCAN_IN), .C2(keyinput72), .A(n6673), .ZN(n6674) );
  NOR4_X1 U7602 ( .A1(n6677), .A2(n6676), .A3(n6675), .A4(n6674), .ZN(n6696)
         );
  AOI22_X1 U7603 ( .A1(LWORD_REG_15__SCAN_IN), .A2(keyinput124), .B1(
        INSTQUEUE_REG_12__0__SCAN_IN), .B2(keyinput78), .ZN(n6678) );
  OAI221_X1 U7604 ( .B1(LWORD_REG_15__SCAN_IN), .B2(keyinput124), .C1(
        INSTQUEUE_REG_12__0__SCAN_IN), .C2(keyinput78), .A(n6678), .ZN(n6685)
         );
  AOI22_X1 U7605 ( .A1(DATAO_REG_13__SCAN_IN), .A2(keyinput117), .B1(
        STATE2_REG_1__SCAN_IN), .B2(keyinput91), .ZN(n6679) );
  OAI221_X1 U7606 ( .B1(DATAO_REG_13__SCAN_IN), .B2(keyinput117), .C1(
        STATE2_REG_1__SCAN_IN), .C2(keyinput91), .A(n6679), .ZN(n6684) );
  AOI22_X1 U7607 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(keyinput96), .B1(
        INSTQUEUE_REG_0__3__SCAN_IN), .B2(keyinput104), .ZN(n6680) );
  OAI221_X1 U7608 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput96), 
        .C1(INSTQUEUE_REG_0__3__SCAN_IN), .C2(keyinput104), .A(n6680), .ZN(
        n6683) );
  AOI22_X1 U7609 ( .A1(DATAI_3_), .A2(keyinput92), .B1(DATAI_27_), .B2(
        keyinput114), .ZN(n6681) );
  OAI221_X1 U7610 ( .B1(DATAI_3_), .B2(keyinput92), .C1(DATAI_27_), .C2(
        keyinput114), .A(n6681), .ZN(n6682) );
  NOR4_X1 U7611 ( .A1(n6685), .A2(n6684), .A3(n6683), .A4(n6682), .ZN(n6695)
         );
  AOI22_X1 U7612 ( .A1(DATAI_28_), .A2(keyinput66), .B1(
        INSTQUEUE_REG_5__0__SCAN_IN), .B2(keyinput122), .ZN(n6686) );
  OAI221_X1 U7613 ( .B1(DATAI_28_), .B2(keyinput66), .C1(
        INSTQUEUE_REG_5__0__SCAN_IN), .C2(keyinput122), .A(n6686), .ZN(n6693)
         );
  AOI22_X1 U7614 ( .A1(REIP_REG_24__SCAN_IN), .A2(keyinput98), .B1(
        INSTQUEUE_REG_9__7__SCAN_IN), .B2(keyinput102), .ZN(n6687) );
  OAI221_X1 U7615 ( .B1(REIP_REG_24__SCAN_IN), .B2(keyinput98), .C1(
        INSTQUEUE_REG_9__7__SCAN_IN), .C2(keyinput102), .A(n6687), .ZN(n6692)
         );
  AOI22_X1 U7616 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(keyinput74), .B1(
        INSTQUEUE_REG_6__5__SCAN_IN), .B2(keyinput86), .ZN(n6688) );
  OAI221_X1 U7617 ( .B1(INSTQUEUE_REG_6__4__SCAN_IN), .B2(keyinput74), .C1(
        INSTQUEUE_REG_6__5__SCAN_IN), .C2(keyinput86), .A(n6688), .ZN(n6691)
         );
  AOI22_X1 U7618 ( .A1(ADDRESS_REG_6__SCAN_IN), .A2(keyinput120), .B1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput123), .ZN(n6689) );
  OAI221_X1 U7619 ( .B1(ADDRESS_REG_6__SCAN_IN), .B2(keyinput120), .C1(
        PHYADDRPOINTER_REG_19__SCAN_IN), .C2(keyinput123), .A(n6689), .ZN(
        n6690) );
  NOR4_X1 U7620 ( .A1(n6693), .A2(n6692), .A3(n6691), .A4(n6690), .ZN(n6694)
         );
  NAND4_X1 U7621 ( .A1(n6697), .A2(n6696), .A3(n6695), .A4(n6694), .ZN(n6800)
         );
  OAI22_X1 U7622 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(keyinput58), .B1(
        keyinput53), .B2(DATAO_REG_13__SCAN_IN), .ZN(n6698) );
  AOI221_X1 U7623 ( .B1(INSTQUEUE_REG_5__0__SCAN_IN), .B2(keyinput58), .C1(
        DATAO_REG_13__SCAN_IN), .C2(keyinput53), .A(n6698), .ZN(n6705) );
  OAI22_X1 U7624 ( .A1(EBX_REG_4__SCAN_IN), .A2(keyinput31), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(keyinput1), .ZN(n6699) );
  AOI221_X1 U7625 ( .B1(EBX_REG_4__SCAN_IN), .B2(keyinput31), .C1(keyinput1), 
        .C2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n6699), .ZN(n6704) );
  OAI22_X1 U7626 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(keyinput20), .B1(
        keyinput41), .B2(ADDRESS_REG_14__SCAN_IN), .ZN(n6700) );
  AOI221_X1 U7627 ( .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(keyinput20), 
        .C1(ADDRESS_REG_14__SCAN_IN), .C2(keyinput41), .A(n6700), .ZN(n6703)
         );
  OAI22_X1 U7628 ( .A1(PHYADDRPOINTER_REG_19__SCAN_IN), .A2(keyinput59), .B1(
        DATAI_11_), .B2(keyinput55), .ZN(n6701) );
  AOI221_X1 U7629 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput59), .C1(
        keyinput55), .C2(DATAI_11_), .A(n6701), .ZN(n6702) );
  NAND4_X1 U7630 ( .A1(n6705), .A2(n6704), .A3(n6703), .A4(n6702), .ZN(n6733)
         );
  OAI22_X1 U7631 ( .A1(EBX_REG_23__SCAN_IN), .A2(keyinput24), .B1(DATAI_28_), 
        .B2(keyinput2), .ZN(n6706) );
  AOI221_X1 U7632 ( .B1(EBX_REG_23__SCAN_IN), .B2(keyinput24), .C1(keyinput2), 
        .C2(DATAI_28_), .A(n6706), .ZN(n6713) );
  OAI22_X1 U7633 ( .A1(INSTQUEUE_REG_4__3__SCAN_IN), .A2(keyinput47), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(keyinput6), .ZN(n6707) );
  AOI221_X1 U7634 ( .B1(INSTQUEUE_REG_4__3__SCAN_IN), .B2(keyinput47), .C1(
        keyinput6), .C2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n6707), .ZN(n6712)
         );
  OAI22_X1 U7635 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(keyinput10), .B1(
        DATAWIDTH_REG_27__SCAN_IN), .B2(keyinput17), .ZN(n6708) );
  AOI221_X1 U7636 ( .B1(INSTQUEUE_REG_6__4__SCAN_IN), .B2(keyinput10), .C1(
        keyinput17), .C2(DATAWIDTH_REG_27__SCAN_IN), .A(n6708), .ZN(n6711) );
  OAI22_X1 U7637 ( .A1(EBX_REG_29__SCAN_IN), .A2(keyinput30), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(keyinput29), .ZN(n6709) );
  AOI221_X1 U7638 ( .B1(EBX_REG_29__SCAN_IN), .B2(keyinput30), .C1(keyinput29), 
        .C2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n6709), .ZN(n6710) );
  NAND4_X1 U7639 ( .A1(n6713), .A2(n6712), .A3(n6711), .A4(n6710), .ZN(n6732)
         );
  OAI22_X1 U7640 ( .A1(DATAI_27_), .A2(keyinput50), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(keyinput19), .ZN(n6714) );
  AOI221_X1 U7641 ( .B1(DATAI_27_), .B2(keyinput50), .C1(keyinput19), .C2(
        ADDRESS_REG_21__SCAN_IN), .A(n6714), .ZN(n6721) );
  OAI22_X1 U7642 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(keyinput5), .B1(
        keyinput9), .B2(DATAO_REG_20__SCAN_IN), .ZN(n6715) );
  AOI221_X1 U7643 ( .B1(INSTQUEUE_REG_13__5__SCAN_IN), .B2(keyinput5), .C1(
        DATAO_REG_20__SCAN_IN), .C2(keyinput9), .A(n6715), .ZN(n6720) );
  OAI22_X1 U7644 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(keyinput22), .B1(
        INSTQUEUE_REG_5__2__SCAN_IN), .B2(keyinput61), .ZN(n6716) );
  AOI221_X1 U7645 ( .B1(INSTQUEUE_REG_6__5__SCAN_IN), .B2(keyinput22), .C1(
        keyinput61), .C2(INSTQUEUE_REG_5__2__SCAN_IN), .A(n6716), .ZN(n6719)
         );
  OAI22_X1 U7646 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(keyinput32), .B1(
        keyinput23), .B2(DATAI_21_), .ZN(n6717) );
  AOI221_X1 U7647 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput32), 
        .C1(DATAI_21_), .C2(keyinput23), .A(n6717), .ZN(n6718) );
  NAND4_X1 U7648 ( .A1(n6721), .A2(n6720), .A3(n6719), .A4(n6718), .ZN(n6731)
         );
  OAI22_X1 U7649 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(keyinput18), .B1(
        keyinput38), .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n6722) );
  AOI221_X1 U7650 ( .B1(INSTQUEUE_REG_9__4__SCAN_IN), .B2(keyinput18), .C1(
        INSTQUEUE_REG_9__7__SCAN_IN), .C2(keyinput38), .A(n6722), .ZN(n6729)
         );
  OAI22_X1 U7651 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(keyinput40), .B1(
        keyinput16), .B2(EBX_REG_15__SCAN_IN), .ZN(n6723) );
  AOI221_X1 U7652 ( .B1(INSTQUEUE_REG_0__3__SCAN_IN), .B2(keyinput40), .C1(
        EBX_REG_15__SCAN_IN), .C2(keyinput16), .A(n6723), .ZN(n6728) );
  OAI22_X1 U7653 ( .A1(MEMORYFETCH_REG_SCAN_IN), .A2(keyinput8), .B1(
        DATAO_REG_1__SCAN_IN), .B2(keyinput4), .ZN(n6724) );
  AOI221_X1 U7654 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(keyinput8), .C1(
        keyinput4), .C2(DATAO_REG_1__SCAN_IN), .A(n6724), .ZN(n6727) );
  OAI22_X1 U7655 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(keyinput48), .B1(
        INSTADDRPOINTER_REG_15__SCAN_IN), .B2(keyinput7), .ZN(n6725) );
  AOI221_X1 U7656 ( .B1(INSTQUEUE_REG_7__7__SCAN_IN), .B2(keyinput48), .C1(
        keyinput7), .C2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n6725), .ZN(n6726) );
  NAND4_X1 U7657 ( .A1(n6729), .A2(n6728), .A3(n6727), .A4(n6726), .ZN(n6730)
         );
  NOR4_X1 U7658 ( .A1(n6733), .A2(n6732), .A3(n6731), .A4(n6730), .ZN(n6799)
         );
  AOI22_X1 U7659 ( .A1(n6736), .A2(keyinput51), .B1(keyinput0), .B2(n6735), 
        .ZN(n6734) );
  OAI221_X1 U7660 ( .B1(n6736), .B2(keyinput51), .C1(n6735), .C2(keyinput0), 
        .A(n6734), .ZN(n6749) );
  AOI22_X1 U7661 ( .A1(n6739), .A2(keyinput56), .B1(n6738), .B2(keyinput21), 
        .ZN(n6737) );
  OAI221_X1 U7662 ( .B1(n6739), .B2(keyinput56), .C1(n6738), .C2(keyinput21), 
        .A(n6737), .ZN(n6748) );
  AOI22_X1 U7663 ( .A1(n6742), .A2(keyinput28), .B1(keyinput46), .B2(n6741), 
        .ZN(n6740) );
  OAI221_X1 U7664 ( .B1(n6742), .B2(keyinput28), .C1(n6741), .C2(keyinput46), 
        .A(n6740), .ZN(n6747) );
  AOI22_X1 U7665 ( .A1(n6745), .A2(keyinput43), .B1(keyinput45), .B2(n6744), 
        .ZN(n6743) );
  OAI221_X1 U7666 ( .B1(n6745), .B2(keyinput43), .C1(n6744), .C2(keyinput45), 
        .A(n6743), .ZN(n6746) );
  NOR4_X1 U7667 ( .A1(n6749), .A2(n6748), .A3(n6747), .A4(n6746), .ZN(n6797)
         );
  AOI22_X1 U7668 ( .A1(n6752), .A2(keyinput12), .B1(keyinput33), .B2(n6751), 
        .ZN(n6750) );
  OAI221_X1 U7669 ( .B1(n6752), .B2(keyinput12), .C1(n6751), .C2(keyinput33), 
        .A(n6750), .ZN(n6763) );
  AOI22_X1 U7670 ( .A1(EBX_REG_20__SCAN_IN), .A2(keyinput15), .B1(n6754), .B2(
        keyinput60), .ZN(n6753) );
  OAI221_X1 U7671 ( .B1(EBX_REG_20__SCAN_IN), .B2(keyinput15), .C1(n6754), 
        .C2(keyinput60), .A(n6753), .ZN(n6762) );
  INV_X1 U7672 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6756) );
  AOI22_X1 U7673 ( .A1(n4390), .A2(keyinput13), .B1(n6756), .B2(keyinput26), 
        .ZN(n6755) );
  OAI221_X1 U7674 ( .B1(n4390), .B2(keyinput13), .C1(n6756), .C2(keyinput26), 
        .A(n6755), .ZN(n6761) );
  AOI22_X1 U7675 ( .A1(n6759), .A2(keyinput57), .B1(n6758), .B2(keyinput49), 
        .ZN(n6757) );
  OAI221_X1 U7676 ( .B1(n6759), .B2(keyinput57), .C1(n6758), .C2(keyinput49), 
        .A(n6757), .ZN(n6760) );
  NOR4_X1 U7677 ( .A1(n6763), .A2(n6762), .A3(n6761), .A4(n6760), .ZN(n6796)
         );
  AOI22_X1 U7678 ( .A1(n6765), .A2(keyinput27), .B1(keyinput11), .B2(n4594), 
        .ZN(n6764) );
  OAI221_X1 U7679 ( .B1(n6765), .B2(keyinput27), .C1(n4594), .C2(keyinput11), 
        .A(n6764), .ZN(n6778) );
  AOI22_X1 U7680 ( .A1(n6768), .A2(keyinput36), .B1(n6767), .B2(keyinput25), 
        .ZN(n6766) );
  OAI221_X1 U7681 ( .B1(n6768), .B2(keyinput36), .C1(n6767), .C2(keyinput25), 
        .A(n6766), .ZN(n6777) );
  AOI22_X1 U7682 ( .A1(n6771), .A2(keyinput52), .B1(n6770), .B2(keyinput63), 
        .ZN(n6769) );
  OAI221_X1 U7683 ( .B1(n6771), .B2(keyinput52), .C1(n6770), .C2(keyinput63), 
        .A(n6769), .ZN(n6776) );
  INV_X1 U7684 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n6774) );
  AOI22_X1 U7685 ( .A1(n6774), .A2(keyinput14), .B1(keyinput54), .B2(n6773), 
        .ZN(n6772) );
  OAI221_X1 U7686 ( .B1(n6774), .B2(keyinput14), .C1(n6773), .C2(keyinput54), 
        .A(n6772), .ZN(n6775) );
  NOR4_X1 U7687 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .ZN(n6795)
         );
  AOI22_X1 U7688 ( .A1(n6781), .A2(keyinput35), .B1(n6780), .B2(keyinput37), 
        .ZN(n6779) );
  OAI221_X1 U7689 ( .B1(n6781), .B2(keyinput35), .C1(n6780), .C2(keyinput37), 
        .A(n6779), .ZN(n6793) );
  AOI22_X1 U7690 ( .A1(n6784), .A2(keyinput62), .B1(n6783), .B2(keyinput34), 
        .ZN(n6782) );
  OAI221_X1 U7691 ( .B1(n6784), .B2(keyinput62), .C1(n6783), .C2(keyinput34), 
        .A(n6782), .ZN(n6792) );
  INV_X1 U7692 ( .A(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n6786) );
  AOI22_X1 U7693 ( .A1(n4399), .A2(keyinput39), .B1(keyinput3), .B2(n6786), 
        .ZN(n6785) );
  OAI221_X1 U7694 ( .B1(n4399), .B2(keyinput39), .C1(n6786), .C2(keyinput3), 
        .A(n6785), .ZN(n6791) );
  AOI22_X1 U7695 ( .A1(n6789), .A2(keyinput44), .B1(n6788), .B2(keyinput42), 
        .ZN(n6787) );
  OAI221_X1 U7696 ( .B1(n6789), .B2(keyinput44), .C1(n6788), .C2(keyinput42), 
        .A(n6787), .ZN(n6790) );
  NOR4_X1 U7697 ( .A1(n6793), .A2(n6792), .A3(n6791), .A4(n6790), .ZN(n6794)
         );
  AND4_X1 U7698 ( .A1(n6797), .A2(n6796), .A3(n6795), .A4(n6794), .ZN(n6798)
         );
  OAI211_X1 U7699 ( .C1(n6801), .C2(n6800), .A(n6799), .B(n6798), .ZN(n6802)
         );
  XNOR2_X1 U7700 ( .A(n6803), .B(n6802), .ZN(U2874) );
  AND2_X2 U3943 ( .A1(n4220), .A2(n4418), .ZN(n3309) );
  AOI22_X1 U3941 ( .A1(n3243), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3308), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3058) );
  AND4_X1 U3947 ( .A1(n3058), .A2(n3057), .A3(n3056), .A4(n3055), .ZN(n3068)
         );
  AND4_X1 U4057 ( .A1(n3172), .A2(n3171), .A3(n3170), .A4(n3169), .ZN(n3183)
         );
  OR2_X1 U3581 ( .A1(n3372), .A2(n3371), .ZN(n3374) );
  INV_X4 U3533 ( .A(n3500), .ZN(n5890) );
  NAND2_X1 U6345 ( .A1(n5511), .A2(n5289), .ZN(n5331) );
  CLKBUF_X1 U3502 ( .A(n3290), .Z(n3273) );
  CLKBUF_X1 U3511 ( .A(n3308), .Z(n5105) );
  XNOR2_X1 U3512 ( .A(n3261), .B(n3260), .ZN(n3372) );
  CLKBUF_X1 U3544 ( .A(n3146), .Z(n3271) );
  CLKBUF_X2 U3575 ( .A(n3187), .Z(n4187) );
  AND2_X1 U3612 ( .A1(n3141), .A2(n3140), .ZN(n3941) );
  CLKBUF_X1 U3667 ( .A(n3983), .Z(n3031) );
  CLKBUF_X1 U3732 ( .A(n3322), .Z(n3323) );
  CLKBUF_X1 U3853 ( .A(n5612), .Z(n5624) );
  CLKBUF_X1 U3873 ( .A(n3563), .Z(n5744) );
  CLKBUF_X1 U4029 ( .A(n6120), .Z(n6131) );
  CLKBUF_X1 U4126 ( .A(n3580), .Z(n5742) );
  CLKBUF_X1 U4135 ( .A(n3569), .Z(n3032) );
endmodule

