

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787;

  INV_X1 U2245 ( .A(n4024), .ZN(n3132) );
  NAND2_X1 U2246 ( .A1(n3599), .A2(IR_REG_31__SCAN_IN), .ZN(n2087) );
  CLKBUF_X1 U2247 ( .A(n3841), .Z(n2003) );
  NOR2_X1 U2248 ( .A1(n2988), .A2(n4737), .ZN(n3841) );
  CLKBUF_X3 U2249 ( .A(n2972), .Z(n3650) );
  INV_X1 U2250 ( .A(n3658), .ZN(n3645) );
  INV_X2 U2251 ( .A(n2347), .ZN(n2758) );
  INV_X1 U2252 ( .A(n2345), .ZN(n2346) );
  NAND2_X1 U2253 ( .A1(n4030), .A2(n2882), .ZN(n2939) );
  AOI21_X1 U2254 ( .B1(n4172), .B2(n3902), .A(n3907), .ZN(n2796) );
  INV_X1 U2255 ( .A(n4018), .ZN(n3338) );
  OR2_X1 U2256 ( .A1(n2747), .A2(n2800), .ZN(n2802) );
  CLKBUF_X3 U2257 ( .A(n2355), .Z(n3510) );
  AND4_X1 U2258 ( .A1(n2371), .A2(n2370), .A3(n2369), .A4(n2368), .ZN(n3160)
         );
  AOI211_X1 U2259 ( .C1(n3114), .C2(n3113), .A(n4114), .B(n3210), .ZN(n3115)
         );
  AND4_X1 U2260 ( .A1(n2341), .A2(n2340), .A3(n2339), .A4(n2338), .ZN(n3068)
         );
  INV_X1 U2261 ( .A(n2705), .ZN(n4687) );
  NAND2_X2 U2262 ( .A1(n2926), .A2(n3123), .ZN(n3552) );
  INV_X1 U2263 ( .A(n3174), .ZN(n3604) );
  INV_X4 U2264 ( .A(n3174), .ZN(n3655) );
  NAND4_X2 U2265 ( .A1(n2351), .A2(n2350), .A3(n2349), .A4(n2348), .ZN(n4024)
         );
  OR2_X1 U2266 ( .A1(n2346), .A2(n3079), .ZN(n2349) );
  NAND2_X2 U2267 ( .A1(n3149), .A2(n3148), .ZN(n3157) );
  AOI22_X2 U2268 ( .A1(n3146), .A2(n3145), .B1(n3144), .B2(n3143), .ZN(n3149)
         );
  NAND2_X2 U2269 ( .A1(n4050), .A2(n2905), .ZN(n2912) );
  INV_X2 U2270 ( .A(n2317), .ZN(n2127) );
  XNOR2_X2 U2271 ( .A(n2156), .B(n2155), .ZN(n4059) );
  XNOR2_X2 U2272 ( .A(n2106), .B(IR_REG_2__SCAN_IN), .ZN(n4697) );
  OAI21_X2 U2273 ( .B1(n3159), .B2(n3158), .A(n3157), .ZN(n3164) );
  NAND2_X1 U2274 ( .A1(n3776), .A2(n3777), .ZN(n3775) );
  NOR2_X1 U2275 ( .A1(n2930), .A2(n2074), .ZN(n2969) );
  NAND2_X1 U2276 ( .A1(n2644), .A2(n2643), .ZN(n2728) );
  NAND3_X2 U2277 ( .A1(n2708), .A2(n2707), .A3(n2844), .ZN(n3123) );
  INV_X1 U2278 ( .A(n2168), .ZN(n4729) );
  OR2_X1 U2279 ( .A1(n2787), .A2(n4782), .ZN(n2791) );
  OR2_X1 U2280 ( .A1(n2787), .A2(n4784), .ZN(n2786) );
  NAND2_X1 U2281 ( .A1(n2160), .A2(n2158), .ZN(n3469) );
  NOR2_X1 U2282 ( .A1(n2128), .A2(n3901), .ZN(n4172) );
  OAI21_X1 U2283 ( .B1(n2165), .B2(n4092), .A(n2047), .ZN(n2159) );
  OAI21_X1 U2284 ( .B1(n2726), .B2(n4139), .A(n2780), .ZN(n4145) );
  OAI22_X1 U2285 ( .A1(n4352), .A2(n2061), .B1(n2062), .B2(n2528), .ZN(n4305)
         );
  NAND2_X1 U2286 ( .A1(n3131), .A2(n3130), .ZN(n3146) );
  NAND2_X1 U2287 ( .A1(n3028), .A2(n2375), .ZN(n2213) );
  OR2_X1 U2288 ( .A1(n2907), .A2(n2177), .ZN(n2176) );
  INV_X2 U2289 ( .A(n3552), .ZN(n3174) );
  INV_X2 U2290 ( .A(n3533), .ZN(n3605) );
  AND2_X1 U2291 ( .A1(n3848), .A2(n3850), .ZN(n3936) );
  NAND2_X1 U2292 ( .A1(n2900), .A2(n2899), .ZN(n2902) );
  CLKBUF_X1 U2293 ( .A(n2334), .Z(n3011) );
  INV_X1 U2294 ( .A(n2334), .ZN(n2975) );
  INV_X2 U2295 ( .A(n2333), .ZN(n2973) );
  INV_X1 U2296 ( .A(n2997), .ZN(n2929) );
  NAND2_X1 U2297 ( .A1(n2885), .A2(REG1_REG_3__SCAN_IN), .ZN(n2900) );
  CLKBUF_X1 U2298 ( .A(n2953), .Z(n4316) );
  OAI21_X1 U2299 ( .B1(n3506), .B2(n2231), .A(n2336), .ZN(n2997) );
  XNOR2_X1 U2300 ( .A(n2898), .B(n2884), .ZN(n2885) );
  NAND2_X1 U2301 ( .A1(n2938), .A2(n2883), .ZN(n2898) );
  OR2_X1 U2302 ( .A1(n2355), .A2(n2871), .ZN(n2126) );
  NAND2_X1 U2303 ( .A1(n2710), .A2(IR_REG_31__SCAN_IN), .ZN(n2696) );
  NAND2_X1 U2304 ( .A1(n2755), .A2(IR_REG_31__SCAN_IN), .ZN(n2703) );
  XNOR2_X1 U2305 ( .A(n2699), .B(n2698), .ZN(n2706) );
  XNOR2_X1 U2306 ( .A(n2655), .B(n2654), .ZN(n4004) );
  OAI21_X1 U2307 ( .B1(n2695), .B2(IR_REG_22__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2709) );
  NAND2_X1 U2308 ( .A1(n2645), .A2(IR_REG_31__SCAN_IN), .ZN(n2647) );
  OR2_X1 U2309 ( .A1(n2636), .A2(n2648), .ZN(n2645) );
  AND3_X1 U2310 ( .A1(n2424), .A2(n2320), .A3(n4576), .ZN(n2107) );
  NOR2_X1 U2311 ( .A1(IR_REG_9__SCAN_IN), .A2(n2436), .ZN(n2524) );
  AND2_X1 U2312 ( .A1(n2650), .A2(n2316), .ZN(n2284) );
  AND3_X1 U2313 ( .A1(n2315), .A2(n2523), .A3(n2314), .ZN(n2650) );
  NAND4_X1 U2314 ( .A1(n2305), .A2(n2307), .A3(n2306), .A4(n4563), .ZN(n2649)
         );
  NAND2_X1 U2315 ( .A1(n2358), .A2(n2310), .ZN(n2311) );
  AND2_X1 U2316 ( .A1(n2423), .A2(n2422), .ZN(n2435) );
  NOR2_X1 U2317 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2306)
         );
  NOR2_X1 U2318 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2315)
         );
  NOR2_X1 U2319 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2305)
         );
  NOR2_X1 U2320 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2307)
         );
  NOR2_X2 U2321 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2322)
         );
  NOR2_X1 U2322 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2523)
         );
  INV_X1 U2323 ( .A(IR_REG_2__SCAN_IN), .ZN(n2309) );
  NOR2_X1 U2324 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2423)
         );
  INV_X1 U2325 ( .A(IR_REG_1__SCAN_IN), .ZN(n2232) );
  INV_X1 U2326 ( .A(IR_REG_3__SCAN_IN), .ZN(n2358) );
  INV_X1 U2327 ( .A(IR_REG_4__SCAN_IN), .ZN(n2310) );
  OR2_X4 U2328 ( .A1(n2127), .A2(n2318), .ZN(n2353) );
  INV_X1 U2329 ( .A(n3533), .ZN(n2004) );
  NAND2_X1 U2330 ( .A1(n2980), .A2(n2981), .ZN(n3131) );
  AND2_X4 U2331 ( .A1(n3660), .A2(n3200), .ZN(n3533) );
  AND2_X2 U2332 ( .A1(n3123), .A2(n2964), .ZN(n3660) );
  NOR2_X4 U2333 ( .A1(n4363), .A2(n4345), .ZN(n4342) );
  OR2_X2 U2334 ( .A1(n3406), .A2(n4361), .ZN(n4363) );
  NAND2_X1 U2335 ( .A1(n4155), .A2(n3670), .ZN(n3912) );
  NAND2_X1 U2336 ( .A1(n3310), .A2(n2220), .ZN(n2069) );
  INV_X1 U2337 ( .A(n2964), .ZN(n2926) );
  NAND2_X1 U2338 ( .A1(n2084), .A2(n2082), .ZN(n2080) );
  OR2_X1 U2339 ( .A1(n2607), .A2(n4647), .ZN(n2628) );
  INV_X1 U2340 ( .A(n2353), .ZN(n2685) );
  AOI21_X1 U2341 ( .B1(n2006), .B2(n2447), .A(n2029), .ZN(n2220) );
  AND2_X1 U2342 ( .A1(n3040), .A2(n2059), .ZN(n2058) );
  AND2_X1 U2343 ( .A1(n2343), .A2(n2060), .ZN(n2059) );
  NAND2_X1 U2344 ( .A1(n3132), .A2(n3135), .ZN(n2060) );
  NAND2_X1 U2345 ( .A1(n3911), .A2(n3912), .ZN(n3989) );
  NAND2_X1 U2346 ( .A1(n2919), .A2(REG2_REG_6__SCAN_IN), .ZN(n2100) );
  OAI21_X1 U2347 ( .B1(n4100), .B2(n3489), .A(n4094), .ZN(n3490) );
  INV_X1 U2348 ( .A(n2159), .ZN(n2158) );
  AND2_X1 U2349 ( .A1(n4183), .A2(n3827), .ZN(n2622) );
  INV_X1 U2350 ( .A(n2217), .ZN(n2216) );
  OAI21_X1 U2351 ( .B1(n4304), .B2(n2218), .A(n2554), .ZN(n2217) );
  NAND2_X1 U2352 ( .A1(n3854), .A2(n3851), .ZN(n2663) );
  AOI21_X1 U2353 ( .B1(n2270), .B2(n2268), .A(n2267), .ZN(n2266) );
  INV_X1 U2354 ( .A(n3811), .ZN(n2267) );
  INV_X1 U2355 ( .A(n2271), .ZN(n2268) );
  INV_X1 U2356 ( .A(n2270), .ZN(n2269) );
  NAND2_X1 U2357 ( .A1(n2397), .A2(REG3_REG_8__SCAN_IN), .ZN(n2416) );
  INV_X1 U2358 ( .A(n2399), .ZN(n2397) );
  INV_X1 U2359 ( .A(n3592), .ZN(n3590) );
  OAI22_X1 U2360 ( .A1(n2973), .A2(n3552), .B1(n2975), .B2(n2972), .ZN(n2974)
         );
  OR3_X1 U2361 ( .A1(n2599), .A2(n3625), .A3(n3770), .ZN(n2607) );
  AND3_X1 U2362 ( .A1(n2952), .A2(n2951), .A3(n2950), .ZN(n2990) );
  NAND2_X1 U2363 ( .A1(n2127), .A2(REG0_REG_1__SCAN_IN), .ZN(n2125) );
  NAND2_X1 U2364 ( .A1(n4053), .A2(n2183), .ZN(n2917) );
  OR2_X1 U2365 ( .A1(n4047), .A2(n2895), .ZN(n2183) );
  AOI21_X1 U2366 ( .B1(n3380), .B2(n2092), .A(n2020), .ZN(n2096) );
  NOR2_X1 U2367 ( .A1(n3381), .A2(n2091), .ZN(n2090) );
  NAND2_X1 U2368 ( .A1(n2130), .A2(n2129), .ZN(n2128) );
  INV_X1 U2369 ( .A(n3925), .ZN(n2129) );
  OAI21_X1 U2370 ( .B1(n4248), .B2(n3976), .A(n3981), .ZN(n2130) );
  NAND2_X1 U2371 ( .A1(n2147), .A2(REG3_REG_23__SCAN_IN), .ZN(n2599) );
  NAND2_X1 U2372 ( .A1(n2148), .A2(REG3_REG_20__SCAN_IN), .ZN(n2573) );
  OAI21_X1 U2373 ( .B1(n4261), .B2(n2563), .A(n2562), .ZN(n4250) );
  AOI21_X1 U2374 ( .B1(n4356), .B2(n2496), .A(n2028), .ZN(n4352) );
  AOI21_X1 U2375 ( .B1(n2007), .B2(n2121), .A(n2038), .ZN(n2117) );
  NAND2_X1 U2376 ( .A1(n3182), .A2(n3864), .ZN(n2666) );
  AND2_X1 U2377 ( .A1(n2767), .A2(n2766), .ZN(n2774) );
  NAND2_X1 U2378 ( .A1(n2684), .A2(n4338), .ZN(n4136) );
  NAND2_X1 U2379 ( .A1(n2795), .A2(n3911), .ZN(n2753) );
  NOR2_X1 U2380 ( .A1(n2642), .A2(n2641), .ZN(n2643) );
  NAND2_X1 U2381 ( .A1(n2692), .A2(n2691), .ZN(n4143) );
  NAND2_X1 U2382 ( .A1(n2619), .A2(n2618), .ZN(n4015) );
  INV_X1 U2383 ( .A(n3864), .ZN(n2120) );
  INV_X1 U2384 ( .A(n3865), .ZN(n2238) );
  AND2_X1 U2385 ( .A1(n2237), .A2(n3886), .ZN(n2236) );
  OR2_X1 U2386 ( .A1(n2239), .A2(n2238), .ZN(n2237) );
  INV_X1 U2387 ( .A(n2636), .ZN(n2321) );
  NOR2_X1 U2388 ( .A1(n2299), .A2(n3236), .ZN(n2289) );
  INV_X1 U2389 ( .A(n3636), .ZN(n3613) );
  NAND2_X1 U2390 ( .A1(n2231), .A2(IR_REG_1__SCAN_IN), .ZN(n2185) );
  NAND2_X1 U2391 ( .A1(n2192), .A2(n2013), .ZN(n3379) );
  OAI211_X1 U2392 ( .C1(n2100), .C2(n2920), .A(n2101), .B(n2099), .ZN(n2192)
         );
  NOR2_X1 U2393 ( .A1(n2196), .A2(n2194), .ZN(n2193) );
  OR2_X1 U2394 ( .A1(n3824), .A2(n4182), .ZN(n3921) );
  OAI21_X1 U2395 ( .B1(n2509), .B2(n2064), .A(n2529), .ZN(n2063) );
  NAND2_X1 U2396 ( .A1(n2213), .A2(n2035), .ZN(n3184) );
  NAND2_X1 U2397 ( .A1(n2242), .A2(n2240), .ZN(n2754) );
  AOI21_X1 U2398 ( .B1(n2243), .B2(n2245), .A(n2241), .ZN(n2240) );
  INV_X1 U2399 ( .A(n3912), .ZN(n2241) );
  AND2_X1 U2400 ( .A1(n4308), .A2(n4329), .ZN(n2256) );
  NAND2_X1 U2401 ( .A1(n3403), .A2(n3929), .ZN(n2252) );
  NAND2_X1 U2402 ( .A1(n2252), .A2(n2250), .ZN(n4359) );
  NOR2_X1 U2403 ( .A1(n4357), .A2(n2251), .ZN(n2250) );
  INV_X1 U2404 ( .A(n3891), .ZN(n2251) );
  NAND2_X1 U2405 ( .A1(n2363), .A2(n2057), .ZN(n3028) );
  INV_X1 U2406 ( .A(n2645), .ZN(n2642) );
  OR2_X1 U2407 ( .A1(n2439), .A2(IR_REG_10__SCAN_IN), .ZN(n2461) );
  INV_X1 U2408 ( .A(IR_REG_6__SCAN_IN), .ZN(n2422) );
  NAND2_X1 U2409 ( .A1(n2232), .A2(IR_REG_31__SCAN_IN), .ZN(n2186) );
  INV_X1 U2410 ( .A(n2148), .ZN(n2555) );
  AND2_X1 U2411 ( .A1(n3642), .A2(n2293), .ZN(n2292) );
  INV_X1 U2412 ( .A(n3820), .ZN(n2293) );
  INV_X1 U2413 ( .A(n2295), .ZN(n2294) );
  OAI21_X1 U2414 ( .B1(n3820), .B2(n2296), .A(n3818), .ZN(n2295) );
  NAND2_X1 U2415 ( .A1(n3799), .A2(n3798), .ZN(n2280) );
  NAND2_X1 U2416 ( .A1(n2283), .A2(n2282), .ZN(n2281) );
  INV_X1 U2417 ( .A(n3798), .ZN(n2282) );
  INV_X1 U2418 ( .A(n3799), .ZN(n2283) );
  OR2_X1 U2419 ( .A1(n2416), .A2(n3107), .ZN(n2429) );
  NAND2_X1 U2420 ( .A1(n3572), .A2(n3571), .ZN(n3573) );
  INV_X1 U2421 ( .A(n3569), .ZN(n3572) );
  NAND2_X1 U2422 ( .A1(n2142), .A2(REG3_REG_10__SCAN_IN), .ZN(n2441) );
  XNOR2_X1 U2423 ( .A(n2966), .B(n3658), .ZN(n3129) );
  OR2_X1 U2424 ( .A1(n3552), .A2(n3068), .ZN(n2963) );
  OR2_X1 U2425 ( .A1(n2021), .A2(n3560), .ZN(n2270) );
  NOR2_X1 U2426 ( .A1(n2021), .A2(n2272), .ZN(n2271) );
  INV_X1 U2427 ( .A(n3553), .ZN(n2272) );
  NAND2_X1 U2428 ( .A1(n3690), .A2(n3539), .ZN(n3545) );
  OR2_X1 U2429 ( .A1(n2480), .A2(n4608), .ZN(n2492) );
  NAND2_X1 U2430 ( .A1(n2491), .A2(REG3_REG_15__SCAN_IN), .ZN(n2501) );
  OAI21_X1 U2431 ( .B1(n3994), .B2(n2139), .A(n2136), .ZN(n2135) );
  AND2_X1 U2432 ( .A1(n3995), .A2(n4120), .ZN(n2139) );
  AND2_X1 U2433 ( .A1(n2138), .A2(n2137), .ZN(n2136) );
  AND2_X1 U2434 ( .A1(n3174), .A2(n2954), .ZN(n4003) );
  INV_X1 U2435 ( .A(n2355), .ZN(n2614) );
  OR2_X1 U2436 ( .A1(n2355), .A2(n2935), .ZN(n2659) );
  INV_X1 U2437 ( .A(n4695), .ZN(n2901) );
  NAND2_X1 U2438 ( .A1(n2100), .A2(n2105), .ZN(n2103) );
  AOI21_X1 U2439 ( .B1(n2173), .B2(n2025), .A(n2172), .ZN(n2174) );
  NAND2_X1 U2440 ( .A1(n2199), .A2(REG2_REG_8__SCAN_IN), .ZN(n2198) );
  AND2_X1 U2441 ( .A1(n2104), .A2(n2011), .ZN(n3104) );
  INV_X1 U2442 ( .A(n3379), .ZN(n2093) );
  XNOR2_X1 U2443 ( .A(n3379), .B(n4691), .ZN(n3380) );
  NAND2_X1 U2444 ( .A1(n2166), .A2(n2165), .ZN(n2164) );
  NAND2_X1 U2445 ( .A1(n4081), .A2(REG1_REG_14__SCAN_IN), .ZN(n2166) );
  NAND2_X1 U2446 ( .A1(n2181), .A2(n2179), .ZN(n4094) );
  AOI21_X1 U2447 ( .B1(n3488), .B2(n4082), .A(n2180), .ZN(n2179) );
  INV_X1 U2448 ( .A(n4095), .ZN(n2180) );
  INV_X1 U2449 ( .A(n3469), .ZN(n3470) );
  NAND2_X1 U2450 ( .A1(n4714), .A2(n2050), .ZN(n2171) );
  NAND2_X1 U2451 ( .A1(n4709), .A2(n2098), .ZN(n4721) );
  NAND2_X1 U2452 ( .A1(n4773), .A2(n2516), .ZN(n2098) );
  NOR2_X1 U2453 ( .A1(n4721), .A2(n4720), .ZN(n4718) );
  OR2_X1 U2454 ( .A1(n2622), .A2(n2621), .ZN(n2793) );
  NAND2_X1 U2455 ( .A1(n2073), .A2(n2597), .ZN(n4176) );
  NAND2_X1 U2456 ( .A1(n2590), .A2(n2022), .ZN(n2073) );
  NAND2_X1 U2457 ( .A1(n2202), .A2(n2203), .ZN(n4203) );
  AOI21_X1 U2458 ( .B1(n2005), .B2(n2571), .A(n2015), .ZN(n2203) );
  NAND2_X1 U2459 ( .A1(n2205), .A2(n2206), .ZN(n2204) );
  INV_X1 U2460 ( .A(n4250), .ZN(n2205) );
  NAND2_X1 U2461 ( .A1(n2230), .A2(n3977), .ZN(n4248) );
  NAND2_X1 U2462 ( .A1(n2215), .A2(n2214), .ZN(n4261) );
  AOI21_X1 U2463 ( .B1(n2216), .B2(n2218), .A(n2030), .ZN(n2214) );
  NAND2_X1 U2464 ( .A1(n4305), .A2(n2216), .ZN(n2215) );
  NAND2_X1 U2465 ( .A1(n2530), .A2(REG3_REG_18__SCAN_IN), .ZN(n2544) );
  INV_X1 U2466 ( .A(n2532), .ZN(n2530) );
  NAND2_X1 U2467 ( .A1(n4352), .A2(n2509), .ZN(n4351) );
  NAND2_X1 U2468 ( .A1(n4359), .A2(n3879), .ZN(n4341) );
  NAND2_X1 U2469 ( .A1(n4341), .A2(n4340), .ZN(n4339) );
  INV_X1 U2470 ( .A(n2067), .ZN(n2066) );
  OAI21_X1 U2471 ( .B1(n2068), .B2(n2210), .A(n2207), .ZN(n2067) );
  AOI21_X1 U2472 ( .B1(n2209), .B2(n2208), .A(n2027), .ZN(n2207) );
  INV_X1 U2473 ( .A(n3449), .ZN(n2212) );
  OR2_X1 U2474 ( .A1(n2469), .A2(n2468), .ZN(n2480) );
  AND2_X1 U2475 ( .A1(n3876), .A2(n2042), .ZN(n2239) );
  NOR2_X1 U2476 ( .A1(n2248), .A2(n2247), .ZN(n2246) );
  INV_X1 U2477 ( .A(n2664), .ZN(n2247) );
  NAND2_X1 U2478 ( .A1(n2377), .A2(n2036), .ZN(n2399) );
  NAND2_X1 U2479 ( .A1(n4023), .A2(n3150), .ZN(n3860) );
  NAND2_X1 U2480 ( .A1(n3063), .A2(n2008), .ZN(n2113) );
  NOR2_X1 U2481 ( .A1(n2070), .A2(n2071), .ZN(n3249) );
  OAI21_X1 U2482 ( .B1(n2353), .B2(n3154), .A(n2072), .ZN(n2071) );
  NAND2_X1 U2483 ( .A1(n3860), .A2(n3857), .ZN(n3040) );
  INV_X1 U2484 ( .A(n2663), .ZN(n3933) );
  NAND2_X1 U2485 ( .A1(n2127), .A2(n2318), .ZN(n2347) );
  NAND2_X1 U2486 ( .A1(n2812), .A2(n2811), .ZN(n2814) );
  INV_X1 U2487 ( .A(n3936), .ZN(n2812) );
  INV_X1 U2488 ( .A(n2982), .ZN(n2986) );
  XNOR2_X1 U2489 ( .A(n4143), .B(n2779), .ZN(n3966) );
  NAND2_X1 U2490 ( .A1(n4239), .A2(n2017), .ZN(n4194) );
  NOR2_X2 U2491 ( .A1(n4295), .A2(n4420), .ZN(n4272) );
  INV_X1 U2492 ( .A(n3806), .ZN(n3427) );
  NAND2_X1 U2493 ( .A1(n2683), .A2(n2682), .ZN(n4338) );
  INV_X1 U2494 ( .A(n4338), .ZN(n4475) );
  AND2_X1 U2495 ( .A1(n2725), .A2(n2724), .ZN(n2951) );
  NAND3_X1 U2496 ( .A1(n2322), .A2(n2308), .A3(n2261), .ZN(n2056) );
  INV_X1 U2497 ( .A(IR_REG_21__SCAN_IN), .ZN(n2646) );
  AND2_X1 U2498 ( .A1(n2485), .A2(IR_REG_31__SCAN_IN), .ZN(n2486) );
  NAND2_X1 U2499 ( .A1(n2488), .A2(n2487), .ZN(n2497) );
  INV_X1 U2500 ( .A(IR_REG_15__SCAN_IN), .ZN(n2487) );
  INV_X1 U2501 ( .A(n2486), .ZN(n2488) );
  INV_X1 U2502 ( .A(IR_REG_11__SCAN_IN), .ZN(n2520) );
  OR2_X1 U2503 ( .A1(n3129), .A2(n3128), .ZN(n3130) );
  INV_X1 U2504 ( .A(n3620), .ZN(n3621) );
  NAND2_X1 U2505 ( .A1(n2079), .A2(n2076), .ZN(n3622) );
  INV_X1 U2506 ( .A(n2743), .ZN(n3827) );
  AND2_X1 U2507 ( .A1(n2628), .A2(n2608), .ZN(n4163) );
  INV_X1 U2508 ( .A(n4155), .ZN(n4014) );
  NAND2_X1 U2509 ( .A1(n2596), .A2(n2595), .ZN(n4016) );
  NAND2_X1 U2510 ( .A1(n2569), .A2(n2568), .ZN(n4230) );
  NAND2_X1 U2511 ( .A1(n2508), .A2(n2507), .ZN(n4456) );
  INV_X1 U2512 ( .A(n3702), .ZN(n4487) );
  INV_X1 U2513 ( .A(n3341), .ZN(n4019) );
  INV_X1 U2514 ( .A(n3160), .ZN(n4022) );
  INV_X1 U2515 ( .A(n3249), .ZN(n4023) );
  NAND2_X1 U2516 ( .A1(n2125), .A2(n2124), .ZN(n2123) );
  XNOR2_X1 U2517 ( .A(n2902), .B(n2901), .ZN(n4042) );
  XNOR2_X1 U2518 ( .A(n2917), .B(n2896), .ZN(n2919) );
  INV_X1 U2519 ( .A(n4694), .ZN(n2896) );
  INV_X1 U2520 ( .A(IR_REG_8__SCAN_IN), .ZN(n2408) );
  INV_X1 U2521 ( .A(n4690), .ZN(n2155) );
  AOI22_X1 U2522 ( .A1(n4060), .A2(REG2_REG_12__SCAN_IN), .B1(n4690), .B2(
        n3484), .ZN(n4070) );
  NAND2_X1 U2523 ( .A1(n2182), .A2(REG2_REG_14__SCAN_IN), .ZN(n4088) );
  INV_X1 U2524 ( .A(n4083), .ZN(n2182) );
  XNOR2_X1 U2525 ( .A(n2739), .B(n3965), .ZN(n4162) );
  OAI21_X1 U2526 ( .B1(n2590), .B2(n2227), .A(n2225), .ZN(n2739) );
  AND2_X1 U2527 ( .A1(n2226), .A2(n2738), .ZN(n2225) );
  OR2_X1 U2528 ( .A1(n2227), .A2(n2022), .ZN(n2226) );
  OR2_X1 U2529 ( .A1(n4745), .A2(n2824), .ZN(n4364) );
  OR2_X1 U2530 ( .A1(n4745), .A2(n3221), .ZN(n4378) );
  AOI21_X1 U2531 ( .B1(n4135), .B2(n4480), .A(n2694), .ZN(n2736) );
  AND2_X1 U2532 ( .A1(n4161), .A2(n2131), .ZN(n2804) );
  AOI21_X1 U2533 ( .B1(n4150), .B2(n4480), .A(n2132), .ZN(n2131) );
  OAI21_X1 U2534 ( .B1(n4155), .B2(n4439), .A(n2798), .ZN(n2132) );
  INV_X2 U2535 ( .A(n4782), .ZN(n4783) );
  OR2_X1 U2536 ( .A1(n2732), .A2(n2951), .ZN(n4782) );
  INV_X1 U2537 ( .A(n3211), .ZN(n2194) );
  NAND2_X1 U2538 ( .A1(n2918), .A2(n2102), .ZN(n2099) );
  AND2_X1 U2539 ( .A1(n2040), .A2(n2011), .ZN(n2101) );
  NOR2_X1 U2540 ( .A1(n4092), .A2(n2162), .ZN(n2161) );
  INV_X1 U2541 ( .A(REG1_REG_14__SCAN_IN), .ZN(n2162) );
  NAND2_X1 U2542 ( .A1(n2333), .A2(n2975), .ZN(n3848) );
  INV_X1 U2543 ( .A(n3911), .ZN(n2245) );
  INV_X1 U2544 ( .A(n2244), .ZN(n2243) );
  OAI21_X1 U2545 ( .B1(n3970), .B2(n2245), .A(n3905), .ZN(n2244) );
  AND2_X1 U2546 ( .A1(n2673), .A2(n3871), .ZN(n2253) );
  INV_X1 U2547 ( .A(n2429), .ZN(n2142) );
  AOI21_X1 U2548 ( .B1(n2278), .B2(n2275), .A(n2274), .ZN(n2273) );
  INV_X1 U2549 ( .A(n3734), .ZN(n2274) );
  INV_X1 U2550 ( .A(n2281), .ZN(n2275) );
  NAND2_X1 U2551 ( .A1(n3997), .A2(n3998), .ZN(n2138) );
  NOR2_X1 U2552 ( .A1(n3996), .A2(n2705), .ZN(n2137) );
  OR2_X1 U2553 ( .A1(n2953), .A2(n4004), .ZN(n2965) );
  OAI21_X1 U2554 ( .B1(n4693), .B2(REG1_REG_7__SCAN_IN), .A(
        REG1_REG_6__SCAN_IN), .ZN(n2177) );
  INV_X1 U2555 ( .A(n2913), .ZN(n2173) );
  NOR2_X1 U2556 ( .A1(n2175), .A2(n2178), .ZN(n2172) );
  INV_X1 U2557 ( .A(n4691), .ZN(n2091) );
  NOR2_X1 U2558 ( .A1(n2544), .A2(n2543), .ZN(n2148) );
  INV_X1 U2559 ( .A(n2542), .ZN(n2218) );
  NOR2_X1 U2560 ( .A1(n2146), .A2(n2145), .ZN(n2144) );
  INV_X1 U2561 ( .A(n2492), .ZN(n2491) );
  INV_X1 U2562 ( .A(n2302), .ZN(n2208) );
  AOI21_X1 U2563 ( .B1(n2220), .B2(n2012), .A(n2034), .ZN(n2068) );
  INV_X1 U2564 ( .A(n2447), .ZN(n2219) );
  AOI21_X1 U2565 ( .B1(n2236), .B2(n2238), .A(n2234), .ZN(n2233) );
  NAND2_X1 U2566 ( .A1(n2236), .A2(n2120), .ZN(n2119) );
  INV_X1 U2567 ( .A(n3883), .ZN(n2234) );
  INV_X1 U2568 ( .A(n2236), .ZN(n2121) );
  INV_X1 U2569 ( .A(n2224), .ZN(n2221) );
  AND2_X1 U2570 ( .A1(n3183), .A2(n2413), .ZN(n2411) );
  INV_X1 U2571 ( .A(n3861), .ZN(n2248) );
  INV_X1 U2572 ( .A(n2379), .ZN(n2377) );
  NAND3_X1 U2573 ( .A1(n2112), .A2(n2111), .A3(n3875), .ZN(n2249) );
  NAND2_X1 U2574 ( .A1(n2114), .A2(n2023), .ZN(n2111) );
  INV_X1 U2575 ( .A(n3860), .ZN(n2116) );
  NOR2_X1 U2576 ( .A1(n2327), .A2(IR_REG_5__SCAN_IN), .ZN(n2260) );
  NAND2_X1 U2577 ( .A1(n2973), .A2(n3011), .ZN(n3850) );
  NOR2_X1 U2578 ( .A1(n2802), .A2(n3670), .ZN(n2778) );
  NOR2_X1 U2579 ( .A1(n4229), .A2(n4210), .ZN(n2258) );
  NAND2_X1 U2580 ( .A1(n3271), .A2(n2257), .ZN(n3355) );
  AND2_X1 U2581 ( .A1(n2010), .A2(n4490), .ZN(n2257) );
  AND2_X1 U2582 ( .A1(n2847), .A2(n4687), .ZN(n2955) );
  AND2_X1 U2583 ( .A1(n2638), .A2(IR_REG_31__SCAN_IN), .ZN(n2639) );
  INV_X1 U2584 ( .A(IR_REG_17__SCAN_IN), .ZN(n2539) );
  INV_X1 U2585 ( .A(n2435), .ZN(n2436) );
  AOI21_X1 U2586 ( .B1(n2287), .B2(n3233), .A(n2289), .ZN(n2286) );
  NAND2_X1 U2587 ( .A1(n2299), .A2(n3236), .ZN(n2287) );
  OR2_X1 U2588 ( .A1(n3530), .A2(n3529), .ZN(n3734) );
  AND2_X1 U2589 ( .A1(n2078), .A2(n2077), .ZN(n2076) );
  NAND2_X1 U2590 ( .A1(n2081), .A2(n3633), .ZN(n2077) );
  NAND2_X1 U2591 ( .A1(n2083), .A2(n2085), .ZN(n2078) );
  NAND2_X1 U2592 ( .A1(n2491), .A2(n2144), .ZN(n2511) );
  INV_X1 U2593 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3107) );
  NOR2_X1 U2594 ( .A1(n2928), .A2(n3552), .ZN(n2074) );
  CLKBUF_X1 U2595 ( .A(n3690), .Z(n3691) );
  NAND2_X1 U2596 ( .A1(n3775), .A2(n2088), .ZN(n2290) );
  AND2_X1 U2597 ( .A1(n2044), .A2(n3779), .ZN(n2088) );
  NAND2_X1 U2598 ( .A1(n2142), .A2(n2140), .ZN(n2453) );
  NOR2_X1 U2599 ( .A1(n3383), .A2(n2141), .ZN(n2140) );
  INV_X1 U2600 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3383) );
  NOR2_X1 U2601 ( .A1(n2628), .A2(n2626), .ZN(n2686) );
  OR2_X1 U2602 ( .A1(n2353), .A2(n2999), .ZN(n2660) );
  NAND2_X1 U2603 ( .A1(n2189), .A2(n2871), .ZN(n2188) );
  OAI211_X1 U2604 ( .C1(n2186), .C2(n2231), .A(n2014), .B(n2185), .ZN(n2187)
         );
  INV_X1 U2605 ( .A(n2191), .ZN(n2189) );
  INV_X1 U2606 ( .A(n4696), .ZN(n2884) );
  OR2_X1 U2607 ( .A1(n2907), .A2(n2376), .ZN(n2914) );
  NAND2_X1 U2608 ( .A1(n3376), .A2(n2154), .ZN(n2150) );
  NOR2_X1 U2609 ( .A1(n3377), .A2(n4673), .ZN(n2154) );
  NAND2_X1 U2610 ( .A1(n2149), .A2(n2152), .ZN(n2151) );
  INV_X1 U2611 ( .A(n3377), .ZN(n2152) );
  INV_X1 U2612 ( .A(n2157), .ZN(n2149) );
  AND2_X1 U2613 ( .A1(n2096), .A2(n2095), .ZN(n3483) );
  NAND2_X1 U2614 ( .A1(n3482), .A2(REG2_REG_11__SCAN_IN), .ZN(n2095) );
  XNOR2_X1 U2615 ( .A(n3486), .B(n4086), .ZN(n4083) );
  NAND2_X1 U2616 ( .A1(n3493), .A2(n3492), .ZN(n4710) );
  INV_X1 U2617 ( .A(n2589), .ZN(n2229) );
  OR2_X1 U2618 ( .A1(n2737), .A2(n2228), .ZN(n2227) );
  INV_X1 U2619 ( .A(n2597), .ZN(n2228) );
  NAND2_X1 U2620 ( .A1(n2491), .A2(n2143), .ZN(n2532) );
  AND2_X1 U2621 ( .A1(n2144), .A2(REG3_REG_17__SCAN_IN), .ZN(n2143) );
  NAND2_X1 U2622 ( .A1(n2510), .A2(n2065), .ZN(n2061) );
  INV_X1 U2623 ( .A(n2063), .ZN(n2062) );
  NAND2_X1 U2624 ( .A1(n4305), .A2(n4304), .ZN(n4303) );
  NAND2_X1 U2625 ( .A1(n2451), .A2(REG3_REG_12__SCAN_IN), .ZN(n2469) );
  INV_X1 U2626 ( .A(n2453), .ZN(n2451) );
  OR2_X1 U2627 ( .A1(n2223), .A2(n2006), .ZN(n3416) );
  NAND2_X1 U2628 ( .A1(n2377), .A2(REG3_REG_6__SCAN_IN), .ZN(n2388) );
  NAND2_X1 U2629 ( .A1(n2249), .A2(n3861), .ZN(n3202) );
  NAND2_X1 U2630 ( .A1(n2956), .A2(n2728), .ZN(n3200) );
  AND2_X1 U2631 ( .A1(n2109), .A2(n3873), .ZN(n2114) );
  NAND2_X1 U2632 ( .A1(n2115), .A2(n2110), .ZN(n2109) );
  NOR2_X1 U2633 ( .A1(n2008), .A2(n2116), .ZN(n2115) );
  AND2_X1 U2634 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2364) );
  NAND2_X1 U2635 ( .A1(n2364), .A2(REG3_REG_5__SCAN_IN), .ZN(n2379) );
  NAND2_X1 U2636 ( .A1(n3063), .A2(n3856), .ZN(n3041) );
  NAND2_X1 U2637 ( .A1(n3936), .A2(n2662), .ZN(n2809) );
  NOR2_X1 U2638 ( .A1(n4119), .A2(n4120), .ZN(n4118) );
  NAND2_X1 U2639 ( .A1(n4239), .A2(n2258), .ZN(n4214) );
  NAND2_X1 U2640 ( .A1(n4239), .A2(n4241), .ZN(n4240) );
  NAND2_X1 U2641 ( .A1(n4342), .A2(n2046), .ZN(n4295) );
  NAND2_X1 U2642 ( .A1(n4342), .A2(n2256), .ZN(n4307) );
  INV_X1 U2643 ( .A(n4436), .ZN(n4329) );
  AND2_X1 U2644 ( .A1(n4342), .A2(n4329), .ZN(n4328) );
  AND2_X1 U2645 ( .A1(n2538), .A2(n2537), .ZN(n4440) );
  INV_X1 U2646 ( .A(n4459), .ZN(n4361) );
  NAND2_X1 U2647 ( .A1(n2252), .A2(n3891), .ZN(n4358) );
  NOR2_X1 U2648 ( .A1(n3355), .A2(n3534), .ZN(n3450) );
  NAND2_X1 U2649 ( .A1(n3271), .A2(n2010), .ZN(n3425) );
  AND2_X1 U2650 ( .A1(n3271), .A2(n3342), .ZN(n3311) );
  NAND2_X1 U2651 ( .A1(n3271), .A2(n2009), .ZN(n3424) );
  OR2_X1 U2652 ( .A1(n3201), .A2(n3204), .ZN(n3198) );
  AND2_X1 U2653 ( .A1(n3220), .A2(n3070), .ZN(n4497) );
  NAND2_X1 U2654 ( .A1(n3099), .A2(n3177), .ZN(n3201) );
  NOR2_X1 U2655 ( .A1(n3075), .A2(n3042), .ZN(n3049) );
  AND2_X1 U2656 ( .A1(n3049), .A2(n3246), .ZN(n3099) );
  NAND2_X1 U2657 ( .A1(n2255), .A2(n2254), .ZN(n3075) );
  INV_X1 U2658 ( .A(n3074), .ZN(n2255) );
  NOR2_X1 U2659 ( .A1(n3073), .A2(n3072), .ZN(n2254) );
  AND2_X1 U2660 ( .A1(n2955), .A2(n2989), .ZN(n4485) );
  INV_X1 U2661 ( .A(n4489), .ZN(n4437) );
  AND2_X1 U2662 ( .A1(n4750), .A2(n4004), .ZN(n4776) );
  NAND2_X1 U2663 ( .A1(n2702), .A2(n2698), .ZN(n2755) );
  NAND2_X1 U2664 ( .A1(n2701), .A2(IR_REG_31__SCAN_IN), .ZN(n2699) );
  OR2_X1 U2665 ( .A1(n2465), .A2(IR_REG_13__SCAN_IN), .ZN(n2477) );
  AND2_X1 U2666 ( .A1(n2435), .A2(n2261), .ZN(n2425) );
  OR2_X1 U2667 ( .A1(n2395), .A2(n2637), .ZN(n2406) );
  NAND2_X1 U2668 ( .A1(n2637), .A2(IR_REG_1__SCAN_IN), .ZN(n2191) );
  OAI21_X1 U2669 ( .B1(IR_REG_0__SCAN_IN), .B2(IR_REG_1__SCAN_IN), .A(n2184), 
        .ZN(n2190) );
  NAND2_X1 U2670 ( .A1(n2186), .A2(IR_REG_0__SCAN_IN), .ZN(n2184) );
  XNOR2_X1 U2671 ( .A(n2628), .B(REG3_REG_27__SCAN_IN), .ZN(n4152) );
  AOI21_X1 U2672 ( .B1(n2266), .B2(n2269), .A(n2264), .ZN(n2263) );
  INV_X1 U2673 ( .A(n3810), .ZN(n2264) );
  AND2_X1 U2674 ( .A1(n3674), .A2(n3668), .ZN(n3669) );
  NAND2_X1 U2675 ( .A1(n2291), .A2(n2031), .ZN(n3681) );
  OR2_X1 U2676 ( .A1(n3797), .A2(n2277), .ZN(n2276) );
  INV_X1 U2677 ( .A(n2280), .ZN(n2277) );
  NAND2_X1 U2678 ( .A1(n3164), .A2(n3163), .ZN(n3172) );
  INV_X1 U2679 ( .A(n4021), .ZN(n3248) );
  AND2_X1 U2680 ( .A1(n2587), .A2(n2586), .ZN(n4233) );
  OR2_X1 U2681 ( .A1(n4217), .A2(n2353), .ZN(n2587) );
  NAND2_X1 U2682 ( .A1(n3710), .A2(n3614), .ZN(n3766) );
  NAND2_X1 U2683 ( .A1(n2075), .A2(n2083), .ZN(n3767) );
  AND4_X1 U2684 ( .A1(n2404), .A2(n2403), .A3(n2402), .A4(n2401), .ZN(n3341)
         );
  AND3_X1 U2685 ( .A1(n2484), .A2(n2483), .A3(n2482), .ZN(n4368) );
  NAND2_X1 U2686 ( .A1(n2290), .A2(n3589), .ZN(n3591) );
  INV_X1 U2687 ( .A(n4017), .ZN(n3802) );
  AND2_X1 U2688 ( .A1(n2977), .A2(n2978), .ZN(n2979) );
  INV_X1 U2689 ( .A(n3128), .ZN(n2968) );
  INV_X1 U2690 ( .A(n4311), .ZN(n4308) );
  NAND2_X1 U2691 ( .A1(n3746), .A2(n2271), .ZN(n2265) );
  INV_X1 U2692 ( .A(n3301), .ZN(n3177) );
  NAND2_X1 U2693 ( .A1(n3127), .A2(n3126), .ZN(n3829) );
  INV_X1 U2694 ( .A(n3783), .ZN(n3843) );
  INV_X1 U2695 ( .A(n3829), .ZN(n3846) );
  NAND2_X1 U2696 ( .A1(n2135), .A2(n2134), .ZN(n2133) );
  NAND2_X1 U2697 ( .A1(n3999), .A2(n2705), .ZN(n2134) );
  NAND2_X1 U2698 ( .A1(n2613), .A2(n2612), .ZN(n4383) );
  NAND2_X1 U2699 ( .A1(n2606), .A2(n2605), .ZN(n3824) );
  OR2_X1 U2700 ( .A1(n3624), .A2(n2353), .ZN(n2606) );
  INV_X1 U2701 ( .A(n4233), .ZN(n4393) );
  NAND2_X1 U2702 ( .A1(n2561), .A2(n2560), .ZN(n4411) );
  OR2_X1 U2703 ( .A1(n3781), .A2(n2353), .ZN(n2561) );
  NAND2_X1 U2704 ( .A1(n2550), .A2(n2549), .ZN(n4421) );
  INV_X1 U2705 ( .A(n4440), .ZN(n4289) );
  INV_X1 U2706 ( .A(n3751), .ZN(n4447) );
  OAI211_X1 U2707 ( .C1(n3510), .C2(n3489), .A(n2495), .B(n2494), .ZN(n4467)
         );
  NAND4_X1 U2708 ( .A1(n2434), .A2(n2433), .A3(n2432), .A4(n2431), .ZN(n3806)
         );
  NAND2_X1 U2709 ( .A1(n4054), .A2(n4055), .ZN(n4053) );
  INV_X1 U2710 ( .A(n2103), .ZN(n2921) );
  XNOR2_X1 U2711 ( .A(n3104), .B(n3110), .ZN(n3106) );
  NAND2_X1 U2712 ( .A1(n3104), .A2(n2198), .ZN(n2195) );
  NAND2_X1 U2713 ( .A1(n2151), .A2(n2150), .ZN(n3465) );
  AND2_X1 U2714 ( .A1(n2153), .A2(n2157), .ZN(n3378) );
  NAND2_X1 U2715 ( .A1(n3376), .A2(REG1_REG_10__SCAN_IN), .ZN(n2153) );
  AND2_X1 U2716 ( .A1(n2094), .A2(n2097), .ZN(n3382) );
  NAND2_X1 U2717 ( .A1(n3380), .A2(REG2_REG_10__SCAN_IN), .ZN(n2094) );
  INV_X1 U2718 ( .A(n4092), .ZN(n2163) );
  INV_X1 U2719 ( .A(n2164), .ZN(n4093) );
  NAND2_X1 U2720 ( .A1(n4088), .A2(n3488), .ZN(n4096) );
  NAND2_X1 U2721 ( .A1(n4710), .A2(n4711), .ZN(n4709) );
  OR2_X1 U2722 ( .A1(n4710), .A2(n4711), .ZN(n2201) );
  OAI22_X1 U2723 ( .A1(n4104), .A2(n2170), .B1(n2171), .B2(n2169), .ZN(n2168)
         );
  INV_X1 U2724 ( .A(n4732), .ZN(n2169) );
  NAND2_X1 U2725 ( .A1(n3473), .A2(n2051), .ZN(n2170) );
  OAI21_X1 U2726 ( .B1(n4104), .B2(n2167), .A(n2171), .ZN(n4731) );
  NAND2_X1 U2727 ( .A1(n3473), .A2(n2050), .ZN(n2167) );
  INV_X1 U2728 ( .A(n4114), .ZN(n4730) );
  INV_X1 U2729 ( .A(n4718), .ZN(n4728) );
  OR2_X1 U2730 ( .A1(n4708), .A2(n4705), .ZN(n4114) );
  OR2_X1 U2731 ( .A1(n4708), .A2(n2989), .ZN(n4735) );
  NOR2_X1 U2732 ( .A1(n4718), .A2(n3497), .ZN(n3499) );
  AND2_X1 U2733 ( .A1(n3496), .A2(REG2_REG_18__SCAN_IN), .ZN(n3497) );
  AND2_X1 U2734 ( .A1(n2634), .A2(n2633), .ZN(n4155) );
  OR2_X1 U2735 ( .A1(n4138), .A2(n2353), .ZN(n2634) );
  OAI21_X1 U2736 ( .B1(n4176), .B2(n2792), .A(n2793), .ZN(n2794) );
  OR2_X1 U2737 ( .A1(n4172), .A2(n4171), .ZN(n4173) );
  INV_X1 U2738 ( .A(n4383), .ZN(n4183) );
  INV_X1 U2739 ( .A(n2128), .ZN(n4189) );
  NAND2_X1 U2740 ( .A1(n2204), .A2(n2005), .ZN(n4236) );
  NAND2_X1 U2741 ( .A1(n2204), .A2(n2570), .ZN(n4238) );
  AND2_X1 U2742 ( .A1(n2579), .A2(n2578), .ZN(n4414) );
  OR2_X1 U2743 ( .A1(n4242), .A2(n2353), .ZN(n2579) );
  INV_X1 U2744 ( .A(n4410), .ZN(n4255) );
  NAND2_X1 U2745 ( .A1(n4351), .A2(n2510), .ZN(n4326) );
  NAND2_X1 U2746 ( .A1(n4339), .A2(n3871), .ZN(n4322) );
  INV_X1 U2747 ( .A(n4467), .ZN(n4350) );
  NAND2_X1 U2748 ( .A1(n2211), .A2(n2209), .ZN(n3404) );
  NAND2_X1 U2749 ( .A1(n2212), .A2(n2302), .ZN(n2211) );
  AND3_X1 U2750 ( .A1(n2475), .A2(n2474), .A3(n2473), .ZN(n3702) );
  INV_X1 U2751 ( .A(n4484), .ZN(n3739) );
  INV_X1 U2752 ( .A(n2667), .ZN(n3397) );
  NAND2_X1 U2753 ( .A1(n2235), .A2(n3865), .ZN(n3309) );
  NAND2_X1 U2754 ( .A1(n2666), .A2(n2239), .ZN(n2235) );
  INV_X1 U2755 ( .A(n3266), .ZN(n3342) );
  NAND2_X1 U2756 ( .A1(n2666), .A2(n3876), .ZN(n3268) );
  NAND4_X1 U2757 ( .A1(n2421), .A2(n2420), .A3(n2419), .A4(n2418), .ZN(n4018)
         );
  OR2_X1 U2758 ( .A1(n3510), .A2(n3325), .ZN(n2418) );
  AND2_X1 U2759 ( .A1(n2213), .A2(n2024), .ZN(n3095) );
  AND4_X1 U2760 ( .A1(n2394), .A2(n2393), .A3(n2392), .A4(n2391), .ZN(n3304)
         );
  NAND2_X1 U2761 ( .A1(n2113), .A2(n3860), .ZN(n3026) );
  INV_X1 U2762 ( .A(n4755), .ZN(n4737) );
  INV_X1 U2763 ( .A(n3073), .ZN(n2967) );
  NAND2_X1 U2764 ( .A1(n2814), .A2(n2337), .ZN(n2830) );
  OR2_X1 U2765 ( .A1(n4745), .A2(n4439), .ZN(n4371) );
  OR2_X1 U2766 ( .A1(n4745), .A2(n4489), .ZN(n4370) );
  AND2_X1 U2767 ( .A1(n4127), .A2(n2777), .ZN(n2787) );
  OAI21_X1 U2768 ( .B1(n4179), .B2(n4182), .A(n4178), .ZN(n4505) );
  NAND2_X1 U2769 ( .A1(n2818), .A2(n2982), .ZN(n4767) );
  AND2_X1 U2770 ( .A1(n2284), .A2(n2285), .ZN(n2108) );
  NAND2_X1 U2771 ( .A1(n2055), .A2(IR_REG_31__SCAN_IN), .ZN(n2086) );
  INV_X1 U2772 ( .A(n4316), .ZN(n3501) );
  NAND2_X1 U2773 ( .A1(n2489), .A2(n2497), .ZN(n4100) );
  XNOR2_X1 U2774 ( .A(n2450), .B(IR_REG_12__SCAN_IN), .ZN(n4690) );
  XNOR2_X1 U2775 ( .A(n2386), .B(IR_REG_6__SCAN_IN), .ZN(n4694) );
  XNOR2_X1 U2776 ( .A(n2373), .B(n2261), .ZN(n4047) );
  XNOR2_X1 U2777 ( .A(n2361), .B(IR_REG_4__SCAN_IN), .ZN(n4695) );
  OAI21_X1 U2778 ( .B1(IR_REG_0__SCAN_IN), .B2(IR_REG_1__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2106) );
  AOI21_X1 U2779 ( .B1(n4147), .B2(n4752), .A(n4146), .ZN(n4148) );
  AND2_X1 U2780 ( .A1(n2734), .A2(n2733), .ZN(n2735) );
  OAI21_X1 U2781 ( .B1(n2804), .B2(n4784), .A(n2016), .ZN(U3545) );
  OR2_X1 U2782 ( .A1(n4151), .A2(n4483), .ZN(n2803) );
  OR2_X1 U2783 ( .A1(n4165), .A2(n4483), .ZN(n2748) );
  AND2_X1 U2784 ( .A1(n2730), .A2(n2729), .ZN(n2731) );
  OR2_X1 U2785 ( .A1(n4151), .A2(n4546), .ZN(n2806) );
  OR2_X1 U2786 ( .A1(n4165), .A2(n4546), .ZN(n2751) );
  AND2_X1 U2787 ( .A1(n2580), .A2(n2570), .ZN(n2005) );
  INV_X1 U2788 ( .A(n3072), .ZN(n3135) );
  OR2_X1 U2789 ( .A1(n3417), .A2(n2221), .ZN(n2006) );
  XNOR2_X1 U2790 ( .A(n2409), .B(n2408), .ZN(n3110) );
  INV_X1 U2791 ( .A(n3110), .ZN(n2199) );
  AND2_X1 U2792 ( .A1(n2233), .A2(n2119), .ZN(n2007) );
  AND2_X1 U2793 ( .A1(n3856), .A2(n3857), .ZN(n2008) );
  AND2_X1 U2794 ( .A1(n3342), .A2(n3397), .ZN(n2009) );
  AND2_X1 U2795 ( .A1(n2009), .A2(n3803), .ZN(n2010) );
  NAND2_X1 U2796 ( .A1(n4693), .A2(REG2_REG_7__SCAN_IN), .ZN(n2011) );
  OR2_X1 U2797 ( .A1(n2438), .A2(n2219), .ZN(n2012) );
  INV_X1 U2798 ( .A(n2082), .ZN(n2081) );
  OAI21_X1 U2799 ( .B1(n3608), .B2(n3633), .A(n3768), .ZN(n2082) );
  OR2_X1 U2800 ( .A1(n2193), .A2(n2298), .ZN(n2013) );
  AND2_X1 U2801 ( .A1(n2191), .A2(REG2_REG_1__SCAN_IN), .ZN(n2014) );
  NAND3_X1 U2802 ( .A1(n2151), .A2(n2048), .A3(n2150), .ZN(n2156) );
  AND2_X1 U2803 ( .A1(n4211), .A2(n4229), .ZN(n2015) );
  AND2_X1 U2804 ( .A1(n2803), .A2(n2043), .ZN(n2016) );
  INV_X1 U2805 ( .A(n2571), .ZN(n2206) );
  AND2_X1 U2806 ( .A1(n2990), .A2(n2984), .ZN(n3838) );
  AND2_X1 U2807 ( .A1(n2258), .A2(n4197), .ZN(n2017) );
  AND2_X1 U2808 ( .A1(n4272), .A2(n4255), .ZN(n4239) );
  NOR2_X1 U2809 ( .A1(n4715), .A2(n4714), .ZN(n2018) );
  NAND2_X1 U2810 ( .A1(n3534), .A2(n4487), .ZN(n2019) );
  AND4_X1 U2811 ( .A1(n2423), .A2(n2313), .A3(n2312), .A4(n2711), .ZN(n2320)
         );
  INV_X1 U2812 ( .A(n2210), .ZN(n2209) );
  NAND2_X1 U2813 ( .A1(n3405), .A2(n2019), .ZN(n2210) );
  AND2_X1 U2814 ( .A1(n2093), .A2(n2090), .ZN(n2020) );
  NAND2_X1 U2815 ( .A1(n2265), .A2(n2270), .ZN(n3812) );
  AND2_X1 U2816 ( .A1(n3559), .A2(n3758), .ZN(n2021) );
  NOR2_X1 U2817 ( .A1(n2229), .A2(n2598), .ZN(n2022) );
  OR2_X1 U2818 ( .A1(n2318), .A2(n2317), .ZN(n2355) );
  NAND2_X1 U2819 ( .A1(n4303), .A2(n2542), .ZN(n4293) );
  OR2_X1 U2820 ( .A1(n3024), .A2(n2116), .ZN(n2023) );
  NAND2_X1 U2821 ( .A1(n3775), .A2(n3779), .ZN(n3723) );
  NAND2_X1 U2822 ( .A1(n2276), .A2(n2281), .ZN(n3732) );
  NAND2_X1 U2823 ( .A1(n4022), .A2(n3029), .ZN(n2024) );
  OR2_X1 U2824 ( .A1(n4693), .A2(REG1_REG_7__SCAN_IN), .ZN(n2025) );
  INV_X1 U2825 ( .A(IR_REG_30__SCAN_IN), .ZN(n3600) );
  OR2_X1 U2826 ( .A1(n3234), .A2(n3233), .ZN(n2026) );
  AND2_X1 U2827 ( .A1(n4470), .A2(n4368), .ZN(n2027) );
  AND2_X1 U2828 ( .A1(n4459), .A2(n4350), .ZN(n2028) );
  AND2_X1 U2829 ( .A1(n3736), .A2(n4017), .ZN(n2029) );
  AND2_X1 U2830 ( .A1(n4313), .A2(n4296), .ZN(n2030) );
  AND2_X1 U2831 ( .A1(n2294), .A2(n3682), .ZN(n2031) );
  AND2_X1 U2832 ( .A1(n2259), .A2(n2326), .ZN(n2032) );
  AND2_X1 U2833 ( .A1(n2790), .A2(n2789), .ZN(n2033) );
  AND2_X1 U2834 ( .A1(n4490), .A2(n3802), .ZN(n2034) );
  AND2_X1 U2835 ( .A1(n2024), .A2(n2387), .ZN(n2035) );
  AND2_X1 U2836 ( .A1(REG3_REG_6__SCAN_IN), .A2(REG3_REG_7__SCAN_IN), .ZN(
        n2036) );
  INV_X1 U2837 ( .A(n2084), .ZN(n2083) );
  AND2_X1 U2838 ( .A1(n3163), .A2(n2026), .ZN(n2037) );
  INV_X1 U2839 ( .A(n2528), .ZN(n2065) );
  OR2_X1 U2840 ( .A1(n3887), .A2(n3889), .ZN(n2038) );
  INV_X1 U2841 ( .A(n2279), .ZN(n2278) );
  NAND2_X1 U2842 ( .A1(n3733), .A2(n2280), .ZN(n2279) );
  INV_X1 U2843 ( .A(n2920), .ZN(n2102) );
  INV_X1 U2844 ( .A(n2510), .ZN(n2064) );
  INV_X1 U2845 ( .A(n2147), .ZN(n2581) );
  NOR2_X1 U2846 ( .A1(n2573), .A2(n2572), .ZN(n2147) );
  XNOR2_X1 U2847 ( .A(n2974), .B(n3658), .ZN(n2977) );
  NAND2_X1 U2848 ( .A1(n4383), .A2(n2743), .ZN(n2039) );
  AND2_X1 U2849 ( .A1(n2198), .A2(n2200), .ZN(n2040) );
  AND2_X1 U2850 ( .A1(n2164), .A2(n2163), .ZN(n2041) );
  INV_X1 U2851 ( .A(IR_REG_29__SCAN_IN), .ZN(n4576) );
  INV_X1 U2852 ( .A(IR_REG_28__SCAN_IN), .ZN(n2316) );
  NAND2_X1 U2853 ( .A1(n4018), .A2(n3342), .ZN(n2042) );
  NOR2_X1 U2854 ( .A1(n3310), .A2(n2438), .ZN(n2223) );
  NAND2_X1 U2855 ( .A1(n2103), .A2(n2102), .ZN(n2104) );
  XNOR2_X1 U2856 ( .A(n2448), .B(n2520), .ZN(n3463) );
  INV_X1 U2857 ( .A(n3024), .ZN(n2110) );
  XNOR2_X1 U2858 ( .A(n2437), .B(IR_REG_10__SCAN_IN), .ZN(n4691) );
  OAI21_X1 U2859 ( .B1(n3265), .B2(n2428), .A(n2427), .ZN(n3310) );
  NAND2_X1 U2860 ( .A1(n3525), .A2(n3524), .ZN(n3797) );
  OAI21_X1 U2861 ( .B1(n2069), .B2(n2210), .A(n2066), .ZN(n4356) );
  NAND2_X1 U2862 ( .A1(n3416), .A2(n2447), .ZN(n3353) );
  NAND2_X1 U2863 ( .A1(n3172), .A2(n2299), .ZN(n3235) );
  NAND2_X1 U2864 ( .A1(n2288), .A2(n2286), .ZN(n3276) );
  OR2_X1 U2865 ( .A1(n4787), .A2(n2799), .ZN(n2043) );
  OR2_X1 U2866 ( .A1(n3725), .A2(n3724), .ZN(n2044) );
  OR2_X1 U2867 ( .A1(n4016), .A2(n4197), .ZN(n3922) );
  INV_X1 U2868 ( .A(REG3_REG_10__SCAN_IN), .ZN(n2141) );
  AND2_X1 U2869 ( .A1(n3590), .A2(n3589), .ZN(n2045) );
  AND2_X1 U2870 ( .A1(n2256), .A2(n4296), .ZN(n2046) );
  NAND3_X1 U2871 ( .A1(n2814), .A2(n2337), .A3(n2663), .ZN(n2831) );
  OR2_X1 U2872 ( .A1(n4100), .A2(n4675), .ZN(n2047) );
  INV_X1 U2873 ( .A(n2298), .ZN(n2200) );
  NAND2_X1 U2874 ( .A1(n2069), .A2(n2068), .ZN(n3449) );
  OR2_X1 U2875 ( .A1(n3463), .A2(n3464), .ZN(n2048) );
  AND2_X1 U2876 ( .A1(n2211), .A2(n2019), .ZN(n2049) );
  INV_X1 U2877 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4651) );
  NAND2_X1 U2878 ( .A1(n2831), .A2(n2343), .ZN(n3036) );
  OR2_X1 U2879 ( .A1(n3495), .A2(REG1_REG_17__SCAN_IN), .ZN(n2050) );
  AND2_X1 U2880 ( .A1(n4732), .A2(n2050), .ZN(n2051) );
  XNOR2_X1 U2881 ( .A(n2977), .B(n2978), .ZN(n3006) );
  INV_X1 U2882 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2145) );
  INV_X1 U2883 ( .A(n2197), .ZN(n2196) );
  NAND2_X1 U2884 ( .A1(n3110), .A2(n3105), .ZN(n2197) );
  OAI22_X1 U2885 ( .A1(n2969), .A2(n2932), .B1(n3123), .B2(n2931), .ZN(n2971)
         );
  AND2_X1 U2886 ( .A1(n2914), .A2(n2913), .ZN(n2052) );
  AND2_X1 U2887 ( .A1(n2195), .A2(n2197), .ZN(n2053) );
  AND2_X1 U2888 ( .A1(n2017), .A2(n4182), .ZN(n2054) );
  XNOR2_X1 U2889 ( .A(n2406), .B(IR_REG_7__SCAN_IN), .ZN(n4693) );
  INV_X1 U2890 ( .A(n4693), .ZN(n2175) );
  XNOR2_X1 U2891 ( .A(n2890), .B(n2884), .ZN(n2889) );
  NAND2_X1 U2892 ( .A1(n2108), .A2(n2107), .ZN(n3599) );
  NAND4_X1 U2893 ( .A1(n2285), .A2(n2284), .A3(n2424), .A4(n2320), .ZN(n2055)
         );
  NOR2_X2 U2894 ( .A1(n2649), .A2(n2056), .ZN(n2285) );
  NAND2_X1 U2895 ( .A1(n2831), .A2(n2058), .ZN(n2057) );
  NAND2_X1 U2896 ( .A1(n2357), .A2(n2356), .ZN(n2070) );
  NAND3_X1 U2897 ( .A1(n2127), .A2(n2318), .A3(REG0_REG_4__SCAN_IN), .ZN(n2072) );
  XNOR2_X2 U2898 ( .A(n2087), .B(n3600), .ZN(n2318) );
  NOR2_X1 U2899 ( .A1(n3007), .A2(n2979), .ZN(n2980) );
  NOR2_X1 U2900 ( .A1(n3008), .A2(n3006), .ZN(n3007) );
  AND4_X2 U2901 ( .A1(n2661), .A2(n2304), .A3(n2659), .A4(n2660), .ZN(n2928)
         );
  OR2_X1 U2902 ( .A1(n3609), .A2(n2085), .ZN(n2075) );
  NAND2_X1 U2903 ( .A1(n3609), .A2(n2080), .ZN(n2079) );
  NAND2_X2 U2904 ( .A1(n3609), .A2(n3608), .ZN(n3710) );
  OAI21_X1 U2905 ( .B1(n3608), .B2(n2085), .A(n3613), .ZN(n2084) );
  INV_X1 U2906 ( .A(n3630), .ZN(n2085) );
  OAI21_X2 U2907 ( .B1(n3797), .B2(n2279), .A(n2273), .ZN(n3690) );
  AND2_X4 U2908 ( .A1(n2318), .A2(n2317), .ZN(n2345) );
  XNOR2_X2 U2909 ( .A(n2086), .B(IR_REG_29__SCAN_IN), .ZN(n2317) );
  NAND2_X1 U2910 ( .A1(n2089), .A2(n2894), .ZN(n4054) );
  NAND2_X1 U2911 ( .A1(n4037), .A2(REG2_REG_4__SCAN_IN), .ZN(n2089) );
  NAND2_X1 U2912 ( .A1(n2093), .A2(n4691), .ZN(n2097) );
  NOR2_X1 U2913 ( .A1(n3381), .A2(n3313), .ZN(n2092) );
  INV_X1 U2914 ( .A(n2096), .ZN(n3481) );
  INV_X1 U2915 ( .A(n2918), .ZN(n2105) );
  INV_X1 U2916 ( .A(n2104), .ZN(n3056) );
  INV_X2 U2917 ( .A(IR_REG_0__SCAN_IN), .ZN(n2231) );
  NAND2_X1 U2918 ( .A1(n2114), .A2(n3063), .ZN(n2112) );
  OAI21_X1 U2919 ( .B1(n3063), .B2(n2023), .A(n2114), .ZN(n3094) );
  OAI21_X1 U2920 ( .B1(n3182), .B2(n2121), .A(n2007), .ZN(n3348) );
  NAND2_X1 U2921 ( .A1(n2118), .A2(n2117), .ZN(n2672) );
  NAND2_X1 U2922 ( .A1(n3182), .A2(n2007), .ZN(n2118) );
  OAI211_X2 U2923 ( .C1(n2353), .C2(n3014), .A(n2126), .B(n2122), .ZN(n2333)
         );
  NAND2_X1 U2924 ( .A1(n2123), .A2(n2318), .ZN(n2122) );
  NAND2_X1 U2925 ( .A1(n2317), .A2(REG1_REG_1__SCAN_IN), .ZN(n2124) );
  INV_X1 U2926 ( .A(n2318), .ZN(n4686) );
  MUX2_X1 U2927 ( .A(n2133), .B(n4001), .S(n2728), .Z(n4002) );
  INV_X1 U2928 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2146) );
  NAND2_X1 U2929 ( .A1(n2939), .A2(n2940), .ZN(n2938) );
  NAND2_X1 U2930 ( .A1(n3375), .A2(n4691), .ZN(n2157) );
  NAND2_X1 U2931 ( .A1(n4081), .A2(n2161), .ZN(n2160) );
  NAND2_X1 U2932 ( .A1(n3468), .A2(n4689), .ZN(n2165) );
  NOR2_X1 U2933 ( .A1(n4104), .A2(n3474), .ZN(n4715) );
  NAND2_X2 U2934 ( .A1(n2176), .A2(n2174), .ZN(n3111) );
  INV_X1 U2935 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2178) );
  NOR2_X4 U2936 ( .A1(n3210), .A2(n2297), .ZN(n3374) );
  XNOR2_X2 U2937 ( .A(n3374), .B(n4691), .ZN(n3376) );
  NAND2_X2 U2938 ( .A1(n4073), .A2(n3467), .ZN(n3468) );
  NAND2_X1 U2939 ( .A1(n4083), .A2(n3488), .ZN(n2181) );
  NAND2_X2 U2940 ( .A1(n2190), .A2(n2191), .ZN(n2870) );
  OAI211_X1 U2941 ( .C1(n2190), .C2(REG2_REG_1__SCAN_IN), .A(n2188), .B(n2187), 
        .ZN(n4029) );
  NAND2_X1 U2942 ( .A1(n4029), .A2(n2872), .ZN(n4028) );
  AOI21_X1 U2943 ( .B1(n2201), .B2(n4709), .A(n4719), .ZN(n4712) );
  NAND2_X1 U2944 ( .A1(n4250), .A2(n2005), .ZN(n2202) );
  NAND2_X1 U2945 ( .A1(n3184), .A2(n2412), .ZN(n2415) );
  INV_X1 U2946 ( .A(n2223), .ZN(n2222) );
  NAND2_X1 U2947 ( .A1(n2222), .A2(n2224), .ZN(n3414) );
  OR2_X1 U2948 ( .A1(n3427), .A2(n3397), .ZN(n2224) );
  NAND2_X1 U2949 ( .A1(n2590), .A2(n2589), .ZN(n4191) );
  INV_X1 U2950 ( .A(n2674), .ZN(n4265) );
  NAND2_X1 U2951 ( .A1(n2674), .A2(n3869), .ZN(n2230) );
  NAND3_X2 U2952 ( .A1(n2231), .A2(n2232), .A3(n2309), .ZN(n2344) );
  NAND2_X1 U2953 ( .A1(n2796), .A2(n2243), .ZN(n2242) );
  NAND2_X1 U2954 ( .A1(n2796), .A2(n3970), .ZN(n2795) );
  NAND2_X1 U2955 ( .A1(n2249), .A2(n2246), .ZN(n2665) );
  NAND2_X1 U2956 ( .A1(n4339), .A2(n2253), .ZN(n4282) );
  AND2_X2 U2957 ( .A1(n4239), .A2(n2054), .ZN(n4177) );
  NAND4_X1 U2958 ( .A1(n2321), .A2(n2320), .A3(n2260), .A4(n2424), .ZN(n2259)
         );
  AND2_X1 U2959 ( .A1(n2424), .A2(n2261), .ZN(n2385) );
  NAND3_X1 U2960 ( .A1(n2321), .A2(n2320), .A3(n2385), .ZN(n2701) );
  INV_X1 U2961 ( .A(n2424), .ZN(n2372) );
  INV_X1 U2962 ( .A(IR_REG_5__SCAN_IN), .ZN(n2261) );
  NAND2_X1 U2963 ( .A1(n3746), .A2(n2266), .ZN(n2262) );
  NAND2_X1 U2964 ( .A1(n2262), .A2(n2263), .ZN(n3716) );
  NAND4_X1 U2965 ( .A1(n2285), .A2(n2424), .A3(n2320), .A4(n2650), .ZN(n2657)
         );
  NOR2_X4 U2966 ( .A1(n2344), .A2(n2311), .ZN(n2424) );
  NAND2_X1 U2967 ( .A1(n3164), .A2(n2037), .ZN(n2288) );
  NAND2_X2 U2968 ( .A1(n2290), .A2(n2045), .ZN(n3609) );
  NAND2_X1 U2969 ( .A1(n3710), .A2(n2292), .ZN(n2291) );
  NAND2_X1 U2970 ( .A1(n2291), .A2(n2294), .ZN(n3683) );
  AOI21_X1 U2971 ( .B1(n3710), .B2(n3642), .A(n3641), .ZN(n3822) );
  INV_X1 U2972 ( .A(n3641), .ZN(n2296) );
  NOR2_X2 U2973 ( .A1(n3114), .A2(n3113), .ZN(n3210) );
  AOI21_X2 U2974 ( .B1(n3112), .B2(REG1_REG_8__SCAN_IN), .A(n2300), .ZN(n3114)
         );
  XNOR2_X2 U2975 ( .A(n3468), .B(n4086), .ZN(n4081) );
  AND2_X1 U2976 ( .A1(n3767), .A2(n3766), .ZN(n3769) );
  AND2_X1 U2977 ( .A1(n2969), .A2(n3645), .ZN(n2970) );
  INV_X1 U2978 ( .A(n2870), .ZN(n2332) );
  OR2_X1 U2979 ( .A1(n2347), .A2(n2335), .ZN(n2661) );
  NAND2_X1 U2980 ( .A1(n3450), .A2(n4470), .ZN(n3406) );
  AND2_X1 U2981 ( .A1(n2385), .A2(n2526), .ZN(n2540) );
  NOR2_X1 U2982 ( .A1(n2971), .A2(n2970), .ZN(n3008) );
  NAND2_X1 U2983 ( .A1(n4177), .A2(n3827), .ZN(n2747) );
  OR2_X1 U2984 ( .A1(n4176), .A2(n2620), .ZN(n2767) );
  NAND2_X1 U2985 ( .A1(n2783), .A2(n2782), .ZN(n2785) );
  NAND2_X1 U2986 ( .A1(n2783), .A2(n2788), .ZN(n2790) );
  INV_X2 U2987 ( .A(n3660), .ZN(n2972) );
  NAND2_X1 U2988 ( .A1(n2342), .A2(n2967), .ZN(n3854) );
  NAND2_X1 U2989 ( .A1(n2778), .A2(n3914), .ZN(n4119) );
  OR2_X1 U2990 ( .A1(n4145), .A2(n4483), .ZN(n2734) );
  INV_X1 U2991 ( .A(n3506), .ZN(n2859) );
  NAND2_X1 U2992 ( .A1(n3506), .A2(DATAI_0_), .ZN(n2336) );
  OAI21_X1 U2993 ( .B1(n3506), .B2(n2332), .A(n2331), .ZN(n2334) );
  AND2_X1 U2994 ( .A1(n4692), .A2(REG1_REG_9__SCAN_IN), .ZN(n2297) );
  AND2_X1 U2995 ( .A1(n4692), .A2(REG2_REG_9__SCAN_IN), .ZN(n2298) );
  INV_X1 U2996 ( .A(n2707), .ZN(n2697) );
  OR2_X1 U2997 ( .A1(n3171), .A2(n3170), .ZN(n2299) );
  AND2_X1 U2998 ( .A1(n3111), .A2(n2199), .ZN(n2300) );
  AND2_X1 U2999 ( .A1(n2785), .A2(n2784), .ZN(n2301) );
  NAND2_X1 U3000 ( .A1(n3792), .A2(n3702), .ZN(n2302) );
  INV_X1 U3001 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3464) );
  INV_X1 U3002 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2880) );
  INV_X1 U3003 ( .A(n4483), .ZN(n2782) );
  INV_X1 U3004 ( .A(n4546), .ZN(n2788) );
  INV_X1 U3005 ( .A(n4237), .ZN(n2580) );
  OR2_X1 U3006 ( .A1(n4771), .A2(n3475), .ZN(n2303) );
  NAND2_X1 U3007 ( .A1(n4119), .A2(n2781), .ZN(n4129) );
  INV_X1 U3008 ( .A(n4129), .ZN(n2783) );
  AND2_X2 U3009 ( .A1(n2823), .A2(n4755), .ZN(n4745) );
  INV_X1 U3010 ( .A(n4745), .ZN(n4752) );
  INV_X1 U3011 ( .A(n3847), .ZN(n2662) );
  INV_X1 U3012 ( .A(IR_REG_31__SCAN_IN), .ZN(n2637) );
  INV_X1 U3013 ( .A(n4075), .ZN(n3466) );
  INV_X1 U3014 ( .A(n3932), .ZN(n3417) );
  NAND2_X1 U3015 ( .A1(n2345), .A2(REG1_REG_0__SCAN_IN), .ZN(n2304) );
  INV_X2 U3016 ( .A(n4784), .ZN(n4787) );
  OR2_X1 U3017 ( .A1(n2821), .A2(n2732), .ZN(n4784) );
  OAI21_X1 U3018 ( .B1(n3788), .B2(n3540), .A(n3695), .ZN(n3538) );
  INV_X1 U3019 ( .A(n3538), .ZN(n3539) );
  INV_X1 U3020 ( .A(IR_REG_27__SCAN_IN), .ZN(n2308) );
  INV_X1 U3021 ( .A(IR_REG_18__SCAN_IN), .ZN(n4563) );
  INV_X1 U3022 ( .A(IR_REG_9__SCAN_IN), .ZN(n2314) );
  INV_X1 U3023 ( .A(n3931), .ZN(n2673) );
  INV_X1 U3024 ( .A(n3570), .ZN(n3571) );
  OR2_X1 U3025 ( .A1(n4047), .A2(n2904), .ZN(n2905) );
  AND2_X1 U3026 ( .A1(n4447), .A2(n4329), .ZN(n3931) );
  AND2_X1 U3027 ( .A1(n3185), .A2(n2411), .ZN(n2412) );
  NOR2_X1 U3028 ( .A1(n2640), .A2(n2639), .ZN(n2641) );
  OR2_X1 U3029 ( .A1(n3279), .A2(n3278), .ZN(n3280) );
  INV_X1 U3030 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4608) );
  NAND2_X1 U3031 ( .A1(n4697), .A2(n2880), .ZN(n2879) );
  AND2_X1 U3032 ( .A1(n2917), .A2(n4694), .ZN(n2918) );
  NAND2_X1 U3033 ( .A1(n3491), .A2(n4106), .ZN(n3492) );
  OR2_X1 U3034 ( .A1(n4016), .A2(n4392), .ZN(n2597) );
  OR2_X1 U3035 ( .A1(n4230), .A2(n4410), .ZN(n2570) );
  NAND2_X1 U3036 ( .A1(n3506), .A2(DATAI_1_), .ZN(n2331) );
  AND2_X1 U3037 ( .A1(n2625), .A2(n2624), .ZN(n2766) );
  INV_X1 U3038 ( .A(n4340), .ZN(n2509) );
  INV_X1 U3039 ( .A(n3792), .ZN(n3534) );
  INV_X1 U3040 ( .A(n3284), .ZN(n3289) );
  NOR2_X1 U3041 ( .A1(n3667), .A2(n3831), .ZN(n3668) );
  INV_X1 U3042 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2468) );
  OAI21_X1 U3043 ( .B1(n4697), .B2(n2880), .A(n2879), .ZN(n2940) );
  INV_X1 U3044 ( .A(n2914), .ZN(n2906) );
  AND2_X1 U3045 ( .A1(n4205), .A2(n2678), .ZN(n4237) );
  INV_X1 U3046 ( .A(n4421), .ZN(n4313) );
  INV_X1 U3047 ( .A(n4449), .ZN(n4345) );
  AND2_X1 U3048 ( .A1(n3856), .A2(n3853), .ZN(n3939) );
  NAND2_X1 U3049 ( .A1(n4784), .A2(REG1_REG_29__SCAN_IN), .ZN(n2784) );
  INV_X1 U3050 ( .A(n4409), .ZN(n4489) );
  AND2_X1 U3051 ( .A1(n3506), .A2(DATAI_20_), .ZN(n4420) );
  INV_X1 U3052 ( .A(n3803), .ZN(n3418) );
  AND2_X1 U3053 ( .A1(n2704), .A2(n2708), .ZN(n2817) );
  INV_X1 U3054 ( .A(IR_REG_23__SCAN_IN), .ZN(n2711) );
  OR2_X1 U3055 ( .A1(n2477), .A2(IR_REG_14__SCAN_IN), .ZN(n2485) );
  AND2_X1 U3056 ( .A1(n2519), .A2(n2518), .ZN(n3751) );
  NAND2_X1 U3057 ( .A1(n4051), .A2(n4052), .ZN(n4050) );
  INV_X1 U3058 ( .A(n4719), .ZN(n4110) );
  AND2_X1 U3059 ( .A1(n3871), .A2(n3979), .ZN(n4340) );
  INV_X1 U3060 ( .A(n4378), .ZN(n4336) );
  INV_X1 U3061 ( .A(n4364), .ZN(n4741) );
  OR2_X1 U3062 ( .A1(n4745), .A2(n4386), .ZN(n4369) );
  INV_X1 U3063 ( .A(n2951), .ZN(n2821) );
  INV_X1 U3064 ( .A(n4229), .ZN(n4241) );
  INV_X1 U3065 ( .A(n4497), .ZN(n4480) );
  INV_X1 U3066 ( .A(n3200), .ZN(n4492) );
  AND2_X1 U3067 ( .A1(n3123), .A2(n4768), .ZN(n2982) );
  XNOR2_X1 U3068 ( .A(n2499), .B(n2498), .ZN(n4106) );
  AND2_X1 U3069 ( .A1(n2877), .A2(n2860), .ZN(n4722) );
  INV_X1 U3070 ( .A(n3838), .ZN(n3831) );
  INV_X1 U3071 ( .A(n4414), .ZN(n4211) );
  INV_X1 U3072 ( .A(n3304), .ZN(n4020) );
  INV_X1 U3073 ( .A(U4043), .ZN(n4025) );
  OR2_X1 U3074 ( .A1(n4708), .A2(n4007), .ZN(n4719) );
  AOI21_X1 U3075 ( .B1(n4728), .B2(n4727), .A(n4726), .ZN(n4734) );
  OR2_X1 U3076 ( .A1(n2822), .A2(n2986), .ZN(n4755) );
  NAND2_X1 U3077 ( .A1(n4787), .A2(n4492), .ZN(n4483) );
  NAND2_X1 U3078 ( .A1(n4783), .A2(n4492), .ZN(n4546) );
  INV_X1 U3079 ( .A(n4767), .ZN(n4766) );
  AND2_X1 U3080 ( .A1(n3122), .A2(STATE_REG_SCAN_IN), .ZN(n4768) );
  INV_X1 U3081 ( .A(n2808), .ZN(U4043) );
  NOR2_X1 U3082 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_22__SCAN_IN), .ZN(n2313)
         );
  NOR2_X1 U3083 ( .A1(IR_REG_6__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2312)
         );
  INV_X1 U3084 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3014) );
  INV_X1 U3085 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4560) );
  INV_X1 U3086 ( .A(n2649), .ZN(n2319) );
  NAND2_X1 U3087 ( .A1(n2319), .A2(n2650), .ZN(n2636) );
  NAND3_X1 U3088 ( .A1(n2701), .A2(IR_REG_27__SCAN_IN), .A3(IR_REG_31__SCAN_IN), .ZN(n2328) );
  NAND2_X1 U3089 ( .A1(n2322), .A2(n2316), .ZN(n2327) );
  INV_X1 U3090 ( .A(n2322), .ZN(n2323) );
  NAND2_X1 U3091 ( .A1(n2323), .A2(IR_REG_27__SCAN_IN), .ZN(n2324) );
  NAND2_X1 U3092 ( .A1(n2324), .A2(IR_REG_31__SCAN_IN), .ZN(n2325) );
  OAI21_X1 U3093 ( .B1(IR_REG_31__SCAN_IN), .B2(n2316), .A(n2325), .ZN(n2326)
         );
  NAND2_X1 U3094 ( .A1(n2328), .A2(n2032), .ZN(n2330) );
  NAND2_X1 U3095 ( .A1(n2316), .A2(IR_REG_27__SCAN_IN), .ZN(n2329) );
  NAND2_X4 U3096 ( .A1(n2330), .A2(n2329), .ZN(n3506) );
  INV_X1 U3097 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2335) );
  INV_X1 U3098 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2935) );
  INV_X1 U3099 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2999) );
  NAND4_X1 U3100 ( .A1(n2661), .A2(n2304), .A3(n2659), .A4(n2660), .ZN(n4026)
         );
  AND2_X1 U3101 ( .A1(n4026), .A2(n2997), .ZN(n2811) );
  NAND2_X1 U3102 ( .A1(n2333), .A2(n3011), .ZN(n2337) );
  NAND2_X1 U3103 ( .A1(n2345), .A2(REG1_REG_2__SCAN_IN), .ZN(n2341) );
  INV_X1 U3104 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2994) );
  OR2_X1 U3105 ( .A1(n2353), .A2(n2994), .ZN(n2340) );
  INV_X1 U3106 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2869) );
  OR2_X1 U3107 ( .A1(n2355), .A2(n2869), .ZN(n2339) );
  INV_X1 U3108 ( .A(REG0_REG_2__SCAN_IN), .ZN(n3021) );
  OR2_X1 U3109 ( .A1(n2347), .A2(n3021), .ZN(n2338) );
  MUX2_X1 U3110 ( .A(n4697), .B(DATAI_2_), .S(n3506), .Z(n3073) );
  NAND2_X1 U3111 ( .A1(n3068), .A2(n3073), .ZN(n3851) );
  INV_X1 U3112 ( .A(n3068), .ZN(n2342) );
  NAND2_X1 U3113 ( .A1(n3068), .A2(n2967), .ZN(n2343) );
  NAND2_X1 U3114 ( .A1(n2344), .A2(IR_REG_31__SCAN_IN), .ZN(n2359) );
  XNOR2_X1 U3115 ( .A(n2359), .B(IR_REG_3__SCAN_IN), .ZN(n4696) );
  MUX2_X1 U3116 ( .A(n4696), .B(DATAI_3_), .S(n3506), .Z(n3072) );
  NAND2_X1 U3117 ( .A1(n2614), .A2(REG2_REG_3__SCAN_IN), .ZN(n2351) );
  OR2_X1 U3118 ( .A1(n2353), .A2(REG3_REG_3__SCAN_IN), .ZN(n2350) );
  INV_X1 U3119 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3079) );
  INV_X1 U3120 ( .A(REG0_REG_3__SCAN_IN), .ZN(n3089) );
  OR2_X1 U3121 ( .A1(n2347), .A2(n3089), .ZN(n2348) );
  NAND2_X1 U3122 ( .A1(n2345), .A2(REG1_REG_4__SCAN_IN), .ZN(n2357) );
  INV_X1 U3123 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2352) );
  XNOR2_X1 U3124 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(n3154) );
  INV_X1 U3125 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2354) );
  OR2_X1 U3126 ( .A1(n2355), .A2(n2354), .ZN(n2356) );
  NAND2_X1 U3127 ( .A1(n2359), .A2(n2358), .ZN(n2360) );
  NAND2_X1 U3128 ( .A1(n2360), .A2(IR_REG_31__SCAN_IN), .ZN(n2361) );
  MUX2_X1 U3129 ( .A(n4695), .B(DATAI_4_), .S(n3506), .Z(n3042) );
  NAND2_X1 U3130 ( .A1(n3249), .A2(n3042), .ZN(n3857) );
  INV_X1 U3131 ( .A(n3042), .ZN(n3150) );
  AND2_X1 U3132 ( .A1(n4024), .A2(n3072), .ZN(n2362) );
  AOI22_X1 U3133 ( .A1(n3040), .A2(n2362), .B1(n3042), .B2(n4023), .ZN(n2363)
         );
  NAND2_X1 U3134 ( .A1(n2758), .A2(REG0_REG_5__SCAN_IN), .ZN(n2371) );
  INV_X1 U3135 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2904) );
  OR2_X1 U3136 ( .A1(n2346), .A2(n2904), .ZN(n2370) );
  INV_X1 U3137 ( .A(n2364), .ZN(n2366) );
  INV_X1 U3138 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2365) );
  NAND2_X1 U3139 ( .A1(n2366), .A2(n2365), .ZN(n2367) );
  NAND2_X1 U3140 ( .A1(n2379), .A2(n2367), .ZN(n3250) );
  OR2_X1 U3141 ( .A1(n2353), .A2(n3250), .ZN(n2369) );
  INV_X1 U3142 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2895) );
  OR2_X1 U3143 ( .A1(n3510), .A2(n2895), .ZN(n2368) );
  NAND2_X1 U3144 ( .A1(n2372), .A2(IR_REG_31__SCAN_IN), .ZN(n2373) );
  INV_X1 U3145 ( .A(DATAI_5_), .ZN(n2374) );
  MUX2_X1 U3146 ( .A(n4047), .B(n2374), .S(n3506), .Z(n3246) );
  NAND2_X1 U3147 ( .A1(n3160), .A2(n3246), .ZN(n2375) );
  INV_X1 U31480 ( .A(n3246), .ZN(n3029) );
  NAND2_X1 U31490 ( .A1(n2758), .A2(REG0_REG_6__SCAN_IN), .ZN(n2384) );
  INV_X1 U3150 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2376) );
  OR2_X1 U3151 ( .A1(n2346), .A2(n2376), .ZN(n2383) );
  INV_X1 U3152 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2378) );
  NAND2_X1 U3153 ( .A1(n2379), .A2(n2378), .ZN(n2380) );
  NAND2_X1 U3154 ( .A1(n2388), .A2(n2380), .ZN(n3297) );
  OR2_X1 U3155 ( .A1(n2353), .A2(n3297), .ZN(n2382) );
  INV_X1 U3156 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3298) );
  OR2_X1 U3157 ( .A1(n3510), .A2(n3298), .ZN(n2381) );
  NAND4_X1 U3158 ( .A1(n2384), .A2(n2383), .A3(n2382), .A4(n2381), .ZN(n4021)
         );
  OR2_X1 U3159 ( .A1(n2385), .A2(n2637), .ZN(n2386) );
  MUX2_X1 U3160 ( .A(n4694), .B(DATAI_6_), .S(n3506), .Z(n3301) );
  NAND2_X1 U3161 ( .A1(n4021), .A2(n3301), .ZN(n2387) );
  NAND2_X1 U3162 ( .A1(n2758), .A2(REG0_REG_7__SCAN_IN), .ZN(n2394) );
  OR2_X1 U3163 ( .A1(n2346), .A2(n2178), .ZN(n2393) );
  INV_X1 U3164 ( .A(REG3_REG_7__SCAN_IN), .ZN(n4562) );
  NAND2_X1 U3165 ( .A1(n2388), .A2(n4562), .ZN(n2389) );
  NAND2_X1 U3166 ( .A1(n2399), .A2(n2389), .ZN(n3260) );
  OR2_X1 U3167 ( .A1(n2353), .A2(n3260), .ZN(n2392) );
  INV_X1 U3168 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2390) );
  OR2_X1 U3169 ( .A1(n3510), .A2(n2390), .ZN(n2391) );
  AND2_X1 U3170 ( .A1(n2385), .A2(n2422), .ZN(n2395) );
  MUX2_X1 U3171 ( .A(n4693), .B(DATAI_7_), .S(n3506), .Z(n3204) );
  NAND2_X1 U3172 ( .A1(n3304), .A2(n3204), .ZN(n2664) );
  INV_X1 U3173 ( .A(n3204), .ZN(n3240) );
  NAND2_X1 U3174 ( .A1(n4020), .A2(n3240), .ZN(n3872) );
  NAND2_X1 U3175 ( .A1(n2664), .A2(n3872), .ZN(n3185) );
  NAND2_X1 U3176 ( .A1(n3248), .A2(n3177), .ZN(n3183) );
  NAND2_X1 U3177 ( .A1(n2758), .A2(REG0_REG_8__SCAN_IN), .ZN(n2404) );
  INV_X1 U3178 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2396) );
  OR2_X1 U3179 ( .A1(n2346), .A2(n2396), .ZN(n2403) );
  INV_X1 U3180 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2398) );
  NAND2_X1 U3181 ( .A1(n2399), .A2(n2398), .ZN(n2400) );
  NAND2_X1 U3182 ( .A1(n2416), .A2(n2400), .ZN(n3225) );
  OR2_X1 U3183 ( .A1(n2353), .A2(n3225), .ZN(n2402) );
  INV_X1 U3184 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3105) );
  OR2_X1 U3185 ( .A1(n3510), .A2(n3105), .ZN(n2401) );
  INV_X1 U3186 ( .A(IR_REG_7__SCAN_IN), .ZN(n2405) );
  NAND2_X1 U3187 ( .A1(n2406), .A2(n2405), .ZN(n2407) );
  NAND2_X1 U3188 ( .A1(n2407), .A2(IR_REG_31__SCAN_IN), .ZN(n2409) );
  INV_X1 U3189 ( .A(DATAI_8_), .ZN(n2410) );
  MUX2_X1 U3190 ( .A(n3110), .B(n2410), .S(n3506), .Z(n3284) );
  NAND2_X1 U3191 ( .A1(n3341), .A2(n3284), .ZN(n2413) );
  AND2_X1 U3192 ( .A1(n4020), .A2(n3204), .ZN(n3186) );
  AOI22_X1 U3193 ( .A1(n2413), .A2(n3186), .B1(n3289), .B2(n4019), .ZN(n2414)
         );
  NAND2_X1 U3194 ( .A1(n2415), .A2(n2414), .ZN(n3265) );
  NAND2_X1 U3195 ( .A1(n2758), .A2(REG0_REG_9__SCAN_IN), .ZN(n2421) );
  INV_X1 U3196 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3321) );
  OR2_X1 U3197 ( .A1(n2346), .A2(n3321), .ZN(n2420) );
  NAND2_X1 U3198 ( .A1(n2416), .A2(n3107), .ZN(n2417) );
  NAND2_X1 U3199 ( .A1(n2429), .A2(n2417), .ZN(n3347) );
  OR2_X1 U3200 ( .A1(n2353), .A2(n3347), .ZN(n2419) );
  INV_X1 U3201 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3325) );
  NAND2_X1 U3202 ( .A1(n2425), .A2(n2424), .ZN(n2648) );
  NAND2_X1 U3203 ( .A1(n2648), .A2(IR_REG_31__SCAN_IN), .ZN(n2426) );
  XNOR2_X1 U3204 ( .A(n2426), .B(IR_REG_9__SCAN_IN), .ZN(n4692) );
  MUX2_X1 U3205 ( .A(n4692), .B(DATAI_9_), .S(n3506), .Z(n3266) );
  AND2_X1 U3206 ( .A1(n4018), .A2(n3266), .ZN(n2428) );
  NAND2_X1 U3207 ( .A1(n3338), .A2(n3342), .ZN(n2427) );
  NAND2_X1 U3208 ( .A1(n2758), .A2(REG0_REG_10__SCAN_IN), .ZN(n2434) );
  INV_X1 U3209 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4673) );
  OR2_X1 U32100 ( .A1(n2346), .A2(n4673), .ZN(n2433) );
  NAND2_X1 U32110 ( .A1(n2429), .A2(n2141), .ZN(n2430) );
  NAND2_X1 U32120 ( .A1(n2441), .A2(n2430), .ZN(n3402) );
  OR2_X1 U32130 ( .A1(n2353), .A2(n3402), .ZN(n2432) );
  INV_X1 U32140 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3313) );
  OR2_X1 U32150 ( .A1(n3510), .A2(n3313), .ZN(n2431) );
  NAND2_X1 U32160 ( .A1(n2524), .A2(n2385), .ZN(n2439) );
  NAND2_X1 U32170 ( .A1(n2439), .A2(IR_REG_31__SCAN_IN), .ZN(n2437) );
  MUX2_X1 U32180 ( .A(n4691), .B(DATAI_10_), .S(n3506), .Z(n2667) );
  NOR2_X1 U32190 ( .A1(n3806), .A2(n2667), .ZN(n2438) );
  NAND2_X1 U32200 ( .A1(n2461), .A2(IR_REG_31__SCAN_IN), .ZN(n2448) );
  INV_X1 U32210 ( .A(DATAI_11_), .ZN(n2440) );
  MUX2_X1 U32220 ( .A(n3463), .B(n2440), .S(n3506), .Z(n3803) );
  NAND2_X1 U32230 ( .A1(n2345), .A2(REG1_REG_11__SCAN_IN), .ZN(n2446) );
  INV_X1 U32240 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3438) );
  OR2_X1 U32250 ( .A1(n2347), .A2(n3438), .ZN(n2445) );
  NAND2_X1 U32260 ( .A1(n2441), .A2(n3383), .ZN(n2442) );
  NAND2_X1 U32270 ( .A1(n2453), .A2(n2442), .ZN(n3809) );
  OR2_X1 U32280 ( .A1(n2353), .A2(n3809), .ZN(n2444) );
  INV_X1 U32290 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3423) );
  OR2_X1 U32300 ( .A1(n3510), .A2(n3423), .ZN(n2443) );
  NAND4_X1 U32310 ( .A1(n2446), .A2(n2445), .A3(n2444), .A4(n2443), .ZN(n4484)
         );
  NAND2_X1 U32320 ( .A1(n3418), .A2(n3739), .ZN(n3349) );
  NAND2_X1 U32330 ( .A1(n3803), .A2(n4484), .ZN(n3351) );
  NAND2_X1 U32340 ( .A1(n3349), .A2(n3351), .ZN(n3932) );
  NAND2_X1 U32350 ( .A1(n3803), .A2(n3739), .ZN(n2447) );
  NAND2_X1 U32360 ( .A1(n2448), .A2(n2520), .ZN(n2449) );
  NAND2_X1 U32370 ( .A1(n2449), .A2(IR_REG_31__SCAN_IN), .ZN(n2450) );
  MUX2_X1 U32380 ( .A(n4690), .B(DATAI_12_), .S(n3506), .Z(n3736) );
  NAND2_X1 U32390 ( .A1(n2758), .A2(REG0_REG_12__SCAN_IN), .ZN(n2460) );
  INV_X1 U32400 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2452) );
  NAND2_X1 U32410 ( .A1(n2453), .A2(n2452), .ZN(n2454) );
  NAND2_X1 U32420 ( .A1(n2469), .A2(n2454), .ZN(n3356) );
  OR2_X1 U32430 ( .A1(n3356), .A2(n2353), .ZN(n2459) );
  INV_X1 U32440 ( .A(REG1_REG_12__SCAN_IN), .ZN(n2455) );
  OR2_X1 U32450 ( .A1(n2346), .A2(n2455), .ZN(n2458) );
  INV_X1 U32460 ( .A(REG2_REG_12__SCAN_IN), .ZN(n2456) );
  OR2_X1 U32470 ( .A1(n3510), .A2(n2456), .ZN(n2457) );
  NAND4_X1 U32480 ( .A1(n2460), .A2(n2459), .A3(n2458), .A4(n2457), .ZN(n4017)
         );
  INV_X1 U32490 ( .A(n3736), .ZN(n4490) );
  INV_X1 U32500 ( .A(DATAI_13_), .ZN(n2467) );
  INV_X1 U32510 ( .A(n2461), .ZN(n2463) );
  NOR2_X1 U32520 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2462) );
  NAND2_X1 U32530 ( .A1(n2463), .A2(n2462), .ZN(n2465) );
  NAND2_X1 U32540 ( .A1(n2465), .A2(IR_REG_31__SCAN_IN), .ZN(n2464) );
  MUX2_X1 U32550 ( .A(IR_REG_31__SCAN_IN), .B(n2464), .S(IR_REG_13__SCAN_IN), 
        .Z(n2466) );
  NAND2_X1 U32560 ( .A1(n2466), .A2(n2477), .ZN(n4075) );
  MUX2_X1 U32570 ( .A(n2467), .B(n4075), .S(n2859), .Z(n3792) );
  NAND2_X1 U32580 ( .A1(n2469), .A2(n2468), .ZN(n2470) );
  NAND2_X1 U32590 ( .A1(n2480), .A2(n2470), .ZN(n3796) );
  OR2_X1 U32600 ( .A1(n3796), .A2(n2353), .ZN(n2475) );
  OR2_X1 U32610 ( .A1(n2347), .A2(n4624), .ZN(n2472) );
  INV_X1 U32620 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4481) );
  OR2_X1 U32630 ( .A1(n2346), .A2(n4481), .ZN(n2471) );
  AND2_X1 U32640 ( .A1(n2472), .A2(n2471), .ZN(n2474) );
  INV_X1 U32650 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3453) );
  OR2_X1 U32660 ( .A1(n3510), .A2(n3453), .ZN(n2473) );
  NAND2_X1 U32670 ( .A1(n2477), .A2(IR_REG_31__SCAN_IN), .ZN(n2476) );
  MUX2_X1 U32680 ( .A(IR_REG_31__SCAN_IN), .B(n2476), .S(IR_REG_14__SCAN_IN), 
        .Z(n2478) );
  NAND2_X1 U32690 ( .A1(n2478), .A2(n2485), .ZN(n4086) );
  INV_X1 U32700 ( .A(DATAI_14_), .ZN(n2479) );
  MUX2_X1 U32710 ( .A(n4086), .B(n2479), .S(n3506), .Z(n4470) );
  INV_X1 U32720 ( .A(n4470), .ZN(n3700) );
  NAND2_X1 U32730 ( .A1(n2480), .A2(n4608), .ZN(n2481) );
  AND2_X1 U32740 ( .A1(n2492), .A2(n2481), .ZN(n3704) );
  NAND2_X1 U32750 ( .A1(n3704), .A2(n2685), .ZN(n2484) );
  AOI22_X1 U32760 ( .A1(n2758), .A2(REG0_REG_14__SCAN_IN), .B1(n2345), .B2(
        REG1_REG_14__SCAN_IN), .ZN(n2483) );
  NAND2_X1 U32770 ( .A1(n2614), .A2(REG2_REG_14__SCAN_IN), .ZN(n2482) );
  NAND2_X1 U32780 ( .A1(n3700), .A2(n4368), .ZN(n3891) );
  INV_X1 U32790 ( .A(n4368), .ZN(n4455) );
  NAND2_X1 U32800 ( .A1(n4470), .A2(n4455), .ZN(n3878) );
  NAND2_X1 U32810 ( .A1(n3891), .A2(n3878), .ZN(n3405) );
  NAND2_X1 U32820 ( .A1(n2486), .A2(IR_REG_15__SCAN_IN), .ZN(n2489) );
  INV_X1 U32830 ( .A(DATAI_15_), .ZN(n2490) );
  MUX2_X1 U32840 ( .A(n4100), .B(n2490), .S(n3506), .Z(n4459) );
  INV_X1 U32850 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3489) );
  NAND2_X1 U32860 ( .A1(n2492), .A2(n2145), .ZN(n2493) );
  NAND2_X1 U32870 ( .A1(n2501), .A2(n2493), .ZN(n4365) );
  OR2_X1 U32880 ( .A1(n4365), .A2(n2353), .ZN(n2495) );
  AOI22_X1 U32890 ( .A1(n2758), .A2(REG0_REG_15__SCAN_IN), .B1(n2345), .B2(
        REG1_REG_15__SCAN_IN), .ZN(n2494) );
  NAND2_X1 U32900 ( .A1(n4361), .A2(n4467), .ZN(n2496) );
  NAND2_X1 U32910 ( .A1(n2497), .A2(IR_REG_31__SCAN_IN), .ZN(n2499) );
  INV_X1 U32920 ( .A(IR_REG_16__SCAN_IN), .ZN(n2498) );
  INV_X1 U32930 ( .A(DATAI_16_), .ZN(n2500) );
  MUX2_X1 U32940 ( .A(n4106), .B(n2500), .S(n3506), .Z(n4449) );
  NAND2_X1 U32950 ( .A1(n2501), .A2(n2146), .ZN(n2502) );
  NAND2_X1 U32960 ( .A1(n2511), .A2(n2502), .ZN(n4346) );
  OR2_X1 U32970 ( .A1(n4346), .A2(n2353), .ZN(n2508) );
  INV_X1 U32980 ( .A(REG2_REG_16__SCAN_IN), .ZN(n2505) );
  NAND2_X1 U32990 ( .A1(n2758), .A2(REG0_REG_16__SCAN_IN), .ZN(n2504) );
  NAND2_X1 U33000 ( .A1(n2345), .A2(REG1_REG_16__SCAN_IN), .ZN(n2503) );
  OAI211_X1 U33010 ( .C1(n2505), .C2(n3510), .A(n2504), .B(n2503), .ZN(n2506)
         );
  INV_X1 U33020 ( .A(n2506), .ZN(n2507) );
  NAND2_X1 U33030 ( .A1(n4449), .A2(n4456), .ZN(n3871) );
  INV_X1 U33040 ( .A(n4456), .ZN(n4372) );
  NAND2_X1 U33050 ( .A1(n4345), .A2(n4372), .ZN(n3979) );
  NAND2_X1 U33060 ( .A1(n4345), .A2(n4456), .ZN(n2510) );
  NAND2_X1 U33070 ( .A1(n2511), .A2(n4651), .ZN(n2512) );
  AND2_X1 U33080 ( .A1(n2532), .A2(n2512), .ZN(n4330) );
  NAND2_X1 U33090 ( .A1(n4330), .A2(n2685), .ZN(n2519) );
  INV_X1 U33100 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2516) );
  NAND2_X1 U33110 ( .A1(n2758), .A2(REG0_REG_17__SCAN_IN), .ZN(n2515) );
  INV_X1 U33120 ( .A(REG1_REG_17__SCAN_IN), .ZN(n2513) );
  OR2_X1 U33130 ( .A1(n2346), .A2(n2513), .ZN(n2514) );
  OAI211_X1 U33140 ( .C1(n2516), .C2(n3510), .A(n2515), .B(n2514), .ZN(n2517)
         );
  INV_X1 U33150 ( .A(n2517), .ZN(n2518) );
  NOR2_X1 U33160 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2522) );
  NOR2_X1 U33170 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2521) );
  AND4_X1 U33180 ( .A1(n2523), .A2(n2522), .A3(n2521), .A4(n2520), .ZN(n2525)
         );
  AND2_X1 U33190 ( .A1(n2525), .A2(n2524), .ZN(n2526) );
  OR2_X1 U33200 ( .A1(n2540), .A2(n2637), .ZN(n2527) );
  XNOR2_X1 U33210 ( .A(n2527), .B(IR_REG_17__SCAN_IN), .ZN(n3495) );
  MUX2_X1 U33220 ( .A(n3495), .B(DATAI_17_), .S(n3506), .Z(n4436) );
  NAND2_X1 U33230 ( .A1(n3751), .A2(n4329), .ZN(n2529) );
  AND2_X1 U33240 ( .A1(n4447), .A2(n4436), .ZN(n2528) );
  INV_X1 U33250 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U33260 ( .A1(n2532), .A2(n2531), .ZN(n2533) );
  NAND2_X1 U33270 ( .A1(n2544), .A2(n2533), .ZN(n4318) );
  OR2_X1 U33280 ( .A1(n4318), .A2(n2353), .ZN(n2538) );
  INV_X1 U33290 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3475) );
  NAND2_X1 U33300 ( .A1(n2758), .A2(REG0_REG_18__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U33310 ( .A1(n2614), .A2(REG2_REG_18__SCAN_IN), .ZN(n2534) );
  OAI211_X1 U33320 ( .C1(n2346), .C2(n3475), .A(n2535), .B(n2534), .ZN(n2536)
         );
  INV_X1 U33330 ( .A(n2536), .ZN(n2537) );
  NAND2_X1 U33340 ( .A1(n2540), .A2(n2539), .ZN(n2551) );
  NAND2_X1 U33350 ( .A1(n2551), .A2(IR_REG_31__SCAN_IN), .ZN(n2541) );
  XNOR2_X1 U33360 ( .A(n2541), .B(IR_REG_18__SCAN_IN), .ZN(n3496) );
  MUX2_X1 U33370 ( .A(DATAI_18_), .B(n3496), .S(n2859), .Z(n4311) );
  NAND2_X1 U33380 ( .A1(n4440), .A2(n4311), .ZN(n4283) );
  NAND2_X1 U33390 ( .A1(n4289), .A2(n4308), .ZN(n4284) );
  NAND2_X1 U33400 ( .A1(n4283), .A2(n4284), .ZN(n4304) );
  NAND2_X1 U33410 ( .A1(n4440), .A2(n4308), .ZN(n2542) );
  INV_X1 U33420 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2543) );
  NAND2_X1 U33430 ( .A1(n2544), .A2(n2543), .ZN(n2545) );
  AND2_X1 U33440 ( .A1(n2555), .A2(n2545), .ZN(n4298) );
  NAND2_X1 U33450 ( .A1(n4298), .A2(n2685), .ZN(n2550) );
  INV_X1 U33460 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4561) );
  NAND2_X1 U33470 ( .A1(n2758), .A2(REG0_REG_19__SCAN_IN), .ZN(n2547) );
  NAND2_X1 U33480 ( .A1(n2345), .A2(REG1_REG_19__SCAN_IN), .ZN(n2546) );
  OAI211_X1 U33490 ( .C1(n4561), .C2(n3510), .A(n2547), .B(n2546), .ZN(n2548)
         );
  INV_X1 U33500 ( .A(n2548), .ZN(n2549) );
  INV_X1 U33510 ( .A(n2551), .ZN(n2552) );
  NAND2_X1 U33520 ( .A1(n2552), .A2(n4563), .ZN(n2635) );
  NAND2_X1 U3353 ( .A1(n2635), .A2(IR_REG_31__SCAN_IN), .ZN(n2553) );
  XNOR2_X1 U33540 ( .A(n2553), .B(IR_REG_19__SCAN_IN), .ZN(n2953) );
  MUX2_X1 U3355 ( .A(DATAI_19_), .B(n4316), .S(n2859), .Z(n4288) );
  NAND2_X1 U3356 ( .A1(n4421), .A2(n4288), .ZN(n2554) );
  INV_X1 U3357 ( .A(n4288), .ZN(n4296) );
  INV_X1 U3358 ( .A(REG3_REG_20__SCAN_IN), .ZN(n3782) );
  NAND2_X1 U3359 ( .A1(n2555), .A2(n3782), .ZN(n2556) );
  NAND2_X1 U3360 ( .A1(n2573), .A2(n2556), .ZN(n3781) );
  INV_X1 U3361 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4582) );
  NAND2_X1 U3362 ( .A1(n2614), .A2(REG2_REG_20__SCAN_IN), .ZN(n2558) );
  NAND2_X1 U3363 ( .A1(n2345), .A2(REG1_REG_20__SCAN_IN), .ZN(n2557) );
  OAI211_X1 U3364 ( .C1(n2347), .C2(n4582), .A(n2558), .B(n2557), .ZN(n2559)
         );
  INV_X1 U3365 ( .A(n2559), .ZN(n2560) );
  NOR2_X1 U3366 ( .A1(n4411), .A2(n4420), .ZN(n2563) );
  NAND2_X1 U3367 ( .A1(n4411), .A2(n4420), .ZN(n2562) );
  XNOR2_X1 U3368 ( .A(n2573), .B(REG3_REG_21__SCAN_IN), .ZN(n4253) );
  NAND2_X1 U3369 ( .A1(n4253), .A2(n2685), .ZN(n2569) );
  INV_X1 U3370 ( .A(REG2_REG_21__SCAN_IN), .ZN(n2566) );
  NAND2_X1 U3371 ( .A1(n2758), .A2(REG0_REG_21__SCAN_IN), .ZN(n2565) );
  NAND2_X1 U3372 ( .A1(n2345), .A2(REG1_REG_21__SCAN_IN), .ZN(n2564) );
  OAI211_X1 U3373 ( .C1(n2566), .C2(n3510), .A(n2565), .B(n2564), .ZN(n2567)
         );
  INV_X1 U3374 ( .A(n2567), .ZN(n2568) );
  AND2_X1 U3375 ( .A1(n3506), .A2(DATAI_21_), .ZN(n4410) );
  AND2_X1 U3376 ( .A1(n4230), .A2(n4410), .ZN(n2571) );
  INV_X1 U3377 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3727) );
  INV_X1 U3378 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3593) );
  OAI21_X1 U3379 ( .B1(n2573), .B2(n3727), .A(n3593), .ZN(n2574) );
  NAND2_X1 U3380 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2572) );
  NAND2_X1 U3381 ( .A1(n2574), .A2(n2581), .ZN(n4242) );
  INV_X1 U3382 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4659) );
  NAND2_X1 U3383 ( .A1(n2758), .A2(REG0_REG_22__SCAN_IN), .ZN(n2576) );
  NAND2_X1 U3384 ( .A1(n2614), .A2(REG2_REG_22__SCAN_IN), .ZN(n2575) );
  OAI211_X1 U3385 ( .C1(n2346), .C2(n4659), .A(n2576), .B(n2575), .ZN(n2577)
         );
  INV_X1 U3386 ( .A(n2577), .ZN(n2578) );
  AND2_X1 U3387 ( .A1(n3506), .A2(DATAI_22_), .ZN(n4229) );
  NAND2_X1 U3388 ( .A1(n4414), .A2(n4229), .ZN(n4205) );
  NAND2_X1 U3389 ( .A1(n4211), .A2(n4241), .ZN(n2678) );
  INV_X1 U3390 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4663) );
  NAND2_X1 U3391 ( .A1(n2581), .A2(n4663), .ZN(n2582) );
  NAND2_X1 U3392 ( .A1(n2599), .A2(n2582), .ZN(n4217) );
  INV_X1 U3393 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4218) );
  NAND2_X1 U3394 ( .A1(n2758), .A2(REG0_REG_23__SCAN_IN), .ZN(n2584) );
  NAND2_X1 U3395 ( .A1(n2345), .A2(REG1_REG_23__SCAN_IN), .ZN(n2583) );
  OAI211_X1 U3396 ( .C1(n4218), .C2(n3510), .A(n2584), .B(n2583), .ZN(n2585)
         );
  INV_X1 U3397 ( .A(n2585), .ZN(n2586) );
  NAND2_X1 U3398 ( .A1(n3506), .A2(DATAI_23_), .ZN(n4215) );
  NAND2_X1 U3399 ( .A1(n4233), .A2(n4215), .ZN(n2588) );
  NAND2_X1 U3400 ( .A1(n4203), .A2(n2588), .ZN(n2590) );
  INV_X1 U3401 ( .A(n4215), .ZN(n4210) );
  NAND2_X1 U3402 ( .A1(n4393), .A2(n4210), .ZN(n2589) );
  XNOR2_X1 U3403 ( .A(n2599), .B(REG3_REG_24__SCAN_IN), .ZN(n4195) );
  NAND2_X1 U3404 ( .A1(n4195), .A2(n2685), .ZN(n2596) );
  INV_X1 U3405 ( .A(REG2_REG_24__SCAN_IN), .ZN(n2593) );
  NAND2_X1 U3406 ( .A1(n2758), .A2(REG0_REG_24__SCAN_IN), .ZN(n2592) );
  NAND2_X1 U3407 ( .A1(n2345), .A2(REG1_REG_24__SCAN_IN), .ZN(n2591) );
  OAI211_X1 U3408 ( .C1(n2593), .C2(n3510), .A(n2592), .B(n2591), .ZN(n2594)
         );
  INV_X1 U3409 ( .A(n2594), .ZN(n2595) );
  AND2_X1 U3410 ( .A1(n3506), .A2(DATAI_24_), .ZN(n4392) );
  AND2_X1 U3411 ( .A1(n4016), .A2(n4392), .ZN(n2598) );
  INV_X1 U3412 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3770) );
  INV_X1 U3413 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3625) );
  OAI21_X1 U3414 ( .B1(n2599), .B2(n3770), .A(n3625), .ZN(n2600) );
  NAND2_X1 U3415 ( .A1(n2600), .A2(n2607), .ZN(n3624) );
  INV_X1 U3416 ( .A(REG2_REG_25__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U3417 ( .A1(n2758), .A2(REG0_REG_25__SCAN_IN), .ZN(n2602) );
  NAND2_X1 U3418 ( .A1(n2345), .A2(REG1_REG_25__SCAN_IN), .ZN(n2601) );
  OAI211_X1 U3419 ( .C1(n2603), .C2(n3510), .A(n2602), .B(n2601), .ZN(n2604)
         );
  INV_X1 U3420 ( .A(n2604), .ZN(n2605) );
  AND2_X1 U3421 ( .A1(n3506), .A2(DATAI_25_), .ZN(n4382) );
  NOR2_X1 U3422 ( .A1(n3824), .A2(n4382), .ZN(n2737) );
  INV_X1 U3423 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4647) );
  NAND2_X1 U3424 ( .A1(n2607), .A2(n4647), .ZN(n2608) );
  NAND2_X1 U3425 ( .A1(n4163), .A2(n2685), .ZN(n2613) );
  INV_X1 U3426 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4634) );
  NAND2_X1 U3427 ( .A1(n2614), .A2(REG2_REG_26__SCAN_IN), .ZN(n2610) );
  NAND2_X1 U3428 ( .A1(n2345), .A2(REG1_REG_26__SCAN_IN), .ZN(n2609) );
  OAI211_X1 U3429 ( .C1(n2347), .C2(n4634), .A(n2610), .B(n2609), .ZN(n2611)
         );
  INV_X1 U3430 ( .A(n2611), .ZN(n2612) );
  AND2_X1 U3431 ( .A1(n3506), .A2(DATAI_26_), .ZN(n2743) );
  OR2_X1 U3432 ( .A1(n2737), .A2(n2622), .ZN(n2792) );
  NAND2_X1 U3433 ( .A1(n4152), .A2(n2685), .ZN(n2619) );
  INV_X1 U3434 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2799) );
  NAND2_X1 U3435 ( .A1(n2758), .A2(REG0_REG_27__SCAN_IN), .ZN(n2616) );
  NAND2_X1 U3436 ( .A1(n2614), .A2(REG2_REG_27__SCAN_IN), .ZN(n2615) );
  OAI211_X1 U3437 ( .C1(n2346), .C2(n2799), .A(n2616), .B(n2615), .ZN(n2617)
         );
  INV_X1 U3438 ( .A(n2617), .ZN(n2618) );
  AND2_X1 U3439 ( .A1(n3506), .A2(DATAI_27_), .ZN(n2800) );
  NOR2_X1 U3440 ( .A1(n4015), .A2(n2800), .ZN(n2623) );
  OR2_X1 U3441 ( .A1(n2792), .A2(n2623), .ZN(n2620) );
  NAND2_X1 U3442 ( .A1(n3824), .A2(n4382), .ZN(n2738) );
  AND2_X1 U3443 ( .A1(n2039), .A2(n2738), .ZN(n2621) );
  OR2_X1 U3444 ( .A1(n2623), .A2(n2793), .ZN(n2625) );
  NAND2_X1 U3445 ( .A1(n4015), .A2(n2800), .ZN(n2624) );
  NAND2_X1 U3446 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .ZN(
        n2626) );
  INV_X1 U3447 ( .A(n2686), .ZN(n4128) );
  INV_X1 U3448 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3685) );
  INV_X1 U3449 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2627) );
  OAI21_X1 U3450 ( .B1(n2628), .B2(n3685), .A(n2627), .ZN(n2629) );
  NAND2_X1 U3451 ( .A1(n4128), .A2(n2629), .ZN(n4138) );
  INV_X1 U3452 ( .A(REG2_REG_28__SCAN_IN), .ZN(n4137) );
  NAND2_X1 U3453 ( .A1(n2758), .A2(REG0_REG_28__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U3454 ( .A1(n2345), .A2(REG1_REG_28__SCAN_IN), .ZN(n2630) );
  OAI211_X1 U3455 ( .C1(n4137), .C2(n3510), .A(n2631), .B(n2630), .ZN(n2632)
         );
  INV_X1 U3456 ( .A(n2632), .ZN(n2633) );
  AND2_X1 U3457 ( .A1(n3506), .A2(DATAI_28_), .ZN(n3670) );
  INV_X1 U34580 ( .A(n3670), .ZN(n4139) );
  NAND2_X1 U34590 ( .A1(n4014), .A2(n4139), .ZN(n3905) );
  NAND2_X1 U3460 ( .A1(n3912), .A2(n3905), .ZN(n3964) );
  XNOR2_X1 U3461 ( .A(n2774), .B(n3964), .ZN(n4135) );
  NAND3_X1 U3462 ( .A1(n2635), .A2(IR_REG_31__SCAN_IN), .A3(IR_REG_20__SCAN_IN), .ZN(n2644) );
  AND2_X1 U3463 ( .A1(n2637), .A2(IR_REG_20__SCAN_IN), .ZN(n2640) );
  NAND2_X1 U3464 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2638) );
  XNOR2_X2 U3465 ( .A(n2647), .B(n2646), .ZN(n2705) );
  NAND2_X2 U3466 ( .A1(n2728), .A2(n4687), .ZN(n2964) );
  INV_X1 U34670 ( .A(n2648), .ZN(n2653) );
  NOR2_X1 U3468 ( .A1(n2649), .A2(IR_REG_21__SCAN_IN), .ZN(n2651) );
  AND2_X1 U34690 ( .A1(n2651), .A2(n2650), .ZN(n2652) );
  NAND2_X1 U3470 ( .A1(n2653), .A2(n2652), .ZN(n2695) );
  NAND2_X1 U34710 ( .A1(n2695), .A2(IR_REG_31__SCAN_IN), .ZN(n2655) );
  INV_X1 U3472 ( .A(IR_REG_22__SCAN_IN), .ZN(n2654) );
  INV_X1 U34730 ( .A(n4004), .ZN(n2847) );
  XNOR2_X1 U3474 ( .A(n2964), .B(n2847), .ZN(n2656) );
  NAND2_X1 U34750 ( .A1(n2656), .A2(n3501), .ZN(n3220) );
  AND2_X1 U3476 ( .A1(n4316), .A2(n2728), .ZN(n4750) );
  INV_X1 U34770 ( .A(n4776), .ZN(n3070) );
  INV_X1 U3478 ( .A(n4015), .ZN(n4140) );
  NAND2_X1 U34790 ( .A1(n2657), .A2(IR_REG_31__SCAN_IN), .ZN(n2658) );
  XNOR2_X1 U3480 ( .A(n2658), .B(n2316), .ZN(n4699) );
  INV_X1 U34810 ( .A(n4699), .ZN(n2989) );
  INV_X1 U3482 ( .A(n4485), .ZN(n4386) );
  NAND2_X1 U34830 ( .A1(n2928), .A2(n2997), .ZN(n3847) );
  NAND2_X1 U3484 ( .A1(n2809), .A2(n3850), .ZN(n2834) );
  NAND2_X1 U34850 ( .A1(n2834), .A2(n3933), .ZN(n2833) );
  NAND2_X1 U3486 ( .A1(n2833), .A2(n3851), .ZN(n3064) );
  NAND2_X1 U34870 ( .A1(n3132), .A2(n3072), .ZN(n3856) );
  NAND2_X1 U3488 ( .A1(n4024), .A2(n3135), .ZN(n3853) );
  NAND2_X1 U34890 ( .A1(n3064), .A2(n3939), .ZN(n3063) );
  AND2_X1 U3490 ( .A1(n4022), .A2(n3246), .ZN(n3024) );
  NAND2_X1 U34910 ( .A1(n3160), .A2(n3029), .ZN(n3873) );
  NAND2_X1 U3492 ( .A1(n4021), .A2(n3177), .ZN(n3875) );
  NAND2_X1 U34930 ( .A1(n3248), .A2(n3301), .ZN(n3861) );
  NAND2_X1 U3494 ( .A1(n2665), .A2(n3872), .ZN(n3182) );
  NAND2_X1 U34950 ( .A1(n3341), .A2(n3289), .ZN(n3864) );
  NAND2_X1 U3496 ( .A1(n4019), .A2(n3284), .ZN(n3876) );
  NAND2_X1 U34970 ( .A1(n3338), .A2(n3266), .ZN(n3865) );
  NAND2_X1 U3498 ( .A1(n3806), .A2(n3397), .ZN(n3886) );
  NAND2_X1 U34990 ( .A1(n3427), .A2(n2667), .ZN(n3883) );
  NAND2_X1 U3500 ( .A1(n4490), .A2(n4017), .ZN(n3441) );
  NAND2_X1 U35010 ( .A1(n3792), .A2(n4487), .ZN(n2668) );
  NAND2_X1 U3502 ( .A1(n3441), .A2(n2668), .ZN(n3887) );
  INV_X1 U35030 ( .A(n3351), .ZN(n3889) );
  INV_X1 U3504 ( .A(n3887), .ZN(n2671) );
  NAND2_X1 U35050 ( .A1(n3736), .A2(n3802), .ZN(n3443) );
  NAND2_X1 U35060 ( .A1(n3443), .A2(n3349), .ZN(n2670) );
  NOR2_X1 U35070 ( .A1(n3792), .A2(n4487), .ZN(n2669) );
  AOI21_X1 U35080 ( .B1(n2671), .B2(n2670), .A(n2669), .ZN(n3893) );
  NAND2_X1 U35090 ( .A1(n2672), .A2(n3893), .ZN(n3403) );
  INV_X1 U35100 ( .A(n3405), .ZN(n3929) );
  NAND2_X1 U35110 ( .A1(n4361), .A2(n4350), .ZN(n3892) );
  NAND2_X1 U35120 ( .A1(n4459), .A2(n4467), .ZN(n3879) );
  NAND2_X1 U35130 ( .A1(n3892), .A2(n3879), .ZN(n4357) );
  NAND2_X1 U35140 ( .A1(n4421), .A2(n4296), .ZN(n3926) );
  NAND2_X1 U35150 ( .A1(n3926), .A2(n4284), .ZN(n3868) );
  NOR2_X1 U35160 ( .A1(n4282), .A2(n3868), .ZN(n2674) );
  INV_X1 U35170 ( .A(n4420), .ZN(n4275) );
  NAND2_X1 U35180 ( .A1(n4411), .A2(n4275), .ZN(n3869) );
  NAND2_X1 U35190 ( .A1(n3751), .A2(n4436), .ZN(n4281) );
  AND2_X1 U35200 ( .A1(n4283), .A2(n4281), .ZN(n2675) );
  OR2_X1 U35210 ( .A1(n2675), .A2(n3868), .ZN(n2676) );
  NAND2_X1 U35220 ( .A1(n4313), .A2(n4288), .ZN(n3927) );
  NAND2_X1 U35230 ( .A1(n2676), .A2(n3927), .ZN(n4263) );
  NOR2_X1 U35240 ( .A1(n4411), .A2(n4275), .ZN(n2677) );
  OAI21_X1 U35250 ( .B1(n4263), .B2(n2677), .A(n3869), .ZN(n3977) );
  OR2_X1 U35260 ( .A1(n4230), .A2(n4255), .ZN(n4223) );
  NAND2_X1 U35270 ( .A1(n4205), .A2(n4223), .ZN(n3976) );
  NAND2_X1 U35280 ( .A1(n4393), .A2(n4215), .ZN(n3923) );
  NAND2_X1 U35290 ( .A1(n3923), .A2(n2678), .ZN(n3903) );
  AND2_X1 U35300 ( .A1(n4230), .A2(n4255), .ZN(n3899) );
  AND2_X1 U35310 ( .A1(n4205), .A2(n3899), .ZN(n2679) );
  NOR2_X1 U35320 ( .A1(n3903), .A2(n2679), .ZN(n3981) );
  NOR2_X1 U35330 ( .A1(n4393), .A2(n4215), .ZN(n3925) );
  INV_X1 U35340 ( .A(n4392), .ZN(n4197) );
  NAND2_X1 U35350 ( .A1(n4183), .A2(n2743), .ZN(n2680) );
  INV_X1 U35360 ( .A(n4382), .ZN(n4182) );
  NAND2_X1 U35370 ( .A1(n2680), .A2(n3921), .ZN(n3988) );
  INV_X1 U35380 ( .A(n3988), .ZN(n3902) );
  NAND2_X1 U35390 ( .A1(n3824), .A2(n4182), .ZN(n3920) );
  NAND2_X1 U35400 ( .A1(n4016), .A2(n4197), .ZN(n4170) );
  AND2_X1 U35410 ( .A1(n3920), .A2(n4170), .ZN(n2740) );
  NAND2_X1 U35420 ( .A1(n4383), .A2(n3827), .ZN(n3969) );
  OAI21_X1 U35430 ( .B1(n3988), .B2(n2740), .A(n3969), .ZN(n3907) );
  XNOR2_X1 U35440 ( .A(n4015), .B(n2800), .ZN(n3970) );
  INV_X1 U35450 ( .A(n2800), .ZN(n4154) );
  OR2_X1 U35460 ( .A1(n4015), .A2(n4154), .ZN(n3911) );
  INV_X1 U35470 ( .A(n3964), .ZN(n2681) );
  XNOR2_X1 U35480 ( .A(n2753), .B(n2681), .ZN(n2684) );
  NAND2_X1 U35490 ( .A1(n4316), .A2(n2847), .ZN(n2683) );
  INV_X1 U35500 ( .A(n2728), .ZN(n4000) );
  NAND2_X1 U35510 ( .A1(n4000), .A2(n4687), .ZN(n2682) );
  NAND2_X1 U35520 ( .A1(n2686), .A2(n2685), .ZN(n2692) );
  INV_X1 U35530 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2689) );
  NAND2_X1 U35540 ( .A1(n2758), .A2(REG0_REG_29__SCAN_IN), .ZN(n2688) );
  NAND2_X1 U35550 ( .A1(n2345), .A2(REG1_REG_29__SCAN_IN), .ZN(n2687) );
  OAI211_X1 U35560 ( .C1(n2689), .C2(n3510), .A(n2688), .B(n2687), .ZN(n2690)
         );
  INV_X1 U35570 ( .A(n2690), .ZN(n2691) );
  NAND2_X1 U35580 ( .A1(n2955), .A2(n4699), .ZN(n4439) );
  INV_X1 U35590 ( .A(n4439), .ZN(n4486) );
  NAND2_X1 U35600 ( .A1(n4004), .A2(n2705), .ZN(n2727) );
  NOR2_X1 U35610 ( .A1(n2728), .A2(n2727), .ZN(n4409) );
  AOI22_X1 U35620 ( .A1(n4143), .A2(n4486), .B1(n4437), .B2(n3670), .ZN(n2693)
         );
  OAI211_X1 U35630 ( .C1(n4140), .C2(n4386), .A(n4136), .B(n2693), .ZN(n2694)
         );
  NAND2_X1 U35640 ( .A1(n2709), .A2(n2711), .ZN(n2710) );
  XNOR2_X2 U35650 ( .A(n2696), .B(IR_REG_24__SCAN_IN), .ZN(n2707) );
  INV_X1 U35660 ( .A(IR_REG_25__SCAN_IN), .ZN(n2698) );
  NAND2_X1 U35670 ( .A1(n2697), .A2(n2706), .ZN(n2700) );
  MUX2_X1 U35680 ( .A(n2697), .B(n2700), .S(B_REG_SCAN_IN), .Z(n2704) );
  INV_X1 U35690 ( .A(n2701), .ZN(n2702) );
  XNOR2_X2 U35700 ( .A(n2703), .B(IR_REG_26__SCAN_IN), .ZN(n2708) );
  INV_X1 U35710 ( .A(D_REG_1__SCAN_IN), .ZN(n2819) );
  NAND2_X1 U35720 ( .A1(n2817), .A2(n2819), .ZN(n2950) );
  INV_X1 U35730 ( .A(n2708), .ZN(n2723) );
  NAND2_X1 U35740 ( .A1(n2723), .A2(n2706), .ZN(n2857) );
  NAND2_X1 U35750 ( .A1(n2950), .A2(n2857), .ZN(n2722) );
  NAND2_X1 U35760 ( .A1(n4776), .A2(n2705), .ZN(n2822) );
  INV_X1 U35770 ( .A(n2706), .ZN(n2844) );
  OAI21_X1 U35780 ( .B1(n2709), .B2(n2711), .A(n2710), .ZN(n3122) );
  NAND2_X1 U35790 ( .A1(n3501), .A2(n2728), .ZN(n2957) );
  NAND2_X1 U35800 ( .A1(n2957), .A2(n2955), .ZN(n2960) );
  AND3_X1 U35810 ( .A1(n2822), .A2(n2982), .A3(n2960), .ZN(n2721) );
  NOR4_X1 U3582 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_21__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n2715) );
  NOR4_X1 U3583 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_8__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2714) );
  NOR4_X1 U3584 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_30__SCAN_IN), .ZN(n2713) );
  NOR4_X1 U3585 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2712) );
  NAND4_X1 U3586 ( .A1(n2715), .A2(n2714), .A3(n2713), .A4(n2712), .ZN(n2720)
         );
  INV_X1 U3587 ( .A(D_REG_11__SCAN_IN), .ZN(n4760) );
  INV_X1 U3588 ( .A(D_REG_22__SCAN_IN), .ZN(n4757) );
  INV_X1 U3589 ( .A(D_REG_6__SCAN_IN), .ZN(n4763) );
  INV_X1 U3590 ( .A(D_REG_9__SCAN_IN), .ZN(n4762) );
  NAND4_X1 U3591 ( .A1(n4760), .A2(n4757), .A3(n4763), .A4(n4762), .ZN(n2716)
         );
  NOR4_X1 U3592 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        D_REG_27__SCAN_IN), .A4(n2716), .ZN(n4551) );
  NOR4_X1 U3593 ( .A1(D_REG_4__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2718) );
  NOR3_X1 U3594 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_19__SCAN_IN), .ZN(n2717) );
  NAND3_X1 U3595 ( .A1(n4551), .A2(n2718), .A3(n2717), .ZN(n2719) );
  OAI21_X1 U3596 ( .B1(n2720), .B2(n2719), .A(n2817), .ZN(n2816) );
  NAND3_X1 U3597 ( .A1(n2722), .A2(n2721), .A3(n2816), .ZN(n2732) );
  INV_X1 U3598 ( .A(D_REG_0__SCAN_IN), .ZN(n3460) );
  NAND2_X1 U3599 ( .A1(n2817), .A2(n3460), .ZN(n2725) );
  NAND2_X1 U3600 ( .A1(n2697), .A2(n2723), .ZN(n2724) );
  NAND2_X1 U3601 ( .A1(n2975), .A2(n2929), .ZN(n3074) );
  NOR2_X4 U3602 ( .A1(n3198), .A2(n3289), .ZN(n3271) );
  INV_X1 U3603 ( .A(n2802), .ZN(n2726) );
  INV_X1 U3604 ( .A(n2778), .ZN(n2780) );
  INV_X1 U3605 ( .A(n2727), .ZN(n2956) );
  OR2_X1 U3606 ( .A1(n4145), .A2(n4546), .ZN(n2730) );
  NAND2_X1 U3607 ( .A1(n4782), .A2(REG0_REG_28__SCAN_IN), .ZN(n2729) );
  OAI21_X1 U3608 ( .B1(n2736), .B2(n4782), .A(n2731), .ZN(U3514) );
  NAND2_X1 U3609 ( .A1(n4784), .A2(REG1_REG_28__SCAN_IN), .ZN(n2733) );
  OAI21_X1 U3610 ( .B1(n2736), .B2(n4784), .A(n2735), .ZN(U3546) );
  INV_X1 U3611 ( .A(REG1_REG_26__SCAN_IN), .ZN(n2746) );
  XNOR2_X1 U3612 ( .A(n4383), .B(n2743), .ZN(n3965) );
  INV_X1 U3613 ( .A(n2740), .ZN(n3984) );
  OAI21_X1 U3614 ( .B1(n4172), .B2(n3984), .A(n3921), .ZN(n2741) );
  XNOR2_X1 U3615 ( .A(n2741), .B(n3965), .ZN(n2742) );
  NAND2_X1 U3616 ( .A1(n2742), .A2(n4338), .ZN(n2745) );
  AOI22_X1 U3617 ( .A1(n3824), .A2(n4485), .B1(n2743), .B2(n4409), .ZN(n2744)
         );
  OAI211_X1 U3618 ( .C1(n4140), .C2(n4439), .A(n2745), .B(n2744), .ZN(n4167)
         );
  AOI21_X1 U3619 ( .B1(n4162), .B2(n4480), .A(n4167), .ZN(n2750) );
  MUX2_X1 U3620 ( .A(n2746), .B(n2750), .S(n4787), .Z(n2749) );
  OAI21_X1 U3621 ( .B1(n4177), .B2(n3827), .A(n2747), .ZN(n4165) );
  NAND2_X1 U3622 ( .A1(n2749), .A2(n2748), .ZN(U3544) );
  MUX2_X1 U3623 ( .A(n4634), .B(n2750), .S(n4783), .Z(n2752) );
  NAND2_X1 U3624 ( .A1(n2752), .A2(n2751), .ZN(U3512) );
  AND2_X1 U3625 ( .A1(n3506), .A2(DATAI_29_), .ZN(n2779) );
  XNOR2_X1 U3626 ( .A(n2754), .B(n3966), .ZN(n2765) );
  NAND2_X1 U3627 ( .A1(n4014), .A2(n4485), .ZN(n2763) );
  OAI21_X1 U3628 ( .B1(n2755), .B2(IR_REG_26__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2756) );
  XNOR2_X1 U3629 ( .A(n2756), .B(IR_REG_27__SCAN_IN), .ZN(n4705) );
  AND2_X1 U3630 ( .A1(n4705), .A2(B_REG_SCAN_IN), .ZN(n2757) );
  NOR2_X1 U3631 ( .A1(n4439), .A2(n2757), .ZN(n3511) );
  INV_X1 U3632 ( .A(REG2_REG_30__SCAN_IN), .ZN(n2761) );
  NAND2_X1 U3633 ( .A1(n2345), .A2(REG1_REG_30__SCAN_IN), .ZN(n2760) );
  NAND2_X1 U3634 ( .A1(n2758), .A2(REG0_REG_30__SCAN_IN), .ZN(n2759) );
  OAI211_X1 U3635 ( .C1(n3510), .C2(n2761), .A(n2760), .B(n2759), .ZN(n4013)
         );
  AOI22_X1 U3636 ( .A1(n3511), .A2(n4013), .B1(n4409), .B2(n2779), .ZN(n2762)
         );
  NAND2_X1 U3637 ( .A1(n2763), .A2(n2762), .ZN(n2764) );
  AOI21_X1 U3638 ( .B1(n2765), .B2(n4338), .A(n2764), .ZN(n4127) );
  NAND2_X1 U3639 ( .A1(n2767), .A2(n2766), .ZN(n2768) );
  NAND2_X1 U3640 ( .A1(n2768), .A2(n3964), .ZN(n4124) );
  NAND2_X1 U3641 ( .A1(n4014), .A2(n3670), .ZN(n4123) );
  AND2_X1 U3642 ( .A1(n3966), .A2(n4123), .ZN(n2773) );
  INV_X1 U3643 ( .A(n2773), .ZN(n2771) );
  INV_X1 U3644 ( .A(n3966), .ZN(n4125) );
  INV_X1 U3645 ( .A(n4123), .ZN(n2769) );
  AOI21_X1 U3646 ( .B1(n4125), .B2(n2769), .A(n4497), .ZN(n2770) );
  OAI21_X1 U3647 ( .B1(n3964), .B2(n2771), .A(n2770), .ZN(n2772) );
  INV_X1 U3648 ( .A(n2772), .ZN(n2776) );
  NAND2_X1 U3649 ( .A1(n2774), .A2(n2773), .ZN(n2775) );
  OAI211_X1 U3650 ( .C1(n4124), .C2(n3966), .A(n2776), .B(n2775), .ZN(n2777)
         );
  INV_X1 U3651 ( .A(n2779), .ZN(n3914) );
  NAND2_X1 U3652 ( .A1(n2780), .A2(n2779), .ZN(n2781) );
  NAND2_X1 U3653 ( .A1(n2786), .A2(n2301), .ZN(U3547) );
  NAND2_X1 U3654 ( .A1(n4782), .A2(REG0_REG_29__SCAN_IN), .ZN(n2789) );
  NAND2_X1 U3655 ( .A1(n2791), .A2(n2033), .ZN(U3515) );
  XNOR2_X1 U3656 ( .A(n2794), .B(n3970), .ZN(n4150) );
  OAI21_X1 U3657 ( .B1(n3970), .B2(n2796), .A(n2795), .ZN(n2797) );
  NAND2_X1 U3658 ( .A1(n2797), .A2(n4338), .ZN(n4161) );
  AOI22_X1 U3659 ( .A1(n4383), .A2(n4485), .B1(n4409), .B2(n2800), .ZN(n2798)
         );
  NAND2_X1 U3660 ( .A1(n2747), .A2(n2800), .ZN(n2801) );
  NAND2_X1 U3661 ( .A1(n2802), .A2(n2801), .ZN(n4151) );
  INV_X1 U3662 ( .A(REG0_REG_27__SCAN_IN), .ZN(n2805) );
  MUX2_X1 U3663 ( .A(n2805), .B(n2804), .S(n4783), .Z(n2807) );
  NAND2_X1 U3664 ( .A1(n2807), .A2(n2806), .ZN(U3513) );
  INV_X1 U3665 ( .A(n4768), .ZN(n3458) );
  OR2_X1 U3666 ( .A1(n3123), .A2(n3458), .ZN(n2808) );
  INV_X1 U3667 ( .A(n2809), .ZN(n2810) );
  AOI21_X1 U3668 ( .B1(n2812), .B2(n3847), .A(n2810), .ZN(n2815) );
  OR2_X1 U3669 ( .A1(n2812), .A2(n2811), .ZN(n2813) );
  NAND2_X1 U3670 ( .A1(n2814), .A2(n2813), .ZN(n3000) );
  OAI22_X1 U3671 ( .A1(n2815), .A2(n4475), .B1(n3220), .B2(n3000), .ZN(n3002)
         );
  AND2_X1 U3672 ( .A1(n2816), .A2(n2857), .ZN(n2952) );
  INV_X1 U3673 ( .A(n2817), .ZN(n2818) );
  OAI21_X1 U3674 ( .B1(n2986), .B2(n2819), .A(n4767), .ZN(n2820) );
  NAND4_X1 U3675 ( .A1(n2821), .A2(n2952), .A3(n2820), .A4(n2960), .ZN(n2823)
         );
  MUX2_X1 U3676 ( .A(n3002), .B(REG2_REG_1__SCAN_IN), .S(n4745), .Z(n2829) );
  OAI22_X1 U3677 ( .A1(n3068), .A2(n4371), .B1(n4370), .B2(n2975), .ZN(n2828)
         );
  NAND2_X1 U3678 ( .A1(n3501), .A2(n4492), .ZN(n2824) );
  NAND2_X1 U3679 ( .A1(n3011), .A2(n2997), .ZN(n2825) );
  NAND2_X1 U3680 ( .A1(n3074), .A2(n2825), .ZN(n3082) );
  OAI22_X1 U3681 ( .A1(n2928), .A2(n4369), .B1(n4364), .B2(n3082), .ZN(n2827)
         );
  NAND2_X1 U3682 ( .A1(n2926), .A2(n4316), .ZN(n3219) );
  OR2_X1 U3683 ( .A1(n4745), .A2(n3219), .ZN(n4738) );
  OAI22_X1 U3684 ( .A1(n4738), .A2(n3000), .B1(n3014), .B2(n4755), .ZN(n2826)
         );
  OR4_X1 U3685 ( .A1(n2829), .A2(n2828), .A3(n2827), .A4(n2826), .ZN(U3289) );
  INV_X1 U3686 ( .A(n2831), .ZN(n2832) );
  AOI21_X1 U3687 ( .B1(n3933), .B2(n2830), .A(n2832), .ZN(n3016) );
  OAI21_X1 U3688 ( .B1(n3933), .B2(n2834), .A(n2833), .ZN(n2835) );
  NAND2_X1 U3689 ( .A1(n2835), .A2(n4338), .ZN(n2836) );
  OAI21_X1 U3690 ( .B1(n3016), .B2(n3220), .A(n2836), .ZN(n3018) );
  MUX2_X1 U3691 ( .A(n3018), .B(REG2_REG_2__SCAN_IN), .S(n4745), .Z(n2840) );
  OAI22_X1 U3692 ( .A1(n3132), .A2(n4371), .B1(n4370), .B2(n2967), .ZN(n2839)
         );
  XNOR2_X1 U3693 ( .A(n3074), .B(n3073), .ZN(n3085) );
  OAI22_X1 U3694 ( .A1(n2973), .A2(n4369), .B1(n4364), .B2(n3085), .ZN(n2838)
         );
  OAI22_X1 U3695 ( .A1(n4738), .A2(n3016), .B1(n2994), .B2(n4755), .ZN(n2837)
         );
  OR4_X1 U3696 ( .A1(n2840), .A2(n2839), .A3(n2838), .A4(n2837), .ZN(U3288) );
  INV_X2 U3697 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  MUX2_X1 U3698 ( .A(n4047), .B(n2374), .S(U3149), .Z(n2841) );
  INV_X1 U3699 ( .A(n2841), .ZN(U3347) );
  INV_X1 U3700 ( .A(DATAI_29_), .ZN(n2843) );
  NAND2_X1 U3701 ( .A1(n2317), .A2(STATE_REG_SCAN_IN), .ZN(n2842) );
  OAI21_X1 U3702 ( .B1(STATE_REG_SCAN_IN), .B2(n2843), .A(n2842), .ZN(U3323)
         );
  INV_X1 U3703 ( .A(DATAI_25_), .ZN(n2846) );
  NAND2_X1 U3704 ( .A1(n2844), .A2(STATE_REG_SCAN_IN), .ZN(n2845) );
  OAI21_X1 U3705 ( .B1(STATE_REG_SCAN_IN), .B2(n2846), .A(n2845), .ZN(U3327)
         );
  INV_X1 U3706 ( .A(DATAI_22_), .ZN(n2849) );
  NAND2_X1 U3707 ( .A1(n2847), .A2(STATE_REG_SCAN_IN), .ZN(n2848) );
  OAI21_X1 U3708 ( .B1(STATE_REG_SCAN_IN), .B2(n2849), .A(n2848), .ZN(U3330)
         );
  MUX2_X1 U3709 ( .A(n2440), .B(n3463), .S(STATE_REG_SCAN_IN), .Z(n2850) );
  INV_X1 U3710 ( .A(n2850), .ZN(U3341) );
  INV_X1 U3711 ( .A(DATAI_20_), .ZN(n2852) );
  NAND2_X1 U3712 ( .A1(n4000), .A2(STATE_REG_SCAN_IN), .ZN(n2851) );
  OAI21_X1 U3713 ( .B1(STATE_REG_SCAN_IN), .B2(n2852), .A(n2851), .ZN(U3332)
         );
  MUX2_X1 U3714 ( .A(n4075), .B(n2467), .S(U3149), .Z(n2853) );
  INV_X1 U3715 ( .A(n2853), .ZN(U3339) );
  INV_X1 U3716 ( .A(DATAI_19_), .ZN(n2854) );
  MUX2_X1 U3717 ( .A(n2854), .B(n3501), .S(STATE_REG_SCAN_IN), .Z(n2855) );
  INV_X1 U3718 ( .A(n2855), .ZN(U3333) );
  MUX2_X1 U3719 ( .A(n4100), .B(n2490), .S(U3149), .Z(n2856) );
  INV_X1 U3720 ( .A(n2856), .ZN(U3337) );
  INV_X1 U3721 ( .A(n2857), .ZN(n2858) );
  AOI22_X1 U3722 ( .A1(n4767), .A2(n2819), .B1(n2858), .B2(n4768), .ZN(U3459)
         );
  OR2_X1 U3723 ( .A1(n3122), .A2(U3149), .ZN(n4010) );
  INV_X1 U3724 ( .A(n4010), .ZN(n4005) );
  OR2_X1 U3725 ( .A1(n2982), .A2(n4005), .ZN(n2877) );
  AOI21_X1 U3726 ( .B1(n3122), .B2(n2955), .A(n2859), .ZN(n2876) );
  INV_X1 U3727 ( .A(n2876), .ZN(n2860) );
  NOR2_X1 U3728 ( .A1(n4722), .A2(U4043), .ZN(U3148) );
  INV_X1 U3729 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n4653) );
  NAND2_X1 U3730 ( .A1(U4043), .A2(n2333), .ZN(n2861) );
  OAI21_X1 U3731 ( .B1(U4043), .B2(n4653), .A(n2861), .ZN(U3551) );
  INV_X1 U3732 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n4612) );
  NAND2_X1 U3733 ( .A1(U4043), .A2(n3806), .ZN(n2862) );
  OAI21_X1 U3734 ( .B1(U4043), .B2(n4612), .A(n2862), .ZN(U3560) );
  INV_X1 U3735 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4626) );
  NAND2_X1 U3736 ( .A1(U4043), .A2(n2342), .ZN(n2863) );
  OAI21_X1 U3737 ( .B1(U4043), .B2(n4626), .A(n2863), .ZN(U3552) );
  NAND2_X1 U3738 ( .A1(n4026), .A2(n2929), .ZN(n3849) );
  AND2_X1 U3739 ( .A1(n3847), .A2(n3849), .ZN(n3946) );
  INV_X1 U3740 ( .A(n3946), .ZN(n4746) );
  NAND2_X1 U3741 ( .A1(n3220), .A2(n4475), .ZN(n2865) );
  NOR2_X1 U3742 ( .A1(n2973), .A2(n4439), .ZN(n2864) );
  AOI21_X1 U3743 ( .B1(n4746), .B2(n2865), .A(n2864), .ZN(n4748) );
  NAND2_X1 U3744 ( .A1(n2956), .A2(n2997), .ZN(n4749) );
  INV_X1 U3745 ( .A(n4749), .ZN(n2866) );
  AOI21_X1 U3746 ( .B1(n4746), .B2(n4776), .A(n2866), .ZN(n2867) );
  AND2_X1 U3747 ( .A1(n4748), .A2(n2867), .ZN(n4775) );
  NAND2_X1 U3748 ( .A1(n4784), .A2(REG1_REG_0__SCAN_IN), .ZN(n2868) );
  OAI21_X1 U3749 ( .B1(n4784), .B2(n4775), .A(n2868), .ZN(U3518) );
  MUX2_X1 U3750 ( .A(REG2_REG_2__SCAN_IN), .B(n2869), .S(n4697), .Z(n2874) );
  INV_X1 U3751 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2871) );
  AND2_X1 U3752 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2872)
         );
  NAND2_X1 U3753 ( .A1(n2870), .A2(REG2_REG_1__SCAN_IN), .ZN(n2941) );
  NAND2_X1 U3754 ( .A1(n4028), .A2(n2941), .ZN(n2873) );
  NAND2_X1 U3755 ( .A1(n2874), .A2(n2873), .ZN(n2944) );
  NAND2_X1 U3756 ( .A1(n4697), .A2(REG2_REG_2__SCAN_IN), .ZN(n2875) );
  NAND2_X1 U3757 ( .A1(n2944), .A2(n2875), .ZN(n2890) );
  XNOR2_X1 U3758 ( .A(n2889), .B(REG2_REG_3__SCAN_IN), .ZN(n2888) );
  NAND2_X1 U3759 ( .A1(n2877), .A2(n2876), .ZN(n4708) );
  NAND2_X1 U3760 ( .A1(n4705), .A2(n2989), .ZN(n4007) );
  INV_X1 U3761 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4736) );
  NOR2_X1 U3762 ( .A1(STATE_REG_SCAN_IN), .A2(n4736), .ZN(n3137) );
  NOR2_X1 U3763 ( .A1(n4735), .A2(n2884), .ZN(n2878) );
  AOI211_X1 U3764 ( .C1(n4722), .C2(ADDR_REG_3__SCAN_IN), .A(n3137), .B(n2878), 
        .ZN(n2887) );
  INV_X1 U3765 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2881) );
  XNOR2_X1 U3766 ( .A(n2870), .B(n2881), .ZN(n4032) );
  NAND2_X1 U3767 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2931) );
  INV_X1 U3768 ( .A(n2931), .ZN(n4031) );
  NAND2_X1 U3769 ( .A1(n4032), .A2(n4031), .ZN(n4030) );
  NAND2_X1 U3770 ( .A1(n2870), .A2(REG1_REG_1__SCAN_IN), .ZN(n2882) );
  NAND2_X1 U3771 ( .A1(n4697), .A2(REG1_REG_2__SCAN_IN), .ZN(n2883) );
  OAI211_X1 U3772 ( .C1(n2885), .C2(REG1_REG_3__SCAN_IN), .A(n4730), .B(n2900), 
        .ZN(n2886) );
  OAI211_X1 U3773 ( .C1(n2888), .C2(n4719), .A(n2887), .B(n2886), .ZN(U3243)
         );
  NAND2_X1 U3774 ( .A1(n2889), .A2(REG2_REG_3__SCAN_IN), .ZN(n2892) );
  NAND2_X1 U3775 ( .A1(n2890), .A2(n4696), .ZN(n2891) );
  NAND2_X1 U3776 ( .A1(n2892), .A2(n2891), .ZN(n2893) );
  XNOR2_X1 U3777 ( .A(n2893), .B(n2901), .ZN(n4037) );
  NAND2_X1 U3778 ( .A1(n2893), .A2(n4695), .ZN(n2894) );
  MUX2_X1 U3779 ( .A(n2895), .B(REG2_REG_5__SCAN_IN), .S(n4047), .Z(n4055) );
  XNOR2_X1 U3780 ( .A(n2919), .B(REG2_REG_6__SCAN_IN), .ZN(n2911) );
  INV_X1 U3781 ( .A(n4735), .ZN(n4065) );
  AND2_X1 U3782 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3179) );
  AOI21_X1 U3783 ( .B1(n4722), .B2(ADDR_REG_6__SCAN_IN), .A(n3179), .ZN(n2897)
         );
  INV_X1 U3784 ( .A(n2897), .ZN(n2909) );
  NAND2_X1 U3785 ( .A1(n2898), .A2(n4696), .ZN(n2899) );
  NAND2_X1 U3786 ( .A1(n4042), .A2(REG1_REG_4__SCAN_IN), .ZN(n4041) );
  NAND2_X1 U3787 ( .A1(n2902), .A2(n4695), .ZN(n2903) );
  NAND2_X1 U3788 ( .A1(n4041), .A2(n2903), .ZN(n4051) );
  MUX2_X1 U3789 ( .A(n2904), .B(REG1_REG_5__SCAN_IN), .S(n4047), .Z(n4052) );
  XNOR2_X1 U3790 ( .A(n2912), .B(n4694), .ZN(n2907) );
  AOI211_X1 U3791 ( .C1(n2907), .C2(n2376), .A(n4114), .B(n2906), .ZN(n2908)
         );
  AOI211_X1 U3792 ( .C1(n4065), .C2(n4694), .A(n2909), .B(n2908), .ZN(n2910)
         );
  OAI21_X1 U3793 ( .B1(n2911), .B2(n4719), .A(n2910), .ZN(U3246) );
  NAND2_X1 U3794 ( .A1(n2912), .A2(n4694), .ZN(n2913) );
  XOR2_X1 U3795 ( .A(REG1_REG_7__SCAN_IN), .B(n4693), .Z(n2915) );
  XNOR2_X1 U3796 ( .A(n2052), .B(n2915), .ZN(n2924) );
  AND2_X1 U3797 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3242) );
  AOI21_X1 U3798 ( .B1(n4722), .B2(ADDR_REG_7__SCAN_IN), .A(n3242), .ZN(n2916)
         );
  OAI21_X1 U3799 ( .B1(n4735), .B2(n2175), .A(n2916), .ZN(n2923) );
  MUX2_X1 U3800 ( .A(n2390), .B(REG2_REG_7__SCAN_IN), .S(n4693), .Z(n2920) );
  AOI211_X1 U3801 ( .C1(n2921), .C2(n2920), .A(n4719), .B(n3056), .ZN(n2922)
         );
  AOI211_X1 U3802 ( .C1(n4730), .C2(n2924), .A(n2923), .B(n2922), .ZN(n2925)
         );
  INV_X1 U3803 ( .A(n2925), .ZN(U3247) );
  NOR2_X1 U3804 ( .A1(n3552), .A2(n2929), .ZN(n2927) );
  AOI21_X1 U3805 ( .B1(n3533), .B2(n4026), .A(n2927), .ZN(n2932) );
  NOR2_X1 U3806 ( .A1(n2972), .A2(n2929), .ZN(n2930) );
  INV_X1 U3807 ( .A(n2971), .ZN(n2934) );
  NOR2_X1 U3808 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4700)
         );
  OAI211_X1 U3809 ( .C1(n4700), .C2(n3123), .A(n2932), .B(n2969), .ZN(n2933)
         );
  NAND2_X1 U3810 ( .A1(n2934), .A2(n2933), .ZN(n2995) );
  NOR2_X1 U3811 ( .A1(n4705), .A2(n4699), .ZN(n2937) );
  AOI21_X1 U3812 ( .B1(n4705), .B2(n2935), .A(n4699), .ZN(n4702) );
  NAND2_X1 U3813 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4027) );
  OAI22_X1 U3814 ( .A1(n4702), .A2(IR_REG_0__SCAN_IN), .B1(n4027), .B2(n4007), 
        .ZN(n2936) );
  AOI211_X1 U3815 ( .C1(n2995), .C2(n2937), .A(n4025), .B(n2936), .ZN(n4038)
         );
  OAI211_X1 U3816 ( .C1(n2940), .C2(n2939), .A(n4730), .B(n2938), .ZN(n2948)
         );
  MUX2_X1 U3817 ( .A(n2869), .B(REG2_REG_2__SCAN_IN), .S(n4697), .Z(n2942) );
  NAND3_X1 U3818 ( .A1(n2942), .A2(n4028), .A3(n2941), .ZN(n2943) );
  NAND3_X1 U3819 ( .A1(n4110), .A2(n2944), .A3(n2943), .ZN(n2947) );
  NAND2_X1 U3820 ( .A1(n4065), .A2(n4697), .ZN(n2946) );
  AOI22_X1 U3821 ( .A1(n4722), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n2945) );
  NAND4_X1 U3822 ( .A1(n2948), .A2(n2947), .A3(n2946), .A4(n2945), .ZN(n2949)
         );
  OR2_X1 U3823 ( .A1(n4038), .A2(n2949), .ZN(U3242) );
  INV_X1 U3824 ( .A(n2990), .ZN(n2987) );
  NOR2_X1 U3825 ( .A1(n3458), .A2(n2965), .ZN(n2954) );
  NAND2_X1 U3826 ( .A1(n2987), .A2(n4003), .ZN(n3126) );
  INV_X1 U3827 ( .A(n3126), .ZN(n2962) );
  AOI21_X1 U3828 ( .B1(n2957), .B2(n2956), .A(n2955), .ZN(n2983) );
  INV_X1 U3829 ( .A(n2983), .ZN(n2958) );
  NAND2_X1 U3830 ( .A1(n2958), .A2(n4489), .ZN(n2959) );
  NAND2_X1 U3831 ( .A1(n2987), .A2(n2959), .ZN(n2961) );
  NAND2_X1 U3832 ( .A1(n2961), .A2(n2960), .ZN(n3125) );
  NOR3_X1 U3833 ( .A1(n2962), .A2(n3125), .A3(n2986), .ZN(n3015) );
  OAI21_X1 U3834 ( .B1(n3650), .B2(n2967), .A(n2963), .ZN(n2966) );
  NAND2_X4 U3835 ( .A1(n2965), .A2(n2964), .ZN(n3658) );
  OAI22_X1 U3836 ( .A1(n3605), .A2(n3068), .B1(n3604), .B2(n2967), .ZN(n3128)
         );
  XNOR2_X1 U3837 ( .A(n3129), .B(n2968), .ZN(n2981) );
  OR2_X1 U3838 ( .A1(n3552), .A2(n2975), .ZN(n2976) );
  OAI21_X1 U3839 ( .B1(n2973), .B2(n2004), .A(n2976), .ZN(n2978) );
  OAI21_X1 U3840 ( .B1(n2981), .B2(n2980), .A(n3131), .ZN(n2985) );
  AND2_X1 U3841 ( .A1(n2983), .A2(n2982), .ZN(n2984) );
  NAND2_X1 U3842 ( .A1(n2985), .A2(n3838), .ZN(n2993) );
  NOR3_X1 U3843 ( .A1(n2987), .A2(n2986), .A3(n4489), .ZN(n2988) );
  INV_X1 U3844 ( .A(n2003), .ZN(n3737) );
  NAND3_X1 U3845 ( .A1(n2990), .A2(n4003), .A3(n4699), .ZN(n3840) );
  NAND3_X1 U3846 ( .A1(n2990), .A2(n4003), .A3(n2989), .ZN(n3783) );
  OAI22_X1 U3847 ( .A1(n3132), .A2(n3840), .B1(n3783), .B2(n2973), .ZN(n2991)
         );
  AOI21_X1 U3848 ( .B1(n3737), .B2(n3073), .A(n2991), .ZN(n2992) );
  OAI211_X1 U3849 ( .C1(n3015), .C2(n2994), .A(n2993), .B(n2992), .ZN(U3234)
         );
  OAI22_X1 U3850 ( .A1(n3831), .A2(n2995), .B1(n3840), .B2(n2973), .ZN(n2996)
         );
  AOI21_X1 U3851 ( .B1(n3737), .B2(n2997), .A(n2996), .ZN(n2998) );
  OAI21_X1 U3852 ( .B1(n3015), .B2(n2999), .A(n2998), .ZN(U3229) );
  INV_X1 U3853 ( .A(n3000), .ZN(n3004) );
  AOI22_X1 U3854 ( .A1(n4437), .A2(n3011), .B1(n4485), .B2(n4026), .ZN(n3001)
         );
  OAI21_X1 U3855 ( .B1(n3068), .B2(n4439), .A(n3001), .ZN(n3003) );
  AOI211_X1 U3856 ( .C1(n4776), .C2(n3004), .A(n3003), .B(n3002), .ZN(n3080)
         );
  MUX2_X1 U3857 ( .A(n4560), .B(n3080), .S(n4783), .Z(n3005) );
  OAI21_X1 U3858 ( .B1(n4546), .B2(n3082), .A(n3005), .ZN(U3469) );
  AOI211_X1 U3859 ( .C1(n3008), .C2(n3006), .A(n3831), .B(n3007), .ZN(n3009)
         );
  INV_X1 U3860 ( .A(n3009), .ZN(n3013) );
  OAI22_X1 U3861 ( .A1(n2928), .A2(n3783), .B1(n3840), .B2(n3068), .ZN(n3010)
         );
  AOI21_X1 U3862 ( .B1(n3737), .B2(n3011), .A(n3010), .ZN(n3012) );
  OAI211_X1 U3863 ( .C1(n3015), .C2(n3014), .A(n3013), .B(n3012), .ZN(U3219)
         );
  INV_X1 U3864 ( .A(n3016), .ZN(n3020) );
  AOI22_X1 U3865 ( .A1(n3073), .A2(n4409), .B1(n2333), .B2(n4485), .ZN(n3017)
         );
  OAI21_X1 U3866 ( .B1(n3132), .B2(n4439), .A(n3017), .ZN(n3019) );
  AOI211_X1 U3867 ( .C1(n4776), .C2(n3020), .A(n3019), .B(n3018), .ZN(n3083)
         );
  MUX2_X1 U3868 ( .A(n3021), .B(n3083), .S(n4783), .Z(n3022) );
  OAI21_X1 U3869 ( .B1(n3085), .B2(n4546), .A(n3022), .ZN(U3471) );
  NOR2_X1 U3870 ( .A1(n3049), .A2(n3246), .ZN(n3023) );
  OR2_X1 U3871 ( .A1(n3099), .A2(n3023), .ZN(n3251) );
  AND2_X1 U3872 ( .A1(n2110), .A2(n3873), .ZN(n3934) );
  INV_X1 U3873 ( .A(n3934), .ZN(n3025) );
  XNOR2_X1 U3874 ( .A(n3026), .B(n3025), .ZN(n3027) );
  NAND2_X1 U3875 ( .A1(n3027), .A2(n4338), .ZN(n3257) );
  XNOR2_X1 U3876 ( .A(n3028), .B(n3934), .ZN(n3245) );
  NAND2_X1 U3877 ( .A1(n4437), .A2(n3029), .ZN(n3031) );
  NAND2_X1 U3878 ( .A1(n4023), .A2(n4485), .ZN(n3030) );
  OAI211_X1 U3879 ( .C1(n3248), .C2(n4439), .A(n3031), .B(n3030), .ZN(n3032)
         );
  AOI21_X1 U3880 ( .B1(n3245), .B2(n4480), .A(n3032), .ZN(n3033) );
  NAND2_X1 U3881 ( .A1(n3257), .A2(n3033), .ZN(n3090) );
  NAND2_X1 U3882 ( .A1(n3090), .A2(n4783), .ZN(n3035) );
  NAND2_X1 U3883 ( .A1(n4782), .A2(REG0_REG_5__SCAN_IN), .ZN(n3034) );
  OAI211_X1 U3884 ( .C1(n3251), .C2(n4546), .A(n3035), .B(n3034), .ZN(U3477)
         );
  OAI21_X1 U3885 ( .B1(n3036), .B2(n3135), .A(n3132), .ZN(n3038) );
  NAND2_X1 U3886 ( .A1(n3036), .A2(n3135), .ZN(n3037) );
  NAND2_X1 U3887 ( .A1(n3038), .A2(n3037), .ZN(n3039) );
  XNOR2_X1 U3888 ( .A(n3040), .B(n3039), .ZN(n4777) );
  INV_X1 U3889 ( .A(n4777), .ZN(n3055) );
  INV_X1 U3890 ( .A(n3220), .ZN(n4262) );
  NAND2_X1 U3891 ( .A1(n4777), .A2(n4262), .ZN(n3048) );
  INV_X1 U3892 ( .A(n3040), .ZN(n3935) );
  XNOR2_X1 U3893 ( .A(n3041), .B(n3935), .ZN(n3046) );
  NAND2_X1 U3894 ( .A1(n4437), .A2(n3042), .ZN(n3044) );
  NAND2_X1 U3895 ( .A1(n4485), .A2(n4024), .ZN(n3043) );
  OAI211_X1 U3896 ( .C1(n3160), .C2(n4439), .A(n3044), .B(n3043), .ZN(n3045)
         );
  AOI21_X1 U3897 ( .B1(n3046), .B2(n4338), .A(n3045), .ZN(n3047) );
  NAND2_X1 U3898 ( .A1(n3048), .A2(n3047), .ZN(n4781) );
  INV_X1 U3899 ( .A(n3075), .ZN(n3051) );
  INV_X1 U3900 ( .A(n3049), .ZN(n3050) );
  OAI211_X1 U3901 ( .C1(n3051), .C2(n3150), .A(n3050), .B(n4492), .ZN(n4778)
         );
  OAI22_X1 U3902 ( .A1(n4755), .A2(n3154), .B1(n4316), .B2(n4778), .ZN(n3052)
         );
  OAI21_X1 U3903 ( .B1(n4781), .B2(n3052), .A(n4752), .ZN(n3054) );
  NAND2_X1 U3904 ( .A1(n4745), .A2(REG2_REG_4__SCAN_IN), .ZN(n3053) );
  OAI211_X1 U3905 ( .C1(n3055), .C2(n4738), .A(n3054), .B(n3053), .ZN(U3286)
         );
  XNOR2_X2 U3906 ( .A(n3111), .B(n3110), .ZN(n3112) );
  XNOR2_X1 U3907 ( .A(n3112), .B(REG1_REG_8__SCAN_IN), .ZN(n3062) );
  NAND2_X1 U3908 ( .A1(U3149), .A2(REG3_REG_8__SCAN_IN), .ZN(n3290) );
  XNOR2_X1 U3909 ( .A(n3106), .B(REG2_REG_8__SCAN_IN), .ZN(n3057) );
  NAND2_X1 U3910 ( .A1(n4110), .A2(n3057), .ZN(n3058) );
  NAND2_X1 U3911 ( .A1(n3290), .A2(n3058), .ZN(n3060) );
  NOR2_X1 U3912 ( .A1(n4735), .A2(n3110), .ZN(n3059) );
  AOI211_X1 U3913 ( .C1(n4722), .C2(ADDR_REG_8__SCAN_IN), .A(n3060), .B(n3059), 
        .ZN(n3061) );
  OAI21_X1 U3914 ( .B1(n3062), .B2(n4114), .A(n3061), .ZN(U3248) );
  XOR2_X1 U3915 ( .A(n3036), .B(n3939), .Z(n4739) );
  INV_X1 U3916 ( .A(n4739), .ZN(n3071) );
  OAI21_X1 U3917 ( .B1(n3939), .B2(n3064), .A(n3063), .ZN(n3065) );
  NAND2_X1 U3918 ( .A1(n3065), .A2(n4338), .ZN(n3067) );
  AOI22_X1 U3919 ( .A1(n4409), .A2(n3072), .B1(n4023), .B2(n4486), .ZN(n3066)
         );
  OAI211_X1 U3920 ( .C1(n3068), .C2(n4386), .A(n3067), .B(n3066), .ZN(n3069)
         );
  AOI21_X1 U3921 ( .B1(n4739), .B2(n4262), .A(n3069), .ZN(n4744) );
  OAI21_X1 U3922 ( .B1(n3071), .B2(n3070), .A(n4744), .ZN(n3086) );
  NAND2_X1 U3923 ( .A1(n3086), .A2(n4787), .ZN(n3078) );
  OAI21_X1 U3924 ( .B1(n3074), .B2(n3073), .A(n3072), .ZN(n3076) );
  AND2_X1 U3925 ( .A1(n3076), .A2(n3075), .ZN(n4740) );
  NAND2_X1 U3926 ( .A1(n2782), .A2(n4740), .ZN(n3077) );
  OAI211_X1 U3927 ( .C1(n4787), .C2(n3079), .A(n3078), .B(n3077), .ZN(U3521)
         );
  MUX2_X1 U3928 ( .A(n2881), .B(n3080), .S(n4787), .Z(n3081) );
  OAI21_X1 U3929 ( .B1(n4483), .B2(n3082), .A(n3081), .ZN(U3519) );
  MUX2_X1 U3930 ( .A(n2880), .B(n3083), .S(n4787), .Z(n3084) );
  OAI21_X1 U3931 ( .B1(n3085), .B2(n4483), .A(n3084), .ZN(U3520) );
  NAND2_X1 U3932 ( .A1(n3086), .A2(n4783), .ZN(n3088) );
  NAND2_X1 U3933 ( .A1(n2788), .A2(n4740), .ZN(n3087) );
  OAI211_X1 U3934 ( .C1(n4783), .C2(n3089), .A(n3088), .B(n3087), .ZN(U3473)
         );
  MUX2_X1 U3935 ( .A(n3090), .B(REG1_REG_5__SCAN_IN), .S(n4784), .Z(n3091) );
  INV_X1 U3936 ( .A(n3091), .ZN(n3092) );
  OAI21_X1 U3937 ( .B1(n4483), .B2(n3251), .A(n3092), .ZN(U3523) );
  INV_X1 U3938 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n4611) );
  NAND2_X1 U3939 ( .A1(n4393), .A2(U4043), .ZN(n3093) );
  OAI21_X1 U3940 ( .B1(n4611), .B2(U4043), .A(n3093), .ZN(U3573) );
  AND2_X1 U3941 ( .A1(n3861), .A2(n3875), .ZN(n3938) );
  XOR2_X1 U3942 ( .A(n3938), .B(n3094), .Z(n3308) );
  XOR2_X1 U3943 ( .A(n3095), .B(n3938), .Z(n3306) );
  AOI22_X1 U3944 ( .A1(n3301), .A2(n4409), .B1(n4020), .B2(n4486), .ZN(n3096)
         );
  OAI21_X1 U3945 ( .B1(n3160), .B2(n4386), .A(n3096), .ZN(n3097) );
  AOI21_X1 U3946 ( .B1(n3306), .B2(n4480), .A(n3097), .ZN(n3098) );
  OAI21_X1 U3947 ( .B1(n3308), .B2(n4475), .A(n3098), .ZN(n3120) );
  OR2_X1 U3948 ( .A1(n3099), .A2(n3177), .ZN(n3100) );
  NAND2_X1 U3949 ( .A1(n3201), .A2(n3100), .ZN(n3296) );
  INV_X1 U3950 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3101) );
  OAI22_X1 U3951 ( .A1(n4546), .A2(n3296), .B1(n4783), .B2(n3101), .ZN(n3102)
         );
  AOI21_X1 U3952 ( .B1(n3120), .B2(n4783), .A(n3102), .ZN(n3103) );
  INV_X1 U3953 ( .A(n3103), .ZN(U3479) );
  XNOR2_X1 U3954 ( .A(n4692), .B(n3325), .ZN(n3211) );
  XOR2_X1 U3955 ( .A(n2053), .B(n3211), .Z(n3117) );
  INV_X1 U3956 ( .A(n4692), .ZN(n3109) );
  NOR2_X1 U3957 ( .A1(n3107), .A2(STATE_REG_SCAN_IN), .ZN(n3344) );
  AOI21_X1 U3958 ( .B1(n4722), .B2(ADDR_REG_9__SCAN_IN), .A(n3344), .ZN(n3108)
         );
  OAI21_X1 U3959 ( .B1(n4735), .B2(n3109), .A(n3108), .ZN(n3116) );
  MUX2_X1 U3960 ( .A(n3321), .B(REG1_REG_9__SCAN_IN), .S(n4692), .Z(n3113) );
  AOI211_X1 U3961 ( .C1(n4110), .C2(n3117), .A(n3116), .B(n3115), .ZN(n3118)
         );
  INV_X1 U3962 ( .A(n3118), .ZN(U3249) );
  OAI22_X1 U3963 ( .A1(n4483), .A2(n3296), .B1(n4787), .B2(n2376), .ZN(n3119)
         );
  AOI21_X1 U3964 ( .B1(n3120), .B2(n4787), .A(n3119), .ZN(n3121) );
  INV_X1 U3965 ( .A(n3121), .ZN(U3524) );
  NAND2_X1 U3966 ( .A1(n3123), .A2(n3122), .ZN(n3124) );
  OAI21_X1 U3967 ( .B1(n3125), .B2(n3124), .A(STATE_REG_SCAN_IN), .ZN(n3127)
         );
  OAI22_X1 U3968 ( .A1(n3605), .A2(n3132), .B1(n3655), .B2(n3135), .ZN(n3142)
         );
  OAI22_X1 U3969 ( .A1(n3132), .A2(n3552), .B1(n3650), .B2(n3135), .ZN(n3133)
         );
  XNOR2_X1 U3970 ( .A(n3133), .B(n3658), .ZN(n3141) );
  XOR2_X1 U3971 ( .A(n3142), .B(n3141), .Z(n3145) );
  XNOR2_X1 U3972 ( .A(n3146), .B(n3145), .ZN(n3134) );
  NAND2_X1 U3973 ( .A1(n3134), .A2(n3838), .ZN(n3139) );
  OAI22_X1 U3974 ( .A1(n2003), .A2(n3135), .B1(n3249), .B2(n3840), .ZN(n3136)
         );
  AOI211_X1 U3975 ( .C1(n3843), .C2(n2342), .A(n3137), .B(n3136), .ZN(n3138)
         );
  OAI211_X1 U3976 ( .C1(REG3_REG_3__SCAN_IN), .C2(n3846), .A(n3139), .B(n3138), 
        .ZN(U3215) );
  INV_X1 U3977 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4671) );
  NAND2_X1 U3978 ( .A1(n3824), .A2(U4043), .ZN(n3140) );
  OAI21_X1 U3979 ( .B1(U4043), .B2(n4671), .A(n3140), .ZN(U3575) );
  INV_X1 U3980 ( .A(n3141), .ZN(n3144) );
  INV_X1 U3981 ( .A(n3142), .ZN(n3143) );
  OAI22_X1 U3982 ( .A1(n3605), .A2(n3249), .B1(n3655), .B2(n3150), .ZN(n3155)
         );
  OAI22_X1 U3983 ( .A1(n3249), .A2(n3655), .B1(n3650), .B2(n3150), .ZN(n3147)
         );
  XNOR2_X1 U3984 ( .A(n3147), .B(n3658), .ZN(n3156) );
  XOR2_X1 U3985 ( .A(n3155), .B(n3156), .Z(n3148) );
  OAI211_X1 U3986 ( .C1(n3149), .C2(n3148), .A(n3157), .B(n3838), .ZN(n3153)
         );
  AND2_X1 U3987 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n4040) );
  OAI22_X1 U3988 ( .A1(n2003), .A2(n3150), .B1(n3160), .B2(n3840), .ZN(n3151)
         );
  AOI211_X1 U3989 ( .C1(n3843), .C2(n4024), .A(n4040), .B(n3151), .ZN(n3152)
         );
  OAI211_X1 U3990 ( .C1(n3846), .C2(n3154), .A(n3153), .B(n3152), .ZN(U3227)
         );
  INV_X1 U3991 ( .A(n3155), .ZN(n3159) );
  INV_X1 U3992 ( .A(n3156), .ZN(n3158) );
  OAI22_X1 U3993 ( .A1(n3605), .A2(n3160), .B1(n3655), .B2(n3246), .ZN(n3169)
         );
  OR2_X1 U3994 ( .A1(n3655), .A2(n3160), .ZN(n3161) );
  OAI21_X1 U3995 ( .B1(n3650), .B2(n3246), .A(n3161), .ZN(n3162) );
  XNOR2_X1 U3996 ( .A(n3162), .B(n3658), .ZN(n3168) );
  XOR2_X1 U3997 ( .A(n3169), .B(n3168), .Z(n3163) );
  OAI211_X1 U3998 ( .C1(n3164), .C2(n3163), .A(n3172), .B(n3838), .ZN(n3167)
         );
  NOR2_X1 U3999 ( .A1(STATE_REG_SCAN_IN), .A2(n2365), .ZN(n4049) );
  OAI22_X1 U4000 ( .A1(n2003), .A2(n3246), .B1(n3248), .B2(n3840), .ZN(n3165)
         );
  AOI211_X1 U4001 ( .C1(n3843), .C2(n4023), .A(n4049), .B(n3165), .ZN(n3166)
         );
  OAI211_X1 U4002 ( .C1(n3846), .C2(n3250), .A(n3167), .B(n3166), .ZN(U3224)
         );
  INV_X1 U4003 ( .A(n3168), .ZN(n3171) );
  INV_X1 U4004 ( .A(n3169), .ZN(n3170) );
  OAI22_X1 U4005 ( .A1(n3248), .A2(n3655), .B1(n3650), .B2(n3177), .ZN(n3173)
         );
  XNOR2_X1 U4006 ( .A(n3173), .B(n3658), .ZN(n3233) );
  OAI22_X1 U4007 ( .A1(n3605), .A2(n3248), .B1(n3655), .B2(n3177), .ZN(n3234)
         );
  XNOR2_X1 U4008 ( .A(n3233), .B(n3234), .ZN(n3175) );
  XNOR2_X1 U4009 ( .A(n3235), .B(n3175), .ZN(n3176) );
  NAND2_X1 U4010 ( .A1(n3176), .A2(n3838), .ZN(n3181) );
  OAI22_X1 U4011 ( .A1(n2003), .A2(n3177), .B1(n3304), .B2(n3840), .ZN(n3178)
         );
  AOI211_X1 U4012 ( .C1(n3843), .C2(n4022), .A(n3179), .B(n3178), .ZN(n3180)
         );
  OAI211_X1 U4013 ( .C1(n3846), .C2(n3297), .A(n3181), .B(n3180), .ZN(U3236)
         );
  AND2_X1 U4014 ( .A1(n3864), .A2(n3876), .ZN(n3937) );
  XOR2_X1 U4015 ( .A(n3182), .B(n3937), .Z(n3223) );
  NAND2_X1 U4016 ( .A1(n3184), .A2(n3183), .ZN(n3197) );
  INV_X1 U4017 ( .A(n3185), .ZN(n3947) );
  NOR2_X1 U4018 ( .A1(n3197), .A2(n3947), .ZN(n3196) );
  NOR2_X1 U4019 ( .A1(n3196), .A2(n3186), .ZN(n3187) );
  XNOR2_X1 U4020 ( .A(n3187), .B(n3937), .ZN(n3232) );
  OAI22_X1 U4021 ( .A1(n4386), .A2(n3304), .B1(n3338), .B2(n4439), .ZN(n3188)
         );
  AOI21_X1 U4022 ( .B1(n3289), .B2(n4437), .A(n3188), .ZN(n3189) );
  OAI21_X1 U4023 ( .B1(n3232), .B2(n4497), .A(n3189), .ZN(n3190) );
  AOI21_X1 U4024 ( .B1(n4338), .B2(n3223), .A(n3190), .ZN(n3195) );
  AND2_X1 U4025 ( .A1(n3198), .A2(n3289), .ZN(n3191) );
  NOR2_X1 U4026 ( .A1(n3271), .A2(n3191), .ZN(n3224) );
  AOI22_X1 U4027 ( .A1(n2788), .A2(n3224), .B1(REG0_REG_8__SCAN_IN), .B2(n4782), .ZN(n3192) );
  OAI21_X1 U4028 ( .B1(n3195), .B2(n4782), .A(n3192), .ZN(U3483) );
  NAND2_X1 U4029 ( .A1(n4784), .A2(REG1_REG_8__SCAN_IN), .ZN(n3194) );
  NAND2_X1 U4030 ( .A1(n2782), .A2(n3224), .ZN(n3193) );
  OAI211_X1 U4031 ( .C1(n3195), .C2(n4784), .A(n3194), .B(n3193), .ZN(U3526)
         );
  AOI21_X1 U4032 ( .B1(n3947), .B2(n3197), .A(n3196), .ZN(n3262) );
  INV_X1 U4033 ( .A(n3198), .ZN(n3199) );
  AOI211_X1 U4034 ( .C1(n3204), .C2(n3201), .A(n3200), .B(n3199), .ZN(n3259)
         );
  XNOR2_X1 U4035 ( .A(n3202), .B(n3947), .ZN(n3203) );
  NAND2_X1 U4036 ( .A1(n3203), .A2(n4338), .ZN(n3206) );
  AOI22_X1 U4037 ( .A1(n4437), .A2(n3204), .B1(n4485), .B2(n4021), .ZN(n3205)
         );
  OAI211_X1 U4038 ( .C1(n3341), .C2(n4439), .A(n3206), .B(n3205), .ZN(n3258)
         );
  AOI211_X1 U4039 ( .C1(n3262), .C2(n4480), .A(n3259), .B(n3258), .ZN(n3209)
         );
  NAND2_X1 U4040 ( .A1(n4784), .A2(REG1_REG_7__SCAN_IN), .ZN(n3207) );
  OAI21_X1 U4041 ( .B1(n3209), .B2(n4784), .A(n3207), .ZN(U3525) );
  NAND2_X1 U4042 ( .A1(n4782), .A2(REG0_REG_7__SCAN_IN), .ZN(n3208) );
  OAI21_X1 U40430 ( .B1(n3209), .B2(n4782), .A(n3208), .ZN(U3481) );
  XNOR2_X1 U4044 ( .A(n3376), .B(REG1_REG_10__SCAN_IN), .ZN(n3217) );
  XOR2_X1 U4045 ( .A(n3380), .B(REG2_REG_10__SCAN_IN), .Z(n3212) );
  NAND2_X1 U4046 ( .A1(n4110), .A2(n3212), .ZN(n3213) );
  NAND2_X1 U4047 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n3396) );
  NAND2_X1 U4048 ( .A1(n3213), .A2(n3396), .ZN(n3214) );
  AOI21_X1 U4049 ( .B1(n4722), .B2(ADDR_REG_10__SCAN_IN), .A(n3214), .ZN(n3216) );
  NAND2_X1 U4050 ( .A1(n4065), .A2(n4691), .ZN(n3215) );
  OAI211_X1 U4051 ( .C1(n3217), .C2(n4114), .A(n3216), .B(n3215), .ZN(U3250)
         );
  INV_X1 U4052 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n4577) );
  NAND2_X1 U4053 ( .A1(n4143), .A2(U4043), .ZN(n3218) );
  OAI21_X1 U4054 ( .B1(U4043), .B2(n4577), .A(n3218), .ZN(U3579) );
  AND2_X1 U4055 ( .A1(n3220), .A2(n3219), .ZN(n3221) );
  OR2_X1 U4056 ( .A1(n4745), .A2(n4475), .ZN(n3413) );
  INV_X1 U4057 ( .A(n3413), .ZN(n3222) );
  NAND2_X1 U4058 ( .A1(n3223), .A2(n3222), .ZN(n3231) );
  INV_X1 U4059 ( .A(n4371), .ZN(n4343) );
  INV_X1 U4060 ( .A(n3224), .ZN(n3227) );
  INV_X1 U4061 ( .A(n3225), .ZN(n3293) );
  AOI22_X1 U4062 ( .A1(n4745), .A2(REG2_REG_8__SCAN_IN), .B1(n3293), .B2(n4737), .ZN(n3226) );
  OAI21_X1 U4063 ( .B1(n4364), .B2(n3227), .A(n3226), .ZN(n3229) );
  OAI22_X1 U4064 ( .A1(n3304), .A2(n4369), .B1(n4370), .B2(n3284), .ZN(n3228)
         );
  AOI211_X1 U4065 ( .C1(n4343), .C2(n4018), .A(n3229), .B(n3228), .ZN(n3230)
         );
  OAI211_X1 U4066 ( .C1(n4378), .C2(n3232), .A(n3231), .B(n3230), .ZN(U3282)
         );
  INV_X1 U4067 ( .A(n3234), .ZN(n3236) );
  OR2_X1 U4068 ( .A1(n3655), .A2(n3304), .ZN(n3237) );
  OAI21_X1 U4069 ( .B1(n3650), .B2(n3240), .A(n3237), .ZN(n3238) );
  XNOR2_X1 U4070 ( .A(n3238), .B(n3645), .ZN(n3279) );
  OAI22_X1 U4071 ( .A1(n3605), .A2(n3304), .B1(n3655), .B2(n3240), .ZN(n3277)
         );
  XNOR2_X1 U4072 ( .A(n3279), .B(n3277), .ZN(n3275) );
  XOR2_X1 U4073 ( .A(n3276), .B(n3275), .Z(n3239) );
  NAND2_X1 U4074 ( .A1(n3239), .A2(n3838), .ZN(n3244) );
  INV_X1 U4075 ( .A(n3840), .ZN(n3823) );
  OAI22_X1 U4076 ( .A1(n2003), .A2(n3240), .B1(n3248), .B2(n3783), .ZN(n3241)
         );
  AOI211_X1 U4077 ( .C1(n3823), .C2(n4019), .A(n3242), .B(n3241), .ZN(n3243)
         );
  OAI211_X1 U4078 ( .C1(n3846), .C2(n3260), .A(n3244), .B(n3243), .ZN(U3210)
         );
  INV_X1 U4079 ( .A(n3245), .ZN(n3247) );
  OAI22_X1 U4080 ( .A1(n4378), .A2(n3247), .B1(n4370), .B2(n3246), .ZN(n3255)
         );
  OAI22_X1 U4081 ( .A1(n3249), .A2(n4369), .B1(n4371), .B2(n3248), .ZN(n3254)
         );
  OAI22_X1 U4082 ( .A1(n4752), .A2(n2895), .B1(n3250), .B2(n4755), .ZN(n3253)
         );
  NOR2_X1 U4083 ( .A1(n4364), .A2(n3251), .ZN(n3252) );
  NOR4_X1 U4084 ( .A1(n3255), .A2(n3254), .A3(n3253), .A4(n3252), .ZN(n3256)
         );
  OAI21_X1 U4085 ( .B1(n4745), .B2(n3257), .A(n3256), .ZN(U3285) );
  AOI21_X1 U4086 ( .B1(n3259), .B2(n3501), .A(n3258), .ZN(n3264) );
  OAI22_X1 U4087 ( .A1(n4752), .A2(n2390), .B1(n3260), .B2(n4755), .ZN(n3261)
         );
  AOI21_X1 U4088 ( .B1(n3262), .B2(n4336), .A(n3261), .ZN(n3263) );
  OAI21_X1 U4089 ( .B1(n3264), .B2(n4745), .A(n3263), .ZN(U3283) );
  AND2_X1 U4090 ( .A1(n2042), .A2(n3865), .ZN(n3940) );
  XNOR2_X1 U4091 ( .A(n3265), .B(n3940), .ZN(n3332) );
  AOI22_X1 U4092 ( .A1(n4437), .A2(n3266), .B1(n4019), .B2(n4485), .ZN(n3267)
         );
  OAI21_X1 U4093 ( .B1(n3427), .B2(n4439), .A(n3267), .ZN(n3270) );
  XNOR2_X1 U4094 ( .A(n3268), .B(n3940), .ZN(n3269) );
  NOR2_X1 U4095 ( .A1(n3269), .A2(n4475), .ZN(n3324) );
  AOI211_X1 U4096 ( .C1(n3332), .C2(n4480), .A(n3270), .B(n3324), .ZN(n3320)
         );
  NAND2_X1 U4097 ( .A1(n4782), .A2(REG0_REG_9__SCAN_IN), .ZN(n3274) );
  NOR2_X1 U4098 ( .A1(n3271), .A2(n3342), .ZN(n3272) );
  OR2_X1 U4099 ( .A1(n3311), .A2(n3272), .ZN(n3323) );
  INV_X1 U4100 ( .A(n3323), .ZN(n3328) );
  NAND2_X1 U4101 ( .A1(n2788), .A2(n3328), .ZN(n3273) );
  OAI211_X1 U4102 ( .C1(n3320), .C2(n4782), .A(n3274), .B(n3273), .ZN(U3485)
         );
  NAND2_X1 U4103 ( .A1(n3276), .A2(n3275), .ZN(n3281) );
  INV_X1 U4104 ( .A(n3277), .ZN(n3278) );
  NAND2_X1 U4105 ( .A1(n3281), .A2(n3280), .ZN(n3337) );
  OR2_X1 U4106 ( .A1(n3655), .A2(n3341), .ZN(n3282) );
  OAI21_X1 U4107 ( .B1(n3650), .B2(n3284), .A(n3282), .ZN(n3283) );
  XNOR2_X1 U4108 ( .A(n3283), .B(n3658), .ZN(n3286) );
  OAI22_X1 U4109 ( .A1(n3605), .A2(n3341), .B1(n3655), .B2(n3284), .ZN(n3285)
         );
  OR2_X1 U4110 ( .A1(n3286), .A2(n3285), .ZN(n3335) );
  INV_X1 U4111 ( .A(n3335), .ZN(n3287) );
  AND2_X1 U4112 ( .A1(n3286), .A2(n3285), .ZN(n3336) );
  NOR2_X1 U4113 ( .A1(n3287), .A2(n3336), .ZN(n3288) );
  XNOR2_X1 U4114 ( .A(n3337), .B(n3288), .ZN(n3295) );
  AOI22_X1 U4115 ( .A1(n3737), .A2(n3289), .B1(n3823), .B2(n4018), .ZN(n3291)
         );
  OAI211_X1 U4116 ( .C1(n3304), .C2(n3783), .A(n3291), .B(n3290), .ZN(n3292)
         );
  AOI21_X1 U4117 ( .B1(n3293), .B2(n3829), .A(n3292), .ZN(n3294) );
  OAI21_X1 U4118 ( .B1(n3295), .B2(n3831), .A(n3294), .ZN(U3218) );
  INV_X1 U4119 ( .A(n3296), .ZN(n3300) );
  OAI22_X1 U4120 ( .A1(n4752), .A2(n3298), .B1(n3297), .B2(n4755), .ZN(n3299)
         );
  AOI21_X1 U4121 ( .B1(n4741), .B2(n3300), .A(n3299), .ZN(n3303) );
  INV_X1 U4122 ( .A(n4370), .ZN(n4344) );
  INV_X1 U4123 ( .A(n4369), .ZN(n3327) );
  AOI22_X1 U4124 ( .A1(n3301), .A2(n4344), .B1(n3327), .B2(n4022), .ZN(n3302)
         );
  OAI211_X1 U4125 ( .C1(n3304), .C2(n4371), .A(n3303), .B(n3302), .ZN(n3305)
         );
  AOI21_X1 U4126 ( .B1(n3306), .B2(n4336), .A(n3305), .ZN(n3307) );
  OAI21_X1 U4127 ( .B1(n3413), .B2(n3308), .A(n3307), .ZN(U3284) );
  AND2_X1 U4128 ( .A1(n3883), .A2(n3886), .ZN(n3945) );
  XOR2_X1 U4129 ( .A(n3309), .B(n3945), .Z(n3367) );
  XOR2_X1 U4130 ( .A(n3310), .B(n3945), .Z(n3365) );
  OAI22_X1 U4131 ( .A1(n3338), .A2(n4369), .B1(n4370), .B2(n3397), .ZN(n3318)
         );
  OR2_X1 U4132 ( .A1(n3311), .A2(n3397), .ZN(n3312) );
  NAND2_X1 U4133 ( .A1(n3424), .A2(n3312), .ZN(n3373) );
  INV_X1 U4134 ( .A(n3373), .ZN(n3315) );
  OAI22_X1 U4135 ( .A1(n4752), .A2(n3313), .B1(n3402), .B2(n4755), .ZN(n3314)
         );
  AOI21_X1 U4136 ( .B1(n4741), .B2(n3315), .A(n3314), .ZN(n3316) );
  OAI21_X1 U4137 ( .B1(n3739), .B2(n4371), .A(n3316), .ZN(n3317) );
  AOI211_X1 U4138 ( .C1(n3365), .C2(n4336), .A(n3318), .B(n3317), .ZN(n3319)
         );
  OAI21_X1 U4139 ( .B1(n3367), .B2(n3413), .A(n3319), .ZN(U3280) );
  MUX2_X1 U4140 ( .A(n3321), .B(n3320), .S(n4787), .Z(n3322) );
  OAI21_X1 U4141 ( .B1(n4483), .B2(n3323), .A(n3322), .ZN(U3527) );
  INV_X1 U4142 ( .A(n3324), .ZN(n3334) );
  OAI22_X1 U4143 ( .A1(n4752), .A2(n3325), .B1(n3347), .B2(n4755), .ZN(n3326)
         );
  AOI21_X1 U4144 ( .B1(n3327), .B2(n4019), .A(n3326), .ZN(n3330) );
  AOI22_X1 U4145 ( .A1(n3328), .A2(n4741), .B1(n4343), .B2(n3806), .ZN(n3329)
         );
  OAI211_X1 U4146 ( .C1(n3342), .C2(n4370), .A(n3330), .B(n3329), .ZN(n3331)
         );
  AOI21_X1 U4147 ( .B1(n4336), .B2(n3332), .A(n3331), .ZN(n3333) );
  OAI21_X1 U4148 ( .B1(n3334), .B2(n4745), .A(n3333), .ZN(U3281) );
  OAI21_X2 U4149 ( .B1(n3337), .B2(n3336), .A(n3335), .ZN(n3392) );
  OAI22_X1 U4150 ( .A1(n3605), .A2(n3338), .B1(n3655), .B2(n3342), .ZN(n3388)
         );
  OAI22_X1 U4151 ( .A1(n3338), .A2(n3655), .B1(n3650), .B2(n3342), .ZN(n3339)
         );
  XNOR2_X1 U4152 ( .A(n3339), .B(n3658), .ZN(n3389) );
  XOR2_X1 U4153 ( .A(n3388), .B(n3389), .Z(n3391) );
  XNOR2_X1 U4154 ( .A(n3392), .B(n3391), .ZN(n3340) );
  NAND2_X1 U4155 ( .A1(n3340), .A2(n3838), .ZN(n3346) );
  OAI22_X1 U4156 ( .A1(n2003), .A2(n3342), .B1(n3341), .B2(n3783), .ZN(n3343)
         );
  AOI211_X1 U4157 ( .C1(n3823), .C2(n3806), .A(n3344), .B(n3343), .ZN(n3345)
         );
  OAI211_X1 U4158 ( .C1(n3846), .C2(n3347), .A(n3346), .B(n3345), .ZN(U3228)
         );
  INV_X1 U4159 ( .A(n3349), .ZN(n3350) );
  AOI21_X1 U4160 ( .B1(n3348), .B2(n3351), .A(n3350), .ZN(n3444) );
  NAND2_X1 U4161 ( .A1(n3441), .A2(n3443), .ZN(n3354) );
  XNOR2_X1 U4162 ( .A(n3444), .B(n3354), .ZN(n3352) );
  NAND2_X1 U4163 ( .A1(n3352), .A2(n4338), .ZN(n4495) );
  INV_X1 U4164 ( .A(n3354), .ZN(n3951) );
  XNOR2_X1 U4165 ( .A(n3353), .B(n3951), .ZN(n4496) );
  INV_X1 U4166 ( .A(n4496), .ZN(n3361) );
  OAI22_X1 U4167 ( .A1(n3702), .A2(n4371), .B1(n4369), .B2(n3739), .ZN(n3360)
         );
  INV_X1 U4168 ( .A(n3355), .ZN(n3452) );
  AOI21_X1 U4169 ( .B1(n3736), .B2(n3425), .A(n3452), .ZN(n4493) );
  NAND2_X1 U4170 ( .A1(n4493), .A2(n4741), .ZN(n3358) );
  INV_X1 U4171 ( .A(n3356), .ZN(n3741) );
  AOI22_X1 U4172 ( .A1(n4745), .A2(REG2_REG_12__SCAN_IN), .B1(n3741), .B2(
        n4737), .ZN(n3357) );
  OAI211_X1 U4173 ( .C1(n4370), .C2(n4490), .A(n3358), .B(n3357), .ZN(n3359)
         );
  AOI211_X1 U4174 ( .C1(n3361), .C2(n4336), .A(n3360), .B(n3359), .ZN(n3362)
         );
  OAI21_X1 U4175 ( .B1(n4495), .B2(n4745), .A(n3362), .ZN(U3278) );
  AOI22_X1 U4176 ( .A1(n4486), .A2(n4484), .B1(n4485), .B2(n4018), .ZN(n3363)
         );
  OAI21_X1 U4177 ( .B1(n4489), .B2(n3397), .A(n3363), .ZN(n3364) );
  AOI21_X1 U4178 ( .B1(n3365), .B2(n4480), .A(n3364), .ZN(n3366) );
  OAI21_X1 U4179 ( .B1(n3367), .B2(n4475), .A(n3366), .ZN(n3370) );
  NAND2_X1 U4180 ( .A1(n3370), .A2(n4787), .ZN(n3369) );
  NAND2_X1 U4181 ( .A1(n4784), .A2(REG1_REG_10__SCAN_IN), .ZN(n3368) );
  OAI211_X1 U4182 ( .C1(n4483), .C2(n3373), .A(n3369), .B(n3368), .ZN(U3528)
         );
  NAND2_X1 U4183 ( .A1(n3370), .A2(n4783), .ZN(n3372) );
  NAND2_X1 U4184 ( .A1(n4782), .A2(REG0_REG_10__SCAN_IN), .ZN(n3371) );
  OAI211_X1 U4185 ( .C1(n3373), .C2(n4546), .A(n3372), .B(n3371), .ZN(U3487)
         );
  INV_X1 U4186 ( .A(n3374), .ZN(n3375) );
  MUX2_X1 U4187 ( .A(REG1_REG_11__SCAN_IN), .B(n3464), .S(n3463), .Z(n3377) );
  AOI211_X1 U4188 ( .C1(n3378), .C2(n3377), .A(n4114), .B(n3465), .ZN(n3387)
         );
  MUX2_X1 U4189 ( .A(REG2_REG_11__SCAN_IN), .B(n3423), .S(n3463), .Z(n3381) );
  AOI211_X1 U4190 ( .C1(n3382), .C2(n3381), .A(n4719), .B(n3481), .ZN(n3386)
         );
  NOR2_X1 U4191 ( .A1(n3383), .A2(STATE_REG_SCAN_IN), .ZN(n3805) );
  AOI21_X1 U4192 ( .B1(n4722), .B2(ADDR_REG_11__SCAN_IN), .A(n3805), .ZN(n3384) );
  OAI21_X1 U4193 ( .B1(n4735), .B2(n3463), .A(n3384), .ZN(n3385) );
  OR3_X1 U4194 ( .A1(n3387), .A2(n3386), .A3(n3385), .ZN(U3251) );
  NOR2_X1 U4195 ( .A1(n3389), .A2(n3388), .ZN(n3390) );
  AOI21_X1 U4196 ( .B1(n3392), .B2(n3391), .A(n3390), .ZN(n3395) );
  OAI22_X1 U4197 ( .A1(n3605), .A2(n3427), .B1(n3604), .B2(n3397), .ZN(n3522)
         );
  OAI22_X1 U4198 ( .A1(n3427), .A2(n3655), .B1(n3650), .B2(n3397), .ZN(n3393)
         );
  XNOR2_X1 U4199 ( .A(n3393), .B(n3658), .ZN(n3523) );
  XOR2_X1 U4200 ( .A(n3522), .B(n3523), .Z(n3394) );
  NAND2_X1 U4201 ( .A1(n3395), .A2(n3394), .ZN(n3525) );
  OAI211_X1 U4202 ( .C1(n3395), .C2(n3394), .A(n3525), .B(n3838), .ZN(n3401)
         );
  INV_X1 U4203 ( .A(n3396), .ZN(n3399) );
  OAI22_X1 U4204 ( .A1(n2003), .A2(n3397), .B1(n3739), .B2(n3840), .ZN(n3398)
         );
  AOI211_X1 U4205 ( .C1(n3843), .C2(n4018), .A(n3399), .B(n3398), .ZN(n3400)
         );
  OAI211_X1 U4206 ( .C1(n3846), .C2(n3402), .A(n3401), .B(n3400), .ZN(U3214)
         );
  XNOR2_X1 U4207 ( .A(n3403), .B(n3405), .ZN(n4474) );
  OAI21_X1 U4208 ( .B1(n2049), .B2(n3405), .A(n3404), .ZN(n4466) );
  OAI22_X1 U4209 ( .A1(n4350), .A2(n4371), .B1(n4369), .B2(n3702), .ZN(n3411)
         );
  OR2_X1 U4210 ( .A1(n3450), .A2(n4470), .ZN(n3407) );
  NAND2_X1 U4211 ( .A1(n3406), .A2(n3407), .ZN(n4543) );
  AOI22_X1 U4212 ( .A1(n4745), .A2(REG2_REG_14__SCAN_IN), .B1(n3704), .B2(
        n4737), .ZN(n3409) );
  NAND2_X1 U4213 ( .A1(n4344), .A2(n3700), .ZN(n3408) );
  OAI211_X1 U4214 ( .C1(n4543), .C2(n4364), .A(n3409), .B(n3408), .ZN(n3410)
         );
  AOI211_X1 U4215 ( .C1(n4466), .C2(n4336), .A(n3411), .B(n3410), .ZN(n3412)
         );
  OAI21_X1 U4216 ( .B1(n4474), .B2(n3413), .A(n3412), .ZN(U3276) );
  NAND2_X1 U4217 ( .A1(n3414), .A2(n3417), .ZN(n3415) );
  NAND2_X1 U4218 ( .A1(n3416), .A2(n3415), .ZN(n3433) );
  INV_X1 U4219 ( .A(n3433), .ZN(n3432) );
  XNOR2_X1 U4220 ( .A(n3348), .B(n3417), .ZN(n3422) );
  NAND2_X1 U4221 ( .A1(n3433), .A2(n4262), .ZN(n3420) );
  AOI22_X1 U4222 ( .A1(n4437), .A2(n3418), .B1(n4486), .B2(n4017), .ZN(n3419)
         );
  NAND2_X1 U4223 ( .A1(n3420), .A2(n3419), .ZN(n3421) );
  AOI21_X1 U4224 ( .B1(n3422), .B2(n4338), .A(n3421), .ZN(n3435) );
  MUX2_X1 U4225 ( .A(n3423), .B(n3435), .S(n4752), .Z(n3431) );
  INV_X1 U4226 ( .A(n3424), .ZN(n3426) );
  OAI21_X1 U4227 ( .B1(n3426), .B2(n3803), .A(n3425), .ZN(n3440) );
  INV_X1 U4228 ( .A(n3440), .ZN(n3429) );
  OAI22_X1 U4229 ( .A1(n4369), .A2(n3427), .B1(n3809), .B2(n4755), .ZN(n3428)
         );
  AOI21_X1 U4230 ( .B1(n3429), .B2(n4741), .A(n3428), .ZN(n3430) );
  OAI211_X1 U4231 ( .C1(n3432), .C2(n4738), .A(n3431), .B(n3430), .ZN(U3279)
         );
  AOI22_X1 U4232 ( .A1(n3433), .A2(n4776), .B1(n4485), .B2(n3806), .ZN(n3434)
         );
  AND2_X1 U4233 ( .A1(n3435), .A2(n3434), .ZN(n3437) );
  MUX2_X1 U4234 ( .A(n3464), .B(n3437), .S(n4787), .Z(n3436) );
  OAI21_X1 U4235 ( .B1(n4483), .B2(n3440), .A(n3436), .ZN(U3529) );
  MUX2_X1 U4236 ( .A(n3438), .B(n3437), .S(n4783), .Z(n3439) );
  OAI21_X1 U4237 ( .B1(n3440), .B2(n4546), .A(n3439), .ZN(U3489) );
  XNOR2_X1 U4238 ( .A(n3792), .B(n3702), .ZN(n3928) );
  INV_X1 U4239 ( .A(n3441), .ZN(n3442) );
  AOI21_X1 U4240 ( .B1(n3444), .B2(n3443), .A(n3442), .ZN(n3445) );
  XOR2_X1 U4241 ( .A(n3928), .B(n3445), .Z(n3448) );
  OAI22_X1 U4242 ( .A1(n4368), .A2(n4439), .B1(n3802), .B2(n4386), .ZN(n3446)
         );
  AOI21_X1 U4243 ( .B1(n3534), .B2(n4437), .A(n3446), .ZN(n3447) );
  OAI21_X1 U4244 ( .B1(n3448), .B2(n4475), .A(n3447), .ZN(n4478) );
  INV_X1 U4245 ( .A(n4478), .ZN(n3457) );
  XOR2_X1 U4246 ( .A(n3928), .B(n3449), .Z(n4479) );
  INV_X1 U4247 ( .A(n3450), .ZN(n3451) );
  OAI21_X1 U4248 ( .B1(n3452), .B2(n3792), .A(n3451), .ZN(n4547) );
  NOR2_X1 U4249 ( .A1(n4547), .A2(n4364), .ZN(n3455) );
  OAI22_X1 U4250 ( .A1(n4752), .A2(n3453), .B1(n3796), .B2(n4755), .ZN(n3454)
         );
  AOI211_X1 U4251 ( .C1(n4479), .C2(n4336), .A(n3455), .B(n3454), .ZN(n3456)
         );
  OAI21_X1 U4252 ( .B1(n3457), .B2(n4745), .A(n3456), .ZN(U3277) );
  NOR3_X1 U4253 ( .A1(n2707), .A2(n3458), .A3(n2708), .ZN(n3459) );
  AOI21_X1 U4254 ( .B1(n4767), .B2(n3460), .A(n3459), .ZN(U3458) );
  INV_X1 U4255 ( .A(DATAI_26_), .ZN(n3462) );
  NAND2_X1 U4256 ( .A1(n2708), .A2(STATE_REG_SCAN_IN), .ZN(n3461) );
  OAI21_X1 U4257 ( .B1(STATE_REG_SCAN_IN), .B2(n3462), .A(n3461), .ZN(U3326)
         );
  INV_X1 U4258 ( .A(n3463), .ZN(n3482) );
  AOI22_X1 U4259 ( .A1(n4059), .A2(REG1_REG_12__SCAN_IN), .B1(n4690), .B2(
        n2156), .ZN(n4072) );
  MUX2_X1 U4260 ( .A(REG1_REG_13__SCAN_IN), .B(n4481), .S(n4075), .Z(n4071) );
  OR2_X2 U4261 ( .A1(n4072), .A2(n4071), .ZN(n4073) );
  NAND2_X1 U4262 ( .A1(n3466), .A2(REG1_REG_13__SCAN_IN), .ZN(n3467) );
  INV_X1 U4263 ( .A(n4086), .ZN(n4689) );
  INV_X1 U4264 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4675) );
  MUX2_X1 U4265 ( .A(REG1_REG_15__SCAN_IN), .B(n4675), .S(n4100), .Z(n4092) );
  INV_X1 U4266 ( .A(n4106), .ZN(n4688) );
  NAND2_X1 U4267 ( .A1(n3469), .A2(n4688), .ZN(n3471) );
  NAND2_X1 U4268 ( .A1(n3470), .A2(n4106), .ZN(n3473) );
  AND2_X2 U4269 ( .A1(n3471), .A2(n3473), .ZN(n4103) );
  INV_X1 U4270 ( .A(REG1_REG_16__SCAN_IN), .ZN(n3472) );
  AND2_X2 U4271 ( .A1(n4103), .A2(n3472), .ZN(n4104) );
  INV_X1 U4272 ( .A(n3473), .ZN(n3474) );
  INV_X1 U4273 ( .A(n3495), .ZN(n4773) );
  AOI22_X1 U4274 ( .A1(n3495), .A2(n2513), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4773), .ZN(n4714) );
  INV_X1 U4275 ( .A(n3496), .ZN(n4771) );
  AOI22_X1 U4276 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3496), .B1(n4771), .B2(
        n3475), .ZN(n4732) );
  NAND2_X1 U4277 ( .A1(n4729), .A2(n2303), .ZN(n3479) );
  INV_X1 U4278 ( .A(REG1_REG_19__SCAN_IN), .ZN(n3476) );
  MUX2_X1 U4279 ( .A(n3476), .B(REG1_REG_19__SCAN_IN), .S(n4316), .Z(n3477) );
  INV_X1 U4280 ( .A(n3477), .ZN(n3478) );
  XNOR2_X1 U4281 ( .A(n3479), .B(n3478), .ZN(n3505) );
  INV_X1 U4282 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3480) );
  AOI22_X1 U4283 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4771), .B1(n3496), .B2(
        n3480), .ZN(n4720) );
  XNOR2_X1 U4284 ( .A(n3483), .B(n4690), .ZN(n4060) );
  INV_X1 U4285 ( .A(n3483), .ZN(n3484) );
  OAI21_X1 U4286 ( .B1(n3453), .B2(n4075), .A(n4070), .ZN(n3485) );
  OAI21_X1 U4287 ( .B1(REG2_REG_13__SCAN_IN), .B2(n3466), .A(n3485), .ZN(n3486) );
  INV_X1 U4288 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4082) );
  INV_X1 U4289 ( .A(n3486), .ZN(n3487) );
  NAND2_X1 U4290 ( .A1(n3487), .A2(n4689), .ZN(n3488) );
  MUX2_X1 U4291 ( .A(n3489), .B(REG2_REG_15__SCAN_IN), .S(n4100), .Z(n4095) );
  XNOR2_X1 U4292 ( .A(n3490), .B(n4106), .ZN(n4109) );
  NAND2_X1 U4293 ( .A1(n4109), .A2(n2505), .ZN(n3493) );
  INV_X1 U4294 ( .A(n3490), .ZN(n3491) );
  NOR2_X1 U4295 ( .A1(n3495), .A2(REG2_REG_17__SCAN_IN), .ZN(n3494) );
  AOI21_X1 U4296 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3495), .A(n3494), .ZN(n4711) );
  MUX2_X1 U4297 ( .A(REG2_REG_19__SCAN_IN), .B(n4561), .S(n4316), .Z(n3498) );
  XNOR2_X1 U4298 ( .A(n3499), .B(n3498), .ZN(n3503) );
  NAND2_X1 U4299 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3718) );
  NAND2_X1 U4300 ( .A1(n4722), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3500) );
  OAI211_X1 U4301 ( .C1(n4735), .C2(n3501), .A(n3718), .B(n3500), .ZN(n3502)
         );
  AOI21_X1 U4302 ( .B1(n3503), .B2(n4110), .A(n3502), .ZN(n3504) );
  OAI21_X1 U4303 ( .B1(n4114), .B2(n3505), .A(n3504), .ZN(U3259) );
  AND2_X1 U4304 ( .A1(n3506), .A2(DATAI_30_), .ZN(n4120) );
  NAND2_X1 U4305 ( .A1(n3506), .A2(DATAI_31_), .ZN(n3968) );
  XNOR2_X1 U4306 ( .A(n4118), .B(n3968), .ZN(n3520) );
  INV_X1 U4307 ( .A(REG2_REG_31__SCAN_IN), .ZN(n3509) );
  NAND2_X1 U4308 ( .A1(n2345), .A2(REG1_REG_31__SCAN_IN), .ZN(n3508) );
  INV_X1 U4309 ( .A(REG0_REG_31__SCAN_IN), .ZN(n3512) );
  OR2_X1 U4310 ( .A1(n2347), .A2(n3512), .ZN(n3507) );
  OAI211_X1 U4311 ( .C1(n3510), .C2(n3509), .A(n3508), .B(n3507), .ZN(n4012)
         );
  NAND2_X1 U4312 ( .A1(n3511), .A2(n4012), .ZN(n4117) );
  OAI21_X1 U4313 ( .B1(n4489), .B2(n3968), .A(n4117), .ZN(n3517) );
  NOR2_X1 U4314 ( .A1(n4783), .A2(n3512), .ZN(n3513) );
  AOI21_X1 U4315 ( .B1(n4783), .B2(n3517), .A(n3513), .ZN(n3514) );
  OAI21_X1 U4316 ( .B1(n3520), .B2(n4546), .A(n3514), .ZN(U3517) );
  NAND2_X1 U4317 ( .A1(n4752), .A2(n3517), .ZN(n3516) );
  NAND2_X1 U4318 ( .A1(n4745), .A2(REG2_REG_31__SCAN_IN), .ZN(n3515) );
  OAI211_X1 U4319 ( .C1(n3520), .C2(n4364), .A(n3516), .B(n3515), .ZN(U3260)
         );
  NAND2_X1 U4320 ( .A1(n4787), .A2(n3517), .ZN(n3519) );
  NAND2_X1 U4321 ( .A1(n4784), .A2(REG1_REG_31__SCAN_IN), .ZN(n3518) );
  OAI211_X1 U4322 ( .C1(n3520), .C2(n4483), .A(n3519), .B(n3518), .ZN(U3549)
         );
  OAI22_X1 U4323 ( .A1(n4414), .A2(n3655), .B1(n3650), .B2(n4241), .ZN(n3521)
         );
  XNOR2_X1 U4324 ( .A(n3521), .B(n3658), .ZN(n3607) );
  OAI22_X1 U4325 ( .A1(n4414), .A2(n3605), .B1(n3655), .B2(n4241), .ZN(n3606)
         );
  XNOR2_X1 U4326 ( .A(n3607), .B(n3606), .ZN(n3592) );
  NAND2_X1 U4327 ( .A1(n3523), .A2(n3522), .ZN(n3524) );
  OAI22_X1 U4328 ( .A1(n3605), .A2(n3739), .B1(n3655), .B2(n3803), .ZN(n3798)
         );
  OAI22_X1 U4329 ( .A1(n3739), .A2(n3655), .B1(n3650), .B2(n3803), .ZN(n3526)
         );
  XNOR2_X1 U4330 ( .A(n3526), .B(n3658), .ZN(n3799) );
  OR2_X1 U4331 ( .A1(n3655), .A2(n3802), .ZN(n3527) );
  OAI21_X1 U4332 ( .B1(n3650), .B2(n4490), .A(n3527), .ZN(n3528) );
  XNOR2_X1 U4333 ( .A(n3528), .B(n3658), .ZN(n3530) );
  OAI22_X1 U4334 ( .A1(n3605), .A2(n3802), .B1(n3655), .B2(n4490), .ZN(n3529)
         );
  NAND2_X1 U4335 ( .A1(n3530), .A2(n3529), .ZN(n3733) );
  OR2_X1 U4336 ( .A1(n3655), .A2(n3702), .ZN(n3531) );
  OAI21_X1 U4337 ( .B1(n3650), .B2(n3792), .A(n3531), .ZN(n3532) );
  XNOR2_X1 U4338 ( .A(n3532), .B(n3645), .ZN(n3788) );
  NAND2_X1 U4339 ( .A1(n3533), .A2(n4487), .ZN(n3536) );
  NAND2_X1 U4340 ( .A1(n3174), .A2(n3534), .ZN(n3535) );
  AND2_X1 U4341 ( .A1(n3536), .A2(n3535), .ZN(n3540) );
  OAI22_X1 U4342 ( .A1(n3650), .A2(n4470), .B1(n3655), .B2(n4368), .ZN(n3537)
         );
  XNOR2_X1 U4343 ( .A(n3537), .B(n3658), .ZN(n3542) );
  OAI22_X1 U4344 ( .A1(n3605), .A2(n4368), .B1(n4470), .B2(n3604), .ZN(n3541)
         );
  NAND2_X1 U4345 ( .A1(n3542), .A2(n3541), .ZN(n3695) );
  INV_X1 U4346 ( .A(n3788), .ZN(n3692) );
  INV_X1 U4347 ( .A(n3540), .ZN(n3789) );
  NOR2_X1 U4348 ( .A1(n3692), .A2(n3789), .ZN(n3543) );
  NOR2_X1 U4349 ( .A1(n3542), .A2(n3541), .ZN(n3697) );
  AOI21_X1 U4350 ( .B1(n3543), .B2(n3695), .A(n3697), .ZN(n3544) );
  NAND2_X1 U4351 ( .A1(n3545), .A2(n3544), .ZN(n3746) );
  NAND2_X1 U4352 ( .A1(n4361), .A2(n3174), .ZN(n3547) );
  NAND2_X1 U4353 ( .A1(n3533), .A2(n4467), .ZN(n3546) );
  NAND2_X1 U4354 ( .A1(n3547), .A2(n3546), .ZN(n3836) );
  OAI22_X1 U4355 ( .A1(n4350), .A2(n3655), .B1(n4459), .B2(n3650), .ZN(n3548)
         );
  XNOR2_X1 U4356 ( .A(n3548), .B(n3658), .ZN(n3747) );
  NAND2_X1 U4357 ( .A1(n4456), .A2(n3174), .ZN(n3549) );
  OAI21_X1 U4358 ( .B1(n4449), .B2(n3650), .A(n3549), .ZN(n3550) );
  XNOR2_X1 U4359 ( .A(n3550), .B(n3658), .ZN(n3745) );
  NAND2_X1 U4360 ( .A1(n3533), .A2(n4456), .ZN(n3551) );
  OAI21_X1 U4361 ( .B1(n4449), .B2(n3604), .A(n3551), .ZN(n3744) );
  AND2_X1 U4362 ( .A1(n3745), .A2(n3744), .ZN(n3556) );
  AOI21_X1 U4363 ( .B1(n3836), .B2(n3747), .A(n3556), .ZN(n3553) );
  OAI22_X1 U4364 ( .A1(n3751), .A2(n3655), .B1(n3650), .B2(n4329), .ZN(n3554)
         );
  XNOR2_X1 U4365 ( .A(n3554), .B(n3645), .ZN(n3759) );
  NOR2_X1 U4366 ( .A1(n3655), .A2(n4329), .ZN(n3555) );
  AOI21_X1 U4367 ( .B1(n4447), .B2(n3533), .A(n3555), .ZN(n3558) );
  NOR2_X1 U4368 ( .A1(n3745), .A2(n3744), .ZN(n3756) );
  NOR3_X1 U4369 ( .A1(n3556), .A2(n3836), .A3(n3747), .ZN(n3557) );
  AOI211_X1 U4370 ( .C1(n3759), .C2(n3558), .A(n3756), .B(n3557), .ZN(n3560)
         );
  INV_X1 U4371 ( .A(n3759), .ZN(n3559) );
  INV_X1 U4372 ( .A(n3558), .ZN(n3758) );
  OAI22_X1 U4373 ( .A1(n4440), .A2(n3655), .B1(n3650), .B2(n4308), .ZN(n3561)
         );
  XNOR2_X1 U4374 ( .A(n3561), .B(n3658), .ZN(n3562) );
  OAI22_X1 U4375 ( .A1(n4440), .A2(n3605), .B1(n3655), .B2(n4308), .ZN(n3563)
         );
  NAND2_X1 U4376 ( .A1(n3562), .A2(n3563), .ZN(n3811) );
  INV_X1 U4377 ( .A(n3562), .ZN(n3565) );
  INV_X1 U4378 ( .A(n3563), .ZN(n3564) );
  NAND2_X1 U4379 ( .A1(n3565), .A2(n3564), .ZN(n3810) );
  OAI22_X1 U4380 ( .A1(n4313), .A2(n3605), .B1(n3655), .B2(n4296), .ZN(n3570)
         );
  NAND2_X1 U4381 ( .A1(n4421), .A2(n3174), .ZN(n3567) );
  NAND2_X1 U4382 ( .A1(n3660), .A2(n4288), .ZN(n3566) );
  NAND2_X1 U4383 ( .A1(n3567), .A2(n3566), .ZN(n3568) );
  XNOR2_X1 U4384 ( .A(n3568), .B(n3658), .ZN(n3569) );
  XOR2_X1 U4385 ( .A(n3570), .B(n3569), .Z(n3717) );
  NAND2_X1 U4386 ( .A1(n3716), .A2(n3717), .ZN(n3574) );
  NAND2_X1 U4387 ( .A1(n3574), .A2(n3573), .ZN(n3776) );
  NAND2_X1 U4388 ( .A1(n4411), .A2(n3174), .ZN(n3576) );
  OR2_X1 U4389 ( .A1(n3650), .A2(n4275), .ZN(n3575) );
  NAND2_X1 U4390 ( .A1(n3576), .A2(n3575), .ZN(n3577) );
  XNOR2_X1 U4391 ( .A(n3577), .B(n3658), .ZN(n3580) );
  NAND2_X1 U4392 ( .A1(n4411), .A2(n3533), .ZN(n3579) );
  NAND2_X1 U4393 ( .A1(n3174), .A2(n4420), .ZN(n3578) );
  NAND2_X1 U4394 ( .A1(n3579), .A2(n3578), .ZN(n3581) );
  NAND2_X1 U4395 ( .A1(n3580), .A2(n3581), .ZN(n3777) );
  INV_X1 U4396 ( .A(n3580), .ZN(n3583) );
  INV_X1 U4397 ( .A(n3581), .ZN(n3582) );
  NAND2_X1 U4398 ( .A1(n3583), .A2(n3582), .ZN(n3779) );
  NAND2_X1 U4399 ( .A1(n4230), .A2(n3174), .ZN(n3585) );
  OR2_X1 U4400 ( .A1(n3650), .A2(n4255), .ZN(n3584) );
  NAND2_X1 U4401 ( .A1(n3585), .A2(n3584), .ZN(n3586) );
  XNOR2_X1 U4402 ( .A(n3586), .B(n3658), .ZN(n3725) );
  NAND2_X1 U4403 ( .A1(n4230), .A2(n3533), .ZN(n3588) );
  NAND2_X1 U4404 ( .A1(n3174), .A2(n4410), .ZN(n3587) );
  NAND2_X1 U4405 ( .A1(n3588), .A2(n3587), .ZN(n3724) );
  NAND2_X1 U4406 ( .A1(n3725), .A2(n3724), .ZN(n3589) );
  INV_X1 U4407 ( .A(n3609), .ZN(n3709) );
  AOI21_X1 U4408 ( .B1(n3592), .B2(n3591), .A(n3709), .ZN(n3598) );
  INV_X1 U4409 ( .A(n4242), .ZN(n3596) );
  INV_X1 U4410 ( .A(n4230), .ZN(n4424) );
  OAI22_X1 U4411 ( .A1(n2003), .A2(n4241), .B1(n4424), .B2(n3783), .ZN(n3595)
         );
  OAI22_X1 U4412 ( .A1(n4233), .A2(n3840), .B1(STATE_REG_SCAN_IN), .B2(n3593), 
        .ZN(n3594) );
  AOI211_X1 U4413 ( .C1(n3596), .C2(n3829), .A(n3595), .B(n3594), .ZN(n3597)
         );
  OAI21_X1 U4414 ( .B1(n3598), .B2(n3831), .A(n3597), .ZN(U3232) );
  NAND3_X1 U4415 ( .A1(n3600), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3602) );
  INV_X1 U4416 ( .A(DATAI_31_), .ZN(n3601) );
  OAI22_X1 U4417 ( .A1(n3599), .A2(n3602), .B1(STATE_REG_SCAN_IN), .B2(n3601), 
        .ZN(U3321) );
  OAI22_X1 U4418 ( .A1(n4233), .A2(n3604), .B1(n3650), .B2(n4215), .ZN(n3603)
         );
  XNOR2_X1 U4419 ( .A(n3603), .B(n3658), .ZN(n3611) );
  OAI22_X1 U4420 ( .A1(n4233), .A2(n3605), .B1(n3655), .B2(n4215), .ZN(n3610)
         );
  XNOR2_X1 U4421 ( .A(n3611), .B(n3610), .ZN(n3707) );
  NOR2_X1 U4422 ( .A1(n3607), .A2(n3606), .ZN(n3708) );
  NOR2_X1 U4423 ( .A1(n3707), .A2(n3708), .ZN(n3608) );
  NAND2_X1 U4424 ( .A1(n3611), .A2(n3610), .ZN(n3630) );
  NOR2_X1 U4425 ( .A1(n3655), .A2(n4197), .ZN(n3612) );
  AOI21_X1 U4426 ( .B1(n4016), .B2(n3533), .A(n3612), .ZN(n3636) );
  NAND2_X1 U4427 ( .A1(n3630), .A2(n3636), .ZN(n3633) );
  INV_X1 U4428 ( .A(n3633), .ZN(n3614) );
  NAND2_X1 U4429 ( .A1(n4016), .A2(n3174), .ZN(n3616) );
  OR2_X1 U4430 ( .A1(n3650), .A2(n4197), .ZN(n3615) );
  NAND2_X1 U4431 ( .A1(n3616), .A2(n3615), .ZN(n3617) );
  XNOR2_X1 U4432 ( .A(n3617), .B(n3645), .ZN(n3635) );
  INV_X1 U4433 ( .A(n3635), .ZN(n3768) );
  NOR2_X1 U4434 ( .A1(n3604), .A2(n4182), .ZN(n3618) );
  AOI21_X1 U4435 ( .B1(n3824), .B2(n3533), .A(n3618), .ZN(n3637) );
  AOI22_X1 U4436 ( .A1(n3824), .A2(n3174), .B1(n3660), .B2(n4382), .ZN(n3619)
         );
  XNOR2_X1 U4437 ( .A(n3619), .B(n3658), .ZN(n3634) );
  NOR2_X1 U4438 ( .A1(n3634), .A2(n3637), .ZN(n3631) );
  AOI21_X1 U4439 ( .B1(n3637), .B2(n3634), .A(n3631), .ZN(n3620) );
  XNOR2_X1 U4440 ( .A(n3622), .B(n3621), .ZN(n3623) );
  NAND2_X1 U4441 ( .A1(n3623), .A2(n3838), .ZN(n3629) );
  INV_X1 U4442 ( .A(n3624), .ZN(n4180) );
  INV_X1 U4443 ( .A(n4016), .ZN(n4387) );
  OAI22_X1 U4444 ( .A1(n4387), .A2(n3783), .B1(STATE_REG_SCAN_IN), .B2(n3625), 
        .ZN(n3627) );
  OAI22_X1 U4445 ( .A1(n4183), .A2(n3840), .B1(n2003), .B2(n4182), .ZN(n3626)
         );
  AOI211_X1 U4446 ( .C1(n4180), .C2(n3829), .A(n3627), .B(n3626), .ZN(n3628)
         );
  NAND2_X1 U4447 ( .A1(n3629), .A2(n3628), .ZN(U3222) );
  NAND2_X1 U4448 ( .A1(n3630), .A2(n3635), .ZN(n3632) );
  AOI21_X1 U4449 ( .B1(n3633), .B2(n3632), .A(n3631), .ZN(n3642) );
  INV_X1 U4450 ( .A(n3634), .ZN(n3640) );
  AOI21_X1 U4451 ( .B1(n3635), .B2(n3636), .A(n3637), .ZN(n3639) );
  NAND2_X1 U4452 ( .A1(n3637), .A2(n3636), .ZN(n3638) );
  OAI22_X1 U4453 ( .A1(n3640), .A2(n3639), .B1(n3768), .B2(n3638), .ZN(n3641)
         );
  NAND2_X1 U4454 ( .A1(n4383), .A2(n3174), .ZN(n3644) );
  OR2_X1 U4455 ( .A1(n3650), .A2(n3827), .ZN(n3643) );
  NAND2_X1 U4456 ( .A1(n3644), .A2(n3643), .ZN(n3646) );
  XNOR2_X1 U4457 ( .A(n3646), .B(n3645), .ZN(n3649) );
  NOR2_X1 U4458 ( .A1(n3604), .A2(n3827), .ZN(n3647) );
  AOI21_X1 U4459 ( .B1(n4383), .B2(n3533), .A(n3647), .ZN(n3648) );
  NOR2_X1 U4460 ( .A1(n3649), .A2(n3648), .ZN(n3820) );
  NAND2_X1 U4461 ( .A1(n3649), .A2(n3648), .ZN(n3818) );
  NAND2_X1 U4462 ( .A1(n4015), .A2(n3174), .ZN(n3652) );
  OR2_X1 U4463 ( .A1(n3650), .A2(n4154), .ZN(n3651) );
  NAND2_X1 U4464 ( .A1(n3652), .A2(n3651), .ZN(n3653) );
  XNOR2_X1 U4465 ( .A(n3653), .B(n3658), .ZN(n3666) );
  NOR2_X1 U4466 ( .A1(n3655), .A2(n4154), .ZN(n3654) );
  AOI21_X1 U4467 ( .B1(n4015), .B2(n3533), .A(n3654), .ZN(n3664) );
  XNOR2_X1 U4468 ( .A(n3666), .B(n3664), .ZN(n3682) );
  NAND2_X1 U4469 ( .A1(n4014), .A2(n3533), .ZN(n3657) );
  OR2_X1 U4470 ( .A1(n3655), .A2(n4139), .ZN(n3656) );
  NAND2_X1 U4471 ( .A1(n3657), .A2(n3656), .ZN(n3659) );
  XNOR2_X1 U4472 ( .A(n3659), .B(n3658), .ZN(n3662) );
  AOI22_X1 U4473 ( .A1(n4014), .A2(n3174), .B1(n3660), .B2(n3670), .ZN(n3661)
         );
  XNOR2_X1 U4474 ( .A(n3662), .B(n3661), .ZN(n3674) );
  INV_X1 U4475 ( .A(n3674), .ZN(n3663) );
  NAND2_X1 U4476 ( .A1(n3663), .A2(n3838), .ZN(n3680) );
  INV_X1 U4477 ( .A(n3664), .ZN(n3665) );
  NAND2_X1 U4478 ( .A1(n3666), .A2(n3665), .ZN(n3673) );
  INV_X1 U4479 ( .A(n3673), .ZN(n3667) );
  NAND2_X1 U4480 ( .A1(n3681), .A2(n3669), .ZN(n3679) );
  INV_X1 U4481 ( .A(n4138), .ZN(n3677) );
  AOI22_X1 U4482 ( .A1(n4143), .A2(n3823), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3672) );
  NAND2_X1 U4483 ( .A1(n3737), .A2(n3670), .ZN(n3671) );
  OAI211_X1 U4484 ( .C1(n4140), .C2(n3783), .A(n3672), .B(n3671), .ZN(n3676)
         );
  NOR3_X1 U4485 ( .A1(n3674), .A2(n3831), .A3(n3673), .ZN(n3675) );
  AOI211_X1 U4486 ( .C1(n3677), .C2(n3829), .A(n3676), .B(n3675), .ZN(n3678)
         );
  OAI211_X1 U4487 ( .C1(n3681), .C2(n3680), .A(n3679), .B(n3678), .ZN(U3217)
         );
  XNOR2_X1 U4488 ( .A(n3683), .B(n3682), .ZN(n3684) );
  NAND2_X1 U4489 ( .A1(n3684), .A2(n3838), .ZN(n3689) );
  OAI22_X1 U4490 ( .A1(n4183), .A2(n3783), .B1(n2003), .B2(n4154), .ZN(n3687)
         );
  OAI22_X1 U4491 ( .A1(n4155), .A2(n3840), .B1(STATE_REG_SCAN_IN), .B2(n3685), 
        .ZN(n3686) );
  AOI211_X1 U4492 ( .C1(n4152), .C2(n3829), .A(n3687), .B(n3686), .ZN(n3688)
         );
  NAND2_X1 U4493 ( .A1(n3689), .A2(n3688), .ZN(U3211) );
  INV_X1 U4494 ( .A(n3691), .ZN(n3693) );
  OAI21_X1 U4495 ( .B1(n3693), .B2(n3692), .A(n3789), .ZN(n3694) );
  OAI21_X1 U4496 ( .B1(n3788), .B2(n3691), .A(n3694), .ZN(n3699) );
  INV_X1 U4497 ( .A(n3695), .ZN(n3696) );
  NOR2_X1 U4498 ( .A1(n3697), .A2(n3696), .ZN(n3698) );
  XNOR2_X1 U4499 ( .A(n3699), .B(n3698), .ZN(n3706) );
  AOI22_X1 U4500 ( .A1(n3737), .A2(n3700), .B1(n3823), .B2(n4467), .ZN(n3701)
         );
  NAND2_X1 U4501 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n4085) );
  OAI211_X1 U4502 ( .C1(n3702), .C2(n3783), .A(n3701), .B(n4085), .ZN(n3703)
         );
  AOI21_X1 U4503 ( .B1(n3704), .B2(n3829), .A(n3703), .ZN(n3705) );
  OAI21_X1 U4504 ( .B1(n3706), .B2(n3831), .A(n3705), .ZN(U3212) );
  OAI21_X1 U4505 ( .B1(n3709), .B2(n3708), .A(n3707), .ZN(n3711) );
  NAND3_X1 U4506 ( .A1(n3711), .A2(n3838), .A3(n3710), .ZN(n3715) );
  OAI22_X1 U4507 ( .A1(n4387), .A2(n3840), .B1(STATE_REG_SCAN_IN), .B2(n4663), 
        .ZN(n3713) );
  OAI22_X1 U4508 ( .A1(n2003), .A2(n4215), .B1(n4414), .B2(n3783), .ZN(n3712)
         );
  NOR2_X1 U4509 ( .A1(n3713), .A2(n3712), .ZN(n3714) );
  OAI211_X1 U4510 ( .C1(n3846), .C2(n4217), .A(n3715), .B(n3714), .ZN(U3213)
         );
  XOR2_X1 U4511 ( .A(n3717), .B(n3716), .Z(n3722) );
  INV_X1 U4512 ( .A(n4411), .ZN(n4292) );
  AOI22_X1 U4513 ( .A1(n3737), .A2(n4288), .B1(n3843), .B2(n4289), .ZN(n3719)
         );
  OAI211_X1 U4514 ( .C1(n4292), .C2(n3840), .A(n3719), .B(n3718), .ZN(n3720)
         );
  AOI21_X1 U4515 ( .B1(n4298), .B2(n3829), .A(n3720), .ZN(n3721) );
  OAI21_X1 U4516 ( .B1(n3722), .B2(n3831), .A(n3721), .ZN(U3216) );
  XNOR2_X1 U4517 ( .A(n3725), .B(n3724), .ZN(n3726) );
  XNOR2_X1 U4518 ( .A(n3723), .B(n3726), .ZN(n3731) );
  OAI22_X1 U4519 ( .A1(n4414), .A2(n3840), .B1(STATE_REG_SCAN_IN), .B2(n3727), 
        .ZN(n3729) );
  OAI22_X1 U4520 ( .A1(n2003), .A2(n4255), .B1(n4292), .B2(n3783), .ZN(n3728)
         );
  AOI211_X1 U4521 ( .C1(n4253), .C2(n3829), .A(n3729), .B(n3728), .ZN(n3730)
         );
  OAI21_X1 U4522 ( .B1(n3731), .B2(n3831), .A(n3730), .ZN(U3220) );
  NAND2_X1 U4523 ( .A1(n3734), .A2(n3733), .ZN(n3735) );
  XNOR2_X1 U4524 ( .A(n3732), .B(n3735), .ZN(n3743) );
  AOI22_X1 U4525 ( .A1(n3737), .A2(n3736), .B1(n3823), .B2(n4487), .ZN(n3738)
         );
  NAND2_X1 U4526 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n4062) );
  OAI211_X1 U4527 ( .C1(n3739), .C2(n3783), .A(n3738), .B(n4062), .ZN(n3740)
         );
  AOI21_X1 U4528 ( .B1(n3741), .B2(n3829), .A(n3740), .ZN(n3742) );
  OAI21_X1 U4529 ( .B1(n3743), .B2(n3831), .A(n3742), .ZN(U3221) );
  XNOR2_X1 U4530 ( .A(n3745), .B(n3744), .ZN(n3755) );
  INV_X1 U4531 ( .A(n3747), .ZN(n3748) );
  NOR2_X1 U4532 ( .A1(n3746), .A2(n3748), .ZN(n3833) );
  NAND2_X1 U4533 ( .A1(n3746), .A2(n3748), .ZN(n3834) );
  OAI21_X1 U4534 ( .B1(n3833), .B2(n3836), .A(n3834), .ZN(n3749) );
  XOR2_X1 U4535 ( .A(n3755), .B(n3749), .Z(n3750) );
  NAND2_X1 U4536 ( .A1(n3750), .A2(n3838), .ZN(n3754) );
  AND2_X1 U4537 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4108) );
  OAI22_X1 U4538 ( .A1(n2003), .A2(n4449), .B1(n3751), .B2(n3840), .ZN(n3752)
         );
  AOI211_X1 U4539 ( .C1(n3843), .C2(n4467), .A(n4108), .B(n3752), .ZN(n3753)
         );
  OAI211_X1 U4540 ( .C1(n3846), .C2(n4346), .A(n3754), .B(n3753), .ZN(U3223)
         );
  AOI211_X1 U4541 ( .C1(n3836), .C2(n3834), .A(n3755), .B(n3833), .ZN(n3757)
         );
  NOR2_X1 U4542 ( .A1(n3757), .A2(n3756), .ZN(n3761) );
  XNOR2_X1 U4543 ( .A(n3759), .B(n3758), .ZN(n3760) );
  XNOR2_X1 U4544 ( .A(n3761), .B(n3760), .ZN(n3765) );
  NOR2_X1 U4545 ( .A1(n4651), .A2(STATE_REG_SCAN_IN), .ZN(n4713) );
  OAI22_X1 U4546 ( .A1(n2003), .A2(n4329), .B1(n4440), .B2(n3840), .ZN(n3762)
         );
  AOI211_X1 U4547 ( .C1(n3843), .C2(n4456), .A(n4713), .B(n3762), .ZN(n3764)
         );
  NAND2_X1 U4548 ( .A1(n3829), .A2(n4330), .ZN(n3763) );
  OAI211_X1 U4549 ( .C1(n3765), .C2(n3831), .A(n3764), .B(n3763), .ZN(U3225)
         );
  XNOR2_X1 U4550 ( .A(n3769), .B(n3768), .ZN(n3774) );
  OAI22_X1 U4551 ( .A1(n4233), .A2(n3783), .B1(STATE_REG_SCAN_IN), .B2(n3770), 
        .ZN(n3772) );
  INV_X1 U4552 ( .A(n3824), .ZN(n4396) );
  OAI22_X1 U4553 ( .A1(n4396), .A2(n3840), .B1(n2003), .B2(n4197), .ZN(n3771)
         );
  AOI211_X1 U4554 ( .C1(n4195), .C2(n3829), .A(n3772), .B(n3771), .ZN(n3773)
         );
  OAI21_X1 U4555 ( .B1(n3774), .B2(n3831), .A(n3773), .ZN(U3226) );
  INV_X1 U4556 ( .A(n3775), .ZN(n3780) );
  AOI21_X1 U4557 ( .B1(n3779), .B2(n3777), .A(n3776), .ZN(n3778) );
  AOI21_X1 U4558 ( .B1(n3780), .B2(n3779), .A(n3778), .ZN(n3787) );
  INV_X1 U4559 ( .A(n3781), .ZN(n4273) );
  OAI22_X1 U4560 ( .A1(n4424), .A2(n3840), .B1(STATE_REG_SCAN_IN), .B2(n3782), 
        .ZN(n3785) );
  OAI22_X1 U4561 ( .A1(n2003), .A2(n4275), .B1(n4313), .B2(n3783), .ZN(n3784)
         );
  AOI211_X1 U4562 ( .C1(n4273), .C2(n3829), .A(n3785), .B(n3784), .ZN(n3786)
         );
  OAI21_X1 U4563 ( .B1(n3787), .B2(n3831), .A(n3786), .ZN(U3230) );
  XNOR2_X1 U4564 ( .A(n3789), .B(n3788), .ZN(n3790) );
  XNOR2_X1 U4565 ( .A(n3691), .B(n3790), .ZN(n3791) );
  NAND2_X1 U4566 ( .A1(n3791), .A2(n3838), .ZN(n3795) );
  AND2_X1 U4567 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4077) );
  OAI22_X1 U4568 ( .A1(n2003), .A2(n3792), .B1(n4368), .B2(n3840), .ZN(n3793)
         );
  AOI211_X1 U4569 ( .C1(n3843), .C2(n4017), .A(n4077), .B(n3793), .ZN(n3794)
         );
  OAI211_X1 U4570 ( .C1(n3846), .C2(n3796), .A(n3795), .B(n3794), .ZN(U3231)
         );
  XNOR2_X1 U4571 ( .A(n3799), .B(n3798), .ZN(n3800) );
  XNOR2_X1 U4572 ( .A(n3797), .B(n3800), .ZN(n3801) );
  NAND2_X1 U4573 ( .A1(n3801), .A2(n3838), .ZN(n3808) );
  OAI22_X1 U4574 ( .A1(n2003), .A2(n3803), .B1(n3802), .B2(n3840), .ZN(n3804)
         );
  AOI211_X1 U4575 ( .C1(n3843), .C2(n3806), .A(n3805), .B(n3804), .ZN(n3807)
         );
  OAI211_X1 U4576 ( .C1(n3846), .C2(n3809), .A(n3808), .B(n3807), .ZN(U3233)
         );
  NAND2_X1 U4577 ( .A1(n3811), .A2(n3810), .ZN(n3813) );
  XOR2_X1 U4578 ( .A(n3813), .B(n3812), .Z(n3814) );
  NAND2_X1 U4579 ( .A1(n3814), .A2(n3838), .ZN(n3817) );
  AND2_X1 U4580 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4723) );
  OAI22_X1 U4581 ( .A1(n2003), .A2(n4308), .B1(n4313), .B2(n3840), .ZN(n3815)
         );
  AOI211_X1 U4582 ( .C1(n3843), .C2(n4447), .A(n4723), .B(n3815), .ZN(n3816)
         );
  OAI211_X1 U4583 ( .C1(n3846), .C2(n4318), .A(n3817), .B(n3816), .ZN(U3235)
         );
  INV_X1 U4584 ( .A(n3818), .ZN(n3819) );
  NOR2_X1 U4585 ( .A1(n3820), .A2(n3819), .ZN(n3821) );
  XNOR2_X1 U4586 ( .A(n3822), .B(n3821), .ZN(n3832) );
  NAND2_X1 U4587 ( .A1(n4015), .A2(n3823), .ZN(n3826) );
  AOI22_X1 U4588 ( .A1(n3824), .A2(n3843), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3825) );
  OAI211_X1 U4589 ( .C1(n2003), .C2(n3827), .A(n3826), .B(n3825), .ZN(n3828)
         );
  AOI21_X1 U4590 ( .B1(n4163), .B2(n3829), .A(n3828), .ZN(n3830) );
  OAI21_X1 U4591 ( .B1(n3832), .B2(n3831), .A(n3830), .ZN(U3237) );
  INV_X1 U4592 ( .A(n3833), .ZN(n3835) );
  NAND2_X1 U4593 ( .A1(n3835), .A2(n3834), .ZN(n3837) );
  XNOR2_X1 U4594 ( .A(n3837), .B(n3836), .ZN(n3839) );
  NAND2_X1 U4595 ( .A1(n3839), .A2(n3838), .ZN(n3845) );
  AND2_X1 U4596 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4097) );
  OAI22_X1 U4597 ( .A1(n2003), .A2(n4459), .B1(n4372), .B2(n3840), .ZN(n3842)
         );
  AOI211_X1 U4598 ( .C1(n3843), .C2(n4455), .A(n4097), .B(n3842), .ZN(n3844)
         );
  OAI211_X1 U4599 ( .C1(n3846), .C2(n4365), .A(n3845), .B(n3844), .ZN(U3238)
         );
  OAI211_X1 U4600 ( .C1(n2662), .C2(n4687), .A(n3849), .B(n3848), .ZN(n3852)
         );
  NAND3_X1 U4601 ( .A1(n3852), .A2(n3851), .A3(n3850), .ZN(n3855) );
  NAND3_X1 U4602 ( .A1(n3855), .A2(n3854), .A3(n3853), .ZN(n3858) );
  NAND3_X1 U4603 ( .A1(n3858), .A2(n3857), .A3(n3856), .ZN(n3859) );
  NAND4_X1 U4604 ( .A1(n3860), .A2(n3859), .A3(n3875), .A4(n2110), .ZN(n3862)
         );
  NAND3_X1 U4605 ( .A1(n3862), .A2(n3947), .A3(n3861), .ZN(n3863) );
  NAND3_X1 U4606 ( .A1(n3863), .A2(n3872), .A3(n3876), .ZN(n3866) );
  NAND3_X1 U4607 ( .A1(n3866), .A2(n3865), .A3(n3864), .ZN(n3867) );
  AND4_X1 U4608 ( .A1(n3867), .A2(n3878), .A3(n3879), .A4(n2042), .ZN(n3885)
         );
  NOR2_X1 U4609 ( .A1(n3868), .A2(n3931), .ZN(n3870) );
  AND2_X1 U4610 ( .A1(n3870), .A2(n3869), .ZN(n3894) );
  AND2_X1 U4611 ( .A1(n3894), .A2(n3871), .ZN(n3975) );
  INV_X1 U4612 ( .A(n3872), .ZN(n3874) );
  NOR2_X1 U4613 ( .A1(n3874), .A2(n3873), .ZN(n3877) );
  NAND4_X1 U4614 ( .A1(n3877), .A2(n2042), .A3(n3876), .A4(n3875), .ZN(n3882)
         );
  NAND2_X1 U4615 ( .A1(n3879), .A2(n3878), .ZN(n3880) );
  NAND2_X1 U4616 ( .A1(n3892), .A2(n3880), .ZN(n3881) );
  NAND2_X1 U4617 ( .A1(n3975), .A2(n3881), .ZN(n3972) );
  AOI21_X1 U4618 ( .B1(n3883), .B2(n3882), .A(n3972), .ZN(n3884) );
  AOI21_X1 U4619 ( .B1(n3885), .B2(n3975), .A(n3884), .ZN(n3890) );
  INV_X1 U4620 ( .A(n3886), .ZN(n3888) );
  NOR4_X1 U4621 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n3898)
         );
  AND2_X1 U4622 ( .A1(n3892), .A2(n3891), .ZN(n3973) );
  AOI21_X1 U4623 ( .B1(n3893), .B2(n3973), .A(n3972), .ZN(n3897) );
  INV_X1 U4624 ( .A(n3894), .ZN(n3895) );
  OAI21_X1 U4625 ( .B1(n3979), .B2(n3895), .A(n3977), .ZN(n3896) );
  OR3_X1 U4626 ( .A1(n3898), .A2(n3897), .A3(n3896), .ZN(n3900) );
  INV_X1 U4627 ( .A(n3899), .ZN(n4204) );
  AOI21_X1 U4628 ( .B1(n3900), .B2(n4204), .A(n3976), .ZN(n3904) );
  INV_X1 U4629 ( .A(n3922), .ZN(n3901) );
  NOR2_X1 U4630 ( .A1(n3901), .A2(n3925), .ZN(n3985) );
  OAI211_X1 U4631 ( .C1(n3904), .C2(n3903), .A(n3902), .B(n3985), .ZN(n3910)
         );
  INV_X1 U4632 ( .A(n3905), .ZN(n3906) );
  AOI21_X1 U4633 ( .B1(n4143), .B2(n3914), .A(n3906), .ZN(n3971) );
  INV_X1 U4634 ( .A(n3971), .ZN(n3908) );
  AOI211_X1 U4635 ( .C1(n4015), .C2(n4154), .A(n3908), .B(n3907), .ZN(n3909)
         );
  NAND2_X1 U4636 ( .A1(n3910), .A2(n3909), .ZN(n3919) );
  NAND2_X1 U4637 ( .A1(n4012), .A2(n3968), .ZN(n3918) );
  INV_X1 U4638 ( .A(n4120), .ZN(n3915) );
  OR2_X1 U4639 ( .A1(n4013), .A2(n3915), .ZN(n3913) );
  AND2_X1 U4640 ( .A1(n3918), .A2(n3913), .ZN(n3941) );
  OAI21_X1 U4641 ( .B1(n4143), .B2(n3914), .A(n3941), .ZN(n3987) );
  AOI21_X1 U4642 ( .B1(n3971), .B2(n3989), .A(n3987), .ZN(n3993) );
  NOR2_X1 U4643 ( .A1(n4012), .A2(n3968), .ZN(n3996) );
  INV_X1 U4644 ( .A(n3996), .ZN(n3917) );
  AND2_X1 U4645 ( .A1(n4013), .A2(n3915), .ZN(n3997) );
  INV_X1 U4646 ( .A(n3997), .ZN(n3916) );
  NAND2_X1 U4647 ( .A1(n3917), .A2(n3916), .ZN(n3943) );
  AOI22_X1 U4648 ( .A1(n3919), .A2(n3993), .B1(n3918), .B2(n3943), .ZN(n4001)
         );
  NAND2_X1 U4649 ( .A1(n3921), .A2(n3920), .ZN(n4175) );
  INV_X1 U4650 ( .A(n4175), .ZN(n3962) );
  NAND2_X1 U4651 ( .A1(n3922), .A2(n4170), .ZN(n4192) );
  INV_X1 U4652 ( .A(n4192), .ZN(n3961) );
  INV_X1 U4653 ( .A(n3923), .ZN(n3924) );
  OR2_X1 U4654 ( .A1(n3925), .A2(n3924), .ZN(n4207) );
  NAND2_X1 U4655 ( .A1(n3927), .A2(n3926), .ZN(n4294) );
  INV_X1 U4656 ( .A(n4294), .ZN(n3930) );
  NAND3_X1 U4657 ( .A1(n3930), .A2(n3929), .A3(n3928), .ZN(n3955) );
  NAND2_X1 U4658 ( .A1(n2673), .A2(n4281), .ZN(n4324) );
  NOR3_X1 U4659 ( .A1(n4324), .A2(n3932), .A3(n4357), .ZN(n3953) );
  INV_X1 U4660 ( .A(n4304), .ZN(n4309) );
  NAND4_X1 U4661 ( .A1(n3936), .A2(n3935), .A3(n3934), .A4(n3933), .ZN(n3950)
         );
  NAND4_X1 U4662 ( .A1(n3940), .A2(n3939), .A3(n3938), .A4(n3937), .ZN(n3949)
         );
  INV_X1 U4663 ( .A(n3941), .ZN(n3942) );
  NOR2_X1 U4664 ( .A1(n3943), .A2(n3942), .ZN(n3944) );
  NAND4_X1 U4665 ( .A1(n3947), .A2(n3946), .A3(n3945), .A4(n3944), .ZN(n3948)
         );
  NOR3_X1 U4666 ( .A1(n3950), .A2(n3949), .A3(n3948), .ZN(n3952) );
  NAND4_X1 U4667 ( .A1(n3953), .A2(n4309), .A3(n3952), .A4(n3951), .ZN(n3954)
         );
  NOR2_X1 U4668 ( .A1(n3955), .A2(n3954), .ZN(n3956) );
  NAND2_X1 U4669 ( .A1(n4237), .A2(n3956), .ZN(n3957) );
  NOR2_X1 U4670 ( .A1(n4207), .A2(n3957), .ZN(n3960) );
  AND2_X1 U4671 ( .A1(n4204), .A2(n4223), .ZN(n4251) );
  XNOR2_X1 U4672 ( .A(n4411), .B(n4275), .ZN(n4266) );
  NOR2_X1 U4673 ( .A1(n4266), .A2(n2509), .ZN(n3958) );
  AND2_X1 U4674 ( .A1(n4251), .A2(n3958), .ZN(n3959) );
  NAND4_X1 U4675 ( .A1(n3962), .A2(n3961), .A3(n3960), .A4(n3959), .ZN(n3963)
         );
  NOR2_X1 U4676 ( .A1(n3964), .A2(n3963), .ZN(n3967) );
  AND4_X1 U4677 ( .A1(n3967), .A2(n3970), .A3(n3966), .A4(n3965), .ZN(n3999)
         );
  INV_X1 U4678 ( .A(n3968), .ZN(n3998) );
  INV_X1 U4679 ( .A(n4012), .ZN(n3995) );
  NAND3_X1 U4680 ( .A1(n3971), .A2(n3970), .A3(n3969), .ZN(n3992) );
  INV_X1 U4681 ( .A(n3403), .ZN(n3974) );
  AOI21_X1 U4682 ( .B1(n3974), .B2(n3973), .A(n3972), .ZN(n3983) );
  INV_X1 U4683 ( .A(n3975), .ZN(n3980) );
  INV_X1 U4684 ( .A(n3976), .ZN(n3978) );
  OAI211_X1 U4685 ( .C1(n3980), .C2(n3979), .A(n3978), .B(n3977), .ZN(n3982)
         );
  OAI21_X1 U4686 ( .B1(n3983), .B2(n3982), .A(n3981), .ZN(n3986) );
  AOI21_X1 U4687 ( .B1(n3986), .B2(n3985), .A(n3984), .ZN(n3990) );
  NOR4_X1 U4688 ( .A1(n3990), .A2(n3989), .A3(n3988), .A4(n3987), .ZN(n3991)
         );
  AOI21_X1 U4689 ( .B1(n3993), .B2(n3992), .A(n3991), .ZN(n3994) );
  XNOR2_X1 U4690 ( .A(n4002), .B(n4316), .ZN(n4011) );
  INV_X1 U4691 ( .A(n4003), .ZN(n4008) );
  NAND2_X1 U4692 ( .A1(n4005), .A2(n4004), .ZN(n4006) );
  OAI211_X1 U4693 ( .C1(n4008), .C2(n4007), .A(B_REG_SCAN_IN), .B(n4006), .ZN(
        n4009) );
  OAI21_X1 U4694 ( .B1(n4011), .B2(n4010), .A(n4009), .ZN(U3239) );
  MUX2_X1 U4695 ( .A(n4012), .B(DATAO_REG_31__SCAN_IN), .S(n2808), .Z(U3581)
         );
  MUX2_X1 U4696 ( .A(n4013), .B(DATAO_REG_30__SCAN_IN), .S(n2808), .Z(U3580)
         );
  MUX2_X1 U4697 ( .A(n4014), .B(DATAO_REG_28__SCAN_IN), .S(n4025), .Z(U3578)
         );
  MUX2_X1 U4698 ( .A(n4015), .B(DATAO_REG_27__SCAN_IN), .S(n2808), .Z(U3577)
         );
  MUX2_X1 U4699 ( .A(n4383), .B(DATAO_REG_26__SCAN_IN), .S(n4025), .Z(U3576)
         );
  MUX2_X1 U4700 ( .A(DATAO_REG_24__SCAN_IN), .B(n4016), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4701 ( .A(n4211), .B(DATAO_REG_22__SCAN_IN), .S(n2808), .Z(U3572)
         );
  MUX2_X1 U4702 ( .A(DATAO_REG_21__SCAN_IN), .B(n4230), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4703 ( .A(n4411), .B(DATAO_REG_20__SCAN_IN), .S(n4025), .Z(U3570)
         );
  MUX2_X1 U4704 ( .A(n4421), .B(DATAO_REG_19__SCAN_IN), .S(n2808), .Z(U3569)
         );
  MUX2_X1 U4705 ( .A(n4289), .B(DATAO_REG_18__SCAN_IN), .S(n4025), .Z(U3568)
         );
  MUX2_X1 U4706 ( .A(n4447), .B(DATAO_REG_17__SCAN_IN), .S(n2808), .Z(U3567)
         );
  MUX2_X1 U4707 ( .A(n4456), .B(DATAO_REG_16__SCAN_IN), .S(n4025), .Z(U3566)
         );
  MUX2_X1 U4708 ( .A(n4467), .B(DATAO_REG_15__SCAN_IN), .S(n2808), .Z(U3565)
         );
  MUX2_X1 U4709 ( .A(n4455), .B(DATAO_REG_14__SCAN_IN), .S(n4025), .Z(U3564)
         );
  MUX2_X1 U4710 ( .A(n4487), .B(DATAO_REG_13__SCAN_IN), .S(n2808), .Z(U3563)
         );
  MUX2_X1 U4711 ( .A(n4017), .B(DATAO_REG_12__SCAN_IN), .S(n4025), .Z(U3562)
         );
  MUX2_X1 U4712 ( .A(n4484), .B(DATAO_REG_11__SCAN_IN), .S(n4025), .Z(U3561)
         );
  MUX2_X1 U4713 ( .A(n4018), .B(DATAO_REG_9__SCAN_IN), .S(n4025), .Z(U3559) );
  MUX2_X1 U4714 ( .A(n4019), .B(DATAO_REG_8__SCAN_IN), .S(n4025), .Z(U3558) );
  MUX2_X1 U4715 ( .A(n4020), .B(DATAO_REG_7__SCAN_IN), .S(n4025), .Z(U3557) );
  MUX2_X1 U4716 ( .A(n4021), .B(DATAO_REG_6__SCAN_IN), .S(n4025), .Z(U3556) );
  MUX2_X1 U4717 ( .A(n4022), .B(DATAO_REG_5__SCAN_IN), .S(n4025), .Z(U3555) );
  MUX2_X1 U4718 ( .A(n4023), .B(DATAO_REG_4__SCAN_IN), .S(n4025), .Z(U3554) );
  MUX2_X1 U4719 ( .A(n4024), .B(DATAO_REG_3__SCAN_IN), .S(n4025), .Z(U3553) );
  MUX2_X1 U4720 ( .A(n4026), .B(DATAO_REG_0__SCAN_IN), .S(n4025), .Z(U3550) );
  OAI211_X1 U4721 ( .C1(n2872), .C2(n4029), .A(n4110), .B(n4028), .ZN(n4036)
         );
  OAI211_X1 U4722 ( .C1(n4032), .C2(n4031), .A(n4730), .B(n4030), .ZN(n4035)
         );
  AOI22_X1 U4723 ( .A1(n4722), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4034) );
  NAND2_X1 U4724 ( .A1(n4065), .A2(n2870), .ZN(n4033) );
  NAND4_X1 U4725 ( .A1(n4036), .A2(n4035), .A3(n4034), .A4(n4033), .ZN(U3241)
         );
  XOR2_X1 U4726 ( .A(n4037), .B(REG2_REG_4__SCAN_IN), .Z(n4039) );
  AOI21_X1 U4727 ( .B1(n4110), .B2(n4039), .A(n4038), .ZN(n4046) );
  AOI21_X1 U4728 ( .B1(n4722), .B2(ADDR_REG_4__SCAN_IN), .A(n4040), .ZN(n4045)
         );
  OAI211_X1 U4729 ( .C1(n4042), .C2(REG1_REG_4__SCAN_IN), .A(n4730), .B(n4041), 
        .ZN(n4044) );
  NAND2_X1 U4730 ( .A1(n4065), .A2(n4695), .ZN(n4043) );
  NAND4_X1 U4731 ( .A1(n4046), .A2(n4045), .A3(n4044), .A4(n4043), .ZN(U3244)
         );
  NOR2_X1 U4732 ( .A1(n4735), .A2(n4047), .ZN(n4048) );
  AOI211_X1 U4733 ( .C1(n4722), .C2(ADDR_REG_5__SCAN_IN), .A(n4049), .B(n4048), 
        .ZN(n4058) );
  OAI211_X1 U4734 ( .C1(n4052), .C2(n4051), .A(n4730), .B(n4050), .ZN(n4057)
         );
  OAI211_X1 U4735 ( .C1(n4055), .C2(n4054), .A(n4110), .B(n4053), .ZN(n4056)
         );
  NAND3_X1 U4736 ( .A1(n4058), .A2(n4057), .A3(n4056), .ZN(U3245) );
  XNOR2_X1 U4737 ( .A(n4059), .B(REG1_REG_12__SCAN_IN), .ZN(n4068) );
  XOR2_X1 U4738 ( .A(REG2_REG_12__SCAN_IN), .B(n4060), .Z(n4061) );
  NAND2_X1 U4739 ( .A1(n4110), .A2(n4061), .ZN(n4063) );
  NAND2_X1 U4740 ( .A1(n4063), .A2(n4062), .ZN(n4064) );
  AOI21_X1 U4741 ( .B1(n4722), .B2(ADDR_REG_12__SCAN_IN), .A(n4064), .ZN(n4067) );
  NAND2_X1 U4742 ( .A1(n4065), .A2(n4690), .ZN(n4066) );
  OAI211_X1 U4743 ( .C1(n4068), .C2(n4114), .A(n4067), .B(n4066), .ZN(U3252)
         );
  XNOR2_X1 U4744 ( .A(n4075), .B(n3453), .ZN(n4069) );
  XNOR2_X1 U4745 ( .A(n4070), .B(n4069), .ZN(n4080) );
  AOI21_X1 U4746 ( .B1(n4072), .B2(n4071), .A(n4114), .ZN(n4074) );
  NAND2_X1 U4747 ( .A1(n4074), .A2(n4073), .ZN(n4079) );
  NOR2_X1 U4748 ( .A1(n4735), .A2(n4075), .ZN(n4076) );
  AOI211_X1 U4749 ( .C1(n4722), .C2(ADDR_REG_13__SCAN_IN), .A(n4077), .B(n4076), .ZN(n4078) );
  OAI211_X1 U4750 ( .C1(n4719), .C2(n4080), .A(n4079), .B(n4078), .ZN(U3253)
         );
  XNOR2_X1 U4751 ( .A(n4081), .B(REG1_REG_14__SCAN_IN), .ZN(n4091) );
  AOI21_X1 U4752 ( .B1(n4083), .B2(n4082), .A(n4719), .ZN(n4089) );
  NAND2_X1 U4753 ( .A1(n4722), .A2(ADDR_REG_14__SCAN_IN), .ZN(n4084) );
  OAI211_X1 U4754 ( .C1(n4735), .C2(n4086), .A(n4085), .B(n4084), .ZN(n4087)
         );
  AOI21_X1 U4755 ( .B1(n4089), .B2(n4088), .A(n4087), .ZN(n4090) );
  OAI21_X1 U4756 ( .B1(n4091), .B2(n4114), .A(n4090), .ZN(U3254) );
  AOI211_X1 U4757 ( .C1(n4093), .C2(n4092), .A(n4114), .B(n2041), .ZN(n4102)
         );
  OAI211_X1 U4758 ( .C1(n4096), .C2(n4095), .A(n4094), .B(n4110), .ZN(n4099)
         );
  AOI21_X1 U4759 ( .B1(n4722), .B2(ADDR_REG_15__SCAN_IN), .A(n4097), .ZN(n4098) );
  OAI211_X1 U4760 ( .C1(n4735), .C2(n4100), .A(n4099), .B(n4098), .ZN(n4101)
         );
  OR2_X1 U4761 ( .A1(n4102), .A2(n4101), .ZN(U3255) );
  INV_X1 U4762 ( .A(n4103), .ZN(n4105) );
  AOI21_X1 U4763 ( .B1(REG1_REG_16__SCAN_IN), .B2(n4105), .A(n4104), .ZN(n4115) );
  NOR2_X1 U4764 ( .A1(n4735), .A2(n4106), .ZN(n4107) );
  AOI211_X1 U4765 ( .C1(n4722), .C2(ADDR_REG_16__SCAN_IN), .A(n4108), .B(n4107), .ZN(n4113) );
  XNOR2_X1 U4766 ( .A(n4109), .B(n2505), .ZN(n4111) );
  NAND2_X1 U4767 ( .A1(n4111), .A2(n4110), .ZN(n4112) );
  OAI211_X1 U4768 ( .C1(n4115), .C2(n4114), .A(n4113), .B(n4112), .ZN(U3256)
         );
  NAND2_X1 U4769 ( .A1(n4437), .A2(n4120), .ZN(n4116) );
  AND2_X1 U4770 ( .A1(n4117), .A2(n4116), .ZN(n4501) );
  AOI21_X1 U4771 ( .B1(n4120), .B2(n4119), .A(n4118), .ZN(n4498) );
  NAND2_X1 U4772 ( .A1(n4498), .A2(n4741), .ZN(n4122) );
  NAND2_X1 U4773 ( .A1(n4745), .A2(REG2_REG_30__SCAN_IN), .ZN(n4121) );
  OAI211_X1 U4774 ( .C1(n4745), .C2(n4501), .A(n4122), .B(n4121), .ZN(U3261)
         );
  NAND2_X1 U4775 ( .A1(n4124), .A2(n4123), .ZN(n4126) );
  XNOR2_X1 U4776 ( .A(n4126), .B(n4125), .ZN(n4134) );
  INV_X1 U4777 ( .A(n4127), .ZN(n4131) );
  OAI22_X1 U4778 ( .A1(n4129), .A2(n4364), .B1(n4128), .B2(n4755), .ZN(n4130)
         );
  OAI21_X1 U4779 ( .B1(n4131), .B2(n4130), .A(n4752), .ZN(n4133) );
  NAND2_X1 U4780 ( .A1(n4745), .A2(REG2_REG_29__SCAN_IN), .ZN(n4132) );
  OAI211_X1 U4781 ( .C1(n4134), .C2(n4378), .A(n4133), .B(n4132), .ZN(U3354)
         );
  INV_X1 U4782 ( .A(n4135), .ZN(n4149) );
  INV_X1 U4783 ( .A(n4136), .ZN(n4147) );
  OAI22_X1 U4784 ( .A1(n4138), .A2(n4755), .B1(n4137), .B2(n4752), .ZN(n4142)
         );
  OAI22_X1 U4785 ( .A1(n4140), .A2(n4369), .B1(n4370), .B2(n4139), .ZN(n4141)
         );
  AOI211_X1 U4786 ( .C1(n4343), .C2(n4143), .A(n4142), .B(n4141), .ZN(n4144)
         );
  OAI21_X1 U4787 ( .B1(n4145), .B2(n4364), .A(n4144), .ZN(n4146) );
  OAI21_X1 U4788 ( .B1(n4149), .B2(n4378), .A(n4148), .ZN(U3262) );
  NAND2_X1 U4789 ( .A1(n4150), .A2(n4336), .ZN(n4160) );
  INV_X1 U4790 ( .A(n4151), .ZN(n4158) );
  AOI22_X1 U4791 ( .A1(n4152), .A2(n4737), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4745), .ZN(n4153) );
  OAI21_X1 U4792 ( .B1(n4183), .B2(n4369), .A(n4153), .ZN(n4157) );
  OAI22_X1 U4793 ( .A1(n4155), .A2(n4371), .B1(n4154), .B2(n4370), .ZN(n4156)
         );
  AOI211_X1 U4794 ( .C1(n4158), .C2(n4741), .A(n4157), .B(n4156), .ZN(n4159)
         );
  OAI211_X1 U4795 ( .C1(n4745), .C2(n4161), .A(n4160), .B(n4159), .ZN(U3263)
         );
  INV_X1 U4796 ( .A(n4162), .ZN(n4169) );
  AOI22_X1 U4797 ( .A1(n4163), .A2(n4737), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4745), .ZN(n4164) );
  OAI21_X1 U4798 ( .B1(n4165), .B2(n4364), .A(n4164), .ZN(n4166) );
  AOI21_X1 U4799 ( .B1(n4167), .B2(n4752), .A(n4166), .ZN(n4168) );
  OAI21_X1 U4800 ( .B1(n4169), .B2(n4378), .A(n4168), .ZN(U3264) );
  INV_X1 U4801 ( .A(n4170), .ZN(n4171) );
  XNOR2_X1 U4802 ( .A(n4173), .B(n4175), .ZN(n4174) );
  NAND2_X1 U4803 ( .A1(n4174), .A2(n4338), .ZN(n4385) );
  XNOR2_X1 U4804 ( .A(n4176), .B(n4175), .ZN(n4389) );
  NAND2_X1 U4805 ( .A1(n4389), .A2(n4336), .ZN(n4188) );
  INV_X1 U4806 ( .A(n4194), .ZN(n4179) );
  INV_X1 U4807 ( .A(n4177), .ZN(n4178) );
  INV_X1 U4808 ( .A(n4505), .ZN(n4186) );
  AOI22_X1 U4809 ( .A1(n4180), .A2(n4737), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4745), .ZN(n4181) );
  OAI21_X1 U4810 ( .B1(n4387), .B2(n4369), .A(n4181), .ZN(n4185) );
  OAI22_X1 U4811 ( .A1(n4183), .A2(n4371), .B1(n4370), .B2(n4182), .ZN(n4184)
         );
  AOI211_X1 U4812 ( .C1(n4186), .C2(n4741), .A(n4185), .B(n4184), .ZN(n4187)
         );
  OAI211_X1 U4813 ( .C1(n4745), .C2(n4385), .A(n4188), .B(n4187), .ZN(U3265)
         );
  XNOR2_X1 U4814 ( .A(n4189), .B(n4192), .ZN(n4190) );
  NAND2_X1 U4815 ( .A1(n4190), .A2(n4338), .ZN(n4395) );
  XOR2_X1 U4816 ( .A(n4192), .B(n4191), .Z(n4398) );
  NAND2_X1 U4817 ( .A1(n4398), .A2(n4336), .ZN(n4202) );
  NAND2_X1 U4818 ( .A1(n4214), .A2(n4392), .ZN(n4193) );
  NAND2_X1 U4819 ( .A1(n4194), .A2(n4193), .ZN(n4509) );
  INV_X1 U4820 ( .A(n4509), .ZN(n4200) );
  AOI22_X1 U4821 ( .A1(n4195), .A2(n4737), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4745), .ZN(n4196) );
  OAI21_X1 U4822 ( .B1(n4233), .B2(n4369), .A(n4196), .ZN(n4199) );
  OAI22_X1 U4823 ( .A1(n4396), .A2(n4371), .B1(n4197), .B2(n4370), .ZN(n4198)
         );
  AOI211_X1 U4824 ( .C1(n4200), .C2(n4741), .A(n4199), .B(n4198), .ZN(n4201)
         );
  OAI211_X1 U4825 ( .C1(n4745), .C2(n4395), .A(n4202), .B(n4201), .ZN(U3266)
         );
  XOR2_X1 U4826 ( .A(n4207), .B(n4203), .Z(n4402) );
  INV_X1 U4827 ( .A(n4402), .ZN(n4222) );
  NAND2_X1 U4828 ( .A1(n4248), .A2(n4204), .ZN(n4226) );
  AOI21_X1 U4829 ( .B1(n4226), .B2(n4223), .A(n2580), .ZN(n4228) );
  INV_X1 U4830 ( .A(n4205), .ZN(n4206) );
  NOR2_X1 U4831 ( .A1(n4228), .A2(n4206), .ZN(n4208) );
  XNOR2_X1 U4832 ( .A(n4208), .B(n4207), .ZN(n4209) );
  NAND2_X1 U4833 ( .A1(n4209), .A2(n4338), .ZN(n4213) );
  AOI22_X1 U4834 ( .A1(n4211), .A2(n4485), .B1(n4409), .B2(n4210), .ZN(n4212)
         );
  OAI211_X1 U4835 ( .C1(n4387), .C2(n4439), .A(n4213), .B(n4212), .ZN(n4401)
         );
  INV_X1 U4836 ( .A(n4240), .ZN(n4216) );
  OAI21_X1 U4837 ( .B1(n4216), .B2(n4215), .A(n4214), .ZN(n4513) );
  NOR2_X1 U4838 ( .A1(n4513), .A2(n4364), .ZN(n4220) );
  OAI22_X1 U4839 ( .A1(n4218), .A2(n4752), .B1(n4217), .B2(n4755), .ZN(n4219)
         );
  AOI211_X1 U4840 ( .C1(n4401), .C2(n4752), .A(n4220), .B(n4219), .ZN(n4221)
         );
  OAI21_X1 U4841 ( .B1(n4222), .B2(n4378), .A(n4221), .ZN(U3267) );
  INV_X1 U4842 ( .A(n4223), .ZN(n4224) );
  NOR2_X1 U4843 ( .A1(n4237), .A2(n4224), .ZN(n4225) );
  AND2_X1 U4844 ( .A1(n4226), .A2(n4225), .ZN(n4227) );
  OR2_X1 U4845 ( .A1(n4228), .A2(n4227), .ZN(n4235) );
  NAND2_X1 U4846 ( .A1(n4437), .A2(n4229), .ZN(n4232) );
  NAND2_X1 U4847 ( .A1(n4230), .A2(n4485), .ZN(n4231) );
  OAI211_X1 U4848 ( .C1(n4233), .C2(n4439), .A(n4232), .B(n4231), .ZN(n4234)
         );
  AOI21_X1 U4849 ( .B1(n4235), .B2(n4338), .A(n4234), .ZN(n4406) );
  NAND2_X1 U4850 ( .A1(n4238), .A2(n4237), .ZN(n4405) );
  NAND3_X1 U4851 ( .A1(n4236), .A2(n4405), .A3(n4336), .ZN(n4247) );
  OAI21_X1 U4852 ( .B1(n4239), .B2(n4241), .A(n4240), .ZN(n4517) );
  INV_X1 U4853 ( .A(n4517), .ZN(n4245) );
  INV_X1 U4854 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4243) );
  OAI22_X1 U4855 ( .A1(n4752), .A2(n4243), .B1(n4242), .B2(n4755), .ZN(n4244)
         );
  AOI21_X1 U4856 ( .B1(n4245), .B2(n4741), .A(n4244), .ZN(n4246) );
  OAI211_X1 U4857 ( .C1(n4745), .C2(n4406), .A(n4247), .B(n4246), .ZN(U3268)
         );
  XNOR2_X1 U4858 ( .A(n4248), .B(n4251), .ZN(n4249) );
  NAND2_X1 U4859 ( .A1(n4249), .A2(n4338), .ZN(n4413) );
  XNOR2_X1 U4860 ( .A(n4250), .B(n4251), .ZN(n4416) );
  NAND2_X1 U4861 ( .A1(n4416), .A2(n4336), .ZN(n4260) );
  INV_X1 U4862 ( .A(n4239), .ZN(n4252) );
  OAI21_X1 U4863 ( .B1(n4272), .B2(n4255), .A(n4252), .ZN(n4521) );
  INV_X1 U4864 ( .A(n4521), .ZN(n4258) );
  AOI22_X1 U4865 ( .A1(n4745), .A2(REG2_REG_21__SCAN_IN), .B1(n4253), .B2(
        n4737), .ZN(n4254) );
  OAI21_X1 U4866 ( .B1(n4369), .B2(n4292), .A(n4254), .ZN(n4257) );
  OAI22_X1 U4867 ( .A1(n4414), .A2(n4371), .B1(n4370), .B2(n4255), .ZN(n4256)
         );
  AOI211_X1 U4868 ( .C1(n4258), .C2(n4741), .A(n4257), .B(n4256), .ZN(n4259)
         );
  OAI211_X1 U4869 ( .C1(n4745), .C2(n4413), .A(n4260), .B(n4259), .ZN(U3269)
         );
  XNOR2_X1 U4870 ( .A(n4261), .B(n4266), .ZN(n4419) );
  INV_X1 U4871 ( .A(n4419), .ZN(n4280) );
  NAND2_X1 U4872 ( .A1(n4419), .A2(n4262), .ZN(n4271) );
  INV_X1 U4873 ( .A(n4263), .ZN(n4264) );
  NAND2_X1 U4874 ( .A1(n4265), .A2(n4264), .ZN(n4268) );
  INV_X1 U4875 ( .A(n4266), .ZN(n4267) );
  XNOR2_X1 U4876 ( .A(n4268), .B(n4267), .ZN(n4269) );
  NAND2_X1 U4877 ( .A1(n4269), .A2(n4338), .ZN(n4270) );
  NAND2_X1 U4878 ( .A1(n4271), .A2(n4270), .ZN(n4426) );
  NAND2_X1 U4879 ( .A1(n4426), .A2(n4752), .ZN(n4279) );
  AOI21_X1 U4880 ( .B1(n4420), .B2(n4295), .A(n4272), .ZN(n4524) );
  AOI22_X1 U4881 ( .A1(n4745), .A2(REG2_REG_20__SCAN_IN), .B1(n4273), .B2(
        n4737), .ZN(n4274) );
  OAI21_X1 U4882 ( .B1(n4369), .B2(n4313), .A(n4274), .ZN(n4277) );
  OAI22_X1 U4883 ( .A1(n4424), .A2(n4371), .B1(n4370), .B2(n4275), .ZN(n4276)
         );
  AOI211_X1 U4884 ( .C1(n4524), .C2(n4741), .A(n4277), .B(n4276), .ZN(n4278)
         );
  OAI211_X1 U4885 ( .C1(n4280), .C2(n4738), .A(n4279), .B(n4278), .ZN(U3270)
         );
  NAND2_X1 U4886 ( .A1(n4282), .A2(n4281), .ZN(n4310) );
  INV_X1 U4887 ( .A(n4283), .ZN(n4285) );
  OAI21_X1 U4888 ( .B1(n4310), .B2(n4285), .A(n4284), .ZN(n4286) );
  XNOR2_X1 U4889 ( .A(n4286), .B(n4294), .ZN(n4287) );
  NAND2_X1 U4890 ( .A1(n4287), .A2(n4338), .ZN(n4291) );
  AOI22_X1 U4891 ( .A1(n4289), .A2(n4485), .B1(n4409), .B2(n4288), .ZN(n4290)
         );
  OAI211_X1 U4892 ( .C1(n4292), .C2(n4439), .A(n4291), .B(n4290), .ZN(n4429)
         );
  INV_X1 U4893 ( .A(n4429), .ZN(n4302) );
  XNOR2_X1 U4894 ( .A(n4293), .B(n4294), .ZN(n4430) );
  INV_X1 U4895 ( .A(n4307), .ZN(n4297) );
  OAI21_X1 U4896 ( .B1(n4297), .B2(n4296), .A(n4295), .ZN(n4529) );
  AOI22_X1 U4897 ( .A1(n4745), .A2(REG2_REG_19__SCAN_IN), .B1(n4298), .B2(
        n4737), .ZN(n4299) );
  OAI21_X1 U4898 ( .B1(n4529), .B2(n4364), .A(n4299), .ZN(n4300) );
  AOI21_X1 U4899 ( .B1(n4430), .B2(n4336), .A(n4300), .ZN(n4301) );
  OAI21_X1 U4900 ( .B1(n4302), .B2(n4745), .A(n4301), .ZN(U3271) );
  OAI21_X1 U4901 ( .B1(n4305), .B2(n4304), .A(n4303), .ZN(n4306) );
  INV_X1 U4902 ( .A(n4306), .ZN(n4434) );
  OAI211_X1 U4903 ( .C1(n4328), .C2(n4308), .A(n4492), .B(n4307), .ZN(n4432)
         );
  XNOR2_X1 U4904 ( .A(n4310), .B(n4309), .ZN(n4315) );
  AOI22_X1 U4905 ( .A1(n4447), .A2(n4485), .B1(n4311), .B2(n4409), .ZN(n4312)
         );
  OAI21_X1 U4906 ( .B1(n4313), .B2(n4439), .A(n4312), .ZN(n4314) );
  AOI21_X1 U4907 ( .B1(n4315), .B2(n4338), .A(n4314), .ZN(n4433) );
  OAI21_X1 U4908 ( .B1(n4316), .B2(n4432), .A(n4433), .ZN(n4317) );
  NAND2_X1 U4909 ( .A1(n4317), .A2(n4752), .ZN(n4321) );
  INV_X1 U4910 ( .A(n4318), .ZN(n4319) );
  AOI22_X1 U4911 ( .A1(n4745), .A2(REG2_REG_18__SCAN_IN), .B1(n4319), .B2(
        n4737), .ZN(n4320) );
  OAI211_X1 U4912 ( .C1(n4434), .C2(n4378), .A(n4321), .B(n4320), .ZN(U3272)
         );
  XNOR2_X1 U4913 ( .A(n4322), .B(n4324), .ZN(n4323) );
  NAND2_X1 U4914 ( .A1(n4323), .A2(n4338), .ZN(n4442) );
  INV_X1 U4915 ( .A(n4324), .ZN(n4325) );
  XNOR2_X1 U4916 ( .A(n4326), .B(n4325), .ZN(n4435) );
  NOR2_X1 U4917 ( .A1(n4342), .A2(n4329), .ZN(n4327) );
  OR2_X1 U4918 ( .A1(n4328), .A2(n4327), .ZN(n4534) );
  OAI22_X1 U4919 ( .A1(n4440), .A2(n4371), .B1(n4370), .B2(n4329), .ZN(n4333)
         );
  AOI22_X1 U4920 ( .A1(n4745), .A2(REG2_REG_17__SCAN_IN), .B1(n4330), .B2(
        n4737), .ZN(n4331) );
  OAI21_X1 U4921 ( .B1(n4369), .B2(n4372), .A(n4331), .ZN(n4332) );
  NOR2_X1 U4922 ( .A1(n4333), .A2(n4332), .ZN(n4334) );
  OAI21_X1 U4923 ( .B1(n4534), .B2(n4364), .A(n4334), .ZN(n4335) );
  AOI21_X1 U4924 ( .B1(n4435), .B2(n4336), .A(n4335), .ZN(n4337) );
  OAI21_X1 U4925 ( .B1(n4745), .B2(n4442), .A(n4337), .ZN(U3273) );
  OAI211_X1 U4926 ( .C1(n4341), .C2(n4340), .A(n4339), .B(n4338), .ZN(n4452)
         );
  AOI21_X1 U4927 ( .B1(n4345), .B2(n4363), .A(n4342), .ZN(n4451) );
  AOI22_X1 U4928 ( .A1(n4345), .A2(n4344), .B1(n4343), .B2(n4447), .ZN(n4349)
         );
  INV_X1 U4929 ( .A(n4346), .ZN(n4347) );
  AOI22_X1 U4930 ( .A1(n4745), .A2(REG2_REG_16__SCAN_IN), .B1(n4347), .B2(
        n4737), .ZN(n4348) );
  OAI211_X1 U4931 ( .C1(n4350), .C2(n4369), .A(n4349), .B(n4348), .ZN(n4354)
         );
  OAI21_X1 U4932 ( .B1(n4352), .B2(n2509), .A(n4351), .ZN(n4454) );
  NOR2_X1 U4933 ( .A1(n4454), .A2(n4378), .ZN(n4353) );
  AOI211_X1 U4934 ( .C1(n4451), .C2(n4741), .A(n4354), .B(n4353), .ZN(n4355)
         );
  OAI21_X1 U4935 ( .B1(n4745), .B2(n4452), .A(n4355), .ZN(U3274) );
  XNOR2_X1 U4936 ( .A(n4356), .B(n4357), .ZN(n4461) );
  INV_X1 U4937 ( .A(n4461), .ZN(n4379) );
  AOI21_X1 U4938 ( .B1(n4358), .B2(n4357), .A(n4475), .ZN(n4360) );
  NAND2_X1 U4939 ( .A1(n4360), .A2(n4359), .ZN(n4458) );
  NOR2_X1 U4940 ( .A1(n4458), .A2(n4745), .ZN(n4376) );
  NAND2_X1 U4941 ( .A1(n3406), .A2(n4361), .ZN(n4362) );
  NAND2_X1 U4942 ( .A1(n4363), .A2(n4362), .ZN(n4539) );
  NOR2_X1 U4943 ( .A1(n4539), .A2(n4364), .ZN(n4375) );
  NOR2_X1 U4944 ( .A1(n4755), .A2(n4365), .ZN(n4366) );
  AOI21_X1 U4945 ( .B1(n4745), .B2(REG2_REG_15__SCAN_IN), .A(n4366), .ZN(n4367) );
  OAI21_X1 U4946 ( .B1(n4369), .B2(n4368), .A(n4367), .ZN(n4374) );
  OAI22_X1 U4947 ( .A1(n4372), .A2(n4371), .B1(n4370), .B2(n4459), .ZN(n4373)
         );
  NOR4_X1 U4948 ( .A1(n4376), .A2(n4375), .A3(n4374), .A4(n4373), .ZN(n4377)
         );
  OAI21_X1 U4949 ( .B1(n4379), .B2(n4378), .A(n4377), .ZN(U3275) );
  NAND2_X1 U4950 ( .A1(n4498), .A2(n2782), .ZN(n4381) );
  NAND2_X1 U4951 ( .A1(n4784), .A2(REG1_REG_30__SCAN_IN), .ZN(n4380) );
  OAI211_X1 U4952 ( .C1(n4501), .C2(n4784), .A(n4381), .B(n4380), .ZN(U3548)
         );
  INV_X1 U4953 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4390) );
  AOI22_X1 U4954 ( .A1(n4383), .A2(n4486), .B1(n4437), .B2(n4382), .ZN(n4384)
         );
  OAI211_X1 U4955 ( .C1(n4387), .C2(n4386), .A(n4385), .B(n4384), .ZN(n4388)
         );
  AOI21_X1 U4956 ( .B1(n4389), .B2(n4480), .A(n4388), .ZN(n4502) );
  MUX2_X1 U4957 ( .A(n4390), .B(n4502), .S(n4787), .Z(n4391) );
  OAI21_X1 U4958 ( .B1(n4483), .B2(n4505), .A(n4391), .ZN(U3543) );
  INV_X1 U4959 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4399) );
  AOI22_X1 U4960 ( .A1(n4393), .A2(n4485), .B1(n4437), .B2(n4392), .ZN(n4394)
         );
  OAI211_X1 U4961 ( .C1(n4396), .C2(n4439), .A(n4395), .B(n4394), .ZN(n4397)
         );
  AOI21_X1 U4962 ( .B1(n4398), .B2(n4480), .A(n4397), .ZN(n4506) );
  MUX2_X1 U4963 ( .A(n4399), .B(n4506), .S(n4787), .Z(n4400) );
  OAI21_X1 U4964 ( .B1(n4483), .B2(n4509), .A(n4400), .ZN(U3542) );
  INV_X1 U4965 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4403) );
  AOI21_X1 U4966 ( .B1(n4402), .B2(n4480), .A(n4401), .ZN(n4510) );
  MUX2_X1 U4967 ( .A(n4403), .B(n4510), .S(n4787), .Z(n4404) );
  OAI21_X1 U4968 ( .B1(n4483), .B2(n4513), .A(n4404), .ZN(U3541) );
  NAND3_X1 U4969 ( .A1(n4236), .A2(n4405), .A3(n4480), .ZN(n4407) );
  AND2_X1 U4970 ( .A1(n4407), .A2(n4406), .ZN(n4514) );
  MUX2_X1 U4971 ( .A(n4659), .B(n4514), .S(n4787), .Z(n4408) );
  OAI21_X1 U4972 ( .B1(n4483), .B2(n4517), .A(n4408), .ZN(U3540) );
  INV_X1 U4973 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4417) );
  AOI22_X1 U4974 ( .A1(n4411), .A2(n4485), .B1(n4410), .B2(n4409), .ZN(n4412)
         );
  OAI211_X1 U4975 ( .C1(n4414), .C2(n4439), .A(n4413), .B(n4412), .ZN(n4415)
         );
  AOI21_X1 U4976 ( .B1(n4416), .B2(n4480), .A(n4415), .ZN(n4518) );
  MUX2_X1 U4977 ( .A(n4417), .B(n4518), .S(n4787), .Z(n4418) );
  OAI21_X1 U4978 ( .B1(n4483), .B2(n4521), .A(n4418), .ZN(U3539) );
  NAND2_X1 U4979 ( .A1(n4419), .A2(n4776), .ZN(n4423) );
  AOI22_X1 U4980 ( .A1(n4421), .A2(n4485), .B1(n4420), .B2(n4437), .ZN(n4422)
         );
  OAI211_X1 U4981 ( .C1(n4424), .C2(n4439), .A(n4423), .B(n4422), .ZN(n4425)
         );
  OR2_X1 U4982 ( .A1(n4426), .A2(n4425), .ZN(n4522) );
  MUX2_X1 U4983 ( .A(REG1_REG_20__SCAN_IN), .B(n4522), .S(n4787), .Z(n4427) );
  AOI21_X1 U4984 ( .B1(n2782), .B2(n4524), .A(n4427), .ZN(n4428) );
  INV_X1 U4985 ( .A(n4428), .ZN(U3538) );
  AOI21_X1 U4986 ( .B1(n4480), .B2(n4430), .A(n4429), .ZN(n4526) );
  MUX2_X1 U4987 ( .A(n3476), .B(n4526), .S(n4787), .Z(n4431) );
  OAI21_X1 U4988 ( .B1(n4483), .B2(n4529), .A(n4431), .ZN(U3537) );
  OAI211_X1 U4989 ( .C1(n4434), .C2(n4497), .A(n4433), .B(n4432), .ZN(n4530)
         );
  MUX2_X1 U4990 ( .A(REG1_REG_18__SCAN_IN), .B(n4530), .S(n4787), .Z(U3536) );
  NAND2_X1 U4991 ( .A1(n4435), .A2(n4480), .ZN(n4444) );
  AOI22_X1 U4992 ( .A1(n4456), .A2(n4485), .B1(n4437), .B2(n4436), .ZN(n4438)
         );
  OAI21_X1 U4993 ( .B1(n4440), .B2(n4439), .A(n4438), .ZN(n4441) );
  INV_X1 U4994 ( .A(n4441), .ZN(n4443) );
  NAND3_X1 U4995 ( .A1(n4444), .A2(n4443), .A3(n4442), .ZN(n4531) );
  MUX2_X1 U4996 ( .A(n4531), .B(REG1_REG_17__SCAN_IN), .S(n4784), .Z(n4445) );
  INV_X1 U4997 ( .A(n4445), .ZN(n4446) );
  OAI21_X1 U4998 ( .B1(n4483), .B2(n4534), .A(n4446), .ZN(U3535) );
  AOI22_X1 U4999 ( .A1(n4447), .A2(n4486), .B1(n4485), .B2(n4467), .ZN(n4448)
         );
  OAI21_X1 U5000 ( .B1(n4449), .B2(n4489), .A(n4448), .ZN(n4450) );
  AOI21_X1 U5001 ( .B1(n4451), .B2(n4492), .A(n4450), .ZN(n4453) );
  OAI211_X1 U5002 ( .C1(n4454), .C2(n4497), .A(n4453), .B(n4452), .ZN(n4535)
         );
  MUX2_X1 U5003 ( .A(REG1_REG_16__SCAN_IN), .B(n4535), .S(n4787), .Z(U3534) );
  AOI22_X1 U5004 ( .A1(n4456), .A2(n4486), .B1(n4455), .B2(n4485), .ZN(n4457)
         );
  OAI211_X1 U5005 ( .C1(n4489), .C2(n4459), .A(n4458), .B(n4457), .ZN(n4460)
         );
  INV_X1 U5006 ( .A(n4460), .ZN(n4463) );
  NAND2_X1 U5007 ( .A1(n4461), .A2(n4480), .ZN(n4462) );
  NAND2_X1 U5008 ( .A1(n4463), .A2(n4462), .ZN(n4536) );
  MUX2_X1 U5009 ( .A(REG1_REG_15__SCAN_IN), .B(n4536), .S(n4787), .Z(n4464) );
  INV_X1 U5010 ( .A(n4464), .ZN(n4465) );
  OAI21_X1 U5011 ( .B1(n4483), .B2(n4539), .A(n4465), .ZN(U3533) );
  NAND2_X1 U5012 ( .A1(n4466), .A2(n4480), .ZN(n4473) );
  NAND2_X1 U5013 ( .A1(n4467), .A2(n4486), .ZN(n4469) );
  NAND2_X1 U5014 ( .A1(n4487), .A2(n4485), .ZN(n4468) );
  OAI211_X1 U5015 ( .C1(n4470), .C2(n4489), .A(n4469), .B(n4468), .ZN(n4471)
         );
  INV_X1 U5016 ( .A(n4471), .ZN(n4472) );
  OAI211_X1 U5017 ( .C1(n4475), .C2(n4474), .A(n4473), .B(n4472), .ZN(n4540)
         );
  MUX2_X1 U5018 ( .A(n4540), .B(REG1_REG_14__SCAN_IN), .S(n4784), .Z(n4476) );
  INV_X1 U5019 ( .A(n4476), .ZN(n4477) );
  OAI21_X1 U5020 ( .B1(n4483), .B2(n4543), .A(n4477), .ZN(U3532) );
  AOI21_X1 U5021 ( .B1(n4480), .B2(n4479), .A(n4478), .ZN(n4544) );
  MUX2_X1 U5022 ( .A(n4481), .B(n4544), .S(n4787), .Z(n4482) );
  OAI21_X1 U5023 ( .B1(n4483), .B2(n4547), .A(n4482), .ZN(U3531) );
  AOI22_X1 U5024 ( .A1(n4487), .A2(n4486), .B1(n4485), .B2(n4484), .ZN(n4488)
         );
  OAI21_X1 U5025 ( .B1(n4490), .B2(n4489), .A(n4488), .ZN(n4491) );
  AOI21_X1 U5026 ( .B1(n4493), .B2(n4492), .A(n4491), .ZN(n4494) );
  OAI211_X1 U5027 ( .C1(n4497), .C2(n4496), .A(n4495), .B(n4494), .ZN(n4548)
         );
  MUX2_X1 U5028 ( .A(REG1_REG_12__SCAN_IN), .B(n4548), .S(n4787), .Z(U3530) );
  NAND2_X1 U5029 ( .A1(n4498), .A2(n2788), .ZN(n4500) );
  NAND2_X1 U5030 ( .A1(n4782), .A2(REG0_REG_30__SCAN_IN), .ZN(n4499) );
  OAI211_X1 U5031 ( .C1(n4501), .C2(n4782), .A(n4500), .B(n4499), .ZN(U3516)
         );
  INV_X1 U5032 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4503) );
  MUX2_X1 U5033 ( .A(n4503), .B(n4502), .S(n4783), .Z(n4504) );
  OAI21_X1 U5034 ( .B1(n4505), .B2(n4546), .A(n4504), .ZN(U3511) );
  INV_X1 U5035 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4507) );
  MUX2_X1 U5036 ( .A(n4507), .B(n4506), .S(n4783), .Z(n4508) );
  OAI21_X1 U5037 ( .B1(n4509), .B2(n4546), .A(n4508), .ZN(U3510) );
  INV_X1 U5038 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4511) );
  MUX2_X1 U5039 ( .A(n4511), .B(n4510), .S(n4783), .Z(n4512) );
  OAI21_X1 U5040 ( .B1(n4513), .B2(n4546), .A(n4512), .ZN(U3509) );
  INV_X1 U5041 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4515) );
  MUX2_X1 U5042 ( .A(n4515), .B(n4514), .S(n4783), .Z(n4516) );
  OAI21_X1 U5043 ( .B1(n4517), .B2(n4546), .A(n4516), .ZN(U3508) );
  INV_X1 U5044 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4519) );
  MUX2_X1 U5045 ( .A(n4519), .B(n4518), .S(n4783), .Z(n4520) );
  OAI21_X1 U5046 ( .B1(n4521), .B2(n4546), .A(n4520), .ZN(U3507) );
  MUX2_X1 U5047 ( .A(REG0_REG_20__SCAN_IN), .B(n4522), .S(n4783), .Z(n4523) );
  AOI21_X1 U5048 ( .B1(n4524), .B2(n2788), .A(n4523), .ZN(n4525) );
  INV_X1 U5049 ( .A(n4525), .ZN(U3506) );
  INV_X1 U5050 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4527) );
  MUX2_X1 U5051 ( .A(n4527), .B(n4526), .S(n4783), .Z(n4528) );
  OAI21_X1 U5052 ( .B1(n4529), .B2(n4546), .A(n4528), .ZN(U3505) );
  MUX2_X1 U5053 ( .A(REG0_REG_18__SCAN_IN), .B(n4530), .S(n4783), .Z(U3503) );
  MUX2_X1 U5054 ( .A(n4531), .B(REG0_REG_17__SCAN_IN), .S(n4782), .Z(n4532) );
  INV_X1 U5055 ( .A(n4532), .ZN(n4533) );
  OAI21_X1 U5056 ( .B1(n4534), .B2(n4546), .A(n4533), .ZN(U3501) );
  MUX2_X1 U5057 ( .A(REG0_REG_16__SCAN_IN), .B(n4535), .S(n4783), .Z(U3499) );
  MUX2_X1 U5058 ( .A(REG0_REG_15__SCAN_IN), .B(n4536), .S(n4783), .Z(n4537) );
  INV_X1 U5059 ( .A(n4537), .ZN(n4538) );
  OAI21_X1 U5060 ( .B1(n4539), .B2(n4546), .A(n4538), .ZN(U3497) );
  MUX2_X1 U5061 ( .A(REG0_REG_14__SCAN_IN), .B(n4540), .S(n4783), .Z(n4541) );
  INV_X1 U5062 ( .A(n4541), .ZN(n4542) );
  OAI21_X1 U5063 ( .B1(n4543), .B2(n4546), .A(n4542), .ZN(U3495) );
  MUX2_X1 U5064 ( .A(n4624), .B(n4544), .S(n4783), .Z(n4545) );
  OAI21_X1 U5065 ( .B1(n4547), .B2(n4546), .A(n4545), .ZN(U3493) );
  MUX2_X1 U5066 ( .A(REG0_REG_12__SCAN_IN), .B(n4548), .S(n4783), .Z(n4685) );
  NOR3_X1 U5067 ( .A1(D_REG_1__SCAN_IN), .A2(DATAO_REG_25__SCAN_IN), .A3(n2178), .ZN(n4550) );
  NOR4_X1 U5068 ( .A1(IR_REG_22__SCAN_IN), .A2(REG1_REG_27__SCAN_IN), .A3(
        REG1_REG_15__SCAN_IN), .A4(REG1_REG_10__SCAN_IN), .ZN(n4549) );
  AND4_X1 U5069 ( .A1(n4551), .A2(REG2_REG_8__SCAN_IN), .A3(n4550), .A4(n4549), 
        .ZN(n4556) );
  NAND4_X1 U5070 ( .A1(IR_REG_16__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        REG2_REG_12__SCAN_IN), .A4(ADDR_REG_7__SCAN_IN), .ZN(n4554) );
  NAND4_X1 U5071 ( .A1(D_REG_4__SCAN_IN), .A2(REG0_REG_17__SCAN_IN), .A3(
        DATAI_9_), .A4(ADDR_REG_8__SCAN_IN), .ZN(n4553) );
  NAND3_X1 U5072 ( .A1(REG3_REG_23__SCAN_IN), .A2(REG1_REG_22__SCAN_IN), .A3(
        REG2_REG_13__SCAN_IN), .ZN(n4552) );
  NOR4_X1 U5073 ( .A1(REG1_REG_5__SCAN_IN), .A2(n4554), .A3(n4553), .A4(n4552), 
        .ZN(n4555) );
  AND2_X1 U5074 ( .A1(n4556), .A2(n4555), .ZN(n4644) );
  NOR4_X1 U5075 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG0_REG_21__SCAN_IN), .A3(
        REG0_REG_11__SCAN_IN), .A4(DATAO_REG_1__SCAN_IN), .ZN(n4559) );
  INV_X1 U5076 ( .A(IR_REG_20__SCAN_IN), .ZN(n4649) );
  NAND4_X1 U5077 ( .A1(REG3_REG_17__SCAN_IN), .A2(DATAI_23_), .A3(
        REG0_REG_4__SCAN_IN), .A4(n4649), .ZN(n4557) );
  NOR4_X1 U5078 ( .A1(DATAI_24_), .A2(DATAI_3_), .A3(n4647), .A4(n4557), .ZN(
        n4558) );
  NAND4_X1 U5079 ( .A1(IR_REG_29__SCAN_IN), .A2(n4559), .A3(n4558), .A4(n2467), 
        .ZN(n4572) );
  NAND4_X1 U5080 ( .A1(REG1_REG_26__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        REG0_REG_26__SCAN_IN), .A4(n3489), .ZN(n4571) );
  NAND4_X1 U5081 ( .A1(n4561), .A2(n4611), .A3(n4560), .A4(DATAI_21_), .ZN(
        n4565) );
  NAND4_X1 U5082 ( .A1(n4563), .A2(n4562), .A3(n2146), .A4(REG3_REG_9__SCAN_IN), .ZN(n4564) );
  NOR2_X1 U5083 ( .A1(n4565), .A2(n4564), .ZN(n4569) );
  NOR4_X1 U5084 ( .A1(IR_REG_9__SCAN_IN), .A2(REG2_REG_21__SCAN_IN), .A3(
        REG0_REG_13__SCAN_IN), .A4(DATAI_7_), .ZN(n4567) );
  AND4_X1 U5085 ( .A1(REG3_REG_14__SCAN_IN), .A2(REG3_REG_5__SCAN_IN), .A3(
        REG0_REG_20__SCAN_IN), .A4(DATAI_30_), .ZN(n4566) );
  AND4_X1 U5086 ( .A1(n2261), .A2(DATAO_REG_2__SCAN_IN), .A3(n4567), .A4(n4566), .ZN(n4568) );
  NAND4_X1 U5087 ( .A1(n4569), .A2(DATAO_REG_10__SCAN_IN), .A3(
        DATAO_REG_29__SCAN_IN), .A4(n4568), .ZN(n4570) );
  NOR3_X1 U5088 ( .A1(n4572), .A2(n4571), .A3(n4570), .ZN(n4643) );
  INV_X1 U5089 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n4574) );
  INV_X1 U5090 ( .A(D_REG_19__SCAN_IN), .ZN(n4758) );
  AOI22_X1 U5091 ( .A1(n4574), .A2(keyinput32), .B1(n4758), .B2(keyinput33), 
        .ZN(n4573) );
  OAI221_X1 U5092 ( .B1(n4574), .B2(keyinput32), .C1(n4758), .C2(keyinput33), 
        .A(n4573), .ZN(n4579) );
  AOI22_X1 U5093 ( .A1(n4577), .A2(keyinput53), .B1(n4576), .B2(keyinput50), 
        .ZN(n4575) );
  OAI221_X1 U5094 ( .B1(n4577), .B2(keyinput53), .C1(n4576), .C2(keyinput50), 
        .A(n4575), .ZN(n4578) );
  NOR2_X1 U5095 ( .A1(n4579), .A2(n4578), .ZN(n4606) );
  AOI22_X1 U5096 ( .A1(n2365), .A2(keyinput10), .B1(n2146), .B2(keyinput13), 
        .ZN(n4580) );
  OAI221_X1 U5097 ( .B1(n2365), .B2(keyinput10), .C1(n2146), .C2(keyinput13), 
        .A(n4580), .ZN(n4584) );
  AOI22_X1 U5098 ( .A1(n4561), .A2(keyinput6), .B1(n4582), .B2(keyinput4), 
        .ZN(n4581) );
  OAI221_X1 U5099 ( .B1(n4561), .B2(keyinput6), .C1(n4582), .C2(keyinput4), 
        .A(n4581), .ZN(n4583) );
  NOR2_X1 U5100 ( .A1(n4584), .A2(n4583), .ZN(n4605) );
  XNOR2_X1 U5101 ( .A(REG3_REG_9__SCAN_IN), .B(keyinput0), .ZN(n4588) );
  XNOR2_X1 U5102 ( .A(IR_REG_18__SCAN_IN), .B(keyinput5), .ZN(n4587) );
  XNOR2_X1 U5103 ( .A(REG1_REG_26__SCAN_IN), .B(keyinput1), .ZN(n4586) );
  XNOR2_X1 U5104 ( .A(IR_REG_9__SCAN_IN), .B(keyinput34), .ZN(n4585) );
  NAND4_X1 U5105 ( .A1(n4588), .A2(n4587), .A3(n4586), .A4(n4585), .ZN(n4594)
         );
  XNOR2_X1 U5106 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput12), .ZN(n4592) );
  XNOR2_X1 U5107 ( .A(IR_REG_16__SCAN_IN), .B(keyinput41), .ZN(n4591) );
  XNOR2_X1 U5108 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput42), .ZN(n4590) );
  XNOR2_X1 U5109 ( .A(IR_REG_5__SCAN_IN), .B(keyinput45), .ZN(n4589) );
  NAND4_X1 U5110 ( .A1(n4592), .A2(n4591), .A3(n4590), .A4(n4589), .ZN(n4593)
         );
  NOR2_X1 U5111 ( .A1(n4594), .A2(n4593), .ZN(n4604) );
  INV_X1 U5112 ( .A(DATAI_24_), .ZN(n4596) );
  AOI22_X1 U5113 ( .A1(n2467), .A2(keyinput49), .B1(keyinput48), .B2(n4596), 
        .ZN(n4595) );
  OAI221_X1 U5114 ( .B1(n2467), .B2(keyinput49), .C1(n4596), .C2(keyinput48), 
        .A(n4595), .ZN(n4602) );
  XNOR2_X1 U5115 ( .A(keyinput40), .B(REG2_REG_12__SCAN_IN), .ZN(n4600) );
  XNOR2_X1 U5116 ( .A(IR_REG_22__SCAN_IN), .B(keyinput44), .ZN(n4599) );
  XNOR2_X1 U5117 ( .A(keyinput46), .B(DATAI_21_), .ZN(n4598) );
  XNOR2_X1 U5118 ( .A(keyinput37), .B(REG2_REG_21__SCAN_IN), .ZN(n4597) );
  NAND4_X1 U5119 ( .A1(n4600), .A2(n4599), .A3(n4598), .A4(n4597), .ZN(n4601)
         );
  NOR2_X1 U5120 ( .A1(n4602), .A2(n4601), .ZN(n4603) );
  AND4_X1 U5121 ( .A1(n4606), .A2(n4605), .A3(n4604), .A4(n4603), .ZN(n4631)
         );
  INV_X1 U5122 ( .A(DATAI_30_), .ZN(n4609) );
  AOI22_X1 U5123 ( .A1(n4609), .A2(keyinput8), .B1(n4608), .B2(keyinput9), 
        .ZN(n4607) );
  OAI221_X1 U5124 ( .B1(n4609), .B2(keyinput8), .C1(n4608), .C2(keyinput9), 
        .A(n4607), .ZN(n4610) );
  INV_X1 U5125 ( .A(n4610), .ZN(n4616) );
  XNOR2_X1 U5126 ( .A(keyinput2), .B(n4611), .ZN(n4614) );
  XNOR2_X1 U5127 ( .A(keyinput14), .B(n4612), .ZN(n4613) );
  NOR2_X1 U5128 ( .A1(n4614), .A2(n4613), .ZN(n4615) );
  NAND2_X1 U5129 ( .A1(n4616), .A2(n4615), .ZN(n4621) );
  INV_X1 U5130 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n4619) );
  INV_X1 U5131 ( .A(DATAI_9_), .ZN(n4618) );
  AOI22_X1 U5132 ( .A1(n4619), .A2(keyinput36), .B1(n4618), .B2(keyinput38), 
        .ZN(n4617) );
  OAI221_X1 U5133 ( .B1(n4619), .B2(keyinput36), .C1(n4618), .C2(keyinput38), 
        .A(n4617), .ZN(n4620) );
  NOR2_X1 U5134 ( .A1(n4621), .A2(n4620), .ZN(n4630) );
  INV_X1 U5135 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4624) );
  INV_X1 U5136 ( .A(DATAI_7_), .ZN(n4623) );
  AOI22_X1 U5137 ( .A1(n4624), .A2(keyinput18), .B1(keyinput21), .B2(n4623), 
        .ZN(n4622) );
  OAI221_X1 U5138 ( .B1(n4624), .B2(keyinput18), .C1(n4623), .C2(keyinput21), 
        .A(n4622), .ZN(n4628) );
  AOI22_X1 U5139 ( .A1(n4757), .A2(keyinput17), .B1(keyinput16), .B2(n4626), 
        .ZN(n4625) );
  OAI221_X1 U5140 ( .B1(n4757), .B2(keyinput17), .C1(n4626), .C2(keyinput16), 
        .A(n4625), .ZN(n4627) );
  NOR2_X1 U5141 ( .A1(n4628), .A2(n4627), .ZN(n4629) );
  NAND3_X1 U5142 ( .A1(n4631), .A2(n4630), .A3(n4629), .ZN(n4642) );
  AOI22_X1 U5143 ( .A1(n4736), .A2(keyinput7), .B1(keyinput3), .B2(n4519), 
        .ZN(n4632) );
  OAI221_X1 U5144 ( .B1(n4736), .B2(keyinput7), .C1(n4519), .C2(keyinput3), 
        .A(n4632), .ZN(n4640) );
  AOI22_X1 U5145 ( .A1(n3489), .A2(keyinput15), .B1(n4634), .B2(keyinput31), 
        .ZN(n4633) );
  OAI221_X1 U5146 ( .B1(n3489), .B2(keyinput15), .C1(n4634), .C2(keyinput31), 
        .A(n4633), .ZN(n4639) );
  INV_X1 U5147 ( .A(D_REG_5__SCAN_IN), .ZN(n4764) );
  INV_X1 U5148 ( .A(D_REG_27__SCAN_IN), .ZN(n4756) );
  AOI22_X1 U5149 ( .A1(n4764), .A2(keyinput63), .B1(keyinput39), .B2(n4756), 
        .ZN(n4635) );
  OAI221_X1 U5150 ( .B1(n4764), .B2(keyinput63), .C1(n4756), .C2(keyinput39), 
        .A(n4635), .ZN(n4638) );
  INV_X1 U5151 ( .A(D_REG_10__SCAN_IN), .ZN(n4761) );
  AOI22_X1 U5152 ( .A1(n4761), .A2(keyinput35), .B1(n4760), .B2(keyinput11), 
        .ZN(n4636) );
  OAI221_X1 U5153 ( .B1(n4761), .B2(keyinput35), .C1(n4760), .C2(keyinput11), 
        .A(n4636), .ZN(n4637) );
  OR4_X1 U5154 ( .A1(n4640), .A2(n4639), .A3(n4638), .A4(n4637), .ZN(n4641) );
  AOI211_X1 U5155 ( .C1(n4644), .C2(n4643), .A(n4642), .B(n4641), .ZN(n4683)
         );
  INV_X1 U5156 ( .A(DATAI_3_), .ZN(n4646) );
  AOI22_X1 U5157 ( .A1(n4647), .A2(keyinput59), .B1(keyinput51), .B2(n4646), 
        .ZN(n4645) );
  OAI221_X1 U5158 ( .B1(n4647), .B2(keyinput59), .C1(n4646), .C2(keyinput51), 
        .A(n4645), .ZN(n4657) );
  INV_X1 U5159 ( .A(DATAI_23_), .ZN(n4769) );
  AOI22_X1 U5160 ( .A1(n4649), .A2(keyinput43), .B1(keyinput55), .B2(n4769), 
        .ZN(n4648) );
  OAI221_X1 U5161 ( .B1(n4649), .B2(keyinput43), .C1(n4769), .C2(keyinput55), 
        .A(n4648), .ZN(n4656) );
  AOI22_X1 U5162 ( .A1(n4651), .A2(keyinput47), .B1(keyinput27), .B2(n2352), 
        .ZN(n4650) );
  OAI221_X1 U5163 ( .B1(n4651), .B2(keyinput47), .C1(n2352), .C2(keyinput27), 
        .A(n4650), .ZN(n4655) );
  AOI22_X1 U5164 ( .A1(n3438), .A2(keyinput19), .B1(keyinput23), .B2(n4653), 
        .ZN(n4652) );
  OAI221_X1 U5165 ( .B1(n3438), .B2(keyinput19), .C1(n4653), .C2(keyinput23), 
        .A(n4652), .ZN(n4654) );
  NOR4_X1 U5166 ( .A1(n4657), .A2(n4656), .A3(n4655), .A4(n4654), .ZN(n4682)
         );
  AOI22_X1 U5167 ( .A1(n4659), .A2(keyinput20), .B1(n4763), .B2(keyinput22), 
        .ZN(n4658) );
  OAI221_X1 U5168 ( .B1(n4659), .B2(keyinput20), .C1(n4763), .C2(keyinput22), 
        .A(n4658), .ZN(n4668) );
  INV_X1 U5169 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4661) );
  INV_X1 U5170 ( .A(D_REG_4__SCAN_IN), .ZN(n4765) );
  AOI22_X1 U5171 ( .A1(n4661), .A2(keyinput25), .B1(n4765), .B2(keyinput24), 
        .ZN(n4660) );
  OAI221_X1 U5172 ( .B1(n4661), .B2(keyinput25), .C1(n4765), .C2(keyinput24), 
        .A(n4660), .ZN(n4667) );
  INV_X1 U5173 ( .A(D_REG_12__SCAN_IN), .ZN(n4759) );
  AOI22_X1 U5174 ( .A1(n4663), .A2(keyinput26), .B1(n4759), .B2(keyinput29), 
        .ZN(n4662) );
  OAI221_X1 U5175 ( .B1(n4663), .B2(keyinput26), .C1(n4759), .C2(keyinput29), 
        .A(n4662), .ZN(n4666) );
  AOI22_X1 U5176 ( .A1(n2904), .A2(keyinput30), .B1(n4762), .B2(keyinput28), 
        .ZN(n4664) );
  OAI221_X1 U5177 ( .B1(n2904), .B2(keyinput30), .C1(n4762), .C2(keyinput28), 
        .A(n4664), .ZN(n4665) );
  NOR4_X1 U5178 ( .A1(n4668), .A2(n4667), .A3(n4666), .A4(n4665), .ZN(n4681)
         );
  AOI22_X1 U5179 ( .A1(n2178), .A2(keyinput54), .B1(n2819), .B2(keyinput52), 
        .ZN(n4669) );
  OAI221_X1 U5180 ( .B1(n2178), .B2(keyinput54), .C1(n2819), .C2(keyinput52), 
        .A(n4669), .ZN(n4679) );
  AOI22_X1 U5181 ( .A1(n3453), .A2(keyinput56), .B1(keyinput57), .B2(n4671), 
        .ZN(n4670) );
  OAI221_X1 U5182 ( .B1(n3453), .B2(keyinput56), .C1(n4671), .C2(keyinput57), 
        .A(n4670), .ZN(n4678) );
  AOI22_X1 U5183 ( .A1(n2799), .A2(keyinput61), .B1(keyinput58), .B2(n4673), 
        .ZN(n4672) );
  OAI221_X1 U5184 ( .B1(n2799), .B2(keyinput61), .C1(n4673), .C2(keyinput58), 
        .A(n4672), .ZN(n4677) );
  AOI22_X1 U5185 ( .A1(n3105), .A2(keyinput60), .B1(n4675), .B2(keyinput62), 
        .ZN(n4674) );
  OAI221_X1 U5186 ( .B1(n3105), .B2(keyinput60), .C1(n4675), .C2(keyinput62), 
        .A(n4674), .ZN(n4676) );
  NOR4_X1 U5187 ( .A1(n4679), .A2(n4678), .A3(n4677), .A4(n4676), .ZN(n4680)
         );
  NAND4_X1 U5188 ( .A1(n4683), .A2(n4682), .A3(n4681), .A4(n4680), .ZN(n4684)
         );
  XNOR2_X1 U5189 ( .A(n4685), .B(n4684), .ZN(U3491) );
  MUX2_X1 U5190 ( .A(DATAI_30_), .B(n4686), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U5191 ( .A(n4705), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U5192 ( .A(DATAI_24_), .B(n2707), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U5193 ( .A(DATAI_21_), .B(n4687), .S(STATE_REG_SCAN_IN), .Z(U3331)
         );
  MUX2_X1 U5194 ( .A(n4688), .B(DATAI_16_), .S(U3149), .Z(U3336) );
  MUX2_X1 U5195 ( .A(n4689), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U5196 ( .A(n4690), .B(DATAI_12_), .S(U3149), .Z(U3340) );
  MUX2_X1 U5197 ( .A(n4691), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5198 ( .A(DATAI_9_), .B(n4692), .S(STATE_REG_SCAN_IN), .Z(U3343) );
  MUX2_X1 U5199 ( .A(DATAI_8_), .B(n2199), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5200 ( .A(n4693), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U5201 ( .A(n4694), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5202 ( .A(DATAI_4_), .B(n4695), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5203 ( .A(DATAI_3_), .B(n4696), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5204 ( .A(n4697), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5205 ( .A(n2870), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U5206 ( .A(DATAI_28_), .ZN(n4698) );
  AOI22_X1 U5207 ( .A1(STATE_REG_SCAN_IN), .A2(n4699), .B1(n4698), .B2(U3149), 
        .ZN(U3324) );
  INV_X1 U5208 ( .A(n4700), .ZN(n4704) );
  OAI21_X1 U5209 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4705), .A(n4702), .ZN(n4701)
         );
  MUX2_X1 U5210 ( .A(n4702), .B(n4701), .S(IR_REG_0__SCAN_IN), .Z(n4703) );
  OAI21_X1 U5211 ( .B1(n4705), .B2(n4704), .A(n4703), .ZN(n4707) );
  AOI22_X1 U5212 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4722), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4706) );
  OAI21_X1 U5213 ( .B1(n4708), .B2(n4707), .A(n4706), .ZN(U3240) );
  AOI211_X1 U5214 ( .C1(n4722), .C2(ADDR_REG_17__SCAN_IN), .A(n4713), .B(n4712), .ZN(n4717) );
  OAI221_X1 U5215 ( .B1(n2018), .B2(n4715), .C1(n2018), .C2(n4714), .A(n4730), 
        .ZN(n4716) );
  OAI211_X1 U5216 ( .C1(n4735), .C2(n4773), .A(n4717), .B(n4716), .ZN(U3257)
         );
  AOI21_X1 U5217 ( .B1(n4721), .B2(n4720), .A(n4719), .ZN(n4727) );
  NAND2_X1 U5218 ( .A1(n4722), .A2(ADDR_REG_18__SCAN_IN), .ZN(n4725) );
  INV_X1 U5219 ( .A(n4723), .ZN(n4724) );
  NAND2_X1 U5220 ( .A1(n4725), .A2(n4724), .ZN(n4726) );
  OAI211_X1 U5221 ( .C1(n4732), .C2(n4731), .A(n4730), .B(n4729), .ZN(n4733)
         );
  OAI211_X1 U5222 ( .C1(n4735), .C2(n4771), .A(n4734), .B(n4733), .ZN(U3258)
         );
  AOI22_X1 U5223 ( .A1(n4745), .A2(REG2_REG_3__SCAN_IN), .B1(n4737), .B2(n4736), .ZN(n4743) );
  INV_X1 U5224 ( .A(n4738), .ZN(n4747) );
  AOI22_X1 U5225 ( .A1(n4741), .A2(n4740), .B1(n4747), .B2(n4739), .ZN(n4742)
         );
  OAI211_X1 U5226 ( .C1(n4745), .C2(n4744), .A(n4743), .B(n4742), .ZN(U3287)
         );
  AOI22_X1 U5227 ( .A1(n4747), .A2(n4746), .B1(REG2_REG_0__SCAN_IN), .B2(n4745), .ZN(n4754) );
  OAI21_X1 U5228 ( .B1(n4750), .B2(n4749), .A(n4748), .ZN(n4751) );
  NAND2_X1 U5229 ( .A1(n4752), .A2(n4751), .ZN(n4753) );
  OAI211_X1 U5230 ( .C1(n4755), .C2(n2999), .A(n4754), .B(n4753), .ZN(U3290)
         );
  AND2_X1 U5231 ( .A1(D_REG_31__SCAN_IN), .A2(n4767), .ZN(U3291) );
  AND2_X1 U5232 ( .A1(D_REG_30__SCAN_IN), .A2(n4767), .ZN(U3292) );
  AND2_X1 U5233 ( .A1(D_REG_29__SCAN_IN), .A2(n4767), .ZN(U3293) );
  AND2_X1 U5234 ( .A1(D_REG_28__SCAN_IN), .A2(n4767), .ZN(U3294) );
  NOR2_X1 U5235 ( .A1(n4766), .A2(n4756), .ZN(U3295) );
  AND2_X1 U5236 ( .A1(D_REG_26__SCAN_IN), .A2(n4767), .ZN(U3296) );
  AND2_X1 U5237 ( .A1(D_REG_25__SCAN_IN), .A2(n4767), .ZN(U3297) );
  AND2_X1 U5238 ( .A1(D_REG_24__SCAN_IN), .A2(n4767), .ZN(U3298) );
  AND2_X1 U5239 ( .A1(D_REG_23__SCAN_IN), .A2(n4767), .ZN(U3299) );
  NOR2_X1 U5240 ( .A1(n4766), .A2(n4757), .ZN(U3300) );
  AND2_X1 U5241 ( .A1(D_REG_21__SCAN_IN), .A2(n4767), .ZN(U3301) );
  AND2_X1 U5242 ( .A1(D_REG_20__SCAN_IN), .A2(n4767), .ZN(U3302) );
  NOR2_X1 U5243 ( .A1(n4766), .A2(n4758), .ZN(U3303) );
  AND2_X1 U5244 ( .A1(D_REG_18__SCAN_IN), .A2(n4767), .ZN(U3304) );
  AND2_X1 U5245 ( .A1(D_REG_17__SCAN_IN), .A2(n4767), .ZN(U3305) );
  AND2_X1 U5246 ( .A1(D_REG_16__SCAN_IN), .A2(n4767), .ZN(U3306) );
  AND2_X1 U5247 ( .A1(D_REG_15__SCAN_IN), .A2(n4767), .ZN(U3307) );
  AND2_X1 U5248 ( .A1(D_REG_14__SCAN_IN), .A2(n4767), .ZN(U3308) );
  AND2_X1 U5249 ( .A1(D_REG_13__SCAN_IN), .A2(n4767), .ZN(U3309) );
  NOR2_X1 U5250 ( .A1(n4766), .A2(n4759), .ZN(U3310) );
  NOR2_X1 U5251 ( .A1(n4766), .A2(n4760), .ZN(U3311) );
  NOR2_X1 U5252 ( .A1(n4766), .A2(n4761), .ZN(U3312) );
  NOR2_X1 U5253 ( .A1(n4766), .A2(n4762), .ZN(U3313) );
  AND2_X1 U5254 ( .A1(D_REG_8__SCAN_IN), .A2(n4767), .ZN(U3314) );
  AND2_X1 U5255 ( .A1(D_REG_7__SCAN_IN), .A2(n4767), .ZN(U3315) );
  NOR2_X1 U5256 ( .A1(n4766), .A2(n4763), .ZN(U3316) );
  NOR2_X1 U5257 ( .A1(n4766), .A2(n4764), .ZN(U3317) );
  NOR2_X1 U5258 ( .A1(n4766), .A2(n4765), .ZN(U3318) );
  AND2_X1 U5259 ( .A1(D_REG_3__SCAN_IN), .A2(n4767), .ZN(U3319) );
  AND2_X1 U5260 ( .A1(D_REG_2__SCAN_IN), .A2(n4767), .ZN(U3320) );
  AOI21_X1 U5261 ( .B1(U3149), .B2(n4769), .A(n4768), .ZN(U3329) );
  INV_X1 U5262 ( .A(DATAI_18_), .ZN(n4770) );
  AOI22_X1 U5263 ( .A1(STATE_REG_SCAN_IN), .A2(n4771), .B1(n4770), .B2(U3149), 
        .ZN(U3334) );
  INV_X1 U5264 ( .A(DATAI_17_), .ZN(n4772) );
  AOI22_X1 U5265 ( .A1(STATE_REG_SCAN_IN), .A2(n4773), .B1(n4772), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5266 ( .A(DATAI_0_), .ZN(n4774) );
  AOI22_X1 U5267 ( .A1(STATE_REG_SCAN_IN), .A2(n2231), .B1(n4774), .B2(U3149), 
        .ZN(U3352) );
  AOI22_X1 U5268 ( .A1(n4783), .A2(n4775), .B1(n2335), .B2(n4782), .ZN(U3467)
         );
  AND2_X1 U5269 ( .A1(n4777), .A2(n4776), .ZN(n4780) );
  INV_X1 U5270 ( .A(n4778), .ZN(n4779) );
  NOR3_X1 U5271 ( .A1(n4781), .A2(n4780), .A3(n4779), .ZN(n4786) );
  AOI22_X1 U5272 ( .A1(n4783), .A2(n4786), .B1(n2352), .B2(n4782), .ZN(U3475)
         );
  INV_X1 U5273 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4785) );
  AOI22_X1 U5274 ( .A1(n4787), .A2(n4786), .B1(n4785), .B2(n4784), .ZN(U3522)
         );
endmodule

