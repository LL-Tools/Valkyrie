

module b20_C_gen_AntiSAT_k_128_7 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, 
        ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, 
        ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, 
        ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, 
        ADD_1068_U5, ADD_1068_U46, U126, U123, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3439, P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, 
        P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, 
        P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, 
        P1_U3501, P1_U3504, P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, 
        P1_U3513, P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, 
        P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, 
        P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, 
        P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, 
        P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, 
        P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, 
        P1_U3559, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, 
        P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, 
        P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, 
        P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, 
        P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, 
        P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, 
        P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, 
        P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, 
        P2_U3264, P2_U3376, P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, 
        P2_U3396, P2_U3399, P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, 
        P2_U3417, P2_U3420, P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, 
        P2_U3438, P2_U3441, P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, 
        P2_U3450, P2_U3451, P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, 
        P2_U3457, P2_U3458, P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, 
        P2_U3464, P2_U3465, P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, 
        P2_U3471, P2_U3472, P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, 
        P2_U3478, P2_U3479, P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, 
        P2_U3485, P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, 
        P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, 
        P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, 
        P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, 
        P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, 
        P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, 
        P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, 
        P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, 
        P2_U3183, P2_U3182, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, 
        P2_U3496, P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, 
        P2_U3503, P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, 
        P2_U3510, P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, 
        P2_U3517, P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, 
        P2_U3181, P2_U3180, P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, 
        P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, 
        P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, 
        P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, 
        P2_U3153, P2_U3151, P2_U3150, P2_U3893 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254;

  OAI21_X1 U4856 ( .B1(n8609), .B2(n8400), .A(n6259), .ZN(n8587) );
  NAND2_X1 U4857 ( .A1(n8193), .A2(n8192), .ZN(n8345) );
  CLKBUF_X2 U4858 ( .A(n5194), .Z(n7596) );
  INV_X1 U4859 ( .A(n5194), .ZN(n5602) );
  INV_X1 U4860 ( .A(n6491), .ZN(n5725) );
  BUF_X1 U4861 ( .A(n6809), .Z(n4449) );
  NAND3_X1 U4863 ( .A1(n5837), .A2(n5836), .A3(n5835), .ZN(n5884) );
  CLKBUF_X1 U4864 ( .A(n8696), .Z(n4350) );
  NOR2_X1 U4865 ( .A1(n6831), .A2(n8708), .ZN(n8696) );
  NAND2_X2 U4866 ( .A1(n5155), .A2(n5752), .ZN(n5361) );
  INV_X1 U4867 ( .A(n6370), .ZN(n7962) );
  INV_X1 U4868 ( .A(n6139), .ZN(n5903) );
  NAND2_X1 U4869 ( .A1(n4471), .A2(n4423), .ZN(n8676) );
  AOI22_X1 U4870 ( .A1(n8702), .A2(n6249), .B1(n8709), .B2(n8173), .ZN(n8690)
         );
  CLKBUF_X2 U4871 ( .A(n5775), .Z(n6341) );
  INV_X1 U4872 ( .A(n6491), .ZN(n6493) );
  NAND2_X1 U4873 ( .A1(n5806), .A2(n7801), .ZN(n6702) );
  OR2_X1 U4874 ( .A1(n6137), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6145) );
  INV_X1 U4875 ( .A(n6474), .ZN(n5601) );
  AND2_X1 U4876 ( .A1(n5115), .A2(n5114), .ZN(n5239) );
  INV_X2 U4877 ( .A(n6139), .ZN(n7003) );
  INV_X1 U4878 ( .A(n8259), .ZN(n8843) );
  INV_X2 U4879 ( .A(n6452), .ZN(n4611) );
  NAND2_X1 U4880 ( .A1(n5290), .A2(n5289), .ZN(n6783) );
  BUF_X1 U4881 ( .A(n6798), .Z(n4354) );
  NAND2_X1 U4882 ( .A1(n4675), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4674) );
  NAND4_X1 U4883 ( .A1(n5266), .A2(n5265), .A3(n5264), .A4(n5263), .ZN(n9040)
         );
  AND2_X1 U4884 ( .A1(n4809), .A2(n4427), .ZN(n4351) );
  NAND2_X2 U4885 ( .A1(n7330), .A2(n7329), .ZN(n7332) );
  OAI21_X2 U4886 ( .B1(n9251), .B2(n7862), .A(n7863), .ZN(n9235) );
  NAND2_X2 U4887 ( .A1(n7861), .A2(n7860), .ZN(n9251) );
  INV_X1 U4888 ( .A(n6274), .ZN(n8389) );
  OAI22_X2 U4889 ( .A1(n5460), .A2(n5048), .B1(SI_13_), .B2(n5458), .ZN(n5484)
         );
  OAI21_X2 U4890 ( .B1(n5430), .B2(n5046), .A(n5045), .ZN(n5460) );
  OAI22_X2 U4891 ( .A1(n9309), .A2(n7854), .B1(n9453), .B2(n9440), .ZN(n9291)
         );
  OAI21_X2 U4892 ( .B1(n9325), .B2(n7852), .A(n7853), .ZN(n9309) );
  OAI22_X2 U4893 ( .A1(n8587), .A2(n6260), .B1(n8605), .B2(n8796), .ZN(n8577)
         );
  OR2_X1 U4894 ( .A1(n7975), .A2(n9627), .ZN(n4809) );
  INV_X1 U4895 ( .A(n8549), .ZN(n8543) );
  NAND2_X1 U4896 ( .A1(n7074), .A2(n7072), .ZN(n6927) );
  OAI21_X1 U4897 ( .B1(n5284), .B2(n4986), .A(n4984), .ZN(n5330) );
  CLKBUF_X2 U4898 ( .A(n5361), .Z(n5325) );
  INV_X1 U4899 ( .A(n6373), .ZN(n9904) );
  INV_X1 U4900 ( .A(n6922), .ZN(n6923) );
  INV_X2 U4901 ( .A(n6337), .ZN(n5775) );
  CLKBUF_X2 U4902 ( .A(n5899), .Z(n6999) );
  INV_X4 U4904 ( .A(n8315), .ZN(n8329) );
  CLKBUF_X2 U4905 ( .A(n5215), .Z(n6495) );
  AND2_X1 U4906 ( .A1(n5869), .A2(n7824), .ZN(n6139) );
  NAND2_X2 U4907 ( .A1(n5869), .A2(n5857), .ZN(n5914) );
  INV_X4 U4908 ( .A(n8389), .ZN(n8856) );
  CLKBUF_X1 U4909 ( .A(n5815), .Z(n4353) );
  NAND2_X1 U4910 ( .A1(n6452), .A2(P1_U3086), .ZN(n9521) );
  NAND2_X1 U4911 ( .A1(n4561), .A2(n4560), .ZN(n9004) );
  AND2_X1 U4912 ( .A1(n4581), .A2(n4580), .ZN(n8388) );
  OAI21_X1 U4913 ( .B1(n6332), .B2(n9970), .A(n6331), .ZN(n6334) );
  NAND2_X2 U4914 ( .A1(n8898), .A2(n8900), .ZN(n8899) );
  OR2_X1 U4915 ( .A1(n9187), .A2(n9186), .ZN(n9379) );
  NAND2_X1 U4916 ( .A1(n7586), .A2(n7585), .ZN(n7982) );
  NOR2_X1 U4917 ( .A1(n9817), .A2(n9816), .ZN(n9815) );
  INV_X1 U4918 ( .A(n7246), .ZN(n7247) );
  NAND2_X1 U4919 ( .A1(n7202), .A2(n7201), .ZN(n7330) );
  NAND2_X1 U4920 ( .A1(n7427), .A2(n5952), .ZN(n7409) );
  NAND2_X1 U4921 ( .A1(n6075), .A2(n6074), .ZN(n8831) );
  NAND2_X1 U4922 ( .A1(n4470), .A2(n8216), .ZN(n7427) );
  NAND2_X2 U4923 ( .A1(n4448), .A2(n6064), .ZN(n8837) );
  XNOR2_X1 U4924 ( .A(n8436), .B(n4769), .ZN(n9728) );
  NAND2_X1 U4925 ( .A1(n6690), .A2(n8316), .ZN(n4448) );
  NAND2_X1 U4926 ( .A1(n5493), .A2(n5492), .ZN(n7444) );
  XNOR2_X1 U4927 ( .A(n5532), .B(n5531), .ZN(n6690) );
  OAI21_X1 U4928 ( .B1(n5514), .B2(n4975), .A(n4974), .ZN(n5532) );
  NAND2_X1 U4929 ( .A1(n6862), .A2(n6861), .ZN(n6860) );
  OR2_X2 U4930 ( .A1(n6936), .A2(n7031), .ZN(n7043) );
  INV_X2 U4931 ( .A(n9342), .ZN(n4352) );
  NAND2_X2 U4932 ( .A1(n6831), .A2(n8706), .ZN(n8710) );
  AND2_X1 U4933 ( .A1(n5256), .A2(n5255), .ZN(n9630) );
  AND2_X1 U4934 ( .A1(n4614), .A2(n8416), .ZN(n7128) );
  INV_X1 U4935 ( .A(n8345), .ZN(n9897) );
  NAND2_X1 U4936 ( .A1(n4616), .A2(n7231), .ZN(n8416) );
  INV_X1 U4937 ( .A(n7997), .ZN(n9912) );
  NAND4_X1 U4938 ( .A1(n5299), .A2(n5298), .A3(n5297), .A4(n5296), .ZN(n6922)
         );
  INV_X1 U4939 ( .A(n9044), .ZN(n6855) );
  XNOR2_X1 U4940 ( .A(n9043), .B(n6798), .ZN(n6630) );
  NAND4_X1 U4941 ( .A1(n5164), .A2(n5163), .A3(n5162), .A4(n5161), .ZN(n9045)
         );
  INV_X2 U4942 ( .A(n8321), .ZN(n8316) );
  OAI211_X1 U4943 ( .C1(n6474), .C2(n6581), .A(n5145), .B(n5144), .ZN(n6809)
         );
  NAND4_X2 U4944 ( .A1(n5219), .A2(n5218), .A3(n5217), .A4(n5216), .ZN(n9042)
         );
  OR2_X1 U4945 ( .A1(n5194), .A2(n6457), .ZN(n5145) );
  CLKBUF_X1 U4946 ( .A(n5805), .Z(n7804) );
  OR2_X1 U4947 ( .A1(n5193), .A2(n6465), .ZN(n5144) );
  INV_X2 U4948 ( .A(n5193), .ZN(n7590) );
  AND2_X1 U4949 ( .A1(n5115), .A2(n9523), .ZN(n5213) );
  NAND2_X2 U4950 ( .A1(n8000), .A2(n5114), .ZN(n6488) );
  XNOR2_X1 U4951 ( .A(n5854), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5857) );
  OR2_X1 U4952 ( .A1(n5581), .A2(n5129), .ZN(n5136) );
  XNOR2_X1 U4953 ( .A(n5112), .B(n5081), .ZN(n5815) );
  NOR2_X1 U4954 ( .A1(n6292), .A2(n4760), .ZN(n4759) );
  XNOR2_X1 U4955 ( .A(n4634), .B(n5110), .ZN(n8000) );
  NAND2_X1 U4956 ( .A1(n7557), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5112) );
  CLKBUF_X3 U4957 ( .A(n4611), .Z(n7550) );
  OAI21_X1 U4958 ( .B1(n7557), .B2(n4412), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n4634) );
  NAND2_X1 U4959 ( .A1(n5895), .A2(n5920), .ZN(n6992) );
  NAND2_X1 U4960 ( .A1(n5080), .A2(n4879), .ZN(n5091) );
  NAND2_X1 U4961 ( .A1(n6214), .A2(n4915), .ZN(n6285) );
  INV_X1 U4962 ( .A(n6450), .ZN(n5038) );
  AND2_X2 U4963 ( .A1(n5070), .A2(n5069), .ZN(n4877) );
  INV_X1 U4964 ( .A(n4998), .ZN(n6452) );
  NOR2_X1 U4965 ( .A1(n4391), .A2(n4917), .ZN(n4916) );
  AND4_X1 U4966 ( .A1(n5079), .A2(n5078), .A3(n5089), .A4(n5077), .ZN(n4374)
         );
  AND2_X1 U4967 ( .A1(n5075), .A2(n5076), .ZN(n4838) );
  AND4_X1 U4968 ( .A1(n5074), .A2(n5073), .A3(n5072), .A4(n5071), .ZN(n5075)
         );
  AND2_X1 U4969 ( .A1(n4882), .A2(n5082), .ZN(n4673) );
  AND2_X1 U4970 ( .A1(n5841), .A2(n5840), .ZN(n4890) );
  NOR2_X1 U4971 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n5071) );
  NOR2_X1 U4972 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n5072) );
  NOR2_X1 U4973 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n5073) );
  NOR2_X1 U4974 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n5074) );
  INV_X1 U4975 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4713) );
  NOR2_X1 U4976 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5189) );
  NOR2_X1 U4977 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5231) );
  NOR2_X1 U4978 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n5840) );
  NOR2_X1 U4979 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5841) );
  INV_X1 U4980 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6056) );
  INV_X1 U4981 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5838) );
  INV_X1 U4982 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6061) );
  INV_X1 U4983 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4691) );
  INV_X1 U4984 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5849) );
  NOR2_X1 U4985 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4632) );
  NOR2_X1 U4986 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4882) );
  OAI21_X2 U4987 ( .B1(n7904), .B2(n6134), .A(n8290), .ZN(n8600) );
  AND2_X1 U4988 ( .A1(n4718), .A2(n4715), .ZN(n8702) );
  OAI21_X2 U4989 ( .B1(n8612), .B2(n6126), .A(n8287), .ZN(n7904) );
  NAND2_X2 U4990 ( .A1(n6117), .A2(n8285), .ZN(n8612) );
  OAI22_X2 U4991 ( .A1(n9206), .A2(n7867), .B1(n9402), .B2(n9495), .ZN(n9191)
         );
  OAI21_X2 U4992 ( .B1(n9221), .B2(n7865), .A(n7866), .ZN(n9206) );
  OAI211_X1 U4993 ( .C1(n6474), .C2(n6580), .A(n5196), .B(n5195), .ZN(n6798)
         );
  NOR2_X4 U4994 ( .A1(n7043), .A2(n7080), .ZN(n7117) );
  AND2_X1 U4995 ( .A1(n8722), .A2(n8396), .ZN(n8379) );
  OR2_X1 U4996 ( .A1(n8327), .A2(n4588), .ZN(n4587) );
  NAND2_X1 U4997 ( .A1(n4590), .A2(n4589), .ZN(n4588) );
  INV_X1 U4998 ( .A(n8326), .ZN(n4589) );
  INV_X1 U4999 ( .A(n8325), .ZN(n4590) );
  NAND2_X1 U5000 ( .A1(n7127), .A2(n7126), .ZN(n4616) );
  OAI21_X2 U5001 ( .B1(n5561), .B2(n5560), .A(n5056), .ZN(n5580) );
  AOI21_X1 U5002 ( .B1(n4489), .B2(n4487), .A(n4439), .ZN(n4486) );
  INV_X1 U5003 ( .A(n7145), .ZN(n4487) );
  OR2_X1 U5004 ( .A1(n7146), .A2(n4488), .ZN(n4485) );
  INV_X1 U5005 ( .A(n4489), .ZN(n4488) );
  NAND2_X1 U5006 ( .A1(n4630), .A2(n4629), .ZN(n4628) );
  INV_X1 U5007 ( .A(n9850), .ZN(n4629) );
  XNOR2_X1 U5008 ( .A(n4627), .B(n8468), .ZN(n9870) );
  XNOR2_X1 U5009 ( .A(n8561), .B(n8305), .ZN(n8555) );
  NAND2_X1 U5010 ( .A1(n4460), .A2(n4457), .ZN(n7743) );
  NAND2_X1 U5011 ( .A1(n7742), .A2(n7747), .ZN(n4460) );
  OR2_X1 U5012 ( .A1(n7741), .A2(n7747), .ZN(n4457) );
  NAND2_X1 U5013 ( .A1(n4928), .A2(n4927), .ZN(n4926) );
  INV_X1 U5014 ( .A(n4930), .ZN(n4927) );
  INV_X1 U5015 ( .A(n4929), .ZN(n4928) );
  NAND2_X1 U5016 ( .A1(n5059), .A2(n10104), .ZN(n5062) );
  INV_X1 U5017 ( .A(n5310), .ZN(n4698) );
  INV_X1 U5018 ( .A(n4910), .ZN(n4909) );
  OAI21_X1 U5019 ( .B1(n8417), .B2(n4766), .A(n4764), .ZN(n7226) );
  INV_X1 U5020 ( .A(n4765), .ZN(n4764) );
  OAI21_X1 U5021 ( .B1(n8416), .B2(n4766), .A(n7225), .ZN(n4765) );
  AND2_X1 U5022 ( .A1(n4620), .A2(n4619), .ZN(n8438) );
  NAND2_X1 U5023 ( .A1(n8481), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4619) );
  NAND2_X1 U5024 ( .A1(n9778), .A2(n8441), .ZN(n8443) );
  NOR2_X1 U5025 ( .A1(n9815), .A2(n4444), .ZN(n8446) );
  OR2_X1 U5026 ( .A1(n8808), .A2(n8125), .ZN(n8287) );
  NAND2_X1 U5027 ( .A1(n4386), .A2(n4363), .ZN(n5847) );
  AND4_X1 U5028 ( .A1(n5846), .A2(n6061), .A3(n6054), .A4(n5845), .ZN(n4363)
         );
  INV_X1 U5029 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5846) );
  NAND4_X1 U5030 ( .A1(n4382), .A2(n4890), .A3(n5839), .A4(n4884), .ZN(n5994)
         );
  NOR2_X1 U5031 ( .A1(n4889), .A2(P2_IR_REG_11__SCAN_IN), .ZN(n4884) );
  AND2_X1 U5032 ( .A1(n4572), .A2(n6774), .ZN(n4571) );
  OAI21_X1 U5033 ( .B1(n8941), .B2(n4381), .A(n5578), .ZN(n4559) );
  NAND2_X1 U5034 ( .A1(n4459), .A2(n4458), .ZN(n7741) );
  OR2_X1 U5035 ( .A1(n4871), .A2(n7468), .ZN(n4870) );
  NAND2_X1 U5036 ( .A1(n4872), .A2(n7445), .ZN(n4871) );
  INV_X1 U5037 ( .A(n4875), .ZN(n4872) );
  AND2_X1 U5038 ( .A1(n7696), .A2(n7692), .ZN(n7624) );
  NOR2_X1 U5039 ( .A1(n4850), .A2(n4357), .ZN(n4849) );
  INV_X1 U5040 ( .A(n7184), .ZN(n4850) );
  INV_X1 U5041 ( .A(n8000), .ZN(n5115) );
  AND2_X1 U5042 ( .A1(n5087), .A2(n5088), .ZN(n4831) );
  INV_X1 U5043 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5088) );
  AND2_X1 U5044 ( .A1(n5717), .A2(n5696), .ZN(n5715) );
  NAND2_X1 U5045 ( .A1(n5693), .A2(n5692), .ZN(n5716) );
  OR2_X1 U5046 ( .A1(n5641), .A2(n5063), .ZN(n5065) );
  AOI21_X1 U5047 ( .B1(n4940), .B2(n4938), .A(n4937), .ZN(n4936) );
  INV_X1 U5048 ( .A(n5062), .ZN(n4937) );
  NAND2_X1 U5049 ( .A1(n4971), .A2(n4970), .ZN(n5561) );
  AOI21_X1 U5050 ( .B1(n4972), .B2(n4975), .A(n4403), .ZN(n4970) );
  NAND2_X1 U5051 ( .A1(n5354), .A2(n4990), .ZN(n5033) );
  OAI21_X2 U5052 ( .B1(n5330), .B2(n5329), .A(n5027), .ZN(n5354) );
  INV_X1 U5053 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4920) );
  OAI22_X1 U5054 ( .A1(n8014), .A2(n4513), .B1(n4515), .B2(n4436), .ZN(n4512)
         );
  NAND2_X1 U5055 ( .A1(n4905), .A2(n7935), .ZN(n4904) );
  NAND2_X1 U5056 ( .A1(n6374), .A2(n7991), .ZN(n4505) );
  AND2_X1 U5057 ( .A1(n4485), .A2(n4420), .ZN(n7316) );
  INV_X1 U5058 ( .A(n6382), .ZN(n4484) );
  AND2_X1 U5059 ( .A1(n6214), .A2(n5848), .ZN(n6217) );
  OAI21_X1 U5060 ( .B1(n4587), .B2(n4586), .A(n4397), .ZN(n4585) );
  INV_X1 U5061 ( .A(n8334), .ZN(n4586) );
  AND4_X1 U5062 ( .A1(n6071), .A2(n6070), .A3(n6069), .A4(n6068), .ZN(n8090)
         );
  AND4_X1 U5063 ( .A1(n6053), .A2(n6052), .A3(n6051), .A4(n6050), .ZN(n8258)
         );
  NAND2_X1 U5064 ( .A1(n4778), .A2(n4774), .ZN(n6985) );
  OAI21_X1 U5065 ( .B1(n7054), .B2(n4779), .A(n4414), .ZN(n4775) );
  OR2_X1 U5066 ( .A1(n9746), .A2(n9745), .ZN(n4620) );
  NAND2_X1 U5067 ( .A1(n4452), .A2(n4451), .ZN(n9778) );
  INV_X1 U5068 ( .A(n9781), .ZN(n4451) );
  NAND2_X1 U5069 ( .A1(n9797), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n4762) );
  OR2_X1 U5070 ( .A1(n9833), .A2(n8694), .ZN(n4773) );
  NAND2_X1 U5071 ( .A1(n4628), .A2(n4446), .ZN(n4627) );
  OR2_X1 U5072 ( .A1(n9870), .A2(n8669), .ZN(n4768) );
  NAND2_X1 U5073 ( .A1(n6167), .A2(n6166), .ZN(n6178) );
  AND4_X1 U5074 ( .A1(n6015), .A2(n6014), .A3(n6013), .A4(n6012), .ZN(n8117)
         );
  XNOR2_X1 U5075 ( .A(n8548), .B(n8558), .ZN(n8549) );
  NAND2_X1 U5076 ( .A1(n4749), .A2(n4751), .ZN(n4747) );
  OR2_X2 U5077 ( .A1(n8565), .A2(n8303), .ZN(n6175) );
  NOR2_X1 U5078 ( .A1(n8678), .A2(n4737), .ZN(n4736) );
  NOR2_X1 U5079 ( .A1(n4739), .A2(n6250), .ZN(n4737) );
  INV_X1 U5080 ( .A(n4716), .ZN(n4715) );
  NOR2_X1 U5081 ( .A1(n4722), .A2(n4720), .ZN(n4719) );
  INV_X1 U5082 ( .A(n8320), .ZN(n6097) );
  NAND2_X1 U5083 ( .A1(n4726), .A2(n4728), .ZN(n4725) );
  INV_X1 U5084 ( .A(n7421), .ZN(n4726) );
  INV_X1 U5085 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5860) );
  NAND2_X1 U5086 ( .A1(n5859), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5861) );
  NOR2_X2 U5087 ( .A1(n5994), .A2(n5847), .ZN(n6214) );
  AND2_X1 U5088 ( .A1(n4551), .A2(n4550), .ZN(n4549) );
  OR2_X1 U5089 ( .A1(n5595), .A2(n4558), .ZN(n4550) );
  INV_X1 U5090 ( .A(n8909), .ZN(n4815) );
  AND2_X1 U5091 ( .A1(n9482), .A2(n9163), .ZN(n7745) );
  NAND2_X1 U5092 ( .A1(n9523), .A2(n8000), .ZN(n5215) );
  INV_X1 U5093 ( .A(n7624), .ZN(n7453) );
  INV_X1 U5094 ( .A(n9647), .ZN(n9672) );
  INV_X1 U5095 ( .A(n9447), .ZN(n9680) );
  NAND2_X1 U5096 ( .A1(n6521), .A2(n4353), .ZN(n9670) );
  AND2_X1 U5097 ( .A1(n6205), .A2(n6193), .ZN(n6203) );
  NAND2_X1 U5098 ( .A1(n5763), .A2(n5762), .ZN(n6188) );
  AND2_X1 U5099 ( .A1(n6189), .A2(n5767), .ZN(n6187) );
  INV_X1 U5100 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5082) );
  AND2_X1 U5101 ( .A1(n6185), .A2(n6184), .ZN(n8305) );
  INV_X1 U5102 ( .A(n8780), .ZN(n8561) );
  NAND2_X1 U5103 ( .A1(n8237), .A2(n8239), .ZN(n4607) );
  AND2_X1 U5104 ( .A1(n8240), .A2(n8329), .ZN(n4606) );
  OR2_X1 U5105 ( .A1(n8244), .A2(n8329), .ZN(n4608) );
  OAI21_X1 U5106 ( .B1(n4409), .B2(n7810), .A(n4672), .ZN(n7695) );
  NAND2_X1 U5107 ( .A1(n7682), .A2(n7810), .ZN(n4672) );
  OAI21_X1 U5108 ( .B1(n8284), .B2(n4575), .A(n4573), .ZN(n4577) );
  OR2_X1 U5109 ( .A1(n4578), .A2(n8283), .ZN(n4575) );
  INV_X1 U5110 ( .A(n4574), .ZN(n4573) );
  AOI21_X1 U5111 ( .B1(n7704), .B2(n7787), .A(n4658), .ZN(n4657) );
  INV_X1 U5112 ( .A(n7716), .ZN(n4655) );
  NAND2_X1 U5113 ( .A1(n7703), .A2(n7705), .ZN(n4656) );
  AOI21_X1 U5114 ( .B1(n4670), .B2(n4669), .A(n4667), .ZN(n7702) );
  NAND2_X1 U5115 ( .A1(n4668), .A2(n7688), .ZN(n4667) );
  NOR2_X1 U5116 ( .A1(n4524), .A2(n4371), .ZN(n4523) );
  NOR2_X1 U5117 ( .A1(n4526), .A2(n4525), .ZN(n4524) );
  NAND2_X1 U5118 ( .A1(n4377), .A2(n7737), .ZN(n4639) );
  INV_X1 U5119 ( .A(n6189), .ZN(n4969) );
  INV_X1 U5120 ( .A(n4968), .ZN(n4967) );
  OAI21_X1 U5121 ( .B1(n6187), .B2(n4969), .A(n6203), .ZN(n4968) );
  INV_X1 U5122 ( .A(n5404), .ZN(n4981) );
  NOR2_X1 U5123 ( .A1(n4537), .A2(n8144), .ZN(n4536) );
  INV_X1 U5124 ( .A(n4540), .ZN(n4537) );
  NOR2_X1 U5125 ( .A1(n8379), .A2(n8328), .ZN(n8337) );
  AND2_X1 U5126 ( .A1(n9862), .A2(n4472), .ZN(n8501) );
  NAND2_X1 U5127 ( .A1(n8499), .A2(n9859), .ZN(n4472) );
  NAND2_X1 U5128 ( .A1(n8543), .A2(n4711), .ZN(n4710) );
  INV_X1 U5129 ( .A(n6186), .ZN(n4711) );
  OR2_X1 U5130 ( .A1(n8311), .A2(n8312), .ZN(n8377) );
  NAND2_X1 U5131 ( .A1(n8226), .A2(n8219), .ZN(n8352) );
  OR2_X1 U5132 ( .A1(n7164), .A2(n6232), .ZN(n7293) );
  NAND2_X1 U5133 ( .A1(n6228), .A2(n4742), .ZN(n4741) );
  INV_X1 U5134 ( .A(n6227), .ZN(n4742) );
  AND2_X1 U5135 ( .A1(n6297), .A2(n6542), .ZN(n6829) );
  AND2_X1 U5136 ( .A1(n6298), .A2(n6540), .ZN(n6366) );
  INV_X1 U5137 ( .A(n6261), .ZN(n4750) );
  OR2_X1 U5138 ( .A1(n8076), .A2(n8589), .ZN(n8298) );
  OR2_X1 U5139 ( .A1(n8101), .A2(n8605), .ZN(n8339) );
  OR2_X1 U5140 ( .A1(n8129), .A2(n8604), .ZN(n8291) );
  OR2_X1 U5141 ( .A1(n8744), .A2(n8656), .ZN(n6254) );
  INV_X1 U5142 ( .A(n4736), .ZN(n4734) );
  INV_X1 U5143 ( .A(n8666), .ZN(n4733) );
  NAND2_X1 U5144 ( .A1(n8831), .A2(n8680), .ZN(n4738) );
  OR2_X1 U5145 ( .A1(n8837), .A2(n8090), .ZN(n8271) );
  NAND2_X1 U5146 ( .A1(n4705), .A2(n6028), .ZN(n4704) );
  INV_X1 U5147 ( .A(n8245), .ZN(n4705) );
  AND2_X1 U5148 ( .A1(n8355), .A2(n8239), .ZN(n4707) );
  NAND2_X1 U5149 ( .A1(n6214), .A2(n4916), .ZN(n6292) );
  INV_X1 U5150 ( .A(n4917), .ZN(n4915) );
  INV_X1 U5151 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6055) );
  INV_X1 U5152 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6054) );
  NAND2_X1 U5153 ( .A1(n5838), .A2(n4713), .ZN(n4889) );
  INV_X1 U5154 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5837) );
  INV_X1 U5155 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5835) );
  INV_X1 U5156 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5836) );
  NOR2_X1 U5157 ( .A1(n9243), .A2(n9260), .ZN(n4680) );
  AND2_X1 U5158 ( .A1(n7880), .A2(n7723), .ZN(n7879) );
  NAND2_X1 U5159 ( .A1(n9253), .A2(n9252), .ZN(n7878) );
  NOR2_X1 U5160 ( .A1(n9303), .A2(n4686), .ZN(n4685) );
  INV_X1 U5161 ( .A(n4687), .ZN(n4686) );
  NOR2_X1 U5162 ( .A1(n9337), .A2(n9453), .ZN(n4687) );
  AND2_X1 U5163 ( .A1(n9293), .A2(n7705), .ZN(n4786) );
  NAND2_X1 U5164 ( .A1(n4794), .A2(n7617), .ZN(n4792) );
  AND2_X1 U5165 ( .A1(n7619), .A2(n7674), .ZN(n4794) );
  NOR2_X1 U5166 ( .A1(n9658), .A2(n9648), .ZN(n4682) );
  OR2_X1 U5167 ( .A1(n6920), .A2(n7647), .ZN(n7755) );
  NAND2_X1 U5168 ( .A1(n6789), .A2(n7761), .ZN(n7648) );
  INV_X1 U5169 ( .A(n6711), .ZN(n4660) );
  NAND2_X1 U5170 ( .A1(n4951), .A2(n4949), .ZN(n5761) );
  AOI21_X1 U5171 ( .B1(n4953), .B2(n4955), .A(n4950), .ZN(n4949) );
  INV_X1 U5172 ( .A(n5736), .ZN(n4950) );
  AND2_X1 U5173 ( .A1(n5762), .A2(n5739), .ZN(n5760) );
  NAND2_X1 U5174 ( .A1(n4925), .A2(n4923), .ZN(n5641) );
  AOI21_X1 U5175 ( .B1(n4929), .B2(n4934), .A(n4924), .ZN(n4923) );
  AND2_X1 U5176 ( .A1(n4930), .A2(n4932), .ZN(n4924) );
  AND2_X1 U5177 ( .A1(n5075), .A2(n4840), .ZN(n4839) );
  AND2_X1 U5178 ( .A1(n5076), .A2(n5085), .ZN(n4840) );
  NOR2_X1 U5179 ( .A1(n5035), .A2(n4983), .ZN(n4982) );
  INV_X1 U5180 ( .A(n5032), .ZN(n4983) );
  INV_X1 U5181 ( .A(n4987), .ZN(n4986) );
  AOI21_X1 U5182 ( .B1(n4987), .B2(n4985), .A(n4411), .ZN(n4984) );
  AOI21_X1 U5183 ( .B1(n5283), .B2(n5019), .A(n4698), .ZN(n4987) );
  NAND2_X1 U5184 ( .A1(n4700), .A2(n4699), .ZN(n5021) );
  NAND2_X1 U5185 ( .A1(n4611), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4699) );
  OR2_X1 U5186 ( .A1(n4611), .A2(n4701), .ZN(n4700) );
  OAI21_X1 U5187 ( .B1(n4998), .B2(n6466), .A(n4450), .ZN(n4995) );
  NAND2_X1 U5188 ( .A1(n4998), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4450) );
  INV_X1 U5189 ( .A(SI_5_), .ZN(n10110) );
  NAND2_X1 U5190 ( .A1(n4502), .A2(n4503), .ZN(n4495) );
  INV_X1 U5191 ( .A(n7967), .ZN(n4895) );
  NAND2_X1 U5192 ( .A1(n8154), .A2(n4901), .ZN(n4900) );
  XNOR2_X1 U5193 ( .A(n6370), .B(n9912), .ZN(n6371) );
  AOI21_X1 U5194 ( .B1(n4911), .B2(n4358), .A(n4392), .ZN(n4910) );
  OR2_X1 U5195 ( .A1(n6048), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U5196 ( .A1(n4445), .A2(n4373), .ZN(n4528) );
  AOI21_X1 U5197 ( .B1(n4445), .B2(n4364), .A(n4516), .ZN(n8113) );
  NAND2_X1 U5198 ( .A1(n4517), .A2(n4438), .ZN(n4516) );
  OAI21_X1 U5199 ( .B1(n4909), .B2(n4531), .A(n4907), .ZN(n4530) );
  NAND2_X1 U5200 ( .A1(n4534), .A2(n4535), .ZN(n4531) );
  AOI21_X1 U5201 ( .B1(n4910), .B2(n4912), .A(n4908), .ZN(n4907) );
  INV_X1 U5202 ( .A(n8053), .ZN(n4908) );
  NOR2_X1 U5203 ( .A1(n4909), .A2(n4533), .ZN(n4532) );
  INV_X1 U5204 ( .A(n4534), .ZN(n4533) );
  NAND2_X1 U5205 ( .A1(n4543), .A2(n4541), .ZN(n4540) );
  INV_X1 U5206 ( .A(n4546), .ZN(n4543) );
  NAND2_X1 U5207 ( .A1(n8088), .A2(n4542), .ZN(n4541) );
  INV_X1 U5208 ( .A(n8080), .ZN(n4542) );
  NOR2_X1 U5209 ( .A1(n4490), .A2(n4492), .ZN(n4489) );
  INV_X1 U5210 ( .A(n7155), .ZN(n4490) );
  AND2_X1 U5211 ( .A1(n4904), .A2(n4442), .ZN(n4902) );
  AND4_X1 U5212 ( .A1(n6125), .A2(n6124), .A3(n6123), .A4(n6122), .ZN(n8125)
         );
  AND4_X1 U5213 ( .A1(n5948), .A2(n5947), .A3(n5946), .A4(n5945), .ZN(n7318)
         );
  OAI21_X1 U5214 ( .B1(n6896), .B2(n6438), .A(n6909), .ZN(n6440) );
  XNOR2_X1 U5215 ( .A(n7062), .B(n6908), .ZN(n7056) );
  AOI21_X1 U5216 ( .B1(n6898), .B2(n7062), .A(n7051), .ZN(n6900) );
  NAND2_X1 U5217 ( .A1(n6981), .A2(n6982), .ZN(n7127) );
  NAND2_X1 U5218 ( .A1(n4618), .A2(n8486), .ZN(n4617) );
  INV_X1 U5219 ( .A(n4772), .ZN(n9704) );
  NOR2_X1 U5220 ( .A1(n9728), .A2(n5973), .ZN(n9727) );
  NOR2_X1 U5221 ( .A1(n9727), .A2(n4621), .ZN(n9746) );
  AND2_X1 U5222 ( .A1(n8436), .A2(n4769), .ZN(n4621) );
  NAND2_X1 U5223 ( .A1(n9735), .A2(n8492), .ZN(n9756) );
  OR2_X1 U5224 ( .A1(n9761), .A2(n8439), .ZN(n4452) );
  XNOR2_X1 U5225 ( .A(n8443), .B(n8475), .ZN(n9796) );
  NAND2_X1 U5226 ( .A1(n9844), .A2(n9845), .ZN(n9843) );
  NAND2_X1 U5227 ( .A1(n4773), .A2(n4385), .ZN(n4630) );
  NAND2_X1 U5228 ( .A1(n8467), .A2(n9860), .ZN(n8515) );
  INV_X1 U5229 ( .A(n6130), .ZN(n6129) );
  AOI21_X1 U5230 ( .B1(n8655), .B2(n6253), .A(n4410), .ZN(n8640) );
  OR2_X1 U5231 ( .A1(n5999), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6010) );
  OR2_X1 U5232 ( .A1(n5903), .A2(n6908), .ZN(n5881) );
  NOR2_X1 U5233 ( .A1(n6262), .A2(n4750), .ZN(n4748) );
  OR2_X1 U5234 ( .A1(n8303), .A2(n8302), .ZN(n8566) );
  OR2_X1 U5235 ( .A1(n8577), .A2(n8582), .ZN(n8575) );
  INV_X1 U5236 ( .A(n9880), .ZN(n9891) );
  NAND2_X1 U5237 ( .A1(n6410), .A2(n8329), .ZN(n9893) );
  INV_X1 U5238 ( .A(n9883), .ZN(n9899) );
  AOI21_X1 U5239 ( .B1(n4736), .B2(n4739), .A(n4370), .ZN(n4735) );
  AND2_X1 U5240 ( .A1(n8843), .A2(n8703), .ZN(n4739) );
  AND2_X2 U5241 ( .A1(n8271), .A2(n8266), .ZN(n8678) );
  NAND2_X1 U5242 ( .A1(n6239), .A2(n7397), .ZN(n6246) );
  AOI21_X1 U5243 ( .B1(n4723), .B2(n6247), .A(n4416), .ZN(n4721) );
  AND2_X1 U5244 ( .A1(n6409), .A2(n8329), .ZN(n9880) );
  NOR2_X1 U5245 ( .A1(n8355), .A2(n4724), .ZN(n4723) );
  INV_X1 U5246 ( .A(n4727), .ZN(n4724) );
  NAND2_X1 U5247 ( .A1(n4725), .A2(n4727), .ZN(n7477) );
  INV_X1 U5248 ( .A(n9893), .ZN(n9878) );
  NAND2_X1 U5249 ( .A1(n6006), .A2(n4707), .ZN(n7483) );
  NAND2_X1 U5250 ( .A1(n6324), .A2(n8382), .ZN(n9883) );
  NAND2_X1 U5251 ( .A1(n4483), .A2(n6296), .ZN(n6506) );
  AND2_X1 U5252 ( .A1(n6214), .A2(n4421), .ZN(n5853) );
  NOR2_X1 U5253 ( .A1(n4760), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n4758) );
  NOR2_X1 U5254 ( .A1(n4889), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n4888) );
  NOR2_X1 U5255 ( .A1(n4887), .A2(n4885), .ZN(n5992) );
  NAND2_X1 U5256 ( .A1(n4382), .A2(n4890), .ZN(n4887) );
  NAND2_X1 U5257 ( .A1(n5839), .A2(n4886), .ZN(n4885) );
  INV_X1 U5258 ( .A(n4889), .ZN(n4886) );
  INV_X1 U5259 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n4623) );
  NAND2_X1 U5260 ( .A1(n5349), .A2(n5352), .ZN(n4837) );
  INV_X1 U5261 ( .A(n5347), .ZN(n5345) );
  INV_X1 U5262 ( .A(n8974), .ZN(n4817) );
  NOR2_X1 U5263 ( .A1(n8952), .A2(n4823), .ZN(n4822) );
  INV_X1 U5264 ( .A(n8874), .ZN(n4824) );
  OR2_X1 U5265 ( .A1(n8952), .A2(n4824), .ZN(n4821) );
  NAND2_X1 U5266 ( .A1(n8899), .A2(n5619), .ZN(n8974) );
  INV_X1 U5267 ( .A(n5606), .ZN(n5108) );
  NAND2_X1 U5268 ( .A1(n4566), .A2(n4564), .ZN(n8982) );
  AOI21_X1 U5269 ( .B1(n4567), .B2(n4813), .A(n4565), .ZN(n4564) );
  INV_X1 U5270 ( .A(n5664), .ZN(n4565) );
  NAND2_X1 U5271 ( .A1(n4559), .A2(n5595), .ZN(n5596) );
  NAND2_X1 U5272 ( .A1(n4556), .A2(n5594), .ZN(n5598) );
  INV_X1 U5273 ( .A(n4559), .ZN(n4556) );
  OR2_X1 U5274 ( .A1(n5586), .A2(n5585), .ZN(n5606) );
  OR2_X1 U5275 ( .A1(n5723), .A2(n8917), .ZN(n5742) );
  NOR2_X1 U5276 ( .A1(n5812), .A2(n7807), .ZN(n5809) );
  NAND2_X1 U5277 ( .A1(n4961), .A2(n7815), .ZN(n4960) );
  INV_X1 U5278 ( .A(n7637), .ZN(n4961) );
  NOR2_X1 U5279 ( .A1(n7750), .A2(n4453), .ZN(n7808) );
  OAI21_X1 U5280 ( .B1(n7749), .B2(n4455), .A(n4454), .ZN(n4453) );
  AOI211_X1 U5281 ( .C1(n9163), .C2(n7893), .A(n7745), .B(n7744), .ZN(n7750)
         );
  NAND2_X1 U5282 ( .A1(n4456), .A2(n7893), .ZN(n4455) );
  NAND2_X1 U5283 ( .A1(n4633), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5151) );
  INV_X1 U5284 ( .A(n4790), .ZN(n4789) );
  OAI21_X1 U5285 ( .B1(n7883), .B2(n7727), .A(n9185), .ZN(n4790) );
  NAND2_X1 U5286 ( .A1(n4651), .A2(n7870), .ZN(n4864) );
  NAND2_X1 U5287 ( .A1(n7887), .A2(n4866), .ZN(n4865) );
  AND2_X1 U5288 ( .A1(n4651), .A2(n4867), .ZN(n4863) );
  INV_X1 U5289 ( .A(n4689), .ZN(n9167) );
  NOR2_X1 U5290 ( .A1(n9185), .A2(n4868), .ZN(n4867) );
  INV_X1 U5291 ( .A(n7868), .ZN(n4868) );
  AND2_X1 U5292 ( .A1(n7731), .A2(n7886), .ZN(n9185) );
  NAND2_X1 U5293 ( .A1(n9218), .A2(n9217), .ZN(n9216) );
  NAND2_X1 U5294 ( .A1(n9265), .A2(n4676), .ZN(n9207) );
  NOR2_X1 U5295 ( .A1(n4677), .A2(n9209), .ZN(n4676) );
  INV_X1 U5296 ( .A(n4678), .ZN(n4677) );
  NAND2_X1 U5297 ( .A1(n9310), .A2(n4786), .ZN(n9292) );
  NAND2_X1 U5298 ( .A1(n9312), .A2(n9311), .ZN(n9310) );
  NOR2_X1 U5299 ( .A1(n7446), .A2(n4876), .ZN(n4875) );
  INV_X1 U5300 ( .A(n7331), .ZN(n4876) );
  INV_X1 U5301 ( .A(n4853), .ZN(n4852) );
  OR2_X1 U5302 ( .A1(n9601), .A2(n9654), .ZN(n7678) );
  AND2_X1 U5303 ( .A1(n7679), .A2(n7772), .ZN(n7620) );
  NAND2_X1 U5304 ( .A1(n7186), .A2(n4794), .ZN(n9593) );
  INV_X1 U5305 ( .A(n7620), .ZN(n7199) );
  NAND2_X1 U5306 ( .A1(n5385), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5440) );
  NAND2_X1 U5307 ( .A1(n7185), .A2(n7184), .ZN(n9591) );
  INV_X1 U5308 ( .A(n7619), .ZN(n9595) );
  BUF_X1 U5309 ( .A(n6488), .Z(n6494) );
  OR2_X1 U5310 ( .A1(n5336), .A2(n5335), .ZN(n5364) );
  NAND2_X1 U5311 ( .A1(n4857), .A2(n4854), .ZN(n7033) );
  NAND2_X1 U5312 ( .A1(n6700), .A2(n6699), .ZN(n6926) );
  NAND2_X1 U5313 ( .A1(n7648), .A2(n7650), .ZN(n6715) );
  INV_X1 U5314 ( .A(n7608), .ZN(n6836) );
  NAND2_X1 U5315 ( .A1(n6836), .A2(n6837), .ZN(n6835) );
  XNOR2_X1 U5316 ( .A(n9623), .B(n9042), .ZN(n7608) );
  OR2_X1 U5317 ( .A1(n6673), .A2(n6548), .ZN(n9348) );
  NAND2_X1 U5318 ( .A1(n5769), .A2(n5768), .ZN(n9193) );
  OR2_X1 U5319 ( .A1(n6673), .A2(n7803), .ZN(n9664) );
  INV_X1 U5320 ( .A(n8891), .ZN(n9623) );
  INV_X1 U5321 ( .A(n9670), .ZN(n9441) );
  NAND2_X1 U5322 ( .A1(n6526), .A2(n7811), .ZN(n9447) );
  NAND2_X1 U5323 ( .A1(n7584), .A2(n7548), .ZN(n7589) );
  XNOR2_X1 U5324 ( .A(n7589), .B(n7588), .ZN(n8317) );
  OR2_X1 U5325 ( .A1(n6206), .A2(SI_29_), .ZN(n7583) );
  NAND2_X1 U5326 ( .A1(n6206), .A2(SI_29_), .ZN(n7584) );
  AND2_X1 U5327 ( .A1(n4632), .A2(n4631), .ZN(n5079) );
  XNOR2_X1 U5328 ( .A(n5092), .B(P1_IR_REG_26__SCAN_IN), .ZN(n5799) );
  XNOR2_X1 U5329 ( .A(n5761), .B(n5760), .ZN(n7522) );
  NAND2_X1 U5330 ( .A1(n4952), .A2(n5717), .ZN(n5735) );
  NAND2_X1 U5331 ( .A1(n5716), .A2(n5715), .ZN(n4952) );
  NAND2_X1 U5332 ( .A1(n5080), .A2(n4374), .ZN(n5093) );
  AOI21_X1 U5333 ( .B1(n4361), .B2(P1_IR_REG_31__SCAN_IN), .A(n4830), .ZN(
        n4829) );
  OAI21_X1 U5334 ( .B1(n5667), .B2(n5666), .A(n5668), .ZN(n5691) );
  AND2_X1 U5335 ( .A1(n5692), .A2(n5672), .ZN(n5690) );
  XNOR2_X1 U5336 ( .A(n5803), .B(P1_IR_REG_23__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U5337 ( .A1(n5802), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5803) );
  NAND2_X1 U5338 ( .A1(n4380), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U5339 ( .A1(n5580), .A2(n4938), .ZN(n4935) );
  OAI21_X1 U5340 ( .B1(n5580), .B2(n4940), .A(n5058), .ZN(n5600) );
  AND2_X2 U5341 ( .A1(n4838), .A2(n4877), .ZN(n5080) );
  NAND2_X1 U5342 ( .A1(n5033), .A2(n5032), .ZN(n5379) );
  NAND2_X1 U5343 ( .A1(n5002), .A2(n5001), .ZN(n5206) );
  OAI21_X1 U5344 ( .B1(n6468), .B2(n8321), .A(n4467), .ZN(n6406) );
  AND2_X1 U5345 ( .A1(n5951), .A2(n4388), .ZN(n4467) );
  NOR2_X1 U5346 ( .A1(n4355), .A2(n8164), .ZN(n4509) );
  NAND2_X1 U5347 ( .A1(n4512), .A2(n4401), .ZN(n4511) );
  INV_X1 U5348 ( .A(n8399), .ZN(n8605) );
  OAI21_X1 U5349 ( .B1(n8258), .B2(n7938), .A(n8166), .ZN(n8082) );
  NAND2_X1 U5350 ( .A1(n7961), .A2(n7960), .ZN(n8156) );
  AND2_X1 U5351 ( .A1(n6047), .A2(n6046), .ZN(n8259) );
  INV_X1 U5352 ( .A(n8692), .ZN(n8173) );
  XNOR2_X1 U5353 ( .A(n6220), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8391) );
  NAND2_X1 U5354 ( .A1(n6217), .A2(n5849), .ZN(n6219) );
  INV_X1 U5355 ( .A(n4585), .ZN(n4584) );
  XNOR2_X1 U5356 ( .A(n6096), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8516) );
  OAI21_X1 U5357 ( .B1(n6095), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6096) );
  INV_X1 U5358 ( .A(n8305), .ZN(n8568) );
  NAND2_X1 U5359 ( .A1(n6174), .A2(n6173), .ZN(n8398) );
  INV_X1 U5360 ( .A(n8589), .ZN(n8569) );
  INV_X1 U5361 ( .A(n8146), .ZN(n8680) );
  INV_X1 U5362 ( .A(n8258), .ZN(n8703) );
  NAND4_X2 U5363 ( .A1(n5893), .A2(n5892), .A3(n5891), .A4(n5890), .ZN(n9881)
         );
  OR2_X1 U5364 ( .A1(n7003), .A2(n5888), .ZN(n5892) );
  NAND2_X1 U5365 ( .A1(n4768), .A2(n4384), .ZN(n4767) );
  INV_X1 U5366 ( .A(n4627), .ZN(n8448) );
  AOI211_X1 U5367 ( .C1(P2_ADDR_REG_18__SCAN_IN), .C2(n9857), .A(n8505), .B(
        n8504), .ZN(n8506) );
  AND2_X1 U5368 ( .A1(n4767), .A2(n4626), .ZN(n8512) );
  INV_X1 U5369 ( .A(n8450), .ZN(n4626) );
  OR2_X1 U5370 ( .A1(n8512), .A2(n4625), .ZN(n4624) );
  NOR2_X1 U5371 ( .A1(n8521), .A2(n8658), .ZN(n4625) );
  INV_X1 U5372 ( .A(n8802), .ZN(n8609) );
  OAI21_X1 U5373 ( .B1(n4359), .B2(n4610), .A(n6281), .ZN(n4609) );
  NAND2_X1 U5374 ( .A1(n6505), .A2(n6404), .ZN(n8706) );
  OAI22_X1 U5375 ( .A1(n8778), .A2(n8734), .B1(n9986), .B2(n8723), .ZN(n4753)
         );
  NOR2_X1 U5376 ( .A1(n9984), .A2(n9962), .ZN(n8762) );
  AND2_X1 U5377 ( .A1(n4756), .A2(n4754), .ZN(n8773) );
  AOI21_X1 U5378 ( .B1(n8545), .B2(n9878), .A(n4755), .ZN(n4754) );
  NAND2_X1 U5379 ( .A1(n4757), .A2(n9883), .ZN(n4756) );
  AND2_X1 U5380 ( .A1(n8568), .A2(n9880), .ZN(n4755) );
  NAND2_X1 U5381 ( .A1(n4708), .A2(n6186), .ZN(n8550) );
  NAND2_X1 U5382 ( .A1(n6175), .A2(n4712), .ZN(n4708) );
  AND2_X1 U5383 ( .A1(n6177), .A2(n6176), .ZN(n8780) );
  NAND2_X1 U5384 ( .A1(n6336), .A2(n6335), .ZN(n9183) );
  AND2_X1 U5385 ( .A1(n5464), .A2(n5463), .ZN(n7381) );
  INV_X1 U5386 ( .A(n9042), .ZN(n8966) );
  INV_X1 U5387 ( .A(n9671), .ZN(n9033) );
  INV_X1 U5388 ( .A(n9654), .ZN(n9036) );
  INV_X1 U5389 ( .A(n7114), .ZN(n9646) );
  NAND3_X2 U5390 ( .A1(n5188), .A2(n5187), .A3(n5186), .ZN(n9043) );
  AND2_X1 U5391 ( .A1(n5185), .A2(n5184), .ZN(n5186) );
  AND2_X1 U5392 ( .A1(n6599), .A2(n6576), .ZN(n9580) );
  NAND2_X1 U5393 ( .A1(n4802), .A2(n4800), .ZN(n7460) );
  OR2_X1 U5394 ( .A1(n5194), .A2(n6454), .ZN(n5195) );
  AND2_X1 U5395 ( .A1(n7598), .A2(n7597), .ZN(n9482) );
  OR2_X1 U5396 ( .A1(n8322), .A2(n5193), .ZN(n7598) );
  INV_X1 U5397 ( .A(n7982), .ZN(n4459) );
  OR2_X1 U5398 ( .A1(n5193), .A2(n6458), .ZN(n5236) );
  OR2_X1 U5399 ( .A1(n7492), .A2(n5799), .ZN(n9520) );
  NAND2_X1 U5400 ( .A1(n4592), .A2(n8329), .ZN(n4591) );
  NAND2_X1 U5401 ( .A1(n4594), .A2(n4593), .ZN(n4592) );
  NOR2_X1 U5402 ( .A1(n8352), .A2(n8205), .ZN(n4593) );
  NAND2_X1 U5403 ( .A1(n8207), .A2(n8206), .ZN(n4594) );
  AND2_X1 U5404 ( .A1(n8220), .A2(n8315), .ZN(n4596) );
  OAI21_X1 U5405 ( .B1(n6715), .B2(n7652), .A(n4665), .ZN(n4664) );
  INV_X1 U5406 ( .A(n7655), .ZN(n4665) );
  NAND2_X1 U5407 ( .A1(n4607), .A2(n4606), .ZN(n4605) );
  NAND2_X1 U5408 ( .A1(n4666), .A2(n4662), .ZN(n7662) );
  NAND2_X1 U5409 ( .A1(n4664), .A2(n4663), .ZN(n4662) );
  NAND2_X1 U5410 ( .A1(n7657), .A2(n7810), .ZN(n4666) );
  NOR2_X1 U5411 ( .A1(n7647), .A2(n7810), .ZN(n4663) );
  INV_X1 U5412 ( .A(n6927), .ZN(n7661) );
  OAI21_X1 U5413 ( .B1(n4578), .B2(n4404), .A(n8287), .ZN(n4574) );
  NAND2_X1 U5414 ( .A1(n8286), .A2(n8285), .ZN(n4578) );
  NAND2_X1 U5415 ( .A1(n7698), .A2(n7699), .ZN(n4668) );
  NAND2_X1 U5416 ( .A1(n4671), .A2(n4395), .ZN(n4670) );
  NAND2_X1 U5417 ( .A1(n7695), .A2(n7776), .ZN(n4671) );
  NOR2_X1 U5418 ( .A1(n7779), .A2(n7697), .ZN(n4669) );
  AOI21_X1 U5419 ( .B1(n8294), .B2(n8293), .A(n8292), .ZN(n4604) );
  INV_X1 U5420 ( .A(n4602), .ZN(n4601) );
  OAI21_X1 U5421 ( .B1(n8295), .B2(n8329), .A(n8339), .ZN(n4602) );
  INV_X1 U5422 ( .A(n8295), .ZN(n4603) );
  NOR2_X1 U5423 ( .A1(n4654), .A2(n7715), .ZN(n4653) );
  AOI21_X1 U5424 ( .B1(n4657), .B2(n4656), .A(n4655), .ZN(n4654) );
  NAND2_X1 U5425 ( .A1(n4600), .A2(n4598), .ZN(n8301) );
  AND2_X1 U5426 ( .A1(n4599), .A2(n8582), .ZN(n4598) );
  OAI21_X1 U5427 ( .B1(n4604), .B2(n4603), .A(n4601), .ZN(n4600) );
  OR2_X1 U5428 ( .A1(n8296), .A2(n8329), .ZN(n4599) );
  INV_X1 U5429 ( .A(n4649), .ZN(n4644) );
  AND2_X1 U5430 ( .A1(n9173), .A2(n7810), .ZN(n4649) );
  OR2_X1 U5431 ( .A1(n7927), .A2(n8059), .ZN(n8236) );
  AOI21_X1 U5432 ( .B1(n4747), .B2(n4745), .A(n4405), .ZN(n4744) );
  INV_X1 U5433 ( .A(n4748), .ZN(n4745) );
  NAND2_X1 U5434 ( .A1(n4417), .A2(n5848), .ZN(n4917) );
  INV_X1 U5435 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n4918) );
  INV_X1 U5436 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5844) );
  AND2_X1 U5437 ( .A1(n5595), .A2(n4558), .ZN(n4557) );
  NAND2_X1 U5438 ( .A1(n6887), .A2(n6888), .ZN(n4572) );
  OR2_X1 U5439 ( .A1(n4650), .A2(n4649), .ZN(n4643) );
  NOR2_X1 U5440 ( .A1(n4379), .A2(n4642), .ZN(n4641) );
  NOR2_X1 U5441 ( .A1(n7739), .A2(n7738), .ZN(n4642) );
  NAND2_X1 U5442 ( .A1(n7886), .A2(n7747), .ZN(n4652) );
  NAND2_X1 U5443 ( .A1(n4646), .A2(n4651), .ZN(n4645) );
  INV_X1 U5444 ( .A(n7743), .ZN(n4646) );
  AND2_X1 U5445 ( .A1(n9353), .A2(n9030), .ZN(n7700) );
  AND2_X1 U5446 ( .A1(n9516), .A2(n9313), .ZN(n7701) );
  AND2_X1 U5447 ( .A1(n8935), .A2(n9031), .ZN(n7687) );
  INV_X1 U5448 ( .A(n5717), .ZN(n4955) );
  INV_X1 U5449 ( .A(n4954), .ZN(n4953) );
  OAI21_X1 U5450 ( .B1(n5715), .B2(n4955), .A(n5734), .ZN(n4954) );
  AOI21_X1 U5451 ( .B1(n4936), .B2(n4931), .A(SI_20_), .ZN(n4930) );
  INV_X1 U5452 ( .A(n4936), .ZN(n4932) );
  AOI21_X1 U5453 ( .B1(n4933), .B2(n4931), .A(n5620), .ZN(n4929) );
  NOR2_X1 U5454 ( .A1(n5052), .A2(n4973), .ZN(n4972) );
  NOR2_X1 U5455 ( .A1(n5530), .A2(SI_16_), .ZN(n5052) );
  INV_X1 U5456 ( .A(n4974), .ZN(n4973) );
  INV_X1 U5457 ( .A(n5019), .ZN(n4985) );
  INV_X1 U5458 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4690) );
  INV_X1 U5459 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4922) );
  INV_X1 U5460 ( .A(SI_18_), .ZN(n10155) );
  OR2_X1 U5461 ( .A1(n4522), .A2(n4518), .ZN(n4517) );
  INV_X1 U5462 ( .A(n7933), .ZN(n4518) );
  AND2_X1 U5463 ( .A1(n4988), .A2(n4523), .ZN(n4522) );
  INV_X1 U5464 ( .A(n8105), .ZN(n4913) );
  OR2_X1 U5465 ( .A1(n8045), .A2(n4358), .ZN(n4914) );
  INV_X1 U5466 ( .A(n8020), .ZN(n4905) );
  OR2_X1 U5467 ( .A1(n4779), .A2(n6911), .ZN(n4776) );
  NAND2_X1 U5468 ( .A1(n8426), .A2(n7236), .ZN(n8453) );
  NAND2_X1 U5469 ( .A1(n9706), .A2(n4770), .ZN(n8436) );
  OR2_X1 U5470 ( .A1(n8489), .A2(n8435), .ZN(n4770) );
  OAI21_X1 U5471 ( .B1(n9734), .B2(n8452), .A(n9738), .ZN(n8458) );
  NAND2_X1 U5472 ( .A1(n8460), .A2(n9769), .ZN(n8461) );
  OAI21_X1 U5473 ( .B1(n9839), .B2(n8754), .A(n9840), .ZN(n8466) );
  AND2_X1 U5474 ( .A1(n8236), .A2(n8221), .ZN(n8224) );
  NAND2_X1 U5475 ( .A1(n7997), .A2(n9892), .ZN(n5876) );
  AND2_X1 U5476 ( .A1(n8338), .A2(n8593), .ZN(n8295) );
  INV_X1 U5477 ( .A(n8252), .ZN(n4720) );
  OAI21_X1 U5478 ( .B1(n4721), .B2(n4720), .A(n4717), .ZN(n4716) );
  OR2_X1 U5479 ( .A1(n9966), .A2(n8402), .ZN(n4727) );
  AND2_X1 U5480 ( .A1(n7296), .A2(n6235), .ZN(n7433) );
  XNOR2_X1 U5481 ( .A(n7476), .B(P2_B_REG_SCAN_IN), .ZN(n4481) );
  NAND2_X1 U5482 ( .A1(n5850), .A2(n4761), .ZN(n4760) );
  INV_X1 U5483 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4761) );
  INV_X1 U5484 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5842) );
  INV_X1 U5485 ( .A(n8995), .ZN(n4558) );
  NOR2_X1 U5486 ( .A1(n4557), .A2(n4555), .ZN(n4554) );
  INV_X1 U5487 ( .A(n5578), .ZN(n4555) );
  OR2_X1 U5488 ( .A1(n4557), .A2(n4552), .ZN(n4551) );
  NAND2_X1 U5489 ( .A1(n4381), .A2(n5578), .ZN(n4552) );
  AND2_X1 U5490 ( .A1(n5102), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n5257) );
  XNOR2_X1 U5491 ( .A(n5223), .B(n5222), .ZN(n5273) );
  AOI21_X1 U5492 ( .B1(n4814), .B2(n4569), .A(n4568), .ZN(n4567) );
  INV_X1 U5493 ( .A(n5619), .ZN(n4569) );
  INV_X1 U5494 ( .A(n4812), .ZN(n4568) );
  AOI21_X1 U5495 ( .B1(n4814), .B2(n8972), .A(n4402), .ZN(n4812) );
  NOR2_X1 U5496 ( .A1(n5467), .A2(n5466), .ZN(n5465) );
  INV_X1 U5497 ( .A(n9482), .ZN(n4456) );
  INV_X1 U5498 ( .A(n6488), .ZN(n4633) );
  NOR2_X1 U5499 ( .A1(n9231), .A2(n4679), .ZN(n4678) );
  INV_X1 U5500 ( .A(n4680), .ZN(n4679) );
  INV_X1 U5501 ( .A(n7700), .ZN(n7783) );
  INV_X1 U5502 ( .A(n7687), .ZN(n7698) );
  OAI21_X1 U5503 ( .B1(n9595), .B2(n4357), .A(n7199), .ZN(n4853) );
  AND2_X1 U5504 ( .A1(n7776), .A2(n7773), .ZN(n7621) );
  AND2_X1 U5505 ( .A1(n5105), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n5385) );
  INV_X1 U5506 ( .A(n6925), .ZN(n4859) );
  NOR2_X1 U5507 ( .A1(n4859), .A2(n4856), .ZN(n4855) );
  INV_X1 U5508 ( .A(n6698), .ZN(n4856) );
  INV_X1 U5509 ( .A(n6695), .ZN(n4847) );
  NOR2_X1 U5510 ( .A1(n4847), .A2(n4846), .ZN(n4845) );
  INV_X1 U5511 ( .A(n6693), .ZN(n4846) );
  OR2_X1 U5512 ( .A1(n5805), .A2(n7844), .ZN(n6523) );
  NAND2_X1 U5513 ( .A1(n9334), .A2(n9516), .ZN(n9335) );
  AOI21_X1 U5514 ( .B1(n4967), .B2(n4969), .A(n4965), .ZN(n4964) );
  INV_X1 U5515 ( .A(n6205), .ZN(n4965) );
  INV_X1 U5516 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5076) );
  XNOR2_X1 U5517 ( .A(n7547), .B(n7545), .ZN(n6206) );
  INV_X1 U5518 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n4631) );
  NAND2_X1 U5519 ( .A1(n5122), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5124) );
  INV_X1 U5520 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5123) );
  NOR2_X1 U5521 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5128) );
  INV_X1 U5522 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5127) );
  INV_X1 U5523 ( .A(n5058), .ZN(n4939) );
  INV_X1 U5524 ( .A(n5579), .ZN(n4940) );
  NAND2_X1 U5525 ( .A1(n5051), .A2(n4976), .ZN(n4974) );
  NOR2_X1 U5526 ( .A1(n5051), .A2(n4976), .ZN(n4975) );
  INV_X1 U5527 ( .A(n4979), .ZN(n4978) );
  OAI21_X1 U5528 ( .B1(n4982), .B2(n4980), .A(n5043), .ZN(n4979) );
  NAND2_X1 U5529 ( .A1(n4981), .A2(n5037), .ZN(n4980) );
  INV_X1 U5530 ( .A(n5010), .ZN(n4942) );
  OAI21_X1 U5531 ( .B1(n5038), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n4461), .ZN(
        n5007) );
  NAND2_X1 U5532 ( .A1(n5038), .A2(n5230), .ZN(n4461) );
  INV_X1 U5533 ( .A(SI_19_), .ZN(n10104) );
  INV_X1 U5534 ( .A(SI_17_), .ZN(n10074) );
  INV_X1 U5535 ( .A(n8154), .ZN(n4513) );
  INV_X1 U5536 ( .A(n4536), .ZN(n4535) );
  AOI21_X1 U5537 ( .B1(n4536), .B2(n4544), .A(n4368), .ZN(n4534) );
  NAND2_X1 U5538 ( .A1(n6065), .A2(n10109), .ZN(n6076) );
  INV_X1 U5539 ( .A(n6066), .ZN(n6065) );
  NOR2_X1 U5540 ( .A1(n4504), .A2(n6735), .ZN(n4501) );
  NAND2_X1 U5541 ( .A1(n4494), .A2(n4505), .ZN(n4499) );
  NAND2_X1 U5542 ( .A1(n8113), .A2(n8112), .ZN(n8111) );
  INV_X1 U5543 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10107) );
  AND2_X1 U5544 ( .A1(n8240), .A2(n8239), .ZN(n8356) );
  NAND2_X1 U5545 ( .A1(n4520), .A2(n4519), .ZN(n8060) );
  OR2_X1 U5546 ( .A1(n4371), .A2(n7922), .ZN(n4519) );
  NAND2_X1 U5547 ( .A1(n4528), .A2(n4521), .ZN(n4520) );
  NOR2_X1 U5548 ( .A1(n4527), .A2(n4371), .ZN(n4521) );
  NAND2_X1 U5549 ( .A1(n6372), .A2(n9892), .ZN(n4506) );
  OR2_X1 U5550 ( .A1(n6076), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6088) );
  NAND2_X1 U5551 ( .A1(n7146), .A2(n7145), .ZN(n4491) );
  OAI21_X1 U5552 ( .B1(n8331), .B2(n8548), .A(n4583), .ZN(n4582) );
  AND2_X1 U5553 ( .A1(n4587), .A2(n4424), .ZN(n4583) );
  OR2_X1 U5554 ( .A1(n6082), .A2(P2_IR_REG_17__SCAN_IN), .ZN(n6095) );
  AND2_X1 U5555 ( .A1(n7007), .A2(n7006), .ZN(n8380) );
  AND2_X1 U5556 ( .A1(n7007), .A2(n6213), .ZN(n8312) );
  OR2_X1 U5557 ( .A1(n5914), .A2(n6431), .ZN(n5864) );
  OR2_X1 U5558 ( .A1(n6109), .A2(n5868), .ZN(n6223) );
  NAND2_X1 U5559 ( .A1(n7059), .A2(n7058), .ZN(n7057) );
  NAND2_X1 U5560 ( .A1(n4615), .A2(n7130), .ZN(n4614) );
  INV_X1 U5561 ( .A(n4616), .ZN(n4615) );
  NAND2_X1 U5562 ( .A1(n7125), .A2(n7124), .ZN(n7232) );
  NOR2_X1 U5563 ( .A1(n7134), .A2(n4462), .ZN(n7137) );
  NOR2_X1 U5564 ( .A1(n4464), .A2(n4463), .ZN(n4462) );
  INV_X1 U5565 ( .A(n7135), .ZN(n4464) );
  INV_X1 U5566 ( .A(n7136), .ZN(n4463) );
  AOI21_X1 U5567 ( .B1(n7223), .B2(n7231), .A(n7222), .ZN(n8413) );
  NAND2_X1 U5568 ( .A1(n4763), .A2(n8415), .ZN(n8419) );
  NAND2_X1 U5569 ( .A1(n8417), .A2(n8416), .ZN(n4763) );
  NAND2_X1 U5570 ( .A1(n4771), .A2(n9703), .ZN(n9706) );
  NAND2_X1 U5571 ( .A1(n4772), .A2(n8434), .ZN(n4771) );
  OR2_X1 U5572 ( .A1(n9698), .A2(n9697), .ZN(n9701) );
  OR2_X1 U5573 ( .A1(n5962), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5966) );
  OAI22_X1 U5574 ( .A1(n9714), .A2(n9713), .B1(n8490), .B2(n9707), .ZN(n9721)
         );
  NAND2_X1 U5575 ( .A1(n9721), .A2(n9720), .ZN(n9719) );
  NAND2_X1 U5576 ( .A1(n9736), .A2(n9737), .ZN(n9735) );
  XNOR2_X1 U5577 ( .A(n8438), .B(n9752), .ZN(n9762) );
  NAND2_X1 U5578 ( .A1(n9773), .A2(n9774), .ZN(n9772) );
  AND2_X1 U5579 ( .A1(n4387), .A2(n4762), .ZN(n9817) );
  NAND2_X1 U5580 ( .A1(n9827), .A2(n9828), .ZN(n9826) );
  NAND2_X1 U5581 ( .A1(n9824), .A2(n8465), .ZN(n9841) );
  NAND2_X1 U5582 ( .A1(n9843), .A2(n8498), .ZN(n9863) );
  NAND2_X1 U5583 ( .A1(n9863), .A2(n9864), .ZN(n9862) );
  NOR2_X1 U5584 ( .A1(n8522), .A2(n8502), .ZN(n8503) );
  NAND2_X1 U5585 ( .A1(n6294), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5862) );
  NAND2_X1 U5586 ( .A1(n4710), .A2(n4383), .ZN(n4709) );
  NAND2_X1 U5587 ( .A1(n6154), .A2(n6153), .ZN(n6168) );
  OR2_X1 U5588 ( .A1(n6145), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6155) );
  OR2_X1 U5589 ( .A1(n6120), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U5590 ( .A1(n6110), .A2(n10124), .ZN(n6120) );
  INV_X1 U5591 ( .A(n6111), .ZN(n6110) );
  OR2_X1 U5592 ( .A1(n6100), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U5593 ( .A1(n6035), .A2(n10129), .ZN(n6048) );
  NAND2_X1 U5594 ( .A1(n6021), .A2(n6020), .ZN(n6036) );
  INV_X1 U5595 ( .A(n6022), .ZN(n6021) );
  OR2_X1 U5596 ( .A1(n6010), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6022) );
  NAND2_X1 U5597 ( .A1(n8238), .A2(n4702), .ZN(n7418) );
  NAND2_X1 U5598 ( .A1(n7390), .A2(n8224), .ZN(n4702) );
  INV_X1 U5599 ( .A(n8356), .ZN(n7926) );
  INV_X1 U5600 ( .A(n5984), .ZN(n5983) );
  OR2_X1 U5601 ( .A1(n7504), .A2(n7503), .ZN(n8354) );
  OR2_X1 U5602 ( .A1(n5971), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5984) );
  AND4_X1 U5603 ( .A1(n5961), .A2(n5960), .A3(n5959), .A4(n5958), .ZN(n7435)
         );
  INV_X1 U5604 ( .A(n8403), .ZN(n8059) );
  INV_X1 U5605 ( .A(n7290), .ZN(n4470) );
  AND2_X1 U5606 ( .A1(n8216), .A2(n8214), .ZN(n8348) );
  NAND2_X1 U5607 ( .A1(n4740), .A2(n4400), .ZN(n9877) );
  INV_X1 U5608 ( .A(n9881), .ZN(n9894) );
  NOR2_X1 U5609 ( .A1(n6465), .A2(n4611), .ZN(n4610) );
  NAND2_X1 U5610 ( .A1(n5876), .A2(n8183), .ZN(n8343) );
  NAND2_X1 U5611 ( .A1(n8343), .A2(n7990), .ZN(n9898) );
  OAI211_X1 U5612 ( .C1(n6829), .C2(n6828), .A(n6827), .B(n6826), .ZN(n6831)
         );
  XNOR2_X1 U5613 ( .A(n8544), .B(n8543), .ZN(n4757) );
  NOR2_X1 U5614 ( .A1(n8555), .A2(n8302), .ZN(n4712) );
  INV_X1 U5615 ( .A(n8566), .ZN(n8564) );
  AND2_X1 U5616 ( .A1(n6133), .A2(n6132), .ZN(n8604) );
  AND2_X1 U5617 ( .A1(n8282), .A2(n8285), .ZN(n8627) );
  INV_X1 U5618 ( .A(n8341), .ZN(n8639) );
  INV_X1 U5619 ( .A(n4738), .ZN(n4729) );
  NAND2_X1 U5620 ( .A1(n4735), .A2(n4738), .ZN(n4730) );
  AOI21_X1 U5621 ( .B1(n4735), .B2(n4734), .A(n4733), .ZN(n4732) );
  AOI21_X1 U5622 ( .B1(n8676), .B2(n6072), .A(n4468), .ZN(n8664) );
  INV_X1 U5623 ( .A(n8266), .ZN(n4468) );
  NAND2_X1 U5624 ( .A1(n4704), .A2(n4389), .ZN(n4703) );
  AND2_X1 U5625 ( .A1(n4707), .A2(n6028), .ZN(n4706) );
  AND2_X1 U5626 ( .A1(n5969), .A2(n5968), .ZN(n9950) );
  INV_X1 U5627 ( .A(n9955), .ZN(n9967) );
  OR3_X1 U5628 ( .A1(n8516), .A2(n6323), .A3(n8315), .ZN(n6821) );
  AND3_X1 U5629 ( .A1(n6389), .A2(n6825), .A3(n6326), .ZN(n6408) );
  NOR2_X1 U5630 ( .A1(n6322), .A2(n6394), .ZN(n6403) );
  OR2_X1 U5631 ( .A1(n5853), .A2(n6059), .ZN(n5854) );
  AND2_X1 U5632 ( .A1(n6295), .A2(n6294), .ZN(n6296) );
  OAI21_X1 U5633 ( .B1(n6285), .B2(P2_IR_REG_23__SCAN_IN), .A(n4362), .ZN(
        n6289) );
  NAND2_X1 U5634 ( .A1(n6312), .A2(n6059), .ZN(n4480) );
  INV_X1 U5635 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6288) );
  XNOR2_X1 U5636 ( .A(n6313), .B(n6312), .ZN(n6420) );
  NAND2_X1 U5637 ( .A1(n6285), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6313) );
  XNOR2_X1 U5638 ( .A(n6270), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8180) );
  NOR2_X1 U5639 ( .A1(n6058), .A2(n6057), .ZN(n6062) );
  NAND2_X1 U5640 ( .A1(n5838), .A2(n5839), .ZN(n5920) );
  CLKBUF_X1 U5641 ( .A(n5155), .Z(n6343) );
  AND2_X1 U5642 ( .A1(n5168), .A2(n5167), .ZN(n5177) );
  INV_X1 U5643 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U5644 ( .A1(n6873), .A2(n6874), .ZN(n6875) );
  OR2_X1 U5645 ( .A1(n5676), .A2(n5675), .ZN(n5701) );
  CLKBUF_X1 U5646 ( .A(n6871), .Z(n6872) );
  INV_X1 U5647 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5466) );
  AND2_X1 U5648 ( .A1(n5202), .A2(n5204), .ZN(n6851) );
  OR2_X1 U5649 ( .A1(n5201), .A2(n5200), .ZN(n5202) );
  NAND2_X1 U5650 ( .A1(n5107), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n5586) );
  INV_X1 U5651 ( .A(n5566), .ZN(n5107) );
  XNOR2_X1 U5652 ( .A(n5268), .B(n5222), .ZN(n6877) );
  NAND2_X1 U5653 ( .A1(n7801), .A2(n7815), .ZN(n6522) );
  INV_X1 U5654 ( .A(n6522), .ZN(n7803) );
  INV_X1 U5655 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5133) );
  NOR2_X1 U5656 ( .A1(n9193), .A2(n9207), .ZN(n9192) );
  NAND2_X1 U5657 ( .A1(n9265), .A2(n4678), .ZN(n9225) );
  NAND2_X1 U5658 ( .A1(n9239), .A2(n4804), .ZN(n9223) );
  AND2_X1 U5659 ( .A1(n9224), .A2(n7880), .ZN(n4804) );
  NAND2_X1 U5660 ( .A1(n7878), .A2(n4805), .ZN(n9239) );
  NOR2_X1 U5661 ( .A1(n9236), .A2(n4806), .ZN(n4805) );
  INV_X1 U5662 ( .A(n7877), .ZN(n4806) );
  NAND2_X1 U5663 ( .A1(n7878), .A2(n7877), .ZN(n9237) );
  AND2_X1 U5664 ( .A1(n5707), .A2(n5706), .ZN(n9258) );
  NAND2_X1 U5665 ( .A1(n9265), .A2(n9507), .ZN(n9254) );
  NAND2_X1 U5666 ( .A1(n5084), .A2(n5083), .ZN(n9266) );
  OAI21_X1 U5667 ( .B1(n9310), .B2(n7643), .A(n4783), .ZN(n7873) );
  AND2_X1 U5668 ( .A1(n4784), .A2(n9279), .ZN(n4783) );
  OR2_X1 U5669 ( .A1(n4786), .A2(n7643), .ZN(n4784) );
  NAND2_X1 U5670 ( .A1(n9334), .A2(n4365), .ZN(n9281) );
  NAND2_X1 U5671 ( .A1(n9334), .A2(n4685), .ZN(n9295) );
  NOR2_X1 U5672 ( .A1(n4785), .A2(n7706), .ZN(n9294) );
  INV_X1 U5673 ( .A(n9310), .ZN(n4785) );
  NAND2_X1 U5674 ( .A1(n9326), .A2(n7640), .ZN(n9312) );
  AND3_X1 U5675 ( .A1(n5590), .A2(n5589), .A3(n5588), .ZN(n9357) );
  NAND2_X1 U5676 ( .A1(n4447), .A2(n7626), .ZN(n9359) );
  INV_X1 U5677 ( .A(n9355), .ZN(n4447) );
  OAI21_X1 U5678 ( .B1(n7332), .B2(n4873), .A(n4413), .ZN(n7471) );
  OR2_X1 U5679 ( .A1(n7468), .A2(n4874), .ZN(n4873) );
  INV_X1 U5680 ( .A(n7445), .ZN(n4874) );
  AOI21_X1 U5681 ( .B1(n4800), .B2(n7683), .A(n4798), .ZN(n4797) );
  AND2_X1 U5682 ( .A1(n7698), .A2(n7688), .ZN(n7625) );
  NAND2_X1 U5683 ( .A1(n4802), .A2(n7693), .ZN(n7454) );
  NOR2_X2 U5684 ( .A1(n7453), .A2(n4801), .ZN(n4800) );
  NAND2_X1 U5685 ( .A1(n7452), .A2(n7451), .ZN(n4802) );
  AND4_X1 U5686 ( .A1(n5544), .A2(n5543), .A3(n5542), .A4(n5541), .ZN(n9356)
         );
  AND2_X1 U5687 ( .A1(n7448), .A2(n9027), .ZN(n7463) );
  NOR2_X1 U5688 ( .A1(n7336), .A2(n7444), .ZN(n7448) );
  NAND2_X1 U5689 ( .A1(n7117), .A2(n4366), .ZN(n7204) );
  OR2_X1 U5690 ( .A1(n7204), .A2(n9676), .ZN(n7336) );
  NAND2_X1 U5691 ( .A1(n4793), .A2(n4791), .ZN(n7198) );
  AND2_X1 U5692 ( .A1(n4792), .A2(n7188), .ZN(n4791) );
  AND4_X1 U5693 ( .A1(n5393), .A2(n5392), .A3(n5391), .A4(n5390), .ZN(n9592)
         );
  NAND2_X1 U5694 ( .A1(n4796), .A2(n4795), .ZN(n7186) );
  NAND2_X1 U5695 ( .A1(n7117), .A2(n7116), .ZN(n7115) );
  INV_X1 U5696 ( .A(n7615), .ZN(n7111) );
  NAND2_X1 U5697 ( .A1(n5314), .A2(n5313), .ZN(n7031) );
  OR2_X1 U5698 ( .A1(n6863), .A2(n6783), .ZN(n6936) );
  NAND2_X1 U5699 ( .A1(n6860), .A2(n6698), .ZN(n6700) );
  AND4_X1 U5700 ( .A1(n5322), .A2(n5321), .A3(n5320), .A4(n5319), .ZN(n7038)
         );
  NOR2_X1 U5701 ( .A1(n6840), .A2(n6788), .ZN(n6864) );
  AND2_X1 U5702 ( .A1(n6714), .A2(n7763), .ZN(n6789) );
  NOR2_X1 U5703 ( .A1(n6713), .A2(n4660), .ZN(n4659) );
  OR2_X1 U5704 ( .A1(n6842), .A2(n9623), .ZN(n6840) );
  NAND2_X1 U5705 ( .A1(n6694), .A2(n6693), .ZN(n6837) );
  NAND2_X1 U5706 ( .A1(n6629), .A2(n6628), .ZN(n6632) );
  OR2_X1 U5707 ( .A1(n6633), .A2(n4354), .ZN(n6842) );
  AND2_X1 U5708 ( .A1(n9163), .A2(n9162), .ZN(n9368) );
  AND2_X1 U5709 ( .A1(n5827), .A2(n5826), .ZN(n9381) );
  NAND2_X1 U5710 ( .A1(n5741), .A2(n5740), .ZN(n9209) );
  AND2_X1 U5711 ( .A1(n5121), .A2(n5120), .ZN(n9417) );
  NAND2_X1 U5712 ( .A1(n5604), .A2(n5603), .ZN(n9453) );
  NAND2_X1 U5713 ( .A1(n5536), .A2(n5535), .ZN(n9468) );
  INV_X1 U5714 ( .A(n9348), .ZN(n9603) );
  INV_X1 U5715 ( .A(n7381), .ZN(n9676) );
  AND4_X1 U5716 ( .A1(n5369), .A2(n5368), .A3(n5367), .A4(n5366), .ZN(n9655)
         );
  AND2_X1 U5717 ( .A1(n6930), .A2(n9634), .ZN(n9627) );
  NAND2_X1 U5718 ( .A1(n5788), .A2(n9520), .ZN(n6668) );
  XNOR2_X1 U5719 ( .A(n6188), .B(n6187), .ZN(n7528) );
  AND2_X1 U5720 ( .A1(n4374), .A2(n4880), .ZN(n4879) );
  INV_X1 U5721 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n4880) );
  NAND2_X1 U5722 ( .A1(n5802), .A2(n5125), .ZN(n5805) );
  OR2_X1 U5723 ( .A1(n5124), .A2(n5123), .ZN(n5125) );
  NAND2_X1 U5724 ( .A1(n4977), .A2(n5037), .ZN(n5405) );
  NAND2_X1 U5725 ( .A1(n5033), .A2(n4982), .ZN(n4977) );
  XNOR2_X1 U5726 ( .A(n5021), .B(n5020), .ZN(n5310) );
  NAND2_X1 U5727 ( .A1(n5017), .A2(n5016), .ZN(n5284) );
  XNOR2_X1 U5728 ( .A(n4995), .B(n4992), .ZN(n5143) );
  NAND2_X1 U5729 ( .A1(n4485), .A2(n4486), .ZN(n6381) );
  NAND2_X1 U5730 ( .A1(n4903), .A2(n4904), .ZN(n8022) );
  AND2_X1 U5731 ( .A1(n4496), .A2(n4495), .ZN(n6944) );
  INV_X1 U5732 ( .A(n4499), .ZN(n4496) );
  NAND2_X1 U5733 ( .A1(n4495), .A2(n4505), .ZN(n6945) );
  OAI21_X1 U5734 ( .B1(n8082), .B2(n4535), .A(n4534), .ZN(n8046) );
  NOR2_X1 U5735 ( .A1(n4899), .A2(n7967), .ZN(n4892) );
  NAND2_X1 U5736 ( .A1(n4896), .A2(n4894), .ZN(n4893) );
  OAI21_X1 U5737 ( .B1(n7967), .B2(n4378), .A(n4898), .ZN(n4896) );
  NAND2_X1 U5738 ( .A1(n4895), .A2(n4899), .ZN(n4894) );
  NAND2_X1 U5739 ( .A1(n7967), .A2(n4378), .ZN(n4897) );
  AND2_X1 U5740 ( .A1(n7317), .A2(n7318), .ZN(n4883) );
  AND4_X1 U5741 ( .A1(n6116), .A2(n6115), .A3(n6114), .A4(n6113), .ZN(n8642)
         );
  NAND2_X1 U5742 ( .A1(n4906), .A2(n4910), .ZN(n8052) );
  NAND2_X1 U5743 ( .A1(n8046), .A2(n4911), .ZN(n4906) );
  NAND2_X1 U5744 ( .A1(n7958), .A2(n7957), .ZN(n8071) );
  NAND2_X1 U5745 ( .A1(n6152), .A2(n6151), .ZN(n8076) );
  AOI21_X1 U5746 ( .B1(n8082), .B2(n8079), .A(n8080), .ZN(n8089) );
  AND3_X1 U5747 ( .A1(n6142), .A2(n6141), .A3(n6140), .ZN(n8590) );
  NAND2_X1 U5748 ( .A1(n6144), .A2(n6143), .ZN(n8101) );
  NAND2_X1 U5749 ( .A1(n7024), .A2(n7023), .ZN(n7022) );
  NAND2_X1 U5750 ( .A1(n4500), .A2(n4497), .ZN(n7024) );
  NAND2_X1 U5751 ( .A1(n4499), .A2(n4498), .ZN(n4497) );
  NAND2_X1 U5752 ( .A1(n4502), .A2(n4501), .ZN(n4500) );
  INV_X1 U5753 ( .A(n4504), .ZN(n4498) );
  NAND2_X1 U5754 ( .A1(n4528), .A2(n4526), .ZN(n7923) );
  AOI21_X1 U5755 ( .B1(n8046), .B2(n8045), .A(n4358), .ZN(n8104) );
  AOI21_X1 U5756 ( .B1(n8082), .B2(n4532), .A(n4530), .ZN(n4529) );
  XNOR2_X1 U5757 ( .A(n6374), .B(n7991), .ZN(n6736) );
  NAND2_X1 U5758 ( .A1(n4538), .A2(n4540), .ZN(n8145) );
  NAND2_X1 U5759 ( .A1(n8082), .A2(n4539), .ZN(n4538) );
  INV_X1 U5760 ( .A(n8172), .ZN(n8157) );
  AND2_X1 U5761 ( .A1(n4491), .A2(n4493), .ZN(n7156) );
  NAND2_X1 U5762 ( .A1(n4491), .A2(n4489), .ZN(n7154) );
  NAND2_X1 U5763 ( .A1(n4903), .A2(n4394), .ZN(n8166) );
  AND2_X1 U5764 ( .A1(n4903), .A2(n4902), .ZN(n8168) );
  INV_X1 U5765 ( .A(n8149), .ZN(n8175) );
  INV_X1 U5766 ( .A(n8380), .ZN(n8536) );
  INV_X1 U5767 ( .A(n8604), .ZN(n8619) );
  INV_X1 U5768 ( .A(n8125), .ZN(n8631) );
  INV_X1 U5769 ( .A(n7435), .ZN(n8405) );
  INV_X1 U5770 ( .A(n7318), .ZN(n8406) );
  OR2_X1 U5771 ( .A1(n6419), .A2(n6362), .ZN(n8408) );
  NAND2_X1 U5772 ( .A1(n6983), .A2(n4778), .ZN(n6912) );
  NOR2_X1 U5773 ( .A1(n6994), .A2(n6995), .ZN(n7134) );
  NAND2_X1 U5774 ( .A1(n4617), .A2(n8434), .ZN(n7227) );
  INV_X1 U5775 ( .A(n4620), .ZN(n9744) );
  INV_X1 U5776 ( .A(n4452), .ZN(n9780) );
  INV_X1 U5777 ( .A(n4762), .ZN(n9799) );
  INV_X1 U5778 ( .A(n4773), .ZN(n9832) );
  INV_X1 U5779 ( .A(n4630), .ZN(n9851) );
  INV_X1 U5780 ( .A(n4628), .ZN(n9849) );
  NAND2_X1 U5781 ( .A1(n6430), .A2(n6429), .ZN(n9858) );
  INV_X1 U5782 ( .A(n4768), .ZN(n9869) );
  NAND2_X1 U5783 ( .A1(n6209), .A2(n6208), .ZN(n8311) );
  AND2_X1 U5784 ( .A1(n4696), .A2(n4694), .ZN(n8010) );
  AOI21_X1 U5785 ( .B1(n6284), .B2(n9883), .A(n4695), .ZN(n4694) );
  OR2_X1 U5786 ( .A1(n8006), .A2(n7992), .ZN(n4696) );
  INV_X1 U5787 ( .A(n6283), .ZN(n4695) );
  NAND2_X1 U5788 ( .A1(n6099), .A2(n6098), .ZN(n8744) );
  AND2_X1 U5789 ( .A1(n8710), .A2(n6969), .ZN(n9888) );
  NAND2_X1 U5790 ( .A1(n9895), .A2(n6227), .ZN(n6965) );
  INV_X1 U5791 ( .A(n8706), .ZN(n9905) );
  NAND2_X1 U5792 ( .A1(n8319), .A2(n8318), .ZN(n8769) );
  NAND2_X1 U5793 ( .A1(n8010), .A2(n4692), .ZN(n6332) );
  NAND2_X1 U5794 ( .A1(n4697), .A2(n4693), .ZN(n4692) );
  INV_X1 U5795 ( .A(n8006), .ZN(n4697) );
  NAND2_X1 U5796 ( .A1(n4743), .A2(n4747), .ZN(n8556) );
  NAND2_X1 U5797 ( .A1(n6175), .A2(n8297), .ZN(n8554) );
  NAND2_X1 U5798 ( .A1(n6165), .A2(n6164), .ZN(n8786) );
  NAND2_X1 U5799 ( .A1(n8575), .A2(n6261), .ZN(n8567) );
  INV_X1 U5800 ( .A(n8076), .ZN(n8791) );
  AND2_X1 U5801 ( .A1(n6136), .A2(n6135), .ZN(n8802) );
  NAND2_X1 U5802 ( .A1(n6128), .A2(n6127), .ZN(n8129) );
  NAND2_X1 U5803 ( .A1(n6119), .A2(n6118), .ZN(n8808) );
  NAND2_X1 U5804 ( .A1(n6108), .A2(n6107), .ZN(n8814) );
  NAND2_X1 U5805 ( .A1(n6085), .A2(n6084), .ZN(n8825) );
  NAND2_X1 U5806 ( .A1(n4731), .A2(n4735), .ZN(n8665) );
  NAND2_X1 U5807 ( .A1(n8690), .A2(n4736), .ZN(n4731) );
  AOI21_X1 U5808 ( .B1(n8690), .B2(n6250), .A(n4739), .ZN(n8679) );
  NAND2_X1 U5809 ( .A1(n4714), .A2(n4721), .ZN(n7530) );
  NAND2_X1 U5810 ( .A1(n7421), .A2(n4723), .ZN(n4714) );
  NAND2_X1 U5811 ( .A1(n7483), .A2(n8245), .ZN(n7534) );
  NAND2_X1 U5812 ( .A1(n4725), .A2(n4723), .ZN(n7479) );
  NAND2_X1 U5813 ( .A1(n6006), .A2(n8239), .ZN(n7485) );
  NOR2_X1 U5814 ( .A1(n9970), .A2(n9962), .ZN(n8851) );
  AND2_X1 U5815 ( .A1(n6420), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6721) );
  INV_X1 U5816 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5851) );
  BUF_X1 U5817 ( .A(n5855), .Z(n8013) );
  INV_X1 U5818 ( .A(n6296), .ZN(n7524) );
  XNOR2_X1 U5819 ( .A(n6287), .B(n6286), .ZN(n7518) );
  INV_X1 U5820 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U5821 ( .A1(n6291), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U5822 ( .A1(n6291), .A2(n6290), .ZN(n7476) );
  OR2_X1 U5823 ( .A1(n6289), .A2(n6288), .ZN(n6290) );
  INV_X1 U5824 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7315) );
  INV_X1 U5825 ( .A(n8180), .ZN(n7180) );
  NAND2_X1 U5826 ( .A1(n6218), .A2(n6269), .ZN(n8324) );
  INV_X1 U5827 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7071) );
  INV_X1 U5828 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6849) );
  INV_X1 U5829 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6533) );
  AND3_X1 U5830 ( .A1(n4890), .A2(n5839), .A3(n4888), .ZN(n5978) );
  INV_X1 U5831 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6502) );
  INV_X1 U5832 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6472) );
  INV_X1 U5833 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6462) );
  NAND2_X1 U5834 ( .A1(n6059), .A2(n4623), .ZN(n4622) );
  NAND2_X1 U5835 ( .A1(n5863), .A2(n4780), .ZN(n6896) );
  AOI22_X1 U5836 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4398), .B1(n6059), .B2(
        n4781), .ZN(n4780) );
  INV_X1 U5837 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4781) );
  NAND2_X1 U5838 ( .A1(n8862), .A2(n4832), .ZN(n8864) );
  NAND2_X1 U5839 ( .A1(n5509), .A2(n5511), .ZN(n4834) );
  AND2_X1 U5840 ( .A1(n4825), .A2(n8983), .ZN(n8876) );
  NAND2_X1 U5841 ( .A1(n5384), .A2(n5383), .ZN(n9658) );
  INV_X1 U5842 ( .A(n4837), .ZN(n4836) );
  NAND2_X1 U5843 ( .A1(n5353), .A2(n5349), .ZN(n6956) );
  NAND2_X1 U5844 ( .A1(n5152), .A2(n5153), .ZN(n4548) );
  AND2_X1 U5845 ( .A1(n5632), .A2(n5631), .ZN(n9316) );
  NAND2_X1 U5846 ( .A1(n4816), .A2(n4814), .ZN(n8907) );
  AND2_X1 U5847 ( .A1(n4816), .A2(n4818), .ZN(n8908) );
  NAND2_X1 U5848 ( .A1(n4817), .A2(n4819), .ZN(n4816) );
  OR2_X1 U5849 ( .A1(n4369), .A2(n8916), .ZN(n4560) );
  AND4_X1 U5850 ( .A1(n5525), .A2(n5524), .A3(n5523), .A4(n5522), .ZN(n8934)
         );
  OAI21_X1 U5851 ( .B1(n8923), .B2(n5554), .A(n5553), .ZN(n5559) );
  NAND2_X1 U5852 ( .A1(n5564), .A2(n5563), .ZN(n9463) );
  AND2_X1 U5853 ( .A1(n4820), .A2(n4824), .ZN(n8953) );
  NAND2_X1 U5854 ( .A1(n4563), .A2(n4821), .ZN(n8951) );
  NAND2_X1 U5855 ( .A1(n5698), .A2(n5697), .ZN(n9243) );
  CLKBUF_X1 U5856 ( .A(n7011), .Z(n7012) );
  AND3_X1 U5857 ( .A1(n5611), .A2(n5610), .A3(n5609), .ZN(n9330) );
  INV_X1 U5858 ( .A(n9266), .ZN(n9426) );
  AND2_X1 U5859 ( .A1(n5653), .A2(n5652), .ZN(n9301) );
  AND4_X1 U5860 ( .A1(n5446), .A2(n5445), .A3(n5444), .A4(n5443), .ZN(n9673)
         );
  AND4_X1 U5861 ( .A1(n5571), .A2(n5570), .A3(n5569), .A4(n5568), .ZN(n9329)
         );
  NAND2_X1 U5862 ( .A1(n4399), .A2(n5598), .ZN(n8993) );
  AND2_X1 U5863 ( .A1(n5598), .A2(n5596), .ZN(n8994) );
  AND2_X1 U5864 ( .A1(n5730), .A2(n5729), .ZN(n9390) );
  AND2_X1 U5865 ( .A1(n5820), .A2(n5743), .ZN(n9210) );
  NAND2_X1 U5866 ( .A1(n5814), .A2(n7819), .ZN(n9022) );
  AND2_X1 U5867 ( .A1(n5809), .A2(n5807), .ZN(n9016) );
  NOR2_X1 U5868 ( .A1(n7636), .A2(n4960), .ZN(n4959) );
  AOI21_X1 U5869 ( .B1(n7802), .B2(n7801), .A(n7819), .ZN(n4957) );
  OR2_X1 U5870 ( .A1(n5169), .A2(n6363), .ZN(n7807) );
  INV_X1 U5871 ( .A(n9390), .ZN(n9211) );
  INV_X1 U5872 ( .A(n9258), .ZN(n9414) );
  INV_X1 U5873 ( .A(n9417), .ZN(n9433) );
  INV_X1 U5874 ( .A(n9316), .ZN(n9432) );
  INV_X1 U5875 ( .A(n9330), .ZN(n9440) );
  INV_X1 U5876 ( .A(n9357), .ZN(n9313) );
  INV_X1 U5877 ( .A(n9329), .ZN(n9030) );
  INV_X1 U5878 ( .A(n9356), .ZN(n9031) );
  INV_X1 U5879 ( .A(n8934), .ZN(n9032) );
  INV_X1 U5880 ( .A(n9592), .ZN(n9037) );
  INV_X1 U5881 ( .A(n9655), .ZN(n9038) );
  INV_X1 U5882 ( .A(n7038), .ZN(n9039) );
  BUF_X1 U5883 ( .A(n5154), .Z(n9044) );
  AND2_X1 U5884 ( .A1(n7835), .A2(n7834), .ZN(n9149) );
  XNOR2_X1 U5885 ( .A(n4688), .B(n9482), .ZN(n9365) );
  NAND2_X1 U5886 ( .A1(n4689), .A2(n4650), .ZN(n4688) );
  NOR2_X1 U5887 ( .A1(n9168), .A2(n9348), .ZN(n9369) );
  AOI21_X1 U5888 ( .B1(n4789), .B2(n7727), .A(n7738), .ZN(n4788) );
  INV_X1 U5889 ( .A(n4862), .ZN(n4861) );
  OAI21_X1 U5890 ( .B1(n4865), .B2(n4867), .A(n4864), .ZN(n4862) );
  AND2_X1 U5891 ( .A1(n7869), .A2(n4867), .ZN(n9187) );
  INV_X1 U5892 ( .A(n9185), .ZN(n4479) );
  AND2_X1 U5893 ( .A1(n5774), .A2(n5773), .ZN(n9391) );
  NAND2_X1 U5894 ( .A1(n9292), .A2(n7871), .ZN(n9280) );
  INV_X1 U5895 ( .A(n9468), .ZN(n8935) );
  NAND2_X1 U5896 ( .A1(n4869), .A2(n7445), .ZN(n7469) );
  NAND2_X1 U5897 ( .A1(n7332), .A2(n4875), .ZN(n4869) );
  NAND2_X1 U5898 ( .A1(n7332), .A2(n7331), .ZN(n7447) );
  AND4_X1 U5899 ( .A1(n5501), .A2(n5500), .A3(n5499), .A4(n5498), .ZN(n9671)
         );
  INV_X1 U5900 ( .A(n9034), .ZN(n8867) );
  AOI21_X1 U5901 ( .B1(n9591), .B2(n9595), .A(n4357), .ZN(n4851) );
  AND4_X1 U5902 ( .A1(n5418), .A2(n5417), .A3(n5416), .A4(n5415), .ZN(n9654)
         );
  AND4_X1 U5903 ( .A1(n5341), .A2(n5340), .A3(n5339), .A4(n5338), .ZN(n7114)
         );
  NAND2_X1 U5904 ( .A1(n6926), .A2(n6925), .ZN(n6928) );
  NOR2_X1 U5905 ( .A1(n4352), .A2(n9680), .ZN(n9307) );
  INV_X1 U5906 ( .A(n6715), .ZN(n7646) );
  NAND2_X1 U5907 ( .A1(n6835), .A2(n6695), .ZN(n6787) );
  NAND2_X1 U5908 ( .A1(n6664), .A2(n6512), .ZN(n7977) );
  INV_X1 U5909 ( .A(n9305), .ZN(n9608) );
  NAND2_X1 U5910 ( .A1(n6712), .A2(n6711), .ZN(n4661) );
  NAND2_X1 U5911 ( .A1(n9342), .A2(n7815), .ZN(n9305) );
  AOI21_X1 U5912 ( .B1(n9365), .B2(n9603), .A(n9368), .ZN(n9479) );
  INV_X1 U5913 ( .A(n9183), .ZN(n9487) );
  NAND2_X1 U5914 ( .A1(n9684), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n4475) );
  INV_X1 U5915 ( .A(n9193), .ZN(n9491) );
  INV_X1 U5916 ( .A(n9209), .ZN(n9495) );
  INV_X1 U5917 ( .A(n9243), .ZN(n9503) );
  OR2_X2 U5918 ( .A1(n6516), .A2(n7807), .ZN(n9621) );
  XNOR2_X1 U5919 ( .A(n7553), .B(n7552), .ZN(n8322) );
  OAI22_X1 U5920 ( .A1(n7589), .A2(n7588), .B1(SI_30_), .B2(n7549), .ZN(n7553)
         );
  INV_X1 U5921 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n7554) );
  XNOR2_X1 U5922 ( .A(n6204), .B(n6203), .ZN(n7901) );
  NAND2_X1 U5923 ( .A1(n4966), .A2(n6189), .ZN(n6204) );
  INV_X1 U5924 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5081) );
  AND2_X1 U5925 ( .A1(n4374), .A2(n4882), .ZN(n4881) );
  AND2_X1 U5926 ( .A1(n5090), .A2(n5093), .ZN(n7492) );
  AOI21_X1 U5927 ( .B1(n4829), .B2(n5408), .A(n4418), .ZN(n4827) );
  INV_X1 U5928 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7313) );
  INV_X1 U5929 ( .A(n5806), .ZN(n7756) );
  INV_X1 U5930 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7567) );
  INV_X1 U5931 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n6847) );
  INV_X1 U5932 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6531) );
  XNOR2_X1 U5933 ( .A(n5310), .B(n5311), .ZN(n6468) );
  OAI21_X1 U5934 ( .B1(n5284), .B2(n5283), .A(n5019), .ZN(n5311) );
  INV_X1 U5935 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U5936 ( .A1(n4948), .A2(n5005), .ZN(n5227) );
  NAND2_X1 U5937 ( .A1(n4511), .A2(n4514), .ZN(n4510) );
  OR2_X1 U5938 ( .A1(n8393), .A2(n8392), .ZN(n4469) );
  AOI21_X1 U5939 ( .B1(n8509), .B2(n9867), .A(n8508), .ZN(n8510) );
  INV_X1 U5940 ( .A(n4767), .ZN(n8449) );
  AOI21_X1 U5941 ( .B1(n8532), .B2(n9867), .A(n8531), .ZN(n8533) );
  XNOR2_X1 U5942 ( .A(n4624), .B(n8519), .ZN(n8534) );
  OAI21_X1 U5943 ( .B1(n8773), .B2(n9984), .A(n4408), .ZN(P2_U3487) );
  INV_X1 U5944 ( .A(n4753), .ZN(n4752) );
  OAI21_X1 U5945 ( .B1(n4351), .B2(n9694), .A(n4807), .ZN(P1_U3551) );
  NOR2_X1 U5946 ( .A1(n4434), .A2(n4808), .ZN(n4807) );
  NOR2_X1 U5947 ( .A1(n9696), .A2(n7897), .ZN(n4808) );
  NAND2_X1 U5948 ( .A1(n4476), .A2(n4473), .ZN(P1_U3518) );
  INV_X1 U5949 ( .A(n4474), .ZN(n4473) );
  NAND2_X1 U5950 ( .A1(n9486), .A2(n9685), .ZN(n4476) );
  OAI21_X1 U5951 ( .B1(n9487), .B2(n9515), .A(n4475), .ZN(n4474) );
  INV_X2 U5952 ( .A(n5647), .ZN(n5442) );
  AND2_X1 U5953 ( .A1(n4512), .A2(n4367), .ZN(n4355) );
  AND2_X1 U5954 ( .A1(n4682), .A2(n4681), .ZN(n4356) );
  INV_X1 U5955 ( .A(n6247), .ZN(n4728) );
  INV_X2 U5956 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6059) );
  INV_X1 U5957 ( .A(n4877), .ZN(n5287) );
  NOR2_X1 U5958 ( .A1(n9601), .A2(n9036), .ZN(n4357) );
  AND2_X1 U5959 ( .A1(n7942), .A2(n7943), .ZN(n4358) );
  INV_X1 U5960 ( .A(n7727), .ZN(n7885) );
  AND2_X1 U5961 ( .A1(n9193), .A2(n9391), .ZN(n7727) );
  AND2_X1 U5962 ( .A1(n4611), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4359) );
  INV_X1 U5963 ( .A(n8014), .ZN(n4515) );
  NOR2_X1 U5964 ( .A1(n4375), .A2(n4815), .ZN(n4814) );
  OR2_X1 U5965 ( .A1(n6437), .A2(n6059), .ZN(n4360) );
  NAND2_X1 U5966 ( .A1(n5089), .A2(n4831), .ZN(n4361) );
  AND2_X1 U5967 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4480), .ZN(n4362) );
  NOR2_X1 U5968 ( .A1(n5599), .A2(n4939), .ZN(n4938) );
  INV_X1 U5969 ( .A(n4938), .ZN(n4931) );
  INV_X1 U5970 ( .A(n6992), .ZN(n4779) );
  AND2_X1 U5971 ( .A1(n7933), .A2(n4437), .ZN(n4364) );
  AND2_X1 U5972 ( .A1(n4685), .A2(n4684), .ZN(n4365) );
  AND2_X1 U5973 ( .A1(n7364), .A2(n4356), .ZN(n4366) );
  AND2_X1 U5974 ( .A1(n7741), .A2(n7601), .ZN(n7887) );
  INV_X1 U5975 ( .A(n7887), .ZN(n4651) );
  AND2_X1 U5976 ( .A1(n9468), .A2(n9356), .ZN(n7786) );
  INV_X1 U5977 ( .A(n7786), .ZN(n7688) );
  OR2_X1 U5978 ( .A1(n8014), .A2(n4901), .ZN(n4367) );
  AND2_X1 U5979 ( .A1(n7941), .A2(n8643), .ZN(n4368) );
  AND2_X1 U5980 ( .A1(n4821), .A2(n5714), .ZN(n4369) );
  NOR2_X1 U5981 ( .A1(n6251), .A2(n8090), .ZN(n4370) );
  AND2_X1 U5982 ( .A1(n7921), .A2(n8404), .ZN(n4371) );
  AND2_X1 U5983 ( .A1(n7117), .A2(n4682), .ZN(n4372) );
  OR2_X1 U5984 ( .A1(n7382), .A2(n8405), .ZN(n4373) );
  AND4_X1 U5985 ( .A1(n5933), .A2(n5932), .A3(n5931), .A4(n5930), .ZN(n7436)
         );
  NAND2_X1 U5986 ( .A1(n6671), .A2(n7977), .ZN(n9342) );
  NAND2_X1 U5987 ( .A1(n5411), .A2(n5410), .ZN(n9601) );
  INV_X1 U5988 ( .A(n9601), .ZN(n4681) );
  INV_X2 U5989 ( .A(n5878), .ZN(n6019) );
  AND2_X2 U5990 ( .A1(n8013), .A2(n5857), .ZN(n5899) );
  NOR2_X1 U5991 ( .A1(n5638), .A2(n5637), .ZN(n4375) );
  AND2_X1 U5992 ( .A1(n9265), .A2(n4680), .ZN(n4376) );
  INV_X1 U5993 ( .A(n7795), .ZN(n4454) );
  INV_X1 U5994 ( .A(n4899), .ZN(n4898) );
  OAI22_X1 U5995 ( .A1(n8014), .A2(n4900), .B1(n7966), .B2(n8305), .ZN(n4899)
         );
  NOR2_X1 U5996 ( .A1(n7743), .A2(n4652), .ZN(n4377) );
  AND2_X1 U5997 ( .A1(n4515), .A2(n8154), .ZN(n4378) );
  OR2_X1 U5998 ( .A1(n7743), .A2(n7747), .ZN(n4379) );
  NAND2_X1 U5999 ( .A1(n5098), .A2(n5087), .ZN(n4380) );
  AND2_X1 U6000 ( .A1(n8943), .A2(n8942), .ZN(n4381) );
  INV_X1 U6001 ( .A(n9474), .ZN(n9027) );
  AND2_X1 U6002 ( .A1(n5921), .A2(n5842), .ZN(n4382) );
  AND3_X1 U6003 ( .A1(n5096), .A2(n5799), .A3(n7492), .ZN(n5169) );
  OR2_X1 U6004 ( .A1(n8548), .A2(n8558), .ZN(n4383) );
  INV_X1 U6005 ( .A(n7693), .ZN(n4801) );
  OR2_X1 U6006 ( .A1(n9859), .A2(n8448), .ZN(n4384) );
  INV_X1 U6007 ( .A(n9337), .ZN(n9516) );
  NAND2_X1 U6008 ( .A1(n5584), .A2(n5583), .ZN(n9337) );
  INV_X1 U6009 ( .A(n4814), .ZN(n4813) );
  OR2_X1 U6010 ( .A1(n9823), .A2(n8446), .ZN(n4385) );
  AND2_X1 U6011 ( .A1(n5674), .A2(n5673), .ZN(n9507) );
  INV_X1 U6012 ( .A(n9507), .ZN(n9260) );
  NAND2_X1 U6013 ( .A1(n7592), .A2(n7591), .ZN(n9173) );
  AND4_X1 U6014 ( .A1(n5844), .A2(n6056), .A3(n6055), .A4(n5843), .ZN(n4386)
         );
  OR2_X1 U6015 ( .A1(n9787), .A2(n8442), .ZN(n4387) );
  OR2_X1 U6016 ( .A1(n6281), .A2(n8454), .ZN(n4388) );
  OR2_X1 U6017 ( .A1(n8249), .A2(n8024), .ZN(n4389) );
  NAND2_X1 U6018 ( .A1(n5624), .A2(n5623), .ZN(n9303) );
  AND2_X1 U6019 ( .A1(n8543), .A2(n4712), .ZN(n4390) );
  INV_X1 U6020 ( .A(n7617), .ZN(n4795) );
  OR3_X1 U6021 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_25__SCAN_IN), .A3(
        P2_IR_REG_24__SCAN_IN), .ZN(n4391) );
  AND2_X1 U6022 ( .A1(n7944), .A2(n8642), .ZN(n4392) );
  OR2_X1 U6023 ( .A1(n6255), .A2(n7943), .ZN(n4393) );
  AND2_X1 U6024 ( .A1(n4902), .A2(n8167), .ZN(n4394) );
  NAND2_X1 U6025 ( .A1(n4553), .A2(n4549), .ZN(n8898) );
  NOR2_X1 U6026 ( .A1(n4801), .A2(n7694), .ZN(n4395) );
  INV_X1 U6027 ( .A(n9231), .ZN(n9499) );
  NAND2_X1 U6028 ( .A1(n5722), .A2(n5721), .ZN(n9231) );
  AND2_X1 U6029 ( .A1(n9239), .A2(n7880), .ZN(n4396) );
  INV_X1 U6030 ( .A(n6262), .ZN(n4751) );
  AND3_X1 U6031 ( .A1(n8336), .A2(n8333), .A3(n8324), .ZN(n4397) );
  INV_X1 U6032 ( .A(n4912), .ZN(n4911) );
  NAND2_X1 U6033 ( .A1(n4914), .A2(n4913), .ZN(n4912) );
  AND2_X1 U6034 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n4398) );
  INV_X1 U6035 ( .A(n4934), .ZN(n4933) );
  NAND2_X1 U6036 ( .A1(n4936), .A2(SI_20_), .ZN(n4934) );
  INV_X1 U6037 ( .A(n4544), .ZN(n4539) );
  OR2_X1 U6038 ( .A1(n4546), .A2(n4545), .ZN(n4544) );
  AND2_X1 U6039 ( .A1(n5596), .A2(n8995), .ZN(n4399) );
  AND2_X1 U6040 ( .A1(n4741), .A2(n6229), .ZN(n4400) );
  OR2_X1 U6041 ( .A1(n4515), .A2(n4513), .ZN(n4401) );
  AND2_X1 U6042 ( .A1(n5660), .A2(n5659), .ZN(n4402) );
  INV_X1 U6043 ( .A(n7626), .ZN(n9354) );
  AND2_X1 U6044 ( .A1(n7783), .A2(n7642), .ZN(n7626) );
  AND2_X1 U6045 ( .A1(n5530), .A2(SI_16_), .ZN(n4403) );
  INV_X1 U6046 ( .A(n7870), .ZN(n4866) );
  AND2_X1 U6047 ( .A1(n9183), .A2(n9028), .ZN(n7870) );
  AND2_X1 U6048 ( .A1(n8282), .A2(n8281), .ZN(n4404) );
  AND2_X1 U6049 ( .A1(n8780), .A2(n8305), .ZN(n4405) );
  AND2_X1 U6050 ( .A1(n9377), .A2(n9378), .ZN(n4406) );
  AND2_X1 U6051 ( .A1(n8298), .A2(n8299), .ZN(n8582) );
  AND2_X1 U6052 ( .A1(n5884), .A2(n4622), .ZN(n4407) );
  AND2_X1 U6053 ( .A1(n8724), .A2(n4752), .ZN(n4408) );
  AND2_X1 U6054 ( .A1(n7672), .A2(n7679), .ZN(n4409) );
  AND2_X1 U6055 ( .A1(n6252), .A2(n8643), .ZN(n4410) );
  AND2_X1 U6056 ( .A1(n5021), .A2(SI_7_), .ZN(n4411) );
  OR2_X1 U6057 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n4412) );
  AND2_X1 U6058 ( .A1(n4870), .A2(n7470), .ZN(n4413) );
  AND2_X1 U6059 ( .A1(n4776), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4414) );
  OR2_X1 U6060 ( .A1(n6281), .A2(n6896), .ZN(n4415) );
  NOR2_X1 U6061 ( .A1(n6248), .A2(n8117), .ZN(n4416) );
  NAND2_X1 U6062 ( .A1(n5436), .A2(n5435), .ZN(n7217) );
  NOR2_X1 U6063 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5089) );
  OAI21_X1 U6064 ( .B1(n8368), .B2(n4750), .A(n6263), .ZN(n4749) );
  AND2_X1 U6065 ( .A1(n5849), .A2(n4918), .ZN(n4417) );
  AND2_X1 U6066 ( .A1(n4830), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4418) );
  OR2_X1 U6067 ( .A1(n6887), .A2(n6888), .ZN(n4419) );
  INV_X1 U6068 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n4830) );
  INV_X1 U6069 ( .A(n8253), .ZN(n4717) );
  AND2_X1 U6070 ( .A1(n4486), .A2(n4484), .ZN(n4420) );
  INV_X1 U6071 ( .A(n8916), .ZN(n4562) );
  AND2_X1 U6072 ( .A1(n4916), .A2(n4758), .ZN(n4421) );
  AND2_X1 U6073 ( .A1(n6911), .A2(n4779), .ZN(n4422) );
  NAND2_X1 U6074 ( .A1(n9027), .A2(n9032), .ZN(n7696) );
  INV_X1 U6075 ( .A(n7696), .ZN(n4798) );
  NAND2_X1 U6076 ( .A1(n8843), .A2(n8258), .ZN(n4423) );
  AND2_X1 U6077 ( .A1(n8337), .A2(n8329), .ZN(n4424) );
  AND2_X1 U6078 ( .A1(n4563), .A2(n4369), .ZN(n4425) );
  AND2_X1 U6079 ( .A1(n8352), .A2(n6235), .ZN(n4426) );
  AND2_X1 U6080 ( .A1(n8245), .A2(n8246), .ZN(n8355) );
  AND2_X1 U6081 ( .A1(n7896), .A2(n7895), .ZN(n4427) );
  AND2_X1 U6082 ( .A1(n4562), .A2(n4822), .ZN(n4428) );
  INV_X1 U6083 ( .A(n9224), .ZN(n9222) );
  AND2_X1 U6084 ( .A1(n7602), .A2(n7881), .ZN(n9224) );
  AND2_X1 U6085 ( .A1(n4645), .A2(n4644), .ZN(n4429) );
  AND2_X1 U6086 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(SI_0_), .ZN(n4430) );
  INV_X2 U6087 ( .A(n5215), .ZN(n5160) );
  XNOR2_X1 U6088 ( .A(n5097), .B(P1_IR_REG_21__SCAN_IN), .ZN(n5806) );
  INV_X1 U6089 ( .A(n9718), .ZN(n4769) );
  NAND2_X1 U6090 ( .A1(n5643), .A2(n5642), .ZN(n9287) );
  INV_X1 U6091 ( .A(n9287), .ZN(n4684) );
  INV_X1 U6092 ( .A(n9372), .ZN(n4458) );
  AND2_X1 U6093 ( .A1(n7432), .A2(n6236), .ZN(n7397) );
  INV_X1 U6094 ( .A(n8153), .ZN(n4901) );
  AND2_X1 U6095 ( .A1(n9334), .A2(n4687), .ZN(n4431) );
  NAND2_X1 U6096 ( .A1(n5075), .A2(n4877), .ZN(n5490) );
  INV_X1 U6097 ( .A(n7991), .ZN(n8409) );
  INV_X1 U6098 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6312) );
  INV_X1 U6099 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n4466) );
  INV_X1 U6100 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4701) );
  INV_X1 U6101 ( .A(n7922), .ZN(n4525) );
  INV_X1 U6102 ( .A(n8873), .ZN(n4823) );
  OR2_X1 U6103 ( .A1(n6333), .A2(n8734), .ZN(n4432) );
  OR2_X1 U6104 ( .A1(n6333), .A2(n8801), .ZN(n4433) );
  OR2_X1 U6105 ( .A1(n9453), .A2(n9330), .ZN(n7705) );
  NOR2_X1 U6106 ( .A1(n4459), .A2(n9461), .ZN(n4434) );
  INV_X1 U6107 ( .A(n5080), .ZN(n5533) );
  NAND2_X1 U6108 ( .A1(n7186), .A2(n7674), .ZN(n4435) );
  AND2_X1 U6109 ( .A1(n4901), .A2(n8154), .ZN(n4436) );
  AND2_X1 U6110 ( .A1(n4373), .A2(n7922), .ZN(n4437) );
  INV_X1 U6111 ( .A(n8548), .ZN(n8778) );
  NAND2_X1 U6112 ( .A1(n6195), .A2(n6194), .ZN(n8548) );
  NAND2_X1 U6113 ( .A1(n7932), .A2(n8401), .ZN(n4438) );
  AND2_X1 U6114 ( .A1(n5759), .A2(n5758), .ZN(n5782) );
  AND2_X1 U6115 ( .A1(n6380), .A2(n8407), .ZN(n4439) );
  AND2_X1 U6116 ( .A1(n4905), .A2(n8112), .ZN(n4440) );
  AND2_X1 U6117 ( .A1(n6296), .A2(n4482), .ZN(n4441) );
  NAND2_X1 U6118 ( .A1(n7936), .A2(n8173), .ZN(n4442) );
  INV_X1 U6119 ( .A(n4375), .ZN(n4818) );
  INV_X2 U6120 ( .A(n9970), .ZN(n9968) );
  INV_X1 U6121 ( .A(n9685), .ZN(n9684) );
  NAND2_X1 U6122 ( .A1(n5309), .A2(n6774), .ZN(n6886) );
  INV_X1 U6123 ( .A(n8079), .ZN(n4545) );
  NAND2_X1 U6124 ( .A1(n4835), .A2(n7302), .ZN(n7245) );
  AND2_X1 U6125 ( .A1(n4836), .A2(n5353), .ZN(n4443) );
  INV_X1 U6126 ( .A(n4723), .ZN(n4722) );
  AND2_X1 U6127 ( .A1(n8473), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n4444) );
  NAND2_X1 U6128 ( .A1(n4837), .A2(n5353), .ZN(n7010) );
  INV_X1 U6129 ( .A(n4527), .ZN(n4526) );
  NOR2_X1 U6130 ( .A1(n7383), .A2(n7435), .ZN(n4527) );
  INV_X1 U6131 ( .A(n4503), .ZN(n6735) );
  NAND2_X1 U6132 ( .A1(n4507), .A2(n4506), .ZN(n4503) );
  NAND2_X1 U6133 ( .A1(n7117), .A2(n4356), .ZN(n4683) );
  INV_X1 U6134 ( .A(SI_20_), .ZN(n10126) );
  NOR2_X1 U6135 ( .A1(n7316), .A2(n4883), .ZN(n4445) );
  INV_X1 U6136 ( .A(n4851), .ZN(n7200) );
  NAND2_X1 U6137 ( .A1(n7804), .A2(n7844), .ZN(n7810) );
  NAND2_X1 U6138 ( .A1(n8391), .A2(n8180), .ZN(n8315) );
  AND2_X2 U6139 ( .A1(n6555), .A2(n6554), .ZN(n9696) );
  AND2_X1 U6140 ( .A1(n6387), .A2(n6386), .ZN(n8164) );
  INV_X1 U6141 ( .A(n8415), .ZN(n4766) );
  OR2_X1 U6142 ( .A1(n9906), .A2(n8391), .ZN(n9957) );
  INV_X1 U6143 ( .A(n9957), .ZN(n4693) );
  AND4_X1 U6144 ( .A1(n6224), .A2(n6223), .A3(n6222), .A4(n6221), .ZN(n6687)
         );
  NAND2_X1 U6145 ( .A1(n8469), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4446) );
  INV_X1 U6146 ( .A(n4493), .ZN(n4492) );
  NAND2_X1 U6147 ( .A1(n6379), .A2(n7026), .ZN(n4493) );
  INV_X1 U6148 ( .A(SI_15_), .ZN(n4976) );
  INV_X1 U6149 ( .A(n4777), .ZN(n6983) );
  NAND2_X1 U6150 ( .A1(n5101), .A2(n4380), .ZN(n7801) );
  INV_X1 U6151 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n4482) );
  NAND2_X1 U6152 ( .A1(n9825), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n9824) );
  NAND2_X1 U6153 ( .A1(n7183), .A2(n7617), .ZN(n7185) );
  OAI21_X1 U6154 ( .B1(n7081), .B2(n9641), .A(n7114), .ZN(n7083) );
  INV_X1 U6155 ( .A(n7609), .ZN(n6699) );
  OAI21_X1 U6156 ( .B1(n9291), .B2(n7856), .A(n7855), .ZN(n9278) );
  NAND2_X1 U6157 ( .A1(n5038), .A2(n4430), .ZN(n4994) );
  AND2_X1 U6158 ( .A1(n7645), .A2(n7654), .ZN(n7609) );
  NAND2_X1 U6159 ( .A1(n4878), .A2(n7851), .ZN(n9325) );
  OAI21_X1 U6160 ( .B1(n9278), .B2(n7857), .A(n7858), .ZN(n9264) );
  INV_X1 U6161 ( .A(n4858), .ZN(n4857) );
  NAND2_X1 U6162 ( .A1(n5038), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n4465) );
  OAI21_X2 U6163 ( .B1(n9379), .B2(n9627), .A(n4406), .ZN(n9486) );
  INV_X1 U6164 ( .A(n6630), .ZN(n6631) );
  AOI21_X1 U6165 ( .B1(n8628), .B2(n8614), .A(n8615), .ZN(n8613) );
  OAI22_X1 U6166 ( .A1(n8690), .A2(n4730), .B1(n4732), .B2(n4729), .ZN(n8655)
         );
  OAI21_X1 U6167 ( .B1(n6699), .B2(n4859), .A(n6927), .ZN(n4858) );
  AOI21_X1 U6168 ( .B1(n8544), .B2(n8549), .A(n6266), .ZN(n6268) );
  NOR2_X1 U6169 ( .A1(n8626), .A2(n8627), .ZN(n6257) );
  NAND2_X1 U6170 ( .A1(n6632), .A2(n6631), .ZN(n6694) );
  NAND2_X1 U6171 ( .A1(n5251), .A2(n5015), .ZN(n5017) );
  NAND2_X1 U6172 ( .A1(n4944), .A2(n4941), .ZN(n5251) );
  OAI22_X1 U6173 ( .A1(n9235), .A2(n7864), .B1(n9503), .B2(n9258), .ZN(n9221)
         );
  AND2_X1 U6174 ( .A1(n6923), .A2(n6783), .ZN(n7647) );
  NAND2_X1 U6175 ( .A1(n7850), .A2(n7849), .ZN(n4878) );
  OAI21_X1 U6176 ( .B1(n6836), .B2(n4847), .A(n7606), .ZN(n4843) );
  XNOR2_X2 U6177 ( .A(n5154), .B(n6809), .ZN(n7604) );
  NAND2_X1 U6178 ( .A1(n6694), .A2(n4845), .ZN(n4844) );
  INV_X1 U6179 ( .A(n9264), .ZN(n7859) );
  NAND2_X1 U6180 ( .A1(n4844), .A2(n4842), .ZN(n6786) );
  XNOR2_X2 U6181 ( .A(n9041), .B(n9615), .ZN(n7606) );
  INV_X1 U6182 ( .A(n4843), .ZN(n4842) );
  XNOR2_X1 U6183 ( .A(n8446), .B(n9823), .ZN(n9833) );
  AOI21_X1 U6184 ( .B1(n7752), .B2(n7751), .A(n7815), .ZN(n4962) );
  NAND2_X1 U6185 ( .A1(n5065), .A2(n5064), .ZN(n5667) );
  NAND2_X1 U6186 ( .A1(n5761), .A2(n5760), .ZN(n5763) );
  NOR2_X2 U6187 ( .A1(n5226), .A2(n4947), .ZN(n4946) );
  OAI21_X1 U6188 ( .B1(n7740), .B2(n7738), .A(n4641), .ZN(n4647) );
  INV_X1 U6189 ( .A(n7701), .ZN(n7640) );
  OAI21_X2 U6190 ( .B1(n5484), .B2(n5050), .A(n5049), .ZN(n5514) );
  NOR2_X1 U6191 ( .A1(n4653), .A2(n7874), .ZN(n7722) );
  OAI21_X1 U6192 ( .B1(n7709), .B2(n7710), .A(n7708), .ZN(n4658) );
  NAND2_X1 U6193 ( .A1(n9755), .A2(n8493), .ZN(n9773) );
  OAI21_X1 U6194 ( .B1(n8613), .B2(n7906), .A(n7905), .ZN(n7908) );
  INV_X1 U6195 ( .A(n5005), .ZN(n4947) );
  OAI21_X1 U6196 ( .B1(n5038), .B2(n4466), .A(n4465), .ZN(n5004) );
  AOI21_X2 U6197 ( .B1(n6006), .B2(n4706), .A(n4703), .ZN(n8714) );
  NAND2_X1 U6198 ( .A1(n6163), .A2(n8298), .ZN(n8565) );
  INV_X1 U6199 ( .A(n8688), .ZN(n4471) );
  OAI21_X1 U6200 ( .B1(n8395), .B2(n8394), .A(n4469), .ZN(P2_U3296) );
  NAND2_X4 U6201 ( .A1(n6281), .A2(n7550), .ZN(n8320) );
  AOI21_X2 U6202 ( .B1(n8378), .B2(n8377), .A(n8376), .ZN(n8381) );
  INV_X1 U6203 ( .A(n4759), .ZN(n5859) );
  NAND2_X1 U6204 ( .A1(n8409), .A2(n9904), .ZN(n8192) );
  NOR2_X1 U6205 ( .A1(n8385), .A2(n8386), .ZN(n4580) );
  OR2_X2 U6206 ( .A1(n9191), .A2(n7883), .ZN(n7869) );
  NAND2_X2 U6207 ( .A1(n7033), .A2(n7032), .ZN(n7081) );
  INV_X1 U6208 ( .A(n4800), .ZN(n4799) );
  NAND2_X1 U6209 ( .A1(n9203), .A2(n7885), .ZN(n9176) );
  NAND2_X1 U6210 ( .A1(n4478), .A2(n4477), .ZN(n9380) );
  NAND2_X1 U6211 ( .A1(n9694), .A2(n5824), .ZN(n4477) );
  OR2_X1 U6212 ( .A1(n9486), .A2(n9694), .ZN(n4478) );
  AOI21_X1 U6213 ( .B1(n7869), .B2(n7868), .A(n4479), .ZN(n9186) );
  NAND2_X1 U6214 ( .A1(n5691), .A2(n5690), .ZN(n5693) );
  NAND2_X1 U6215 ( .A1(n4641), .A2(n7738), .ZN(n4640) );
  NAND2_X1 U6216 ( .A1(n4638), .A2(n4643), .ZN(n4635) );
  OAI21_X1 U6217 ( .B1(n4962), .B2(n4959), .A(n6548), .ZN(n4958) );
  NAND2_X1 U6218 ( .A1(n4958), .A2(n4957), .ZN(n4956) );
  NAND2_X1 U6219 ( .A1(n7518), .A2(n4481), .ZN(n4483) );
  NAND2_X1 U6220 ( .A1(n4483), .A2(n4441), .ZN(n6298) );
  INV_X1 U6221 ( .A(n6946), .ZN(n4494) );
  INV_X1 U6222 ( .A(n6736), .ZN(n4502) );
  AND2_X1 U6223 ( .A1(n6375), .A2(n9881), .ZN(n4504) );
  NAND2_X1 U6224 ( .A1(n6720), .A2(n6719), .ZN(n4507) );
  NAND2_X1 U6225 ( .A1(n8156), .A2(n4509), .ZN(n4508) );
  OAI211_X1 U6226 ( .C1(n8156), .C2(n4510), .A(n8018), .B(n4508), .ZN(P2_U3154) );
  INV_X1 U6227 ( .A(n8164), .ZN(n4514) );
  INV_X1 U6228 ( .A(n4529), .ZN(n7947) );
  AND2_X1 U6229 ( .A1(n7940), .A2(n8146), .ZN(n4546) );
  NAND2_X1 U6230 ( .A1(n5157), .A2(n4547), .ZN(n4811) );
  INV_X1 U6231 ( .A(n5158), .ZN(n4547) );
  XNOR2_X1 U6232 ( .A(n4548), .B(n5222), .ZN(n5158) );
  NAND2_X1 U6233 ( .A1(n8941), .A2(n4554), .ZN(n4553) );
  NAND3_X1 U6234 ( .A1(n4826), .A2(n4428), .A3(n4825), .ZN(n4561) );
  NAND3_X1 U6235 ( .A1(n4826), .A2(n4825), .A3(n4822), .ZN(n4563) );
  OAI21_X1 U6236 ( .B1(n8899), .B2(n4813), .A(n4567), .ZN(n5665) );
  NAND2_X1 U6237 ( .A1(n8899), .A2(n4567), .ZN(n4566) );
  NAND2_X1 U6238 ( .A1(n5309), .A2(n4571), .ZN(n4570) );
  NAND2_X1 U6239 ( .A1(n4570), .A2(n4419), .ZN(n5346) );
  INV_X1 U6240 ( .A(n5346), .ZN(n5348) );
  OR2_X2 U6241 ( .A1(n5169), .A2(n6702), .ZN(n6337) );
  NAND2_X1 U6242 ( .A1(n8288), .A2(n8329), .ZN(n4579) );
  NAND2_X1 U6243 ( .A1(n4579), .A2(n4576), .ZN(n8289) );
  NAND2_X1 U6244 ( .A1(n4577), .A2(n8315), .ZN(n4576) );
  NAND3_X1 U6245 ( .A1(n8387), .A2(n4584), .A3(n4582), .ZN(n4581) );
  MUX2_X1 U6246 ( .A(n8315), .B(n8188), .S(n5876), .Z(n8189) );
  NAND2_X1 U6247 ( .A1(n7988), .A2(n5876), .ZN(n9890) );
  NAND3_X1 U6248 ( .A1(n4595), .A2(n8225), .A3(n4591), .ZN(n8235) );
  NAND3_X1 U6249 ( .A1(n4597), .A2(n8219), .A3(n4596), .ZN(n4595) );
  NAND3_X1 U6250 ( .A1(n8218), .A2(n8216), .A3(n8217), .ZN(n4597) );
  NAND3_X1 U6251 ( .A1(n4608), .A2(n8355), .A3(n4605), .ZN(n8248) );
  NAND2_X2 U6252 ( .A1(n6452), .A2(n6281), .ZN(n8321) );
  NAND2_X1 U6253 ( .A1(n4415), .A2(n4609), .ZN(n7997) );
  NAND3_X1 U6254 ( .A1(n4613), .A2(n4916), .A3(n4612), .ZN(n6294) );
  NOR2_X1 U6255 ( .A1(n5847), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n4612) );
  INV_X1 U6256 ( .A(n5994), .ZN(n4613) );
  NAND3_X1 U6257 ( .A1(n4617), .A2(n8434), .A3(P2_REG2_REG_7__SCAN_IN), .ZN(
        n4772) );
  INV_X1 U6258 ( .A(n7226), .ZN(n4618) );
  OAI21_X2 U6259 ( .B1(n4360), .B2(n4623), .A(n4407), .ZN(n7062) );
  OAI21_X1 U6260 ( .B1(n7732), .B2(n7737), .A(n4377), .ZN(n4648) );
  NAND3_X1 U6261 ( .A1(n4637), .A2(n4636), .A3(n4635), .ZN(n7744) );
  NAND3_X1 U6262 ( .A1(n7740), .A2(n4643), .A3(n4641), .ZN(n4636) );
  NAND3_X1 U6263 ( .A1(n7732), .A2(n4377), .A3(n4643), .ZN(n4637) );
  NAND3_X1 U6264 ( .A1(n4640), .A2(n4429), .A3(n4639), .ZN(n4638) );
  NAND3_X1 U6265 ( .A1(n4647), .A2(n4648), .A3(n4645), .ZN(n7746) );
  INV_X1 U6266 ( .A(n9173), .ZN(n4650) );
  NAND2_X1 U6267 ( .A1(n6712), .A2(n4659), .ZN(n6714) );
  XNOR2_X1 U6268 ( .A(n7608), .B(n4661), .ZN(n6839) );
  NAND4_X2 U6269 ( .A1(n4838), .A2(n4877), .A3(n4673), .A4(n4374), .ZN(n7557)
         );
  XNOR2_X2 U6270 ( .A(n4674), .B(n5082), .ZN(n7891) );
  NAND2_X1 U6271 ( .A1(n5080), .A2(n4881), .ZN(n4675) );
  INV_X1 U6272 ( .A(n4683), .ZN(n9602) );
  NOR2_X2 U6273 ( .A1(n9177), .A2(n7982), .ZN(n4689) );
  NAND3_X1 U6274 ( .A1(n4922), .A2(n4691), .A3(n4690), .ZN(n4921) );
  AOI21_X2 U6275 ( .B1(n6175), .B2(n4390), .A(n4709), .ZN(n8378) );
  NAND2_X1 U6276 ( .A1(n5937), .A2(n4713), .ZN(n5962) );
  MUX2_X1 U6277 ( .A(n6059), .B(n5935), .S(P2_IR_REG_6__SCAN_IN), .Z(n5936) );
  NAND2_X1 U6278 ( .A1(n7421), .A2(n4719), .ZN(n4718) );
  NAND3_X1 U6279 ( .A1(n6226), .A2(n8345), .A3(n6228), .ZN(n4740) );
  NAND2_X1 U6280 ( .A1(n6226), .A2(n8345), .ZN(n9895) );
  AND4_X2 U6281 ( .A1(n5864), .A2(n5867), .A3(n5865), .A4(n5866), .ZN(n9892)
         );
  OR2_X1 U6282 ( .A1(n5878), .A2(n5858), .ZN(n5866) );
  NAND2_X2 U6283 ( .A1(n8013), .A2(n7824), .ZN(n5878) );
  NAND2_X1 U6284 ( .A1(n8577), .A2(n4748), .ZN(n4743) );
  OAI21_X1 U6285 ( .B1(n8577), .B2(n4746), .A(n4744), .ZN(n6265) );
  INV_X1 U6286 ( .A(n4747), .ZN(n4746) );
  NAND2_X1 U6287 ( .A1(n7296), .A2(n4426), .ZN(n7432) );
  INV_X2 U6288 ( .A(n5884), .ZN(n5839) );
  INV_X1 U6289 ( .A(n4775), .ZN(n4774) );
  AOI21_X1 U6290 ( .B1(n7054), .B2(n6911), .A(n4779), .ZN(n4777) );
  NAND2_X1 U6291 ( .A1(n7054), .A2(n4422), .ZN(n4778) );
  NAND2_X1 U6292 ( .A1(n4782), .A2(n6630), .ZN(n6712) );
  XNOR2_X1 U6293 ( .A(n4782), .B(n6630), .ZN(n6797) );
  NAND2_X1 U6294 ( .A1(n6627), .A2(n6626), .ZN(n4782) );
  NAND2_X1 U6295 ( .A1(n7884), .A2(n4789), .ZN(n4787) );
  NAND2_X1 U6296 ( .A1(n4787), .A2(n4788), .ZN(n7888) );
  NAND2_X1 U6297 ( .A1(n7884), .A2(n7883), .ZN(n9203) );
  NAND2_X1 U6298 ( .A1(n7079), .A2(n4794), .ZN(n4793) );
  INV_X1 U6299 ( .A(n7079), .ZN(n4796) );
  OAI21_X1 U6300 ( .B1(n7452), .B2(n4799), .A(n4797), .ZN(n4803) );
  INV_X1 U6301 ( .A(n4803), .ZN(n7461) );
  OAI21_X1 U6302 ( .B1(n5157), .B2(n5158), .A(n6852), .ZN(n6727) );
  NAND2_X1 U6303 ( .A1(n5158), .A2(n5157), .ZN(n6852) );
  NAND2_X1 U6304 ( .A1(n4811), .A2(n4810), .ZN(n5181) );
  NAND2_X1 U6305 ( .A1(n5158), .A2(n5156), .ZN(n4810) );
  NAND3_X1 U6306 ( .A1(n6359), .A2(n6361), .A3(n6360), .ZN(P1_U3220) );
  INV_X1 U6307 ( .A(n8972), .ZN(n4819) );
  NAND3_X1 U6308 ( .A1(n4825), .A2(n8983), .A3(n8873), .ZN(n4820) );
  NAND2_X1 U6309 ( .A1(n8982), .A2(n8984), .ZN(n4825) );
  INV_X1 U6310 ( .A(n8981), .ZN(n4826) );
  NAND2_X1 U6311 ( .A1(n5098), .A2(n4831), .ZN(n5122) );
  NAND2_X1 U6312 ( .A1(n4828), .A2(n4827), .ZN(n5090) );
  NAND2_X1 U6313 ( .A1(n5098), .A2(n4829), .ZN(n4828) );
  NAND3_X1 U6314 ( .A1(n5509), .A2(n5511), .A3(n8863), .ZN(n8862) );
  NAND2_X1 U6315 ( .A1(n4834), .A2(n4833), .ZN(n4832) );
  INV_X1 U6316 ( .A(n8863), .ZN(n4833) );
  NAND3_X1 U6317 ( .A1(n4835), .A2(n7302), .A3(n5403), .ZN(n7246) );
  NAND2_X1 U6318 ( .A1(n5400), .A2(n5399), .ZN(n7302) );
  NAND2_X1 U6319 ( .A1(n5398), .A2(n5397), .ZN(n4835) );
  NAND2_X1 U6320 ( .A1(n4877), .A2(n4839), .ZN(n5126) );
  NAND3_X1 U6321 ( .A1(n5189), .A2(n5231), .A3(n4841), .ZN(n5285) );
  NOR2_X1 U6322 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n4841) );
  NAND2_X1 U6323 ( .A1(n4848), .A2(n4852), .ZN(n7202) );
  NAND2_X1 U6324 ( .A1(n7185), .A2(n4849), .ZN(n4848) );
  NAND2_X1 U6325 ( .A1(n6860), .A2(n4855), .ZN(n4854) );
  NAND2_X1 U6326 ( .A1(n7869), .A2(n4863), .ZN(n4860) );
  OAI211_X1 U6327 ( .C1(n7869), .C2(n4865), .A(n4861), .B(n4860), .ZN(n7975)
         );
  NAND2_X1 U6328 ( .A1(n8156), .A2(n4892), .ZN(n4891) );
  OAI211_X1 U6329 ( .C1(n8156), .C2(n4897), .A(n4893), .B(n4891), .ZN(n7974)
         );
  NAND2_X1 U6330 ( .A1(n8113), .A2(n4440), .ZN(n4903) );
  NAND2_X2 U6331 ( .A1(n4921), .A2(n4919), .ZN(n4998) );
  NAND3_X1 U6332 ( .A1(n4920), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4919) );
  NAND2_X1 U6333 ( .A1(n5580), .A2(n4926), .ZN(n4925) );
  NAND2_X1 U6334 ( .A1(n4935), .A2(n4936), .ZN(n5622) );
  NAND2_X1 U6335 ( .A1(n4948), .A2(n4946), .ZN(n5229) );
  NAND2_X1 U6336 ( .A1(n5206), .A2(n5205), .ZN(n4948) );
  AOI21_X1 U6337 ( .B1(n4946), .B2(n4943), .A(n4942), .ZN(n4941) );
  INV_X1 U6338 ( .A(n5205), .ZN(n4943) );
  NAND2_X1 U6339 ( .A1(n4945), .A2(n4946), .ZN(n4944) );
  INV_X1 U6340 ( .A(n5206), .ZN(n4945) );
  NAND3_X1 U6341 ( .A1(n7583), .A2(n7584), .A3(n7590), .ZN(n7586) );
  NAND2_X1 U6342 ( .A1(n5716), .A2(n4953), .ZN(n4951) );
  NAND3_X1 U6343 ( .A1(n7817), .A2(n7818), .A3(n4956), .ZN(P1_U3242) );
  NAND2_X1 U6344 ( .A1(n6188), .A2(n4967), .ZN(n4963) );
  NAND2_X1 U6345 ( .A1(n4963), .A2(n4964), .ZN(n7547) );
  NAND2_X1 U6346 ( .A1(n6188), .A2(n6187), .ZN(n4966) );
  NAND2_X1 U6347 ( .A1(n5514), .A2(n4972), .ZN(n4971) );
  OAI21_X2 U6348 ( .B1(n5033), .B2(n4980), .A(n4978), .ZN(n5430) );
  INV_X1 U6349 ( .A(n6366), .ZN(n6825) );
  NAND2_X1 U6350 ( .A1(n6829), .A2(n6366), .ZN(n6394) );
  INV_X1 U6351 ( .A(n8769), .ZN(n8722) );
  NAND2_X1 U6352 ( .A1(n7293), .A2(n6234), .ZN(n7296) );
  OR2_X1 U6353 ( .A1(n6506), .A2(n6309), .ZN(n6391) );
  OR2_X1 U6354 ( .A1(n6506), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U6355 ( .A1(n7986), .A2(n9447), .ZN(n7896) );
  INV_X1 U6356 ( .A(n9001), .ZN(n9006) );
  OAI21_X1 U6357 ( .B1(n9001), .B2(n5782), .A(n5783), .ZN(n5784) );
  NAND2_X1 U6358 ( .A1(n7859), .A2(n4991), .ZN(n7861) );
  NAND2_X1 U6359 ( .A1(n7899), .A2(n7898), .ZN(n7900) );
  OR2_X1 U6360 ( .A1(n6488), .A2(n5182), .ZN(n5188) );
  OR2_X1 U6361 ( .A1(n6488), .A2(n5159), .ZN(n5164) );
  NAND2_X1 U6362 ( .A1(n4351), .A2(n9685), .ZN(n7899) );
  NAND2_X1 U6363 ( .A1(n6289), .A2(n6288), .ZN(n6291) );
  OR2_X1 U6364 ( .A1(n7547), .A2(n7546), .ZN(n7548) );
  CLKBUF_X1 U6365 ( .A(n5994), .Z(n6016) );
  NOR2_X2 U6366 ( .A1(n9004), .A2(n5756), .ZN(n9001) );
  NOR3_X2 U6367 ( .A1(n9001), .A2(n5782), .A3(n5783), .ZN(n6358) );
  AND2_X1 U6368 ( .A1(n8134), .A2(n7924), .ZN(n4988) );
  AND2_X2 U6369 ( .A1(n6827), .A2(n6318), .ZN(n9986) );
  AND2_X1 U6370 ( .A1(n8924), .A2(n5551), .ZN(n4989) );
  AND2_X1 U6371 ( .A1(n5032), .A2(n5031), .ZN(n4990) );
  OR3_X1 U6372 ( .A1(n5828), .A2(n9672), .A3(n6522), .ZN(n8988) );
  OR2_X1 U6373 ( .A1(n9266), .A2(n9433), .ZN(n4991) );
  INV_X1 U6374 ( .A(n5239), .ZN(n5647) );
  INV_X1 U6375 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5845) );
  INV_X1 U6376 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5843) );
  OR2_X1 U6377 ( .A1(n8035), .A2(n8059), .ZN(n7924) );
  INV_X1 U6378 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5850) );
  INV_X1 U6379 ( .A(n7248), .ZN(n5403) );
  INV_X1 U6380 ( .A(n6730), .ZN(n5180) );
  INV_X1 U6381 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5069) );
  INV_X1 U6382 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10124) );
  INV_X1 U6383 ( .A(n6088), .ZN(n6087) );
  NOR2_X1 U6384 ( .A1(n5552), .A2(n4989), .ZN(n5553) );
  INV_X1 U6385 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n5335) );
  INV_X1 U6386 ( .A(SI_26_), .ZN(n10143) );
  INV_X1 U6387 ( .A(SI_13_), .ZN(n10156) );
  INV_X1 U6388 ( .A(SI_9_), .ZN(n10171) );
  INV_X1 U6389 ( .A(n6155), .ZN(n6154) );
  NAND2_X1 U6390 ( .A1(n6087), .A2(n6086), .ZN(n6100) );
  NAND2_X1 U6391 ( .A1(n5983), .A2(n8037), .ZN(n5999) );
  INV_X1 U6392 ( .A(n8324), .ZN(n6323) );
  INV_X1 U6393 ( .A(n6315), .ZN(n6828) );
  OAI21_X1 U6394 ( .B1(n9877), .B2(n6231), .A(n6230), .ZN(n7164) );
  INV_X1 U6395 ( .A(n6829), .ZN(n6389) );
  INV_X1 U6396 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5848) );
  INV_X1 U6397 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U6398 ( .A1(n5108), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5625) );
  INV_X1 U6399 ( .A(n5645), .ZN(n5109) );
  OR2_X1 U6400 ( .A1(n9002), .A2(n9003), .ZN(n5756) );
  AND2_X1 U6401 ( .A1(n7978), .A2(n5821), .ZN(n9178) );
  INV_X1 U6402 ( .A(n7684), .ZN(n7776) );
  INV_X1 U6403 ( .A(n7894), .ZN(n7895) );
  AND2_X1 U6404 ( .A1(n7678), .A2(n7675), .ZN(n7619) );
  INV_X1 U6405 ( .A(n7801), .ZN(n6548) );
  INV_X1 U6406 ( .A(n6473), .ZN(n5804) );
  INV_X1 U6407 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5087) );
  NAND2_X1 U6408 ( .A1(n5053), .A2(n10074), .ZN(n5056) );
  INV_X1 U6409 ( .A(SI_12_), .ZN(n10072) );
  OR2_X1 U6410 ( .A1(n6419), .A2(n6418), .ZN(n6424) );
  OR2_X1 U6411 ( .A1(n5942), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5956) );
  INV_X1 U6412 ( .A(n8402), .ZN(n8063) );
  INV_X1 U6413 ( .A(n8656), .ZN(n7943) );
  AND2_X1 U6414 ( .A1(n6411), .A2(n6410), .ZN(n8170) );
  INV_X1 U6415 ( .A(n8170), .ZN(n8160) );
  INV_X1 U6416 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10095) );
  INV_X1 U6417 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n8037) );
  INV_X1 U6418 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10129) );
  INV_X1 U6419 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10109) );
  INV_X1 U6420 ( .A(n6424), .ZN(n6428) );
  OR2_X1 U6421 ( .A1(n6432), .A2(n7821), .ZN(n6609) );
  OR2_X1 U6422 ( .A1(n6178), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6197) );
  NAND2_X1 U6423 ( .A1(n6129), .A2(n10107), .ZN(n6137) );
  INV_X1 U6424 ( .A(n8667), .ZN(n8643) );
  AND2_X1 U6425 ( .A1(n6391), .A2(n6505), .ZN(n6326) );
  INV_X1 U6426 ( .A(n8398), .ZN(n8579) );
  AND2_X1 U6427 ( .A1(n8281), .A2(n8280), .ZN(n8341) );
  AND2_X1 U6428 ( .A1(n4717), .A2(n8252), .ZN(n8359) );
  NAND2_X1 U6429 ( .A1(n6272), .A2(n6821), .ZN(n7992) );
  AND2_X1 U6430 ( .A1(n8209), .A2(n8213), .ZN(n7166) );
  INV_X1 U6431 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n7560) );
  OR2_X1 U6432 ( .A1(n5440), .A2(n5439), .ZN(n5467) );
  OR2_X1 U6433 ( .A1(n5539), .A2(n5538), .ZN(n5566) );
  OR2_X1 U6434 ( .A1(n5625), .A2(n8976), .ZN(n5645) );
  NAND2_X1 U6435 ( .A1(n5109), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5676) );
  OR2_X1 U6436 ( .A1(n5742), .A2(n9007), .ZN(n5820) );
  NOR2_X1 U6437 ( .A1(n9634), .A2(n5806), .ZN(n6512) );
  OR2_X1 U6438 ( .A1(n9226), .A2(n5647), .ZN(n5730) );
  AND2_X1 U6439 ( .A1(n7281), .A2(n7271), .ZN(n7272) );
  INV_X1 U6440 ( .A(n7879), .ZN(n9236) );
  INV_X1 U6441 ( .A(n9424), .ZN(n9270) );
  OR2_X1 U6442 ( .A1(n7804), .A2(n7756), .ZN(n7599) );
  AND2_X1 U6443 ( .A1(n5736), .A2(n5720), .ZN(n5734) );
  NAND2_X1 U6444 ( .A1(n5124), .A2(n5123), .ZN(n5802) );
  INV_X1 U6445 ( .A(n6281), .ZN(n6422) );
  NAND2_X1 U6446 ( .A1(n6405), .A2(n8706), .ZN(n8162) );
  AND2_X1 U6447 ( .A1(n6162), .A2(n6161), .ZN(n8589) );
  AND4_X1 U6448 ( .A1(n6081), .A2(n6080), .A3(n6079), .A4(n6078), .ZN(n8146)
         );
  NAND2_X1 U6449 ( .A1(n6311), .A2(n6310), .ZN(n6419) );
  OR2_X1 U6450 ( .A1(n8408), .A2(n6444), .ZN(n8529) );
  INV_X1 U6451 ( .A(n8479), .ZN(n9752) );
  INV_X1 U6452 ( .A(n8529), .ZN(n9866) );
  INV_X1 U6453 ( .A(n8734), .ZN(n8761) );
  AND2_X1 U6454 ( .A1(n6394), .A2(n6326), .ZN(n6827) );
  NAND2_X1 U6455 ( .A1(n8182), .A2(n7180), .ZN(n9955) );
  INV_X1 U6456 ( .A(n8101), .ZN(n8796) );
  AND2_X1 U6457 ( .A1(n8287), .A2(n8286), .ZN(n8615) );
  INV_X1 U6458 ( .A(n8801), .ZN(n8850) );
  AND2_X1 U6459 ( .A1(n6419), .A2(n6721), .ZN(n6505) );
  AND2_X1 U6460 ( .A1(n6044), .A2(n6032), .ZN(n9805) );
  INV_X1 U6461 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5921) );
  INV_X1 U6462 ( .A(n7561), .ZN(n6535) );
  INV_X1 U6463 ( .A(n9008), .ZN(n9018) );
  OR3_X1 U6464 ( .A1(n5828), .A2(n6522), .A3(n9670), .ZN(n9008) );
  INV_X1 U6465 ( .A(n7745), .ZN(n7816) );
  AND2_X1 U6466 ( .A1(n5748), .A2(n5747), .ZN(n9402) );
  INV_X1 U6467 ( .A(n9584), .ZN(n9564) );
  INV_X1 U6468 ( .A(n9528), .ZN(n9575) );
  AND2_X1 U6469 ( .A1(n7719), .A2(n7877), .ZN(n9252) );
  AND2_X1 U6470 ( .A1(n7705), .A2(n7787), .ZN(n9311) );
  INV_X1 U6471 ( .A(n7621), .ZN(n7329) );
  AND2_X1 U6472 ( .A1(n7668), .A2(n7673), .ZN(n7615) );
  INV_X1 U6473 ( .A(n9664), .ZN(n9677) );
  INV_X1 U6474 ( .A(n9627), .ZN(n9682) );
  AND3_X1 U6475 ( .A1(n6519), .A2(n6518), .A3(n6517), .ZN(n6555) );
  AND2_X1 U6476 ( .A1(n5461), .A2(n5434), .ZN(n6654) );
  AND2_X1 U6477 ( .A1(n7550), .A2(P1_U3086), .ZN(n7367) );
  AND2_X1 U6478 ( .A1(n6722), .A2(n8394), .ZN(n8149) );
  INV_X1 U6479 ( .A(n8312), .ZN(n8545) );
  INV_X1 U6480 ( .A(n8590), .ZN(n8400) );
  INV_X1 U6481 ( .A(n8090), .ZN(n8691) );
  NAND2_X1 U6482 ( .A1(n6441), .A2(n8389), .ZN(n9872) );
  INV_X1 U6483 ( .A(n9888), .ZN(n8699) );
  INV_X1 U6484 ( .A(n8710), .ZN(n9910) );
  NAND2_X1 U6485 ( .A1(n9986), .A2(n9967), .ZN(n8734) );
  INV_X1 U6486 ( .A(n8762), .ZN(n8747) );
  INV_X1 U6487 ( .A(n9986), .ZN(n9984) );
  OR2_X1 U6488 ( .A1(n9970), .A2(n9955), .ZN(n8801) );
  INV_X1 U6489 ( .A(n8851), .ZN(n8821) );
  AND2_X1 U6490 ( .A1(n6329), .A2(n6328), .ZN(n9970) );
  NAND2_X1 U6491 ( .A1(n6506), .A2(n6505), .ZN(n6539) );
  INV_X1 U6492 ( .A(n5857), .ZN(n7824) );
  INV_X1 U6493 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7366) );
  NAND2_X1 U6494 ( .A1(n4611), .A2(P2_U3151), .ZN(n7561) );
  OR2_X1 U6495 ( .A1(n6358), .A2(n6357), .ZN(n6359) );
  INV_X1 U6496 ( .A(n7217), .ZN(n7364) );
  INV_X1 U6497 ( .A(n9303), .ZN(n9445) );
  AND2_X1 U6498 ( .A1(n5810), .A2(n7977), .ZN(n9026) );
  INV_X1 U6499 ( .A(n9402), .ZN(n9194) );
  INV_X1 U6500 ( .A(n9301), .ZN(n9442) );
  NAND2_X1 U6501 ( .A1(n6480), .A2(n6478), .ZN(n9590) );
  INV_X1 U6502 ( .A(n9600), .ZN(n9614) );
  AND2_X1 U6503 ( .A1(n7042), .A2(n7041), .ZN(n9645) );
  NAND2_X1 U6504 ( .A1(n9342), .A2(n6703), .ZN(n9364) );
  NAND2_X1 U6505 ( .A1(n9696), .A2(n9677), .ZN(n9461) );
  INV_X1 U6506 ( .A(n9696), .ZN(n9694) );
  NAND2_X1 U6507 ( .A1(n9685), .A2(n9677), .ZN(n9515) );
  AND2_X1 U6508 ( .A1(n9645), .A2(n9644), .ZN(n9689) );
  AND2_X2 U6509 ( .A1(n6555), .A2(n6668), .ZN(n9685) );
  INV_X1 U6510 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7902) );
  INV_X1 U6511 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7495) );
  INV_X2 U6512 ( .A(n8408), .ZN(P2_U3893) );
  INV_X1 U6513 ( .A(SI_1_), .ZN(n4992) );
  INV_X1 U6514 ( .A(n4998), .ZN(n6450) );
  AND2_X1 U6515 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4993) );
  NAND2_X1 U6516 ( .A1(n6450), .A2(n4993), .ZN(n5874) );
  NAND2_X1 U6517 ( .A1(n4994), .A2(n5874), .ZN(n5142) );
  NAND2_X1 U6518 ( .A1(n5143), .A2(n5142), .ZN(n4997) );
  NAND2_X1 U6519 ( .A1(n4995), .A2(SI_1_), .ZN(n4996) );
  NAND2_X1 U6520 ( .A1(n4997), .A2(n4996), .ZN(n5192) );
  MUX2_X1 U6521 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4998), .Z(n5000) );
  INV_X1 U6522 ( .A(SI_2_), .ZN(n4999) );
  XNOR2_X1 U6523 ( .A(n5000), .B(n4999), .ZN(n5191) );
  NAND2_X1 U6524 ( .A1(n5192), .A2(n5191), .ZN(n5002) );
  NAND2_X1 U6525 ( .A1(n5000), .A2(SI_2_), .ZN(n5001) );
  INV_X1 U6526 ( .A(SI_3_), .ZN(n5003) );
  XNOR2_X1 U6527 ( .A(n5004), .B(n5003), .ZN(n5205) );
  NAND2_X1 U6528 ( .A1(n5004), .A2(SI_3_), .ZN(n5005) );
  INV_X1 U6529 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6459) );
  INV_X1 U6530 ( .A(SI_4_), .ZN(n5006) );
  NAND2_X1 U6531 ( .A1(n5007), .A2(n5006), .ZN(n5010) );
  INV_X1 U6532 ( .A(n5007), .ZN(n5008) );
  NAND2_X1 U6533 ( .A1(n5008), .A2(SI_4_), .ZN(n5009) );
  NAND2_X1 U6534 ( .A1(n5010), .A2(n5009), .ZN(n5226) );
  INV_X1 U6535 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n5011) );
  MUX2_X1 U6536 ( .A(n6462), .B(n5011), .S(n4611), .Z(n5012) );
  NAND2_X1 U6537 ( .A1(n5012), .A2(n10110), .ZN(n5016) );
  INV_X1 U6538 ( .A(n5012), .ZN(n5013) );
  NAND2_X1 U6539 ( .A1(n5013), .A2(SI_5_), .ZN(n5014) );
  NAND2_X1 U6540 ( .A1(n5016), .A2(n5014), .ZN(n5250) );
  INV_X1 U6541 ( .A(n5250), .ZN(n5015) );
  MUX2_X1 U6542 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4611), .Z(n5018) );
  XNOR2_X1 U6543 ( .A(n5018), .B(SI_6_), .ZN(n5283) );
  NAND2_X1 U6544 ( .A1(n5018), .A2(SI_6_), .ZN(n5019) );
  INV_X1 U6545 ( .A(SI_7_), .ZN(n5020) );
  INV_X1 U6546 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n5022) );
  MUX2_X1 U6547 ( .A(n6472), .B(n5022), .S(n4611), .Z(n5024) );
  INV_X1 U6548 ( .A(SI_8_), .ZN(n5023) );
  NAND2_X1 U6549 ( .A1(n5024), .A2(n5023), .ZN(n5027) );
  INV_X1 U6550 ( .A(n5024), .ZN(n5025) );
  NAND2_X1 U6551 ( .A1(n5025), .A2(SI_8_), .ZN(n5026) );
  NAND2_X1 U6552 ( .A1(n5027), .A2(n5026), .ZN(n5329) );
  INV_X1 U6553 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n5028) );
  MUX2_X1 U6554 ( .A(n6502), .B(n5028), .S(n4611), .Z(n5029) );
  NAND2_X1 U6555 ( .A1(n5029), .A2(n10171), .ZN(n5032) );
  INV_X1 U6556 ( .A(n5029), .ZN(n5030) );
  NAND2_X1 U6557 ( .A1(n5030), .A2(SI_9_), .ZN(n5031) );
  MUX2_X1 U6558 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n4611), .Z(n5036) );
  INV_X1 U6559 ( .A(SI_10_), .ZN(n5034) );
  XNOR2_X1 U6560 ( .A(n5036), .B(n5034), .ZN(n5378) );
  INV_X1 U6561 ( .A(n5378), .ZN(n5035) );
  NAND2_X1 U6562 ( .A1(n5036), .A2(SI_10_), .ZN(n5037) );
  MUX2_X1 U6563 ( .A(n6533), .B(n6531), .S(n7550), .Z(n5040) );
  INV_X1 U6564 ( .A(SI_11_), .ZN(n5039) );
  NAND2_X1 U6565 ( .A1(n5040), .A2(n5039), .ZN(n5043) );
  INV_X1 U6566 ( .A(n5040), .ZN(n5041) );
  NAND2_X1 U6567 ( .A1(n5041), .A2(SI_11_), .ZN(n5042) );
  NAND2_X1 U6568 ( .A1(n5043), .A2(n5042), .ZN(n5404) );
  MUX2_X1 U6569 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n7550), .Z(n5044) );
  XNOR2_X1 U6570 ( .A(n5044), .B(n10072), .ZN(n5429) );
  INV_X1 U6571 ( .A(n5429), .ZN(n5046) );
  NAND2_X1 U6572 ( .A1(n5044), .A2(SI_12_), .ZN(n5045) );
  MUX2_X1 U6573 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n7550), .Z(n5458) );
  INV_X1 U6574 ( .A(n5458), .ZN(n5047) );
  NOR2_X1 U6575 ( .A1(n5047), .A2(n10156), .ZN(n5048) );
  MUX2_X1 U6576 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n7550), .Z(n5482) );
  NOR2_X1 U6577 ( .A1(n5482), .A2(SI_14_), .ZN(n5050) );
  NAND2_X1 U6578 ( .A1(n5482), .A2(SI_14_), .ZN(n5049) );
  MUX2_X1 U6579 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n7550), .Z(n5512) );
  INV_X1 U6580 ( .A(n5512), .ZN(n5051) );
  MUX2_X1 U6581 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n7550), .Z(n5530) );
  MUX2_X1 U6582 ( .A(n6849), .B(n6847), .S(n7550), .Z(n5053) );
  INV_X1 U6583 ( .A(n5053), .ZN(n5054) );
  NAND2_X1 U6584 ( .A1(n5054), .A2(SI_17_), .ZN(n5055) );
  NAND2_X1 U6585 ( .A1(n5056), .A2(n5055), .ZN(n5560) );
  MUX2_X1 U6586 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7550), .Z(n5057) );
  XNOR2_X1 U6587 ( .A(n5057), .B(n10155), .ZN(n5579) );
  NAND2_X1 U6588 ( .A1(n5057), .A2(SI_18_), .ZN(n5058) );
  MUX2_X1 U6589 ( .A(n7071), .B(n7567), .S(n7550), .Z(n5059) );
  INV_X1 U6590 ( .A(n5059), .ZN(n5060) );
  NAND2_X1 U6591 ( .A1(n5060), .A2(SI_19_), .ZN(n5061) );
  NAND2_X1 U6592 ( .A1(n5062), .A2(n5061), .ZN(n5599) );
  MUX2_X1 U6593 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n7550), .Z(n5620) );
  MUX2_X1 U6594 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n7550), .Z(n5639) );
  NOR2_X1 U6595 ( .A1(n5639), .A2(SI_21_), .ZN(n5063) );
  NAND2_X1 U6596 ( .A1(n5639), .A2(SI_21_), .ZN(n5064) );
  MUX2_X1 U6597 ( .A(n7315), .B(n7313), .S(n7550), .Z(n5066) );
  INV_X1 U6598 ( .A(SI_22_), .ZN(n10087) );
  NAND2_X1 U6599 ( .A1(n5066), .A2(n10087), .ZN(n5668) );
  INV_X1 U6600 ( .A(n5066), .ZN(n5067) );
  NAND2_X1 U6601 ( .A1(n5067), .A2(SI_22_), .ZN(n5068) );
  NAND2_X1 U6602 ( .A1(n5668), .A2(n5068), .ZN(n5666) );
  XNOR2_X1 U6603 ( .A(n5667), .B(n5666), .ZN(n7312) );
  INV_X1 U6604 ( .A(n5285), .ZN(n5070) );
  NOR2_X1 U6605 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5078) );
  NOR2_X1 U6606 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5077) );
  NAND2_X2 U6607 ( .A1(n5815), .A2(n7891), .ZN(n6474) );
  NAND2_X2 U6608 ( .A1(n6474), .A2(n4611), .ZN(n5193) );
  NAND2_X1 U6609 ( .A1(n7312), .A2(n7590), .ZN(n5084) );
  NAND2_X2 U6610 ( .A1(n6450), .A2(n6474), .ZN(n5194) );
  OR2_X1 U6611 ( .A1(n7596), .A2(n7313), .ZN(n5083) );
  INV_X1 U6612 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5085) );
  NAND2_X1 U6613 ( .A1(n5128), .A2(n5127), .ZN(n5086) );
  NOR2_X2 U6614 ( .A1(n5126), .A2(n5086), .ZN(n5098) );
  NAND2_X1 U6615 ( .A1(n5091), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5092) );
  NAND2_X1 U6616 ( .A1(n5093), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5094) );
  MUX2_X1 U6617 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5094), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5095) );
  NAND2_X1 U6618 ( .A1(n5095), .A2(n5091), .ZN(n7520) );
  INV_X1 U6619 ( .A(n7520), .ZN(n5096) );
  INV_X1 U6620 ( .A(n5098), .ZN(n5099) );
  NAND2_X1 U6621 ( .A1(n5099), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5100) );
  MUX2_X1 U6622 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5100), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n5101) );
  NAND2_X1 U6623 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n5259) );
  INV_X1 U6624 ( .A(n5259), .ZN(n5102) );
  NAND2_X1 U6625 ( .A1(n5257), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5317) );
  INV_X1 U6626 ( .A(n5317), .ZN(n5103) );
  NAND2_X1 U6627 ( .A1(n5103), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5336) );
  INV_X1 U6628 ( .A(n5364), .ZN(n5104) );
  NAND2_X1 U6629 ( .A1(n5104), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n5387) );
  INV_X1 U6630 ( .A(n5387), .ZN(n5105) );
  NAND2_X1 U6631 ( .A1(n5465), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5520) );
  INV_X1 U6632 ( .A(n5520), .ZN(n5106) );
  NAND2_X1 U6633 ( .A1(n5106), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5539) );
  INV_X1 U6634 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5585) );
  INV_X1 U6635 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n8976) );
  XNOR2_X1 U6636 ( .A(n5676), .B(P1_REG3_REG_22__SCAN_IN), .ZN(n9267) );
  INV_X1 U6637 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5110) );
  NAND2_X1 U6638 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_28__SCAN_IN), 
        .ZN(n5111) );
  NAND2_X1 U6639 ( .A1(n5112), .A2(n5111), .ZN(n5113) );
  XNOR2_X2 U6640 ( .A(n5113), .B(n7554), .ZN(n5114) );
  NAND2_X1 U6641 ( .A1(n9267), .A2(n5442), .ZN(n5121) );
  INV_X1 U6642 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5118) );
  INV_X1 U6643 ( .A(n5114), .ZN(n9523) );
  NAND2_X1 U6644 ( .A1(n5160), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5117) );
  NAND2_X1 U6645 ( .A1(n6493), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5116) );
  OAI211_X1 U6646 ( .C1(n6494), .C2(n5118), .A(n5117), .B(n5116), .ZN(n5119)
         );
  INV_X1 U6647 ( .A(n5119), .ZN(n5120) );
  NAND2_X1 U6648 ( .A1(n5126), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5562) );
  NAND2_X1 U6649 ( .A1(n5562), .A2(n5127), .ZN(n5581) );
  INV_X1 U6650 ( .A(n5128), .ZN(n5129) );
  AND2_X1 U6651 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n5130) );
  NAND2_X1 U6652 ( .A1(n5581), .A2(n5130), .ZN(n5135) );
  NAND2_X1 U6653 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n5131) );
  NAND2_X1 U6654 ( .A1(n5131), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5132) );
  OAI21_X1 U6655 ( .B1(n5133), .B2(P1_IR_REG_31__SCAN_IN), .A(n5132), .ZN(
        n5134) );
  AND3_X2 U6656 ( .A1(n5136), .A2(n5135), .A3(n5134), .ZN(n7844) );
  INV_X2 U6657 ( .A(n7844), .ZN(n7815) );
  NAND2_X1 U6658 ( .A1(n6522), .A2(n6702), .ZN(n5137) );
  NAND2_X1 U6659 ( .A1(n6523), .A2(n5137), .ZN(n5138) );
  INV_X1 U6660 ( .A(n5169), .ZN(n5172) );
  NAND2_X1 U6661 ( .A1(n5138), .A2(n5172), .ZN(n5155) );
  OAI22_X1 U6662 ( .A1(n9426), .A2(n6337), .B1(n9417), .B2(n6343), .ZN(n8984)
         );
  NAND2_X1 U6663 ( .A1(n6523), .A2(n6702), .ZN(n5139) );
  OR2_X4 U6664 ( .A1(n5169), .A2(n5139), .ZN(n5752) );
  INV_X1 U6665 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6666 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5140) );
  XNOR2_X1 U6667 ( .A(n5141), .B(n5140), .ZN(n6581) );
  INV_X1 U6668 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6457) );
  XNOR2_X1 U6669 ( .A(n5143), .B(n5142), .ZN(n6465) );
  NAND2_X1 U6670 ( .A1(n5361), .A2(n4449), .ZN(n5153) );
  INV_X1 U6671 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n5146) );
  INV_X1 U6672 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5147) );
  OR2_X1 U6673 ( .A1(n5215), .A2(n5147), .ZN(n5150) );
  NAND2_X1 U6674 ( .A1(n5213), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6675 ( .A1(n5239), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n5148) );
  NAND4_X1 U6676 ( .A1(n5151), .A2(n5150), .A3(n5149), .A4(n5148), .ZN(n5154)
         );
  NAND2_X1 U6677 ( .A1(n5154), .A2(n5775), .ZN(n5152) );
  INV_X2 U6678 ( .A(n5752), .ZN(n5222) );
  INV_X1 U6679 ( .A(n5155), .ZN(n5174) );
  AOI22_X1 U6680 ( .A1(n5154), .A2(n5174), .B1(n5775), .B2(n4449), .ZN(n5157)
         );
  INV_X1 U6681 ( .A(n5157), .ZN(n5156) );
  INV_X1 U6682 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U6683 ( .A1(n5160), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5163) );
  NAND2_X1 U6684 ( .A1(n5213), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n5162) );
  NAND2_X1 U6685 ( .A1(n5239), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5161) );
  NAND2_X1 U6686 ( .A1(n9045), .A2(n5775), .ZN(n5168) );
  INV_X1 U6687 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5171) );
  NAND2_X1 U6688 ( .A1(n4611), .A2(SI_0_), .ZN(n5166) );
  INV_X1 U6689 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5165) );
  XNOR2_X1 U6690 ( .A(n5166), .B(n5165), .ZN(n9526) );
  MUX2_X1 U6691 ( .A(n5171), .B(n9526), .S(n6474), .Z(n6549) );
  INV_X1 U6692 ( .A(n6549), .ZN(n6680) );
  NAND2_X1 U6693 ( .A1(n6680), .A2(n5361), .ZN(n5167) );
  NAND2_X1 U6694 ( .A1(n5169), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6695 ( .A1(n5177), .A2(n5170), .ZN(n6616) );
  OAI22_X1 U6696 ( .A1(n6549), .A2(n6337), .B1(n5172), .B2(n5171), .ZN(n5173)
         );
  INV_X1 U6697 ( .A(n5173), .ZN(n5176) );
  NAND2_X1 U6698 ( .A1(n9045), .A2(n5174), .ZN(n5175) );
  NAND2_X1 U6699 ( .A1(n5176), .A2(n5175), .ZN(n6615) );
  NAND2_X1 U6700 ( .A1(n6616), .A2(n6615), .ZN(n5179) );
  NAND2_X1 U6701 ( .A1(n5177), .A2(n5222), .ZN(n5178) );
  NAND2_X1 U6702 ( .A1(n5179), .A2(n5178), .ZN(n6730) );
  NAND2_X1 U6703 ( .A1(n5181), .A2(n5180), .ZN(n6728) );
  NAND2_X1 U6704 ( .A1(n6728), .A2(n6852), .ZN(n5203) );
  INV_X1 U6705 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n5182) );
  INV_X1 U6706 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5183) );
  OR2_X1 U6707 ( .A1(n5215), .A2(n5183), .ZN(n5187) );
  NAND2_X1 U6708 ( .A1(n5239), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5185) );
  NAND2_X1 U6709 ( .A1(n5213), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5184) );
  NAND2_X1 U6710 ( .A1(n9043), .A2(n5775), .ZN(n5198) );
  OR2_X1 U6711 ( .A1(n5189), .A2(n5408), .ZN(n5233) );
  INV_X1 U6712 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U6713 ( .A1(n5233), .A2(n5190), .ZN(n5207) );
  OAI21_X1 U6714 ( .B1(n5233), .B2(n5190), .A(n5207), .ZN(n6580) );
  XNOR2_X1 U6715 ( .A(n5192), .B(n5191), .ZN(n6453) );
  OR2_X1 U6716 ( .A1(n5193), .A2(n6453), .ZN(n5196) );
  INV_X1 U6717 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6454) );
  NAND2_X1 U6718 ( .A1(n5361), .A2(n4354), .ZN(n5197) );
  NAND2_X1 U6719 ( .A1(n5198), .A2(n5197), .ZN(n5199) );
  XNOR2_X1 U6720 ( .A(n5199), .B(n5222), .ZN(n5201) );
  AOI22_X1 U6721 ( .A1(n9043), .A2(n5174), .B1(n5775), .B2(n4354), .ZN(n5200)
         );
  NAND2_X1 U6722 ( .A1(n5201), .A2(n5200), .ZN(n5204) );
  NAND2_X1 U6723 ( .A1(n5203), .A2(n6851), .ZN(n6850) );
  NAND2_X1 U6724 ( .A1(n6850), .A2(n5204), .ZN(n8885) );
  XNOR2_X1 U6725 ( .A(n5205), .B(n5206), .ZN(n6455) );
  OR2_X1 U6726 ( .A1(n5193), .A2(n6455), .ZN(n5212) );
  INV_X1 U6727 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6456) );
  OR2_X1 U6728 ( .A1(n5194), .A2(n6456), .ZN(n5211) );
  NAND2_X1 U6729 ( .A1(n5207), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5209) );
  INV_X1 U6730 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5208) );
  XNOR2_X1 U6731 ( .A(n5209), .B(n5208), .ZN(n6585) );
  OR2_X1 U6732 ( .A1(n6474), .A2(n6585), .ZN(n5210) );
  AND3_X2 U6733 ( .A1(n5212), .A2(n5211), .A3(n5210), .ZN(n8891) );
  NAND2_X1 U6734 ( .A1(n9623), .A2(n5325), .ZN(n5221) );
  INV_X1 U6735 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8893) );
  NAND2_X1 U6736 ( .A1(n5239), .A2(n8893), .ZN(n5219) );
  NAND2_X1 U6737 ( .A1(n5213), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5218) );
  INV_X1 U6738 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6584) );
  OR2_X1 U6739 ( .A1(n6488), .A2(n6584), .ZN(n5217) );
  INV_X1 U6740 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5214) );
  OR2_X1 U6741 ( .A1(n5215), .A2(n5214), .ZN(n5216) );
  NAND2_X1 U6742 ( .A1(n9042), .A2(n5775), .ZN(n5220) );
  NAND2_X1 U6743 ( .A1(n5221), .A2(n5220), .ZN(n5223) );
  NAND2_X1 U6744 ( .A1(n9042), .A2(n5174), .ZN(n5225) );
  OR2_X1 U6745 ( .A1(n6337), .A2(n8891), .ZN(n5224) );
  NAND2_X1 U6746 ( .A1(n5225), .A2(n5224), .ZN(n5271) );
  XNOR2_X1 U6747 ( .A(n5273), .B(n5271), .ZN(n8886) );
  NAND2_X1 U6748 ( .A1(n8885), .A2(n8886), .ZN(n6871) );
  NAND2_X1 U6749 ( .A1(n5227), .A2(n5226), .ZN(n5228) );
  AND2_X1 U6750 ( .A1(n5229), .A2(n5228), .ZN(n6458) );
  OR2_X1 U6751 ( .A1(n7596), .A2(n5230), .ZN(n5235) );
  OR2_X1 U6752 ( .A1(n5231), .A2(n5408), .ZN(n5232) );
  NAND2_X1 U6753 ( .A1(n5233), .A2(n5232), .ZN(n5253) );
  XNOR2_X1 U6754 ( .A(n5253), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6587) );
  OR2_X1 U6755 ( .A1(n6474), .A2(n6587), .ZN(n5234) );
  AND3_X2 U6756 ( .A1(n5236), .A2(n5235), .A3(n5234), .ZN(n9615) );
  INV_X1 U6757 ( .A(n5361), .ZN(n5683) );
  NAND2_X1 U6758 ( .A1(n5725), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n5245) );
  INV_X1 U6759 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6760 ( .A1(n8893), .A2(n5237), .ZN(n5238) );
  AND2_X1 U6761 ( .A1(n5238), .A2(n5259), .ZN(n9611) );
  NAND2_X1 U6762 ( .A1(n5239), .A2(n9611), .ZN(n5244) );
  INV_X1 U6763 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5240) );
  OR2_X1 U6764 ( .A1(n6488), .A2(n5240), .ZN(n5243) );
  INV_X1 U6765 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5241) );
  OR2_X1 U6766 ( .A1(n6495), .A2(n5241), .ZN(n5242) );
  NAND4_X2 U6767 ( .A1(n5245), .A2(n5244), .A3(n5243), .A4(n5242), .ZN(n9041)
         );
  NAND2_X1 U6768 ( .A1(n9041), .A2(n5775), .ZN(n5246) );
  OAI21_X1 U6769 ( .B1(n9615), .B2(n5683), .A(n5246), .ZN(n5247) );
  XNOR2_X1 U6770 ( .A(n5247), .B(n5752), .ZN(n6873) );
  NAND2_X1 U6771 ( .A1(n9041), .A2(n5174), .ZN(n5249) );
  OR2_X1 U6772 ( .A1(n9615), .A2(n6337), .ZN(n5248) );
  NAND2_X1 U6773 ( .A1(n5249), .A2(n5248), .ZN(n6874) );
  XNOR2_X1 U6774 ( .A(n5251), .B(n5250), .ZN(n6461) );
  INV_X1 U6775 ( .A(n6461), .ZN(n5252) );
  NAND2_X1 U6776 ( .A1(n5252), .A2(n7590), .ZN(n5256) );
  OAI21_X1 U6777 ( .B1(n5253), .B2(P1_IR_REG_4__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5254) );
  XNOR2_X1 U6778 ( .A(n5254), .B(P1_IR_REG_5__SCAN_IN), .ZN(n9110) );
  AOI22_X1 U6779 ( .A1(n5602), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5601), .B2(
        n9110), .ZN(n5255) );
  INV_X1 U6780 ( .A(n5257), .ZN(n5292) );
  INV_X1 U6781 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5258) );
  NAND2_X1 U6782 ( .A1(n5259), .A2(n5258), .ZN(n5260) );
  AND2_X1 U6783 ( .A1(n5292), .A2(n5260), .ZN(n6882) );
  NAND2_X1 U6784 ( .A1(n5239), .A2(n6882), .ZN(n5266) );
  NAND2_X1 U6785 ( .A1(n5725), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5265) );
  INV_X1 U6786 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5261) );
  OR2_X1 U6787 ( .A1(n6495), .A2(n5261), .ZN(n5264) );
  INV_X1 U6788 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n5262) );
  OR2_X1 U6789 ( .A1(n6494), .A2(n5262), .ZN(n5263) );
  NAND2_X1 U6790 ( .A1(n9040), .A2(n5775), .ZN(n5267) );
  OAI21_X1 U6791 ( .B1(n9630), .B2(n5683), .A(n5267), .ZN(n5268) );
  OR2_X1 U6792 ( .A1(n9630), .A2(n6337), .ZN(n5270) );
  NAND2_X1 U6793 ( .A1(n9040), .A2(n5174), .ZN(n5269) );
  AND2_X1 U6794 ( .A1(n5270), .A2(n5269), .ZN(n5277) );
  NAND2_X1 U6795 ( .A1(n6877), .A2(n5277), .ZN(n5274) );
  INV_X1 U6796 ( .A(n5271), .ZN(n5272) );
  NAND2_X1 U6797 ( .A1(n5273), .A2(n5272), .ZN(n8962) );
  OAI211_X1 U6798 ( .C1(n6873), .C2(n6874), .A(n5274), .B(n8962), .ZN(n5275)
         );
  INV_X1 U6799 ( .A(n5275), .ZN(n5276) );
  NAND2_X1 U6800 ( .A1(n6871), .A2(n5276), .ZN(n5282) );
  INV_X1 U6801 ( .A(n6877), .ZN(n5280) );
  NAND2_X1 U6802 ( .A1(n6875), .A2(n5277), .ZN(n5279) );
  INV_X1 U6803 ( .A(n6875), .ZN(n5278) );
  INV_X1 U6804 ( .A(n5277), .ZN(n6876) );
  AOI22_X1 U6805 ( .A1(n5280), .A2(n5279), .B1(n5278), .B2(n6876), .ZN(n5281)
         );
  NAND2_X1 U6806 ( .A1(n5282), .A2(n5281), .ZN(n6775) );
  XNOR2_X1 U6807 ( .A(n5284), .B(n5283), .ZN(n6464) );
  OR2_X1 U6808 ( .A1(n6464), .A2(n5193), .ZN(n5290) );
  NAND2_X1 U6809 ( .A1(n5285), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5286) );
  MUX2_X1 U6810 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5286), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n5288) );
  AND2_X1 U6811 ( .A1(n5288), .A2(n5287), .ZN(n9563) );
  AOI22_X1 U6812 ( .A1(n5602), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5601), .B2(
        n9563), .ZN(n5289) );
  NAND2_X1 U6813 ( .A1(n6783), .A2(n5325), .ZN(n5301) );
  INV_X1 U6814 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5291) );
  NAND2_X1 U6815 ( .A1(n5292), .A2(n5291), .ZN(n5293) );
  AND2_X1 U6816 ( .A1(n5317), .A2(n5293), .ZN(n6778) );
  NAND2_X1 U6817 ( .A1(n5239), .A2(n6778), .ZN(n5299) );
  NAND2_X1 U6818 ( .A1(n5725), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5298) );
  INV_X1 U6819 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5294) );
  OR2_X1 U6820 ( .A1(n6495), .A2(n5294), .ZN(n5297) );
  INV_X1 U6821 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5295) );
  OR2_X1 U6822 ( .A1(n6488), .A2(n5295), .ZN(n5296) );
  NAND2_X1 U6823 ( .A1(n6922), .A2(n6341), .ZN(n5300) );
  NAND2_X1 U6824 ( .A1(n5301), .A2(n5300), .ZN(n5302) );
  XNOR2_X1 U6825 ( .A(n5302), .B(n5222), .ZN(n5305) );
  NAND2_X1 U6826 ( .A1(n6783), .A2(n6341), .ZN(n5304) );
  NAND2_X1 U6827 ( .A1(n6922), .A2(n5174), .ZN(n5303) );
  AND2_X1 U6828 ( .A1(n5304), .A2(n5303), .ZN(n5306) );
  NAND2_X1 U6829 ( .A1(n5305), .A2(n5306), .ZN(n6773) );
  NAND2_X1 U6830 ( .A1(n6775), .A2(n6773), .ZN(n5309) );
  INV_X1 U6831 ( .A(n5305), .ZN(n5308) );
  INV_X1 U6832 ( .A(n5306), .ZN(n5307) );
  NAND2_X1 U6833 ( .A1(n5308), .A2(n5307), .ZN(n6774) );
  OR2_X1 U6834 ( .A1(n6468), .A2(n5193), .ZN(n5314) );
  NAND2_X1 U6835 ( .A1(n5287), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5312) );
  XNOR2_X1 U6836 ( .A(n5312), .B(P1_IR_REG_7__SCAN_IN), .ZN(n9123) );
  AOI22_X1 U6837 ( .A1(n5602), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5601), .B2(
        n9123), .ZN(n5313) );
  NAND2_X1 U6838 ( .A1(n7031), .A2(n6341), .ZN(n5324) );
  INV_X1 U6839 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n5315) );
  OR2_X1 U6840 ( .A1(n6495), .A2(n5315), .ZN(n5322) );
  INV_X1 U6841 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6591) );
  OR2_X1 U6842 ( .A1(n6488), .A2(n6591), .ZN(n5321) );
  INV_X1 U6843 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5316) );
  NAND2_X1 U6844 ( .A1(n5317), .A2(n5316), .ZN(n5318) );
  AND2_X1 U6845 ( .A1(n5336), .A2(n5318), .ZN(n6938) );
  NAND2_X1 U6846 ( .A1(n5442), .A2(n6938), .ZN(n5320) );
  NAND2_X1 U6847 ( .A1(n6493), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5319) );
  NAND2_X1 U6848 ( .A1(n9039), .A2(n5174), .ZN(n5323) );
  NAND2_X1 U6849 ( .A1(n5324), .A2(n5323), .ZN(n6888) );
  NAND2_X1 U6850 ( .A1(n7031), .A2(n5325), .ZN(n5327) );
  NAND2_X1 U6851 ( .A1(n9039), .A2(n6341), .ZN(n5326) );
  NAND2_X1 U6852 ( .A1(n5327), .A2(n5326), .ZN(n5328) );
  XNOR2_X1 U6853 ( .A(n5328), .B(n5752), .ZN(n6887) );
  XNOR2_X1 U6854 ( .A(n5330), .B(n5329), .ZN(n6469) );
  NAND2_X1 U6855 ( .A1(n6469), .A2(n7590), .ZN(n5332) );
  NOR2_X1 U6856 ( .A1(n5287), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5381) );
  INV_X1 U6857 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5408) );
  OR2_X1 U6858 ( .A1(n5381), .A2(n5408), .ZN(n5356) );
  XNOR2_X1 U6859 ( .A(n5356), .B(P1_IR_REG_8__SCAN_IN), .ZN(n9550) );
  AOI22_X1 U6860 ( .A1(n5602), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5601), .B2(
        n9550), .ZN(n5331) );
  NAND2_X1 U6861 ( .A1(n5332), .A2(n5331), .ZN(n7080) );
  NAND2_X1 U6862 ( .A1(n7080), .A2(n5325), .ZN(n5343) );
  INV_X1 U6863 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n5333) );
  OR2_X1 U6864 ( .A1(n6494), .A2(n5333), .ZN(n5341) );
  INV_X1 U6865 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5334) );
  OR2_X1 U6866 ( .A1(n6495), .A2(n5334), .ZN(n5340) );
  NAND2_X1 U6867 ( .A1(n6493), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6868 ( .A1(n5336), .A2(n5335), .ZN(n5337) );
  AND2_X1 U6869 ( .A1(n5364), .A2(n5337), .ZN(n7046) );
  NAND2_X1 U6870 ( .A1(n5239), .A2(n7046), .ZN(n5338) );
  NAND2_X1 U6871 ( .A1(n9646), .A2(n5775), .ZN(n5342) );
  NAND2_X1 U6872 ( .A1(n5343), .A2(n5342), .ZN(n5344) );
  XNOR2_X1 U6873 ( .A(n5344), .B(n5752), .ZN(n5347) );
  NAND2_X1 U6874 ( .A1(n5346), .A2(n5345), .ZN(n5353) );
  NAND2_X1 U6875 ( .A1(n5348), .A2(n5347), .ZN(n5349) );
  NAND2_X1 U6876 ( .A1(n7080), .A2(n6341), .ZN(n5351) );
  NAND2_X1 U6877 ( .A1(n9646), .A2(n5174), .ZN(n5350) );
  NAND2_X1 U6878 ( .A1(n5351), .A2(n5350), .ZN(n6957) );
  INV_X1 U6879 ( .A(n6957), .ZN(n5352) );
  XNOR2_X1 U6880 ( .A(n5354), .B(n4990), .ZN(n6485) );
  NAND2_X1 U6881 ( .A1(n6485), .A2(n7590), .ZN(n5360) );
  INV_X1 U6882 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n5355) );
  NAND2_X1 U6883 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  NAND2_X1 U6884 ( .A1(n5357), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5358) );
  XNOR2_X1 U6885 ( .A(n5358), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9142) );
  AOI22_X1 U6886 ( .A1(n5602), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5601), .B2(
        n9142), .ZN(n5359) );
  NAND2_X1 U6887 ( .A1(n5360), .A2(n5359), .ZN(n9648) );
  NAND2_X1 U6888 ( .A1(n9648), .A2(n5325), .ZN(n5371) );
  INV_X1 U6889 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n5362) );
  OR2_X1 U6890 ( .A1(n6488), .A2(n5362), .ZN(n5369) );
  INV_X1 U6891 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n5363) );
  OR2_X1 U6892 ( .A1(n6495), .A2(n5363), .ZN(n5368) );
  NAND2_X1 U6893 ( .A1(n6493), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n5367) );
  INV_X1 U6894 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7015) );
  NAND2_X1 U6895 ( .A1(n5364), .A2(n7015), .ZN(n5365) );
  AND2_X1 U6896 ( .A1(n5387), .A2(n5365), .ZN(n7112) );
  NAND2_X1 U6897 ( .A1(n5442), .A2(n7112), .ZN(n5366) );
  NAND2_X1 U6898 ( .A1(n9038), .A2(n6341), .ZN(n5370) );
  NAND2_X1 U6899 ( .A1(n5371), .A2(n5370), .ZN(n5372) );
  XNOR2_X1 U6900 ( .A(n5372), .B(n5752), .ZN(n5374) );
  NOR2_X1 U6901 ( .A1(n9655), .A2(n6343), .ZN(n5373) );
  AOI21_X1 U6902 ( .B1(n9648), .B2(n6341), .A(n5373), .ZN(n5375) );
  XNOR2_X1 U6903 ( .A(n5374), .B(n5375), .ZN(n7013) );
  NAND2_X1 U6904 ( .A1(n7010), .A2(n7013), .ZN(n7011) );
  INV_X1 U6905 ( .A(n5374), .ZN(n5376) );
  NAND2_X1 U6906 ( .A1(n5376), .A2(n5375), .ZN(n5377) );
  NAND2_X1 U6907 ( .A1(n7011), .A2(n5377), .ZN(n5400) );
  INV_X1 U6908 ( .A(n5400), .ZN(n5398) );
  XNOR2_X1 U6909 ( .A(n5379), .B(n5378), .ZN(n6503) );
  NAND2_X1 U6910 ( .A1(n6503), .A2(n7590), .ZN(n5384) );
  NOR2_X1 U6911 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5380) );
  AND2_X1 U6912 ( .A1(n5381), .A2(n5380), .ZN(n5407) );
  OR2_X1 U6913 ( .A1(n5407), .A2(n5408), .ZN(n5382) );
  XNOR2_X1 U6914 ( .A(n5382), .B(P1_IR_REG_10__SCAN_IN), .ZN(n9538) );
  AOI22_X1 U6915 ( .A1(n5602), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5601), .B2(
        n9538), .ZN(n5383) );
  NAND2_X1 U6916 ( .A1(n9658), .A2(n5325), .ZN(n5395) );
  NAND2_X1 U6917 ( .A1(n5608), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5393) );
  INV_X1 U6918 ( .A(n5385), .ZN(n5413) );
  INV_X1 U6919 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U6920 ( .A1(n5387), .A2(n5386), .ZN(n5388) );
  AND2_X1 U6921 ( .A1(n5413), .A2(n5388), .ZN(n7250) );
  NAND2_X1 U6922 ( .A1(n5442), .A2(n7250), .ZN(n5392) );
  INV_X1 U6923 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5389) );
  OR2_X1 U6924 ( .A1(n6495), .A2(n5389), .ZN(n5391) );
  NAND2_X1 U6925 ( .A1(n6493), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6926 ( .A1(n9037), .A2(n6341), .ZN(n5394) );
  NAND2_X1 U6927 ( .A1(n5395), .A2(n5394), .ZN(n5396) );
  XNOR2_X1 U6928 ( .A(n5396), .B(n5222), .ZN(n5399) );
  INV_X1 U6929 ( .A(n5399), .ZN(n5397) );
  NAND2_X1 U6930 ( .A1(n9658), .A2(n6341), .ZN(n5402) );
  NAND2_X1 U6931 ( .A1(n9037), .A2(n5174), .ZN(n5401) );
  NAND2_X1 U6932 ( .A1(n5402), .A2(n5401), .ZN(n7248) );
  NAND2_X1 U6933 ( .A1(n7246), .A2(n7302), .ZN(n5428) );
  XNOR2_X1 U6934 ( .A(n5405), .B(n5404), .ZN(n6530) );
  NAND2_X1 U6935 ( .A1(n6530), .A2(n7590), .ZN(n5411) );
  INV_X1 U6936 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5406) );
  AND2_X1 U6937 ( .A1(n5407), .A2(n5406), .ZN(n5432) );
  OR2_X1 U6938 ( .A1(n5432), .A2(n5408), .ZN(n5409) );
  XNOR2_X1 U6939 ( .A(n5409), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6596) );
  AOI22_X1 U6940 ( .A1(n5602), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5601), .B2(
        n6596), .ZN(n5410) );
  NAND2_X1 U6941 ( .A1(n9601), .A2(n5325), .ZN(n5420) );
  INV_X1 U6942 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n5412) );
  OR2_X1 U6943 ( .A1(n6495), .A2(n5412), .ZN(n5418) );
  INV_X1 U6944 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n6595) );
  OR2_X1 U6945 ( .A1(n6488), .A2(n6595), .ZN(n5417) );
  INV_X1 U6946 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7307) );
  NAND2_X1 U6947 ( .A1(n5413), .A2(n7307), .ZN(n5414) );
  AND2_X1 U6948 ( .A1(n5440), .A2(n5414), .ZN(n9599) );
  NAND2_X1 U6949 ( .A1(n5442), .A2(n9599), .ZN(n5416) );
  NAND2_X1 U6950 ( .A1(n6493), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6951 ( .A1(n9036), .A2(n6341), .ZN(n5419) );
  NAND2_X1 U6952 ( .A1(n5420), .A2(n5419), .ZN(n5421) );
  XNOR2_X1 U6953 ( .A(n5421), .B(n5222), .ZN(n5423) );
  NOR2_X1 U6954 ( .A1(n9654), .A2(n6343), .ZN(n5422) );
  AOI21_X1 U6955 ( .B1(n9601), .B2(n6341), .A(n5422), .ZN(n5424) );
  NAND2_X1 U6956 ( .A1(n5423), .A2(n5424), .ZN(n7351) );
  INV_X1 U6957 ( .A(n5423), .ZN(n5426) );
  INV_X1 U6958 ( .A(n5424), .ZN(n5425) );
  NAND2_X1 U6959 ( .A1(n5426), .A2(n5425), .ZN(n5427) );
  AND2_X1 U6960 ( .A1(n7351), .A2(n5427), .ZN(n7303) );
  NAND2_X1 U6961 ( .A1(n5428), .A2(n7303), .ZN(n7305) );
  NAND2_X1 U6962 ( .A1(n7305), .A2(n7351), .ZN(n5456) );
  XNOR2_X1 U6963 ( .A(n5430), .B(n5429), .ZN(n6534) );
  NAND2_X1 U6964 ( .A1(n6534), .A2(n7590), .ZN(n5436) );
  INV_X1 U6965 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5431) );
  NAND2_X1 U6966 ( .A1(n5432), .A2(n5431), .ZN(n5488) );
  NAND2_X1 U6967 ( .A1(n5488), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5433) );
  INV_X1 U6968 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5486) );
  NAND2_X1 U6969 ( .A1(n5433), .A2(n5486), .ZN(n5461) );
  OR2_X1 U6970 ( .A1(n5433), .A2(n5486), .ZN(n5434) );
  AOI22_X1 U6971 ( .A1(n5602), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5601), .B2(
        n6654), .ZN(n5435) );
  NAND2_X1 U6972 ( .A1(n7217), .A2(n5325), .ZN(n5448) );
  INV_X1 U6973 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5437) );
  OR2_X1 U6974 ( .A1(n6495), .A2(n5437), .ZN(n5446) );
  INV_X1 U6975 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n5438) );
  OR2_X1 U6976 ( .A1(n6494), .A2(n5438), .ZN(n5445) );
  NAND2_X1 U6977 ( .A1(n5440), .A2(n5439), .ZN(n5441) );
  AND2_X1 U6978 ( .A1(n5467), .A2(n5441), .ZN(n7361) );
  NAND2_X1 U6979 ( .A1(n5442), .A2(n7361), .ZN(n5444) );
  NAND2_X1 U6980 ( .A1(n6493), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5443) );
  INV_X1 U6981 ( .A(n9673), .ZN(n9035) );
  NAND2_X1 U6982 ( .A1(n9035), .A2(n6341), .ZN(n5447) );
  NAND2_X1 U6983 ( .A1(n5448), .A2(n5447), .ZN(n5449) );
  XNOR2_X1 U6984 ( .A(n5449), .B(n5222), .ZN(n5451) );
  NOR2_X1 U6985 ( .A1(n9673), .A2(n6343), .ZN(n5450) );
  AOI21_X1 U6986 ( .B1(n7217), .B2(n6341), .A(n5450), .ZN(n5452) );
  NAND2_X1 U6987 ( .A1(n5451), .A2(n5452), .ZN(n5457) );
  INV_X1 U6988 ( .A(n5451), .ZN(n5454) );
  INV_X1 U6989 ( .A(n5452), .ZN(n5453) );
  NAND2_X1 U6990 ( .A1(n5454), .A2(n5453), .ZN(n5455) );
  AND2_X1 U6991 ( .A1(n5457), .A2(n5455), .ZN(n7352) );
  NAND2_X1 U6992 ( .A1(n5456), .A2(n7352), .ZN(n7355) );
  NAND2_X1 U6993 ( .A1(n7355), .A2(n5457), .ZN(n7372) );
  XNOR2_X1 U6994 ( .A(n5458), .B(SI_13_), .ZN(n5459) );
  XNOR2_X1 U6995 ( .A(n5460), .B(n5459), .ZN(n6621) );
  NAND2_X1 U6996 ( .A1(n6621), .A2(n7590), .ZN(n5464) );
  NAND2_X1 U6997 ( .A1(n5461), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5462) );
  XNOR2_X1 U6998 ( .A(n5462), .B(P1_IR_REG_13__SCAN_IN), .ZN(n6747) );
  AOI22_X1 U6999 ( .A1(n5602), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5601), .B2(
        n6747), .ZN(n5463) );
  INV_X1 U7000 ( .A(n5465), .ZN(n5496) );
  NAND2_X1 U7001 ( .A1(n5467), .A2(n5466), .ZN(n5468) );
  AND2_X1 U7002 ( .A1(n5496), .A2(n5468), .ZN(n7378) );
  NAND2_X1 U7003 ( .A1(n5442), .A2(n7378), .ZN(n5474) );
  NAND2_X1 U7004 ( .A1(n5725), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5473) );
  INV_X1 U7005 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5469) );
  OR2_X1 U7006 ( .A1(n6495), .A2(n5469), .ZN(n5472) );
  INV_X1 U7007 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n5470) );
  OR2_X1 U7008 ( .A1(n6488), .A2(n5470), .ZN(n5471) );
  NAND4_X1 U7009 ( .A1(n5474), .A2(n5473), .A3(n5472), .A4(n5471), .ZN(n9034)
         );
  OAI22_X1 U7010 ( .A1(n7381), .A2(n5683), .B1(n8867), .B2(n6337), .ZN(n5475)
         );
  XNOR2_X1 U7011 ( .A(n5475), .B(n5222), .ZN(n5480) );
  OR2_X1 U7012 ( .A1(n7381), .A2(n6337), .ZN(n5477) );
  NAND2_X1 U7013 ( .A1(n9034), .A2(n5174), .ZN(n5476) );
  NAND2_X1 U7014 ( .A1(n5477), .A2(n5476), .ZN(n5478) );
  XNOR2_X1 U7015 ( .A(n5480), .B(n5478), .ZN(n7373) );
  NAND2_X1 U7016 ( .A1(n7372), .A2(n7373), .ZN(n7371) );
  INV_X1 U7017 ( .A(n5478), .ZN(n5479) );
  NAND2_X1 U7018 ( .A1(n5480), .A2(n5479), .ZN(n5481) );
  NAND2_X1 U7019 ( .A1(n7371), .A2(n5481), .ZN(n5508) );
  INV_X1 U7020 ( .A(n5508), .ZN(n5506) );
  INV_X1 U7021 ( .A(SI_14_), .ZN(n10081) );
  XNOR2_X1 U7022 ( .A(n5482), .B(n10081), .ZN(n5483) );
  XNOR2_X1 U7023 ( .A(n5484), .B(n5483), .ZN(n6644) );
  NAND2_X1 U7024 ( .A1(n6644), .A2(n7590), .ZN(n5493) );
  INV_X1 U7025 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U7026 ( .A1(n5486), .A2(n5485), .ZN(n5487) );
  OAI21_X1 U7027 ( .B1(n5488), .B2(n5487), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5489) );
  MUX2_X1 U7028 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5489), .S(
        P1_IR_REG_14__SCAN_IN), .Z(n5491) );
  AND2_X1 U7029 ( .A1(n5491), .A2(n5490), .ZN(n7099) );
  AOI22_X1 U7030 ( .A1(n5602), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5601), .B2(
        n7099), .ZN(n5492) );
  NAND2_X1 U7031 ( .A1(n7444), .A2(n5325), .ZN(n5503) );
  INV_X1 U7032 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5494) );
  OR2_X1 U7033 ( .A1(n6495), .A2(n5494), .ZN(n5501) );
  INV_X1 U7034 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6748) );
  OR2_X1 U7035 ( .A1(n6488), .A2(n6748), .ZN(n5500) );
  INV_X1 U7036 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5495) );
  NAND2_X1 U7037 ( .A1(n5496), .A2(n5495), .ZN(n5497) );
  AND2_X1 U7038 ( .A1(n5520), .A2(n5497), .ZN(n8869) );
  NAND2_X1 U7039 ( .A1(n5442), .A2(n8869), .ZN(n5499) );
  NAND2_X1 U7040 ( .A1(n6493), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5498) );
  NAND2_X1 U7041 ( .A1(n9033), .A2(n6341), .ZN(n5502) );
  NAND2_X1 U7042 ( .A1(n5503), .A2(n5502), .ZN(n5504) );
  XNOR2_X1 U7043 ( .A(n5504), .B(n5222), .ZN(n5507) );
  INV_X1 U7044 ( .A(n5507), .ZN(n5505) );
  NAND2_X1 U7045 ( .A1(n5506), .A2(n5505), .ZN(n5509) );
  NAND2_X1 U7046 ( .A1(n5508), .A2(n5507), .ZN(n5511) );
  NOR2_X1 U7047 ( .A1(n9671), .A2(n6343), .ZN(n5510) );
  AOI21_X1 U7048 ( .B1(n7444), .B2(n6341), .A(n5510), .ZN(n8863) );
  NAND2_X1 U7049 ( .A1(n8862), .A2(n5511), .ZN(n8923) );
  XNOR2_X1 U7050 ( .A(n5512), .B(SI_15_), .ZN(n5513) );
  XNOR2_X1 U7051 ( .A(n5514), .B(n5513), .ZN(n6683) );
  NAND2_X1 U7052 ( .A1(n6683), .A2(n7590), .ZN(n5517) );
  NAND2_X1 U7053 ( .A1(n5490), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5515) );
  XNOR2_X1 U7054 ( .A(n5515), .B(P1_IR_REG_15__SCAN_IN), .ZN(n7094) );
  AOI22_X1 U7055 ( .A1(n5602), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n5601), .B2(
        n7094), .ZN(n5516) );
  NAND2_X2 U7056 ( .A1(n5517), .A2(n5516), .ZN(n9474) );
  NAND2_X1 U7057 ( .A1(n9474), .A2(n5325), .ZN(n5527) );
  INV_X1 U7058 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7101) );
  OR2_X1 U7059 ( .A1(n6494), .A2(n7101), .ZN(n5525) );
  INV_X1 U7060 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5518) );
  OR2_X1 U7061 ( .A1(n6495), .A2(n5518), .ZN(n5524) );
  NAND2_X1 U7062 ( .A1(n5725), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5523) );
  INV_X1 U7063 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U7064 ( .A1(n5520), .A2(n5519), .ZN(n5521) );
  AND2_X1 U7065 ( .A1(n5539), .A2(n5521), .ZN(n9023) );
  NAND2_X1 U7066 ( .A1(n5442), .A2(n9023), .ZN(n5522) );
  NAND2_X1 U7067 ( .A1(n9032), .A2(n6341), .ZN(n5526) );
  NAND2_X1 U7068 ( .A1(n5527), .A2(n5526), .ZN(n5528) );
  XNOR2_X1 U7069 ( .A(n5528), .B(n5222), .ZN(n5550) );
  NOR2_X1 U7070 ( .A1(n8934), .A2(n6343), .ZN(n5529) );
  AOI21_X1 U7071 ( .B1(n9474), .B2(n6341), .A(n5529), .ZN(n9015) );
  AND2_X1 U7072 ( .A1(n5550), .A2(n9015), .ZN(n5554) );
  INV_X1 U7073 ( .A(SI_16_), .ZN(n10123) );
  XNOR2_X1 U7074 ( .A(n5530), .B(n10123), .ZN(n5531) );
  NAND2_X1 U7075 ( .A1(n6690), .A2(n7590), .ZN(n5536) );
  NAND2_X1 U7076 ( .A1(n5533), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5534) );
  XNOR2_X1 U7077 ( .A(n5534), .B(P1_IR_REG_16__SCAN_IN), .ZN(n7287) );
  AOI22_X1 U7078 ( .A1(n5602), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5601), .B2(
        n7287), .ZN(n5535) );
  NAND2_X1 U7079 ( .A1(n9468), .A2(n5361), .ZN(n5546) );
  NAND2_X1 U7080 ( .A1(n5160), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5544) );
  INV_X1 U7081 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n5537) );
  OR2_X1 U7082 ( .A1(n6488), .A2(n5537), .ZN(n5543) );
  NAND2_X1 U7083 ( .A1(n5539), .A2(n5538), .ZN(n5540) );
  AND2_X1 U7084 ( .A1(n5566), .A2(n5540), .ZN(n8938) );
  NAND2_X1 U7085 ( .A1(n5442), .A2(n8938), .ZN(n5542) );
  NAND2_X1 U7086 ( .A1(n5725), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5541) );
  NAND2_X1 U7087 ( .A1(n9031), .A2(n6341), .ZN(n5545) );
  NAND2_X1 U7088 ( .A1(n5546), .A2(n5545), .ZN(n5547) );
  XNOR2_X1 U7089 ( .A(n5547), .B(n5752), .ZN(n5555) );
  NAND2_X1 U7090 ( .A1(n9468), .A2(n6341), .ZN(n5549) );
  NAND2_X1 U7091 ( .A1(n9031), .A2(n5174), .ZN(n5548) );
  NAND2_X1 U7092 ( .A1(n5549), .A2(n5548), .ZN(n5556) );
  NAND2_X1 U7093 ( .A1(n5555), .A2(n5556), .ZN(n8929) );
  INV_X1 U7094 ( .A(n8929), .ZN(n5552) );
  INV_X1 U7095 ( .A(n5550), .ZN(n8924) );
  INV_X1 U7096 ( .A(n9015), .ZN(n5551) );
  INV_X1 U7097 ( .A(n5555), .ZN(n5558) );
  INV_X1 U7098 ( .A(n5556), .ZN(n5557) );
  NAND2_X1 U7099 ( .A1(n5558), .A2(n5557), .ZN(n8928) );
  NAND2_X1 U7100 ( .A1(n5559), .A2(n8928), .ZN(n8941) );
  XNOR2_X1 U7101 ( .A(n5561), .B(n5560), .ZN(n6846) );
  NAND2_X1 U7102 ( .A1(n6846), .A2(n7590), .ZN(n5564) );
  XNOR2_X1 U7103 ( .A(n5562), .B(P1_IR_REG_17__SCAN_IN), .ZN(n7833) );
  AOI22_X1 U7104 ( .A1(n5602), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5601), .B2(
        n7833), .ZN(n5563) );
  NAND2_X1 U7105 ( .A1(n9463), .A2(n5325), .ZN(n5573) );
  INV_X1 U7106 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5565) );
  NAND2_X1 U7107 ( .A1(n5566), .A2(n5565), .ZN(n5567) );
  NAND2_X1 U7108 ( .A1(n5586), .A2(n5567), .ZN(n9350) );
  OR2_X1 U7109 ( .A1(n5647), .A2(n9350), .ZN(n5571) );
  NAND2_X1 U7110 ( .A1(n5160), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n5570) );
  INV_X1 U7111 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n7827) );
  OR2_X1 U7112 ( .A1(n6494), .A2(n7827), .ZN(n5569) );
  NAND2_X1 U7113 ( .A1(n6493), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7114 ( .A1(n9030), .A2(n6341), .ZN(n5572) );
  NAND2_X1 U7115 ( .A1(n5573), .A2(n5572), .ZN(n5574) );
  XNOR2_X1 U7116 ( .A(n5574), .B(n5222), .ZN(n8943) );
  NOR2_X1 U7117 ( .A1(n9329), .A2(n6343), .ZN(n5575) );
  AOI21_X1 U7118 ( .B1(n9463), .B2(n6341), .A(n5575), .ZN(n8942) );
  INV_X1 U7119 ( .A(n8943), .ZN(n5577) );
  INV_X1 U7120 ( .A(n8942), .ZN(n5576) );
  NAND2_X1 U7121 ( .A1(n5577), .A2(n5576), .ZN(n5578) );
  XNOR2_X1 U7122 ( .A(n5580), .B(n5579), .ZN(n6952) );
  NAND2_X1 U7123 ( .A1(n6952), .A2(n7590), .ZN(n5584) );
  NAND2_X1 U7124 ( .A1(n5581), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5582) );
  XNOR2_X1 U7125 ( .A(n5582), .B(P1_IR_REG_18__SCAN_IN), .ZN(n7836) );
  AOI22_X1 U7126 ( .A1(n5602), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5601), .B2(
        n7836), .ZN(n5583) );
  NAND2_X1 U7127 ( .A1(n9337), .A2(n5325), .ZN(n5592) );
  NAND2_X1 U7128 ( .A1(n5586), .A2(n5585), .ZN(n5587) );
  AND2_X1 U7129 ( .A1(n5606), .A2(n5587), .ZN(n9338) );
  NAND2_X1 U7130 ( .A1(n9338), .A2(n5442), .ZN(n5590) );
  INV_X1 U7131 ( .A(n6488), .ZN(n5608) );
  AOI22_X1 U7132 ( .A1(n5608), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n5160), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5589) );
  NAND2_X1 U7133 ( .A1(n5725), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7134 ( .A1(n9313), .A2(n6341), .ZN(n5591) );
  NAND2_X1 U7135 ( .A1(n5592), .A2(n5591), .ZN(n5593) );
  XNOR2_X1 U7136 ( .A(n5593), .B(n5752), .ZN(n5595) );
  INV_X1 U7137 ( .A(n5595), .ZN(n5594) );
  NOR2_X1 U7138 ( .A1(n9357), .A2(n6343), .ZN(n5597) );
  AOI21_X1 U7139 ( .B1(n9337), .B2(n6341), .A(n5597), .ZN(n8995) );
  XNOR2_X1 U7140 ( .A(n5600), .B(n5599), .ZN(n7070) );
  NAND2_X1 U7141 ( .A1(n7070), .A2(n7590), .ZN(n5604) );
  AOI22_X1 U7142 ( .A1(n5602), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7844), .B2(
        n5601), .ZN(n5603) );
  NAND2_X1 U7143 ( .A1(n9453), .A2(n5361), .ZN(n5613) );
  INV_X1 U7144 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5605) );
  NAND2_X1 U7145 ( .A1(n5606), .A2(n5605), .ZN(n5607) );
  NAND2_X1 U7146 ( .A1(n5625), .A2(n5607), .ZN(n9317) );
  OR2_X1 U7147 ( .A1(n9317), .A2(n5647), .ZN(n5611) );
  AOI22_X1 U7148 ( .A1(n5608), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n5160), .B2(
        P1_REG0_REG_19__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U7149 ( .A1(n6493), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7150 ( .A1(n9440), .A2(n6341), .ZN(n5612) );
  NAND2_X1 U7151 ( .A1(n5613), .A2(n5612), .ZN(n5614) );
  XNOR2_X1 U7152 ( .A(n5614), .B(n5752), .ZN(n5616) );
  NOR2_X1 U7153 ( .A1(n9330), .A2(n6343), .ZN(n5615) );
  AOI21_X1 U7154 ( .B1(n9453), .B2(n6341), .A(n5615), .ZN(n5617) );
  XNOR2_X1 U7155 ( .A(n5616), .B(n5617), .ZN(n8900) );
  INV_X1 U7156 ( .A(n5616), .ZN(n5618) );
  NAND2_X1 U7157 ( .A1(n5618), .A2(n5617), .ZN(n5619) );
  XNOR2_X1 U7158 ( .A(n5620), .B(n10126), .ZN(n5621) );
  XNOR2_X1 U7159 ( .A(n5622), .B(n5621), .ZN(n7143) );
  NAND2_X1 U7160 ( .A1(n7143), .A2(n7590), .ZN(n5624) );
  INV_X1 U7161 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7153) );
  OR2_X1 U7162 ( .A1(n7596), .A2(n7153), .ZN(n5623) );
  NAND2_X1 U7163 ( .A1(n9303), .A2(n5325), .ZN(n5634) );
  NAND2_X1 U7164 ( .A1(n5625), .A2(n8976), .ZN(n5626) );
  AND2_X1 U7165 ( .A1(n5645), .A2(n5626), .ZN(n9297) );
  NAND2_X1 U7166 ( .A1(n9297), .A2(n5442), .ZN(n5632) );
  INV_X1 U7167 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5629) );
  NAND2_X1 U7168 ( .A1(n5160), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5628) );
  NAND2_X1 U7169 ( .A1(n5725), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5627) );
  OAI211_X1 U7170 ( .C1(n6494), .C2(n5629), .A(n5628), .B(n5627), .ZN(n5630)
         );
  INV_X1 U7171 ( .A(n5630), .ZN(n5631) );
  OR2_X1 U7172 ( .A1(n9316), .A2(n6337), .ZN(n5633) );
  NAND2_X1 U7173 ( .A1(n5634), .A2(n5633), .ZN(n5635) );
  XNOR2_X1 U7174 ( .A(n5635), .B(n5222), .ZN(n5638) );
  NOR2_X1 U7175 ( .A1(n9316), .A2(n6343), .ZN(n5636) );
  AOI21_X1 U7176 ( .B1(n9303), .B2(n6341), .A(n5636), .ZN(n5637) );
  AND2_X1 U7177 ( .A1(n5638), .A2(n5637), .ZN(n8972) );
  INV_X1 U7178 ( .A(SI_21_), .ZN(n10170) );
  XNOR2_X1 U7179 ( .A(n5639), .B(n10170), .ZN(n5640) );
  XNOR2_X1 U7180 ( .A(n5641), .B(n5640), .ZN(n7178) );
  NAND2_X1 U7181 ( .A1(n7178), .A2(n7590), .ZN(n5643) );
  INV_X1 U7182 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n7179) );
  OR2_X1 U7183 ( .A1(n7596), .A2(n7179), .ZN(n5642) );
  NAND2_X1 U7184 ( .A1(n9287), .A2(n5325), .ZN(n5655) );
  INV_X1 U7185 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n5644) );
  NAND2_X1 U7186 ( .A1(n5645), .A2(n5644), .ZN(n5646) );
  NAND2_X1 U7187 ( .A1(n5676), .A2(n5646), .ZN(n8911) );
  OR2_X1 U7188 ( .A1(n8911), .A2(n5647), .ZN(n5653) );
  INV_X1 U7189 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5650) );
  NAND2_X1 U7190 ( .A1(n5160), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5649) );
  NAND2_X1 U7191 ( .A1(n6493), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5648) );
  OAI211_X1 U7192 ( .C1(n6488), .C2(n5650), .A(n5649), .B(n5648), .ZN(n5651)
         );
  INV_X1 U7193 ( .A(n5651), .ZN(n5652) );
  OR2_X1 U7194 ( .A1(n9301), .A2(n6337), .ZN(n5654) );
  NAND2_X1 U7195 ( .A1(n5655), .A2(n5654), .ZN(n5656) );
  XNOR2_X1 U7196 ( .A(n5656), .B(n5752), .ZN(n5658) );
  NOR2_X1 U7197 ( .A1(n9301), .A2(n6343), .ZN(n5657) );
  AOI21_X1 U7198 ( .B1(n9287), .B2(n5775), .A(n5657), .ZN(n5659) );
  XNOR2_X1 U7199 ( .A(n5658), .B(n5659), .ZN(n8909) );
  INV_X1 U7200 ( .A(n5658), .ZN(n5660) );
  NAND2_X1 U7201 ( .A1(n9266), .A2(n5361), .ZN(n5662) );
  OR2_X1 U7202 ( .A1(n9417), .A2(n6337), .ZN(n5661) );
  NAND2_X1 U7203 ( .A1(n5662), .A2(n5661), .ZN(n5663) );
  XNOR2_X1 U7204 ( .A(n5663), .B(n5222), .ZN(n5664) );
  NOR2_X1 U7205 ( .A1(n5665), .A2(n5664), .ZN(n8981) );
  INV_X1 U7206 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7370) );
  MUX2_X1 U7207 ( .A(n7366), .B(n7370), .S(n4611), .Z(n5670) );
  INV_X1 U7208 ( .A(SI_23_), .ZN(n5669) );
  NAND2_X1 U7209 ( .A1(n5670), .A2(n5669), .ZN(n5692) );
  INV_X1 U7210 ( .A(n5670), .ZN(n5671) );
  NAND2_X1 U7211 ( .A1(n5671), .A2(SI_23_), .ZN(n5672) );
  XNOR2_X1 U7212 ( .A(n5691), .B(n5690), .ZN(n7368) );
  NAND2_X1 U7213 ( .A1(n7368), .A2(n7590), .ZN(n5674) );
  OR2_X1 U7214 ( .A1(n7596), .A2(n7370), .ZN(n5673) );
  INV_X1 U7215 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8987) );
  INV_X1 U7216 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n8877) );
  OAI21_X1 U7217 ( .B1(n5676), .B2(n8987), .A(n8877), .ZN(n5677) );
  NAND2_X1 U7218 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n5675) );
  NAND2_X1 U7219 ( .A1(n5677), .A2(n5701), .ZN(n8879) );
  OR2_X1 U7220 ( .A1(n8879), .A2(n5647), .ZN(n5682) );
  INV_X1 U7221 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n9422) );
  NAND2_X1 U7222 ( .A1(n5160), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5679) );
  NAND2_X1 U7223 ( .A1(n6493), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5678) );
  OAI211_X1 U7224 ( .C1(n6488), .C2(n9422), .A(n5679), .B(n5678), .ZN(n5680)
         );
  INV_X1 U7225 ( .A(n5680), .ZN(n5681) );
  NAND2_X1 U7226 ( .A1(n5682), .A2(n5681), .ZN(n9424) );
  OAI22_X1 U7227 ( .A1(n9507), .A2(n5683), .B1(n9270), .B2(n6337), .ZN(n5684)
         );
  XNOR2_X1 U7228 ( .A(n5684), .B(n5222), .ZN(n5689) );
  INV_X1 U7229 ( .A(n5689), .ZN(n5687) );
  AND2_X1 U7230 ( .A1(n9424), .A2(n5174), .ZN(n5685) );
  AOI21_X1 U7231 ( .B1(n9260), .B2(n6341), .A(n5685), .ZN(n5688) );
  INV_X1 U7232 ( .A(n5688), .ZN(n5686) );
  NAND2_X1 U7233 ( .A1(n5687), .A2(n5686), .ZN(n8873) );
  AND2_X1 U7234 ( .A1(n5689), .A2(n5688), .ZN(n8874) );
  INV_X1 U7235 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7475) );
  MUX2_X1 U7236 ( .A(n7475), .B(n7495), .S(n7550), .Z(n5694) );
  INV_X1 U7237 ( .A(SI_24_), .ZN(n10167) );
  NAND2_X1 U7238 ( .A1(n5694), .A2(n10167), .ZN(n5717) );
  INV_X1 U7239 ( .A(n5694), .ZN(n5695) );
  NAND2_X1 U7240 ( .A1(n5695), .A2(SI_24_), .ZN(n5696) );
  XNOR2_X1 U7241 ( .A(n5716), .B(n5715), .ZN(n7474) );
  NAND2_X1 U7242 ( .A1(n7474), .A2(n7590), .ZN(n5698) );
  OR2_X1 U7243 ( .A1(n7596), .A2(n7495), .ZN(n5697) );
  NAND2_X1 U7244 ( .A1(n9243), .A2(n5361), .ZN(n5709) );
  INV_X1 U7245 ( .A(n5701), .ZN(n5699) );
  NAND2_X1 U7246 ( .A1(n5699), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n5723) );
  INV_X1 U7247 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5700) );
  NAND2_X1 U7248 ( .A1(n5701), .A2(n5700), .ZN(n5702) );
  NAND2_X1 U7249 ( .A1(n5723), .A2(n5702), .ZN(n9244) );
  OR2_X1 U7250 ( .A1(n9244), .A2(n5647), .ZN(n5707) );
  INV_X1 U7251 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n9412) );
  NAND2_X1 U7252 ( .A1(n5160), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5704) );
  NAND2_X1 U7253 ( .A1(n6493), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5703) );
  OAI211_X1 U7254 ( .C1(n6494), .C2(n9412), .A(n5704), .B(n5703), .ZN(n5705)
         );
  INV_X1 U7255 ( .A(n5705), .ZN(n5706) );
  NAND2_X1 U7256 ( .A1(n9414), .A2(n6341), .ZN(n5708) );
  NAND2_X1 U7257 ( .A1(n5709), .A2(n5708), .ZN(n5710) );
  XNOR2_X1 U7258 ( .A(n5710), .B(n5222), .ZN(n5713) );
  NOR2_X1 U7259 ( .A1(n9258), .A2(n6343), .ZN(n5711) );
  AOI21_X1 U7260 ( .B1(n9243), .B2(n5775), .A(n5711), .ZN(n5712) );
  NAND2_X1 U7261 ( .A1(n5713), .A2(n5712), .ZN(n5714) );
  OAI21_X1 U7262 ( .B1(n5713), .B2(n5712), .A(n5714), .ZN(n8952) );
  INV_X1 U7263 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7517) );
  INV_X1 U7264 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7521) );
  MUX2_X1 U7265 ( .A(n7517), .B(n7521), .S(n7550), .Z(n5718) );
  INV_X1 U7266 ( .A(SI_25_), .ZN(n10165) );
  NAND2_X1 U7267 ( .A1(n5718), .A2(n10165), .ZN(n5736) );
  INV_X1 U7268 ( .A(n5718), .ZN(n5719) );
  NAND2_X1 U7269 ( .A1(n5719), .A2(SI_25_), .ZN(n5720) );
  XNOR2_X1 U7270 ( .A(n5735), .B(n5734), .ZN(n7516) );
  NAND2_X1 U7271 ( .A1(n7516), .A2(n7590), .ZN(n5722) );
  OR2_X1 U7272 ( .A1(n7596), .A2(n7521), .ZN(n5721) );
  NAND2_X1 U7273 ( .A1(n9231), .A2(n5361), .ZN(n5732) );
  INV_X1 U7274 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8917) );
  NAND2_X1 U7275 ( .A1(n5723), .A2(n8917), .ZN(n5724) );
  NAND2_X1 U7276 ( .A1(n5742), .A2(n5724), .ZN(n9226) );
  INV_X1 U7277 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n9407) );
  NAND2_X1 U7278 ( .A1(n5160), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5727) );
  NAND2_X1 U7279 ( .A1(n5725), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5726) );
  OAI211_X1 U7280 ( .C1(n6488), .C2(n9407), .A(n5727), .B(n5726), .ZN(n5728)
         );
  INV_X1 U7281 ( .A(n5728), .ZN(n5729) );
  NAND2_X1 U7282 ( .A1(n9211), .A2(n6341), .ZN(n5731) );
  NAND2_X1 U7283 ( .A1(n5732), .A2(n5731), .ZN(n5733) );
  XNOR2_X1 U7284 ( .A(n5733), .B(n5752), .ZN(n5755) );
  OAI22_X1 U7285 ( .A1(n9499), .A2(n6337), .B1(n9390), .B2(n6343), .ZN(n5754)
         );
  XNOR2_X1 U7286 ( .A(n5755), .B(n5754), .ZN(n8916) );
  INV_X1 U7287 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7523) );
  INV_X1 U7288 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7527) );
  MUX2_X1 U7289 ( .A(n7523), .B(n7527), .S(n7550), .Z(n5737) );
  NAND2_X1 U7290 ( .A1(n5737), .A2(n10143), .ZN(n5762) );
  INV_X1 U7291 ( .A(n5737), .ZN(n5738) );
  NAND2_X1 U7292 ( .A1(n5738), .A2(SI_26_), .ZN(n5739) );
  NAND2_X1 U7293 ( .A1(n7522), .A2(n7590), .ZN(n5741) );
  OR2_X1 U7294 ( .A1(n7596), .A2(n7527), .ZN(n5740) );
  INV_X1 U7295 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n9007) );
  NAND2_X1 U7296 ( .A1(n5742), .A2(n9007), .ZN(n5743) );
  NAND2_X1 U7297 ( .A1(n9210), .A2(n5442), .ZN(n5748) );
  INV_X1 U7298 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n9398) );
  NAND2_X1 U7299 ( .A1(n5160), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5745) );
  NAND2_X1 U7300 ( .A1(n6493), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n5744) );
  OAI211_X1 U7301 ( .C1(n6494), .C2(n9398), .A(n5745), .B(n5744), .ZN(n5746)
         );
  INV_X1 U7302 ( .A(n5746), .ZN(n5747) );
  NOR2_X1 U7303 ( .A1(n9402), .A2(n6343), .ZN(n5749) );
  AOI21_X1 U7304 ( .B1(n9209), .B2(n6341), .A(n5749), .ZN(n5757) );
  NAND2_X1 U7305 ( .A1(n9209), .A2(n5361), .ZN(n5751) );
  NAND2_X1 U7306 ( .A1(n9194), .A2(n6341), .ZN(n5750) );
  NAND2_X1 U7307 ( .A1(n5751), .A2(n5750), .ZN(n5753) );
  XNOR2_X1 U7308 ( .A(n5753), .B(n5752), .ZN(n5759) );
  XOR2_X1 U7309 ( .A(n5757), .B(n5759), .Z(n9002) );
  NOR2_X1 U7310 ( .A1(n5755), .A2(n5754), .ZN(n9003) );
  INV_X1 U7311 ( .A(n5757), .ZN(n5758) );
  INV_X1 U7312 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8859) );
  INV_X1 U7313 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n7529) );
  MUX2_X1 U7314 ( .A(n8859), .B(n7529), .S(n7550), .Z(n5765) );
  INV_X1 U7315 ( .A(SI_27_), .ZN(n5764) );
  NAND2_X1 U7316 ( .A1(n5765), .A2(n5764), .ZN(n6189) );
  INV_X1 U7317 ( .A(n5765), .ZN(n5766) );
  NAND2_X1 U7318 ( .A1(n5766), .A2(SI_27_), .ZN(n5767) );
  NAND2_X1 U7319 ( .A1(n7528), .A2(n7590), .ZN(n5769) );
  OR2_X1 U7320 ( .A1(n7596), .A2(n7529), .ZN(n5768) );
  NAND2_X1 U7321 ( .A1(n9193), .A2(n5361), .ZN(n5777) );
  XNOR2_X1 U7322 ( .A(n5820), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9195) );
  NAND2_X1 U7323 ( .A1(n9195), .A2(n5442), .ZN(n5774) );
  INV_X1 U7324 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n9388) );
  NAND2_X1 U7325 ( .A1(n5160), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5771) );
  NAND2_X1 U7326 ( .A1(n6493), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5770) );
  OAI211_X1 U7327 ( .C1(n6488), .C2(n9388), .A(n5771), .B(n5770), .ZN(n5772)
         );
  INV_X1 U7328 ( .A(n5772), .ZN(n5773) );
  INV_X1 U7329 ( .A(n9391), .ZN(n9029) );
  NAND2_X1 U7330 ( .A1(n9029), .A2(n5775), .ZN(n5776) );
  NAND2_X1 U7331 ( .A1(n5777), .A2(n5776), .ZN(n5778) );
  XNOR2_X1 U7332 ( .A(n5778), .B(n5222), .ZN(n5781) );
  NOR2_X1 U7333 ( .A1(n9391), .A2(n6343), .ZN(n5779) );
  AOI21_X1 U7334 ( .B1(n9193), .B2(n6341), .A(n5779), .ZN(n5780) );
  NAND2_X1 U7335 ( .A1(n5781), .A2(n5780), .ZN(n6355) );
  OAI21_X1 U7336 ( .B1(n5781), .B2(n5780), .A(n6355), .ZN(n5783) );
  INV_X1 U7337 ( .A(n5784), .ZN(n5808) );
  NAND2_X1 U7338 ( .A1(n7520), .A2(P1_B_REG_SCAN_IN), .ZN(n5785) );
  MUX2_X1 U7339 ( .A(n5785), .B(P1_B_REG_SCAN_IN), .S(n7492), .Z(n5786) );
  AND2_X1 U7340 ( .A1(n5786), .A2(n5799), .ZN(n6516) );
  INV_X1 U7341 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n5787) );
  NAND2_X1 U7342 ( .A1(n6516), .A2(n5787), .ZN(n5788) );
  INV_X1 U7343 ( .A(n6516), .ZN(n5800) );
  NOR4_X1 U7344 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5792) );
  NOR4_X1 U7345 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n5791) );
  NOR4_X1 U7346 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5790) );
  NOR4_X1 U7347 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5789) );
  NAND4_X1 U7348 ( .A1(n5792), .A2(n5791), .A3(n5790), .A4(n5789), .ZN(n5798)
         );
  NOR2_X1 U7349 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n5796) );
  NOR4_X1 U7350 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n5795) );
  NOR4_X1 U7351 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n5794) );
  NOR4_X1 U7352 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n5793) );
  NAND4_X1 U7353 ( .A1(n5796), .A2(n5795), .A3(n5794), .A4(n5793), .ZN(n5797)
         );
  NOR2_X1 U7354 ( .A1(n5798), .A2(n5797), .ZN(n6514) );
  AND2_X1 U7355 ( .A1(n6514), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6663) );
  INV_X1 U7356 ( .A(n5799), .ZN(n7526) );
  NAND2_X1 U7357 ( .A1(n7526), .A2(n7520), .ZN(n6666) );
  OAI21_X1 U7358 ( .B1(n5800), .B2(n6663), .A(n6666), .ZN(n5801) );
  OR2_X1 U7359 ( .A1(n6668), .A2(n5801), .ZN(n5812) );
  NAND2_X1 U7360 ( .A1(n5804), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6363) );
  NAND2_X1 U7361 ( .A1(n7804), .A2(n7756), .ZN(n6673) );
  AND2_X1 U7362 ( .A1(n9664), .A2(n7599), .ZN(n5807) );
  OAI21_X1 U7363 ( .B1(n6358), .B2(n5808), .A(n9016), .ZN(n5834) );
  INV_X1 U7364 ( .A(n5809), .ZN(n5828) );
  OR2_X1 U7365 ( .A1(n6673), .A2(n7801), .ZN(n6679) );
  OR2_X1 U7366 ( .A1(n5828), .A2(n6679), .ZN(n5810) );
  INV_X1 U7367 ( .A(n7807), .ZN(n6664) );
  OR2_X1 U7368 ( .A1(n7810), .A2(n6548), .ZN(n9634) );
  INV_X1 U7369 ( .A(n6512), .ZN(n5811) );
  NAND2_X1 U7370 ( .A1(n5812), .A2(n5811), .ZN(n5813) );
  INV_X1 U7371 ( .A(n7599), .ZN(n6521) );
  NAND2_X1 U7372 ( .A1(n6521), .A2(n6522), .ZN(n6667) );
  NAND2_X1 U7373 ( .A1(n5813), .A2(n6667), .ZN(n6617) );
  OAI21_X1 U7374 ( .B1(n6617), .B2(n5169), .A(P1_STATE_REG_SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7375 ( .A1(n6473), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7819) );
  NOR2_X2 U7376 ( .A1(n7599), .A2(n4353), .ZN(n9647) );
  INV_X1 U7377 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5819) );
  OAI22_X1 U7378 ( .A1(n9402), .A2(n8988), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n5819), .ZN(n5830) );
  INV_X1 U7379 ( .A(n5820), .ZN(n5817) );
  AND2_X1 U7380 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5816) );
  NAND2_X1 U7381 ( .A1(n5817), .A2(n5816), .ZN(n7978) );
  INV_X1 U7382 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5818) );
  OAI21_X1 U7383 ( .B1(n5820), .B2(n5819), .A(n5818), .ZN(n5821) );
  NAND2_X1 U7384 ( .A1(n9178), .A2(n5442), .ZN(n5827) );
  INV_X1 U7385 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7386 ( .A1(n5160), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5823) );
  NAND2_X1 U7387 ( .A1(n6493), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n5822) );
  OAI211_X1 U7388 ( .C1(n6488), .C2(n5824), .A(n5823), .B(n5822), .ZN(n5825)
         );
  INV_X1 U7389 ( .A(n5825), .ZN(n5826) );
  NOR2_X1 U7390 ( .A1(n9381), .A2(n9008), .ZN(n5829) );
  AOI211_X1 U7391 ( .C1(n9195), .C2(n9022), .A(n5830), .B(n5829), .ZN(n5831)
         );
  OAI21_X1 U7392 ( .B1(n9491), .B2(n9026), .A(n5831), .ZN(n5832) );
  INV_X1 U7393 ( .A(n5832), .ZN(n5833) );
  NAND2_X1 U7394 ( .A1(n5834), .A2(n5833), .ZN(P1_U3214) );
  NAND2_X1 U7395 ( .A1(n5853), .A2(n5851), .ZN(n7563) );
  NAND2_X1 U7396 ( .A1(n7563), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5852) );
  XNOR2_X1 U7397 ( .A(n5852), .B(n7560), .ZN(n5855) );
  INV_X1 U7398 ( .A(n5855), .ZN(n5869) );
  INV_X1 U7399 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6431) );
  NAND2_X1 U7400 ( .A1(n5899), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5867) );
  INV_X1 U7401 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n7996) );
  NOR2_X1 U7402 ( .A1(n5857), .A2(n7996), .ZN(n5856) );
  NAND2_X1 U7403 ( .A1(n5869), .A2(n5856), .ZN(n5865) );
  INV_X1 U7404 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5858) );
  XNOR2_X2 U7405 ( .A(n5861), .B(n5860), .ZN(n6273) );
  XNOR2_X2 U7406 ( .A(n5862), .B(n5850), .ZN(n6274) );
  NAND2_X4 U7407 ( .A1(n6273), .A2(n6274), .ZN(n6281) );
  INV_X1 U7408 ( .A(n6437), .ZN(n5863) );
  INV_X1 U7409 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6466) );
  NAND4_X1 U7410 ( .A1(n5867), .A2(n5866), .A3(n5865), .A4(n5864), .ZN(n8410)
         );
  NAND2_X1 U7411 ( .A1(n8410), .A2(n9912), .ZN(n8183) );
  INV_X2 U7412 ( .A(n5914), .ZN(n6202) );
  NAND2_X1 U7413 ( .A1(n6202), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n6224) );
  INV_X1 U7414 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5868) );
  INV_X1 U7415 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n5870) );
  OR2_X1 U7416 ( .A1(n5903), .A2(n5870), .ZN(n6222) );
  INV_X1 U7417 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5871) );
  OR2_X1 U7418 ( .A1(n5878), .A2(n5871), .ZN(n6221) );
  NAND2_X1 U7419 ( .A1(n6452), .A2(SI_0_), .ZN(n5873) );
  INV_X1 U7420 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U7421 ( .A1(n5873), .A2(n5872), .ZN(n5875) );
  AND2_X1 U7422 ( .A1(n5875), .A2(n5874), .ZN(n8861) );
  MUX2_X1 U7423 ( .A(P2_IR_REG_0__SCAN_IN), .B(n8861), .S(n6281), .Z(n6832) );
  NAND2_X1 U7424 ( .A1(n6687), .A2(n6832), .ZN(n8187) );
  OR2_X1 U7425 ( .A1(n8343), .A2(n8187), .ZN(n7988) );
  NAND2_X1 U7426 ( .A1(n5899), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5883) );
  INV_X1 U7427 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n5877) );
  OR2_X1 U7428 ( .A1(n5878), .A2(n5877), .ZN(n5882) );
  INV_X1 U7429 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6908) );
  INV_X1 U7430 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n5879) );
  OR2_X1 U7431 ( .A1(n5914), .A2(n5879), .ZN(n5880) );
  AND4_X2 U7432 ( .A1(n5883), .A2(n5882), .A3(n5881), .A4(n5880), .ZN(n7991)
         );
  INV_X1 U7433 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6451) );
  OR2_X1 U7434 ( .A1(n8320), .A2(n6451), .ZN(n5886) );
  OR2_X1 U7435 ( .A1(n8321), .A2(n6453), .ZN(n5885) );
  OAI211_X1 U7436 ( .C1(n6281), .C2(n7062), .A(n5886), .B(n5885), .ZN(n6373)
         );
  NAND2_X1 U7437 ( .A1(n7991), .A2(n6373), .ZN(n8193) );
  NAND2_X1 U7438 ( .A1(n9890), .A2(n9897), .ZN(n5887) );
  NAND2_X1 U7439 ( .A1(n5887), .A2(n8193), .ZN(n6967) );
  NAND2_X1 U7440 ( .A1(n6999), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5893) );
  INV_X1 U7441 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n5888) );
  INV_X1 U7442 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n5889) );
  OR2_X1 U7443 ( .A1(n5878), .A2(n5889), .ZN(n5891) );
  OR2_X1 U7444 ( .A1(n5914), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7445 ( .A1(n5884), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5894) );
  MUX2_X1 U7446 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5894), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n5895) );
  OR2_X1 U7447 ( .A1(n8320), .A2(n4466), .ZN(n5897) );
  OR2_X1 U7448 ( .A1(n8321), .A2(n6455), .ZN(n5896) );
  OAI211_X1 U7449 ( .C1(n6281), .C2(n6992), .A(n5897), .B(n5896), .ZN(n9920)
         );
  XNOR2_X1 U7450 ( .A(n9881), .B(n9920), .ZN(n8347) );
  NAND2_X1 U7451 ( .A1(n6967), .A2(n8347), .ZN(n5898) );
  NAND2_X1 U7452 ( .A1(n9894), .A2(n9920), .ZN(n8200) );
  NAND2_X1 U7453 ( .A1(n5898), .A2(n8200), .ZN(n9885) );
  NAND2_X1 U7454 ( .A1(n6019), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5907) );
  INV_X2 U7455 ( .A(n5899), .ZN(n6109) );
  INV_X1 U7456 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6973) );
  OR2_X1 U7457 ( .A1(n6109), .A2(n6973), .ZN(n5906) );
  INV_X1 U7458 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n5901) );
  INV_X1 U7459 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5900) );
  NAND2_X1 U7460 ( .A1(n5901), .A2(n5900), .ZN(n5925) );
  NAND2_X1 U7461 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5902) );
  AND2_X1 U7462 ( .A1(n5925), .A2(n5902), .ZN(n9886) );
  OR2_X1 U7463 ( .A1(n5914), .A2(n9886), .ZN(n5905) );
  INV_X1 U7464 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6980) );
  OR2_X1 U7465 ( .A1(n7003), .A2(n6980), .ZN(n5904) );
  NAND4_X1 U7466 ( .A1(n5907), .A2(n5906), .A3(n5905), .A4(n5904), .ZN(n8202)
         );
  NAND2_X1 U7467 ( .A1(n5920), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5909) );
  INV_X1 U7468 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5908) );
  XNOR2_X1 U7469 ( .A(n5909), .B(n5908), .ZN(n7135) );
  OR2_X1 U7470 ( .A1(n8320), .A2(n6459), .ZN(n5911) );
  OR2_X1 U7471 ( .A1(n8321), .A2(n6458), .ZN(n5910) );
  OAI211_X1 U7472 ( .C1(n6281), .C2(n7135), .A(n5911), .B(n5910), .ZN(n9924)
         );
  XNOR2_X1 U7473 ( .A(n8202), .B(n9924), .ZN(n9884) );
  NAND2_X1 U7474 ( .A1(n9885), .A2(n9884), .ZN(n5912) );
  INV_X1 U7475 ( .A(n8202), .ZN(n7168) );
  NAND2_X1 U7476 ( .A1(n7168), .A2(n9924), .ZN(n8210) );
  NAND2_X1 U7477 ( .A1(n5912), .A2(n8210), .ZN(n7167) );
  NAND2_X1 U7478 ( .A1(n6019), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5919) );
  INV_X1 U7479 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n5913) );
  OR2_X1 U7480 ( .A1(n6109), .A2(n5913), .ZN(n5918) );
  INV_X1 U7481 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10168) );
  XNOR2_X1 U7482 ( .A(n5925), .B(n10168), .ZN(n7173) );
  OR2_X1 U7483 ( .A1(n5914), .A2(n7173), .ZN(n5917) );
  INV_X1 U7484 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5915) );
  OR2_X1 U7485 ( .A1(n7003), .A2(n5915), .ZN(n5916) );
  NAND4_X1 U7486 ( .A1(n5919), .A2(n5918), .A3(n5917), .A4(n5916), .ZN(n9879)
         );
  INV_X1 U7487 ( .A(n9879), .ZN(n7026) );
  OR2_X1 U7488 ( .A1(n5920), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n5934) );
  NAND2_X1 U7489 ( .A1(n5934), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5922) );
  XNOR2_X1 U7490 ( .A(n5922), .B(n5921), .ZN(n7231) );
  OR2_X1 U7491 ( .A1(n8321), .A2(n6461), .ZN(n5924) );
  OR2_X1 U7492 ( .A1(n8320), .A2(n6462), .ZN(n5923) );
  OAI211_X1 U7493 ( .C1(n6281), .C2(n7231), .A(n5924), .B(n5923), .ZN(n6378)
         );
  NAND2_X1 U7494 ( .A1(n7026), .A2(n6378), .ZN(n8209) );
  INV_X1 U7495 ( .A(n6378), .ZN(n9929) );
  NAND2_X1 U7496 ( .A1(n9879), .A2(n9929), .ZN(n8213) );
  NAND2_X1 U7497 ( .A1(n7167), .A2(n7166), .ZN(n7165) );
  NAND2_X1 U7498 ( .A1(n7165), .A2(n8209), .ZN(n7290) );
  NAND2_X1 U7499 ( .A1(n6019), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5933) );
  INV_X1 U7500 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7235) );
  OR2_X1 U7501 ( .A1(n6109), .A2(n7235), .ZN(n5932) );
  OAI21_X1 U7502 ( .B1(n5925), .B2(P2_REG3_REG_5__SCAN_IN), .A(
        P2_REG3_REG_6__SCAN_IN), .ZN(n5928) );
  INV_X1 U7503 ( .A(n5925), .ZN(n5927) );
  NOR2_X1 U7504 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_REG3_REG_5__SCAN_IN), 
        .ZN(n5926) );
  NAND2_X1 U7505 ( .A1(n5927), .A2(n5926), .ZN(n5942) );
  AND2_X1 U7506 ( .A1(n5928), .A2(n5942), .ZN(n7291) );
  OR2_X1 U7507 ( .A1(n5914), .A2(n7291), .ZN(n5931) );
  INV_X1 U7508 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5929) );
  OR2_X1 U7509 ( .A1(n7003), .A2(n5929), .ZN(n5930) );
  NOR2_X1 U7510 ( .A1(n5934), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5937) );
  NOR2_X1 U7511 ( .A1(n5937), .A2(n6059), .ZN(n5935) );
  INV_X1 U7512 ( .A(n5936), .ZN(n5938) );
  NAND2_X1 U7513 ( .A1(n5938), .A2(n5962), .ZN(n8420) );
  INV_X1 U7514 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5939) );
  OR2_X1 U7515 ( .A1(n8320), .A2(n5939), .ZN(n5941) );
  OR2_X1 U7516 ( .A1(n8321), .A2(n6464), .ZN(n5940) );
  OAI211_X1 U7517 ( .C1(n6281), .C2(n8420), .A(n5941), .B(n5940), .ZN(n7157)
         );
  NAND2_X1 U7518 ( .A1(n7436), .A2(n7157), .ZN(n8216) );
  INV_X1 U7519 ( .A(n7436), .ZN(n8407) );
  INV_X1 U7520 ( .A(n7157), .ZN(n9934) );
  NAND2_X1 U7521 ( .A1(n8407), .A2(n9934), .ZN(n8214) );
  NAND2_X1 U7522 ( .A1(n6019), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5948) );
  OR2_X1 U7523 ( .A1(n6109), .A2(n9979), .ZN(n5947) );
  NAND2_X1 U7524 ( .A1(n5942), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5943) );
  AND2_X1 U7525 ( .A1(n5956), .A2(n5943), .ZN(n7431) );
  OR2_X1 U7526 ( .A1(n5914), .A2(n7431), .ZN(n5946) );
  INV_X1 U7527 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5944) );
  OR2_X1 U7528 ( .A1(n7003), .A2(n5944), .ZN(n5945) );
  NAND2_X1 U7529 ( .A1(n5962), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5950) );
  INV_X1 U7530 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5949) );
  XNOR2_X1 U7531 ( .A(n5950), .B(n5949), .ZN(n8454) );
  OR2_X1 U7532 ( .A1(n8320), .A2(n4701), .ZN(n5951) );
  INV_X1 U7533 ( .A(n6406), .ZN(n9939) );
  NAND2_X1 U7534 ( .A1(n8406), .A2(n9939), .ZN(n8219) );
  AND2_X1 U7535 ( .A1(n8214), .A2(n8219), .ZN(n5952) );
  INV_X1 U7536 ( .A(n8219), .ZN(n5953) );
  NAND2_X1 U7537 ( .A1(n7318), .A2(n6406), .ZN(n8226) );
  INV_X1 U7538 ( .A(n8352), .ZN(n8217) );
  OR2_X1 U7539 ( .A1(n5953), .A2(n8217), .ZN(n7408) );
  NAND2_X1 U7540 ( .A1(n6019), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5961) );
  INV_X1 U7541 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n5954) );
  OR2_X1 U7542 ( .A1(n6109), .A2(n5954), .ZN(n5960) );
  INV_X1 U7543 ( .A(n5956), .ZN(n5955) );
  NAND2_X1 U7544 ( .A1(n5955), .A2(n10095), .ZN(n5971) );
  NAND2_X1 U7545 ( .A1(n5956), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5957) );
  AND2_X1 U7546 ( .A1(n5971), .A2(n5957), .ZN(n7411) );
  OR2_X1 U7547 ( .A1(n5914), .A2(n7411), .ZN(n5959) );
  INV_X1 U7548 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8435) );
  OR2_X1 U7549 ( .A1(n7003), .A2(n8435), .ZN(n5958) );
  NAND2_X1 U7550 ( .A1(n5966), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5963) );
  XNOR2_X1 U7551 ( .A(n5963), .B(P2_IR_REG_8__SCAN_IN), .ZN(n8489) );
  AOI22_X1 U7552 ( .A1(n6097), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6422), .B2(
        n8489), .ZN(n5965) );
  NAND2_X1 U7553 ( .A1(n6469), .A2(n8316), .ZN(n5964) );
  NAND2_X1 U7554 ( .A1(n5965), .A2(n5964), .ZN(n7323) );
  NAND2_X1 U7555 ( .A1(n7435), .A2(n7323), .ZN(n8227) );
  AND2_X1 U7556 ( .A1(n7408), .A2(n8227), .ZN(n7392) );
  NAND2_X1 U7557 ( .A1(n6485), .A2(n8316), .ZN(n5969) );
  OAI21_X1 U7558 ( .B1(n5966), .B2(P2_IR_REG_8__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5967) );
  XNOR2_X1 U7559 ( .A(n5967), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9718) );
  AOI22_X1 U7560 ( .A1(n6097), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6422), .B2(
        n9718), .ZN(n5968) );
  NAND2_X1 U7561 ( .A1(n6019), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5977) );
  INV_X1 U7562 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n5970) );
  OR2_X1 U7563 ( .A1(n6109), .A2(n5970), .ZN(n5976) );
  NAND2_X1 U7564 ( .A1(n5971), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n5972) );
  AND2_X1 U7565 ( .A1(n5984), .A2(n5972), .ZN(n7403) );
  OR2_X1 U7566 ( .A1(n5914), .A2(n7403), .ZN(n5975) );
  INV_X1 U7567 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n5973) );
  OR2_X1 U7568 ( .A1(n7003), .A2(n5973), .ZN(n5974) );
  NAND4_X1 U7569 ( .A1(n5977), .A2(n5976), .A3(n5975), .A4(n5974), .ZN(n8404)
         );
  NAND2_X1 U7570 ( .A1(n9950), .A2(n8404), .ZN(n8221) );
  INV_X1 U7571 ( .A(n8404), .ZN(n7509) );
  INV_X1 U7572 ( .A(n9950), .ZN(n7405) );
  NAND2_X1 U7573 ( .A1(n7509), .A2(n7405), .ZN(n8228) );
  NAND2_X1 U7574 ( .A1(n8221), .A2(n8228), .ZN(n8351) );
  INV_X1 U7575 ( .A(n8351), .ZN(n5991) );
  AND2_X1 U7576 ( .A1(n7392), .A2(n5991), .ZN(n7389) );
  NAND2_X1 U7577 ( .A1(n6503), .A2(n8316), .ZN(n5982) );
  NOR2_X1 U7578 ( .A1(n5978), .A2(n6059), .ZN(n5979) );
  MUX2_X1 U7579 ( .A(n6059), .B(n5979), .S(P2_IR_REG_10__SCAN_IN), .Z(n5980)
         );
  OR2_X1 U7580 ( .A1(n5980), .A2(n5992), .ZN(n8481) );
  INV_X1 U7581 ( .A(n8481), .ZN(n9734) );
  AOI22_X1 U7582 ( .A1(n6097), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6422), .B2(
        n9734), .ZN(n5981) );
  NAND2_X1 U7583 ( .A1(n5982), .A2(n5981), .ZN(n7927) );
  NAND2_X1 U7584 ( .A1(n6019), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5989) );
  INV_X1 U7585 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8452) );
  OR2_X1 U7586 ( .A1(n6109), .A2(n8452), .ZN(n5988) );
  NAND2_X1 U7587 ( .A1(n5984), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n5985) );
  AND2_X1 U7588 ( .A1(n5999), .A2(n5985), .ZN(n8040) );
  OR2_X1 U7589 ( .A1(n5914), .A2(n8040), .ZN(n5987) );
  INV_X1 U7590 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8437) );
  OR2_X1 U7591 ( .A1(n7003), .A2(n8437), .ZN(n5986) );
  NAND4_X1 U7592 ( .A1(n5989), .A2(n5988), .A3(n5987), .A4(n5986), .ZN(n8403)
         );
  NAND2_X1 U7593 ( .A1(n7927), .A2(n8059), .ZN(n8238) );
  AND2_X1 U7594 ( .A1(n7389), .A2(n8238), .ZN(n5990) );
  NAND2_X1 U7595 ( .A1(n7409), .A2(n5990), .ZN(n7419) );
  INV_X1 U7596 ( .A(n7323), .ZN(n9944) );
  NAND2_X1 U7597 ( .A1(n8405), .A2(n9944), .ZN(n8220) );
  INV_X1 U7598 ( .A(n8220), .ZN(n7393) );
  NAND2_X1 U7599 ( .A1(n5991), .A2(n7393), .ZN(n7390) );
  NAND2_X1 U7600 ( .A1(n6530), .A2(n8316), .ZN(n5997) );
  NOR2_X1 U7601 ( .A1(n5992), .A2(n6059), .ZN(n5993) );
  MUX2_X1 U7602 ( .A(n6059), .B(n5993), .S(P2_IR_REG_11__SCAN_IN), .Z(n5995)
         );
  OR2_X1 U7603 ( .A1(n5995), .A2(n4613), .ZN(n8479) );
  AOI22_X1 U7604 ( .A1(n6097), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6422), .B2(
        n9752), .ZN(n5996) );
  NAND2_X1 U7605 ( .A1(n5997), .A2(n5996), .ZN(n9966) );
  NAND2_X1 U7606 ( .A1(n6019), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6004) );
  INV_X1 U7607 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n5998) );
  OR2_X1 U7608 ( .A1(n6109), .A2(n5998), .ZN(n6003) );
  NAND2_X1 U7609 ( .A1(n5999), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6000) );
  AND2_X1 U7610 ( .A1(n6010), .A2(n6000), .ZN(n8139) );
  OR2_X1 U7611 ( .A1(n5914), .A2(n8139), .ZN(n6002) );
  INV_X1 U7612 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7423) );
  OR2_X1 U7613 ( .A1(n7003), .A2(n7423), .ZN(n6001) );
  NAND4_X1 U7614 ( .A1(n6004), .A2(n6003), .A3(n6002), .A4(n6001), .ZN(n8402)
         );
  OR2_X1 U7615 ( .A1(n9966), .A2(n8063), .ZN(n8240) );
  NAND2_X1 U7616 ( .A1(n9966), .A2(n8063), .ZN(n8239) );
  AND2_X1 U7617 ( .A1(n7418), .A2(n8356), .ZN(n6005) );
  NAND2_X1 U7618 ( .A1(n7419), .A2(n6005), .ZN(n6006) );
  NAND2_X1 U7619 ( .A1(n6534), .A2(n8316), .ZN(n6009) );
  NAND2_X1 U7620 ( .A1(n6016), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6007) );
  XNOR2_X1 U7621 ( .A(n6007), .B(P2_IR_REG_12__SCAN_IN), .ZN(n9768) );
  AOI22_X1 U7622 ( .A1(n6097), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6422), .B2(
        n9768), .ZN(n6008) );
  NAND2_X1 U7623 ( .A1(n6009), .A2(n6008), .ZN(n8068) );
  NAND2_X1 U7624 ( .A1(n6999), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n6015) );
  INV_X1 U7625 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8440) );
  OR2_X1 U7626 ( .A1(n7003), .A2(n8440), .ZN(n6014) );
  NAND2_X1 U7627 ( .A1(n6010), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6011) );
  AND2_X1 U7628 ( .A1(n6022), .A2(n6011), .ZN(n8066) );
  OR2_X1 U7629 ( .A1(n5914), .A2(n8066), .ZN(n6013) );
  INV_X1 U7630 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n7482) );
  OR2_X1 U7631 ( .A1(n5878), .A2(n7482), .ZN(n6012) );
  OR2_X1 U7632 ( .A1(n8068), .A2(n8117), .ZN(n8245) );
  NAND2_X1 U7633 ( .A1(n8068), .A2(n8117), .ZN(n8246) );
  INV_X1 U7634 ( .A(n8355), .ZN(n7486) );
  NAND2_X1 U7635 ( .A1(n6621), .A2(n8316), .ZN(n6018) );
  OR2_X1 U7636 ( .A1(n6016), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U7637 ( .A1(n6058), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6029) );
  XNOR2_X1 U7638 ( .A(n6029), .B(P2_IR_REG_13__SCAN_IN), .ZN(n9787) );
  AOI22_X1 U7639 ( .A1(n6097), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6422), .B2(
        n9787), .ZN(n6017) );
  NAND2_X1 U7640 ( .A1(n6018), .A2(n6017), .ZN(n8249) );
  NAND2_X1 U7641 ( .A1(n6019), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6027) );
  INV_X1 U7642 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n7541) );
  OR2_X1 U7643 ( .A1(n6109), .A2(n7541), .ZN(n6026) );
  INV_X1 U7644 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U7645 ( .A1(n6022), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6023) );
  AND2_X1 U7646 ( .A1(n6036), .A2(n6023), .ZN(n8115) );
  OR2_X1 U7647 ( .A1(n5914), .A2(n8115), .ZN(n6025) );
  INV_X1 U7648 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8444) );
  OR2_X1 U7649 ( .A1(n7003), .A2(n8444), .ZN(n6024) );
  NAND4_X1 U7650 ( .A1(n6027), .A2(n6026), .A3(n6025), .A4(n6024), .ZN(n8704)
         );
  INV_X1 U7651 ( .A(n8704), .ZN(n8024) );
  NAND2_X1 U7652 ( .A1(n8249), .A2(n8024), .ZN(n6028) );
  NAND2_X1 U7653 ( .A1(n6644), .A2(n8316), .ZN(n6034) );
  NAND2_X1 U7654 ( .A1(n6029), .A2(n6055), .ZN(n6030) );
  NAND2_X1 U7655 ( .A1(n6030), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7656 ( .A1(n6031), .A2(n6056), .ZN(n6044) );
  OR2_X1 U7657 ( .A1(n6031), .A2(n6056), .ZN(n6032) );
  AOI22_X1 U7658 ( .A1(n6097), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6422), .B2(
        n9805), .ZN(n6033) );
  NAND2_X1 U7659 ( .A1(n6034), .A2(n6033), .ZN(n8849) );
  NAND2_X1 U7660 ( .A1(n6019), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6042) );
  INV_X1 U7661 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n8760) );
  OR2_X1 U7662 ( .A1(n6109), .A2(n8760), .ZN(n6041) );
  INV_X1 U7663 ( .A(n6036), .ZN(n6035) );
  NAND2_X1 U7664 ( .A1(n6036), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6037) );
  AND2_X1 U7665 ( .A1(n6048), .A2(n6037), .ZN(n8707) );
  OR2_X1 U7666 ( .A1(n5914), .A2(n8707), .ZN(n6040) );
  INV_X1 U7667 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n6038) );
  OR2_X1 U7668 ( .A1(n7003), .A2(n6038), .ZN(n6039) );
  NAND4_X1 U7669 ( .A1(n6042), .A2(n6041), .A3(n6040), .A4(n6039), .ZN(n8692)
         );
  OR2_X1 U7670 ( .A1(n8849), .A2(n8173), .ZN(n8260) );
  NAND2_X1 U7671 ( .A1(n8714), .A2(n8260), .ZN(n6043) );
  NAND2_X1 U7672 ( .A1(n8849), .A2(n8173), .ZN(n8261) );
  NAND2_X1 U7673 ( .A1(n6043), .A2(n8261), .ZN(n8688) );
  NAND2_X1 U7674 ( .A1(n6683), .A2(n8316), .ZN(n6047) );
  NAND2_X1 U7675 ( .A1(n6044), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6045) );
  XNOR2_X1 U7676 ( .A(n6045), .B(P2_IR_REG_15__SCAN_IN), .ZN(n9823) );
  AOI22_X1 U7677 ( .A1(n6097), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6422), .B2(
        n9823), .ZN(n6046) );
  NAND2_X1 U7678 ( .A1(n6019), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6053) );
  INV_X1 U7679 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8757) );
  OR2_X1 U7680 ( .A1(n6109), .A2(n8757), .ZN(n6052) );
  NAND2_X1 U7681 ( .A1(n6048), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6049) );
  AND2_X1 U7682 ( .A1(n6066), .A2(n6049), .ZN(n8169) );
  OR2_X1 U7683 ( .A1(n5914), .A2(n8169), .ZN(n6051) );
  INV_X1 U7684 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8694) );
  OR2_X1 U7685 ( .A1(n7003), .A2(n8694), .ZN(n6050) );
  OR2_X1 U7686 ( .A1(n8843), .A2(n8258), .ZN(n8675) );
  NAND3_X1 U7687 ( .A1(n6056), .A2(n6055), .A3(n6054), .ZN(n6057) );
  OR2_X1 U7688 ( .A1(n6062), .A2(n6059), .ZN(n6060) );
  MUX2_X1 U7689 ( .A(n6060), .B(P2_IR_REG_31__SCAN_IN), .S(n6061), .Z(n6063)
         );
  NAND2_X1 U7690 ( .A1(n6062), .A2(n6061), .ZN(n6082) );
  NAND2_X1 U7691 ( .A1(n6063), .A2(n6082), .ZN(n8469) );
  INV_X1 U7692 ( .A(n8469), .ZN(n9839) );
  AOI22_X1 U7693 ( .A1(n6097), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6422), .B2(
        n9839), .ZN(n6064) );
  NAND2_X1 U7694 ( .A1(n6019), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6071) );
  INV_X1 U7695 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8754) );
  OR2_X1 U7696 ( .A1(n6109), .A2(n8754), .ZN(n6070) );
  NAND2_X1 U7697 ( .A1(n6066), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6067) );
  AND2_X1 U7698 ( .A1(n6076), .A2(n6067), .ZN(n8683) );
  OR2_X1 U7699 ( .A1(n5914), .A2(n8683), .ZN(n6069) );
  INV_X1 U7700 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8682) );
  OR2_X1 U7701 ( .A1(n7003), .A2(n8682), .ZN(n6068) );
  AND2_X1 U7702 ( .A1(n8675), .A2(n8271), .ZN(n6072) );
  NAND2_X1 U7703 ( .A1(n8837), .A2(n8090), .ZN(n8266) );
  NAND2_X1 U7704 ( .A1(n6846), .A2(n8316), .ZN(n6075) );
  NAND2_X1 U7705 ( .A1(n6082), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6073) );
  XNOR2_X1 U7706 ( .A(n6073), .B(P2_IR_REG_17__SCAN_IN), .ZN(n9859) );
  AOI22_X1 U7707 ( .A1(n6097), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6422), .B2(
        n9859), .ZN(n6074) );
  NAND2_X1 U7708 ( .A1(n6019), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6081) );
  INV_X1 U7709 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8751) );
  OR2_X1 U7710 ( .A1(n6109), .A2(n8751), .ZN(n6080) );
  NAND2_X1 U7711 ( .A1(n6076), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6077) );
  AND2_X1 U7712 ( .A1(n6088), .A2(n6077), .ZN(n8670) );
  OR2_X1 U7713 ( .A1(n5914), .A2(n8670), .ZN(n6079) );
  INV_X1 U7714 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8669) );
  OR2_X1 U7715 ( .A1(n7003), .A2(n8669), .ZN(n6078) );
  NAND2_X1 U7716 ( .A1(n8831), .A2(n8146), .ZN(n8272) );
  NAND2_X1 U7717 ( .A1(n8664), .A2(n8272), .ZN(n8650) );
  NAND2_X1 U7718 ( .A1(n6952), .A2(n8316), .ZN(n6085) );
  NAND2_X1 U7719 ( .A1(n6095), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6083) );
  XNOR2_X1 U7720 ( .A(n6083), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8521) );
  AOI22_X1 U7721 ( .A1(n6097), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6422), .B2(
        n8521), .ZN(n6084) );
  NAND2_X1 U7722 ( .A1(n6019), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n6093) );
  INV_X1 U7723 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8748) );
  OR2_X1 U7724 ( .A1(n6109), .A2(n8748), .ZN(n6092) );
  INV_X1 U7725 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6086) );
  NAND2_X1 U7726 ( .A1(n6088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6089) );
  AND2_X1 U7727 ( .A1(n6100), .A2(n6089), .ZN(n8659) );
  OR2_X1 U7728 ( .A1(n5914), .A2(n8659), .ZN(n6091) );
  INV_X1 U7729 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8658) );
  OR2_X1 U7730 ( .A1(n7003), .A2(n8658), .ZN(n6090) );
  NAND4_X1 U7731 ( .A1(n6093), .A2(n6092), .A3(n6091), .A4(n6090), .ZN(n8667)
         );
  OR2_X1 U7732 ( .A1(n8825), .A2(n8643), .ZN(n8652) );
  OR2_X1 U7733 ( .A1(n8831), .A2(n8146), .ZN(n8649) );
  AND2_X1 U7734 ( .A1(n8652), .A2(n8649), .ZN(n8362) );
  NAND2_X1 U7735 ( .A1(n8650), .A2(n8362), .ZN(n6094) );
  NAND2_X1 U7736 ( .A1(n8825), .A2(n8643), .ZN(n8651) );
  NAND2_X1 U7737 ( .A1(n6094), .A2(n8651), .ZN(n8638) );
  NAND2_X1 U7738 ( .A1(n7070), .A2(n8316), .ZN(n6099) );
  AOI22_X1 U7739 ( .A1(n6097), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8516), .B2(
        n6422), .ZN(n6098) );
  NAND2_X1 U7740 ( .A1(n6019), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6105) );
  INV_X1 U7741 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8745) );
  OR2_X1 U7742 ( .A1(n6109), .A2(n8745), .ZN(n6104) );
  INV_X1 U7743 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8645) );
  OR2_X1 U7744 ( .A1(n7003), .A2(n8645), .ZN(n6103) );
  NAND2_X1 U7745 ( .A1(n6100), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6101) );
  AND2_X1 U7746 ( .A1(n6111), .A2(n6101), .ZN(n8644) );
  OR2_X1 U7747 ( .A1(n5914), .A2(n8644), .ZN(n6102) );
  NAND4_X1 U7748 ( .A1(n6105), .A2(n6104), .A3(n6103), .A4(n6102), .ZN(n8656)
         );
  OR2_X1 U7749 ( .A1(n8744), .A2(n7943), .ZN(n8281) );
  NAND2_X1 U7750 ( .A1(n8744), .A2(n7943), .ZN(n8280) );
  NAND2_X1 U7751 ( .A1(n8638), .A2(n8341), .ZN(n6106) );
  NAND2_X1 U7752 ( .A1(n6106), .A2(n8280), .ZN(n8625) );
  NAND2_X1 U7753 ( .A1(n7143), .A2(n8316), .ZN(n6108) );
  INV_X1 U7754 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7144) );
  OR2_X1 U7755 ( .A1(n8320), .A2(n7144), .ZN(n6107) );
  NAND2_X1 U7756 ( .A1(n6019), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6116) );
  INV_X1 U7757 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8740) );
  OR2_X1 U7758 ( .A1(n6109), .A2(n8740), .ZN(n6115) );
  NAND2_X1 U7759 ( .A1(n6111), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6112) );
  AND2_X1 U7760 ( .A1(n6120), .A2(n6112), .ZN(n8634) );
  OR2_X1 U7761 ( .A1(n5914), .A2(n8634), .ZN(n6114) );
  INV_X1 U7762 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8633) );
  OR2_X1 U7763 ( .A1(n7003), .A2(n8633), .ZN(n6113) );
  OR2_X1 U7764 ( .A1(n8814), .A2(n8642), .ZN(n8282) );
  NAND2_X1 U7765 ( .A1(n8814), .A2(n8642), .ZN(n8285) );
  NAND2_X1 U7766 ( .A1(n8625), .A2(n8627), .ZN(n6117) );
  NAND2_X1 U7767 ( .A1(n7178), .A2(n8316), .ZN(n6119) );
  INV_X1 U7768 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7182) );
  OR2_X1 U7769 ( .A1(n8320), .A2(n7182), .ZN(n6118) );
  NAND2_X1 U7770 ( .A1(n6120), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7771 ( .A1(n6130), .A2(n6121), .ZN(n8622) );
  NAND2_X1 U7772 ( .A1(n6202), .A2(n8622), .ZN(n6125) );
  INV_X1 U7773 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n8807) );
  OR2_X1 U7774 ( .A1(n5878), .A2(n8807), .ZN(n6124) );
  INV_X1 U7775 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8737) );
  OR2_X1 U7776 ( .A1(n6109), .A2(n8737), .ZN(n6123) );
  INV_X1 U7777 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n8621) );
  OR2_X1 U7778 ( .A1(n7003), .A2(n8621), .ZN(n6122) );
  NAND2_X1 U7779 ( .A1(n8808), .A2(n8125), .ZN(n8286) );
  INV_X1 U7780 ( .A(n8286), .ZN(n6126) );
  NAND2_X1 U7781 ( .A1(n7312), .A2(n8316), .ZN(n6128) );
  OR2_X1 U7782 ( .A1(n8320), .A2(n7315), .ZN(n6127) );
  NAND2_X1 U7783 ( .A1(n6130), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7784 ( .A1(n6137), .A2(n6131), .ZN(n8128) );
  AOI22_X1 U7785 ( .A1(n8128), .A2(n6202), .B1(n6139), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n6133) );
  AOI22_X1 U7786 ( .A1(n6019), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n6999), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n6132) );
  INV_X1 U7787 ( .A(n8291), .ZN(n6134) );
  NAND2_X1 U7788 ( .A1(n8129), .A2(n8604), .ZN(n8290) );
  NAND2_X1 U7789 ( .A1(n7368), .A2(n8316), .ZN(n6136) );
  OR2_X1 U7790 ( .A1(n8320), .A2(n7366), .ZN(n6135) );
  NAND2_X1 U7791 ( .A1(n6137), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6138) );
  NAND2_X1 U7792 ( .A1(n6145), .A2(n6138), .ZN(n8608) );
  NAND2_X1 U7793 ( .A1(n8608), .A2(n6202), .ZN(n6142) );
  AOI22_X1 U7794 ( .A1(n6019), .A2(P2_REG0_REG_23__SCAN_IN), .B1(n6999), .B2(
        P2_REG1_REG_23__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7795 ( .A1(n6139), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6140) );
  NAND2_X1 U7796 ( .A1(n8802), .A2(n8400), .ZN(n8340) );
  NAND2_X1 U7797 ( .A1(n8600), .A2(n8340), .ZN(n8594) );
  NAND2_X1 U7798 ( .A1(n7474), .A2(n8316), .ZN(n6144) );
  OR2_X1 U7799 ( .A1(n8320), .A2(n7475), .ZN(n6143) );
  INV_X1 U7800 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6149) );
  NAND2_X1 U7801 ( .A1(n6145), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6146) );
  NAND2_X1 U7802 ( .A1(n6155), .A2(n6146), .ZN(n8592) );
  NAND2_X1 U7803 ( .A1(n8592), .A2(n6202), .ZN(n6148) );
  AOI22_X1 U7804 ( .A1(n6019), .A2(P2_REG0_REG_24__SCAN_IN), .B1(n6999), .B2(
        P2_REG1_REG_24__SCAN_IN), .ZN(n6147) );
  OAI211_X1 U7805 ( .C1(n7003), .C2(n6149), .A(n6148), .B(n6147), .ZN(n8399)
         );
  NAND2_X1 U7806 ( .A1(n8101), .A2(n8605), .ZN(n8338) );
  NAND2_X1 U7807 ( .A1(n8609), .A2(n8590), .ZN(n8593) );
  NAND2_X1 U7808 ( .A1(n8594), .A2(n8295), .ZN(n6150) );
  NAND2_X1 U7809 ( .A1(n6150), .A2(n8339), .ZN(n8583) );
  NAND2_X1 U7810 ( .A1(n7516), .A2(n8316), .ZN(n6152) );
  OR2_X1 U7811 ( .A1(n8320), .A2(n7517), .ZN(n6151) );
  INV_X1 U7812 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6153) );
  NAND2_X1 U7813 ( .A1(n6155), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6156) );
  NAND2_X1 U7814 ( .A1(n6168), .A2(n6156), .ZN(n8581) );
  NAND2_X1 U7815 ( .A1(n8581), .A2(n6202), .ZN(n6162) );
  INV_X1 U7816 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n6159) );
  NAND2_X1 U7817 ( .A1(n6999), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U7818 ( .A1(n6019), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6157) );
  OAI211_X1 U7819 ( .C1(n6159), .C2(n7003), .A(n6158), .B(n6157), .ZN(n6160)
         );
  INV_X1 U7820 ( .A(n6160), .ZN(n6161) );
  NAND2_X1 U7821 ( .A1(n8076), .A2(n8589), .ZN(n8299) );
  NAND2_X1 U7822 ( .A1(n8583), .A2(n8299), .ZN(n6163) );
  NAND2_X1 U7823 ( .A1(n7522), .A2(n8316), .ZN(n6165) );
  OR2_X1 U7824 ( .A1(n8320), .A2(n7523), .ZN(n6164) );
  INV_X1 U7825 ( .A(n6168), .ZN(n6167) );
  INV_X1 U7826 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n6166) );
  NAND2_X1 U7827 ( .A1(n6168), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7828 ( .A1(n6178), .A2(n6169), .ZN(n8572) );
  NAND2_X1 U7829 ( .A1(n8572), .A2(n6202), .ZN(n6174) );
  INV_X1 U7830 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8571) );
  NAND2_X1 U7831 ( .A1(n6019), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6171) );
  NAND2_X1 U7832 ( .A1(n6999), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6170) );
  OAI211_X1 U7833 ( .C1(n8571), .C2(n7003), .A(n6171), .B(n6170), .ZN(n6172)
         );
  INV_X1 U7834 ( .A(n6172), .ZN(n6173) );
  NOR2_X1 U7835 ( .A1(n8786), .A2(n8579), .ZN(n8303) );
  NAND2_X1 U7836 ( .A1(n8786), .A2(n8579), .ZN(n8297) );
  NAND2_X1 U7837 ( .A1(n7528), .A2(n8316), .ZN(n6177) );
  OR2_X1 U7838 ( .A1(n8320), .A2(n8859), .ZN(n6176) );
  NAND2_X1 U7839 ( .A1(n6178), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6179) );
  NAND2_X1 U7840 ( .A1(n6197), .A2(n6179), .ZN(n8560) );
  NAND2_X1 U7841 ( .A1(n8560), .A2(n6202), .ZN(n6185) );
  INV_X1 U7842 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n6182) );
  NAND2_X1 U7843 ( .A1(n6019), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7844 ( .A1(n6999), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6180) );
  OAI211_X1 U7845 ( .C1(n6182), .C2(n7003), .A(n6181), .B(n6180), .ZN(n6183)
         );
  INV_X1 U7846 ( .A(n6183), .ZN(n6184) );
  OR2_X1 U7847 ( .A1(n8561), .A2(n8305), .ZN(n6186) );
  INV_X1 U7848 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7823) );
  MUX2_X1 U7849 ( .A(n7823), .B(n7902), .S(n7550), .Z(n6191) );
  INV_X1 U7850 ( .A(SI_28_), .ZN(n6190) );
  NAND2_X1 U7851 ( .A1(n6191), .A2(n6190), .ZN(n6205) );
  INV_X1 U7852 ( .A(n6191), .ZN(n6192) );
  NAND2_X1 U7853 ( .A1(n6192), .A2(SI_28_), .ZN(n6193) );
  NAND2_X1 U7854 ( .A1(n7901), .A2(n8316), .ZN(n6195) );
  OR2_X1 U7855 ( .A1(n8320), .A2(n7823), .ZN(n6194) );
  INV_X1 U7856 ( .A(n6197), .ZN(n6196) );
  INV_X1 U7857 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n7968) );
  NAND2_X1 U7858 ( .A1(n6196), .A2(n7968), .ZN(n8002) );
  NAND2_X1 U7859 ( .A1(n6197), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6198) );
  NAND2_X1 U7860 ( .A1(n8002), .A2(n6198), .ZN(n8547) );
  INV_X1 U7861 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n8546) );
  NAND2_X1 U7862 ( .A1(n6019), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6200) );
  NAND2_X1 U7863 ( .A1(n6999), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6199) );
  OAI211_X1 U7864 ( .C1(n8546), .C2(n5903), .A(n6200), .B(n6199), .ZN(n6201)
         );
  AOI21_X1 U7865 ( .B1(n8547), .B2(n6202), .A(n6201), .ZN(n8558) );
  MUX2_X1 U7866 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n7550), .Z(n7545) );
  INV_X1 U7867 ( .A(SI_29_), .ZN(n6207) );
  NAND2_X1 U7868 ( .A1(n7584), .A2(n7583), .ZN(n9524) );
  OR2_X1 U7869 ( .A1(n9524), .A2(n8321), .ZN(n6209) );
  INV_X1 U7870 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7825) );
  OR2_X1 U7871 ( .A1(n8320), .A2(n7825), .ZN(n6208) );
  OR2_X1 U7872 ( .A1(n8002), .A2(n5914), .ZN(n7007) );
  INV_X1 U7873 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8004) );
  NAND2_X1 U7874 ( .A1(n6019), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6211) );
  NAND2_X1 U7875 ( .A1(n6999), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6210) );
  OAI211_X1 U7876 ( .C1(n8004), .C2(n5903), .A(n6211), .B(n6210), .ZN(n6212)
         );
  INV_X1 U7877 ( .A(n6212), .ZN(n6213) );
  NAND2_X1 U7878 ( .A1(n8311), .A2(n8312), .ZN(n8332) );
  NAND2_X1 U7879 ( .A1(n8377), .A2(n8332), .ZN(n6267) );
  XNOR2_X1 U7880 ( .A(n8378), .B(n6267), .ZN(n8006) );
  INV_X1 U7881 ( .A(n6214), .ZN(n6215) );
  NAND2_X1 U7882 ( .A1(n6215), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6216) );
  MUX2_X1 U7883 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6216), .S(
        P2_IR_REG_20__SCAN_IN), .Z(n6218) );
  INV_X1 U7884 ( .A(n6217), .ZN(n6269) );
  NAND2_X1 U7885 ( .A1(n8516), .A2(n8324), .ZN(n9906) );
  NAND2_X1 U7886 ( .A1(n6219), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6220) );
  INV_X1 U7887 ( .A(n8068), .ZN(n6248) );
  NAND4_X1 U7888 ( .A1(n6224), .A2(n6223), .A3(n6222), .A4(n6221), .ZN(n6225)
         );
  NAND2_X1 U7889 ( .A1(n6225), .A2(n6832), .ZN(n7990) );
  NAND2_X1 U7890 ( .A1(n9892), .A2(n9912), .ZN(n9896) );
  NAND2_X1 U7891 ( .A1(n9898), .A2(n9896), .ZN(n6226) );
  NAND2_X1 U7892 ( .A1(n7991), .A2(n9904), .ZN(n6227) );
  NAND2_X1 U7893 ( .A1(n9881), .A2(n9920), .ZN(n6228) );
  INV_X1 U7894 ( .A(n9920), .ZN(n8191) );
  NAND2_X1 U7895 ( .A1(n9894), .A2(n8191), .ZN(n6229) );
  NOR2_X1 U7896 ( .A1(n8202), .A2(n9924), .ZN(n6231) );
  NAND2_X1 U7897 ( .A1(n8202), .A2(n9924), .ZN(n6230) );
  AND2_X1 U7898 ( .A1(n9879), .A2(n6378), .ZN(n6232) );
  INV_X1 U7899 ( .A(n8348), .ZN(n6233) );
  NAND2_X1 U7900 ( .A1(n7026), .A2(n9929), .ZN(n7292) );
  AND2_X1 U7901 ( .A1(n6233), .A2(n7292), .ZN(n6234) );
  NAND2_X1 U7902 ( .A1(n8407), .A2(n7157), .ZN(n6235) );
  NAND2_X1 U7903 ( .A1(n7318), .A2(n9939), .ZN(n6236) );
  NAND2_X1 U7904 ( .A1(n8227), .A2(n8220), .ZN(n8350) );
  NAND2_X1 U7905 ( .A1(n7927), .A2(n8403), .ZN(n6241) );
  INV_X1 U7906 ( .A(n6241), .ZN(n7503) );
  NOR2_X1 U7907 ( .A1(n7927), .A2(n8403), .ZN(n7504) );
  INV_X1 U7908 ( .A(n7504), .ZN(n6237) );
  NAND2_X1 U7909 ( .A1(n9950), .A2(n7509), .ZN(n7506) );
  AND2_X1 U7910 ( .A1(n6237), .A2(n7506), .ZN(n6238) );
  OR2_X1 U7911 ( .A1(n7503), .A2(n6238), .ZN(n6240) );
  AND2_X1 U7912 ( .A1(n8350), .A2(n6240), .ZN(n6239) );
  INV_X1 U7913 ( .A(n6240), .ZN(n6244) );
  AND2_X1 U7914 ( .A1(n8351), .A2(n6241), .ZN(n6242) );
  NAND2_X1 U7915 ( .A1(n8405), .A2(n7323), .ZN(n7398) );
  AND2_X1 U7916 ( .A1(n6242), .A2(n7398), .ZN(n6243) );
  OR2_X1 U7917 ( .A1(n6244), .A2(n6243), .ZN(n6245) );
  NAND2_X1 U7918 ( .A1(n6246), .A2(n6245), .ZN(n7421) );
  AND2_X1 U7919 ( .A1(n9966), .A2(n8402), .ZN(n6247) );
  OR2_X1 U7920 ( .A1(n8249), .A2(n8704), .ZN(n8252) );
  AND2_X1 U7921 ( .A1(n8249), .A2(n8704), .ZN(n8253) );
  NAND2_X1 U7922 ( .A1(n8849), .A2(n8692), .ZN(n6249) );
  INV_X1 U7923 ( .A(n8849), .ZN(n8709) );
  NAND2_X1 U7924 ( .A1(n8259), .A2(n8258), .ZN(n6250) );
  INV_X1 U7925 ( .A(n8837), .ZN(n6251) );
  NAND2_X1 U7926 ( .A1(n8649), .A2(n8272), .ZN(n8666) );
  NAND2_X1 U7927 ( .A1(n8825), .A2(n8667), .ZN(n6253) );
  INV_X1 U7928 ( .A(n8825), .ZN(n6252) );
  NAND2_X1 U7929 ( .A1(n8640), .A2(n6254), .ZN(n6256) );
  INV_X1 U7930 ( .A(n8744), .ZN(n6255) );
  NAND2_X1 U7931 ( .A1(n6256), .A2(n4393), .ZN(n8626) );
  INV_X1 U7932 ( .A(n6257), .ZN(n8628) );
  INV_X1 U7933 ( .A(n8814), .ZN(n6258) );
  NAND2_X1 U7934 ( .A1(n6258), .A2(n8642), .ZN(n8614) );
  NOR2_X1 U7935 ( .A1(n8808), .A2(n8631), .ZN(n7906) );
  NAND2_X1 U7936 ( .A1(n8291), .A2(n8290), .ZN(n7905) );
  OAI21_X1 U7937 ( .B1(n8619), .B2(n8129), .A(n7908), .ZN(n8601) );
  OAI21_X1 U7938 ( .B1(n8590), .B2(n8802), .A(n8601), .ZN(n6259) );
  NOR2_X1 U7939 ( .A1(n8101), .A2(n8399), .ZN(n6260) );
  NAND2_X1 U7940 ( .A1(n8791), .A2(n8589), .ZN(n6261) );
  NAND2_X1 U7941 ( .A1(n8786), .A2(n8398), .ZN(n6263) );
  NOR2_X1 U7942 ( .A1(n8786), .A2(n8398), .ZN(n6262) );
  NAND2_X1 U7943 ( .A1(n8561), .A2(n8568), .ZN(n6264) );
  NAND2_X1 U7944 ( .A1(n6265), .A2(n6264), .ZN(n8544) );
  NOR2_X1 U7945 ( .A1(n8778), .A2(n8558), .ZN(n6266) );
  XNOR2_X1 U7946 ( .A(n6268), .B(n6267), .ZN(n6284) );
  NAND2_X1 U7947 ( .A1(n8516), .A2(n8391), .ZN(n6324) );
  NAND2_X1 U7948 ( .A1(n6269), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U7949 ( .A1(n8180), .A2(n6323), .ZN(n8382) );
  INV_X1 U7950 ( .A(n8391), .ZN(n8182) );
  OAI21_X1 U7951 ( .B1(n8391), .B2(n8324), .A(n9955), .ZN(n6271) );
  NOR2_X1 U7952 ( .A1(n8516), .A2(n6271), .ZN(n6272) );
  INV_X1 U7953 ( .A(n8558), .ZN(n8397) );
  INV_X1 U7954 ( .A(n6273), .ZN(n6444) );
  NAND2_X1 U7955 ( .A1(n6444), .A2(n8389), .ZN(n6275) );
  NAND2_X1 U7956 ( .A1(n6281), .A2(n6275), .ZN(n6410) );
  INV_X1 U7957 ( .A(n6410), .ZN(n6409) );
  INV_X1 U7958 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6278) );
  NAND2_X1 U7959 ( .A1(n6019), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U7960 ( .A1(n6999), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n6276) );
  OAI211_X1 U7961 ( .C1(n6278), .C2(n5903), .A(n6277), .B(n6276), .ZN(n6279)
         );
  INV_X1 U7962 ( .A(n6279), .ZN(n6280) );
  NAND2_X1 U7963 ( .A1(n7007), .A2(n6280), .ZN(n8396) );
  AND2_X1 U7964 ( .A1(n6281), .A2(P2_B_REG_SCAN_IN), .ZN(n6282) );
  NOR2_X1 U7965 ( .A1(n9893), .A2(n6282), .ZN(n8535) );
  AOI22_X1 U7966 ( .A1(n8397), .A2(n9880), .B1(n8396), .B2(n8535), .ZN(n6283)
         );
  NAND2_X1 U7967 ( .A1(n6292), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6293) );
  MUX2_X1 U7968 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6293), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6295) );
  NAND2_X1 U7969 ( .A1(n7518), .A2(n7524), .ZN(n6542) );
  NAND2_X1 U7970 ( .A1(n7524), .A2(n7476), .ZN(n6540) );
  NOR2_X1 U7971 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6302) );
  NOR4_X1 U7972 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6301) );
  NOR4_X1 U7973 ( .A1(P2_D_REG_12__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6300) );
  NOR4_X1 U7974 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_26__SCAN_IN), .ZN(n6299) );
  NAND4_X1 U7975 ( .A1(n6302), .A2(n6301), .A3(n6300), .A4(n6299), .ZN(n6308)
         );
  NOR4_X1 U7976 ( .A1(P2_D_REG_14__SCAN_IN), .A2(P2_D_REG_13__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6306) );
  NOR4_X1 U7977 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_9__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_15__SCAN_IN), .ZN(n6305) );
  NOR4_X1 U7978 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6304) );
  NOR4_X1 U7979 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6303) );
  NAND4_X1 U7980 ( .A1(n6306), .A2(n6305), .A3(n6304), .A4(n6303), .ZN(n6307)
         );
  NOR2_X1 U7981 ( .A1(n6308), .A2(n6307), .ZN(n6309) );
  INV_X1 U7982 ( .A(n7518), .ZN(n6311) );
  NOR2_X1 U7983 ( .A1(n7524), .A2(n7476), .ZN(n6310) );
  NOR2_X1 U7984 ( .A1(n9957), .A2(n8180), .ZN(n6404) );
  INV_X1 U7985 ( .A(n8516), .ZN(n8526) );
  NAND3_X1 U7986 ( .A1(n8526), .A2(n8391), .A3(n6323), .ZN(n6314) );
  AND2_X1 U7987 ( .A1(n6314), .A2(n8315), .ZN(n6315) );
  OAI21_X1 U7988 ( .B1(n6825), .B2(n6404), .A(n6315), .ZN(n6317) );
  AOI21_X1 U7989 ( .B1(n8526), .B2(n8324), .A(n8315), .ZN(n6824) );
  AOI21_X1 U7990 ( .B1(n6389), .B2(n6828), .A(n6824), .ZN(n6316) );
  AND2_X1 U7991 ( .A1(n6317), .A2(n6316), .ZN(n6318) );
  INV_X1 U7992 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6319) );
  NAND2_X1 U7993 ( .A1(n9984), .A2(n6319), .ZN(n6320) );
  OAI21_X1 U7994 ( .B1(n6332), .B2(n9984), .A(n6320), .ZN(n6321) );
  INV_X1 U7995 ( .A(n8311), .ZN(n6333) );
  NAND2_X1 U7996 ( .A1(n6321), .A2(n4432), .ZN(P2_U3488) );
  INV_X1 U7997 ( .A(n6326), .ZN(n6322) );
  NAND2_X1 U7998 ( .A1(n7180), .A2(n6323), .ZN(n8374) );
  OR2_X1 U7999 ( .A1(n6324), .A2(n8374), .ZN(n6385) );
  NAND2_X1 U8000 ( .A1(n6385), .A2(n6821), .ZN(n6325) );
  NAND2_X1 U8001 ( .A1(n6403), .A2(n6325), .ZN(n6329) );
  AND2_X1 U8002 ( .A1(n8315), .A2(n9955), .ZN(n6327) );
  NAND2_X1 U8003 ( .A1(n6385), .A2(n6327), .ZN(n6383) );
  NAND2_X1 U8004 ( .A1(n9906), .A2(n9967), .ZN(n8708) );
  NAND2_X1 U8005 ( .A1(n6383), .A2(n8708), .ZN(n6392) );
  NAND2_X1 U8006 ( .A1(n6408), .A2(n6392), .ZN(n6328) );
  INV_X1 U8007 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6330) );
  NAND2_X1 U8008 ( .A1(n9970), .A2(n6330), .ZN(n6331) );
  NAND2_X1 U8009 ( .A1(n6334), .A2(n4433), .ZN(P2_U3456) );
  INV_X2 U8010 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NAND2_X1 U8011 ( .A1(n7901), .A2(n7590), .ZN(n6336) );
  OR2_X1 U8012 ( .A1(n7596), .A2(n7902), .ZN(n6335) );
  NAND2_X1 U8013 ( .A1(n9183), .A2(n5361), .ZN(n6339) );
  OR2_X1 U8014 ( .A1(n9381), .A2(n6337), .ZN(n6338) );
  NAND2_X1 U8015 ( .A1(n6339), .A2(n6338), .ZN(n6340) );
  XNOR2_X1 U8016 ( .A(n6340), .B(n5222), .ZN(n6345) );
  NAND2_X1 U8017 ( .A1(n9183), .A2(n6341), .ZN(n6342) );
  OAI21_X1 U8018 ( .B1(n9381), .B2(n6343), .A(n6342), .ZN(n6344) );
  XNOR2_X1 U8019 ( .A(n6345), .B(n6344), .ZN(n6352) );
  NAND3_X1 U8020 ( .A1(n6358), .A2(n6352), .A3(n9016), .ZN(n6361) );
  INV_X1 U8021 ( .A(n9026), .ZN(n8958) );
  INV_X1 U8022 ( .A(n7978), .ZN(n6349) );
  INV_X1 U8023 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n7897) );
  NAND2_X1 U8024 ( .A1(n5160), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6347) );
  NAND2_X1 U8025 ( .A1(n6493), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n6346) );
  OAI211_X1 U8026 ( .C1(n6494), .C2(n7897), .A(n6347), .B(n6346), .ZN(n6348)
         );
  AOI21_X1 U8027 ( .B1(n6349), .B2(n5442), .A(n6348), .ZN(n9372) );
  AOI22_X1 U8028 ( .A1(n4458), .A2(n9018), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n6351) );
  NAND2_X1 U8029 ( .A1(n9178), .A2(n9022), .ZN(n6350) );
  OAI211_X1 U8030 ( .C1(n9391), .C2(n8988), .A(n6351), .B(n6350), .ZN(n6354)
         );
  INV_X1 U8031 ( .A(n6352), .ZN(n6356) );
  INV_X1 U8032 ( .A(n9016), .ZN(n8960) );
  NOR3_X1 U8033 ( .A1(n6356), .A2(n6355), .A3(n8960), .ZN(n6353) );
  AOI211_X1 U8034 ( .C1(n9183), .C2(n8958), .A(n6354), .B(n6353), .ZN(n6360)
         );
  NAND3_X1 U8035 ( .A1(n6356), .A2(n9016), .A3(n6355), .ZN(n6357) );
  INV_X1 U8036 ( .A(n6721), .ZN(n6362) );
  INV_X2 U8037 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  INV_X1 U8038 ( .A(n6363), .ZN(n6364) );
  AND2_X2 U8039 ( .A1(n6364), .A2(n5169), .ZN(P1_U3973) );
  INV_X1 U8040 ( .A(n8374), .ZN(n6365) );
  NAND2_X1 U8041 ( .A1(n6366), .A2(n6365), .ZN(n6369) );
  NAND2_X1 U8042 ( .A1(n8516), .A2(n7180), .ZN(n6367) );
  NAND2_X1 U8043 ( .A1(n6367), .A2(n8324), .ZN(n6368) );
  NAND2_X2 U8044 ( .A1(n6369), .A2(n6368), .ZN(n6370) );
  XNOR2_X1 U8045 ( .A(n6370), .B(n6406), .ZN(n7317) );
  XNOR2_X1 U8046 ( .A(n7317), .B(n7318), .ZN(n6382) );
  XNOR2_X1 U8047 ( .A(n9934), .B(n6370), .ZN(n6380) );
  XNOR2_X1 U8048 ( .A(n6370), .B(n9924), .ZN(n6376) );
  INV_X1 U8049 ( .A(n6376), .ZN(n6377) );
  XNOR2_X1 U8050 ( .A(n8191), .B(n6370), .ZN(n6375) );
  XNOR2_X1 U8051 ( .A(n6371), .B(n9892), .ZN(n6719) );
  OAI21_X1 U8052 ( .B1(n6832), .B2(n6370), .A(n8187), .ZN(n6720) );
  INV_X1 U8053 ( .A(n6371), .ZN(n6372) );
  XNOR2_X1 U8054 ( .A(n6370), .B(n6373), .ZN(n6374) );
  XNOR2_X1 U8055 ( .A(n6375), .B(n9881), .ZN(n6946) );
  XNOR2_X1 U8056 ( .A(n6376), .B(n8202), .ZN(n7023) );
  OAI21_X1 U8057 ( .B1(n6377), .B2(n8202), .A(n7022), .ZN(n7146) );
  XNOR2_X1 U8058 ( .A(n6370), .B(n6378), .ZN(n6379) );
  XNOR2_X1 U8059 ( .A(n6379), .B(n9879), .ZN(n7145) );
  XNOR2_X1 U8060 ( .A(n6380), .B(n7436), .ZN(n7155) );
  AOI21_X1 U8061 ( .B1(n6382), .B2(n6381), .A(n7316), .ZN(n6388) );
  INV_X1 U8062 ( .A(n6383), .ZN(n6384) );
  NAND2_X1 U8063 ( .A1(n6403), .A2(n6384), .ZN(n6387) );
  INV_X1 U8064 ( .A(n6385), .ZN(n6390) );
  NAND2_X1 U8065 ( .A1(n6408), .A2(n6390), .ZN(n6386) );
  NOR2_X1 U8066 ( .A1(n6388), .A2(n8164), .ZN(n6417) );
  NAND3_X1 U8067 ( .A1(n6389), .A2(n6825), .A3(n6391), .ZN(n6400) );
  NAND2_X1 U8068 ( .A1(n6400), .A2(n6390), .ZN(n6397) );
  INV_X1 U8069 ( .A(n6824), .ZN(n6396) );
  INV_X1 U8070 ( .A(n6391), .ZN(n6393) );
  OAI21_X1 U8071 ( .B1(n6394), .B2(n6393), .A(n6392), .ZN(n6395) );
  NAND4_X1 U8072 ( .A1(n6397), .A2(n6419), .A3(n6396), .A4(n6395), .ZN(n6398)
         );
  NAND2_X1 U8073 ( .A1(n6398), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6402) );
  INV_X1 U8074 ( .A(n6821), .ZN(n6407) );
  NAND2_X1 U8075 ( .A1(n6505), .A2(n6407), .ZN(n8390) );
  INV_X1 U8076 ( .A(n8390), .ZN(n6399) );
  NAND2_X1 U8077 ( .A1(n6400), .A2(n6399), .ZN(n6401) );
  AND2_X1 U8078 ( .A1(n6402), .A2(n6401), .ZN(n6722) );
  OR2_X1 U8079 ( .A1(n6420), .A2(P2_U3151), .ZN(n8394) );
  NOR2_X1 U8080 ( .A1(n8149), .A2(n7431), .ZN(n6416) );
  NAND2_X1 U8081 ( .A1(n6403), .A2(n9967), .ZN(n6405) );
  AND2_X1 U8082 ( .A1(n8162), .A2(n6406), .ZN(n6415) );
  AND2_X1 U8083 ( .A1(n6408), .A2(n6407), .ZN(n6411) );
  NAND2_X1 U8084 ( .A1(n6411), .A2(n6409), .ZN(n8172) );
  NAND2_X1 U8085 ( .A1(n8170), .A2(n8405), .ZN(n6413) );
  INV_X1 U8086 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10127) );
  NOR2_X1 U8087 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10127), .ZN(n7229) );
  INV_X1 U8088 ( .A(n7229), .ZN(n6412) );
  OAI211_X1 U8089 ( .C1(n7436), .C2(n8172), .A(n6413), .B(n6412), .ZN(n6414)
         );
  OR4_X1 U8090 ( .A1(n6417), .A2(n6416), .A3(n6415), .A4(n6414), .ZN(P2_U3153)
         );
  INV_X1 U8091 ( .A(n6420), .ZN(n6418) );
  NAND2_X1 U8092 ( .A1(n8329), .A2(n6420), .ZN(n6421) );
  NAND2_X1 U8093 ( .A1(n6424), .A2(n6421), .ZN(n6432) );
  OR2_X1 U8094 ( .A1(n6432), .A2(n6422), .ZN(n6423) );
  NAND2_X1 U8095 ( .A1(n6423), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NOR2_X2 U8096 ( .A1(P2_U3150), .A2(n6428), .ZN(n9857) );
  INV_X1 U8097 ( .A(n9857), .ZN(n7067) );
  INV_X1 U8098 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n9990) );
  NOR2_X1 U8099 ( .A1(n7067), .A2(n9990), .ZN(n6449) );
  NOR2_X1 U8100 ( .A1(n6274), .A2(P2_U3151), .ZN(n6425) );
  NAND2_X1 U8101 ( .A1(n6425), .A2(n6273), .ZN(n6426) );
  OR2_X1 U8102 ( .A1(n6432), .A2(n6426), .ZN(n6430) );
  OR2_X1 U8103 ( .A1(n6273), .A2(P2_U3151), .ZN(n7821) );
  INV_X1 U8104 ( .A(n7821), .ZN(n6427) );
  NAND2_X1 U8105 ( .A1(n6428), .A2(n6427), .ZN(n6429) );
  INV_X1 U8106 ( .A(n9858), .ZN(n9708) );
  OAI22_X1 U8107 ( .A1(n9708), .A2(n6896), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6431), .ZN(n6448) );
  NOR2_X2 U8108 ( .A1(n6609), .A2(n8389), .ZN(n9867) );
  INV_X1 U8109 ( .A(n9867), .ZN(n9699) );
  NAND2_X1 U8110 ( .A1(n6437), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6904) );
  NAND2_X1 U8111 ( .A1(n6896), .A2(n6904), .ZN(n6435) );
  INV_X1 U8112 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6436) );
  NAND2_X1 U8113 ( .A1(n6436), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6433) );
  OR2_X1 U8114 ( .A1(n6433), .A2(n6437), .ZN(n6434) );
  NAND2_X1 U8115 ( .A1(n6435), .A2(n6434), .ZN(n6903) );
  XOR2_X1 U8116 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6903), .Z(n6443) );
  AND2_X1 U8117 ( .A1(n6436), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6438) );
  NAND2_X1 U8118 ( .A1(n6437), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6909) );
  OR2_X1 U8119 ( .A1(n6440), .A2(n7996), .ZN(n6910) );
  INV_X1 U8120 ( .A(n6910), .ZN(n6439) );
  AOI21_X1 U8121 ( .B1(n7996), .B2(n6440), .A(n6439), .ZN(n6442) );
  INV_X1 U8122 ( .A(n6609), .ZN(n6441) );
  OAI22_X1 U8123 ( .A1(n9699), .A2(n6443), .B1(n6442), .B2(n9872), .ZN(n6447)
         );
  MUX2_X1 U8124 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n6274), .Z(n6897) );
  XNOR2_X1 U8125 ( .A(n6897), .B(n6896), .ZN(n6445) );
  MUX2_X1 U8126 ( .A(n5870), .B(n5868), .S(n6274), .Z(n6608) );
  AND2_X1 U8127 ( .A1(n6608), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6606) );
  NOR2_X1 U8128 ( .A1(n6445), .A2(n6606), .ZN(n6895) );
  AOI211_X1 U8129 ( .C1(n6445), .C2(n6606), .A(n8529), .B(n6895), .ZN(n6446)
         );
  OR4_X1 U8130 ( .A1(n6449), .A2(n6448), .A3(n6447), .A4(n6446), .ZN(P2_U3183)
         );
  AND2_X1 U8131 ( .A1(n6452), .A2(P2_U3151), .ZN(n7820) );
  INV_X2 U8132 ( .A(n7820), .ZN(n8858) );
  OAI222_X1 U8133 ( .A1(n7561), .A2(n6451), .B1(n8858), .B2(n6453), .C1(
        P2_U3151), .C2(n7062), .ZN(P2_U3293) );
  OAI222_X1 U8134 ( .A1(n7561), .A2(n4466), .B1(n8858), .B2(n6455), .C1(
        P2_U3151), .C2(n6992), .ZN(P2_U3292) );
  INV_X2 U8135 ( .A(n7367), .ZN(n9525) );
  OAI222_X1 U8136 ( .A1(n9521), .A2(n6454), .B1(n9525), .B2(n6453), .C1(
        P1_U3086), .C2(n6580), .ZN(P1_U3353) );
  OAI222_X1 U8137 ( .A1(n9521), .A2(n6456), .B1(n9525), .B2(n6455), .C1(
        P1_U3086), .C2(n6585), .ZN(P1_U3352) );
  OAI222_X1 U8138 ( .A1(n9521), .A2(n6457), .B1(n9525), .B2(n6465), .C1(
        P1_U3086), .C2(n6581), .ZN(P1_U3354) );
  OAI222_X1 U8139 ( .A1(n9521), .A2(n5230), .B1(n9525), .B2(n6458), .C1(
        P1_U3086), .C2(n6587), .ZN(P1_U3351) );
  OAI222_X1 U8140 ( .A1(n7561), .A2(n6459), .B1(n8858), .B2(n6458), .C1(
        P2_U3151), .C2(n7135), .ZN(P2_U3291) );
  INV_X1 U8141 ( .A(n9521), .ZN(n6691) );
  AOI22_X1 U8142 ( .A1(n9110), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n6691), .ZN(n6460) );
  OAI21_X1 U8143 ( .B1(n6461), .B2(n9525), .A(n6460), .ZN(P1_U3350) );
  OAI222_X1 U8144 ( .A1(n7561), .A2(n6462), .B1(n8858), .B2(n6461), .C1(n7231), 
        .C2(P2_U3151), .ZN(P2_U3290) );
  AOI22_X1 U8145 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9563), .B1(n6691), .B2(
        P2_DATAO_REG_6__SCAN_IN), .ZN(n6463) );
  OAI21_X1 U8146 ( .B1(n6464), .B2(n9525), .A(n6463), .ZN(P1_U3349) );
  OAI222_X1 U8147 ( .A1(P2_U3151), .A2(n8420), .B1(n7561), .B2(n5939), .C1(
        n6464), .C2(n8858), .ZN(P2_U3289) );
  INV_X1 U8148 ( .A(n6535), .ZN(n8860) );
  OAI222_X1 U8149 ( .A1(n8860), .A2(n6466), .B1(n8858), .B2(n6465), .C1(
        P2_U3151), .C2(n6896), .ZN(P2_U3294) );
  AOI22_X1 U8150 ( .A1(n9123), .A2(P1_STATE_REG_SCAN_IN), .B1(n6691), .B2(
        P2_DATAO_REG_7__SCAN_IN), .ZN(n6467) );
  OAI21_X1 U8151 ( .B1(n6468), .B2(n9525), .A(n6467), .ZN(P1_U3348) );
  OAI222_X1 U8152 ( .A1(n7561), .A2(n4701), .B1(n8858), .B2(n6468), .C1(
        P2_U3151), .C2(n8454), .ZN(P2_U3288) );
  INV_X1 U8153 ( .A(n6469), .ZN(n6471) );
  AOI22_X1 U8154 ( .A1(n9550), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n6691), .ZN(n6470) );
  OAI21_X1 U8155 ( .B1(n6471), .B2(n9525), .A(n6470), .ZN(P1_U3347) );
  INV_X1 U8156 ( .A(n8489), .ZN(n9707) );
  OAI222_X1 U8157 ( .A1(n7561), .A2(n6472), .B1(n8858), .B2(n6471), .C1(
        P2_U3151), .C2(n9707), .ZN(P2_U3287) );
  NAND2_X1 U8158 ( .A1(n7807), .A2(n7819), .ZN(n6480) );
  OR2_X1 U8159 ( .A1(n7599), .A2(n6473), .ZN(n6475) );
  NAND2_X1 U8160 ( .A1(n6475), .A2(n6474), .ZN(n6478) );
  INV_X1 U8161 ( .A(n9590), .ZN(n9154) );
  NOR2_X1 U8162 ( .A1(n9154), .A2(P1_U3973), .ZN(P1_U3085) );
  INV_X1 U8163 ( .A(n9621), .ZN(n6477) );
  INV_X1 U8164 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6509) );
  NAND2_X1 U8165 ( .A1(n6477), .A2(n6666), .ZN(n6476) );
  OAI21_X1 U8166 ( .B1(n6477), .B2(n6509), .A(n6476), .ZN(P1_U3440) );
  INV_X1 U8167 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6484) );
  INV_X1 U8168 ( .A(n6478), .ZN(n6479) );
  AND2_X1 U8169 ( .A1(n6480), .A2(n6479), .ZN(n6599) );
  INV_X1 U8170 ( .A(n7891), .ZN(n9058) );
  INV_X1 U8171 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6672) );
  AOI21_X1 U8172 ( .B1(n9058), .B2(n6672), .A(n4353), .ZN(n9065) );
  OAI21_X1 U8173 ( .B1(n9058), .B2(P1_REG1_REG_0__SCAN_IN), .A(n9065), .ZN(
        n6481) );
  XNOR2_X1 U8174 ( .A(n6481), .B(P1_IR_REG_0__SCAN_IN), .ZN(n6482) );
  AOI22_X1 U8175 ( .A1(n6599), .A2(n6482), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n6483) );
  OAI21_X1 U8176 ( .B1(n9590), .B2(n6484), .A(n6483), .ZN(P1_U3243) );
  INV_X1 U8177 ( .A(n6485), .ZN(n6501) );
  AOI22_X1 U8178 ( .A1(n9142), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n6691), .ZN(n6486) );
  OAI21_X1 U8179 ( .B1(n6501), .B2(n9525), .A(n6486), .ZN(P1_U3346) );
  NAND2_X1 U8180 ( .A1(n6922), .A2(P1_U3973), .ZN(n6487) );
  OAI21_X1 U8181 ( .B1(P1_U3973), .B2(n5939), .A(n6487), .ZN(P1_U3560) );
  INV_X1 U8182 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8011) );
  INV_X1 U8183 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9171) );
  INV_X1 U8184 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n9370) );
  OR2_X1 U8185 ( .A1(n6488), .A2(n9370), .ZN(n6490) );
  INV_X1 U8186 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n9484) );
  OR2_X1 U8187 ( .A1(n6495), .A2(n9484), .ZN(n6489) );
  OAI211_X1 U8188 ( .C1(n6491), .C2(n9171), .A(n6490), .B(n6489), .ZN(n7893)
         );
  NAND2_X1 U8189 ( .A1(n7893), .A2(P1_U3973), .ZN(n6492) );
  OAI21_X1 U8190 ( .B1(n8011), .B2(P1_U3973), .A(n6492), .ZN(P1_U3584) );
  INV_X1 U8191 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6500) );
  INV_X1 U8192 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6498) );
  INV_X1 U8193 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9366) );
  OR2_X1 U8194 ( .A1(n6494), .A2(n9366), .ZN(n6497) );
  INV_X1 U8195 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9480) );
  OR2_X1 U8196 ( .A1(n6495), .A2(n9480), .ZN(n6496) );
  OAI211_X1 U8197 ( .C1(n6491), .C2(n6498), .A(n6497), .B(n6496), .ZN(n9163)
         );
  NAND2_X1 U8198 ( .A1(n9163), .A2(P1_U3973), .ZN(n6499) );
  OAI21_X1 U8199 ( .B1(P1_U3973), .B2(n6500), .A(n6499), .ZN(P1_U3585) );
  OAI222_X1 U8200 ( .A1(n7561), .A2(n6502), .B1(n8858), .B2(n6501), .C1(n4769), 
        .C2(P2_U3151), .ZN(P2_U3286) );
  INV_X1 U8201 ( .A(n6503), .ZN(n6507) );
  AOI22_X1 U8202 ( .A1(n9538), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n6691), .ZN(n6504) );
  OAI21_X1 U8203 ( .B1(n6507), .B2(n9525), .A(n6504), .ZN(P1_U3345) );
  AND2_X1 U8204 ( .A1(n6539), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U8205 ( .A1(n6539), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U8206 ( .A1(n6539), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U8207 ( .A1(n6539), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U8208 ( .A1(n6539), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U8209 ( .A1(n6539), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U8210 ( .A1(n6539), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U8211 ( .A1(n6539), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  AND2_X1 U8212 ( .A1(n6539), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U8213 ( .A1(n6539), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U8214 ( .A1(n6539), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U8215 ( .A1(n6539), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U8216 ( .A1(n6539), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  INV_X1 U8217 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6508) );
  OAI222_X1 U8218 ( .A1(n7561), .A2(n6508), .B1(n8858), .B2(n6507), .C1(n8481), 
        .C2(P2_U3151), .ZN(P2_U3285) );
  NAND2_X1 U8219 ( .A1(n6516), .A2(n6509), .ZN(n6510) );
  NAND2_X1 U8220 ( .A1(n6510), .A2(n6666), .ZN(n6519) );
  INV_X1 U8221 ( .A(n6667), .ZN(n6511) );
  OR2_X1 U8222 ( .A1(n6512), .A2(n6511), .ZN(n6513) );
  NOR2_X1 U8223 ( .A1(n6513), .A2(n7807), .ZN(n6518) );
  INV_X1 U8224 ( .A(n6514), .ZN(n6515) );
  NAND2_X1 U8225 ( .A1(n6516), .A2(n6515), .ZN(n6517) );
  INV_X1 U8226 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6529) );
  NOR2_X1 U8227 ( .A1(n9045), .A2(n6549), .ZN(n6625) );
  INV_X1 U8228 ( .A(n6625), .ZN(n6520) );
  NAND2_X1 U8229 ( .A1(n9045), .A2(n6549), .ZN(n7759) );
  AND2_X1 U8230 ( .A1(n6520), .A2(n7759), .ZN(n7605) );
  NAND2_X1 U8231 ( .A1(n6521), .A2(n7803), .ZN(n6674) );
  NAND2_X1 U8232 ( .A1(n6523), .A2(n6522), .ZN(n6524) );
  AND2_X1 U8233 ( .A1(n6524), .A2(n6673), .ZN(n6525) );
  NAND2_X1 U8234 ( .A1(n6674), .A2(n6525), .ZN(n6930) );
  OR2_X1 U8235 ( .A1(n7804), .A2(n7815), .ZN(n6526) );
  NAND2_X1 U8236 ( .A1(n5806), .A2(n6548), .ZN(n7811) );
  NOR2_X1 U8237 ( .A1(n9682), .A2(n9447), .ZN(n6527) );
  OAI222_X1 U8238 ( .A1(n6549), .A2(n6673), .B1(n7605), .B2(n6527), .C1(n9670), 
        .C2(n6855), .ZN(n9478) );
  NAND2_X1 U8239 ( .A1(n9478), .A2(n9685), .ZN(n6528) );
  OAI21_X1 U8240 ( .B1(n9685), .B2(n6529), .A(n6528), .ZN(P1_U3453) );
  INV_X1 U8241 ( .A(n6530), .ZN(n6532) );
  INV_X1 U8242 ( .A(n6596), .ZN(n9583) );
  OAI222_X1 U8243 ( .A1(n9521), .A2(n6531), .B1(n9525), .B2(n6532), .C1(
        P1_U3086), .C2(n9583), .ZN(P1_U3344) );
  OAI222_X1 U8244 ( .A1(n7561), .A2(n6533), .B1(n8858), .B2(n6532), .C1(
        P2_U3151), .C2(n8479), .ZN(P2_U3284) );
  INV_X1 U8245 ( .A(n6534), .ZN(n6538) );
  AOI22_X1 U8246 ( .A1(n9768), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n6535), .ZN(n6536) );
  OAI21_X1 U8247 ( .B1(n6538), .B2(n8858), .A(n6536), .ZN(P2_U3283) );
  INV_X1 U8248 ( .A(n6654), .ZN(n6601) );
  INV_X1 U8249 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6537) );
  OAI222_X1 U8250 ( .A1(n9525), .A2(n6538), .B1(n6601), .B2(P1_U3086), .C1(
        n6537), .C2(n9521), .ZN(P1_U3343) );
  INV_X1 U8251 ( .A(n6540), .ZN(n6541) );
  AOI22_X1 U8252 ( .A1(n6539), .A2(n4482), .B1(n6721), .B2(n6541), .ZN(
        P2_U3376) );
  INV_X1 U8253 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6544) );
  INV_X1 U8254 ( .A(n6542), .ZN(n6543) );
  AOI22_X1 U8255 ( .A1(n6539), .A2(n6544), .B1(n6721), .B2(n6543), .ZN(
        P2_U3377) );
  INV_X1 U8256 ( .A(n7604), .ZN(n6546) );
  NAND2_X1 U8257 ( .A1(n9045), .A2(n6680), .ZN(n6545) );
  NAND2_X1 U8258 ( .A1(n6546), .A2(n6545), .ZN(n6629) );
  OAI21_X1 U8259 ( .B1(n6546), .B2(n6545), .A(n6629), .ZN(n6818) );
  NAND2_X1 U8260 ( .A1(n6818), .A2(n9682), .ZN(n6551) );
  AOI22_X1 U8261 ( .A1(n9441), .A2(n9043), .B1(n9045), .B2(n9647), .ZN(n6550)
         );
  XNOR2_X1 U8262 ( .A(n7604), .B(n6625), .ZN(n6547) );
  NAND2_X1 U8263 ( .A1(n6547), .A2(n9447), .ZN(n6820) );
  INV_X2 U8264 ( .A(n4449), .ZN(n7757) );
  NAND2_X1 U8265 ( .A1(n7757), .A2(n6549), .ZN(n6633) );
  OAI211_X1 U8266 ( .C1(n7757), .C2(n6549), .A(n9603), .B(n6633), .ZN(n6814)
         );
  AND4_X1 U8267 ( .A1(n6551), .A2(n6550), .A3(n6820), .A4(n6814), .ZN(n6557)
         );
  OAI22_X1 U8268 ( .A1(n9515), .A2(n7757), .B1(n9685), .B2(n5147), .ZN(n6552)
         );
  INV_X1 U8269 ( .A(n6552), .ZN(n6553) );
  OAI21_X1 U8270 ( .B1(n6557), .B2(n9684), .A(n6553), .ZN(P1_U3456) );
  INV_X1 U8271 ( .A(n6668), .ZN(n6554) );
  INV_X1 U8272 ( .A(n9461), .ZN(n7193) );
  AOI22_X1 U8273 ( .A1(n7193), .A2(n4449), .B1(n9694), .B2(
        P1_REG1_REG_1__SCAN_IN), .ZN(n6556) );
  OAI21_X1 U8274 ( .B1(n6557), .B2(n9694), .A(n6556), .ZN(P1_U3523) );
  AND2_X1 U8275 ( .A1(n6539), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U8276 ( .A1(n6539), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U8277 ( .A1(n6539), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U8278 ( .A1(n6539), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U8279 ( .A1(n6539), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U8280 ( .A1(n6539), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U8281 ( .A1(n6539), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U8282 ( .A1(n6539), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U8283 ( .A1(n6539), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U8284 ( .A1(n6539), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U8285 ( .A1(n6539), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U8286 ( .A1(n6539), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U8287 ( .A1(n6539), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U8288 ( .A1(n6539), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U8289 ( .A1(n6539), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U8290 ( .A1(n6539), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U8291 ( .A1(n6539), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  INV_X1 U8292 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6558) );
  AOI22_X1 U8293 ( .A1(n6654), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n6558), .B2(
        n6601), .ZN(n6575) );
  NAND2_X1 U8294 ( .A1(n9538), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6559) );
  OAI21_X1 U8295 ( .B1(n9538), .B2(P1_REG2_REG_10__SCAN_IN), .A(n6559), .ZN(
        n9534) );
  NOR2_X1 U8296 ( .A1(n9142), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6560) );
  AOI21_X1 U8297 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n9142), .A(n6560), .ZN(
        n9135) );
  INV_X1 U8298 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6799) );
  MUX2_X1 U8299 ( .A(n6799), .B(P1_REG2_REG_2__SCAN_IN), .S(n6580), .Z(n9075)
         );
  INV_X1 U8300 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n6810) );
  MUX2_X1 U8301 ( .A(n6810), .B(P1_REG2_REG_1__SCAN_IN), .S(n6581), .Z(n9051)
         );
  AND2_X1 U8302 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n9059) );
  NAND2_X1 U8303 ( .A1(n9051), .A2(n9059), .ZN(n9050) );
  INV_X1 U8304 ( .A(n6581), .ZN(n9049) );
  NAND2_X1 U8305 ( .A1(n9049), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U8306 ( .A1(n9050), .A2(n6561), .ZN(n9074) );
  NAND2_X1 U8307 ( .A1(n9075), .A2(n9074), .ZN(n9073) );
  INV_X1 U8308 ( .A(n6580), .ZN(n9069) );
  NAND2_X1 U8309 ( .A1(n9069), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6562) );
  NAND2_X1 U8310 ( .A1(n9073), .A2(n6562), .ZN(n9087) );
  INV_X1 U8311 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6563) );
  MUX2_X1 U8312 ( .A(n6563), .B(P1_REG2_REG_3__SCAN_IN), .S(n6585), .Z(n9088)
         );
  NAND2_X1 U8313 ( .A1(n9087), .A2(n9088), .ZN(n9086) );
  INV_X1 U8314 ( .A(n6585), .ZN(n9082) );
  NAND2_X1 U8315 ( .A1(n9082), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6564) );
  NAND2_X1 U8316 ( .A1(n9086), .A2(n6564), .ZN(n9099) );
  XNOR2_X1 U8317 ( .A(n6587), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9098) );
  NAND2_X1 U8318 ( .A1(n9099), .A2(n9098), .ZN(n9097) );
  INV_X1 U8319 ( .A(n6587), .ZN(n9096) );
  NAND2_X1 U8320 ( .A1(n9096), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6565) );
  NAND2_X1 U8321 ( .A1(n9097), .A2(n6565), .ZN(n9115) );
  INV_X1 U8322 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6566) );
  MUX2_X1 U8323 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n6566), .S(n9110), .Z(n9116)
         );
  NAND2_X1 U8324 ( .A1(n9115), .A2(n9116), .ZN(n9114) );
  NAND2_X1 U8325 ( .A1(n9110), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6567) );
  NAND2_X1 U8326 ( .A1(n9114), .A2(n6567), .ZN(n9561) );
  INV_X1 U8327 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6705) );
  MUX2_X1 U8328 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n6705), .S(n9563), .Z(n9562)
         );
  NAND2_X1 U8329 ( .A1(n9561), .A2(n9562), .ZN(n9560) );
  NAND2_X1 U8330 ( .A1(n9563), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6568) );
  NAND2_X1 U8331 ( .A1(n9560), .A2(n6568), .ZN(n9128) );
  INV_X1 U8332 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6569) );
  XNOR2_X1 U8333 ( .A(n9123), .B(n6569), .ZN(n9129) );
  NAND2_X1 U8334 ( .A1(n9128), .A2(n9129), .ZN(n9127) );
  NAND2_X1 U8335 ( .A1(n9123), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6570) );
  NAND2_X1 U8336 ( .A1(n9127), .A2(n6570), .ZN(n9548) );
  OR2_X1 U8337 ( .A1(n9550), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6572) );
  NAND2_X1 U8338 ( .A1(n9550), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6571) );
  AND2_X1 U8339 ( .A1(n6572), .A2(n6571), .ZN(n9549) );
  AND2_X1 U8340 ( .A1(n9548), .A2(n9549), .ZN(n9546) );
  AOI21_X1 U8341 ( .B1(P1_REG2_REG_8__SCAN_IN), .B2(n9550), .A(n9546), .ZN(
        n9134) );
  NAND2_X1 U8342 ( .A1(n9135), .A2(n9134), .ZN(n9133) );
  OAI21_X1 U8343 ( .B1(n9142), .B2(P1_REG2_REG_9__SCAN_IN), .A(n9133), .ZN(
        n9535) );
  NOR2_X1 U8344 ( .A1(n9534), .A2(n9535), .ZN(n9533) );
  AOI21_X1 U8345 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(n9538), .A(n9533), .ZN(
        n9577) );
  INV_X1 U8346 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6573) );
  AOI22_X1 U8347 ( .A1(n6596), .A2(n6573), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n9583), .ZN(n9578) );
  NOR2_X1 U8348 ( .A1(n9577), .A2(n9578), .ZN(n9576) );
  AOI21_X1 U8349 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6596), .A(n9576), .ZN(
        n6574) );
  NAND2_X1 U8350 ( .A1(n6575), .A2(n6574), .ZN(n6649) );
  OAI21_X1 U8351 ( .B1(n6575), .B2(n6574), .A(n6649), .ZN(n6577) );
  NOR2_X1 U8352 ( .A1(n4353), .A2(n7891), .ZN(n6576) );
  NAND2_X1 U8353 ( .A1(n6577), .A2(n9580), .ZN(n6605) );
  NAND2_X1 U8354 ( .A1(n9538), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6578) );
  OAI21_X1 U8355 ( .B1(n9538), .B2(P1_REG1_REG_10__SCAN_IN), .A(n6578), .ZN(
        n9530) );
  NOR2_X1 U8356 ( .A1(n9142), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6579) );
  AOI21_X1 U8357 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n9142), .A(n6579), .ZN(
        n9139) );
  MUX2_X1 U8358 ( .A(n5182), .B(P1_REG1_REG_2__SCAN_IN), .S(n6580), .Z(n9072)
         );
  MUX2_X1 U8359 ( .A(n5146), .B(P1_REG1_REG_1__SCAN_IN), .S(n6581), .Z(n9054)
         );
  AND2_X1 U8360 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n9053) );
  NAND2_X1 U8361 ( .A1(n9054), .A2(n9053), .ZN(n9052) );
  NAND2_X1 U8362 ( .A1(n9049), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6582) );
  NAND2_X1 U8363 ( .A1(n9052), .A2(n6582), .ZN(n9071) );
  NAND2_X1 U8364 ( .A1(n9072), .A2(n9071), .ZN(n9070) );
  NAND2_X1 U8365 ( .A1(n9069), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6583) );
  NAND2_X1 U8366 ( .A1(n9070), .A2(n6583), .ZN(n9084) );
  MUX2_X1 U8367 ( .A(n6584), .B(P1_REG1_REG_3__SCAN_IN), .S(n6585), .Z(n9085)
         );
  NAND2_X1 U8368 ( .A1(n9084), .A2(n9085), .ZN(n9083) );
  OR2_X1 U8369 ( .A1(n6585), .A2(n6584), .ZN(n6586) );
  NAND2_X1 U8370 ( .A1(n9083), .A2(n6586), .ZN(n9102) );
  XNOR2_X1 U8371 ( .A(n6587), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n9101) );
  NAND2_X1 U8372 ( .A1(n9102), .A2(n9101), .ZN(n9100) );
  NAND2_X1 U8373 ( .A1(n9096), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6588) );
  NAND2_X1 U8374 ( .A1(n9100), .A2(n6588), .ZN(n9112) );
  MUX2_X1 U8375 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n5262), .S(n9110), .Z(n9113)
         );
  NAND2_X1 U8376 ( .A1(n9112), .A2(n9113), .ZN(n9111) );
  NAND2_X1 U8377 ( .A1(n9110), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6589) );
  NAND2_X1 U8378 ( .A1(n9111), .A2(n6589), .ZN(n9558) );
  MUX2_X1 U8379 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n5295), .S(n9563), .Z(n9559)
         );
  NAND2_X1 U8380 ( .A1(n9558), .A2(n9559), .ZN(n9557) );
  NAND2_X1 U8381 ( .A1(n9563), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6590) );
  NAND2_X1 U8382 ( .A1(n9557), .A2(n6590), .ZN(n9125) );
  XNOR2_X1 U8383 ( .A(n9123), .B(n6591), .ZN(n9126) );
  NAND2_X1 U8384 ( .A1(n9125), .A2(n9126), .ZN(n9124) );
  NAND2_X1 U8385 ( .A1(n9123), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6592) );
  NAND2_X1 U8386 ( .A1(n9124), .A2(n6592), .ZN(n9544) );
  OR2_X1 U8387 ( .A1(n9550), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6594) );
  NAND2_X1 U8388 ( .A1(n9550), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6593) );
  AND2_X1 U8389 ( .A1(n6594), .A2(n6593), .ZN(n9545) );
  AND2_X1 U8390 ( .A1(n9544), .A2(n9545), .ZN(n9542) );
  AOI21_X1 U8391 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n9550), .A(n9542), .ZN(
        n9138) );
  NAND2_X1 U8392 ( .A1(n9139), .A2(n9138), .ZN(n9137) );
  OAI21_X1 U8393 ( .B1(n9142), .B2(P1_REG1_REG_9__SCAN_IN), .A(n9137), .ZN(
        n9531) );
  NOR2_X1 U8394 ( .A1(n9530), .A2(n9531), .ZN(n9529) );
  AOI21_X1 U8395 ( .B1(n9538), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9529), .ZN(
        n9572) );
  MUX2_X1 U8396 ( .A(n6595), .B(P1_REG1_REG_11__SCAN_IN), .S(n6596), .Z(n9573)
         );
  NOR2_X1 U8397 ( .A1(n9572), .A2(n9573), .ZN(n9571) );
  AOI21_X1 U8398 ( .B1(P1_REG1_REG_11__SCAN_IN), .B2(n6596), .A(n9571), .ZN(
        n6598) );
  AOI22_X1 U8399 ( .A1(n6654), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n5438), .B2(
        n6601), .ZN(n6597) );
  NAND2_X1 U8400 ( .A1(n6598), .A2(n6597), .ZN(n6653) );
  OAI21_X1 U8401 ( .B1(n6598), .B2(n6597), .A(n6653), .ZN(n6603) );
  NAND2_X1 U8402 ( .A1(n6599), .A2(n7891), .ZN(n9528) );
  NAND2_X1 U8403 ( .A1(n6599), .A2(n4353), .ZN(n9584) );
  NAND2_X1 U8404 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7358) );
  NAND2_X1 U8405 ( .A1(n9154), .A2(P1_ADDR_REG_12__SCAN_IN), .ZN(n6600) );
  OAI211_X1 U8406 ( .C1(n9584), .C2(n6601), .A(n7358), .B(n6600), .ZN(n6602)
         );
  AOI21_X1 U8407 ( .B1(n6603), .B2(n9575), .A(n6602), .ZN(n6604) );
  NAND2_X1 U8408 ( .A1(n6605), .A2(n6604), .ZN(P1_U3255) );
  INV_X1 U8409 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n6614) );
  INV_X1 U8410 ( .A(n6606), .ZN(n6607) );
  OAI21_X1 U8411 ( .B1(P2_IR_REG_0__SCAN_IN), .B2(n6608), .A(n6607), .ZN(n6611) );
  NAND2_X1 U8412 ( .A1(n6609), .A2(n8529), .ZN(n6610) );
  AOI22_X1 U8413 ( .A1(n6611), .A2(n6610), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        P2_U3151), .ZN(n6613) );
  NAND2_X1 U8414 ( .A1(n9858), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n6612) );
  OAI211_X1 U8415 ( .C1(n7067), .C2(n6614), .A(n6613), .B(n6612), .ZN(P2_U3182) );
  XNOR2_X1 U8416 ( .A(n6616), .B(n6615), .ZN(n9060) );
  NOR2_X1 U8417 ( .A1(n6617), .A2(n7807), .ZN(n6856) );
  INV_X1 U8418 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6618) );
  OAI22_X1 U8419 ( .A1(n6856), .A2(n6618), .B1(n9008), .B2(n6855), .ZN(n6619)
         );
  AOI21_X1 U8420 ( .B1(n6680), .B2(n8958), .A(n6619), .ZN(n6620) );
  OAI21_X1 U8421 ( .B1(n8960), .B2(n9060), .A(n6620), .ZN(P1_U3232) );
  INV_X1 U8422 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6622) );
  INV_X1 U8423 ( .A(n6621), .ZN(n6623) );
  INV_X1 U8424 ( .A(n6747), .ZN(n6658) );
  OAI222_X1 U8425 ( .A1(n9521), .A2(n6622), .B1(n9525), .B2(n6623), .C1(
        P1_U3086), .C2(n6658), .ZN(P1_U3342) );
  INV_X1 U8426 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6624) );
  INV_X1 U8427 ( .A(n9787), .ZN(n8475) );
  OAI222_X1 U8428 ( .A1(n7561), .A2(n6624), .B1(n8858), .B2(n6623), .C1(
        P2_U3151), .C2(n8475), .ZN(P2_U3282) );
  NAND2_X1 U8429 ( .A1(n7604), .A2(n6625), .ZN(n6627) );
  NAND2_X1 U8430 ( .A1(n6855), .A2(n4449), .ZN(n6626) );
  NAND2_X1 U8431 ( .A1(n6855), .A2(n7757), .ZN(n6628) );
  OAI21_X1 U8432 ( .B1(n6632), .B2(n6631), .A(n6694), .ZN(n6806) );
  INV_X1 U8433 ( .A(n6806), .ZN(n6636) );
  AOI22_X1 U8434 ( .A1(n9647), .A2(n9044), .B1(n9042), .B2(n9441), .ZN(n6635)
         );
  AOI21_X1 U8435 ( .B1(n6633), .B2(n4354), .A(n9348), .ZN(n6634) );
  NAND2_X1 U8436 ( .A1(n6634), .A2(n6842), .ZN(n6803) );
  OAI211_X1 U8437 ( .C1(n6636), .C2(n9627), .A(n6635), .B(n6803), .ZN(n6637)
         );
  AOI21_X1 U8438 ( .B1(n9447), .B2(n6797), .A(n6637), .ZN(n6641) );
  INV_X1 U8439 ( .A(n4354), .ZN(n7758) );
  OAI22_X1 U8440 ( .A1(n9515), .A2(n7758), .B1(n9685), .B2(n5183), .ZN(n6638)
         );
  INV_X1 U8441 ( .A(n6638), .ZN(n6639) );
  OAI21_X1 U8442 ( .B1(n6641), .B2(n9684), .A(n6639), .ZN(P1_U3459) );
  AOI22_X1 U8443 ( .A1(n7193), .A2(n4354), .B1(n9694), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6640) );
  OAI21_X1 U8444 ( .B1(n6641), .B2(n9694), .A(n6640), .ZN(P1_U3524) );
  NAND2_X1 U8445 ( .A1(n8202), .A2(P2_U3893), .ZN(n6642) );
  OAI21_X1 U8446 ( .B1(P2_U3893), .B2(n5230), .A(n6642), .ZN(P2_U3495) );
  NAND2_X1 U8447 ( .A1(n6225), .A2(P2_U3893), .ZN(n6643) );
  OAI21_X1 U8448 ( .B1(P2_U3893), .B2(n5165), .A(n6643), .ZN(P2_U3491) );
  INV_X1 U8449 ( .A(n6644), .ZN(n6646) );
  INV_X1 U8450 ( .A(n7099), .ZN(n6752) );
  INV_X1 U8451 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6645) );
  OAI222_X1 U8452 ( .A1(n9525), .A2(n6646), .B1(n6752), .B2(P1_U3086), .C1(
        n6645), .C2(n9521), .ZN(P1_U3341) );
  INV_X1 U8453 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6647) );
  INV_X1 U8454 ( .A(n9805), .ZN(n8473) );
  OAI222_X1 U8455 ( .A1(n8860), .A2(n6647), .B1(n8858), .B2(n6646), .C1(n8473), 
        .C2(P2_U3151), .ZN(P2_U3281) );
  INV_X1 U8456 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6648) );
  AOI22_X1 U8457 ( .A1(n6747), .A2(n6648), .B1(P1_REG2_REG_13__SCAN_IN), .B2(
        n6658), .ZN(n6651) );
  OAI21_X1 U8458 ( .B1(n6654), .B2(P1_REG2_REG_12__SCAN_IN), .A(n6649), .ZN(
        n6650) );
  NOR2_X1 U8459 ( .A1(n6651), .A2(n6650), .ZN(n6741) );
  AOI21_X1 U8460 ( .B1(n6651), .B2(n6650), .A(n6741), .ZN(n6652) );
  NAND2_X1 U8461 ( .A1(n6652), .A2(n9580), .ZN(n6662) );
  AOI22_X1 U8462 ( .A1(n6747), .A2(n5470), .B1(P1_REG1_REG_13__SCAN_IN), .B2(
        n6658), .ZN(n6656) );
  OAI21_X1 U8463 ( .B1(n6654), .B2(P1_REG1_REG_12__SCAN_IN), .A(n6653), .ZN(
        n6655) );
  NOR2_X1 U8464 ( .A1(n6656), .A2(n6655), .ZN(n6746) );
  AOI21_X1 U8465 ( .B1(n6656), .B2(n6655), .A(n6746), .ZN(n6660) );
  NAND2_X1 U8466 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7375) );
  NAND2_X1 U8467 ( .A1(n9154), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n6657) );
  OAI211_X1 U8468 ( .C1(n9584), .C2(n6658), .A(n7375), .B(n6657), .ZN(n6659)
         );
  AOI21_X1 U8469 ( .B1(n6660), .B2(n9575), .A(n6659), .ZN(n6661) );
  NAND2_X1 U8470 ( .A1(n6662), .A2(n6661), .ZN(P1_U3256) );
  NAND2_X1 U8471 ( .A1(n6664), .A2(n6663), .ZN(n6665) );
  NAND2_X1 U8472 ( .A1(n9621), .A2(n6665), .ZN(n6670) );
  AND2_X1 U8473 ( .A1(n6667), .A2(n6666), .ZN(n6669) );
  NAND3_X1 U8474 ( .A1(n6670), .A2(n6669), .A3(n6668), .ZN(n6671) );
  NAND2_X1 U8475 ( .A1(n9342), .A2(n9441), .ZN(n9300) );
  INV_X2 U8476 ( .A(n7977), .ZN(n9610) );
  NOR2_X1 U8477 ( .A1(n9342), .A2(n6672), .ZN(n6678) );
  INV_X1 U8478 ( .A(n6673), .ZN(n6676) );
  INV_X1 U8479 ( .A(n6674), .ZN(n6675) );
  NOR4_X1 U8480 ( .A1(n4352), .A2(n7605), .A3(n6676), .A4(n6675), .ZN(n6677)
         );
  AOI211_X1 U8481 ( .C1(n9610), .C2(P1_REG3_REG_0__SCAN_IN), .A(n6678), .B(
        n6677), .ZN(n6682) );
  NOR2_X1 U8482 ( .A1(n9305), .A2(n9348), .ZN(n9161) );
  NOR2_X2 U8483 ( .A1(n4352), .A2(n6679), .ZN(n9600) );
  OAI21_X1 U8484 ( .B1(n9161), .B2(n9600), .A(n6680), .ZN(n6681) );
  OAI211_X1 U8485 ( .C1(n6855), .C2(n9300), .A(n6682), .B(n6681), .ZN(P1_U3293) );
  INV_X1 U8486 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6684) );
  INV_X1 U8487 ( .A(n6683), .ZN(n6685) );
  INV_X1 U8488 ( .A(n7094), .ZN(n7264) );
  OAI222_X1 U8489 ( .A1(n9521), .A2(n6684), .B1(n9525), .B2(n6685), .C1(
        P1_U3086), .C2(n7264), .ZN(P1_U3340) );
  INV_X1 U8490 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6686) );
  INV_X1 U8491 ( .A(n9823), .ZN(n8471) );
  OAI222_X1 U8492 ( .A1(n8860), .A2(n6686), .B1(n8858), .B2(n6685), .C1(
        P2_U3151), .C2(n8471), .ZN(P2_U3280) );
  INV_X1 U8493 ( .A(n6832), .ZN(n6769) );
  AND2_X1 U8494 ( .A1(n7992), .A2(n9957), .ZN(n9962) );
  INV_X1 U8495 ( .A(n9962), .ZN(n9948) );
  NAND2_X1 U8496 ( .A1(n6225), .A2(n6769), .ZN(n8181) );
  NAND2_X1 U8497 ( .A1(n8187), .A2(n8181), .ZN(n8344) );
  OAI21_X1 U8498 ( .B1(n9883), .B2(n9948), .A(n8344), .ZN(n6688) );
  OR2_X1 U8499 ( .A1(n9892), .A2(n9893), .ZN(n6822) );
  OAI211_X1 U8500 ( .C1(n9955), .C2(n6769), .A(n6688), .B(n6822), .ZN(n8765)
         );
  NAND2_X1 U8501 ( .A1(n8765), .A2(n9968), .ZN(n6689) );
  OAI21_X1 U8502 ( .B1(n5871), .B2(n9968), .A(n6689), .ZN(P2_U3390) );
  INV_X1 U8503 ( .A(n6690), .ZN(n6757) );
  AOI22_X1 U8504 ( .A1(n7287), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n6691), .ZN(n6692) );
  OAI21_X1 U8505 ( .B1(n6757), .B2(n9525), .A(n6692), .ZN(P1_U3339) );
  INV_X1 U8506 ( .A(n9043), .ZN(n6813) );
  NAND2_X1 U8507 ( .A1(n6813), .A2(n7758), .ZN(n6693) );
  NAND2_X1 U8508 ( .A1(n8966), .A2(n8891), .ZN(n6695) );
  INV_X1 U8509 ( .A(n9041), .ZN(n8890) );
  NAND2_X1 U8510 ( .A1(n8890), .A2(n9615), .ZN(n6696) );
  NAND2_X1 U8511 ( .A1(n6786), .A2(n6696), .ZN(n6862) );
  INV_X1 U8512 ( .A(n9040), .ZN(n6697) );
  INV_X1 U8513 ( .A(n9630), .ZN(n6865) );
  NAND2_X1 U8514 ( .A1(n6697), .A2(n6865), .ZN(n7649) );
  NAND2_X1 U8515 ( .A1(n9630), .A2(n9040), .ZN(n7764) );
  AND2_X1 U8516 ( .A1(n7649), .A2(n7764), .ZN(n7610) );
  INV_X1 U8517 ( .A(n7610), .ZN(n6861) );
  NAND2_X1 U8518 ( .A1(n6697), .A2(n9630), .ZN(n6698) );
  INV_X1 U8519 ( .A(n6783), .ZN(n6924) );
  NAND2_X1 U8520 ( .A1(n6924), .A2(n6922), .ZN(n7645) );
  INV_X1 U8521 ( .A(n7647), .ZN(n7654) );
  OAI21_X1 U8522 ( .B1(n6700), .B2(n6699), .A(n6926), .ZN(n6701) );
  INV_X1 U8523 ( .A(n6701), .ZN(n6761) );
  OR2_X1 U8524 ( .A1(n6702), .A2(n7815), .ZN(n6934) );
  NAND2_X1 U8525 ( .A1(n6930), .A2(n6934), .ZN(n6703) );
  NAND2_X1 U8526 ( .A1(n9342), .A2(n9647), .ZN(n9181) );
  INV_X1 U8527 ( .A(n9181), .ZN(n9296) );
  INV_X1 U8528 ( .A(n6778), .ZN(n6704) );
  OAI22_X1 U8529 ( .A1(n9342), .A2(n6705), .B1(n6704), .B2(n7977), .ZN(n6706)
         );
  AOI21_X1 U8530 ( .B1(n9296), .B2(n9040), .A(n6706), .ZN(n6707) );
  OAI21_X1 U8531 ( .B1(n7038), .B2(n9300), .A(n6707), .ZN(n6710) );
  INV_X1 U8532 ( .A(n9615), .ZN(n6788) );
  NAND2_X1 U8533 ( .A1(n6864), .A2(n9630), .ZN(n6863) );
  AOI21_X1 U8534 ( .B1(n6863), .B2(n6783), .A(n9348), .ZN(n6708) );
  NAND2_X1 U8535 ( .A1(n6708), .A2(n6936), .ZN(n6759) );
  NOR2_X1 U8536 ( .A1(n6759), .A2(n9305), .ZN(n6709) );
  AOI211_X1 U8537 ( .C1(n9600), .C2(n6783), .A(n6710), .B(n6709), .ZN(n6718)
         );
  NAND2_X1 U8538 ( .A1(n6813), .A2(n4354), .ZN(n6711) );
  NOR2_X1 U8539 ( .A1(n9042), .A2(n8891), .ZN(n6713) );
  NAND2_X1 U8540 ( .A1(n9042), .A2(n8891), .ZN(n7763) );
  NAND2_X1 U8541 ( .A1(n9041), .A2(n9615), .ZN(n7761) );
  NAND2_X1 U8542 ( .A1(n8890), .A2(n6788), .ZN(n7650) );
  NAND2_X1 U8543 ( .A1(n6715), .A2(n7764), .ZN(n6716) );
  NAND2_X1 U8544 ( .A1(n6716), .A2(n7649), .ZN(n6920) );
  XNOR2_X1 U8545 ( .A(n7609), .B(n6920), .ZN(n6763) );
  NAND2_X1 U8546 ( .A1(n6763), .A2(n9307), .ZN(n6717) );
  OAI211_X1 U8547 ( .C1(n6761), .C2(n9364), .A(n6718), .B(n6717), .ZN(P1_U3287) );
  XOR2_X1 U8548 ( .A(n6720), .B(n6719), .Z(n6726) );
  NAND2_X1 U8549 ( .A1(n6722), .A2(n6721), .ZN(n6768) );
  INV_X1 U8550 ( .A(n8162), .ZN(n8178) );
  AOI22_X1 U8551 ( .A1(n8157), .A2(n6225), .B1(n8170), .B2(n8409), .ZN(n6723)
         );
  OAI21_X1 U8552 ( .B1(n9912), .B2(n8178), .A(n6723), .ZN(n6724) );
  AOI21_X1 U8553 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n6768), .A(n6724), .ZN(
        n6725) );
  OAI21_X1 U8554 ( .B1(n8164), .B2(n6726), .A(n6725), .ZN(P2_U3162) );
  INV_X1 U8555 ( .A(n6728), .ZN(n6729) );
  AOI21_X1 U8556 ( .B1(n6730), .B2(n6727), .A(n6729), .ZN(n6734) );
  INV_X1 U8557 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9046) );
  OAI22_X1 U8558 ( .A1(n9026), .A2(n7757), .B1(n6856), .B2(n9046), .ZN(n6732)
         );
  INV_X1 U8559 ( .A(n9045), .ZN(n6815) );
  OAI22_X1 U8560 ( .A1(n6813), .A2(n9008), .B1(n8988), .B2(n6815), .ZN(n6731)
         );
  NOR2_X1 U8561 ( .A1(n6732), .A2(n6731), .ZN(n6733) );
  OAI21_X1 U8562 ( .B1(n6734), .B2(n8960), .A(n6733), .ZN(P1_U3222) );
  XOR2_X1 U8563 ( .A(n6736), .B(n6735), .Z(n6740) );
  AOI22_X1 U8564 ( .A1(n8157), .A2(n8410), .B1(n8170), .B2(n9881), .ZN(n6737)
         );
  OAI21_X1 U8565 ( .B1(n9904), .B2(n8178), .A(n6737), .ZN(n6738) );
  AOI21_X1 U8566 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n6768), .A(n6738), .ZN(
        n6739) );
  OAI21_X1 U8567 ( .B1(n6740), .B2(n8164), .A(n6739), .ZN(P2_U3177) );
  AOI21_X1 U8568 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n6747), .A(n6741), .ZN(
        n6744) );
  INV_X1 U8569 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6742) );
  AOI22_X1 U8570 ( .A1(n7099), .A2(n6742), .B1(P1_REG2_REG_14__SCAN_IN), .B2(
        n6752), .ZN(n6743) );
  NOR2_X1 U8571 ( .A1(n6744), .A2(n6743), .ZN(n7093) );
  AOI21_X1 U8572 ( .B1(n6744), .B2(n6743), .A(n7093), .ZN(n6745) );
  NAND2_X1 U8573 ( .A1(n6745), .A2(n9580), .ZN(n6756) );
  AOI21_X1 U8574 ( .B1(P1_REG1_REG_13__SCAN_IN), .B2(n6747), .A(n6746), .ZN(
        n6750) );
  AOI22_X1 U8575 ( .A1(n7099), .A2(n6748), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n6752), .ZN(n6749) );
  NOR2_X1 U8576 ( .A1(n6750), .A2(n6749), .ZN(n7098) );
  AOI21_X1 U8577 ( .B1(n6750), .B2(n6749), .A(n7098), .ZN(n6754) );
  NAND2_X1 U8578 ( .A1(P1_U3086), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n8865) );
  NAND2_X1 U8579 ( .A1(n9154), .A2(P1_ADDR_REG_14__SCAN_IN), .ZN(n6751) );
  OAI211_X1 U8580 ( .C1(n9584), .C2(n6752), .A(n8865), .B(n6751), .ZN(n6753)
         );
  AOI21_X1 U8581 ( .B1(n6754), .B2(n9575), .A(n6753), .ZN(n6755) );
  NAND2_X1 U8582 ( .A1(n6756), .A2(n6755), .ZN(P1_U3257) );
  INV_X1 U8583 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n6758) );
  OAI222_X1 U8584 ( .A1(n7561), .A2(n6758), .B1(n8858), .B2(n6757), .C1(n8469), 
        .C2(P2_U3151), .ZN(P2_U3279) );
  AOI22_X1 U8585 ( .A1(n9039), .A2(n9441), .B1(n9647), .B2(n9040), .ZN(n6760)
         );
  OAI211_X1 U8586 ( .C1(n6761), .C2(n9627), .A(n6760), .B(n6759), .ZN(n6762)
         );
  AOI21_X1 U8587 ( .B1(n6763), .B2(n9447), .A(n6762), .ZN(n6767) );
  AOI22_X1 U8588 ( .A1(n7193), .A2(n6783), .B1(n9694), .B2(
        P1_REG1_REG_6__SCAN_IN), .ZN(n6764) );
  OAI21_X1 U8589 ( .B1(n6767), .B2(n9694), .A(n6764), .ZN(P1_U3528) );
  OAI22_X1 U8590 ( .A1(n9515), .A2(n6924), .B1(n9685), .B2(n5294), .ZN(n6765)
         );
  INV_X1 U8591 ( .A(n6765), .ZN(n6766) );
  OAI21_X1 U8592 ( .B1(n6767), .B2(n9684), .A(n6766), .ZN(P1_U3471) );
  INV_X1 U8593 ( .A(n6768), .ZN(n6772) );
  INV_X1 U8594 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10082) );
  OAI22_X1 U8595 ( .A1(n8160), .A2(n9892), .B1(n8178), .B2(n6769), .ZN(n6770)
         );
  AOI21_X1 U8596 ( .B1(n8344), .B2(n4514), .A(n6770), .ZN(n6771) );
  OAI21_X1 U8597 ( .B1(n6772), .B2(n10082), .A(n6771), .ZN(P2_U3172) );
  NAND2_X1 U8598 ( .A1(n6774), .A2(n6773), .ZN(n6776) );
  XOR2_X1 U8599 ( .A(n6776), .B(n6775), .Z(n6785) );
  INV_X1 U8600 ( .A(n8988), .ZN(n8889) );
  NAND2_X1 U8601 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n9568) );
  INV_X1 U8602 ( .A(n9568), .ZN(n6777) );
  AOI21_X1 U8603 ( .B1(n8889), .B2(n9040), .A(n6777), .ZN(n6781) );
  NAND2_X1 U8604 ( .A1(n9022), .A2(n6778), .ZN(n6780) );
  NAND2_X1 U8605 ( .A1(n9018), .A2(n9039), .ZN(n6779) );
  NAND3_X1 U8606 ( .A1(n6781), .A2(n6780), .A3(n6779), .ZN(n6782) );
  AOI21_X1 U8607 ( .B1(n6783), .B2(n8958), .A(n6782), .ZN(n6784) );
  OAI21_X1 U8608 ( .B1(n6785), .B2(n8960), .A(n6784), .ZN(P1_U3239) );
  OAI21_X1 U8609 ( .B1(n6787), .B2(n7606), .A(n6786), .ZN(n9617) );
  AOI211_X1 U8610 ( .C1(n6788), .C2(n6840), .A(n9348), .B(n6864), .ZN(n9609)
         );
  XOR2_X1 U8611 ( .A(n7606), .B(n6789), .Z(n6790) );
  AOI222_X1 U8612 ( .A1(n9447), .A2(n6790), .B1(n9040), .B2(n9441), .C1(n9042), 
        .C2(n9647), .ZN(n9620) );
  INV_X1 U8613 ( .A(n9620), .ZN(n6791) );
  AOI211_X1 U8614 ( .C1(n9682), .C2(n9617), .A(n9609), .B(n6791), .ZN(n6796)
         );
  OAI22_X1 U8615 ( .A1(n9515), .A2(n9615), .B1(n9685), .B2(n5241), .ZN(n6792)
         );
  INV_X1 U8616 ( .A(n6792), .ZN(n6793) );
  OAI21_X1 U8617 ( .B1(n6796), .B2(n9684), .A(n6793), .ZN(P1_U3465) );
  OAI22_X1 U8618 ( .A1(n9461), .A2(n9615), .B1(n9696), .B2(n5240), .ZN(n6794)
         );
  INV_X1 U8619 ( .A(n6794), .ZN(n6795) );
  OAI21_X1 U8620 ( .B1(n6796), .B2(n9694), .A(n6795), .ZN(P1_U3526) );
  INV_X1 U8621 ( .A(n6797), .ZN(n6808) );
  INV_X1 U8622 ( .A(n9307), .ZN(n7220) );
  INV_X1 U8623 ( .A(n9364), .ZN(n9618) );
  NAND2_X1 U8624 ( .A1(n9600), .A2(n4354), .ZN(n6802) );
  INV_X1 U8625 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n9066) );
  NOR2_X1 U8626 ( .A1(n7977), .A2(n9066), .ZN(n6800) );
  AOI21_X1 U8627 ( .B1(n4352), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6800), .ZN(
        n6801) );
  OAI211_X1 U8628 ( .C1(n9300), .C2(n8966), .A(n6802), .B(n6801), .ZN(n6805)
         );
  OAI22_X1 U8629 ( .A1(n6855), .A2(n9181), .B1(n9305), .B2(n6803), .ZN(n6804)
         );
  AOI211_X1 U8630 ( .C1(n9618), .C2(n6806), .A(n6805), .B(n6804), .ZN(n6807)
         );
  OAI21_X1 U8631 ( .B1(n6808), .B2(n7220), .A(n6807), .ZN(P1_U3291) );
  NAND2_X1 U8632 ( .A1(n9600), .A2(n4449), .ZN(n6812) );
  AOI22_X1 U8633 ( .A1(n4352), .A2(P1_REG2_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(n9610), .ZN(n6811) );
  OAI211_X1 U8634 ( .C1(n9300), .C2(n6813), .A(n6812), .B(n6811), .ZN(n6817)
         );
  OAI22_X1 U8635 ( .A1(n6815), .A2(n9181), .B1(n9305), .B2(n6814), .ZN(n6816)
         );
  AOI211_X1 U8636 ( .C1(n9618), .C2(n6818), .A(n6817), .B(n6816), .ZN(n6819)
         );
  OAI21_X1 U8637 ( .B1(n4352), .B2(n6820), .A(n6819), .ZN(P1_U3292) );
  NAND3_X1 U8638 ( .A1(n8344), .A2(n6821), .A3(n9955), .ZN(n6823) );
  OAI211_X1 U8639 ( .C1(n10082), .C2(n8706), .A(n6823), .B(n6822), .ZN(n6830)
         );
  AOI21_X1 U8640 ( .B1(n6825), .B2(n6828), .A(n6824), .ZN(n6826) );
  NAND2_X1 U8641 ( .A1(n6830), .A2(n8710), .ZN(n6834) );
  AOI22_X1 U8642 ( .A1(P2_REG2_REG_0__SCAN_IN), .A2(n9910), .B1(n4350), .B2(
        n6832), .ZN(n6833) );
  NAND2_X1 U8643 ( .A1(n6834), .A2(n6833), .ZN(P2_U3233) );
  OAI21_X1 U8644 ( .B1(n6837), .B2(n6836), .A(n6835), .ZN(n6838) );
  INV_X1 U8645 ( .A(n6838), .ZN(n9626) );
  AOI222_X1 U8646 ( .A1(n9447), .A2(n6839), .B1(n9041), .B2(n9441), .C1(n9043), 
        .C2(n9647), .ZN(n9625) );
  MUX2_X1 U8647 ( .A(n6563), .B(n9625), .S(n9342), .Z(n6845) );
  INV_X1 U8648 ( .A(n6840), .ZN(n6841) );
  AOI211_X1 U8649 ( .C1(n9623), .C2(n6842), .A(n9348), .B(n6841), .ZN(n9622)
         );
  OAI22_X1 U8650 ( .A1(n9614), .A2(n8891), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n7977), .ZN(n6843) );
  AOI21_X1 U8651 ( .B1(n9608), .B2(n9622), .A(n6843), .ZN(n6844) );
  OAI211_X1 U8652 ( .C1(n9626), .C2(n9364), .A(n6845), .B(n6844), .ZN(P1_U3290) );
  INV_X1 U8653 ( .A(n6846), .ZN(n6848) );
  INV_X1 U8654 ( .A(n7833), .ZN(n7826) );
  OAI222_X1 U8655 ( .A1(n9521), .A2(n6847), .B1(n9525), .B2(n6848), .C1(
        P1_U3086), .C2(n7826), .ZN(P1_U3338) );
  INV_X1 U8656 ( .A(n9859), .ZN(n8468) );
  OAI222_X1 U8657 ( .A1(n8860), .A2(n6849), .B1(n8858), .B2(n6848), .C1(
        P2_U3151), .C2(n8468), .ZN(P2_U3278) );
  INV_X1 U8658 ( .A(n6851), .ZN(n6853) );
  NAND3_X1 U8659 ( .A1(n6853), .A2(n6728), .A3(n6852), .ZN(n6854) );
  AOI21_X1 U8660 ( .B1(n6850), .B2(n6854), .A(n8960), .ZN(n6859) );
  OAI22_X1 U8661 ( .A1(n6855), .A2(n8988), .B1(n9008), .B2(n8966), .ZN(n6858)
         );
  OAI22_X1 U8662 ( .A1(n9026), .A2(n7758), .B1(n6856), .B2(n9066), .ZN(n6857)
         );
  OR3_X1 U8663 ( .A1(n6859), .A2(n6858), .A3(n6857), .ZN(P1_U3237) );
  OAI21_X1 U8664 ( .B1(n6862), .B2(n6861), .A(n6860), .ZN(n9633) );
  OAI211_X1 U8665 ( .C1(n6864), .C2(n9630), .A(n6863), .B(n9603), .ZN(n9629)
         );
  AOI22_X1 U8666 ( .A1(n9600), .A2(n6865), .B1(n9610), .B2(n6882), .ZN(n6866)
         );
  OAI21_X1 U8667 ( .B1(n9629), .B2(n9305), .A(n6866), .ZN(n6869) );
  XNOR2_X1 U8668 ( .A(n7646), .B(n7610), .ZN(n6867) );
  OAI222_X1 U8669 ( .A1(n9670), .A2(n6923), .B1(n9672), .B2(n8890), .C1(n6867), 
        .C2(n9680), .ZN(n9631) );
  MUX2_X1 U8670 ( .A(n9631), .B(P1_REG2_REG_5__SCAN_IN), .S(n4352), .Z(n6868)
         );
  AOI211_X1 U8671 ( .C1(n9618), .C2(n9633), .A(n6869), .B(n6868), .ZN(n6870)
         );
  INV_X1 U8672 ( .A(n6870), .ZN(P1_U3288) );
  XOR2_X1 U8673 ( .A(n6874), .B(n6873), .Z(n8964) );
  NAND3_X1 U8674 ( .A1(n6872), .A2(n8964), .A3(n8962), .ZN(n8963) );
  NAND2_X1 U8675 ( .A1(n8963), .A2(n6875), .ZN(n6879) );
  XNOR2_X1 U8676 ( .A(n6877), .B(n6876), .ZN(n6878) );
  XNOR2_X1 U8677 ( .A(n6879), .B(n6878), .ZN(n6885) );
  OAI22_X1 U8678 ( .A1(n9026), .A2(n9630), .B1(n8890), .B2(n8988), .ZN(n6881)
         );
  NAND2_X1 U8679 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n9107) );
  OAI21_X1 U8680 ( .B1(n9008), .B2(n6923), .A(n9107), .ZN(n6880) );
  NOR2_X1 U8681 ( .A1(n6881), .A2(n6880), .ZN(n6884) );
  NAND2_X1 U8682 ( .A1(n9022), .A2(n6882), .ZN(n6883) );
  OAI211_X1 U8683 ( .C1(n6885), .C2(n8960), .A(n6884), .B(n6883), .ZN(P1_U3227) );
  XOR2_X1 U8684 ( .A(n6888), .B(n6887), .Z(n6889) );
  XNOR2_X1 U8685 ( .A(n6886), .B(n6889), .ZN(n6894) );
  NAND2_X1 U8686 ( .A1(n9018), .A2(n9646), .ZN(n6890) );
  NAND2_X1 U8687 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n9120) );
  OAI211_X1 U8688 ( .C1(n6923), .C2(n8988), .A(n6890), .B(n9120), .ZN(n6892)
         );
  INV_X1 U8689 ( .A(n7031), .ZN(n9636) );
  NOR2_X1 U8690 ( .A1(n9026), .A2(n9636), .ZN(n6891) );
  AOI211_X1 U8691 ( .C1(n6938), .C2(n9022), .A(n6892), .B(n6891), .ZN(n6893)
         );
  OAI21_X1 U8692 ( .B1(n6894), .B2(n8960), .A(n6893), .ZN(P1_U3213) );
  INV_X1 U8693 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n6919) );
  MUX2_X1 U8694 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n8856), .Z(n6898) );
  AOI21_X1 U8695 ( .B1(n6897), .B2(n6896), .A(n6895), .ZN(n7052) );
  XNOR2_X1 U8696 ( .A(n6898), .B(n7062), .ZN(n7053) );
  NOR2_X1 U8697 ( .A1(n7052), .A2(n7053), .ZN(n7051) );
  MUX2_X1 U8698 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n8856), .Z(n6993) );
  XNOR2_X1 U8699 ( .A(n6993), .B(n4779), .ZN(n6899) );
  NAND2_X1 U8700 ( .A1(n6900), .A2(n6899), .ZN(n6991) );
  OAI21_X1 U8701 ( .B1(n6900), .B2(n6899), .A(n6991), .ZN(n6901) );
  NAND2_X1 U8702 ( .A1(n6901), .A2(n9866), .ZN(n6918) );
  INV_X1 U8703 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6902) );
  MUX2_X1 U8704 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6902), .S(n7062), .Z(n7059)
         );
  NAND2_X1 U8705 ( .A1(n6903), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6905) );
  NAND2_X1 U8706 ( .A1(n6905), .A2(n6904), .ZN(n7058) );
  NAND2_X1 U8707 ( .A1(n7062), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6906) );
  NAND2_X1 U8708 ( .A1(n7057), .A2(n6906), .ZN(n6975) );
  XNOR2_X1 U8709 ( .A(n6975), .B(n4779), .ZN(n6974) );
  XNOR2_X1 U8710 ( .A(n6974), .B(P2_REG1_REG_3__SCAN_IN), .ZN(n6916) );
  NOR2_X1 U8711 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5901), .ZN(n6949) );
  INV_X1 U8712 ( .A(n6949), .ZN(n6907) );
  OAI21_X1 U8713 ( .B1(n9708), .B2(n6992), .A(n6907), .ZN(n6915) );
  NAND2_X1 U8714 ( .A1(n6910), .A2(n6909), .ZN(n7055) );
  NAND2_X1 U8715 ( .A1(n7056), .A2(n7055), .ZN(n7054) );
  NAND2_X1 U8716 ( .A1(n7062), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6911) );
  NAND2_X1 U8717 ( .A1(n6912), .A2(n5888), .ZN(n6913) );
  AOI21_X1 U8718 ( .B1(n6985), .B2(n6913), .A(n9872), .ZN(n6914) );
  AOI211_X1 U8719 ( .C1(n9867), .C2(n6916), .A(n6915), .B(n6914), .ZN(n6917)
         );
  OAI211_X1 U8720 ( .C1(n7067), .C2(n6919), .A(n6918), .B(n6917), .ZN(P2_U3185) );
  OR2_X1 U8721 ( .A1(n7031), .A2(n7038), .ZN(n7074) );
  NAND2_X1 U8722 ( .A1(n7031), .A2(n7038), .ZN(n7072) );
  NAND2_X1 U8723 ( .A1(n7755), .A2(n7645), .ZN(n6921) );
  NOR2_X1 U8724 ( .A1(n6921), .A2(n6927), .ZN(n7108) );
  AOI21_X1 U8725 ( .B1(n6927), .B2(n6921), .A(n7108), .ZN(n6933) );
  AOI22_X1 U8726 ( .A1(n9646), .A2(n9441), .B1(n9647), .B2(n6922), .ZN(n6932)
         );
  NAND2_X1 U8727 ( .A1(n6924), .A2(n6923), .ZN(n6925) );
  OR2_X1 U8728 ( .A1(n6928), .A2(n6927), .ZN(n6929) );
  NAND2_X1 U8729 ( .A1(n7033), .A2(n6929), .ZN(n9639) );
  INV_X1 U8730 ( .A(n6930), .ZN(n9598) );
  NAND2_X1 U8731 ( .A1(n9639), .A2(n9598), .ZN(n6931) );
  OAI211_X1 U8732 ( .C1(n6933), .C2(n9680), .A(n6932), .B(n6931), .ZN(n9637)
         );
  INV_X1 U8733 ( .A(n9637), .ZN(n6943) );
  INV_X1 U8734 ( .A(n6934), .ZN(n6935) );
  AND2_X1 U8735 ( .A1(n9342), .A2(n6935), .ZN(n9605) );
  AOI21_X1 U8736 ( .B1(n6936), .B2(n7031), .A(n9348), .ZN(n6937) );
  NAND2_X1 U8737 ( .A1(n6937), .A2(n7043), .ZN(n9635) );
  AOI22_X1 U8738 ( .A1(n4352), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n6938), .B2(
        n9610), .ZN(n6940) );
  NAND2_X1 U8739 ( .A1(n9600), .A2(n7031), .ZN(n6939) );
  OAI211_X1 U8740 ( .C1(n9635), .C2(n9305), .A(n6940), .B(n6939), .ZN(n6941)
         );
  AOI21_X1 U8741 ( .B1(n9639), .B2(n9605), .A(n6941), .ZN(n6942) );
  OAI21_X1 U8742 ( .B1(n6943), .B2(n4352), .A(n6942), .ZN(P1_U3286) );
  AOI211_X1 U8743 ( .C1(n6946), .C2(n6945), .A(n8164), .B(n6944), .ZN(n6947)
         );
  INV_X1 U8744 ( .A(n6947), .ZN(n6951) );
  OAI22_X1 U8745 ( .A1(n8160), .A2(n7168), .B1(n8191), .B2(n8178), .ZN(n6948)
         );
  AOI211_X1 U8746 ( .C1(n8157), .C2(n8409), .A(n6949), .B(n6948), .ZN(n6950)
         );
  OAI211_X1 U8747 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8149), .A(n6951), .B(
        n6950), .ZN(P2_U3158) );
  INV_X1 U8748 ( .A(n8521), .ZN(n8513) );
  INV_X1 U8749 ( .A(n6952), .ZN(n6954) );
  INV_X1 U8750 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6953) );
  OAI222_X1 U8751 ( .A1(P2_U3151), .A2(n8513), .B1(n8858), .B2(n6954), .C1(
        n6953), .C2(n8860), .ZN(P2_U3277) );
  INV_X1 U8752 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6955) );
  INV_X1 U8753 ( .A(n7836), .ZN(n9151) );
  OAI222_X1 U8754 ( .A1(n9521), .A2(n6955), .B1(n9151), .B2(P1_U3086), .C1(
        n9525), .C2(n6954), .ZN(P1_U3337) );
  AOI21_X1 U8755 ( .B1(n6957), .B2(n6956), .A(n4443), .ZN(n6964) );
  NAND2_X1 U8756 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n9554) );
  INV_X1 U8757 ( .A(n9554), .ZN(n6958) );
  AOI21_X1 U8758 ( .B1(n8889), .B2(n9039), .A(n6958), .ZN(n6961) );
  NAND2_X1 U8759 ( .A1(n9022), .A2(n7046), .ZN(n6960) );
  NAND2_X1 U8760 ( .A1(n9018), .A2(n9038), .ZN(n6959) );
  NAND3_X1 U8761 ( .A1(n6961), .A2(n6960), .A3(n6959), .ZN(n6962) );
  AOI21_X1 U8762 ( .B1(n7080), .B2(n8958), .A(n6962), .ZN(n6963) );
  OAI21_X1 U8763 ( .B1(n6964), .B2(n8960), .A(n6963), .ZN(P1_U3221) );
  XOR2_X1 U8764 ( .A(n6965), .B(n8347), .Z(n6966) );
  AOI222_X1 U8765 ( .A1(n9883), .A2(n6966), .B1(n8202), .B2(n9878), .C1(n8409), 
        .C2(n9880), .ZN(n9923) );
  XNOR2_X1 U8766 ( .A(n6967), .B(n8347), .ZN(n9921) );
  NOR2_X1 U8767 ( .A1(n9906), .A2(n7180), .ZN(n7172) );
  INV_X1 U8768 ( .A(n7172), .ZN(n6968) );
  NAND2_X1 U8769 ( .A1(n6968), .A2(n7992), .ZN(n6969) );
  AOI22_X1 U8770 ( .A1(n4350), .A2(n9920), .B1(n5901), .B2(n9905), .ZN(n6970)
         );
  OAI21_X1 U8771 ( .B1(n5888), .B2(n8710), .A(n6970), .ZN(n6971) );
  AOI21_X1 U8772 ( .B1(n9921), .B2(n9888), .A(n6971), .ZN(n6972) );
  OAI21_X1 U8773 ( .B1(n9923), .B2(n9910), .A(n6972), .ZN(P2_U3230) );
  MUX2_X1 U8774 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6973), .S(n7135), .Z(n6979)
         );
  NAND2_X1 U8775 ( .A1(n6974), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6977) );
  NAND2_X1 U8776 ( .A1(n6975), .A2(n6992), .ZN(n6976) );
  NAND2_X1 U8777 ( .A1(n6977), .A2(n6976), .ZN(n6978) );
  NAND2_X1 U8778 ( .A1(n6978), .A2(n6979), .ZN(n7125) );
  OAI21_X1 U8779 ( .B1(n6979), .B2(n6978), .A(n7125), .ZN(n6988) );
  NAND2_X1 U8780 ( .A1(n6985), .A2(n6983), .ZN(n6981) );
  XNOR2_X1 U8781 ( .A(n7135), .B(n6980), .ZN(n6982) );
  INV_X1 U8782 ( .A(n6982), .ZN(n6984) );
  NAND3_X1 U8783 ( .A1(n6985), .A2(n6984), .A3(n6983), .ZN(n6986) );
  AOI21_X1 U8784 ( .B1(n7127), .B2(n6986), .A(n9872), .ZN(n6987) );
  AOI21_X1 U8785 ( .B1(n9867), .B2(n6988), .A(n6987), .ZN(n6990) );
  NOR2_X1 U8786 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5900), .ZN(n7028) );
  INV_X1 U8787 ( .A(n7028), .ZN(n6989) );
  OAI211_X1 U8788 ( .C1(n9708), .C2(n7135), .A(n6990), .B(n6989), .ZN(n6997)
         );
  MUX2_X1 U8789 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n8856), .Z(n7136) );
  XNOR2_X1 U8790 ( .A(n7136), .B(n7135), .ZN(n6995) );
  OAI21_X1 U8791 ( .B1(n6993), .B2(n6992), .A(n6991), .ZN(n6994) );
  AOI211_X1 U8792 ( .C1(n6995), .C2(n6994), .A(n8529), .B(n7134), .ZN(n6996)
         );
  AOI211_X1 U8793 ( .C1(n9857), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6997), .B(
        n6996), .ZN(n6998) );
  INV_X1 U8794 ( .A(n6998), .ZN(P2_U3186) );
  INV_X1 U8795 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n7009) );
  INV_X1 U8796 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7004) );
  NAND2_X1 U8797 ( .A1(n6999), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n7002) );
  INV_X1 U8798 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n7000) );
  OR2_X1 U8799 ( .A1(n5878), .A2(n7000), .ZN(n7001) );
  OAI211_X1 U8800 ( .C1(n7004), .C2(n7003), .A(n7002), .B(n7001), .ZN(n7005)
         );
  INV_X1 U8801 ( .A(n7005), .ZN(n7006) );
  NAND2_X1 U8802 ( .A1(n8536), .A2(P2_U3893), .ZN(n7008) );
  OAI21_X1 U8803 ( .B1(P2_U3893), .B2(n7009), .A(n7008), .ZN(P2_U3522) );
  OAI21_X1 U8804 ( .B1(n7013), .B2(n7010), .A(n7012), .ZN(n7014) );
  NAND2_X1 U8805 ( .A1(n7014), .A2(n9016), .ZN(n7021) );
  NAND2_X1 U8806 ( .A1(n8889), .A2(n9646), .ZN(n7017) );
  NOR2_X1 U8807 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7015), .ZN(n9141) );
  INV_X1 U8808 ( .A(n9141), .ZN(n7016) );
  OAI211_X1 U8809 ( .C1(n9592), .C2(n9008), .A(n7017), .B(n7016), .ZN(n7019)
         );
  INV_X1 U8810 ( .A(n9648), .ZN(n7116) );
  NOR2_X1 U8811 ( .A1(n7116), .A2(n9026), .ZN(n7018) );
  AOI211_X1 U8812 ( .C1(n7112), .C2(n9022), .A(n7019), .B(n7018), .ZN(n7020)
         );
  NAND2_X1 U8813 ( .A1(n7021), .A2(n7020), .ZN(P1_U3231) );
  OAI21_X1 U8814 ( .B1(n7024), .B2(n7023), .A(n7022), .ZN(n7025) );
  NAND2_X1 U8815 ( .A1(n7025), .A2(n4514), .ZN(n7030) );
  INV_X1 U8816 ( .A(n9924), .ZN(n8201) );
  OAI22_X1 U8817 ( .A1(n8160), .A2(n7026), .B1(n8201), .B2(n8178), .ZN(n7027)
         );
  AOI211_X1 U8818 ( .C1(n8157), .C2(n9881), .A(n7028), .B(n7027), .ZN(n7029)
         );
  OAI211_X1 U8819 ( .C1(n9886), .C2(n8149), .A(n7030), .B(n7029), .ZN(P2_U3170) );
  OR2_X1 U8820 ( .A1(n7031), .A2(n9039), .ZN(n7032) );
  XNOR2_X1 U8821 ( .A(n7080), .B(n7114), .ZN(n7035) );
  XNOR2_X1 U8822 ( .A(n7081), .B(n7035), .ZN(n9643) );
  NAND2_X1 U8823 ( .A1(n9643), .A2(n9598), .ZN(n7042) );
  INV_X1 U8824 ( .A(n7072), .ZN(n7034) );
  OR2_X1 U8825 ( .A1(n7108), .A2(n7034), .ZN(n7037) );
  INV_X1 U8826 ( .A(n7035), .ZN(n7036) );
  XNOR2_X1 U8827 ( .A(n7037), .B(n7036), .ZN(n7040) );
  OAI22_X1 U8828 ( .A1(n7038), .A2(n9672), .B1(n9655), .B2(n9670), .ZN(n7039)
         );
  AOI21_X1 U8829 ( .B1(n7040), .B2(n9447), .A(n7039), .ZN(n7041) );
  INV_X1 U8830 ( .A(n7117), .ZN(n7045) );
  AOI21_X1 U8831 ( .B1(n7043), .B2(n7080), .A(n9348), .ZN(n7044) );
  NAND2_X1 U8832 ( .A1(n7045), .A2(n7044), .ZN(n9640) );
  AOI22_X1 U8833 ( .A1(n4352), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n7046), .B2(
        n9610), .ZN(n7048) );
  NAND2_X1 U8834 ( .A1(n9600), .A2(n7080), .ZN(n7047) );
  OAI211_X1 U8835 ( .C1(n9640), .C2(n9305), .A(n7048), .B(n7047), .ZN(n7049)
         );
  AOI21_X1 U8836 ( .B1(n9643), .B2(n9605), .A(n7049), .ZN(n7050) );
  OAI21_X1 U8837 ( .B1(n9645), .B2(n4352), .A(n7050), .ZN(P1_U3285) );
  AOI211_X1 U8838 ( .C1(n7053), .C2(n7052), .A(n8529), .B(n7051), .ZN(n7069)
         );
  INV_X1 U8839 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7066) );
  INV_X1 U8840 ( .A(n9872), .ZN(n9798) );
  OAI21_X1 U8841 ( .B1(n7056), .B2(n7055), .A(n7054), .ZN(n7061) );
  OAI21_X1 U8842 ( .B1(n7059), .B2(n7058), .A(n7057), .ZN(n7060) );
  AOI22_X1 U8843 ( .A1(n9798), .A2(n7061), .B1(n9867), .B2(n7060), .ZN(n7065)
         );
  INV_X1 U8844 ( .A(n7062), .ZN(n7063) );
  AOI22_X1 U8845 ( .A1(n9858), .A2(n7063), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n7064) );
  OAI211_X1 U8846 ( .C1(n7067), .C2(n7066), .A(n7065), .B(n7064), .ZN(n7068)
         );
  OR2_X1 U8847 ( .A1(n7069), .A2(n7068), .ZN(P2_U3184) );
  INV_X1 U8848 ( .A(n7070), .ZN(n7566) );
  OAI222_X1 U8849 ( .A1(n8860), .A2(n7071), .B1(n8858), .B2(n7566), .C1(
        P2_U3151), .C2(n8526), .ZN(P2_U3276) );
  OR2_X1 U8850 ( .A1(n9658), .A2(n9592), .ZN(n7680) );
  NAND2_X1 U8851 ( .A1(n9658), .A2(n9592), .ZN(n7674) );
  NAND2_X1 U8852 ( .A1(n7680), .A2(n7674), .ZN(n7617) );
  NAND2_X1 U8853 ( .A1(n9648), .A2(n9655), .ZN(n7673) );
  NAND2_X1 U8854 ( .A1(n7080), .A2(n7114), .ZN(n7663) );
  NAND2_X1 U8855 ( .A1(n7663), .A2(n7072), .ZN(n7658) );
  INV_X1 U8856 ( .A(n7658), .ZN(n7614) );
  NAND2_X1 U8857 ( .A1(n7673), .A2(n7614), .ZN(n7077) );
  OR2_X1 U8858 ( .A1(n9648), .A2(n9655), .ZN(n7668) );
  OR2_X1 U8859 ( .A1(n7080), .A2(n7114), .ZN(n7107) );
  NAND2_X1 U8860 ( .A1(n7668), .A2(n7107), .ZN(n7665) );
  OR2_X1 U8861 ( .A1(n7665), .A2(n7614), .ZN(n7073) );
  AND2_X1 U8862 ( .A1(n7073), .A2(n7673), .ZN(n7767) );
  NAND2_X1 U8863 ( .A1(n7107), .A2(n7074), .ZN(n7659) );
  INV_X1 U8864 ( .A(n7659), .ZN(n7075) );
  NAND3_X1 U8865 ( .A1(n7668), .A2(n7075), .A3(n7645), .ZN(n7076) );
  NAND2_X1 U8866 ( .A1(n7767), .A2(n7076), .ZN(n7770) );
  OAI21_X1 U8867 ( .B1(n7755), .B2(n7077), .A(n7770), .ZN(n7079) );
  INV_X1 U8868 ( .A(n7186), .ZN(n7078) );
  AOI21_X1 U8869 ( .B1(n7617), .B2(n7079), .A(n7078), .ZN(n9660) );
  INV_X1 U8870 ( .A(n7080), .ZN(n9641) );
  NAND2_X1 U8871 ( .A1(n7081), .A2(n9641), .ZN(n7082) );
  NAND2_X1 U8872 ( .A1(n7083), .A2(n7082), .ZN(n7110) );
  NAND2_X1 U8873 ( .A1(n7110), .A2(n7111), .ZN(n7085) );
  OR2_X1 U8874 ( .A1(n9648), .A2(n9038), .ZN(n7084) );
  NAND2_X1 U8875 ( .A1(n7085), .A2(n7084), .ZN(n7183) );
  XNOR2_X1 U8876 ( .A(n7183), .B(n7617), .ZN(n9662) );
  NAND2_X1 U8877 ( .A1(n9662), .A2(n9618), .ZN(n7092) );
  AOI211_X1 U8878 ( .C1(n9658), .C2(n7115), .A(n9348), .B(n4372), .ZN(n9656)
         );
  INV_X1 U8879 ( .A(n9658), .ZN(n7086) );
  NOR2_X1 U8880 ( .A1(n7086), .A2(n9614), .ZN(n7090) );
  NAND2_X1 U8881 ( .A1(n9296), .A2(n9038), .ZN(n7088) );
  AOI22_X1 U8882 ( .A1(n4352), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n7250), .B2(
        n9610), .ZN(n7087) );
  OAI211_X1 U8883 ( .C1(n9654), .C2(n9300), .A(n7088), .B(n7087), .ZN(n7089)
         );
  AOI211_X1 U8884 ( .C1(n9656), .C2(n9608), .A(n7090), .B(n7089), .ZN(n7091)
         );
  OAI211_X1 U8885 ( .C1(n9660), .C2(n7220), .A(n7092), .B(n7091), .ZN(P1_U3283) );
  INV_X1 U8886 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7096) );
  AOI21_X1 U8887 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7099), .A(n7093), .ZN(
        n7265) );
  XOR2_X1 U8888 ( .A(n7094), .B(n7265), .Z(n7095) );
  NOR2_X1 U8889 ( .A1(n7096), .A2(n7095), .ZN(n7266) );
  AOI21_X1 U8890 ( .B1(n7096), .B2(n7095), .A(n7266), .ZN(n7097) );
  NAND2_X1 U8891 ( .A1(n7097), .A2(n9580), .ZN(n7106) );
  AOI21_X1 U8892 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n7099), .A(n7098), .ZN(
        n7257) );
  XNOR2_X1 U8893 ( .A(n7264), .B(n7257), .ZN(n7100) );
  NOR2_X1 U8894 ( .A1(n7101), .A2(n7100), .ZN(n7258) );
  AOI21_X1 U8895 ( .B1(n7101), .B2(n7100), .A(n7258), .ZN(n7104) );
  NAND2_X1 U8896 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9019) );
  NAND2_X1 U8897 ( .A1(n9154), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n7102) );
  OAI211_X1 U8898 ( .C1(n9584), .C2(n7264), .A(n9019), .B(n7102), .ZN(n7103)
         );
  AOI21_X1 U8899 ( .B1(n7104), .B2(n9575), .A(n7103), .ZN(n7105) );
  NAND2_X1 U8900 ( .A1(n7106), .A2(n7105), .ZN(P1_U3258) );
  OAI21_X1 U8901 ( .B1(n7108), .B2(n7658), .A(n7107), .ZN(n7109) );
  XNOR2_X1 U8902 ( .A(n7109), .B(n7615), .ZN(n9651) );
  XNOR2_X1 U8903 ( .A(n7110), .B(n7111), .ZN(n9653) );
  NAND2_X1 U8904 ( .A1(n9653), .A2(n9618), .ZN(n7123) );
  AOI22_X1 U8905 ( .A1(n4352), .A2(P1_REG2_REG_9__SCAN_IN), .B1(n7112), .B2(
        n9610), .ZN(n7113) );
  OAI21_X1 U8906 ( .B1(n9181), .B2(n7114), .A(n7113), .ZN(n7121) );
  OAI211_X1 U8907 ( .C1(n7117), .C2(n7116), .A(n7115), .B(n9603), .ZN(n7119)
         );
  NAND2_X1 U8908 ( .A1(n9037), .A2(n9441), .ZN(n7118) );
  AND2_X1 U8909 ( .A1(n7119), .A2(n7118), .ZN(n9650) );
  NOR2_X1 U8910 ( .A1(n9650), .A2(n9305), .ZN(n7120) );
  AOI211_X1 U8911 ( .C1(n9600), .C2(n9648), .A(n7121), .B(n7120), .ZN(n7122)
         );
  OAI211_X1 U8912 ( .C1(n9651), .C2(n7220), .A(n7123), .B(n7122), .ZN(P1_U3284) );
  NAND2_X1 U8913 ( .A1(n7135), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7124) );
  INV_X1 U8914 ( .A(n7231), .ZN(n7130) );
  XNOR2_X1 U8915 ( .A(n7232), .B(n7130), .ZN(n7230) );
  XNOR2_X1 U8916 ( .A(n7230), .B(P2_REG1_REG_5__SCAN_IN), .ZN(n7141) );
  NAND2_X1 U8917 ( .A1(n7135), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n7126) );
  NAND2_X1 U8918 ( .A1(n7128), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n8417) );
  OAI21_X1 U8919 ( .B1(n7128), .B2(P2_REG2_REG_5__SCAN_IN), .A(n8417), .ZN(
        n7129) );
  INV_X1 U8920 ( .A(n7129), .ZN(n7133) );
  NAND2_X1 U8921 ( .A1(n9857), .A2(P2_ADDR_REG_5__SCAN_IN), .ZN(n7132) );
  NOR2_X1 U8922 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10168), .ZN(n7149) );
  AOI21_X1 U8923 ( .B1(n9858), .B2(n7130), .A(n7149), .ZN(n7131) );
  OAI211_X1 U8924 ( .C1(n7133), .C2(n9872), .A(n7132), .B(n7131), .ZN(n7140)
         );
  MUX2_X1 U8925 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n8856), .Z(n7223) );
  XNOR2_X1 U8926 ( .A(n7223), .B(n7231), .ZN(n7138) );
  NOR2_X1 U8927 ( .A1(n7137), .A2(n7138), .ZN(n7222) );
  AOI211_X1 U8928 ( .C1(n7138), .C2(n7137), .A(n8529), .B(n7222), .ZN(n7139)
         );
  AOI211_X1 U8929 ( .C1(n9867), .C2(n7141), .A(n7140), .B(n7139), .ZN(n7142)
         );
  INV_X1 U8930 ( .A(n7142), .ZN(P2_U3187) );
  INV_X1 U8931 ( .A(n7143), .ZN(n7152) );
  OAI222_X1 U8932 ( .A1(P2_U3151), .A2(n8324), .B1(n8858), .B2(n7152), .C1(
        n7144), .C2(n8860), .ZN(P2_U3275) );
  XNOR2_X1 U8933 ( .A(n7146), .B(n7145), .ZN(n7147) );
  NAND2_X1 U8934 ( .A1(n7147), .A2(n4514), .ZN(n7151) );
  OAI22_X1 U8935 ( .A1(n8160), .A2(n7436), .B1(n9929), .B2(n8178), .ZN(n7148)
         );
  AOI211_X1 U8936 ( .C1(n8157), .C2(n8202), .A(n7149), .B(n7148), .ZN(n7150)
         );
  OAI211_X1 U8937 ( .C1(n8149), .C2(n7173), .A(n7151), .B(n7150), .ZN(P2_U3167) );
  OAI222_X1 U8938 ( .A1(n9521), .A2(n7153), .B1(n7801), .B2(P1_U3086), .C1(
        n9525), .C2(n7152), .ZN(P1_U3335) );
  OAI211_X1 U8939 ( .C1(n7156), .C2(n7155), .A(n7154), .B(n4514), .ZN(n7163)
         );
  NAND2_X1 U8940 ( .A1(n8157), .A2(n9879), .ZN(n7161) );
  NAND2_X1 U8941 ( .A1(n8162), .A2(n7157), .ZN(n7160) );
  NAND2_X1 U8942 ( .A1(n8170), .A2(n8406), .ZN(n7159) );
  INV_X1 U8943 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7158) );
  OR2_X1 U8944 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7158), .ZN(n8423) );
  AND4_X1 U8945 ( .A1(n7161), .A2(n7160), .A3(n7159), .A4(n8423), .ZN(n7162)
         );
  OAI211_X1 U8946 ( .C1(n7291), .C2(n8149), .A(n7163), .B(n7162), .ZN(P2_U3179) );
  INV_X1 U8947 ( .A(n7166), .ZN(n8346) );
  XNOR2_X1 U8948 ( .A(n7164), .B(n8346), .ZN(n7171) );
  OAI21_X1 U8949 ( .B1(n7167), .B2(n7166), .A(n7165), .ZN(n9932) );
  INV_X1 U8950 ( .A(n7992), .ZN(n9903) );
  OAI22_X1 U8951 ( .A1(n7168), .A2(n9891), .B1(n7436), .B2(n9893), .ZN(n7169)
         );
  AOI21_X1 U8952 ( .B1(n9932), .B2(n9903), .A(n7169), .ZN(n7170) );
  OAI21_X1 U8953 ( .B1(n9899), .B2(n7171), .A(n7170), .ZN(n9930) );
  INV_X1 U8954 ( .A(n9930), .ZN(n7177) );
  NAND2_X1 U8955 ( .A1(n8710), .A2(n7172), .ZN(n8005) );
  INV_X1 U8956 ( .A(n8005), .ZN(n9907) );
  NOR2_X1 U8957 ( .A1(n8710), .A2(n5915), .ZN(n7175) );
  INV_X1 U8958 ( .A(n4350), .ZN(n8542) );
  OAI22_X1 U8959 ( .A1(n8542), .A2(n9929), .B1(n8706), .B2(n7173), .ZN(n7174)
         );
  AOI211_X1 U8960 ( .C1(n9932), .C2(n9907), .A(n7175), .B(n7174), .ZN(n7176)
         );
  OAI21_X1 U8961 ( .B1(n7177), .B2(n9910), .A(n7176), .ZN(P2_U3228) );
  INV_X1 U8962 ( .A(n7178), .ZN(n7181) );
  OAI222_X1 U8963 ( .A1(n9525), .A2(n7181), .B1(n7756), .B2(P1_U3086), .C1(
        n7179), .C2(n9521), .ZN(P1_U3334) );
  OAI222_X1 U8964 ( .A1(n8860), .A2(n7182), .B1(n8858), .B2(n7181), .C1(n7180), 
        .C2(P2_U3151), .ZN(P2_U3274) );
  OR2_X1 U8965 ( .A1(n9658), .A2(n9037), .ZN(n7184) );
  NAND2_X1 U8966 ( .A1(n9601), .A2(n9654), .ZN(n7675) );
  OR2_X1 U8967 ( .A1(n7217), .A2(n9673), .ZN(n7679) );
  NAND2_X1 U8968 ( .A1(n7217), .A2(n9673), .ZN(n7772) );
  XNOR2_X1 U8969 ( .A(n7200), .B(n7199), .ZN(n7211) );
  INV_X1 U8970 ( .A(n7678), .ZN(n7187) );
  NOR2_X1 U8971 ( .A1(n7199), .A2(n7187), .ZN(n7188) );
  INV_X1 U8972 ( .A(n7198), .ZN(n7190) );
  AOI21_X1 U8973 ( .B1(n9593), .B2(n7678), .A(n7620), .ZN(n7189) );
  NOR2_X1 U8974 ( .A1(n7190), .A2(n7189), .ZN(n7221) );
  AOI22_X1 U8975 ( .A1(n9036), .A2(n9647), .B1(n9441), .B2(n9034), .ZN(n7191)
         );
  OAI211_X1 U8976 ( .C1(n9602), .C2(n7364), .A(n7204), .B(n9603), .ZN(n7214)
         );
  OAI211_X1 U8977 ( .C1(n7221), .C2(n9680), .A(n7191), .B(n7214), .ZN(n7192)
         );
  AOI21_X1 U8978 ( .B1(n7211), .B2(n9682), .A(n7192), .ZN(n7197) );
  AOI22_X1 U8979 ( .A1(n7217), .A2(n7193), .B1(n9694), .B2(
        P1_REG1_REG_12__SCAN_IN), .ZN(n7194) );
  OAI21_X1 U8980 ( .B1(n7197), .B2(n9694), .A(n7194), .ZN(P1_U3534) );
  OAI22_X1 U8981 ( .A1(n7364), .A2(n9515), .B1(n9685), .B2(n5437), .ZN(n7195)
         );
  INV_X1 U8982 ( .A(n7195), .ZN(n7196) );
  OAI21_X1 U8983 ( .B1(n7197), .B2(n9684), .A(n7196), .ZN(P1_U3489) );
  NAND2_X1 U8984 ( .A1(n7198), .A2(n7772), .ZN(n7326) );
  AND2_X1 U8985 ( .A1(n7381), .A2(n9034), .ZN(n7684) );
  NAND2_X1 U8986 ( .A1(n9676), .A2(n8867), .ZN(n7773) );
  XNOR2_X1 U8987 ( .A(n7326), .B(n7329), .ZN(n9679) );
  OR2_X1 U8988 ( .A1(n7217), .A2(n9035), .ZN(n7201) );
  XNOR2_X1 U8989 ( .A(n7330), .B(n7329), .ZN(n9683) );
  NAND2_X1 U8990 ( .A1(n9683), .A2(n9618), .ZN(n7210) );
  INV_X1 U8991 ( .A(n7336), .ZN(n7203) );
  AOI211_X1 U8992 ( .C1(n9676), .C2(n7204), .A(n9348), .B(n7203), .ZN(n9674)
         );
  NOR2_X1 U8993 ( .A1(n7381), .A2(n9614), .ZN(n7208) );
  NAND2_X1 U8994 ( .A1(n9296), .A2(n9035), .ZN(n7206) );
  AOI22_X1 U8995 ( .A1(n4352), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7378), .B2(
        n9610), .ZN(n7205) );
  OAI211_X1 U8996 ( .C1(n9671), .C2(n9300), .A(n7206), .B(n7205), .ZN(n7207)
         );
  AOI211_X1 U8997 ( .C1(n9674), .C2(n9608), .A(n7208), .B(n7207), .ZN(n7209)
         );
  OAI211_X1 U8998 ( .C1(n9679), .C2(n7220), .A(n7210), .B(n7209), .ZN(P1_U3280) );
  NAND2_X1 U8999 ( .A1(n7211), .A2(n9618), .ZN(n7219) );
  NAND2_X1 U9000 ( .A1(n9296), .A2(n9036), .ZN(n7213) );
  AOI22_X1 U9001 ( .A1(n4352), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7361), .B2(
        n9610), .ZN(n7212) );
  OAI211_X1 U9002 ( .C1(n8867), .C2(n9300), .A(n7213), .B(n7212), .ZN(n7216)
         );
  NOR2_X1 U9003 ( .A1(n7214), .A2(n9305), .ZN(n7215) );
  AOI211_X1 U9004 ( .C1(n9600), .C2(n7217), .A(n7216), .B(n7215), .ZN(n7218)
         );
  OAI211_X1 U9005 ( .C1(n7221), .C2(n7220), .A(n7219), .B(n7218), .ZN(P1_U3281) );
  MUX2_X1 U9006 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n8856), .Z(n7224) );
  XOR2_X1 U9007 ( .A(n8420), .B(n7224), .Z(n8412) );
  NAND2_X1 U9008 ( .A1(n8413), .A2(n8412), .ZN(n8411) );
  OAI21_X1 U9009 ( .B1(n7224), .B2(n8420), .A(n8411), .ZN(n8488) );
  MUX2_X1 U9010 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n8856), .Z(n8484) );
  INV_X1 U9011 ( .A(n8454), .ZN(n8486) );
  XNOR2_X1 U9012 ( .A(n8484), .B(n8486), .ZN(n8487) );
  XNOR2_X1 U9013 ( .A(n8488), .B(n8487), .ZN(n7243) );
  NAND2_X1 U9014 ( .A1(n9857), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7241) );
  MUX2_X1 U9015 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n5929), .S(n8420), .Z(n8415)
         );
  NAND2_X1 U9016 ( .A1(n8420), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n7225) );
  NAND2_X1 U9017 ( .A1(n7226), .A2(n8454), .ZN(n8434) );
  AND2_X1 U9018 ( .A1(n7227), .A2(n5944), .ZN(n7228) );
  OAI21_X1 U9019 ( .B1(n9704), .B2(n7228), .A(n9798), .ZN(n7240) );
  AOI21_X1 U9020 ( .B1(n9858), .B2(n8486), .A(n7229), .ZN(n7239) );
  NAND2_X1 U9021 ( .A1(n7230), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7234) );
  NAND2_X1 U9022 ( .A1(n7232), .A2(n7231), .ZN(n7233) );
  NAND2_X1 U9023 ( .A1(n7234), .A2(n7233), .ZN(n8427) );
  MUX2_X1 U9024 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7235), .S(n8420), .Z(n8428)
         );
  NAND2_X1 U9025 ( .A1(n8427), .A2(n8428), .ZN(n8426) );
  NAND2_X1 U9026 ( .A1(n8420), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n7236) );
  XNOR2_X1 U9027 ( .A(n8453), .B(n8486), .ZN(n8455) );
  XNOR2_X1 U9028 ( .A(n8455), .B(P2_REG1_REG_7__SCAN_IN), .ZN(n7237) );
  NAND2_X1 U9029 ( .A1(n7237), .A2(n9867), .ZN(n7238) );
  NAND4_X1 U9030 ( .A1(n7241), .A2(n7240), .A3(n7239), .A4(n7238), .ZN(n7242)
         );
  AOI21_X1 U9031 ( .B1(n7243), .B2(n9866), .A(n7242), .ZN(n7244) );
  INV_X1 U9032 ( .A(n7244), .ZN(P2_U3189) );
  AOI21_X1 U9033 ( .B1(n7248), .B2(n7245), .A(n7247), .ZN(n7256) );
  NAND2_X1 U9034 ( .A1(P1_U3086), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n9539) );
  INV_X1 U9035 ( .A(n9539), .ZN(n7249) );
  AOI21_X1 U9036 ( .B1(n8889), .B2(n9038), .A(n7249), .ZN(n7253) );
  NAND2_X1 U9037 ( .A1(n9022), .A2(n7250), .ZN(n7252) );
  NAND2_X1 U9038 ( .A1(n9018), .A2(n9036), .ZN(n7251) );
  NAND3_X1 U9039 ( .A1(n7253), .A2(n7252), .A3(n7251), .ZN(n7254) );
  AOI21_X1 U9040 ( .B1(n9658), .B2(n8958), .A(n7254), .ZN(n7255) );
  OAI21_X1 U9041 ( .B1(n7256), .B2(n8960), .A(n7255), .ZN(P1_U3217) );
  XNOR2_X1 U9042 ( .A(n7833), .B(n7827), .ZN(n7828) );
  NOR2_X1 U9043 ( .A1(n7257), .A2(n7264), .ZN(n7259) );
  NOR2_X1 U9044 ( .A1(n7259), .A2(n7258), .ZN(n7279) );
  INV_X1 U9045 ( .A(n7279), .ZN(n7260) );
  XNOR2_X1 U9046 ( .A(n7287), .B(P1_REG1_REG_16__SCAN_IN), .ZN(n7278) );
  OAI22_X1 U9047 ( .A1(n7260), .A2(n7278), .B1(n7287), .B2(
        P1_REG1_REG_16__SCAN_IN), .ZN(n7829) );
  XOR2_X1 U9048 ( .A(n7828), .B(n7829), .Z(n7277) );
  INV_X1 U9049 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n7261) );
  NAND2_X1 U9050 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n8945) );
  OAI21_X1 U9051 ( .B1(n9590), .B2(n7261), .A(n8945), .ZN(n7262) );
  AOI21_X1 U9052 ( .B1(n9564), .B2(n7833), .A(n7262), .ZN(n7276) );
  INV_X1 U9053 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n7263) );
  XNOR2_X1 U9054 ( .A(n7833), .B(n7263), .ZN(n7273) );
  NOR2_X1 U9055 ( .A1(n7265), .A2(n7264), .ZN(n7267) );
  NOR2_X1 U9056 ( .A1(n7267), .A2(n7266), .ZN(n7283) );
  INV_X1 U9057 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7268) );
  OR2_X1 U9058 ( .A1(n7287), .A2(n7268), .ZN(n7270) );
  NAND2_X1 U9059 ( .A1(n7287), .A2(n7268), .ZN(n7269) );
  AND2_X1 U9060 ( .A1(n7270), .A2(n7269), .ZN(n7284) );
  OR2_X1 U9061 ( .A1(n7283), .A2(n7284), .ZN(n7281) );
  NAND2_X1 U9062 ( .A1(n7287), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n7271) );
  NAND2_X1 U9063 ( .A1(n7272), .A2(n7273), .ZN(n7835) );
  OAI21_X1 U9064 ( .B1(n7273), .B2(n7272), .A(n7835), .ZN(n7274) );
  NAND2_X1 U9065 ( .A1(n7274), .A2(n9580), .ZN(n7275) );
  OAI211_X1 U9066 ( .C1(n7277), .C2(n9528), .A(n7276), .B(n7275), .ZN(P1_U3260) );
  XNOR2_X1 U9067 ( .A(n7279), .B(n7278), .ZN(n7289) );
  INV_X1 U9068 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7280) );
  NAND2_X1 U9069 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8932) );
  OAI21_X1 U9070 ( .B1(n9590), .B2(n7280), .A(n8932), .ZN(n7286) );
  INV_X1 U9071 ( .A(n9580), .ZN(n9532) );
  INV_X1 U9072 ( .A(n7281), .ZN(n7282) );
  AOI211_X1 U9073 ( .C1(n7284), .C2(n7283), .A(n9532), .B(n7282), .ZN(n7285)
         );
  AOI211_X1 U9074 ( .C1(n9564), .C2(n7287), .A(n7286), .B(n7285), .ZN(n7288)
         );
  OAI21_X1 U9075 ( .B1(n7289), .B2(n9528), .A(n7288), .ZN(P1_U3259) );
  XNOR2_X1 U9076 ( .A(n7290), .B(n8348), .ZN(n9937) );
  OAI22_X1 U9077 ( .A1(n8542), .A2(n9934), .B1(n7291), .B2(n8706), .ZN(n7300)
         );
  NAND2_X1 U9078 ( .A1(n7293), .A2(n7292), .ZN(n7294) );
  NAND2_X1 U9079 ( .A1(n7294), .A2(n8348), .ZN(n7295) );
  NAND3_X1 U9080 ( .A1(n7296), .A2(n9883), .A3(n7295), .ZN(n7298) );
  AOI22_X1 U9081 ( .A1(n8406), .A2(n9878), .B1(n9880), .B2(n9879), .ZN(n7297)
         );
  NAND2_X1 U9082 ( .A1(n7298), .A2(n7297), .ZN(n9935) );
  MUX2_X1 U9083 ( .A(n9935), .B(P2_REG2_REG_6__SCAN_IN), .S(n9910), .Z(n7299)
         );
  AOI211_X1 U9084 ( .C1(n9888), .C2(n9937), .A(n7300), .B(n7299), .ZN(n7301)
         );
  INV_X1 U9085 ( .A(n7301), .ZN(P2_U3227) );
  INV_X1 U9086 ( .A(n7302), .ZN(n7304) );
  NOR3_X1 U9087 ( .A1(n7247), .A2(n7304), .A3(n7303), .ZN(n7306) );
  INV_X1 U9088 ( .A(n7305), .ZN(n7354) );
  OAI21_X1 U9089 ( .B1(n7306), .B2(n7354), .A(n9016), .ZN(n7311) );
  NOR2_X1 U9090 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7307), .ZN(n9586) );
  AOI21_X1 U9091 ( .B1(n8889), .B2(n9037), .A(n9586), .ZN(n7308) );
  OAI21_X1 U9092 ( .B1(n9673), .B2(n9008), .A(n7308), .ZN(n7309) );
  AOI21_X1 U9093 ( .B1(n9599), .B2(n9022), .A(n7309), .ZN(n7310) );
  OAI211_X1 U9094 ( .C1(n4681), .C2(n9026), .A(n7311), .B(n7310), .ZN(P1_U3236) );
  INV_X1 U9095 ( .A(n7312), .ZN(n7314) );
  OAI222_X1 U9096 ( .A1(n9521), .A2(n7313), .B1(n9525), .B2(n7314), .C1(
        P1_U3086), .C2(n7804), .ZN(P1_U3333) );
  OAI222_X1 U9097 ( .A1(n8860), .A2(n7315), .B1(n8858), .B2(n7314), .C1(
        P2_U3151), .C2(n8182), .ZN(P2_U3273) );
  XNOR2_X1 U9098 ( .A(n7962), .B(n7323), .ZN(n7382) );
  XNOR2_X1 U9099 ( .A(n7382), .B(n7435), .ZN(n7319) );
  XNOR2_X1 U9100 ( .A(n4445), .B(n7319), .ZN(n7325) );
  NOR2_X1 U9101 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10095), .ZN(n9710) );
  AOI21_X1 U9102 ( .B1(n8157), .B2(n8406), .A(n9710), .ZN(n7321) );
  NAND2_X1 U9103 ( .A1(n8170), .A2(n8404), .ZN(n7320) );
  OAI211_X1 U9104 ( .C1(n8149), .C2(n7411), .A(n7321), .B(n7320), .ZN(n7322)
         );
  AOI21_X1 U9105 ( .B1(n7323), .B2(n8162), .A(n7322), .ZN(n7324) );
  OAI21_X1 U9106 ( .B1(n7325), .B2(n8164), .A(n7324), .ZN(P2_U3161) );
  NAND2_X1 U9107 ( .A1(n7326), .A2(n7621), .ZN(n7327) );
  NAND2_X1 U9108 ( .A1(n7327), .A2(n7773), .ZN(n7452) );
  OR2_X1 U9109 ( .A1(n7444), .A2(n9671), .ZN(n7777) );
  NAND2_X1 U9110 ( .A1(n7444), .A2(n9671), .ZN(n7693) );
  NAND2_X1 U9111 ( .A1(n7777), .A2(n7693), .ZN(n7683) );
  INV_X1 U9112 ( .A(n7683), .ZN(n7451) );
  XNOR2_X1 U9113 ( .A(n7452), .B(n7451), .ZN(n7328) );
  AND2_X1 U9114 ( .A1(n7328), .A2(n9447), .ZN(n7346) );
  INV_X1 U9115 ( .A(n7346), .ZN(n7342) );
  NAND2_X1 U9116 ( .A1(n7381), .A2(n8867), .ZN(n7331) );
  XNOR2_X1 U9117 ( .A(n7447), .B(n7683), .ZN(n7347) );
  NAND2_X1 U9118 ( .A1(n7347), .A2(n9618), .ZN(n7341) );
  NAND2_X1 U9119 ( .A1(n9296), .A2(n9034), .ZN(n7334) );
  AOI22_X1 U9120 ( .A1(n4352), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8869), .B2(
        n9610), .ZN(n7333) );
  OAI211_X1 U9121 ( .C1(n8934), .C2(n9300), .A(n7334), .B(n7333), .ZN(n7339)
         );
  NAND2_X1 U9122 ( .A1(n7336), .A2(n7444), .ZN(n7335) );
  NAND2_X1 U9123 ( .A1(n7335), .A2(n9603), .ZN(n7337) );
  OR2_X1 U9124 ( .A1(n7337), .A2(n7448), .ZN(n7344) );
  NOR2_X1 U9125 ( .A1(n7344), .A2(n9305), .ZN(n7338) );
  AOI211_X1 U9126 ( .C1(n9600), .C2(n7444), .A(n7339), .B(n7338), .ZN(n7340)
         );
  OAI211_X1 U9127 ( .C1(n4352), .C2(n7342), .A(n7341), .B(n7340), .ZN(P1_U3279) );
  INV_X1 U9128 ( .A(n7444), .ZN(n8872) );
  AOI22_X1 U9129 ( .A1(n9032), .A2(n9441), .B1(n9647), .B2(n9034), .ZN(n7343)
         );
  OAI211_X1 U9130 ( .C1(n8872), .C2(n9664), .A(n7344), .B(n7343), .ZN(n7345)
         );
  AOI211_X1 U9131 ( .C1(n7347), .C2(n9682), .A(n7346), .B(n7345), .ZN(n7350)
         );
  NAND2_X1 U9132 ( .A1(n9694), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7348) );
  OAI21_X1 U9133 ( .B1(n7350), .B2(n9694), .A(n7348), .ZN(P1_U3536) );
  NAND2_X1 U9134 ( .A1(n9684), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7349) );
  OAI21_X1 U9135 ( .B1(n7350), .B2(n9684), .A(n7349), .ZN(P1_U3495) );
  INV_X1 U9136 ( .A(n7351), .ZN(n7353) );
  NOR3_X1 U9137 ( .A1(n7354), .A2(n7353), .A3(n7352), .ZN(n7357) );
  INV_X1 U9138 ( .A(n7355), .ZN(n7356) );
  OAI21_X1 U9139 ( .B1(n7357), .B2(n7356), .A(n9016), .ZN(n7363) );
  NAND2_X1 U9140 ( .A1(n9018), .A2(n9034), .ZN(n7359) );
  OAI211_X1 U9141 ( .C1(n9654), .C2(n8988), .A(n7359), .B(n7358), .ZN(n7360)
         );
  AOI21_X1 U9142 ( .B1(n7361), .B2(n9022), .A(n7360), .ZN(n7362) );
  OAI211_X1 U9143 ( .C1(n7364), .C2(n9026), .A(n7363), .B(n7362), .ZN(P1_U3224) );
  NAND2_X1 U9144 ( .A1(n7368), .A2(n7820), .ZN(n7365) );
  OAI211_X1 U9145 ( .C1(n7366), .C2(n7561), .A(n7365), .B(n8394), .ZN(P2_U3272) );
  NAND2_X1 U9146 ( .A1(n7368), .A2(n7367), .ZN(n7369) );
  OAI211_X1 U9147 ( .C1(n7370), .C2(n9521), .A(n7369), .B(n7819), .ZN(P1_U3332) );
  OAI21_X1 U9148 ( .B1(n7373), .B2(n7372), .A(n7371), .ZN(n7374) );
  NAND2_X1 U9149 ( .A1(n7374), .A2(n9016), .ZN(n7380) );
  NAND2_X1 U9150 ( .A1(n9018), .A2(n9033), .ZN(n7376) );
  OAI211_X1 U9151 ( .C1(n9673), .C2(n8988), .A(n7376), .B(n7375), .ZN(n7377)
         );
  AOI21_X1 U9152 ( .B1(n7378), .B2(n9022), .A(n7377), .ZN(n7379) );
  OAI211_X1 U9153 ( .C1(n7381), .C2(n9026), .A(n7380), .B(n7379), .ZN(P1_U3234) );
  INV_X1 U9154 ( .A(n7382), .ZN(n7383) );
  XNOR2_X1 U9155 ( .A(n9950), .B(n6370), .ZN(n7921) );
  XNOR2_X1 U9156 ( .A(n7921), .B(n7509), .ZN(n7922) );
  XNOR2_X1 U9157 ( .A(n7923), .B(n7922), .ZN(n7388) );
  INV_X1 U9158 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n10222) );
  NOR2_X1 U9159 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10222), .ZN(n9726) );
  AOI21_X1 U9160 ( .B1(n8157), .B2(n8405), .A(n9726), .ZN(n7385) );
  NAND2_X1 U9161 ( .A1(n8170), .A2(n8403), .ZN(n7384) );
  OAI211_X1 U9162 ( .C1(n8149), .C2(n7403), .A(n7385), .B(n7384), .ZN(n7386)
         );
  AOI21_X1 U9163 ( .B1(n7405), .B2(n8162), .A(n7386), .ZN(n7387) );
  OAI21_X1 U9164 ( .B1(n7388), .B2(n8164), .A(n7387), .ZN(P2_U3171) );
  NAND2_X1 U9165 ( .A1(n7409), .A2(n7389), .ZN(n7391) );
  AND2_X1 U9166 ( .A1(n7391), .A2(n7390), .ZN(n7502) );
  AND2_X1 U9167 ( .A1(n7409), .A2(n7392), .ZN(n7394) );
  NOR2_X1 U9168 ( .A1(n7394), .A2(n7393), .ZN(n7395) );
  NAND2_X1 U9169 ( .A1(n7395), .A2(n8351), .ZN(n7396) );
  NAND2_X1 U9170 ( .A1(n7502), .A2(n7396), .ZN(n9951) );
  NAND2_X1 U9171 ( .A1(n7397), .A2(n8350), .ZN(n7412) );
  AND2_X1 U9172 ( .A1(n7412), .A2(n7398), .ZN(n7399) );
  NAND2_X1 U9173 ( .A1(n7399), .A2(n8351), .ZN(n7507) );
  OAI21_X1 U9174 ( .B1(n7399), .B2(n8351), .A(n7507), .ZN(n7401) );
  OAI22_X1 U9175 ( .A1(n8059), .A2(n9893), .B1(n7435), .B2(n9891), .ZN(n7400)
         );
  AOI21_X1 U9176 ( .B1(n7401), .B2(n9883), .A(n7400), .ZN(n7402) );
  OAI21_X1 U9177 ( .B1(n7992), .B2(n9951), .A(n7402), .ZN(n9953) );
  NAND2_X1 U9178 ( .A1(n9953), .A2(n8710), .ZN(n7407) );
  OAI22_X1 U9179 ( .A1(n8710), .A2(n5973), .B1(n7403), .B2(n8706), .ZN(n7404)
         );
  AOI21_X1 U9180 ( .B1(n4350), .B2(n7405), .A(n7404), .ZN(n7406) );
  OAI211_X1 U9181 ( .C1(n9951), .C2(n8005), .A(n7407), .B(n7406), .ZN(P2_U3224) );
  AND2_X1 U9182 ( .A1(n7409), .A2(n7408), .ZN(n7410) );
  XNOR2_X1 U9183 ( .A(n7410), .B(n8350), .ZN(n9947) );
  OAI22_X1 U9184 ( .A1(n8542), .A2(n9944), .B1(n7411), .B2(n8706), .ZN(n7416)
         );
  OAI211_X1 U9185 ( .C1(n7397), .C2(n8350), .A(n7412), .B(n9883), .ZN(n7414)
         );
  AOI22_X1 U9186 ( .A1(n8406), .A2(n9880), .B1(n9878), .B2(n8404), .ZN(n7413)
         );
  NAND2_X1 U9187 ( .A1(n7414), .A2(n7413), .ZN(n9945) );
  MUX2_X1 U9188 ( .A(n9945), .B(P2_REG2_REG_8__SCAN_IN), .S(n9910), .Z(n7415)
         );
  AOI211_X1 U9189 ( .C1(n9888), .C2(n9947), .A(n7416), .B(n7415), .ZN(n7417)
         );
  INV_X1 U9190 ( .A(n7417), .ZN(P2_U3225) );
  AND2_X1 U9191 ( .A1(n7419), .A2(n7418), .ZN(n7420) );
  XNOR2_X1 U9192 ( .A(n7420), .B(n7926), .ZN(n9963) );
  XNOR2_X1 U9193 ( .A(n7421), .B(n7926), .ZN(n7422) );
  OAI222_X1 U9194 ( .A1(n9893), .A2(n8117), .B1(n9891), .B2(n8059), .C1(n7422), 
        .C2(n9899), .ZN(n9964) );
  NAND2_X1 U9195 ( .A1(n9964), .A2(n8710), .ZN(n7426) );
  OAI22_X1 U9196 ( .A1(n8710), .A2(n7423), .B1(n8139), .B2(n8706), .ZN(n7424)
         );
  AOI21_X1 U9197 ( .B1(n4350), .B2(n9966), .A(n7424), .ZN(n7425) );
  OAI211_X1 U9198 ( .C1(n8699), .C2(n9963), .A(n7426), .B(n7425), .ZN(P2_U3222) );
  NAND2_X1 U9199 ( .A1(n7427), .A2(n8214), .ZN(n7428) );
  NAND2_X1 U9200 ( .A1(n7428), .A2(n8217), .ZN(n7430) );
  OR2_X1 U9201 ( .A1(n7428), .A2(n8217), .ZN(n7429) );
  NAND2_X1 U9202 ( .A1(n7430), .A2(n7429), .ZN(n9940) );
  INV_X1 U9203 ( .A(n9940), .ZN(n7442) );
  OAI22_X1 U9204 ( .A1(n8542), .A2(n9939), .B1(n7431), .B2(n8706), .ZN(n7441)
         );
  OAI21_X1 U9205 ( .B1(n7433), .B2(n8352), .A(n7432), .ZN(n7434) );
  NAND2_X1 U9206 ( .A1(n7434), .A2(n9883), .ZN(n7439) );
  OAI22_X1 U9207 ( .A1(n7436), .A2(n9891), .B1(n7435), .B2(n9893), .ZN(n7437)
         );
  INV_X1 U9208 ( .A(n7437), .ZN(n7438) );
  OAI211_X1 U9209 ( .C1(n9940), .C2(n7992), .A(n7439), .B(n7438), .ZN(n9942)
         );
  MUX2_X1 U9210 ( .A(n9942), .B(P2_REG2_REG_7__SCAN_IN), .S(n9910), .Z(n7440)
         );
  AOI211_X1 U9211 ( .C1(n7442), .C2(n9907), .A(n7441), .B(n7440), .ZN(n7443)
         );
  INV_X1 U9212 ( .A(n7443), .ZN(P2_U3226) );
  NOR2_X1 U9213 ( .A1(n7444), .A2(n9033), .ZN(n7446) );
  NAND2_X1 U9214 ( .A1(n7444), .A2(n9033), .ZN(n7445) );
  NAND2_X1 U9215 ( .A1(n9474), .A2(n8934), .ZN(n7692) );
  XNOR2_X1 U9216 ( .A(n7469), .B(n7453), .ZN(n9477) );
  INV_X1 U9217 ( .A(n7448), .ZN(n7449) );
  AOI211_X1 U9218 ( .C1(n9474), .C2(n7449), .A(n9348), .B(n7463), .ZN(n9473)
         );
  AOI22_X1 U9219 ( .A1(n4352), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n9023), .B2(
        n9610), .ZN(n7450) );
  OAI21_X1 U9220 ( .B1(n9027), .B2(n9614), .A(n7450), .ZN(n7458) );
  AOI21_X1 U9221 ( .B1(n7454), .B2(n7453), .A(n9680), .ZN(n7456) );
  OAI22_X1 U9222 ( .A1(n9356), .A2(n9670), .B1(n9671), .B2(n9672), .ZN(n7455)
         );
  AOI21_X1 U9223 ( .B1(n7456), .B2(n7460), .A(n7455), .ZN(n9476) );
  NOR2_X1 U9224 ( .A1(n9476), .A2(n4352), .ZN(n7457) );
  AOI211_X1 U9225 ( .C1(n9473), .C2(n9608), .A(n7458), .B(n7457), .ZN(n7459)
         );
  OAI21_X1 U9226 ( .B1(n9364), .B2(n9477), .A(n7459), .ZN(P1_U3278) );
  NAND2_X1 U9227 ( .A1(n7461), .A2(n7625), .ZN(n7574) );
  OAI21_X1 U9228 ( .B1(n7625), .B2(n7461), .A(n7574), .ZN(n7462) );
  AOI222_X1 U9229 ( .A1(n9447), .A2(n7462), .B1(n9030), .B2(n9441), .C1(n9032), 
        .C2(n9647), .ZN(n9471) );
  INV_X1 U9230 ( .A(n7463), .ZN(n7465) );
  NAND2_X1 U9231 ( .A1(n8935), .A2(n7463), .ZN(n9349) );
  INV_X1 U9232 ( .A(n9349), .ZN(n7464) );
  AOI21_X1 U9233 ( .B1(n9468), .B2(n7465), .A(n7464), .ZN(n9469) );
  AOI22_X1 U9234 ( .A1(n4352), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n8938), .B2(
        n9610), .ZN(n7466) );
  OAI21_X1 U9235 ( .B1(n8935), .B2(n9614), .A(n7466), .ZN(n7467) );
  AOI21_X1 U9236 ( .B1(n9469), .B2(n9161), .A(n7467), .ZN(n7473) );
  AND2_X1 U9237 ( .A1(n9474), .A2(n9032), .ZN(n7468) );
  OR2_X1 U9238 ( .A1(n9474), .A2(n9032), .ZN(n7470) );
  OR2_X2 U9239 ( .A1(n7471), .A2(n7625), .ZN(n7850) );
  NAND2_X1 U9240 ( .A1(n7471), .A2(n7625), .ZN(n9467) );
  NAND3_X1 U9241 ( .A1(n7850), .A2(n9467), .A3(n9618), .ZN(n7472) );
  OAI211_X1 U9242 ( .C1(n9471), .C2(n4352), .A(n7473), .B(n7472), .ZN(P1_U3277) );
  INV_X1 U9243 ( .A(n7474), .ZN(n7493) );
  OAI222_X1 U9244 ( .A1(n7476), .A2(P2_U3151), .B1(n8858), .B2(n7493), .C1(
        n7475), .C2(n8860), .ZN(P2_U3271) );
  NAND2_X1 U9245 ( .A1(n7477), .A2(n8355), .ZN(n7478) );
  NAND3_X1 U9246 ( .A1(n7479), .A2(n9883), .A3(n7478), .ZN(n7481) );
  AOI22_X1 U9247 ( .A1(n9880), .A2(n8402), .B1(n8704), .B2(n9878), .ZN(n7480)
         );
  AND2_X1 U9248 ( .A1(n7481), .A2(n7480), .ZN(n7497) );
  MUX2_X1 U9249 ( .A(n7497), .B(n7482), .S(n9970), .Z(n7488) );
  INV_X1 U9250 ( .A(n7483), .ZN(n7484) );
  AOI21_X1 U9251 ( .B1(n7486), .B2(n7485), .A(n7484), .ZN(n7496) );
  AOI22_X1 U9252 ( .A1(n7496), .A2(n8851), .B1(n8850), .B2(n8068), .ZN(n7487)
         );
  NAND2_X1 U9253 ( .A1(n7488), .A2(n7487), .ZN(P2_U3426) );
  INV_X1 U9254 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7489) );
  MUX2_X1 U9255 ( .A(n7489), .B(n7497), .S(n9986), .Z(n7491) );
  AOI22_X1 U9256 ( .A1(n7496), .A2(n8762), .B1(n8761), .B2(n8068), .ZN(n7490)
         );
  NAND2_X1 U9257 ( .A1(n7491), .A2(n7490), .ZN(P2_U3471) );
  INV_X1 U9258 ( .A(n7492), .ZN(n7494) );
  OAI222_X1 U9259 ( .A1(n9521), .A2(n7495), .B1(n7494), .B2(P1_U3086), .C1(
        n9525), .C2(n7493), .ZN(P1_U3331) );
  INV_X1 U9260 ( .A(n7496), .ZN(n7501) );
  MUX2_X1 U9261 ( .A(n7497), .B(n8440), .S(n9910), .Z(n7500) );
  INV_X1 U9262 ( .A(n8066), .ZN(n7498) );
  AOI22_X1 U9263 ( .A1(n8068), .A2(n4350), .B1(n9905), .B2(n7498), .ZN(n7499)
         );
  OAI211_X1 U9264 ( .C1(n7501), .C2(n8699), .A(n7500), .B(n7499), .ZN(P2_U3221) );
  NAND2_X1 U9265 ( .A1(n7502), .A2(n8221), .ZN(n7505) );
  XNOR2_X1 U9266 ( .A(n7505), .B(n8354), .ZN(n9958) );
  NAND2_X1 U9267 ( .A1(n7507), .A2(n7506), .ZN(n7508) );
  XOR2_X1 U9268 ( .A(n8354), .B(n7508), .Z(n7511) );
  OAI22_X1 U9269 ( .A1(n7509), .A2(n9891), .B1(n8063), .B2(n9893), .ZN(n7510)
         );
  AOI21_X1 U9270 ( .B1(n7511), .B2(n9883), .A(n7510), .ZN(n7512) );
  OAI21_X1 U9271 ( .B1(n7992), .B2(n9958), .A(n7512), .ZN(n9960) );
  NAND2_X1 U9272 ( .A1(n9960), .A2(n8710), .ZN(n7515) );
  OAI22_X1 U9273 ( .A1(n8710), .A2(n8437), .B1(n8040), .B2(n8706), .ZN(n7513)
         );
  AOI21_X1 U9274 ( .B1(n4350), .B2(n7927), .A(n7513), .ZN(n7514) );
  OAI211_X1 U9275 ( .C1(n9958), .C2(n8005), .A(n7515), .B(n7514), .ZN(P2_U3223) );
  INV_X1 U9276 ( .A(n7516), .ZN(n7519) );
  OAI222_X1 U9277 ( .A1(n7518), .A2(P2_U3151), .B1(n8858), .B2(n7519), .C1(
        n7517), .C2(n8860), .ZN(P2_U3270) );
  OAI222_X1 U9278 ( .A1(n9521), .A2(n7521), .B1(n7520), .B2(P1_U3086), .C1(
        n9525), .C2(n7519), .ZN(P1_U3330) );
  INV_X1 U9279 ( .A(n7522), .ZN(n7525) );
  OAI222_X1 U9280 ( .A1(n7524), .A2(P2_U3151), .B1(n8858), .B2(n7525), .C1(
        n7523), .C2(n8860), .ZN(P2_U3269) );
  OAI222_X1 U9281 ( .A1(n9521), .A2(n7527), .B1(n7526), .B2(P1_U3086), .C1(
        n9525), .C2(n7525), .ZN(P1_U3329) );
  INV_X1 U9282 ( .A(n7528), .ZN(n8857) );
  OAI222_X1 U9283 ( .A1(n9525), .A2(n8857), .B1(n7891), .B2(P1_U3086), .C1(
        n7529), .C2(n9521), .ZN(P1_U3328) );
  XOR2_X1 U9284 ( .A(n7530), .B(n8359), .Z(n7531) );
  INV_X1 U9285 ( .A(n8117), .ZN(n8401) );
  AOI222_X1 U9286 ( .A1(n9883), .A2(n7531), .B1(n8692), .B2(n9878), .C1(n8401), 
        .C2(n9880), .ZN(n7540) );
  INV_X1 U9287 ( .A(n7540), .ZN(n7533) );
  INV_X1 U9288 ( .A(n8249), .ZN(n8122) );
  OAI22_X1 U9289 ( .A1(n8122), .A2(n8708), .B1(n8115), .B2(n8706), .ZN(n7532)
         );
  OAI21_X1 U9290 ( .B1(n7533), .B2(n7532), .A(n8710), .ZN(n7536) );
  XNOR2_X1 U9291 ( .A(n7534), .B(n8359), .ZN(n7542) );
  AOI22_X1 U9292 ( .A1(n7542), .A2(n9888), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n9910), .ZN(n7535) );
  NAND2_X1 U9293 ( .A1(n7536), .A2(n7535), .ZN(P2_U3220) );
  INV_X1 U9294 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7537) );
  MUX2_X1 U9295 ( .A(n7537), .B(n7540), .S(n9968), .Z(n7539) );
  AOI22_X1 U9296 ( .A1(n7542), .A2(n8851), .B1(n8850), .B2(n8249), .ZN(n7538)
         );
  NAND2_X1 U9297 ( .A1(n7539), .A2(n7538), .ZN(P2_U3429) );
  MUX2_X1 U9298 ( .A(n7541), .B(n7540), .S(n9986), .Z(n7544) );
  AOI22_X1 U9299 ( .A1(n7542), .A2(n8762), .B1(n8761), .B2(n8249), .ZN(n7543)
         );
  NAND2_X1 U9300 ( .A1(n7544), .A2(n7543), .ZN(P2_U3472) );
  INV_X1 U9301 ( .A(n7545), .ZN(n7546) );
  MUX2_X1 U9302 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7550), .Z(n7549) );
  XNOR2_X1 U9303 ( .A(n7549), .B(SI_30_), .ZN(n7588) );
  MUX2_X1 U9304 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7550), .Z(n7551) );
  XNOR2_X1 U9305 ( .A(n7551), .B(SI_31_), .ZN(n7552) );
  NOR2_X1 U9306 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_30__SCAN_IN), .ZN(
        n7555) );
  NAND4_X1 U9307 ( .A1(n7555), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .A4(n7554), .ZN(n7556) );
  OAI22_X1 U9308 ( .A1(n7557), .A2(n7556), .B1(n7009), .B2(n9521), .ZN(n7558)
         );
  INV_X1 U9309 ( .A(n7558), .ZN(n7559) );
  OAI21_X1 U9310 ( .B1(n8322), .B2(n9525), .A(n7559), .ZN(P1_U3324) );
  NAND3_X1 U9311 ( .A1(n7560), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n7562) );
  OAI22_X1 U9312 ( .A1(n7563), .A2(n7562), .B1(n6500), .B2(n7561), .ZN(n7564)
         );
  INV_X1 U9313 ( .A(n7564), .ZN(n7565) );
  OAI21_X1 U9314 ( .B1(n8322), .B2(n8858), .A(n7565), .ZN(P2_U3264) );
  OAI222_X1 U9315 ( .A1(n9521), .A2(n7567), .B1(n9525), .B2(n7566), .C1(
        P1_U3086), .C2(n7815), .ZN(P1_U3336) );
  OR2_X1 U9316 ( .A1(n9209), .A2(n9402), .ZN(n7728) );
  NOR2_X1 U9317 ( .A1(n9231), .A2(n9390), .ZN(n7726) );
  INV_X1 U9318 ( .A(n7726), .ZN(n7602) );
  NAND2_X1 U9319 ( .A1(n7728), .A2(n7602), .ZN(n7735) );
  NAND2_X1 U9320 ( .A1(n9507), .A2(n9424), .ZN(n7719) );
  OR2_X1 U9321 ( .A1(n9266), .A2(n9417), .ZN(n7603) );
  NAND2_X1 U9322 ( .A1(n7719), .A2(n7603), .ZN(n7718) );
  NAND2_X1 U9323 ( .A1(n9260), .A2(n9270), .ZN(n7877) );
  NAND2_X1 U9324 ( .A1(n7718), .A2(n7877), .ZN(n7568) );
  OR2_X1 U9325 ( .A1(n9243), .A2(n9258), .ZN(n7880) );
  NAND2_X1 U9326 ( .A1(n7568), .A2(n7880), .ZN(n7569) );
  NAND2_X1 U9327 ( .A1(n9243), .A2(n9258), .ZN(n7723) );
  AND2_X1 U9328 ( .A1(n7569), .A2(n7723), .ZN(n7570) );
  NOR2_X1 U9329 ( .A1(n7735), .A2(n7570), .ZN(n7578) );
  INV_X1 U9330 ( .A(n7578), .ZN(n7573) );
  OR2_X1 U9331 ( .A1(n9287), .A2(n9301), .ZN(n7575) );
  NOR2_X1 U9332 ( .A1(n9303), .A2(n9316), .ZN(n7707) );
  INV_X1 U9333 ( .A(n7707), .ZN(n7571) );
  AND2_X1 U9334 ( .A1(n7575), .A2(n7571), .ZN(n7711) );
  INV_X1 U9335 ( .A(n7711), .ZN(n7572) );
  NOR2_X1 U9336 ( .A1(n7573), .A2(n7572), .ZN(n7789) );
  NAND2_X1 U9337 ( .A1(n7574), .A2(n7688), .ZN(n9355) );
  INV_X1 U9338 ( .A(n9463), .ZN(n9353) );
  AND2_X1 U9339 ( .A1(n9463), .A2(n9329), .ZN(n7690) );
  INV_X1 U9340 ( .A(n7690), .ZN(n7642) );
  NAND2_X1 U9341 ( .A1(n9359), .A2(n7783), .ZN(n9327) );
  AND2_X1 U9342 ( .A1(n9337), .A2(n9357), .ZN(n7689) );
  INV_X1 U9343 ( .A(n7689), .ZN(n7641) );
  NAND2_X1 U9344 ( .A1(n7640), .A2(n7641), .ZN(n9324) );
  INV_X1 U9345 ( .A(n9324), .ZN(n9328) );
  NAND2_X1 U9346 ( .A1(n9327), .A2(n9328), .ZN(n9326) );
  NAND2_X1 U9347 ( .A1(n9453), .A2(n9330), .ZN(n7787) );
  OR2_X1 U9348 ( .A1(n9193), .A2(n9391), .ZN(n7730) );
  INV_X1 U9349 ( .A(n7728), .ZN(n7580) );
  NAND2_X1 U9350 ( .A1(n9231), .A2(n9390), .ZN(n7881) );
  INV_X1 U9351 ( .A(n7575), .ZN(n7714) );
  NAND2_X1 U9352 ( .A1(n9287), .A2(n9301), .ZN(n7872) );
  AND2_X1 U9353 ( .A1(n9303), .A2(n9316), .ZN(n7643) );
  INV_X1 U9354 ( .A(n7643), .ZN(n7871) );
  AND2_X1 U9355 ( .A1(n7872), .A2(n7871), .ZN(n7712) );
  NAND2_X1 U9356 ( .A1(n9266), .A2(n9417), .ZN(n7875) );
  NAND2_X1 U9357 ( .A1(n7877), .A2(n7875), .ZN(n7717) );
  INV_X1 U9358 ( .A(n7717), .ZN(n7576) );
  OAI211_X1 U9359 ( .C1(n7714), .C2(n7712), .A(n7723), .B(n7576), .ZN(n7577)
         );
  NAND2_X1 U9360 ( .A1(n7578), .A2(n7577), .ZN(n7579) );
  OAI21_X1 U9361 ( .B1(n7580), .B2(n7881), .A(n7579), .ZN(n7581) );
  NAND2_X1 U9362 ( .A1(n9183), .A2(n9381), .ZN(n7886) );
  INV_X1 U9363 ( .A(n7886), .ZN(n7738) );
  AOI211_X1 U9364 ( .C1(n7730), .C2(n7581), .A(n7727), .B(n7738), .ZN(n7582)
         );
  NAND2_X1 U9365 ( .A1(n9209), .A2(n9402), .ZN(n9201) );
  NAND2_X1 U9366 ( .A1(n7582), .A2(n9201), .ZN(n7753) );
  AOI21_X1 U9367 ( .B1(n7789), .B2(n9294), .A(n7753), .ZN(n7593) );
  INV_X1 U9368 ( .A(n7582), .ZN(n7587) );
  INV_X1 U9369 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9522) );
  OR2_X1 U9370 ( .A1(n7596), .A2(n9522), .ZN(n7585) );
  OR2_X1 U9371 ( .A1(n9183), .A2(n9381), .ZN(n7731) );
  OAI211_X1 U9372 ( .C1(n7587), .C2(n7730), .A(n7741), .B(n7731), .ZN(n7792)
         );
  NAND2_X1 U9373 ( .A1(n8317), .A2(n7590), .ZN(n7592) );
  INV_X1 U9374 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8001) );
  OR2_X1 U9375 ( .A1(n7596), .A2(n8001), .ZN(n7591) );
  OAI22_X1 U9376 ( .A1(n7593), .A2(n7792), .B1(n4650), .B2(n9163), .ZN(n7595)
         );
  INV_X1 U9377 ( .A(n7893), .ZN(n7748) );
  NAND2_X1 U9378 ( .A1(n9173), .A2(n7748), .ZN(n7633) );
  AND2_X1 U9379 ( .A1(n7982), .A2(n9372), .ZN(n7742) );
  INV_X1 U9380 ( .A(n7742), .ZN(n7601) );
  NAND2_X1 U9381 ( .A1(n7633), .A2(n7601), .ZN(n7797) );
  INV_X1 U9382 ( .A(n9163), .ZN(n7594) );
  NOR2_X1 U9383 ( .A1(n9173), .A2(n7748), .ZN(n7634) );
  INV_X1 U9384 ( .A(n7634), .ZN(n7796) );
  OAI22_X1 U9385 ( .A1(n7595), .A2(n7797), .B1(n7594), .B2(n7796), .ZN(n7600)
         );
  OR2_X1 U9386 ( .A1(n7596), .A2(n7009), .ZN(n7597) );
  NOR2_X1 U9387 ( .A1(n9482), .A2(n9163), .ZN(n7795) );
  AOI211_X1 U9388 ( .C1(n7600), .C2(n7816), .A(n7795), .B(n7599), .ZN(n7637)
         );
  NAND2_X1 U9389 ( .A1(n7730), .A2(n7885), .ZN(n9200) );
  XNOR2_X1 U9390 ( .A(n9209), .B(n9402), .ZN(n7882) );
  NAND2_X1 U9391 ( .A1(n7603), .A2(n7875), .ZN(n7874) );
  XNOR2_X1 U9392 ( .A(n9287), .B(n9301), .ZN(n9277) );
  XNOR2_X1 U9393 ( .A(n9303), .B(n9432), .ZN(n9293) );
  NAND4_X1 U9394 ( .A1(n7605), .A2(n7604), .A3(n6630), .A4(n7756), .ZN(n7607)
         );
  NOR2_X1 U9395 ( .A1(n7607), .A2(n7606), .ZN(n7611) );
  NAND4_X1 U9396 ( .A1(n7611), .A2(n7610), .A3(n7609), .A4(n7608), .ZN(n7612)
         );
  NOR2_X1 U9397 ( .A1(n7612), .A2(n7659), .ZN(n7613) );
  NAND3_X1 U9398 ( .A1(n7615), .A2(n7614), .A3(n7613), .ZN(n7616) );
  NOR2_X1 U9399 ( .A1(n7617), .A2(n7616), .ZN(n7618) );
  NAND4_X1 U9400 ( .A1(n7621), .A2(n7620), .A3(n7619), .A4(n7618), .ZN(n7622)
         );
  NOR2_X1 U9401 ( .A1(n7683), .A2(n7622), .ZN(n7623) );
  NAND4_X1 U9402 ( .A1(n7624), .A2(n7625), .A3(n7626), .A4(n7623), .ZN(n7627)
         );
  NOR2_X1 U9403 ( .A1(n9324), .A2(n7627), .ZN(n7628) );
  NAND3_X1 U9404 ( .A1(n9293), .A2(n9311), .A3(n7628), .ZN(n7629) );
  NOR3_X1 U9405 ( .A1(n7874), .A2(n9277), .A3(n7629), .ZN(n7630) );
  NAND4_X1 U9406 ( .A1(n9224), .A2(n7879), .A3(n9252), .A4(n7630), .ZN(n7631)
         );
  NOR3_X1 U9407 ( .A1(n9200), .A2(n7882), .A3(n7631), .ZN(n7632) );
  NAND4_X1 U9408 ( .A1(n7633), .A2(n7887), .A3(n9185), .A4(n7632), .ZN(n7635)
         );
  OR4_X1 U9409 ( .A1(n7635), .A2(n7745), .A3(n7795), .A4(n7634), .ZN(n7751) );
  INV_X1 U9410 ( .A(n7751), .ZN(n7636) );
  NOR2_X1 U9411 ( .A1(n7700), .A2(n9313), .ZN(n7638) );
  OAI22_X1 U9412 ( .A1(n7638), .A2(n9337), .B1(n9357), .B2(n7783), .ZN(n7639)
         );
  AOI21_X1 U9413 ( .B1(n7639), .B2(n7787), .A(n7810), .ZN(n7710) );
  NAND2_X1 U9414 ( .A1(n7705), .A2(n7640), .ZN(n7782) );
  AOI21_X1 U9415 ( .B1(n7642), .B2(n7641), .A(n7782), .ZN(n7791) );
  INV_X1 U9416 ( .A(n7787), .ZN(n7644) );
  INV_X1 U9417 ( .A(n7810), .ZN(n7747) );
  NOR4_X1 U9418 ( .A1(n7791), .A2(n7644), .A3(n7643), .A4(n7747), .ZN(n7709)
         );
  NAND2_X1 U9419 ( .A1(n7645), .A2(n7764), .ZN(n7655) );
  INV_X1 U9420 ( .A(n7648), .ZN(n7653) );
  INV_X1 U9421 ( .A(n7649), .ZN(n7652) );
  INV_X1 U9422 ( .A(n7650), .ZN(n7651) );
  NOR3_X1 U9423 ( .A1(n7653), .A2(n7652), .A3(n7651), .ZN(n7656) );
  OAI21_X1 U9424 ( .B1(n7656), .B2(n7655), .A(n7654), .ZN(n7657) );
  MUX2_X1 U9425 ( .A(n7659), .B(n7658), .S(n7810), .Z(n7660) );
  AOI21_X1 U9426 ( .B1(n7662), .B2(n7661), .A(n7660), .ZN(n7667) );
  NAND2_X1 U9427 ( .A1(n7673), .A2(n7663), .ZN(n7664) );
  MUX2_X1 U9428 ( .A(n7665), .B(n7664), .S(n7747), .Z(n7666) );
  NOR2_X1 U9429 ( .A1(n7667), .A2(n7666), .ZN(n7677) );
  INV_X1 U9430 ( .A(n7668), .ZN(n7669) );
  OAI21_X1 U9431 ( .B1(n7677), .B2(n7669), .A(n7674), .ZN(n7670) );
  NAND3_X1 U9432 ( .A1(n7670), .A2(n7680), .A3(n7678), .ZN(n7671) );
  NAND3_X1 U9433 ( .A1(n7671), .A2(n7675), .A3(n7772), .ZN(n7672) );
  INV_X1 U9434 ( .A(n7673), .ZN(n7676) );
  NAND2_X1 U9435 ( .A1(n7675), .A2(n7674), .ZN(n7769) );
  NOR3_X1 U9436 ( .A1(n7677), .A2(n7676), .A3(n7769), .ZN(n7681) );
  OAI211_X1 U9437 ( .C1(n7769), .C2(n7680), .A(n7679), .B(n7678), .ZN(n7774)
         );
  OAI21_X1 U9438 ( .B1(n7681), .B2(n7774), .A(n7772), .ZN(n7682) );
  AOI211_X1 U9439 ( .C1(n7695), .C2(n7773), .A(n7684), .B(n7683), .ZN(n7685)
         );
  NAND2_X1 U9440 ( .A1(n7692), .A2(n7693), .ZN(n7754) );
  NOR3_X1 U9441 ( .A1(n7685), .A2(n7786), .A3(n7754), .ZN(n7686) );
  AOI211_X1 U9442 ( .C1(n4798), .C2(n7688), .A(n7687), .B(n7686), .ZN(n7691)
         );
  NOR4_X1 U9443 ( .A1(n7691), .A2(n7690), .A3(n7689), .A4(n7810), .ZN(n7704)
         );
  INV_X1 U9444 ( .A(n7692), .ZN(n7699) );
  INV_X1 U9445 ( .A(n7773), .ZN(n7694) );
  INV_X1 U9446 ( .A(n7777), .ZN(n7697) );
  NAND2_X1 U9447 ( .A1(n7698), .A2(n7696), .ZN(n7779) );
  NOR4_X1 U9448 ( .A1(n7702), .A2(n7701), .A3(n7700), .A4(n7747), .ZN(n7703)
         );
  INV_X1 U9449 ( .A(n7705), .ZN(n7706) );
  OAI21_X1 U9450 ( .B1(n7707), .B2(n7706), .A(n7747), .ZN(n7708) );
  MUX2_X1 U9451 ( .A(n7712), .B(n7711), .S(n7810), .Z(n7716) );
  INV_X1 U9452 ( .A(n7872), .ZN(n7713) );
  MUX2_X1 U9453 ( .A(n7714), .B(n7713), .S(n7810), .Z(n7715) );
  MUX2_X1 U9454 ( .A(n7718), .B(n7717), .S(n7810), .Z(n7721) );
  MUX2_X1 U9455 ( .A(n7877), .B(n7719), .S(n7810), .Z(n7720) );
  OAI211_X1 U9456 ( .C1(n7722), .C2(n7721), .A(n7879), .B(n7720), .ZN(n7725)
         );
  MUX2_X1 U9457 ( .A(n7880), .B(n7723), .S(n7810), .Z(n7724) );
  NAND2_X1 U9458 ( .A1(n7725), .A2(n7724), .ZN(n7734) );
  OAI211_X1 U9459 ( .C1(n7734), .C2(n7726), .A(n7881), .B(n9201), .ZN(n7729)
         );
  AOI21_X1 U9460 ( .B1(n7729), .B2(n7728), .A(n7727), .ZN(n7732) );
  NAND2_X1 U9461 ( .A1(n7731), .A2(n7730), .ZN(n7737) );
  INV_X1 U9462 ( .A(n7881), .ZN(n7733) );
  NOR2_X1 U9463 ( .A1(n7734), .A2(n7733), .ZN(n7736) );
  OAI211_X1 U9464 ( .C1(n7736), .C2(n7735), .A(n7885), .B(n9201), .ZN(n7740)
         );
  INV_X1 U9465 ( .A(n7737), .ZN(n7739) );
  MUX2_X1 U9466 ( .A(n7747), .B(n7746), .S(n9173), .Z(n7749) );
  OAI21_X1 U9467 ( .B1(n7808), .B2(n7804), .A(n5806), .ZN(n7752) );
  INV_X1 U9468 ( .A(n7753), .ZN(n7794) );
  INV_X1 U9469 ( .A(n7754), .ZN(n7781) );
  INV_X1 U9470 ( .A(n7755), .ZN(n7768) );
  AOI21_X1 U9471 ( .B1(n9044), .B2(n7757), .A(n7756), .ZN(n7762) );
  NAND2_X1 U9472 ( .A1(n9043), .A2(n7758), .ZN(n7760) );
  AND4_X1 U9473 ( .A1(n7762), .A2(n7761), .A3(n7760), .A4(n7759), .ZN(n7765)
         );
  NAND3_X1 U9474 ( .A1(n7765), .A2(n7764), .A3(n7763), .ZN(n7766) );
  NAND3_X1 U9475 ( .A1(n7768), .A2(n7767), .A3(n7766), .ZN(n7771) );
  AOI21_X1 U9476 ( .B1(n7771), .B2(n7770), .A(n7769), .ZN(n7775) );
  OAI211_X1 U9477 ( .C1(n7775), .C2(n7774), .A(n7773), .B(n7772), .ZN(n7778)
         );
  NAND3_X1 U9478 ( .A1(n7778), .A2(n7777), .A3(n7776), .ZN(n7780) );
  AOI21_X1 U9479 ( .B1(n7781), .B2(n7780), .A(n7779), .ZN(n7785) );
  INV_X1 U9480 ( .A(n7782), .ZN(n7784) );
  OAI211_X1 U9481 ( .C1(n7786), .C2(n7785), .A(n7784), .B(n7783), .ZN(n7788)
         );
  NAND2_X1 U9482 ( .A1(n7788), .A2(n7787), .ZN(n7790) );
  OAI21_X1 U9483 ( .B1(n7791), .B2(n7790), .A(n7789), .ZN(n7793) );
  AOI21_X1 U9484 ( .B1(n7794), .B2(n7793), .A(n7792), .ZN(n7798) );
  OAI211_X1 U9485 ( .C1(n7798), .C2(n7797), .A(n7796), .B(n4454), .ZN(n7799)
         );
  NAND2_X1 U9486 ( .A1(n7799), .A2(n7816), .ZN(n7800) );
  XNOR2_X1 U9487 ( .A(n7800), .B(n7844), .ZN(n7802) );
  NAND3_X1 U9488 ( .A1(n9647), .A2(n9058), .A3(n7803), .ZN(n7806) );
  INV_X1 U9489 ( .A(n7804), .ZN(n7805) );
  OR2_X1 U9490 ( .A1(n7819), .A2(n7805), .ZN(n7812) );
  OAI211_X1 U9491 ( .C1(n7807), .C2(n7806), .A(P1_B_REG_SCAN_IN), .B(n7812), 
        .ZN(n7818) );
  INV_X1 U9492 ( .A(n7808), .ZN(n7809) );
  OAI21_X1 U9493 ( .B1(n7810), .B2(n4454), .A(n7809), .ZN(n7814) );
  NOR2_X1 U9494 ( .A1(n7812), .A2(n7811), .ZN(n7813) );
  OAI211_X1 U9495 ( .C1(n7816), .C2(n7815), .A(n7814), .B(n7813), .ZN(n7817)
         );
  NAND2_X1 U9496 ( .A1(n7901), .A2(n7820), .ZN(n7822) );
  OAI211_X1 U9497 ( .C1(n8860), .C2(n7823), .A(n7822), .B(n7821), .ZN(P2_U3267) );
  OAI222_X1 U9498 ( .A1(n8860), .A2(n7825), .B1(n8858), .B2(n9524), .C1(n7824), 
        .C2(P2_U3151), .ZN(P2_U3266) );
  AOI22_X1 U9499 ( .A1(n7829), .A2(n7828), .B1(n7827), .B2(n7826), .ZN(n9157)
         );
  INV_X1 U9500 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9459) );
  AND2_X1 U9501 ( .A1(n7836), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n7830) );
  AOI21_X1 U9502 ( .B1(n9459), .B2(n9151), .A(n7830), .ZN(n9156) );
  NAND2_X1 U9503 ( .A1(n9157), .A2(n9156), .ZN(n9155) );
  INV_X1 U9504 ( .A(n7830), .ZN(n7831) );
  NAND2_X1 U9505 ( .A1(n9155), .A2(n7831), .ZN(n7832) );
  XOR2_X1 U9506 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n7832), .Z(n7841) );
  OR2_X1 U9507 ( .A1(n7833), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n7834) );
  NAND2_X1 U9508 ( .A1(n7836), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7838) );
  OR2_X1 U9509 ( .A1(n7836), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n7837) );
  AND2_X1 U9510 ( .A1(n7838), .A2(n7837), .ZN(n9148) );
  NAND2_X1 U9511 ( .A1(n9149), .A2(n9148), .ZN(n9147) );
  NAND2_X1 U9512 ( .A1(n9147), .A2(n7838), .ZN(n7839) );
  XNOR2_X1 U9513 ( .A(n7839), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n7843) );
  INV_X1 U9514 ( .A(n7843), .ZN(n7840) );
  AOI22_X1 U9515 ( .A1(n7841), .A2(n9575), .B1(n9580), .B2(n7840), .ZN(n7846)
         );
  OAI21_X1 U9516 ( .B1(n7841), .B2(n9528), .A(n9584), .ZN(n7842) );
  AOI21_X1 U9517 ( .B1(n7843), .B2(n9580), .A(n7842), .ZN(n7845) );
  MUX2_X1 U9518 ( .A(n7846), .B(n7845), .S(n7844), .Z(n7847) );
  NAND2_X1 U9519 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8902) );
  OAI211_X1 U9520 ( .C1(n4691), .C2(n9590), .A(n7847), .B(n8902), .ZN(P1_U3262) );
  NAND2_X1 U9521 ( .A1(n9468), .A2(n9031), .ZN(n9345) );
  NAND2_X1 U9522 ( .A1(n9463), .A2(n9030), .ZN(n7848) );
  AND2_X1 U9523 ( .A1(n9345), .A2(n7848), .ZN(n7849) );
  OR2_X1 U9524 ( .A1(n9463), .A2(n9030), .ZN(n7851) );
  NOR2_X1 U9525 ( .A1(n9337), .A2(n9313), .ZN(n7852) );
  NAND2_X1 U9526 ( .A1(n9337), .A2(n9313), .ZN(n7853) );
  AND2_X1 U9527 ( .A1(n9453), .A2(n9440), .ZN(n7854) );
  NOR2_X1 U9528 ( .A1(n9303), .A2(n9432), .ZN(n7856) );
  NAND2_X1 U9529 ( .A1(n9303), .A2(n9432), .ZN(n7855) );
  AND2_X1 U9530 ( .A1(n9287), .A2(n9442), .ZN(n7857) );
  OR2_X1 U9531 ( .A1(n9287), .A2(n9442), .ZN(n7858) );
  NAND2_X1 U9532 ( .A1(n9266), .A2(n9433), .ZN(n7860) );
  NOR2_X1 U9533 ( .A1(n9507), .A2(n9270), .ZN(n7862) );
  NAND2_X1 U9534 ( .A1(n9507), .A2(n9270), .ZN(n7863) );
  NOR2_X1 U9535 ( .A1(n9243), .A2(n9414), .ZN(n7864) );
  AND2_X1 U9536 ( .A1(n9231), .A2(n9211), .ZN(n7865) );
  OR2_X1 U9537 ( .A1(n9231), .A2(n9211), .ZN(n7866) );
  NOR2_X1 U9538 ( .A1(n9209), .A2(n9194), .ZN(n7867) );
  INV_X1 U9539 ( .A(n9200), .ZN(n7883) );
  OR2_X1 U9540 ( .A1(n9193), .A2(n9029), .ZN(n7868) );
  INV_X1 U9541 ( .A(n9381), .ZN(n9028) );
  INV_X1 U9542 ( .A(n9277), .ZN(n9279) );
  NAND2_X1 U9543 ( .A1(n7873), .A2(n7872), .ZN(n9274) );
  INV_X1 U9544 ( .A(n7874), .ZN(n9273) );
  NAND2_X1 U9545 ( .A1(n9274), .A2(n9273), .ZN(n7876) );
  NAND2_X1 U9546 ( .A1(n7876), .A2(n7875), .ZN(n9253) );
  NAND2_X1 U9547 ( .A1(n9223), .A2(n7881), .ZN(n9218) );
  INV_X1 U9548 ( .A(n7882), .ZN(n9217) );
  NAND2_X1 U9549 ( .A1(n9216), .A2(n9201), .ZN(n7884) );
  XNOR2_X1 U9550 ( .A(n7888), .B(n7887), .ZN(n7986) );
  NOR2_X2 U9551 ( .A1(n9349), .A2(n9463), .ZN(n9334) );
  NOR2_X2 U9552 ( .A1(n9266), .A2(n9281), .ZN(n9265) );
  NAND2_X1 U9553 ( .A1(n9487), .A2(n9192), .ZN(n9177) );
  AOI21_X1 U9554 ( .B1(n7982), .B2(n9177), .A(n9348), .ZN(n7889) );
  NAND2_X1 U9555 ( .A1(n7889), .A2(n9167), .ZN(n7984) );
  INV_X1 U9556 ( .A(P1_B_REG_SCAN_IN), .ZN(n7890) );
  NOR2_X1 U9557 ( .A1(n7891), .A2(n7890), .ZN(n7892) );
  NOR2_X1 U9558 ( .A1(n9670), .A2(n7892), .ZN(n9162) );
  NAND2_X1 U9559 ( .A1(n7893), .A2(n9162), .ZN(n7976) );
  OAI211_X1 U9560 ( .C1(n9381), .C2(n9672), .A(n7984), .B(n7976), .ZN(n7894)
         );
  OR2_X1 U9561 ( .A1(n9685), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n7898) );
  OAI21_X1 U9562 ( .B1(n4459), .B2(n9515), .A(n7900), .ZN(P1_U3519) );
  INV_X1 U9563 ( .A(n7901), .ZN(n7903) );
  OAI222_X1 U9564 ( .A1(n9525), .A2(n7903), .B1(n4353), .B2(P1_U3086), .C1(
        n7902), .C2(n9521), .ZN(P1_U3327) );
  INV_X1 U9565 ( .A(n7905), .ZN(n8366) );
  XNOR2_X1 U9566 ( .A(n7904), .B(n8366), .ZN(n7920) );
  INV_X1 U9567 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n7910) );
  OR3_X1 U9568 ( .A1(n8613), .A2(n7906), .A3(n7905), .ZN(n7907) );
  NAND2_X1 U9569 ( .A1(n7908), .A2(n7907), .ZN(n7909) );
  AOI222_X1 U9570 ( .A1(n9883), .A2(n7909), .B1(n8400), .B2(n9878), .C1(n8631), 
        .C2(n9880), .ZN(n7916) );
  MUX2_X1 U9571 ( .A(n7910), .B(n7916), .S(n9968), .Z(n7912) );
  NAND2_X1 U9572 ( .A1(n8129), .A2(n8850), .ZN(n7911) );
  OAI211_X1 U9573 ( .C1(n7920), .C2(n8821), .A(n7912), .B(n7911), .ZN(P2_U3449) );
  INV_X1 U9574 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n7913) );
  MUX2_X1 U9575 ( .A(n7913), .B(n7916), .S(n9986), .Z(n7915) );
  NAND2_X1 U9576 ( .A1(n8129), .A2(n8761), .ZN(n7914) );
  OAI211_X1 U9577 ( .C1(n7920), .C2(n8747), .A(n7915), .B(n7914), .ZN(P2_U3481) );
  INV_X1 U9578 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n7917) );
  MUX2_X1 U9579 ( .A(n7917), .B(n7916), .S(n8710), .Z(n7919) );
  AOI22_X1 U9580 ( .A1(n8129), .A2(n4350), .B1(n9905), .B2(n8128), .ZN(n7918)
         );
  OAI211_X1 U9581 ( .C1(n7920), .C2(n8699), .A(n7919), .B(n7918), .ZN(P2_U3211) );
  XNOR2_X1 U9582 ( .A(n8259), .B(n6370), .ZN(n7937) );
  INV_X1 U9583 ( .A(n7937), .ZN(n7938) );
  XNOR2_X1 U9584 ( .A(n8849), .B(n6370), .ZN(n7936) );
  XNOR2_X1 U9585 ( .A(n8356), .B(n6370), .ZN(n8134) );
  XNOR2_X1 U9586 ( .A(n7927), .B(n6370), .ZN(n8035) );
  INV_X1 U9587 ( .A(n7927), .ZN(n9956) );
  NAND3_X1 U9588 ( .A1(n9956), .A2(n8059), .A3(n7962), .ZN(n7925) );
  OAI211_X1 U9589 ( .C1(n7962), .C2(n8402), .A(n7926), .B(n7925), .ZN(n7930)
         );
  NAND3_X1 U9590 ( .A1(n7927), .A2(n8059), .A3(n6370), .ZN(n7928) );
  OAI211_X1 U9591 ( .C1(n8402), .C2(n6370), .A(n8356), .B(n7928), .ZN(n7929)
         );
  XNOR2_X1 U9592 ( .A(n8068), .B(n6370), .ZN(n7931) );
  XNOR2_X1 U9593 ( .A(n7931), .B(n8117), .ZN(n8062) );
  AOI21_X1 U9594 ( .B1(n7930), .B2(n7929), .A(n8062), .ZN(n7933) );
  INV_X1 U9595 ( .A(n7931), .ZN(n7932) );
  XNOR2_X1 U9596 ( .A(n8249), .B(n7962), .ZN(n7934) );
  NOR2_X1 U9597 ( .A1(n7934), .A2(n8704), .ZN(n7935) );
  AOI21_X1 U9598 ( .B1(n7934), .B2(n8704), .A(n7935), .ZN(n8112) );
  INV_X1 U9599 ( .A(n7935), .ZN(n8019) );
  XNOR2_X1 U9600 ( .A(n7936), .B(n8173), .ZN(n8020) );
  XNOR2_X1 U9601 ( .A(n7937), .B(n8258), .ZN(n8167) );
  XNOR2_X1 U9602 ( .A(n8837), .B(n6370), .ZN(n7939) );
  NAND2_X1 U9603 ( .A1(n7939), .A2(n8090), .ZN(n8079) );
  NOR2_X1 U9604 ( .A1(n7939), .A2(n8090), .ZN(n8080) );
  XNOR2_X1 U9605 ( .A(n8831), .B(n6370), .ZN(n7940) );
  XNOR2_X1 U9606 ( .A(n7940), .B(n8680), .ZN(n8088) );
  XNOR2_X1 U9607 ( .A(n8825), .B(n6370), .ZN(n7941) );
  XNOR2_X1 U9608 ( .A(n7941), .B(n8643), .ZN(n8144) );
  XNOR2_X1 U9609 ( .A(n8744), .B(n6370), .ZN(n7942) );
  XNOR2_X1 U9610 ( .A(n7942), .B(n8656), .ZN(n8045) );
  XNOR2_X1 U9611 ( .A(n8814), .B(n6370), .ZN(n7944) );
  XNOR2_X1 U9612 ( .A(n7944), .B(n8642), .ZN(n8105) );
  XNOR2_X1 U9613 ( .A(n8808), .B(n6370), .ZN(n7945) );
  XNOR2_X1 U9614 ( .A(n7945), .B(n8631), .ZN(n8053) );
  NAND2_X1 U9615 ( .A1(n7945), .A2(n8125), .ZN(n7946) );
  NAND2_X1 U9616 ( .A1(n7947), .A2(n7946), .ZN(n8123) );
  XOR2_X1 U9617 ( .A(n6370), .B(n8129), .Z(n7949) );
  INV_X1 U9618 ( .A(n7949), .ZN(n7948) );
  XNOR2_X1 U9619 ( .A(n7948), .B(n8619), .ZN(n8124) );
  NOR2_X1 U9620 ( .A1(n7949), .A2(n8619), .ZN(n7950) );
  AOI21_X1 U9621 ( .B1(n8123), .B2(n8124), .A(n7950), .ZN(n7953) );
  XNOR2_X1 U9622 ( .A(n8802), .B(n7962), .ZN(n7951) );
  XNOR2_X1 U9623 ( .A(n7953), .B(n7951), .ZN(n8029) );
  NAND2_X1 U9624 ( .A1(n8029), .A2(n8590), .ZN(n7955) );
  INV_X1 U9625 ( .A(n7951), .ZN(n7952) );
  OR2_X1 U9626 ( .A1(n7953), .A2(n7952), .ZN(n7954) );
  NAND2_X1 U9627 ( .A1(n7955), .A2(n7954), .ZN(n8096) );
  XNOR2_X1 U9628 ( .A(n8101), .B(n6370), .ZN(n7956) );
  XNOR2_X1 U9629 ( .A(n7956), .B(n8399), .ZN(n8097) );
  NAND2_X1 U9630 ( .A1(n8096), .A2(n8097), .ZN(n7958) );
  NAND2_X1 U9631 ( .A1(n7956), .A2(n8605), .ZN(n7957) );
  XNOR2_X1 U9632 ( .A(n8076), .B(n6370), .ZN(n7959) );
  XNOR2_X1 U9633 ( .A(n7959), .B(n8569), .ZN(n8072) );
  NAND2_X1 U9634 ( .A1(n8071), .A2(n8072), .ZN(n7961) );
  NAND2_X1 U9635 ( .A1(n7959), .A2(n8589), .ZN(n7960) );
  XNOR2_X1 U9636 ( .A(n8786), .B(n7962), .ZN(n7963) );
  NAND2_X1 U9637 ( .A1(n7963), .A2(n8398), .ZN(n8153) );
  INV_X1 U9638 ( .A(n7963), .ZN(n7964) );
  NAND2_X1 U9639 ( .A1(n7964), .A2(n8579), .ZN(n8154) );
  XNOR2_X1 U9640 ( .A(n8780), .B(n6370), .ZN(n7965) );
  XNOR2_X1 U9641 ( .A(n7965), .B(n8568), .ZN(n8014) );
  INV_X1 U9642 ( .A(n7965), .ZN(n7966) );
  XNOR2_X1 U9643 ( .A(n8543), .B(n6370), .ZN(n7967) );
  INV_X1 U9644 ( .A(n8547), .ZN(n7971) );
  OAI22_X1 U9645 ( .A1(n8305), .A2(n8172), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7968), .ZN(n7969) );
  AOI21_X1 U9646 ( .B1(n8545), .B2(n8170), .A(n7969), .ZN(n7970) );
  OAI21_X1 U9647 ( .B1(n7971), .B2(n8149), .A(n7970), .ZN(n7972) );
  AOI21_X1 U9648 ( .B1(n8548), .B2(n8162), .A(n7972), .ZN(n7973) );
  OAI21_X1 U9649 ( .B1(n7974), .B2(n8164), .A(n7973), .ZN(P2_U3160) );
  OAI22_X1 U9650 ( .A1(n7978), .A2(n7977), .B1(n4352), .B2(n7976), .ZN(n7979)
         );
  AOI21_X1 U9651 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n4352), .A(n7979), .ZN(
        n7980) );
  OAI21_X1 U9652 ( .B1(n9381), .B2(n9181), .A(n7980), .ZN(n7981) );
  AOI21_X1 U9653 ( .B1(n7982), .B2(n9600), .A(n7981), .ZN(n7983) );
  OAI21_X1 U9654 ( .B1(n7984), .B2(n9305), .A(n7983), .ZN(n7985) );
  AOI21_X1 U9655 ( .B1(n7986), .B2(n9307), .A(n7985), .ZN(n7987) );
  OAI21_X1 U9656 ( .B1(n7975), .B2(n9364), .A(n7987), .ZN(P1_U3356) );
  INV_X1 U9657 ( .A(n7988), .ZN(n7989) );
  AOI21_X1 U9658 ( .B1(n8187), .B2(n8343), .A(n7989), .ZN(n9913) );
  OAI21_X1 U9659 ( .B1(n7990), .B2(n8343), .A(n9898), .ZN(n7995) );
  OAI22_X1 U9660 ( .A1(n6687), .A2(n9891), .B1(n7991), .B2(n9893), .ZN(n7994)
         );
  NOR2_X1 U9661 ( .A1(n9913), .A2(n7992), .ZN(n7993) );
  AOI211_X1 U9662 ( .C1(n9883), .C2(n7995), .A(n7994), .B(n7993), .ZN(n9911)
         );
  MUX2_X1 U9663 ( .A(n7996), .B(n9911), .S(n8710), .Z(n7999) );
  AOI22_X1 U9664 ( .A1(n4350), .A2(n7997), .B1(n9905), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n7998) );
  OAI211_X1 U9665 ( .C1(n9913), .C2(n8005), .A(n7999), .B(n7998), .ZN(P2_U3232) );
  INV_X1 U9666 ( .A(n8317), .ZN(n8012) );
  OAI222_X1 U9667 ( .A1(n9521), .A2(n8001), .B1(n9525), .B2(n8012), .C1(
        P1_U3086), .C2(n8000), .ZN(P1_U3325) );
  INV_X1 U9668 ( .A(n8002), .ZN(n8003) );
  NAND2_X1 U9669 ( .A1(n8003), .A2(n9905), .ZN(n8537) );
  OAI21_X1 U9670 ( .B1(n8710), .B2(n8004), .A(n8537), .ZN(n8008) );
  NOR2_X1 U9671 ( .A1(n8006), .A2(n8005), .ZN(n8007) );
  AOI211_X1 U9672 ( .C1(n4350), .C2(n8311), .A(n8008), .B(n8007), .ZN(n8009)
         );
  OAI21_X1 U9673 ( .B1(n8010), .B2(n9910), .A(n8009), .ZN(P2_U3204) );
  OAI222_X1 U9674 ( .A1(P2_U3151), .A2(n8013), .B1(n8858), .B2(n8012), .C1(
        n8860), .C2(n8011), .ZN(P2_U3265) );
  AOI22_X1 U9675 ( .A1(n8398), .A2(n8157), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8016) );
  NAND2_X1 U9676 ( .A1(n8175), .A2(n8560), .ZN(n8015) );
  OAI211_X1 U9677 ( .C1(n8558), .C2(n8160), .A(n8016), .B(n8015), .ZN(n8017)
         );
  AOI21_X1 U9678 ( .B1(n8561), .B2(n8162), .A(n8017), .ZN(n8018) );
  AND3_X1 U9679 ( .A1(n8111), .A2(n8020), .A3(n8019), .ZN(n8021) );
  OAI21_X1 U9680 ( .B1(n8022), .B2(n8021), .A(n4514), .ZN(n8028) );
  INV_X1 U9681 ( .A(n8707), .ZN(n8026) );
  NOR2_X1 U9682 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10129), .ZN(n9814) );
  AOI21_X1 U9683 ( .B1(n8170), .B2(n8703), .A(n9814), .ZN(n8023) );
  OAI21_X1 U9684 ( .B1(n8024), .B2(n8172), .A(n8023), .ZN(n8025) );
  AOI21_X1 U9685 ( .B1(n8026), .B2(n8175), .A(n8025), .ZN(n8027) );
  OAI211_X1 U9686 ( .C1(n8709), .C2(n8178), .A(n8028), .B(n8027), .ZN(P2_U3155) );
  XNOR2_X1 U9687 ( .A(n8029), .B(n8400), .ZN(n8034) );
  INV_X1 U9688 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10043) );
  OAI22_X1 U9689 ( .A1(n8172), .A2(n8604), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10043), .ZN(n8031) );
  NOR2_X1 U9690 ( .A1(n8160), .A2(n8605), .ZN(n8030) );
  AOI211_X1 U9691 ( .C1(n8608), .C2(n8175), .A(n8031), .B(n8030), .ZN(n8033)
         );
  NAND2_X1 U9692 ( .A1(n8609), .A2(n8162), .ZN(n8032) );
  OAI211_X1 U9693 ( .C1(n8034), .C2(n8164), .A(n8033), .B(n8032), .ZN(P2_U3156) );
  XNOR2_X1 U9694 ( .A(n8060), .B(n8403), .ZN(n8036) );
  NAND2_X1 U9695 ( .A1(n8036), .A2(n8035), .ZN(n8136) );
  OAI21_X1 U9696 ( .B1(n8036), .B2(n8035), .A(n8136), .ZN(n8043) );
  NOR2_X1 U9697 ( .A1(n9956), .A2(n8178), .ZN(n8042) );
  NOR2_X1 U9698 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8037), .ZN(n9743) );
  AOI21_X1 U9699 ( .B1(n8157), .B2(n8404), .A(n9743), .ZN(n8039) );
  NAND2_X1 U9700 ( .A1(n8170), .A2(n8402), .ZN(n8038) );
  OAI211_X1 U9701 ( .C1(n8149), .C2(n8040), .A(n8039), .B(n8038), .ZN(n8041)
         );
  AOI211_X1 U9702 ( .C1(n8043), .C2(n4514), .A(n8042), .B(n8041), .ZN(n8044)
         );
  INV_X1 U9703 ( .A(n8044), .ZN(P2_U3157) );
  XOR2_X1 U9704 ( .A(n8046), .B(n8045), .Z(n8051) );
  INV_X1 U9705 ( .A(n8642), .ZN(n8618) );
  AOI22_X1 U9706 ( .A1(n8170), .A2(n8618), .B1(P2_REG3_REG_19__SCAN_IN), .B2(
        P2_U3151), .ZN(n8048) );
  NAND2_X1 U9707 ( .A1(n8157), .A2(n8667), .ZN(n8047) );
  OAI211_X1 U9708 ( .C1(n8149), .C2(n8644), .A(n8048), .B(n8047), .ZN(n8049)
         );
  AOI21_X1 U9709 ( .B1(n8744), .B2(n8162), .A(n8049), .ZN(n8050) );
  OAI21_X1 U9710 ( .B1(n8051), .B2(n8164), .A(n8050), .ZN(P2_U3159) );
  XOR2_X1 U9711 ( .A(n8053), .B(n8052), .Z(n8058) );
  NAND2_X1 U9712 ( .A1(n8175), .A2(n8622), .ZN(n8055) );
  AOI22_X1 U9713 ( .A1(n8170), .A2(n8619), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8054) );
  OAI211_X1 U9714 ( .C1(n8642), .C2(n8172), .A(n8055), .B(n8054), .ZN(n8056)
         );
  AOI21_X1 U9715 ( .B1(n8808), .B2(n8162), .A(n8056), .ZN(n8057) );
  OAI21_X1 U9716 ( .B1(n8058), .B2(n8164), .A(n8057), .ZN(P2_U3163) );
  NAND2_X1 U9717 ( .A1(n8060), .A2(n8059), .ZN(n8135) );
  NAND3_X1 U9718 ( .A1(n8136), .A2(n8134), .A3(n8135), .ZN(n8133) );
  OAI21_X1 U9719 ( .B1(n8063), .B2(n8134), .A(n8133), .ZN(n8061) );
  XOR2_X1 U9720 ( .A(n8062), .B(n8061), .Z(n8070) );
  INV_X1 U9721 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10141) );
  NOR2_X1 U9722 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10141), .ZN(n9777) );
  NOR2_X1 U9723 ( .A1(n8172), .A2(n8063), .ZN(n8064) );
  AOI211_X1 U9724 ( .C1(n8170), .C2(n8704), .A(n9777), .B(n8064), .ZN(n8065)
         );
  OAI21_X1 U9725 ( .B1(n8066), .B2(n8149), .A(n8065), .ZN(n8067) );
  AOI21_X1 U9726 ( .B1(n8068), .B2(n8162), .A(n8067), .ZN(n8069) );
  OAI21_X1 U9727 ( .B1(n8070), .B2(n8164), .A(n8069), .ZN(P2_U3164) );
  XOR2_X1 U9728 ( .A(n8072), .B(n8071), .Z(n8078) );
  AOI22_X1 U9729 ( .A1(n8398), .A2(n8170), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8074) );
  NAND2_X1 U9730 ( .A1(n8175), .A2(n8581), .ZN(n8073) );
  OAI211_X1 U9731 ( .C1(n8605), .C2(n8172), .A(n8074), .B(n8073), .ZN(n8075)
         );
  AOI21_X1 U9732 ( .B1(n8076), .B2(n8162), .A(n8075), .ZN(n8077) );
  OAI21_X1 U9733 ( .B1(n8078), .B2(n8164), .A(n8077), .ZN(P2_U3165) );
  NOR2_X1 U9734 ( .A1(n8080), .A2(n4545), .ZN(n8081) );
  XNOR2_X1 U9735 ( .A(n8082), .B(n8081), .ZN(n8087) );
  NOR2_X1 U9736 ( .A1(n10109), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9848) );
  NOR2_X1 U9737 ( .A1(n8172), .A2(n8258), .ZN(n8083) );
  AOI211_X1 U9738 ( .C1(n8170), .C2(n8680), .A(n9848), .B(n8083), .ZN(n8084)
         );
  OAI21_X1 U9739 ( .B1(n8683), .B2(n8149), .A(n8084), .ZN(n8085) );
  AOI21_X1 U9740 ( .B1(n8837), .B2(n8162), .A(n8085), .ZN(n8086) );
  OAI21_X1 U9741 ( .B1(n8087), .B2(n8164), .A(n8086), .ZN(P2_U3166) );
  XOR2_X1 U9742 ( .A(n8089), .B(n8088), .Z(n8095) );
  AOI22_X1 U9743 ( .A1(n8170), .A2(n8667), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3151), .ZN(n8092) );
  NAND2_X1 U9744 ( .A1(n8157), .A2(n8691), .ZN(n8091) );
  OAI211_X1 U9745 ( .C1(n8149), .C2(n8670), .A(n8092), .B(n8091), .ZN(n8093)
         );
  AOI21_X1 U9746 ( .B1(n8831), .B2(n8162), .A(n8093), .ZN(n8094) );
  OAI21_X1 U9747 ( .B1(n8095), .B2(n8164), .A(n8094), .ZN(P2_U3168) );
  XOR2_X1 U9748 ( .A(n8097), .B(n8096), .Z(n8103) );
  AOI22_X1 U9749 ( .A1(n8569), .A2(n8170), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8099) );
  NAND2_X1 U9750 ( .A1(n8175), .A2(n8592), .ZN(n8098) );
  OAI211_X1 U9751 ( .C1(n8590), .C2(n8172), .A(n8099), .B(n8098), .ZN(n8100)
         );
  AOI21_X1 U9752 ( .B1(n8101), .B2(n8162), .A(n8100), .ZN(n8102) );
  OAI21_X1 U9753 ( .B1(n8103), .B2(n8164), .A(n8102), .ZN(P2_U3169) );
  XOR2_X1 U9754 ( .A(n8105), .B(n8104), .Z(n8110) );
  AOI22_X1 U9755 ( .A1(n8170), .A2(n8631), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8107) );
  NAND2_X1 U9756 ( .A1(n8157), .A2(n8656), .ZN(n8106) );
  OAI211_X1 U9757 ( .C1(n8149), .C2(n8634), .A(n8107), .B(n8106), .ZN(n8108)
         );
  AOI21_X1 U9758 ( .B1(n8814), .B2(n8162), .A(n8108), .ZN(n8109) );
  OAI21_X1 U9759 ( .B1(n8110), .B2(n8164), .A(n8109), .ZN(P2_U3173) );
  OAI21_X1 U9760 ( .B1(n8113), .B2(n8112), .A(n8111), .ZN(n8114) );
  NAND2_X1 U9761 ( .A1(n8114), .A2(n4514), .ZN(n8121) );
  INV_X1 U9762 ( .A(n8115), .ZN(n8119) );
  NOR2_X1 U9763 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6020), .ZN(n9795) );
  AOI21_X1 U9764 ( .B1(n8170), .B2(n8692), .A(n9795), .ZN(n8116) );
  OAI21_X1 U9765 ( .B1(n8117), .B2(n8172), .A(n8116), .ZN(n8118) );
  AOI21_X1 U9766 ( .B1(n8119), .B2(n8175), .A(n8118), .ZN(n8120) );
  OAI211_X1 U9767 ( .C1(n8122), .C2(n8178), .A(n8121), .B(n8120), .ZN(P2_U3174) );
  XOR2_X1 U9768 ( .A(n8124), .B(n8123), .Z(n8132) );
  OAI22_X1 U9769 ( .A1(n8172), .A2(n8125), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10107), .ZN(n8127) );
  NOR2_X1 U9770 ( .A1(n8160), .A2(n8590), .ZN(n8126) );
  AOI211_X1 U9771 ( .C1(n8128), .C2(n8175), .A(n8127), .B(n8126), .ZN(n8131)
         );
  NAND2_X1 U9772 ( .A1(n8129), .A2(n8162), .ZN(n8130) );
  OAI211_X1 U9773 ( .C1(n8132), .C2(n8164), .A(n8131), .B(n8130), .ZN(P2_U3175) );
  NAND2_X1 U9774 ( .A1(n8133), .A2(n4514), .ZN(n8143) );
  AOI21_X1 U9775 ( .B1(n8136), .B2(n8135), .A(n8134), .ZN(n8142) );
  INV_X1 U9776 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n10191) );
  NOR2_X1 U9777 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10191), .ZN(n9760) );
  AOI21_X1 U9778 ( .B1(n8157), .B2(n8403), .A(n9760), .ZN(n8138) );
  NAND2_X1 U9779 ( .A1(n8170), .A2(n8401), .ZN(n8137) );
  OAI211_X1 U9780 ( .C1(n8149), .C2(n8139), .A(n8138), .B(n8137), .ZN(n8140)
         );
  AOI21_X1 U9781 ( .B1(n9966), .B2(n8162), .A(n8140), .ZN(n8141) );
  OAI21_X1 U9782 ( .B1(n8143), .B2(n8142), .A(n8141), .ZN(P2_U3176) );
  XOR2_X1 U9783 ( .A(n8145), .B(n8144), .Z(n8152) );
  AND2_X1 U9784 ( .A1(P2_U3151), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8505) );
  NOR2_X1 U9785 ( .A1(n8172), .A2(n8146), .ZN(n8147) );
  AOI211_X1 U9786 ( .C1(n8170), .C2(n8656), .A(n8505), .B(n8147), .ZN(n8148)
         );
  OAI21_X1 U9787 ( .B1(n8659), .B2(n8149), .A(n8148), .ZN(n8150) );
  AOI21_X1 U9788 ( .B1(n8825), .B2(n8162), .A(n8150), .ZN(n8151) );
  OAI21_X1 U9789 ( .B1(n8152), .B2(n8164), .A(n8151), .ZN(P2_U3178) );
  NAND2_X1 U9790 ( .A1(n8154), .A2(n8153), .ZN(n8155) );
  XNOR2_X1 U9791 ( .A(n8156), .B(n8155), .ZN(n8165) );
  AOI22_X1 U9792 ( .A1(n8569), .A2(n8157), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8159) );
  NAND2_X1 U9793 ( .A1(n8175), .A2(n8572), .ZN(n8158) );
  OAI211_X1 U9794 ( .C1(n8305), .C2(n8160), .A(n8159), .B(n8158), .ZN(n8161)
         );
  AOI21_X1 U9795 ( .B1(n8786), .B2(n8162), .A(n8161), .ZN(n8163) );
  OAI21_X1 U9796 ( .B1(n8165), .B2(n8164), .A(n8163), .ZN(P2_U3180) );
  OAI211_X1 U9797 ( .C1(n8168), .C2(n8167), .A(n8166), .B(n4514), .ZN(n8177)
         );
  INV_X1 U9798 ( .A(n8169), .ZN(n8695) );
  INV_X1 U9799 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10149) );
  NOR2_X1 U9800 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10149), .ZN(n9831) );
  AOI21_X1 U9801 ( .B1(n8170), .B2(n8691), .A(n9831), .ZN(n8171) );
  OAI21_X1 U9802 ( .B1(n8173), .B2(n8172), .A(n8171), .ZN(n8174) );
  AOI21_X1 U9803 ( .B1(n8695), .B2(n8175), .A(n8174), .ZN(n8176) );
  OAI211_X1 U9804 ( .C1(n8259), .C2(n8178), .A(n8177), .B(n8176), .ZN(P2_U3181) );
  INV_X1 U9805 ( .A(n8340), .ZN(n8292) );
  INV_X1 U9806 ( .A(n8339), .ZN(n8179) );
  AOI21_X1 U9807 ( .B1(n8292), .B2(n8295), .A(n8179), .ZN(n8296) );
  NAND2_X1 U9808 ( .A1(n8181), .A2(n8180), .ZN(n8186) );
  NOR2_X1 U9809 ( .A1(n8186), .A2(n8182), .ZN(n8184) );
  MUX2_X1 U9810 ( .A(n8315), .B(n8184), .S(n8183), .Z(n8185) );
  INV_X1 U9811 ( .A(n8185), .ZN(n8190) );
  NAND3_X1 U9812 ( .A1(n8187), .A2(n8186), .A3(n8315), .ZN(n8188) );
  NAND3_X1 U9813 ( .A1(n8190), .A2(n9897), .A3(n8189), .ZN(n8198) );
  NAND2_X1 U9814 ( .A1(n9881), .A2(n8191), .ZN(n8208) );
  NAND2_X1 U9815 ( .A1(n8208), .A2(n8192), .ZN(n8195) );
  NAND2_X1 U9816 ( .A1(n8193), .A2(n8200), .ZN(n8194) );
  MUX2_X1 U9817 ( .A(n8195), .B(n8194), .S(n8315), .Z(n8196) );
  INV_X1 U9818 ( .A(n8196), .ZN(n8197) );
  NAND2_X1 U9819 ( .A1(n8198), .A2(n8197), .ZN(n8199) );
  NAND2_X1 U9820 ( .A1(n8199), .A2(n9884), .ZN(n8212) );
  INV_X1 U9821 ( .A(n8200), .ZN(n8204) );
  NAND2_X1 U9822 ( .A1(n8202), .A2(n8201), .ZN(n8203) );
  OAI211_X1 U9823 ( .C1(n8212), .C2(n8204), .A(n8203), .B(n8213), .ZN(n8207)
         );
  AND2_X1 U9824 ( .A1(n8209), .A2(n8216), .ZN(n8206) );
  INV_X1 U9825 ( .A(n8214), .ZN(n8205) );
  INV_X1 U9826 ( .A(n8208), .ZN(n8211) );
  OAI211_X1 U9827 ( .C1(n8212), .C2(n8211), .A(n8210), .B(n8209), .ZN(n8215)
         );
  NAND3_X1 U9828 ( .A1(n8215), .A2(n8214), .A3(n8213), .ZN(n8218) );
  AND2_X1 U9829 ( .A1(n8221), .A2(n8220), .ZN(n8223) );
  AND2_X1 U9830 ( .A1(n8227), .A2(n8228), .ZN(n8222) );
  MUX2_X1 U9831 ( .A(n8223), .B(n8222), .S(n8315), .Z(n8225) );
  INV_X1 U9832 ( .A(n8224), .ZN(n8232) );
  INV_X1 U9833 ( .A(n8225), .ZN(n8230) );
  AND2_X1 U9834 ( .A1(n8227), .A2(n8226), .ZN(n8229) );
  OAI211_X1 U9835 ( .C1(n8230), .C2(n8229), .A(n8228), .B(n8238), .ZN(n8231)
         );
  MUX2_X1 U9836 ( .A(n8232), .B(n8231), .S(n8329), .Z(n8233) );
  INV_X1 U9837 ( .A(n8233), .ZN(n8234) );
  NAND2_X1 U9838 ( .A1(n8235), .A2(n8234), .ZN(n8243) );
  NAND2_X1 U9839 ( .A1(n8243), .A2(n8236), .ZN(n8237) );
  AND2_X1 U9840 ( .A1(n8239), .A2(n8238), .ZN(n8242) );
  INV_X1 U9841 ( .A(n8240), .ZN(n8241) );
  AOI21_X1 U9842 ( .B1(n8243), .B2(n8242), .A(n8241), .ZN(n8244) );
  MUX2_X1 U9843 ( .A(n8246), .B(n8245), .S(n8329), .Z(n8247) );
  NAND2_X1 U9844 ( .A1(n8248), .A2(n8247), .ZN(n8254) );
  MUX2_X1 U9845 ( .A(n8704), .B(n8249), .S(n8329), .Z(n8250) );
  INV_X1 U9846 ( .A(n8250), .ZN(n8251) );
  OAI21_X1 U9847 ( .B1(n8254), .B2(n8252), .A(n8251), .ZN(n8256) );
  NAND2_X1 U9848 ( .A1(n8254), .A2(n8253), .ZN(n8255) );
  NAND2_X1 U9849 ( .A1(n8256), .A2(n8255), .ZN(n8257) );
  AND2_X1 U9850 ( .A1(n8260), .A2(n8261), .ZN(n8713) );
  NAND2_X1 U9851 ( .A1(n8257), .A2(n8713), .ZN(n8263) );
  XNOR2_X1 U9852 ( .A(n8259), .B(n8258), .ZN(n8689) );
  MUX2_X1 U9853 ( .A(n8261), .B(n8260), .S(n8329), .Z(n8262) );
  NAND3_X1 U9854 ( .A1(n8263), .A2(n8689), .A3(n8262), .ZN(n8265) );
  MUX2_X1 U9855 ( .A(n8675), .B(n4423), .S(n8329), .Z(n8264) );
  NAND3_X1 U9856 ( .A1(n8265), .A2(n8678), .A3(n8264), .ZN(n8269) );
  NOR2_X1 U9857 ( .A1(n8266), .A2(n8329), .ZN(n8267) );
  NOR2_X1 U9858 ( .A1(n8666), .A2(n8267), .ZN(n8268) );
  NAND2_X1 U9859 ( .A1(n8269), .A2(n8268), .ZN(n8274) );
  NAND2_X1 U9860 ( .A1(n8274), .A2(n8362), .ZN(n8270) );
  NAND2_X1 U9861 ( .A1(n8270), .A2(n8651), .ZN(n8277) );
  INV_X1 U9862 ( .A(n8271), .ZN(n8273) );
  AND2_X1 U9863 ( .A1(n8651), .A2(n8272), .ZN(n8342) );
  OAI21_X1 U9864 ( .B1(n8274), .B2(n8273), .A(n8342), .ZN(n8275) );
  NAND3_X1 U9865 ( .A1(n8275), .A2(n8652), .A3(n8281), .ZN(n8276) );
  MUX2_X1 U9866 ( .A(n8277), .B(n8276), .S(n8329), .Z(n8284) );
  NAND3_X1 U9867 ( .A1(n8284), .A2(n8280), .A3(n8285), .ZN(n8278) );
  NAND3_X1 U9868 ( .A1(n8278), .A2(n8287), .A3(n8282), .ZN(n8279) );
  NAND2_X1 U9869 ( .A1(n8279), .A2(n8286), .ZN(n8288) );
  INV_X1 U9870 ( .A(n8280), .ZN(n8283) );
  NAND2_X1 U9871 ( .A1(n8289), .A2(n8366), .ZN(n8294) );
  MUX2_X1 U9872 ( .A(n8291), .B(n8290), .S(n8329), .Z(n8293) );
  INV_X1 U9873 ( .A(n8297), .ZN(n8302) );
  MUX2_X1 U9874 ( .A(n8299), .B(n8298), .S(n8329), .Z(n8300) );
  NAND3_X1 U9875 ( .A1(n8301), .A2(n8564), .A3(n8300), .ZN(n8310) );
  MUX2_X1 U9876 ( .A(n8303), .B(n8302), .S(n8329), .Z(n8304) );
  NOR2_X1 U9877 ( .A1(n8555), .A2(n8304), .ZN(n8309) );
  AND2_X1 U9878 ( .A1(n8305), .A2(n8315), .ZN(n8307) );
  NOR2_X1 U9879 ( .A1(n8305), .A2(n8315), .ZN(n8306) );
  MUX2_X1 U9880 ( .A(n8307), .B(n8306), .S(n8780), .Z(n8308) );
  AOI21_X1 U9881 ( .B1(n8310), .B2(n8309), .A(n8308), .ZN(n8327) );
  NAND2_X1 U9882 ( .A1(n8311), .A2(n8329), .ZN(n8314) );
  NOR2_X1 U9883 ( .A1(n8312), .A2(n8315), .ZN(n8313) );
  AOI21_X1 U9884 ( .B1(n8377), .B2(n8314), .A(n8313), .ZN(n8325) );
  MUX2_X1 U9885 ( .A(n8558), .B(n8778), .S(n8315), .Z(n8326) );
  NAND2_X1 U9886 ( .A1(n8317), .A2(n8316), .ZN(n8319) );
  OR2_X1 U9887 ( .A1(n8320), .A2(n8011), .ZN(n8318) );
  NOR2_X1 U9888 ( .A1(n8379), .A2(n8329), .ZN(n8334) );
  OAI22_X1 U9889 ( .A1(n8322), .A2(n8321), .B1(n8320), .B2(n6500), .ZN(n8766)
         );
  INV_X1 U9890 ( .A(n8766), .ZN(n8539) );
  NAND2_X1 U9891 ( .A1(n8539), .A2(n8536), .ZN(n8336) );
  INV_X1 U9892 ( .A(n8396), .ZN(n8323) );
  NAND2_X1 U9893 ( .A1(n8769), .A2(n8323), .ZN(n8333) );
  AOI21_X1 U9894 ( .B1(n8327), .B2(n8326), .A(n8325), .ZN(n8330) );
  INV_X1 U9895 ( .A(n8377), .ZN(n8328) );
  INV_X1 U9896 ( .A(n8330), .ZN(n8331) );
  NOR2_X1 U9897 ( .A1(n8331), .A2(n8397), .ZN(n8335) );
  NAND2_X1 U9898 ( .A1(n8333), .A2(n8332), .ZN(n8376) );
  OAI21_X1 U9899 ( .B1(n8335), .B2(n8376), .A(n8334), .ZN(n8387) );
  INV_X1 U9900 ( .A(n8336), .ZN(n8373) );
  INV_X1 U9901 ( .A(n8337), .ZN(n8372) );
  INV_X1 U9902 ( .A(n8582), .ZN(n8368) );
  NAND2_X1 U9903 ( .A1(n8339), .A2(n8338), .ZN(n8595) );
  NAND2_X1 U9904 ( .A1(n8340), .A2(n8593), .ZN(n8602) );
  INV_X1 U9905 ( .A(n8342), .ZN(n8364) );
  INV_X1 U9906 ( .A(n8689), .ZN(n8360) );
  INV_X1 U9907 ( .A(n8713), .ZN(n8701) );
  NOR4_X1 U9908 ( .A1(n8346), .A2(n8345), .A3(n8344), .A4(n8343), .ZN(n8349)
         );
  NAND4_X1 U9909 ( .A1(n8349), .A2(n8348), .A3(n9884), .A4(n8347), .ZN(n8353)
         );
  NOR4_X1 U9910 ( .A1(n8353), .A2(n8352), .A3(n8351), .A4(n8350), .ZN(n8357)
         );
  NAND4_X1 U9911 ( .A1(n8357), .A2(n8356), .A3(n8355), .A4(n8354), .ZN(n8358)
         );
  NOR4_X1 U9912 ( .A1(n8360), .A2(n8359), .A3(n8701), .A4(n8358), .ZN(n8361)
         );
  NAND3_X1 U9913 ( .A1(n8362), .A2(n8678), .A3(n8361), .ZN(n8363) );
  NOR3_X1 U9914 ( .A1(n8639), .A2(n8364), .A3(n8363), .ZN(n8365) );
  NAND4_X1 U9915 ( .A1(n8366), .A2(n8627), .A3(n8615), .A4(n8365), .ZN(n8367)
         );
  NOR4_X1 U9916 ( .A1(n8368), .A2(n8595), .A3(n8602), .A4(n8367), .ZN(n8370)
         );
  INV_X1 U9917 ( .A(n8555), .ZN(n8369) );
  NAND4_X1 U9918 ( .A1(n8543), .A2(n8564), .A3(n8370), .A4(n8369), .ZN(n8371)
         );
  NOR4_X1 U9919 ( .A1(n8373), .A2(n8372), .A3(n8376), .A4(n8371), .ZN(n8375)
         );
  OAI22_X1 U9920 ( .A1(n8375), .A2(n8374), .B1(n8539), .B2(n8536), .ZN(n8386)
         );
  OAI21_X1 U9921 ( .B1(n8381), .B2(n8379), .A(n8766), .ZN(n8384) );
  NAND3_X1 U9922 ( .A1(n8381), .A2(n8722), .A3(n8380), .ZN(n8383) );
  AOI21_X1 U9923 ( .B1(n8384), .B2(n8383), .A(n8382), .ZN(n8385) );
  XNOR2_X1 U9924 ( .A(n8388), .B(n8516), .ZN(n8395) );
  NOR3_X1 U9925 ( .A1(n8390), .A2(n8389), .A3(n6273), .ZN(n8393) );
  OAI21_X1 U9926 ( .B1(n8394), .B2(n8391), .A(P2_B_REG_SCAN_IN), .ZN(n8392) );
  MUX2_X1 U9927 ( .A(n8396), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8408), .Z(
        P2_U3521) );
  MUX2_X1 U9928 ( .A(n8545), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8408), .Z(
        P2_U3520) );
  MUX2_X1 U9929 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8397), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U9930 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8568), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U9931 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8398), .S(P2_U3893), .Z(
        P2_U3517) );
  MUX2_X1 U9932 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8569), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U9933 ( .A(n8399), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8408), .Z(
        P2_U3515) );
  MUX2_X1 U9934 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n8400), .S(P2_U3893), .Z(
        P2_U3514) );
  MUX2_X1 U9935 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n8619), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U9936 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n8631), .S(P2_U3893), .Z(
        P2_U3512) );
  MUX2_X1 U9937 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n8618), .S(P2_U3893), .Z(
        P2_U3511) );
  MUX2_X1 U9938 ( .A(n8656), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8408), .Z(
        P2_U3510) );
  MUX2_X1 U9939 ( .A(n8667), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8408), .Z(
        P2_U3509) );
  MUX2_X1 U9940 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n8680), .S(P2_U3893), .Z(
        P2_U3508) );
  MUX2_X1 U9941 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n8691), .S(P2_U3893), .Z(
        P2_U3507) );
  MUX2_X1 U9942 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n8703), .S(P2_U3893), .Z(
        P2_U3506) );
  MUX2_X1 U9943 ( .A(n8692), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8408), .Z(
        P2_U3505) );
  MUX2_X1 U9944 ( .A(n8704), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8408), .Z(
        P2_U3504) );
  MUX2_X1 U9945 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n8401), .S(P2_U3893), .Z(
        P2_U3503) );
  MUX2_X1 U9946 ( .A(n8402), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8408), .Z(
        P2_U3502) );
  MUX2_X1 U9947 ( .A(n8403), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8408), .Z(
        P2_U3501) );
  MUX2_X1 U9948 ( .A(n8404), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8408), .Z(
        P2_U3500) );
  MUX2_X1 U9949 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n8405), .S(P2_U3893), .Z(
        P2_U3499) );
  MUX2_X1 U9950 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8406), .S(P2_U3893), .Z(
        P2_U3498) );
  MUX2_X1 U9951 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n8407), .S(P2_U3893), .Z(
        P2_U3497) );
  MUX2_X1 U9952 ( .A(n9879), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8408), .Z(
        P2_U3496) );
  MUX2_X1 U9953 ( .A(n9881), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8408), .Z(
        P2_U3494) );
  MUX2_X1 U9954 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n8409), .S(P2_U3893), .Z(
        P2_U3493) );
  MUX2_X1 U9955 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8410), .S(P2_U3893), .Z(
        P2_U3492) );
  OAI21_X1 U9956 ( .B1(n8413), .B2(n8412), .A(n8411), .ZN(n8414) );
  NAND2_X1 U9957 ( .A1(n8414), .A2(n9866), .ZN(n8432) );
  NAND3_X1 U9958 ( .A1(n8417), .A2(n4766), .A3(n8416), .ZN(n8418) );
  AND2_X1 U9959 ( .A1(n8419), .A2(n8418), .ZN(n8424) );
  INV_X1 U9960 ( .A(n8420), .ZN(n8421) );
  NAND2_X1 U9961 ( .A1(n9858), .A2(n8421), .ZN(n8422) );
  OAI211_X1 U9962 ( .C1(n9872), .C2(n8424), .A(n8423), .B(n8422), .ZN(n8425)
         );
  AOI21_X1 U9963 ( .B1(n9857), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n8425), .ZN(
        n8431) );
  OAI21_X1 U9964 ( .B1(n8428), .B2(n8427), .A(n8426), .ZN(n8429) );
  NAND2_X1 U9965 ( .A1(n9867), .A2(n8429), .ZN(n8430) );
  NAND3_X1 U9966 ( .A1(n8432), .A2(n8431), .A3(n8430), .ZN(P2_U3188) );
  NOR2_X1 U9967 ( .A1(n8513), .A2(n8658), .ZN(n8433) );
  AOI21_X1 U9968 ( .B1(n8658), .B2(n8513), .A(n8433), .ZN(n8450) );
  INV_X1 U9969 ( .A(n8434), .ZN(n9702) );
  MUX2_X1 U9970 ( .A(n8435), .B(P2_REG2_REG_8__SCAN_IN), .S(n8489), .Z(n9703)
         );
  MUX2_X1 U9971 ( .A(n8437), .B(P2_REG2_REG_10__SCAN_IN), .S(n8481), .Z(n9745)
         );
  NOR2_X1 U9972 ( .A1(n9752), .A2(n8438), .ZN(n8439) );
  NOR2_X1 U9973 ( .A1(n7423), .A2(n9762), .ZN(n9761) );
  XNOR2_X1 U9974 ( .A(n9768), .B(n8440), .ZN(n9781) );
  OR2_X1 U9975 ( .A1(n9768), .A2(n8440), .ZN(n8441) );
  INV_X1 U9976 ( .A(n8443), .ZN(n8442) );
  NAND2_X1 U9977 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n8473), .ZN(n8445) );
  OAI21_X1 U9978 ( .B1(n8473), .B2(P2_REG2_REG_14__SCAN_IN), .A(n8445), .ZN(
        n9816) );
  NAND2_X1 U9979 ( .A1(P2_REG2_REG_16__SCAN_IN), .A2(n8469), .ZN(n8447) );
  OAI21_X1 U9980 ( .B1(n8469), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8447), .ZN(
        n9850) );
  AOI21_X1 U9981 ( .B1(n8450), .B2(n8449), .A(n8512), .ZN(n8511) );
  AOI22_X1 U9982 ( .A1(P2_REG1_REG_16__SCAN_IN), .A2(n8469), .B1(n9839), .B2(
        n8754), .ZN(n9842) );
  NAND2_X1 U9983 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8473), .ZN(n8463) );
  AOI22_X1 U9984 ( .A1(P2_REG1_REG_14__SCAN_IN), .A2(n8473), .B1(n9805), .B2(
        n8760), .ZN(n9808) );
  INV_X1 U9985 ( .A(n9768), .ZN(n8451) );
  NAND2_X1 U9986 ( .A1(n8451), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n8460) );
  XNOR2_X1 U9987 ( .A(n9768), .B(P2_REG1_REG_12__SCAN_IN), .ZN(n9770) );
  MUX2_X1 U9988 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n8452), .S(n8481), .Z(n9739)
         );
  AOI22_X1 U9989 ( .A1(n8455), .A2(P2_REG1_REG_7__SCAN_IN), .B1(n8454), .B2(
        n8453), .ZN(n9698) );
  MUX2_X1 U9990 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n5954), .S(n8489), .Z(n9697)
         );
  OAI21_X1 U9991 ( .B1(n8489), .B2(n5954), .A(n9701), .ZN(n8456) );
  NAND2_X1 U9992 ( .A1(n4769), .A2(n8456), .ZN(n8457) );
  XNOR2_X1 U9993 ( .A(n8456), .B(n9718), .ZN(n9723) );
  NAND2_X1 U9994 ( .A1(P2_REG1_REG_9__SCAN_IN), .A2(n9723), .ZN(n9722) );
  NAND2_X1 U9995 ( .A1(n8457), .A2(n9722), .ZN(n9740) );
  NAND2_X1 U9996 ( .A1(n9739), .A2(n9740), .ZN(n9738) );
  NAND2_X1 U9997 ( .A1(n8479), .A2(n8458), .ZN(n8459) );
  XNOR2_X1 U9998 ( .A(n8458), .B(n9752), .ZN(n9754) );
  NAND2_X1 U9999 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n9754), .ZN(n9753) );
  NAND2_X1 U10000 ( .A1(n8459), .A2(n9753), .ZN(n9771) );
  NAND2_X1 U10001 ( .A1(n9770), .A2(n9771), .ZN(n9769) );
  NAND2_X1 U10002 ( .A1(n8475), .A2(n8461), .ZN(n8462) );
  XNOR2_X1 U10003 ( .A(n8461), .B(n9787), .ZN(n9789) );
  NAND2_X1 U10004 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n9789), .ZN(n9788) );
  NAND2_X1 U10005 ( .A1(n8462), .A2(n9788), .ZN(n9807) );
  NAND2_X1 U10006 ( .A1(n9808), .A2(n9807), .ZN(n9806) );
  NAND2_X1 U10007 ( .A1(n8463), .A2(n9806), .ZN(n8464) );
  NAND2_X1 U10008 ( .A1(n8471), .A2(n8464), .ZN(n8465) );
  XOR2_X1 U10009 ( .A(n8471), .B(n8464), .Z(n9825) );
  NAND2_X1 U10010 ( .A1(n9842), .A2(n9841), .ZN(n9840) );
  NAND2_X1 U10011 ( .A1(n8468), .A2(n8466), .ZN(n8467) );
  XOR2_X1 U10012 ( .A(n8468), .B(n8466), .Z(n9861) );
  NAND2_X1 U10013 ( .A1(P2_REG1_REG_17__SCAN_IN), .A2(n9861), .ZN(n9860) );
  XNOR2_X1 U10014 ( .A(n8521), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8514) );
  XNOR2_X1 U10015 ( .A(n8515), .B(n8514), .ZN(n8509) );
  MUX2_X1 U10016 ( .A(n8669), .B(n8751), .S(n8856), .Z(n8499) );
  XNOR2_X1 U10017 ( .A(n8499), .B(n8468), .ZN(n9864) );
  MUX2_X1 U10018 ( .A(P2_REG2_REG_16__SCAN_IN), .B(P2_REG1_REG_16__SCAN_IN), 
        .S(n8856), .Z(n8470) );
  OR2_X1 U10019 ( .A1(n8470), .A2(n8469), .ZN(n8498) );
  XNOR2_X1 U10020 ( .A(n8470), .B(n9839), .ZN(n9845) );
  MUX2_X1 U10021 ( .A(P2_REG2_REG_15__SCAN_IN), .B(P2_REG1_REG_15__SCAN_IN), 
        .S(n8856), .Z(n8472) );
  OR2_X1 U10022 ( .A1(n8472), .A2(n8471), .ZN(n8497) );
  XNOR2_X1 U10023 ( .A(n8472), .B(n9823), .ZN(n9828) );
  MUX2_X1 U10024 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n8856), .Z(n8474) );
  OR2_X1 U10025 ( .A1(n8474), .A2(n8473), .ZN(n8496) );
  XNOR2_X1 U10026 ( .A(n8474), .B(n9805), .ZN(n9811) );
  MUX2_X1 U10027 ( .A(P2_REG2_REG_13__SCAN_IN), .B(P2_REG1_REG_13__SCAN_IN), 
        .S(n8856), .Z(n8476) );
  OR2_X1 U10028 ( .A1(n8476), .A2(n8475), .ZN(n8495) );
  XNOR2_X1 U10029 ( .A(n8476), .B(n9787), .ZN(n9792) );
  MUX2_X1 U10030 ( .A(P2_REG2_REG_12__SCAN_IN), .B(P2_REG1_REG_12__SCAN_IN), 
        .S(n8856), .Z(n8478) );
  INV_X1 U10031 ( .A(n8478), .ZN(n8477) );
  NAND2_X1 U10032 ( .A1(n9768), .A2(n8477), .ZN(n8494) );
  XNOR2_X1 U10033 ( .A(n8478), .B(n9768), .ZN(n9774) );
  MUX2_X1 U10034 ( .A(P2_REG2_REG_11__SCAN_IN), .B(P2_REG1_REG_11__SCAN_IN), 
        .S(n8856), .Z(n8480) );
  OR2_X1 U10035 ( .A1(n8480), .A2(n8479), .ZN(n8493) );
  XNOR2_X1 U10036 ( .A(n8480), .B(n9752), .ZN(n9757) );
  MUX2_X1 U10037 ( .A(P2_REG2_REG_10__SCAN_IN), .B(P2_REG1_REG_10__SCAN_IN), 
        .S(n8856), .Z(n8482) );
  OR2_X1 U10038 ( .A1(n8482), .A2(n8481), .ZN(n8492) );
  XNOR2_X1 U10039 ( .A(n8482), .B(n9734), .ZN(n9737) );
  MUX2_X1 U10040 ( .A(P2_REG2_REG_9__SCAN_IN), .B(P2_REG1_REG_9__SCAN_IN), .S(
        n8856), .Z(n8483) );
  OR2_X1 U10041 ( .A1(n8483), .A2(n4769), .ZN(n8491) );
  XNOR2_X1 U10042 ( .A(n8483), .B(n9718), .ZN(n9720) );
  INV_X1 U10043 ( .A(n8484), .ZN(n8485) );
  AOI22_X1 U10044 ( .A1(n8488), .A2(n8487), .B1(n8486), .B2(n8485), .ZN(n9714)
         );
  MUX2_X1 U10045 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n8856), .Z(n8490) );
  XOR2_X1 U10046 ( .A(n8489), .B(n8490), .Z(n9713) );
  NAND2_X1 U10047 ( .A1(n8491), .A2(n9719), .ZN(n9736) );
  NAND2_X1 U10048 ( .A1(n9757), .A2(n9756), .ZN(n9755) );
  NAND2_X1 U10049 ( .A1(n8494), .A2(n9772), .ZN(n9791) );
  NAND2_X1 U10050 ( .A1(n9792), .A2(n9791), .ZN(n9790) );
  NAND2_X1 U10051 ( .A1(n8495), .A2(n9790), .ZN(n9810) );
  NAND2_X1 U10052 ( .A1(n9811), .A2(n9810), .ZN(n9809) );
  NAND2_X1 U10053 ( .A1(n8496), .A2(n9809), .ZN(n9827) );
  NAND2_X1 U10054 ( .A1(n8497), .A2(n9826), .ZN(n9844) );
  MUX2_X1 U10055 ( .A(P2_REG2_REG_18__SCAN_IN), .B(P2_REG1_REG_18__SCAN_IN), 
        .S(n8856), .Z(n8500) );
  NOR2_X1 U10056 ( .A1(n8501), .A2(n8500), .ZN(n8522) );
  NAND2_X1 U10057 ( .A1(n8501), .A2(n8500), .ZN(n8520) );
  INV_X1 U10058 ( .A(n8520), .ZN(n8502) );
  AOI21_X1 U10059 ( .B1(n8503), .B2(P2_U3893), .A(n9858), .ZN(n8507) );
  NOR3_X1 U10060 ( .A1(n8503), .A2(n8521), .A3(n8529), .ZN(n8504) );
  OAI21_X1 U10061 ( .B1(n8507), .B2(n8513), .A(n8506), .ZN(n8508) );
  OAI21_X1 U10062 ( .B1(n8511), .B2(n9872), .A(n8510), .ZN(P2_U3200) );
  MUX2_X1 U10063 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8645), .S(n8516), .Z(n8519) );
  AOI22_X1 U10064 ( .A1(n8515), .A2(n8514), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8513), .ZN(n8517) );
  XNOR2_X1 U10065 ( .A(n8516), .B(n8745), .ZN(n8518) );
  XNOR2_X1 U10066 ( .A(n8517), .B(n8518), .ZN(n8532) );
  MUX2_X1 U10067 ( .A(n8519), .B(n8518), .S(n6274), .Z(n8524) );
  OAI21_X1 U10068 ( .B1(n8522), .B2(n8521), .A(n8520), .ZN(n8523) );
  XOR2_X1 U10069 ( .A(n8524), .B(n8523), .Z(n8530) );
  NAND2_X1 U10070 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3151), .ZN(n8525) );
  OAI21_X1 U10071 ( .B1(n9708), .B2(n8526), .A(n8525), .ZN(n8527) );
  AOI21_X1 U10072 ( .B1(P2_ADDR_REG_19__SCAN_IN), .B2(n9857), .A(n8527), .ZN(
        n8528) );
  OAI21_X1 U10073 ( .B1(n8530), .B2(n8529), .A(n8528), .ZN(n8531) );
  OAI21_X1 U10074 ( .B1(n8534), .B2(n9872), .A(n8533), .ZN(P2_U3201) );
  NAND2_X1 U10075 ( .A1(n8536), .A2(n8535), .ZN(n8717) );
  AOI21_X1 U10076 ( .B1(n8537), .B2(n8717), .A(n9910), .ZN(n8540) );
  AOI21_X1 U10077 ( .B1(n9910), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8540), .ZN(
        n8538) );
  OAI21_X1 U10078 ( .B1(n8539), .B2(n8542), .A(n8538), .ZN(P2_U3202) );
  AOI21_X1 U10079 ( .B1(n9910), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8540), .ZN(
        n8541) );
  OAI21_X1 U10080 ( .B1(n8722), .B2(n8542), .A(n8541), .ZN(P2_U3203) );
  MUX2_X1 U10081 ( .A(n8546), .B(n8773), .S(n8710), .Z(n8553) );
  AOI22_X1 U10082 ( .A1(n8548), .A2(n4350), .B1(n9905), .B2(n8547), .ZN(n8552)
         );
  XNOR2_X1 U10083 ( .A(n8550), .B(n8549), .ZN(n8775) );
  NAND2_X1 U10084 ( .A1(n8775), .A2(n9888), .ZN(n8551) );
  NAND3_X1 U10085 ( .A1(n8553), .A2(n8552), .A3(n8551), .ZN(P2_U3205) );
  XNOR2_X1 U10086 ( .A(n8554), .B(n8555), .ZN(n8781) );
  XNOR2_X1 U10087 ( .A(n8556), .B(n8555), .ZN(n8557) );
  OAI222_X1 U10088 ( .A1(n9893), .A2(n8558), .B1(n9891), .B2(n8579), .C1(n8557), .C2(n9899), .ZN(n8779) );
  MUX2_X1 U10089 ( .A(P2_REG2_REG_27__SCAN_IN), .B(n8779), .S(n8710), .Z(n8559) );
  INV_X1 U10090 ( .A(n8559), .ZN(n8563) );
  AOI22_X1 U10091 ( .A1(n8561), .A2(n4350), .B1(n9905), .B2(n8560), .ZN(n8562)
         );
  OAI211_X1 U10092 ( .C1(n8781), .C2(n8699), .A(n8563), .B(n8562), .ZN(
        P2_U3206) );
  XNOR2_X1 U10093 ( .A(n8565), .B(n8564), .ZN(n8789) );
  XNOR2_X1 U10094 ( .A(n8567), .B(n8566), .ZN(n8570) );
  AOI222_X1 U10095 ( .A1(n9883), .A2(n8570), .B1(n8569), .B2(n9880), .C1(n8568), .C2(n9878), .ZN(n8784) );
  MUX2_X1 U10096 ( .A(n8571), .B(n8784), .S(n8710), .Z(n8574) );
  AOI22_X1 U10097 ( .A1(n8786), .A2(n4350), .B1(n9905), .B2(n8572), .ZN(n8573)
         );
  OAI211_X1 U10098 ( .C1(n8789), .C2(n8699), .A(n8574), .B(n8573), .ZN(
        P2_U3207) );
  NOR2_X1 U10099 ( .A1(n8791), .A2(n8708), .ZN(n8580) );
  INV_X1 U10100 ( .A(n8575), .ZN(n8576) );
  AOI21_X1 U10101 ( .B1(n8582), .B2(n8577), .A(n8576), .ZN(n8578) );
  OAI222_X1 U10102 ( .A1(n9891), .A2(n8605), .B1(n9893), .B2(n8579), .C1(n9899), .C2(n8578), .ZN(n8790) );
  AOI211_X1 U10103 ( .C1(n9905), .C2(n8581), .A(n8580), .B(n8790), .ZN(n8586)
         );
  XNOR2_X1 U10104 ( .A(n8583), .B(n8582), .ZN(n8792) );
  INV_X1 U10105 ( .A(n8792), .ZN(n8584) );
  AOI22_X1 U10106 ( .A1(n8584), .A2(n9888), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n9910), .ZN(n8585) );
  OAI21_X1 U10107 ( .B1(n8586), .B2(n9910), .A(n8585), .ZN(P2_U3208) );
  NOR2_X1 U10108 ( .A1(n8796), .A2(n8708), .ZN(n8591) );
  XOR2_X1 U10109 ( .A(n8595), .B(n8587), .Z(n8588) );
  OAI222_X1 U10110 ( .A1(n9891), .A2(n8590), .B1(n9893), .B2(n8589), .C1(n9899), .C2(n8588), .ZN(n8795) );
  AOI211_X1 U10111 ( .C1(n9905), .C2(n8592), .A(n8591), .B(n8795), .ZN(n8599)
         );
  NAND2_X1 U10112 ( .A1(n8594), .A2(n8593), .ZN(n8596) );
  XNOR2_X1 U10113 ( .A(n8596), .B(n8595), .ZN(n8797) );
  INV_X1 U10114 ( .A(n8797), .ZN(n8597) );
  AOI22_X1 U10115 ( .A1(n8597), .A2(n9888), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9910), .ZN(n8598) );
  OAI21_X1 U10116 ( .B1(n8599), .B2(n9910), .A(n8598), .ZN(P2_U3209) );
  XNOR2_X1 U10117 ( .A(n8600), .B(n8602), .ZN(n8803) );
  INV_X1 U10118 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n8607) );
  XOR2_X1 U10119 ( .A(n8602), .B(n8601), .Z(n8603) );
  OAI222_X1 U10120 ( .A1(n9893), .A2(n8605), .B1(n9891), .B2(n8604), .C1(n9899), .C2(n8603), .ZN(n8800) );
  INV_X1 U10121 ( .A(n8800), .ZN(n8606) );
  MUX2_X1 U10122 ( .A(n8607), .B(n8606), .S(n8710), .Z(n8611) );
  AOI22_X1 U10123 ( .A1(n8609), .A2(n4350), .B1(n9905), .B2(n8608), .ZN(n8610)
         );
  OAI211_X1 U10124 ( .C1(n8803), .C2(n8699), .A(n8611), .B(n8610), .ZN(
        P2_U3210) );
  XOR2_X1 U10125 ( .A(n8615), .B(n8612), .Z(n8811) );
  INV_X1 U10126 ( .A(n8613), .ZN(n8617) );
  NAND3_X1 U10127 ( .A1(n8628), .A2(n8615), .A3(n8614), .ZN(n8616) );
  NAND2_X1 U10128 ( .A1(n8617), .A2(n8616), .ZN(n8620) );
  AOI222_X1 U10129 ( .A1(n9883), .A2(n8620), .B1(n8619), .B2(n9878), .C1(n8618), .C2(n9880), .ZN(n8806) );
  MUX2_X1 U10130 ( .A(n8621), .B(n8806), .S(n8710), .Z(n8624) );
  AOI22_X1 U10131 ( .A1(n8808), .A2(n4350), .B1(n9905), .B2(n8622), .ZN(n8623)
         );
  OAI211_X1 U10132 ( .C1(n8811), .C2(n8699), .A(n8624), .B(n8623), .ZN(
        P2_U3212) );
  XOR2_X1 U10133 ( .A(n8625), .B(n8627), .Z(n8817) );
  INV_X1 U10134 ( .A(n8626), .ZN(n8630) );
  INV_X1 U10135 ( .A(n8627), .ZN(n8629) );
  OAI21_X1 U10136 ( .B1(n8630), .B2(n8629), .A(n8628), .ZN(n8632) );
  AOI222_X1 U10137 ( .A1(n9883), .A2(n8632), .B1(n8631), .B2(n9878), .C1(n8656), .C2(n9880), .ZN(n8812) );
  MUX2_X1 U10138 ( .A(n8633), .B(n8812), .S(n8710), .Z(n8637) );
  INV_X1 U10139 ( .A(n8634), .ZN(n8635) );
  AOI22_X1 U10140 ( .A1(n8814), .A2(n4350), .B1(n9905), .B2(n8635), .ZN(n8636)
         );
  OAI211_X1 U10141 ( .C1(n8817), .C2(n8699), .A(n8637), .B(n8636), .ZN(
        P2_U3213) );
  XNOR2_X1 U10142 ( .A(n8638), .B(n8639), .ZN(n8822) );
  XNOR2_X1 U10143 ( .A(n8640), .B(n8639), .ZN(n8641) );
  OAI222_X1 U10144 ( .A1(n9891), .A2(n8643), .B1(n9893), .B2(n8642), .C1(n9899), .C2(n8641), .ZN(n8743) );
  NAND2_X1 U10145 ( .A1(n8743), .A2(n8710), .ZN(n8648) );
  OAI22_X1 U10146 ( .A1(n8710), .A2(n8645), .B1(n8644), .B2(n8706), .ZN(n8646)
         );
  AOI21_X1 U10147 ( .B1(n8744), .B2(n4350), .A(n8646), .ZN(n8647) );
  OAI211_X1 U10148 ( .C1(n8822), .C2(n8699), .A(n8648), .B(n8647), .ZN(
        P2_U3214) );
  NAND2_X1 U10149 ( .A1(n8650), .A2(n8649), .ZN(n8653) );
  NAND2_X1 U10150 ( .A1(n8652), .A2(n8651), .ZN(n8654) );
  XNOR2_X1 U10151 ( .A(n8653), .B(n8654), .ZN(n8826) );
  INV_X1 U10152 ( .A(n8826), .ZN(n8663) );
  XNOR2_X1 U10153 ( .A(n8655), .B(n8654), .ZN(n8657) );
  AOI222_X1 U10154 ( .A1(n9883), .A2(n8657), .B1(n8656), .B2(n9878), .C1(n8680), .C2(n9880), .ZN(n8823) );
  MUX2_X1 U10155 ( .A(n8658), .B(n8823), .S(n8710), .Z(n8662) );
  INV_X1 U10156 ( .A(n8659), .ZN(n8660) );
  AOI22_X1 U10157 ( .A1(n8825), .A2(n4350), .B1(n9905), .B2(n8660), .ZN(n8661)
         );
  OAI211_X1 U10158 ( .C1(n8663), .C2(n8699), .A(n8662), .B(n8661), .ZN(
        P2_U3215) );
  XNOR2_X1 U10159 ( .A(n8664), .B(n8666), .ZN(n8832) );
  INV_X1 U10160 ( .A(n8832), .ZN(n8674) );
  XOR2_X1 U10161 ( .A(n8666), .B(n8665), .Z(n8668) );
  AOI222_X1 U10162 ( .A1(n9883), .A2(n8668), .B1(n8667), .B2(n9878), .C1(n8691), .C2(n9880), .ZN(n8829) );
  MUX2_X1 U10163 ( .A(n8669), .B(n8829), .S(n8710), .Z(n8673) );
  INV_X1 U10164 ( .A(n8670), .ZN(n8671) );
  AOI22_X1 U10165 ( .A1(n8831), .A2(n4350), .B1(n9905), .B2(n8671), .ZN(n8672)
         );
  OAI211_X1 U10166 ( .C1(n8674), .C2(n8699), .A(n8673), .B(n8672), .ZN(
        P2_U3216) );
  NAND2_X1 U10167 ( .A1(n8676), .A2(n8675), .ZN(n8677) );
  XOR2_X1 U10168 ( .A(n8678), .B(n8677), .Z(n8838) );
  INV_X1 U10169 ( .A(n8838), .ZN(n8687) );
  XOR2_X1 U10170 ( .A(n8679), .B(n8678), .Z(n8681) );
  AOI222_X1 U10171 ( .A1(n9883), .A2(n8681), .B1(n8680), .B2(n9878), .C1(n8703), .C2(n9880), .ZN(n8835) );
  MUX2_X1 U10172 ( .A(n8682), .B(n8835), .S(n8710), .Z(n8686) );
  INV_X1 U10173 ( .A(n8683), .ZN(n8684) );
  AOI22_X1 U10174 ( .A1(n8837), .A2(n4350), .B1(n9905), .B2(n8684), .ZN(n8685)
         );
  OAI211_X1 U10175 ( .C1(n8687), .C2(n8699), .A(n8686), .B(n8685), .ZN(
        P2_U3217) );
  XNOR2_X1 U10176 ( .A(n8688), .B(n8689), .ZN(n8844) );
  INV_X1 U10177 ( .A(n8844), .ZN(n8700) );
  XNOR2_X1 U10178 ( .A(n8690), .B(n8689), .ZN(n8693) );
  AOI222_X1 U10179 ( .A1(n9883), .A2(n8693), .B1(n8692), .B2(n9880), .C1(n8691), .C2(n9878), .ZN(n8841) );
  MUX2_X1 U10180 ( .A(n8694), .B(n8841), .S(n8710), .Z(n8698) );
  AOI22_X1 U10181 ( .A1(n8843), .A2(n4350), .B1(n9905), .B2(n8695), .ZN(n8697)
         );
  OAI211_X1 U10182 ( .C1(n8700), .C2(n8699), .A(n8698), .B(n8697), .ZN(
        P2_U3218) );
  XNOR2_X1 U10183 ( .A(n8702), .B(n8701), .ZN(n8705) );
  AOI222_X1 U10184 ( .A1(n9883), .A2(n8705), .B1(n8704), .B2(n9880), .C1(n8703), .C2(n9878), .ZN(n8847) );
  INV_X1 U10185 ( .A(n8847), .ZN(n8712) );
  OAI22_X1 U10186 ( .A1(n8709), .A2(n8708), .B1(n8707), .B2(n8706), .ZN(n8711)
         );
  OAI21_X1 U10187 ( .B1(n8712), .B2(n8711), .A(n8710), .ZN(n8716) );
  XNOR2_X1 U10188 ( .A(n8714), .B(n8713), .ZN(n8852) );
  AOI22_X1 U10189 ( .A1(n8852), .A2(n9888), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n9910), .ZN(n8715) );
  NAND2_X1 U10190 ( .A1(n8716), .A2(n8715), .ZN(P2_U3219) );
  INV_X1 U10191 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8719) );
  NAND2_X1 U10192 ( .A1(n8766), .A2(n8761), .ZN(n8718) );
  INV_X1 U10193 ( .A(n8717), .ZN(n8767) );
  NAND2_X1 U10194 ( .A1(n8767), .A2(n9986), .ZN(n8720) );
  OAI211_X1 U10195 ( .C1(n9986), .C2(n8719), .A(n8718), .B(n8720), .ZN(
        P2_U3490) );
  NAND2_X1 U10196 ( .A1(n9984), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8721) );
  OAI211_X1 U10197 ( .C1(n8722), .C2(n8734), .A(n8721), .B(n8720), .ZN(
        P2_U3489) );
  INV_X1 U10198 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U10199 ( .A1(n8775), .A2(n8762), .ZN(n8724) );
  MUX2_X1 U10200 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8779), .S(n9986), .Z(n8726) );
  OAI22_X1 U10201 ( .A1(n8781), .A2(n8747), .B1(n8780), .B2(n8734), .ZN(n8725)
         );
  OR2_X1 U10202 ( .A1(n8726), .A2(n8725), .ZN(P2_U3486) );
  INV_X1 U10203 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n8727) );
  MUX2_X1 U10204 ( .A(n8727), .B(n8784), .S(n9986), .Z(n8729) );
  NAND2_X1 U10205 ( .A1(n8786), .A2(n8761), .ZN(n8728) );
  OAI211_X1 U10206 ( .C1(n8789), .C2(n8747), .A(n8729), .B(n8728), .ZN(
        P2_U3485) );
  MUX2_X1 U10207 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8790), .S(n9986), .Z(n8731) );
  OAI22_X1 U10208 ( .A1(n8792), .A2(n8747), .B1(n8791), .B2(n8734), .ZN(n8730)
         );
  OR2_X1 U10209 ( .A1(n8731), .A2(n8730), .ZN(P2_U3484) );
  MUX2_X1 U10210 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8795), .S(n9986), .Z(n8733) );
  OAI22_X1 U10211 ( .A1(n8797), .A2(n8747), .B1(n8796), .B2(n8734), .ZN(n8732)
         );
  OR2_X1 U10212 ( .A1(n8733), .A2(n8732), .ZN(P2_U3483) );
  MUX2_X1 U10213 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8800), .S(n9986), .Z(n8736) );
  OAI22_X1 U10214 ( .A1(n8803), .A2(n8747), .B1(n8802), .B2(n8734), .ZN(n8735)
         );
  OR2_X1 U10215 ( .A1(n8736), .A2(n8735), .ZN(P2_U3482) );
  MUX2_X1 U10216 ( .A(n8737), .B(n8806), .S(n9986), .Z(n8739) );
  NAND2_X1 U10217 ( .A1(n8808), .A2(n8761), .ZN(n8738) );
  OAI211_X1 U10218 ( .C1(n8747), .C2(n8811), .A(n8739), .B(n8738), .ZN(
        P2_U3480) );
  MUX2_X1 U10219 ( .A(n8740), .B(n8812), .S(n9986), .Z(n8742) );
  NAND2_X1 U10220 ( .A1(n8814), .A2(n8761), .ZN(n8741) );
  OAI211_X1 U10221 ( .C1(n8747), .C2(n8817), .A(n8742), .B(n8741), .ZN(
        P2_U3479) );
  AOI21_X1 U10222 ( .B1(n9967), .B2(n8744), .A(n8743), .ZN(n8818) );
  MUX2_X1 U10223 ( .A(n8745), .B(n8818), .S(n9986), .Z(n8746) );
  OAI21_X1 U10224 ( .B1(n8747), .B2(n8822), .A(n8746), .ZN(P2_U3478) );
  MUX2_X1 U10225 ( .A(n8748), .B(n8823), .S(n9986), .Z(n8750) );
  AOI22_X1 U10226 ( .A1(n8826), .A2(n8762), .B1(n8761), .B2(n8825), .ZN(n8749)
         );
  NAND2_X1 U10227 ( .A1(n8750), .A2(n8749), .ZN(P2_U3477) );
  MUX2_X1 U10228 ( .A(n8751), .B(n8829), .S(n9986), .Z(n8753) );
  AOI22_X1 U10229 ( .A1(n8832), .A2(n8762), .B1(n8761), .B2(n8831), .ZN(n8752)
         );
  NAND2_X1 U10230 ( .A1(n8753), .A2(n8752), .ZN(P2_U3476) );
  MUX2_X1 U10231 ( .A(n8754), .B(n8835), .S(n9986), .Z(n8756) );
  AOI22_X1 U10232 ( .A1(n8838), .A2(n8762), .B1(n8761), .B2(n8837), .ZN(n8755)
         );
  NAND2_X1 U10233 ( .A1(n8756), .A2(n8755), .ZN(P2_U3475) );
  MUX2_X1 U10234 ( .A(n8757), .B(n8841), .S(n9986), .Z(n8759) );
  AOI22_X1 U10235 ( .A1(n8844), .A2(n8762), .B1(n8761), .B2(n8843), .ZN(n8758)
         );
  NAND2_X1 U10236 ( .A1(n8759), .A2(n8758), .ZN(P2_U3474) );
  MUX2_X1 U10237 ( .A(n8760), .B(n8847), .S(n9986), .Z(n8764) );
  AOI22_X1 U10238 ( .A1(n8852), .A2(n8762), .B1(n8761), .B2(n8849), .ZN(n8763)
         );
  NAND2_X1 U10239 ( .A1(n8764), .A2(n8763), .ZN(P2_U3473) );
  MUX2_X1 U10240 ( .A(P2_REG1_REG_0__SCAN_IN), .B(n8765), .S(n9986), .Z(
        P2_U3459) );
  NAND2_X1 U10241 ( .A1(n8766), .A2(n8850), .ZN(n8768) );
  NAND2_X1 U10242 ( .A1(n8767), .A2(n9968), .ZN(n8770) );
  OAI211_X1 U10243 ( .C1(n7000), .C2(n9968), .A(n8768), .B(n8770), .ZN(
        P2_U3458) );
  INV_X1 U10244 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8772) );
  NAND2_X1 U10245 ( .A1(n8769), .A2(n8850), .ZN(n8771) );
  OAI211_X1 U10246 ( .C1(n8772), .C2(n9968), .A(n8771), .B(n8770), .ZN(
        P2_U3457) );
  INV_X1 U10247 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n8774) );
  MUX2_X1 U10248 ( .A(n8774), .B(n8773), .S(n9968), .Z(n8777) );
  NAND2_X1 U10249 ( .A1(n8775), .A2(n8851), .ZN(n8776) );
  OAI211_X1 U10250 ( .C1(n8778), .C2(n8801), .A(n8777), .B(n8776), .ZN(
        P2_U3455) );
  MUX2_X1 U10251 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8779), .S(n9968), .Z(n8783) );
  OAI22_X1 U10252 ( .A1(n8781), .A2(n8821), .B1(n8780), .B2(n8801), .ZN(n8782)
         );
  OR2_X1 U10253 ( .A1(n8783), .A2(n8782), .ZN(P2_U3454) );
  INV_X1 U10254 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n8785) );
  MUX2_X1 U10255 ( .A(n8785), .B(n8784), .S(n9968), .Z(n8788) );
  NAND2_X1 U10256 ( .A1(n8786), .A2(n8850), .ZN(n8787) );
  OAI211_X1 U10257 ( .C1(n8789), .C2(n8821), .A(n8788), .B(n8787), .ZN(
        P2_U3453) );
  MUX2_X1 U10258 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8790), .S(n9968), .Z(n8794) );
  OAI22_X1 U10259 ( .A1(n8792), .A2(n8821), .B1(n8791), .B2(n8801), .ZN(n8793)
         );
  OR2_X1 U10260 ( .A1(n8794), .A2(n8793), .ZN(P2_U3452) );
  MUX2_X1 U10261 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8795), .S(n9968), .Z(n8799) );
  OAI22_X1 U10262 ( .A1(n8797), .A2(n8821), .B1(n8796), .B2(n8801), .ZN(n8798)
         );
  OR2_X1 U10263 ( .A1(n8799), .A2(n8798), .ZN(P2_U3451) );
  MUX2_X1 U10264 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8800), .S(n9968), .Z(n8805) );
  OAI22_X1 U10265 ( .A1(n8803), .A2(n8821), .B1(n8802), .B2(n8801), .ZN(n8804)
         );
  OR2_X1 U10266 ( .A1(n8805), .A2(n8804), .ZN(P2_U3450) );
  MUX2_X1 U10267 ( .A(n8807), .B(n8806), .S(n9968), .Z(n8810) );
  NAND2_X1 U10268 ( .A1(n8808), .A2(n8850), .ZN(n8809) );
  OAI211_X1 U10269 ( .C1(n8811), .C2(n8821), .A(n8810), .B(n8809), .ZN(
        P2_U3448) );
  INV_X1 U10270 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n8813) );
  MUX2_X1 U10271 ( .A(n8813), .B(n8812), .S(n9968), .Z(n8816) );
  NAND2_X1 U10272 ( .A1(n8814), .A2(n8850), .ZN(n8815) );
  OAI211_X1 U10273 ( .C1(n8817), .C2(n8821), .A(n8816), .B(n8815), .ZN(
        P2_U3447) );
  INV_X1 U10274 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n8819) );
  MUX2_X1 U10275 ( .A(n8819), .B(n8818), .S(n9968), .Z(n8820) );
  OAI21_X1 U10276 ( .B1(n8822), .B2(n8821), .A(n8820), .ZN(P2_U3446) );
  INV_X1 U10277 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n8824) );
  MUX2_X1 U10278 ( .A(n8824), .B(n8823), .S(n9968), .Z(n8828) );
  AOI22_X1 U10279 ( .A1(n8826), .A2(n8851), .B1(n8850), .B2(n8825), .ZN(n8827)
         );
  NAND2_X1 U10280 ( .A1(n8828), .A2(n8827), .ZN(P2_U3444) );
  INV_X1 U10281 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8830) );
  MUX2_X1 U10282 ( .A(n8830), .B(n8829), .S(n9968), .Z(n8834) );
  AOI22_X1 U10283 ( .A1(n8832), .A2(n8851), .B1(n8850), .B2(n8831), .ZN(n8833)
         );
  NAND2_X1 U10284 ( .A1(n8834), .A2(n8833), .ZN(P2_U3441) );
  INV_X1 U10285 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n8836) );
  MUX2_X1 U10286 ( .A(n8836), .B(n8835), .S(n9968), .Z(n8840) );
  AOI22_X1 U10287 ( .A1(n8838), .A2(n8851), .B1(n8850), .B2(n8837), .ZN(n8839)
         );
  NAND2_X1 U10288 ( .A1(n8840), .A2(n8839), .ZN(P2_U3438) );
  INV_X1 U10289 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8842) );
  MUX2_X1 U10290 ( .A(n8842), .B(n8841), .S(n9968), .Z(n8846) );
  AOI22_X1 U10291 ( .A1(n8844), .A2(n8851), .B1(n8850), .B2(n8843), .ZN(n8845)
         );
  NAND2_X1 U10292 ( .A1(n8846), .A2(n8845), .ZN(P2_U3435) );
  INV_X1 U10293 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n8848) );
  MUX2_X1 U10294 ( .A(n8848), .B(n8847), .S(n9968), .Z(n8854) );
  AOI22_X1 U10295 ( .A1(n8852), .A2(n8851), .B1(n8850), .B2(n8849), .ZN(n8853)
         );
  NAND2_X1 U10296 ( .A1(n8854), .A2(n8853), .ZN(P2_U3432) );
  OAI222_X1 U10297 ( .A1(n8860), .A2(n8859), .B1(n8858), .B2(n8857), .C1(n8856), .C2(P2_U3151), .ZN(P2_U3268) );
  MUX2_X1 U10298 ( .A(n8861), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3295) );
  NAND2_X1 U10299 ( .A1(n8864), .A2(n9016), .ZN(n8871) );
  NAND2_X1 U10300 ( .A1(n9018), .A2(n9032), .ZN(n8866) );
  OAI211_X1 U10301 ( .C1(n8867), .C2(n8988), .A(n8866), .B(n8865), .ZN(n8868)
         );
  AOI21_X1 U10302 ( .B1(n8869), .B2(n9022), .A(n8868), .ZN(n8870) );
  OAI211_X1 U10303 ( .C1(n8872), .C2(n9026), .A(n8871), .B(n8870), .ZN(
        P1_U3215) );
  NOR2_X1 U10304 ( .A1(n4823), .A2(n8874), .ZN(n8875) );
  XNOR2_X1 U10305 ( .A(n8876), .B(n8875), .ZN(n8883) );
  OAI22_X1 U10306 ( .A1(n9417), .A2(n8988), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8877), .ZN(n8878) );
  AOI21_X1 U10307 ( .B1(n9414), .B2(n9018), .A(n8878), .ZN(n8881) );
  INV_X1 U10308 ( .A(n8879), .ZN(n9255) );
  NAND2_X1 U10309 ( .A1(n9022), .A2(n9255), .ZN(n8880) );
  OAI211_X1 U10310 ( .C1(n9507), .C2(n9026), .A(n8881), .B(n8880), .ZN(n8882)
         );
  AOI21_X1 U10311 ( .B1(n8883), .B2(n9016), .A(n8882), .ZN(n8884) );
  INV_X1 U10312 ( .A(n8884), .ZN(P1_U3216) );
  OAI21_X1 U10313 ( .B1(n8886), .B2(n8885), .A(n6872), .ZN(n8887) );
  NAND2_X1 U10314 ( .A1(n8887), .A2(n9016), .ZN(n8897) );
  NAND2_X1 U10315 ( .A1(P1_U3086), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9079) );
  INV_X1 U10316 ( .A(n9079), .ZN(n8888) );
  AOI21_X1 U10317 ( .B1(n8889), .B2(n9043), .A(n8888), .ZN(n8896) );
  OAI22_X1 U10318 ( .A1(n9026), .A2(n8891), .B1(n8890), .B2(n9008), .ZN(n8892)
         );
  INV_X1 U10319 ( .A(n8892), .ZN(n8895) );
  NAND2_X1 U10320 ( .A1(n9022), .A2(n8893), .ZN(n8894) );
  NAND4_X1 U10321 ( .A1(n8897), .A2(n8896), .A3(n8895), .A4(n8894), .ZN(
        P1_U3218) );
  INV_X1 U10322 ( .A(n9453), .ZN(n9321) );
  OAI21_X1 U10323 ( .B1(n8900), .B2(n8898), .A(n8899), .ZN(n8901) );
  NAND2_X1 U10324 ( .A1(n8901), .A2(n9016), .ZN(n8906) );
  OAI21_X1 U10325 ( .B1(n8988), .B2(n9357), .A(n8902), .ZN(n8904) );
  INV_X1 U10326 ( .A(n9022), .ZN(n8954) );
  NOR2_X1 U10327 ( .A1(n8954), .A2(n9317), .ZN(n8903) );
  AOI211_X1 U10328 ( .C1(n9018), .C2(n9432), .A(n8904), .B(n8903), .ZN(n8905)
         );
  OAI211_X1 U10329 ( .C1(n9321), .C2(n9026), .A(n8906), .B(n8905), .ZN(
        P1_U3219) );
  OAI21_X1 U10330 ( .B1(n8909), .B2(n8908), .A(n8907), .ZN(n8910) );
  NAND2_X1 U10331 ( .A1(n8910), .A2(n9016), .ZN(n8915) );
  INV_X1 U10332 ( .A(n8911), .ZN(n9283) );
  AOI22_X1 U10333 ( .A1(n9433), .A2(n9018), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3086), .ZN(n8912) );
  OAI21_X1 U10334 ( .B1(n9316), .B2(n8988), .A(n8912), .ZN(n8913) );
  AOI21_X1 U10335 ( .B1(n9283), .B2(n9022), .A(n8913), .ZN(n8914) );
  OAI211_X1 U10336 ( .C1(n4684), .C2(n9026), .A(n8915), .B(n8914), .ZN(
        P1_U3223) );
  AOI21_X1 U10337 ( .B1(n4425), .B2(n8916), .A(n9004), .ZN(n8922) );
  OAI22_X1 U10338 ( .A1(n9258), .A2(n8988), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8917), .ZN(n8918) );
  AOI21_X1 U10339 ( .B1(n9194), .B2(n9018), .A(n8918), .ZN(n8919) );
  OAI21_X1 U10340 ( .B1(n8954), .B2(n9226), .A(n8919), .ZN(n8920) );
  AOI21_X1 U10341 ( .B1(n9231), .B2(n8958), .A(n8920), .ZN(n8921) );
  OAI21_X1 U10342 ( .B1(n8922), .B2(n8960), .A(n8921), .ZN(P1_U3225) );
  INV_X1 U10343 ( .A(n8923), .ZN(n8925) );
  NOR2_X1 U10344 ( .A1(n8925), .A2(n8924), .ZN(n8926) );
  AOI21_X1 U10345 ( .B1(n8925), .B2(n8924), .A(n8926), .ZN(n9014) );
  NAND2_X1 U10346 ( .A1(n9014), .A2(n9015), .ZN(n9013) );
  INV_X1 U10347 ( .A(n8926), .ZN(n8927) );
  NAND2_X1 U10348 ( .A1(n9013), .A2(n8927), .ZN(n8931) );
  NAND2_X1 U10349 ( .A1(n8929), .A2(n8928), .ZN(n8930) );
  XNOR2_X1 U10350 ( .A(n8931), .B(n8930), .ZN(n8940) );
  NAND2_X1 U10351 ( .A1(n9018), .A2(n9030), .ZN(n8933) );
  OAI211_X1 U10352 ( .C1(n8934), .C2(n8988), .A(n8933), .B(n8932), .ZN(n8937)
         );
  NOR2_X1 U10353 ( .A1(n8935), .A2(n9026), .ZN(n8936) );
  AOI211_X1 U10354 ( .C1(n8938), .C2(n9022), .A(n8937), .B(n8936), .ZN(n8939)
         );
  OAI21_X1 U10355 ( .B1(n8940), .B2(n8960), .A(n8939), .ZN(P1_U3226) );
  XNOR2_X1 U10356 ( .A(n8943), .B(n8942), .ZN(n8944) );
  XNOR2_X1 U10357 ( .A(n8941), .B(n8944), .ZN(n8950) );
  OAI21_X1 U10358 ( .B1(n8988), .B2(n9356), .A(n8945), .ZN(n8946) );
  AOI21_X1 U10359 ( .B1(n9018), .B2(n9313), .A(n8946), .ZN(n8947) );
  OAI21_X1 U10360 ( .B1(n8954), .B2(n9350), .A(n8947), .ZN(n8948) );
  AOI21_X1 U10361 ( .B1(n9463), .B2(n8958), .A(n8948), .ZN(n8949) );
  OAI21_X1 U10362 ( .B1(n8950), .B2(n8960), .A(n8949), .ZN(P1_U3228) );
  AOI21_X1 U10363 ( .B1(n8953), .B2(n8952), .A(n8951), .ZN(n8961) );
  NOR2_X1 U10364 ( .A1(n8954), .A2(n9244), .ZN(n8957) );
  AOI22_X1 U10365 ( .A1(n9211), .A2(n9018), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3086), .ZN(n8955) );
  OAI21_X1 U10366 ( .B1(n9270), .B2(n8988), .A(n8955), .ZN(n8956) );
  AOI211_X1 U10367 ( .C1(n9243), .C2(n8958), .A(n8957), .B(n8956), .ZN(n8959)
         );
  OAI21_X1 U10368 ( .B1(n8961), .B2(n8960), .A(n8959), .ZN(P1_U3229) );
  AND2_X1 U10369 ( .A1(n6872), .A2(n8962), .ZN(n8965) );
  OAI211_X1 U10370 ( .C1(n8965), .C2(n8964), .A(n9016), .B(n8963), .ZN(n8971)
         );
  AND2_X1 U10371 ( .A1(P1_U3086), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9092) );
  AOI21_X1 U10372 ( .B1(n9018), .B2(n9040), .A(n9092), .ZN(n8970) );
  OAI22_X1 U10373 ( .A1(n9026), .A2(n9615), .B1(n8966), .B2(n8988), .ZN(n8967)
         );
  INV_X1 U10374 ( .A(n8967), .ZN(n8969) );
  NAND2_X1 U10375 ( .A1(n9022), .A2(n9611), .ZN(n8968) );
  NAND4_X1 U10376 ( .A1(n8971), .A2(n8970), .A3(n8969), .A4(n8968), .ZN(
        P1_U3230) );
  NOR2_X1 U10377 ( .A1(n4375), .A2(n8972), .ZN(n8973) );
  XNOR2_X1 U10378 ( .A(n8974), .B(n8973), .ZN(n8975) );
  NAND2_X1 U10379 ( .A1(n8975), .A2(n9016), .ZN(n8980) );
  OAI22_X1 U10380 ( .A1(n8988), .A2(n9330), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8976), .ZN(n8978) );
  NOR2_X1 U10381 ( .A1(n9301), .A2(n9008), .ZN(n8977) );
  AOI211_X1 U10382 ( .C1(n9297), .C2(n9022), .A(n8978), .B(n8977), .ZN(n8979)
         );
  OAI211_X1 U10383 ( .C1(n9445), .C2(n9026), .A(n8980), .B(n8979), .ZN(
        P1_U3233) );
  INV_X1 U10384 ( .A(n8981), .ZN(n8983) );
  NAND2_X1 U10385 ( .A1(n8983), .A2(n8982), .ZN(n8985) );
  XNOR2_X1 U10386 ( .A(n8985), .B(n8984), .ZN(n8986) );
  NAND2_X1 U10387 ( .A1(n8986), .A2(n9016), .ZN(n8992) );
  OAI22_X1 U10388 ( .A1(n9301), .A2(n8988), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8987), .ZN(n8990) );
  NOR2_X1 U10389 ( .A1(n9270), .A2(n9008), .ZN(n8989) );
  AOI211_X1 U10390 ( .C1(n9267), .C2(n9022), .A(n8990), .B(n8989), .ZN(n8991)
         );
  OAI211_X1 U10391 ( .C1(n9426), .C2(n9026), .A(n8992), .B(n8991), .ZN(
        P1_U3235) );
  OAI21_X1 U10392 ( .B1(n8995), .B2(n8994), .A(n8993), .ZN(n8996) );
  NAND2_X1 U10393 ( .A1(n8996), .A2(n9016), .ZN(n9000) );
  NAND2_X1 U10394 ( .A1(n9018), .A2(n9440), .ZN(n8997) );
  NAND2_X1 U10395 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9150) );
  OAI211_X1 U10396 ( .C1(n9329), .C2(n8988), .A(n8997), .B(n9150), .ZN(n8998)
         );
  AOI21_X1 U10397 ( .B1(n9338), .B2(n9022), .A(n8998), .ZN(n8999) );
  OAI211_X1 U10398 ( .C1(n9516), .C2(n9026), .A(n9000), .B(n8999), .ZN(
        P1_U3238) );
  OAI21_X1 U10399 ( .B1(n9004), .B2(n9003), .A(n9002), .ZN(n9005) );
  NAND3_X1 U10400 ( .A1(n9006), .A2(n9016), .A3(n9005), .ZN(n9012) );
  OAI22_X1 U10401 ( .A1(n9390), .A2(n8988), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9007), .ZN(n9010) );
  NOR2_X1 U10402 ( .A1(n9391), .A2(n9008), .ZN(n9009) );
  AOI211_X1 U10403 ( .C1(n9210), .C2(n9022), .A(n9010), .B(n9009), .ZN(n9011)
         );
  OAI211_X1 U10404 ( .C1(n9495), .C2(n9026), .A(n9012), .B(n9011), .ZN(
        P1_U3240) );
  OAI21_X1 U10405 ( .B1(n9015), .B2(n9014), .A(n9013), .ZN(n9017) );
  NAND2_X1 U10406 ( .A1(n9017), .A2(n9016), .ZN(n9025) );
  NAND2_X1 U10407 ( .A1(n9018), .A2(n9031), .ZN(n9020) );
  OAI211_X1 U10408 ( .C1(n9671), .C2(n8988), .A(n9020), .B(n9019), .ZN(n9021)
         );
  AOI21_X1 U10409 ( .B1(n9023), .B2(n9022), .A(n9021), .ZN(n9024) );
  OAI211_X1 U10410 ( .C1(n9027), .C2(n9026), .A(n9025), .B(n9024), .ZN(
        P1_U3241) );
  MUX2_X1 U10411 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n4458), .S(P1_U3973), .Z(
        P1_U3583) );
  MUX2_X1 U10412 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9028), .S(P1_U3973), .Z(
        P1_U3582) );
  MUX2_X1 U10413 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9029), .S(P1_U3973), .Z(
        P1_U3581) );
  MUX2_X1 U10414 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9194), .S(P1_U3973), .Z(
        P1_U3580) );
  MUX2_X1 U10415 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9211), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10416 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9414), .S(P1_U3973), .Z(
        P1_U3578) );
  MUX2_X1 U10417 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9424), .S(P1_U3973), .Z(
        P1_U3577) );
  MUX2_X1 U10418 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9433), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10419 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9442), .S(P1_U3973), .Z(
        P1_U3575) );
  MUX2_X1 U10420 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9432), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10421 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9440), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10422 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9313), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10423 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9030), .S(P1_U3973), .Z(
        P1_U3571) );
  MUX2_X1 U10424 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9031), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10425 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9032), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10426 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9033), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10427 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9034), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10428 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9035), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10429 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9036), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10430 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9037), .S(P1_U3973), .Z(
        P1_U3564) );
  MUX2_X1 U10431 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9038), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10432 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9646), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10433 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9039), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10434 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9040), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10435 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9041), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10436 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9042), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10437 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9043), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10438 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9044), .S(P1_U3973), .Z(
        P1_U3555) );
  MUX2_X1 U10439 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9045), .S(P1_U3973), .Z(
        P1_U3554) );
  INV_X1 U10440 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9047) );
  OAI22_X1 U10441 ( .A1(n9590), .A2(n9047), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9046), .ZN(n9048) );
  AOI21_X1 U10442 ( .B1(n9564), .B2(n9049), .A(n9048), .ZN(n9057) );
  OAI211_X1 U10443 ( .C1(n9051), .C2(n9059), .A(n9580), .B(n9050), .ZN(n9056)
         );
  OAI211_X1 U10444 ( .C1(n9054), .C2(n9053), .A(n9575), .B(n9052), .ZN(n9055)
         );
  NAND3_X1 U10445 ( .A1(n9057), .A2(n9056), .A3(n9055), .ZN(P1_U3244) );
  MUX2_X1 U10446 ( .A(n9060), .B(n9059), .S(n9058), .Z(n9062) );
  INV_X1 U10447 ( .A(n4353), .ZN(n9061) );
  NAND2_X1 U10448 ( .A1(n9062), .A2(n9061), .ZN(n9064) );
  OAI211_X1 U10449 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n9065), .A(n9064), .B(
        P1_U3973), .ZN(n9106) );
  INV_X1 U10450 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9067) );
  OAI22_X1 U10451 ( .A1(n9590), .A2(n9067), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9066), .ZN(n9068) );
  AOI21_X1 U10452 ( .B1(n9564), .B2(n9069), .A(n9068), .ZN(n9078) );
  OAI211_X1 U10453 ( .C1(n9072), .C2(n9071), .A(n9575), .B(n9070), .ZN(n9077)
         );
  OAI211_X1 U10454 ( .C1(n9075), .C2(n9074), .A(n9580), .B(n9073), .ZN(n9076)
         );
  NAND4_X1 U10455 ( .A1(n9106), .A2(n9078), .A3(n9077), .A4(n9076), .ZN(
        P1_U3245) );
  INV_X1 U10456 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9080) );
  OAI21_X1 U10457 ( .B1(n9590), .B2(n9080), .A(n9079), .ZN(n9081) );
  AOI21_X1 U10458 ( .B1(n9564), .B2(n9082), .A(n9081), .ZN(n9091) );
  OAI211_X1 U10459 ( .C1(n9085), .C2(n9084), .A(n9575), .B(n9083), .ZN(n9090)
         );
  OAI211_X1 U10460 ( .C1(n9088), .C2(n9087), .A(n9580), .B(n9086), .ZN(n9089)
         );
  NAND3_X1 U10461 ( .A1(n9091), .A2(n9090), .A3(n9089), .ZN(P1_U3246) );
  INV_X1 U10462 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9094) );
  INV_X1 U10463 ( .A(n9092), .ZN(n9093) );
  OAI21_X1 U10464 ( .B1(n9590), .B2(n9094), .A(n9093), .ZN(n9095) );
  AOI21_X1 U10465 ( .B1(n9564), .B2(n9096), .A(n9095), .ZN(n9105) );
  OAI211_X1 U10466 ( .C1(n9099), .C2(n9098), .A(n9580), .B(n9097), .ZN(n9104)
         );
  OAI211_X1 U10467 ( .C1(n9102), .C2(n9101), .A(n9575), .B(n9100), .ZN(n9103)
         );
  NAND4_X1 U10468 ( .A1(n9106), .A2(n9105), .A3(n9104), .A4(n9103), .ZN(
        P1_U3247) );
  INV_X1 U10469 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n9108) );
  OAI21_X1 U10470 ( .B1(n9590), .B2(n9108), .A(n9107), .ZN(n9109) );
  AOI21_X1 U10471 ( .B1(n9564), .B2(n9110), .A(n9109), .ZN(n9119) );
  OAI211_X1 U10472 ( .C1(n9113), .C2(n9112), .A(n9575), .B(n9111), .ZN(n9118)
         );
  OAI211_X1 U10473 ( .C1(n9116), .C2(n9115), .A(n9580), .B(n9114), .ZN(n9117)
         );
  NAND3_X1 U10474 ( .A1(n9119), .A2(n9118), .A3(n9117), .ZN(P1_U3248) );
  INV_X1 U10475 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n9121) );
  OAI21_X1 U10476 ( .B1(n9590), .B2(n9121), .A(n9120), .ZN(n9122) );
  AOI21_X1 U10477 ( .B1(n9564), .B2(n9123), .A(n9122), .ZN(n9132) );
  OAI211_X1 U10478 ( .C1(n9126), .C2(n9125), .A(n9575), .B(n9124), .ZN(n9131)
         );
  OAI211_X1 U10479 ( .C1(n9129), .C2(n9128), .A(n9580), .B(n9127), .ZN(n9130)
         );
  NAND3_X1 U10480 ( .A1(n9132), .A2(n9131), .A3(n9130), .ZN(P1_U3250) );
  OAI21_X1 U10481 ( .B1(n9135), .B2(n9134), .A(n9133), .ZN(n9136) );
  NAND2_X1 U10482 ( .A1(n9136), .A2(n9580), .ZN(n9146) );
  OAI21_X1 U10483 ( .B1(n9139), .B2(n9138), .A(n9137), .ZN(n9140) );
  NAND2_X1 U10484 ( .A1(n9140), .A2(n9575), .ZN(n9145) );
  AOI21_X1 U10485 ( .B1(n9154), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n9141), .ZN(
        n9144) );
  NAND2_X1 U10486 ( .A1(n9564), .A2(n9142), .ZN(n9143) );
  NAND4_X1 U10487 ( .A1(n9146), .A2(n9145), .A3(n9144), .A4(n9143), .ZN(
        P1_U3252) );
  OAI211_X1 U10488 ( .C1(n9149), .C2(n9148), .A(n9147), .B(n9580), .ZN(n9160)
         );
  INV_X1 U10489 ( .A(n9150), .ZN(n9153) );
  NOR2_X1 U10490 ( .A1(n9584), .A2(n9151), .ZN(n9152) );
  AOI211_X1 U10491 ( .C1(n9154), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9153), .B(
        n9152), .ZN(n9159) );
  OAI211_X1 U10492 ( .C1(n9157), .C2(n9156), .A(n9155), .B(n9575), .ZN(n9158)
         );
  NAND3_X1 U10493 ( .A1(n9160), .A2(n9159), .A3(n9158), .ZN(P1_U3261) );
  NAND2_X1 U10494 ( .A1(n9365), .A2(n9161), .ZN(n9166) );
  INV_X1 U10495 ( .A(n9368), .ZN(n9164) );
  NOR2_X1 U10496 ( .A1(n4352), .A2(n9164), .ZN(n9169) );
  AOI21_X1 U10497 ( .B1(n4352), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9169), .ZN(
        n9165) );
  OAI211_X1 U10498 ( .C1(n9482), .C2(n9614), .A(n9166), .B(n9165), .ZN(
        P1_U3263) );
  XNOR2_X1 U10499 ( .A(n9167), .B(n9173), .ZN(n9168) );
  INV_X1 U10500 ( .A(n9369), .ZN(n9175) );
  INV_X1 U10501 ( .A(n9169), .ZN(n9170) );
  OAI21_X1 U10502 ( .B1(n9342), .B2(n9171), .A(n9170), .ZN(n9172) );
  AOI21_X1 U10503 ( .B1(n9173), .B2(n9600), .A(n9172), .ZN(n9174) );
  OAI21_X1 U10504 ( .B1(n9175), .B2(n9305), .A(n9174), .ZN(P1_U3264) );
  XNOR2_X1 U10505 ( .A(n9176), .B(n9185), .ZN(n9376) );
  OAI211_X1 U10506 ( .C1(n9487), .C2(n9192), .A(n9603), .B(n9177), .ZN(n9375)
         );
  AOI22_X1 U10507 ( .A1(n9178), .A2(n9610), .B1(P1_REG2_REG_28__SCAN_IN), .B2(
        n4352), .ZN(n9180) );
  OR2_X1 U10508 ( .A1(n9372), .A2(n9300), .ZN(n9179) );
  OAI211_X1 U10509 ( .C1(n9391), .C2(n9181), .A(n9180), .B(n9179), .ZN(n9182)
         );
  AOI21_X1 U10510 ( .B1(n9183), .B2(n9600), .A(n9182), .ZN(n9184) );
  OAI21_X1 U10511 ( .B1(n9375), .B2(n9305), .A(n9184), .ZN(n9189) );
  NOR2_X1 U10512 ( .A1(n9379), .A2(n9364), .ZN(n9188) );
  AOI211_X1 U10513 ( .C1(n9307), .C2(n9376), .A(n9189), .B(n9188), .ZN(n9190)
         );
  INV_X1 U10514 ( .A(n9190), .ZN(P1_U3265) );
  XNOR2_X1 U10515 ( .A(n9191), .B(n9200), .ZN(n9386) );
  AOI211_X1 U10516 ( .C1(n9193), .C2(n9207), .A(n9348), .B(n9192), .ZN(n9382)
         );
  NOR2_X1 U10517 ( .A1(n9491), .A2(n9614), .ZN(n9199) );
  AOI22_X1 U10518 ( .A1(n9194), .A2(n9296), .B1(n4352), .B2(
        P1_REG2_REG_27__SCAN_IN), .ZN(n9197) );
  NAND2_X1 U10519 ( .A1(n9195), .A2(n9610), .ZN(n9196) );
  OAI211_X1 U10520 ( .C1(n9381), .C2(n9300), .A(n9197), .B(n9196), .ZN(n9198)
         );
  AOI211_X1 U10521 ( .C1(n9382), .C2(n9608), .A(n9199), .B(n9198), .ZN(n9205)
         );
  NAND3_X1 U10522 ( .A1(n9216), .A2(n9201), .A3(n9200), .ZN(n9202) );
  NAND2_X1 U10523 ( .A1(n9203), .A2(n9202), .ZN(n9384) );
  NAND2_X1 U10524 ( .A1(n9384), .A2(n9307), .ZN(n9204) );
  OAI211_X1 U10525 ( .C1(n9386), .C2(n9364), .A(n9205), .B(n9204), .ZN(
        P1_U3266) );
  XNOR2_X1 U10526 ( .A(n9206), .B(n9217), .ZN(n9396) );
  INV_X1 U10527 ( .A(n9207), .ZN(n9208) );
  AOI211_X1 U10528 ( .C1(n9209), .C2(n9225), .A(n9348), .B(n9208), .ZN(n9392)
         );
  NOR2_X1 U10529 ( .A1(n9495), .A2(n9614), .ZN(n9215) );
  AOI22_X1 U10530 ( .A1(n9210), .A2(n9610), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n4352), .ZN(n9213) );
  NAND2_X1 U10531 ( .A1(n9211), .A2(n9296), .ZN(n9212) );
  OAI211_X1 U10532 ( .C1(n9391), .C2(n9300), .A(n9213), .B(n9212), .ZN(n9214)
         );
  AOI211_X1 U10533 ( .C1(n9392), .C2(n9608), .A(n9215), .B(n9214), .ZN(n9220)
         );
  OAI21_X1 U10534 ( .B1(n9218), .B2(n9217), .A(n9216), .ZN(n9394) );
  NAND2_X1 U10535 ( .A1(n9394), .A2(n9307), .ZN(n9219) );
  OAI211_X1 U10536 ( .C1(n9396), .C2(n9364), .A(n9220), .B(n9219), .ZN(
        P1_U3267) );
  XNOR2_X1 U10537 ( .A(n9221), .B(n9222), .ZN(n9403) );
  OAI21_X1 U10538 ( .B1(n4396), .B2(n9224), .A(n9223), .ZN(n9406) );
  OAI211_X1 U10539 ( .C1(n9499), .C2(n4376), .A(n9603), .B(n9225), .ZN(n9401)
         );
  INV_X1 U10540 ( .A(n9226), .ZN(n9227) );
  AOI22_X1 U10541 ( .A1(n9227), .A2(n9610), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n4352), .ZN(n9229) );
  NAND2_X1 U10542 ( .A1(n9414), .A2(n9296), .ZN(n9228) );
  OAI211_X1 U10543 ( .C1(n9402), .C2(n9300), .A(n9229), .B(n9228), .ZN(n9230)
         );
  AOI21_X1 U10544 ( .B1(n9231), .B2(n9600), .A(n9230), .ZN(n9232) );
  OAI21_X1 U10545 ( .B1(n9401), .B2(n9305), .A(n9232), .ZN(n9233) );
  AOI21_X1 U10546 ( .B1(n9406), .B2(n9307), .A(n9233), .ZN(n9234) );
  OAI21_X1 U10547 ( .B1(n9403), .B2(n9364), .A(n9234), .ZN(P1_U3268) );
  XNOR2_X1 U10548 ( .A(n9235), .B(n9236), .ZN(n9411) );
  INV_X1 U10549 ( .A(n9411), .ZN(n9250) );
  NAND2_X1 U10550 ( .A1(n9237), .A2(n9236), .ZN(n9238) );
  NAND3_X1 U10551 ( .A1(n9239), .A2(n9447), .A3(n9238), .ZN(n9242) );
  OAI22_X1 U10552 ( .A1(n9390), .A2(n9670), .B1(n9270), .B2(n9672), .ZN(n9240)
         );
  INV_X1 U10553 ( .A(n9240), .ZN(n9241) );
  NAND2_X1 U10554 ( .A1(n9242), .A2(n9241), .ZN(n9409) );
  AOI211_X1 U10555 ( .C1(n9243), .C2(n9254), .A(n9348), .B(n4376), .ZN(n9410)
         );
  NAND2_X1 U10556 ( .A1(n9410), .A2(n9608), .ZN(n9247) );
  INV_X1 U10557 ( .A(n9244), .ZN(n9245) );
  AOI22_X1 U10558 ( .A1(n9245), .A2(n9610), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n4352), .ZN(n9246) );
  OAI211_X1 U10559 ( .C1(n9503), .C2(n9614), .A(n9247), .B(n9246), .ZN(n9248)
         );
  AOI21_X1 U10560 ( .B1(n9342), .B2(n9409), .A(n9248), .ZN(n9249) );
  OAI21_X1 U10561 ( .B1(n9250), .B2(n9364), .A(n9249), .ZN(P1_U3269) );
  XOR2_X1 U10562 ( .A(n9251), .B(n9252), .Z(n9418) );
  XNOR2_X1 U10563 ( .A(n9253), .B(n9252), .ZN(n9421) );
  OAI211_X1 U10564 ( .C1(n9507), .C2(n9265), .A(n9603), .B(n9254), .ZN(n9416)
         );
  AOI22_X1 U10565 ( .A1(n9255), .A2(n9610), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n4352), .ZN(n9257) );
  NAND2_X1 U10566 ( .A1(n9433), .A2(n9296), .ZN(n9256) );
  OAI211_X1 U10567 ( .C1(n9258), .C2(n9300), .A(n9257), .B(n9256), .ZN(n9259)
         );
  AOI21_X1 U10568 ( .B1(n9260), .B2(n9600), .A(n9259), .ZN(n9261) );
  OAI21_X1 U10569 ( .B1(n9416), .B2(n9305), .A(n9261), .ZN(n9262) );
  AOI21_X1 U10570 ( .B1(n9421), .B2(n9307), .A(n9262), .ZN(n9263) );
  OAI21_X1 U10571 ( .B1(n9418), .B2(n9364), .A(n9263), .ZN(P1_U3270) );
  XNOR2_X1 U10572 ( .A(n9264), .B(n9273), .ZN(n9431) );
  AOI211_X1 U10573 ( .C1(n9266), .C2(n9281), .A(n9348), .B(n9265), .ZN(n9427)
         );
  NOR2_X1 U10574 ( .A1(n9426), .A2(n9614), .ZN(n9272) );
  AOI22_X1 U10575 ( .A1(n9267), .A2(n9610), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n4352), .ZN(n9269) );
  NAND2_X1 U10576 ( .A1(n9442), .A2(n9296), .ZN(n9268) );
  OAI211_X1 U10577 ( .C1(n9270), .C2(n9300), .A(n9269), .B(n9268), .ZN(n9271)
         );
  AOI211_X1 U10578 ( .C1(n9427), .C2(n9608), .A(n9272), .B(n9271), .ZN(n9276)
         );
  XNOR2_X1 U10579 ( .A(n9274), .B(n9273), .ZN(n9429) );
  NAND2_X1 U10580 ( .A1(n9429), .A2(n9307), .ZN(n9275) );
  OAI211_X1 U10581 ( .C1(n9431), .C2(n9364), .A(n9276), .B(n9275), .ZN(
        P1_U3271) );
  XNOR2_X1 U10582 ( .A(n9278), .B(n9277), .ZN(n9439) );
  XNOR2_X1 U10583 ( .A(n9280), .B(n9279), .ZN(n9437) );
  INV_X1 U10584 ( .A(n9295), .ZN(n9282) );
  OAI211_X1 U10585 ( .C1(n4684), .C2(n9282), .A(n9603), .B(n9281), .ZN(n9435)
         );
  AOI22_X1 U10586 ( .A1(n9283), .A2(n9610), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n4352), .ZN(n9285) );
  NAND2_X1 U10587 ( .A1(n9296), .A2(n9432), .ZN(n9284) );
  OAI211_X1 U10588 ( .C1(n9417), .C2(n9300), .A(n9285), .B(n9284), .ZN(n9286)
         );
  AOI21_X1 U10589 ( .B1(n9287), .B2(n9600), .A(n9286), .ZN(n9288) );
  OAI21_X1 U10590 ( .B1(n9435), .B2(n9305), .A(n9288), .ZN(n9289) );
  AOI21_X1 U10591 ( .B1(n9437), .B2(n9307), .A(n9289), .ZN(n9290) );
  OAI21_X1 U10592 ( .B1(n9439), .B2(n9364), .A(n9290), .ZN(P1_U3272) );
  XNOR2_X1 U10593 ( .A(n9291), .B(n9293), .ZN(n9450) );
  OAI21_X1 U10594 ( .B1(n9294), .B2(n9293), .A(n9292), .ZN(n9448) );
  OAI211_X1 U10595 ( .C1(n9445), .C2(n4431), .A(n9603), .B(n9295), .ZN(n9444)
         );
  NAND2_X1 U10596 ( .A1(n9296), .A2(n9440), .ZN(n9299) );
  AOI22_X1 U10597 ( .A1(n4352), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9297), .B2(
        n9610), .ZN(n9298) );
  OAI211_X1 U10598 ( .C1(n9301), .C2(n9300), .A(n9299), .B(n9298), .ZN(n9302)
         );
  AOI21_X1 U10599 ( .B1(n9303), .B2(n9600), .A(n9302), .ZN(n9304) );
  OAI21_X1 U10600 ( .B1(n9444), .B2(n9305), .A(n9304), .ZN(n9306) );
  AOI21_X1 U10601 ( .B1(n9448), .B2(n9307), .A(n9306), .ZN(n9308) );
  OAI21_X1 U10602 ( .B1(n9450), .B2(n9364), .A(n9308), .ZN(P1_U3273) );
  XOR2_X1 U10603 ( .A(n9309), .B(n9311), .Z(n9455) );
  OAI211_X1 U10604 ( .C1(n9312), .C2(n9311), .A(n9310), .B(n9447), .ZN(n9315)
         );
  NAND2_X1 U10605 ( .A1(n9313), .A2(n9647), .ZN(n9314) );
  OAI211_X1 U10606 ( .C1(n9316), .C2(n9670), .A(n9315), .B(n9314), .ZN(n9451)
         );
  AOI211_X1 U10607 ( .C1(n9453), .C2(n9335), .A(n9348), .B(n4431), .ZN(n9452)
         );
  NAND2_X1 U10608 ( .A1(n9452), .A2(n9608), .ZN(n9320) );
  INV_X1 U10609 ( .A(n9317), .ZN(n9318) );
  AOI22_X1 U10610 ( .A1(n4352), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9318), .B2(
        n9610), .ZN(n9319) );
  OAI211_X1 U10611 ( .C1(n9321), .C2(n9614), .A(n9320), .B(n9319), .ZN(n9322)
         );
  AOI21_X1 U10612 ( .B1(n9451), .B2(n9342), .A(n9322), .ZN(n9323) );
  OAI21_X1 U10613 ( .B1(n9455), .B2(n9364), .A(n9323), .ZN(P1_U3274) );
  XNOR2_X1 U10614 ( .A(n9325), .B(n9324), .ZN(n9458) );
  INV_X1 U10615 ( .A(n9458), .ZN(n9344) );
  OAI211_X1 U10616 ( .C1(n9328), .C2(n9327), .A(n9326), .B(n9447), .ZN(n9333)
         );
  OAI22_X1 U10617 ( .A1(n9330), .A2(n9670), .B1(n9329), .B2(n9672), .ZN(n9331)
         );
  INV_X1 U10618 ( .A(n9331), .ZN(n9332) );
  NAND2_X1 U10619 ( .A1(n9333), .A2(n9332), .ZN(n9456) );
  INV_X1 U10620 ( .A(n9334), .ZN(n9347) );
  INV_X1 U10621 ( .A(n9335), .ZN(n9336) );
  AOI211_X1 U10622 ( .C1(n9337), .C2(n9347), .A(n9348), .B(n9336), .ZN(n9457)
         );
  NAND2_X1 U10623 ( .A1(n9457), .A2(n9608), .ZN(n9340) );
  AOI22_X1 U10624 ( .A1(n4352), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9338), .B2(
        n9610), .ZN(n9339) );
  OAI211_X1 U10625 ( .C1(n9516), .C2(n9614), .A(n9340), .B(n9339), .ZN(n9341)
         );
  AOI21_X1 U10626 ( .B1(n9456), .B2(n9342), .A(n9341), .ZN(n9343) );
  OAI21_X1 U10627 ( .B1(n9344), .B2(n9364), .A(n9343), .ZN(P1_U3275) );
  NAND2_X1 U10628 ( .A1(n7850), .A2(n9345), .ZN(n9346) );
  XNOR2_X1 U10629 ( .A(n9346), .B(n9354), .ZN(n9466) );
  AOI211_X1 U10630 ( .C1(n9463), .C2(n9349), .A(n9348), .B(n9334), .ZN(n9462)
         );
  INV_X1 U10631 ( .A(n9350), .ZN(n9351) );
  AOI22_X1 U10632 ( .A1(n4352), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9351), .B2(
        n9610), .ZN(n9352) );
  OAI21_X1 U10633 ( .B1(n9353), .B2(n9614), .A(n9352), .ZN(n9362) );
  AOI21_X1 U10634 ( .B1(n9355), .B2(n9354), .A(n9680), .ZN(n9360) );
  OAI22_X1 U10635 ( .A1(n9357), .A2(n9670), .B1(n9356), .B2(n9672), .ZN(n9358)
         );
  AOI21_X1 U10636 ( .B1(n9360), .B2(n9359), .A(n9358), .ZN(n9465) );
  NOR2_X1 U10637 ( .A1(n9465), .A2(n4352), .ZN(n9361) );
  AOI211_X1 U10638 ( .C1(n9462), .C2(n9608), .A(n9362), .B(n9361), .ZN(n9363)
         );
  OAI21_X1 U10639 ( .B1(n9364), .B2(n9466), .A(n9363), .ZN(P1_U3276) );
  MUX2_X1 U10640 ( .A(n9366), .B(n9479), .S(n9696), .Z(n9367) );
  OAI21_X1 U10641 ( .B1(n9482), .B2(n9461), .A(n9367), .ZN(P1_U3553) );
  NOR2_X1 U10642 ( .A1(n9369), .A2(n9368), .ZN(n9483) );
  MUX2_X1 U10643 ( .A(n9370), .B(n9483), .S(n9696), .Z(n9371) );
  OAI21_X1 U10644 ( .B1(n4650), .B2(n9461), .A(n9371), .ZN(P1_U3552) );
  OAI22_X1 U10645 ( .A1(n9391), .A2(n9672), .B1(n9372), .B2(n9670), .ZN(n9373)
         );
  INV_X1 U10646 ( .A(n9373), .ZN(n9374) );
  AND2_X1 U10647 ( .A1(n9375), .A2(n9374), .ZN(n9378) );
  NAND2_X1 U10648 ( .A1(n9376), .A2(n9447), .ZN(n9377) );
  OAI21_X1 U10649 ( .B1(n9487), .B2(n9461), .A(n9380), .ZN(P1_U3550) );
  OAI22_X1 U10650 ( .A1(n9381), .A2(n9670), .B1(n9402), .B2(n9672), .ZN(n9383)
         );
  AOI211_X1 U10651 ( .C1(n9384), .C2(n9447), .A(n9383), .B(n9382), .ZN(n9385)
         );
  OAI21_X1 U10652 ( .B1(n9386), .B2(n9627), .A(n9385), .ZN(n9488) );
  INV_X1 U10653 ( .A(n9488), .ZN(n9387) );
  MUX2_X1 U10654 ( .A(n9388), .B(n9387), .S(n9696), .Z(n9389) );
  OAI21_X1 U10655 ( .B1(n9491), .B2(n9461), .A(n9389), .ZN(P1_U3549) );
  OAI22_X1 U10656 ( .A1(n9391), .A2(n9670), .B1(n9390), .B2(n9672), .ZN(n9393)
         );
  AOI211_X1 U10657 ( .C1(n9394), .C2(n9447), .A(n9393), .B(n9392), .ZN(n9395)
         );
  OAI21_X1 U10658 ( .B1(n9396), .B2(n9627), .A(n9395), .ZN(n9397) );
  INV_X1 U10659 ( .A(n9397), .ZN(n9492) );
  MUX2_X1 U10660 ( .A(n9398), .B(n9492), .S(n9696), .Z(n9399) );
  OAI21_X1 U10661 ( .B1(n9495), .B2(n9461), .A(n9399), .ZN(P1_U3548) );
  NAND2_X1 U10662 ( .A1(n9414), .A2(n9647), .ZN(n9400) );
  OAI211_X1 U10663 ( .C1(n9402), .C2(n9670), .A(n9401), .B(n9400), .ZN(n9405)
         );
  NOR2_X1 U10664 ( .A1(n9403), .A2(n9627), .ZN(n9404) );
  AOI211_X1 U10665 ( .C1(n9447), .C2(n9406), .A(n9405), .B(n9404), .ZN(n9496)
         );
  MUX2_X1 U10666 ( .A(n9407), .B(n9496), .S(n9696), .Z(n9408) );
  OAI21_X1 U10667 ( .B1(n9499), .B2(n9461), .A(n9408), .ZN(P1_U3547) );
  AOI211_X1 U10668 ( .C1(n9411), .C2(n9682), .A(n9410), .B(n9409), .ZN(n9500)
         );
  MUX2_X1 U10669 ( .A(n9412), .B(n9500), .S(n9696), .Z(n9413) );
  OAI21_X1 U10670 ( .B1(n9503), .B2(n9461), .A(n9413), .ZN(P1_U3546) );
  NAND2_X1 U10671 ( .A1(n9414), .A2(n9441), .ZN(n9415) );
  OAI211_X1 U10672 ( .C1(n9417), .C2(n9672), .A(n9416), .B(n9415), .ZN(n9420)
         );
  NOR2_X1 U10673 ( .A1(n9418), .A2(n9627), .ZN(n9419) );
  AOI211_X1 U10674 ( .C1(n9421), .C2(n9447), .A(n9420), .B(n9419), .ZN(n9504)
         );
  MUX2_X1 U10675 ( .A(n9422), .B(n9504), .S(n9696), .Z(n9423) );
  OAI21_X1 U10676 ( .B1(n9507), .B2(n9461), .A(n9423), .ZN(P1_U3545) );
  AOI22_X1 U10677 ( .A1(n9441), .A2(n9424), .B1(n9442), .B2(n9647), .ZN(n9425)
         );
  OAI21_X1 U10678 ( .B1(n9426), .B2(n9664), .A(n9425), .ZN(n9428) );
  AOI211_X1 U10679 ( .C1(n9429), .C2(n9447), .A(n9428), .B(n9427), .ZN(n9430)
         );
  OAI21_X1 U10680 ( .B1(n9431), .B2(n9627), .A(n9430), .ZN(n9508) );
  MUX2_X1 U10681 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9508), .S(n9696), .Z(
        P1_U3544) );
  AOI22_X1 U10682 ( .A1(n9433), .A2(n9441), .B1(n9647), .B2(n9432), .ZN(n9434)
         );
  OAI211_X1 U10683 ( .C1(n4684), .C2(n9664), .A(n9435), .B(n9434), .ZN(n9436)
         );
  AOI21_X1 U10684 ( .B1(n9437), .B2(n9447), .A(n9436), .ZN(n9438) );
  OAI21_X1 U10685 ( .B1(n9439), .B2(n9627), .A(n9438), .ZN(n9509) );
  MUX2_X1 U10686 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9509), .S(n9696), .Z(
        P1_U3543) );
  AOI22_X1 U10687 ( .A1(n9442), .A2(n9441), .B1(n9647), .B2(n9440), .ZN(n9443)
         );
  OAI211_X1 U10688 ( .C1(n9445), .C2(n9664), .A(n9444), .B(n9443), .ZN(n9446)
         );
  AOI21_X1 U10689 ( .B1(n9448), .B2(n9447), .A(n9446), .ZN(n9449) );
  OAI21_X1 U10690 ( .B1(n9450), .B2(n9627), .A(n9449), .ZN(n9510) );
  MUX2_X1 U10691 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9510), .S(n9696), .Z(
        P1_U3542) );
  AOI211_X1 U10692 ( .C1(n9677), .C2(n9453), .A(n9452), .B(n9451), .ZN(n9454)
         );
  OAI21_X1 U10693 ( .B1(n9455), .B2(n9627), .A(n9454), .ZN(n9511) );
  MUX2_X1 U10694 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9511), .S(n9696), .Z(
        P1_U3541) );
  AOI211_X1 U10695 ( .C1(n9458), .C2(n9682), .A(n9457), .B(n9456), .ZN(n9512)
         );
  MUX2_X1 U10696 ( .A(n9459), .B(n9512), .S(n9696), .Z(n9460) );
  OAI21_X1 U10697 ( .B1(n9516), .B2(n9461), .A(n9460), .ZN(P1_U3540) );
  AOI21_X1 U10698 ( .B1(n9677), .B2(n9463), .A(n9462), .ZN(n9464) );
  OAI211_X1 U10699 ( .C1(n9466), .C2(n9627), .A(n9465), .B(n9464), .ZN(n9517)
         );
  MUX2_X1 U10700 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9517), .S(n9696), .Z(
        P1_U3539) );
  NAND3_X1 U10701 ( .A1(n7850), .A2(n9467), .A3(n9682), .ZN(n9472) );
  AOI22_X1 U10702 ( .A1(n9469), .A2(n9603), .B1(n9677), .B2(n9468), .ZN(n9470)
         );
  NAND3_X1 U10703 ( .A1(n9472), .A2(n9471), .A3(n9470), .ZN(n9518) );
  MUX2_X1 U10704 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9518), .S(n9696), .Z(
        P1_U3538) );
  AOI21_X1 U10705 ( .B1(n9677), .B2(n9474), .A(n9473), .ZN(n9475) );
  OAI211_X1 U10706 ( .C1(n9477), .C2(n9627), .A(n9476), .B(n9475), .ZN(n9519)
         );
  MUX2_X1 U10707 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9519), .S(n9696), .Z(
        P1_U3537) );
  MUX2_X1 U10708 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9478), .S(n9696), .Z(
        P1_U3522) );
  MUX2_X1 U10709 ( .A(n9480), .B(n9479), .S(n9685), .Z(n9481) );
  OAI21_X1 U10710 ( .B1(n9482), .B2(n9515), .A(n9481), .ZN(P1_U3521) );
  MUX2_X1 U10711 ( .A(n9484), .B(n9483), .S(n9685), .Z(n9485) );
  OAI21_X1 U10712 ( .B1(n4650), .B2(n9515), .A(n9485), .ZN(P1_U3520) );
  MUX2_X1 U10713 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9488), .S(n9685), .Z(n9489) );
  INV_X1 U10714 ( .A(n9489), .ZN(n9490) );
  OAI21_X1 U10715 ( .B1(n9491), .B2(n9515), .A(n9490), .ZN(P1_U3517) );
  INV_X1 U10716 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n9493) );
  MUX2_X1 U10717 ( .A(n9493), .B(n9492), .S(n9685), .Z(n9494) );
  OAI21_X1 U10718 ( .B1(n9495), .B2(n9515), .A(n9494), .ZN(P1_U3516) );
  INV_X1 U10719 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9497) );
  MUX2_X1 U10720 ( .A(n9497), .B(n9496), .S(n9685), .Z(n9498) );
  OAI21_X1 U10721 ( .B1(n9499), .B2(n9515), .A(n9498), .ZN(P1_U3515) );
  INV_X1 U10722 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9501) );
  MUX2_X1 U10723 ( .A(n9501), .B(n9500), .S(n9685), .Z(n9502) );
  OAI21_X1 U10724 ( .B1(n9503), .B2(n9515), .A(n9502), .ZN(P1_U3514) );
  INV_X1 U10725 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n9505) );
  MUX2_X1 U10726 ( .A(n9505), .B(n9504), .S(n9685), .Z(n9506) );
  OAI21_X1 U10727 ( .B1(n9507), .B2(n9515), .A(n9506), .ZN(P1_U3513) );
  MUX2_X1 U10728 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9508), .S(n9685), .Z(
        P1_U3512) );
  MUX2_X1 U10729 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9509), .S(n9685), .Z(
        P1_U3511) );
  MUX2_X1 U10730 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9510), .S(n9685), .Z(
        P1_U3510) );
  MUX2_X1 U10731 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9511), .S(n9685), .Z(
        P1_U3509) );
  INV_X1 U10732 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n9513) );
  MUX2_X1 U10733 ( .A(n9513), .B(n9512), .S(n9685), .Z(n9514) );
  OAI21_X1 U10734 ( .B1(n9516), .B2(n9515), .A(n9514), .ZN(P1_U3507) );
  MUX2_X1 U10735 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9517), .S(n9685), .Z(
        P1_U3504) );
  MUX2_X1 U10736 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9518), .S(n9685), .Z(
        P1_U3501) );
  MUX2_X1 U10737 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9519), .S(n9685), .Z(
        P1_U3498) );
  MUX2_X1 U10738 ( .A(n9520), .B(P1_D_REG_0__SCAN_IN), .S(n9621), .Z(P1_U3439)
         );
  OAI222_X1 U10739 ( .A1(n9525), .A2(n9524), .B1(P1_U3086), .B2(n9523), .C1(
        n9522), .C2(n9521), .ZN(P1_U3326) );
  INV_X1 U10740 ( .A(n9526), .ZN(n9527) );
  MUX2_X1 U10741 ( .A(n9527), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U10742 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9541) );
  AOI211_X1 U10743 ( .C1(n9531), .C2(n9530), .A(n9529), .B(n9528), .ZN(n9537)
         );
  AOI211_X1 U10744 ( .C1(n9535), .C2(n9534), .A(n9533), .B(n9532), .ZN(n9536)
         );
  AOI211_X1 U10745 ( .C1(n9564), .C2(n9538), .A(n9537), .B(n9536), .ZN(n9540)
         );
  OAI211_X1 U10746 ( .C1(n9590), .C2(n9541), .A(n9540), .B(n9539), .ZN(
        P1_U3253) );
  INV_X1 U10747 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9556) );
  INV_X1 U10748 ( .A(n9542), .ZN(n9543) );
  OAI211_X1 U10749 ( .C1(n9545), .C2(n9544), .A(n9575), .B(n9543), .ZN(n9553)
         );
  INV_X1 U10750 ( .A(n9546), .ZN(n9547) );
  OAI211_X1 U10751 ( .C1(n9549), .C2(n9548), .A(n9580), .B(n9547), .ZN(n9552)
         );
  NAND2_X1 U10752 ( .A1(n9564), .A2(n9550), .ZN(n9551) );
  AND3_X1 U10753 ( .A1(n9553), .A2(n9552), .A3(n9551), .ZN(n9555) );
  OAI211_X1 U10754 ( .C1(n9590), .C2(n9556), .A(n9555), .B(n9554), .ZN(
        P1_U3251) );
  XNOR2_X1 U10755 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10756 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10757 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n9570) );
  OAI211_X1 U10758 ( .C1(n9559), .C2(n9558), .A(n9575), .B(n9557), .ZN(n9567)
         );
  OAI211_X1 U10759 ( .C1(n9562), .C2(n9561), .A(n9580), .B(n9560), .ZN(n9566)
         );
  NAND2_X1 U10760 ( .A1(n9564), .A2(n9563), .ZN(n9565) );
  AND3_X1 U10761 ( .A1(n9567), .A2(n9566), .A3(n9565), .ZN(n9569) );
  OAI211_X1 U10762 ( .C1(n9590), .C2(n9570), .A(n9569), .B(n9568), .ZN(
        P1_U3249) );
  INV_X1 U10763 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n9589) );
  AOI21_X1 U10764 ( .B1(n9573), .B2(n9572), .A(n9571), .ZN(n9574) );
  NAND2_X1 U10765 ( .A1(n9575), .A2(n9574), .ZN(n9582) );
  AOI21_X1 U10766 ( .B1(n9578), .B2(n9577), .A(n9576), .ZN(n9579) );
  NAND2_X1 U10767 ( .A1(n9580), .A2(n9579), .ZN(n9581) );
  OAI211_X1 U10768 ( .C1(n9584), .C2(n9583), .A(n9582), .B(n9581), .ZN(n9585)
         );
  INV_X1 U10769 ( .A(n9585), .ZN(n9588) );
  INV_X1 U10770 ( .A(n9586), .ZN(n9587) );
  OAI211_X1 U10771 ( .C1(n9590), .C2(n9589), .A(n9588), .B(n9587), .ZN(
        P1_U3254) );
  XNOR2_X1 U10772 ( .A(n9591), .B(n9595), .ZN(n9668) );
  OAI22_X1 U10773 ( .A1(n9592), .A2(n9672), .B1(n9673), .B2(n9670), .ZN(n9597)
         );
  INV_X1 U10774 ( .A(n9593), .ZN(n9594) );
  AOI211_X1 U10775 ( .C1(n9595), .C2(n4435), .A(n9680), .B(n9594), .ZN(n9596)
         );
  AOI211_X1 U10776 ( .C1(n9668), .C2(n9598), .A(n9597), .B(n9596), .ZN(n9665)
         );
  AOI222_X1 U10777 ( .A1(n9601), .A2(n9600), .B1(P1_REG2_REG_11__SCAN_IN), 
        .B2(n4352), .C1(n9599), .C2(n9610), .ZN(n9607) );
  OAI211_X1 U10778 ( .C1(n4681), .C2(n4372), .A(n4683), .B(n9603), .ZN(n9663)
         );
  INV_X1 U10779 ( .A(n9663), .ZN(n9604) );
  AOI22_X1 U10780 ( .A1(n9668), .A2(n9605), .B1(n9608), .B2(n9604), .ZN(n9606)
         );
  OAI211_X1 U10781 ( .C1(n4352), .C2(n9665), .A(n9607), .B(n9606), .ZN(
        P1_U3282) );
  NAND2_X1 U10782 ( .A1(n9609), .A2(n9608), .ZN(n9613) );
  AOI22_X1 U10783 ( .A1(n4352), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n9611), .B2(
        n9610), .ZN(n9612) );
  OAI211_X1 U10784 ( .C1(n9615), .C2(n9614), .A(n9613), .B(n9612), .ZN(n9616)
         );
  AOI21_X1 U10785 ( .B1(n9618), .B2(n9617), .A(n9616), .ZN(n9619) );
  OAI21_X1 U10786 ( .B1(n4352), .B2(n9620), .A(n9619), .ZN(P1_U3289) );
  AND2_X1 U10787 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9621), .ZN(P1_U3294) );
  AND2_X1 U10788 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9621), .ZN(P1_U3295) );
  AND2_X1 U10789 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9621), .ZN(P1_U3296) );
  AND2_X1 U10790 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9621), .ZN(P1_U3297) );
  AND2_X1 U10791 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9621), .ZN(P1_U3298) );
  AND2_X1 U10792 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9621), .ZN(P1_U3299) );
  AND2_X1 U10793 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9621), .ZN(P1_U3300) );
  AND2_X1 U10794 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9621), .ZN(P1_U3301) );
  AND2_X1 U10795 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9621), .ZN(P1_U3302) );
  AND2_X1 U10796 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9621), .ZN(P1_U3303) );
  AND2_X1 U10797 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9621), .ZN(P1_U3304) );
  AND2_X1 U10798 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9621), .ZN(P1_U3305) );
  AND2_X1 U10799 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9621), .ZN(P1_U3306) );
  AND2_X1 U10800 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9621), .ZN(P1_U3307) );
  AND2_X1 U10801 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9621), .ZN(P1_U3308) );
  AND2_X1 U10802 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9621), .ZN(P1_U3309) );
  AND2_X1 U10803 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9621), .ZN(P1_U3310) );
  AND2_X1 U10804 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9621), .ZN(P1_U3311) );
  AND2_X1 U10805 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9621), .ZN(P1_U3312) );
  AND2_X1 U10806 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9621), .ZN(P1_U3313) );
  AND2_X1 U10807 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9621), .ZN(P1_U3314) );
  AND2_X1 U10808 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9621), .ZN(P1_U3315) );
  AND2_X1 U10809 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9621), .ZN(P1_U3316) );
  AND2_X1 U10810 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9621), .ZN(P1_U3317) );
  AND2_X1 U10811 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9621), .ZN(P1_U3318) );
  AND2_X1 U10812 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9621), .ZN(P1_U3319) );
  AND2_X1 U10813 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9621), .ZN(P1_U3320) );
  AND2_X1 U10814 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9621), .ZN(P1_U3321) );
  AND2_X1 U10815 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9621), .ZN(P1_U3322) );
  AND2_X1 U10816 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9621), .ZN(P1_U3323) );
  AOI21_X1 U10817 ( .B1(n9677), .B2(n9623), .A(n9622), .ZN(n9624) );
  OAI211_X1 U10818 ( .C1(n9627), .C2(n9626), .A(n9625), .B(n9624), .ZN(n9628)
         );
  INV_X1 U10819 ( .A(n9628), .ZN(n9686) );
  AOI22_X1 U10820 ( .A1(n9685), .A2(n9686), .B1(n5214), .B2(n9684), .ZN(
        P1_U3462) );
  OAI21_X1 U10821 ( .B1(n9630), .B2(n9664), .A(n9629), .ZN(n9632) );
  AOI211_X1 U10822 ( .C1(n9682), .C2(n9633), .A(n9632), .B(n9631), .ZN(n9687)
         );
  AOI22_X1 U10823 ( .A1(n9685), .A2(n9687), .B1(n5261), .B2(n9684), .ZN(
        P1_U3468) );
  INV_X1 U10824 ( .A(n9634), .ZN(n9669) );
  OAI21_X1 U10825 ( .B1(n9636), .B2(n9664), .A(n9635), .ZN(n9638) );
  AOI211_X1 U10826 ( .C1(n9669), .C2(n9639), .A(n9638), .B(n9637), .ZN(n9688)
         );
  AOI22_X1 U10827 ( .A1(n9685), .A2(n9688), .B1(n5315), .B2(n9684), .ZN(
        P1_U3474) );
  OAI21_X1 U10828 ( .B1(n9641), .B2(n9664), .A(n9640), .ZN(n9642) );
  AOI21_X1 U10829 ( .B1(n9643), .B2(n9669), .A(n9642), .ZN(n9644) );
  AOI22_X1 U10830 ( .A1(n9685), .A2(n9689), .B1(n5334), .B2(n9684), .ZN(
        P1_U3477) );
  AOI22_X1 U10831 ( .A1(n9648), .A2(n9677), .B1(n9647), .B2(n9646), .ZN(n9649)
         );
  OAI211_X1 U10832 ( .C1(n9651), .C2(n9680), .A(n9650), .B(n9649), .ZN(n9652)
         );
  AOI21_X1 U10833 ( .B1(n9682), .B2(n9653), .A(n9652), .ZN(n9690) );
  AOI22_X1 U10834 ( .A1(n9685), .A2(n9690), .B1(n5363), .B2(n9684), .ZN(
        P1_U3480) );
  OAI22_X1 U10835 ( .A1(n9655), .A2(n9672), .B1(n9654), .B2(n9670), .ZN(n9657)
         );
  AOI211_X1 U10836 ( .C1(n9677), .C2(n9658), .A(n9657), .B(n9656), .ZN(n9659)
         );
  OAI21_X1 U10837 ( .B1(n9680), .B2(n9660), .A(n9659), .ZN(n9661) );
  AOI21_X1 U10838 ( .B1(n9682), .B2(n9662), .A(n9661), .ZN(n9692) );
  AOI22_X1 U10839 ( .A1(n9685), .A2(n9692), .B1(n5389), .B2(n9684), .ZN(
        P1_U3483) );
  OAI21_X1 U10840 ( .B1(n4681), .B2(n9664), .A(n9663), .ZN(n9667) );
  INV_X1 U10841 ( .A(n9665), .ZN(n9666) );
  AOI211_X1 U10842 ( .C1(n9669), .C2(n9668), .A(n9667), .B(n9666), .ZN(n9693)
         );
  AOI22_X1 U10843 ( .A1(n9685), .A2(n9693), .B1(n5412), .B2(n9684), .ZN(
        P1_U3486) );
  OAI22_X1 U10844 ( .A1(n9673), .A2(n9672), .B1(n9671), .B2(n9670), .ZN(n9675)
         );
  AOI211_X1 U10845 ( .C1(n9677), .C2(n9676), .A(n9675), .B(n9674), .ZN(n9678)
         );
  OAI21_X1 U10846 ( .B1(n9680), .B2(n9679), .A(n9678), .ZN(n9681) );
  AOI21_X1 U10847 ( .B1(n9683), .B2(n9682), .A(n9681), .ZN(n9695) );
  AOI22_X1 U10848 ( .A1(n9685), .A2(n9695), .B1(n5469), .B2(n9684), .ZN(
        P1_U3492) );
  AOI22_X1 U10849 ( .A1(n9696), .A2(n9686), .B1(n6584), .B2(n9694), .ZN(
        P1_U3525) );
  AOI22_X1 U10850 ( .A1(n9696), .A2(n9687), .B1(n5262), .B2(n9694), .ZN(
        P1_U3527) );
  AOI22_X1 U10851 ( .A1(n9696), .A2(n9688), .B1(n6591), .B2(n9694), .ZN(
        P1_U3529) );
  AOI22_X1 U10852 ( .A1(n9696), .A2(n9689), .B1(n5333), .B2(n9694), .ZN(
        P1_U3530) );
  AOI22_X1 U10853 ( .A1(n9696), .A2(n9690), .B1(n5362), .B2(n9694), .ZN(
        P1_U3531) );
  INV_X1 U10854 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n9691) );
  AOI22_X1 U10855 ( .A1(n9696), .A2(n9692), .B1(n9691), .B2(n9694), .ZN(
        P1_U3532) );
  AOI22_X1 U10856 ( .A1(n9696), .A2(n9693), .B1(n6595), .B2(n9694), .ZN(
        P1_U3533) );
  AOI22_X1 U10857 ( .A1(n9696), .A2(n9695), .B1(n5470), .B2(n9694), .ZN(
        P1_U3535) );
  NAND2_X1 U10858 ( .A1(n9698), .A2(n9697), .ZN(n9700) );
  AOI21_X1 U10859 ( .B1(n9701), .B2(n9700), .A(n9699), .ZN(n9712) );
  OR3_X1 U10860 ( .A1(n9704), .A2(n9703), .A3(n9702), .ZN(n9705) );
  AOI21_X1 U10861 ( .B1(n9706), .B2(n9705), .A(n9872), .ZN(n9711) );
  NOR2_X1 U10862 ( .A1(n9708), .A2(n9707), .ZN(n9709) );
  NOR4_X1 U10863 ( .A1(n9712), .A2(n9711), .A3(n9710), .A4(n9709), .ZN(n9717)
         );
  XNOR2_X1 U10864 ( .A(n9714), .B(n9713), .ZN(n9715) );
  AOI22_X1 U10865 ( .A1(n9715), .A2(n9866), .B1(n9857), .B2(
        P2_ADDR_REG_8__SCAN_IN), .ZN(n9716) );
  NAND2_X1 U10866 ( .A1(n9717), .A2(n9716), .ZN(P2_U3190) );
  AOI22_X1 U10867 ( .A1(n9718), .A2(n9858), .B1(n9857), .B2(
        P2_ADDR_REG_9__SCAN_IN), .ZN(n9733) );
  OAI21_X1 U10868 ( .B1(n9721), .B2(n9720), .A(n9719), .ZN(n9725) );
  OAI21_X1 U10869 ( .B1(n9723), .B2(P2_REG1_REG_9__SCAN_IN), .A(n9722), .ZN(
        n9724) );
  AOI22_X1 U10870 ( .A1(n9725), .A2(n9866), .B1(n9867), .B2(n9724), .ZN(n9732)
         );
  INV_X1 U10871 ( .A(n9726), .ZN(n9731) );
  AOI21_X1 U10872 ( .B1(n5973), .B2(n9728), .A(n9727), .ZN(n9729) );
  OR2_X1 U10873 ( .A1(n9729), .A2(n9872), .ZN(n9730) );
  NAND4_X1 U10874 ( .A1(n9733), .A2(n9732), .A3(n9731), .A4(n9730), .ZN(
        P2_U3191) );
  AOI22_X1 U10875 ( .A1(n9857), .A2(P2_ADDR_REG_10__SCAN_IN), .B1(n9734), .B2(
        n9858), .ZN(n9751) );
  OAI21_X1 U10876 ( .B1(n9737), .B2(n9736), .A(n9735), .ZN(n9742) );
  OAI21_X1 U10877 ( .B1(n9740), .B2(n9739), .A(n9738), .ZN(n9741) );
  AOI22_X1 U10878 ( .A1(n9866), .A2(n9742), .B1(n9867), .B2(n9741), .ZN(n9750)
         );
  INV_X1 U10879 ( .A(n9743), .ZN(n9749) );
  AOI21_X1 U10880 ( .B1(n9746), .B2(n9745), .A(n9744), .ZN(n9747) );
  OR2_X1 U10881 ( .A1(n9747), .A2(n9872), .ZN(n9748) );
  NAND4_X1 U10882 ( .A1(n9751), .A2(n9750), .A3(n9749), .A4(n9748), .ZN(
        P2_U3192) );
  AOI22_X1 U10883 ( .A1(n9752), .A2(n9858), .B1(n9857), .B2(
        P2_ADDR_REG_11__SCAN_IN), .ZN(n9767) );
  OAI21_X1 U10884 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n9754), .A(n9753), .ZN(
        n9759) );
  OAI21_X1 U10885 ( .B1(n9757), .B2(n9756), .A(n9755), .ZN(n9758) );
  AOI22_X1 U10886 ( .A1(n9759), .A2(n9867), .B1(n9866), .B2(n9758), .ZN(n9766)
         );
  INV_X1 U10887 ( .A(n9760), .ZN(n9765) );
  AOI21_X1 U10888 ( .B1(n9762), .B2(n7423), .A(n9761), .ZN(n9763) );
  OR2_X1 U10889 ( .A1(n9763), .A2(n9872), .ZN(n9764) );
  NAND4_X1 U10890 ( .A1(n9767), .A2(n9766), .A3(n9765), .A4(n9764), .ZN(
        P2_U3193) );
  AOI22_X1 U10891 ( .A1(n9857), .A2(P2_ADDR_REG_12__SCAN_IN), .B1(n9768), .B2(
        n9858), .ZN(n9786) );
  OAI21_X1 U10892 ( .B1(n9771), .B2(n9770), .A(n9769), .ZN(n9776) );
  OAI21_X1 U10893 ( .B1(n9774), .B2(n9773), .A(n9772), .ZN(n9775) );
  AOI22_X1 U10894 ( .A1(n9776), .A2(n9867), .B1(n9866), .B2(n9775), .ZN(n9785)
         );
  INV_X1 U10895 ( .A(n9777), .ZN(n9784) );
  INV_X1 U10896 ( .A(n9778), .ZN(n9779) );
  AOI21_X1 U10897 ( .B1(n9781), .B2(n9780), .A(n9779), .ZN(n9782) );
  OR2_X1 U10898 ( .A1(n9782), .A2(n9872), .ZN(n9783) );
  NAND4_X1 U10899 ( .A1(n9786), .A2(n9785), .A3(n9784), .A4(n9783), .ZN(
        P2_U3194) );
  AOI22_X1 U10900 ( .A1(n9787), .A2(n9858), .B1(n9857), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n9804) );
  OAI21_X1 U10901 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n9789), .A(n9788), .ZN(
        n9794) );
  OAI21_X1 U10902 ( .B1(n9792), .B2(n9791), .A(n9790), .ZN(n9793) );
  AOI22_X1 U10903 ( .A1(n9794), .A2(n9867), .B1(n9866), .B2(n9793), .ZN(n9803)
         );
  INV_X1 U10904 ( .A(n9795), .ZN(n9802) );
  INV_X1 U10905 ( .A(n9796), .ZN(n9797) );
  NOR2_X1 U10906 ( .A1(n9797), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n9800) );
  OAI21_X1 U10907 ( .B1(n9800), .B2(n9799), .A(n9798), .ZN(n9801) );
  NAND4_X1 U10908 ( .A1(n9804), .A2(n9803), .A3(n9802), .A4(n9801), .ZN(
        P2_U3195) );
  AOI22_X1 U10909 ( .A1(n9805), .A2(n9858), .B1(n9857), .B2(
        P2_ADDR_REG_14__SCAN_IN), .ZN(n9822) );
  OAI21_X1 U10910 ( .B1(n9808), .B2(n9807), .A(n9806), .ZN(n9813) );
  OAI21_X1 U10911 ( .B1(n9811), .B2(n9810), .A(n9809), .ZN(n9812) );
  AOI22_X1 U10912 ( .A1(n9813), .A2(n9867), .B1(n9866), .B2(n9812), .ZN(n9821)
         );
  INV_X1 U10913 ( .A(n9814), .ZN(n9820) );
  AOI21_X1 U10914 ( .B1(n9817), .B2(n9816), .A(n9815), .ZN(n9818) );
  OR2_X1 U10915 ( .A1(n9818), .A2(n9872), .ZN(n9819) );
  NAND4_X1 U10916 ( .A1(n9822), .A2(n9821), .A3(n9820), .A4(n9819), .ZN(
        P2_U3196) );
  AOI22_X1 U10917 ( .A1(n9823), .A2(n9858), .B1(n9857), .B2(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n9838) );
  OAI21_X1 U10918 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n9825), .A(n9824), .ZN(
        n9830) );
  OAI21_X1 U10919 ( .B1(n9828), .B2(n9827), .A(n9826), .ZN(n9829) );
  AOI22_X1 U10920 ( .A1(n9830), .A2(n9867), .B1(n9866), .B2(n9829), .ZN(n9837)
         );
  INV_X1 U10921 ( .A(n9831), .ZN(n9836) );
  AOI21_X1 U10922 ( .B1(n9833), .B2(n8694), .A(n9832), .ZN(n9834) );
  OR2_X1 U10923 ( .A1(n9872), .A2(n9834), .ZN(n9835) );
  NAND4_X1 U10924 ( .A1(n9838), .A2(n9837), .A3(n9836), .A4(n9835), .ZN(
        P2_U3197) );
  AOI22_X1 U10925 ( .A1(n9839), .A2(n9858), .B1(n9857), .B2(
        P2_ADDR_REG_16__SCAN_IN), .ZN(n9856) );
  OAI21_X1 U10926 ( .B1(n9842), .B2(n9841), .A(n9840), .ZN(n9847) );
  OAI21_X1 U10927 ( .B1(n9845), .B2(n9844), .A(n9843), .ZN(n9846) );
  AOI22_X1 U10928 ( .A1(n9847), .A2(n9867), .B1(n9866), .B2(n9846), .ZN(n9855)
         );
  INV_X1 U10929 ( .A(n9848), .ZN(n9854) );
  AOI21_X1 U10930 ( .B1(n9851), .B2(n9850), .A(n9849), .ZN(n9852) );
  OR2_X1 U10931 ( .A1(n9852), .A2(n9872), .ZN(n9853) );
  NAND4_X1 U10932 ( .A1(n9856), .A2(n9855), .A3(n9854), .A4(n9853), .ZN(
        P2_U3198) );
  AOI22_X1 U10933 ( .A1(n9859), .A2(n9858), .B1(n9857), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n9876) );
  OAI21_X1 U10934 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n9861), .A(n9860), .ZN(
        n9868) );
  OAI21_X1 U10935 ( .B1(n9864), .B2(n9863), .A(n9862), .ZN(n9865) );
  AOI22_X1 U10936 ( .A1(n9868), .A2(n9867), .B1(n9866), .B2(n9865), .ZN(n9875)
         );
  NAND2_X1 U10937 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3151), .ZN(n9874) );
  AOI21_X1 U10938 ( .B1(n9870), .B2(n8669), .A(n9869), .ZN(n9871) );
  OR2_X1 U10939 ( .A1(n9872), .A2(n9871), .ZN(n9873) );
  NAND4_X1 U10940 ( .A1(n9876), .A2(n9875), .A3(n9874), .A4(n9873), .ZN(
        P2_U3199) );
  XOR2_X1 U10941 ( .A(n9877), .B(n9884), .Z(n9882) );
  AOI222_X1 U10942 ( .A1(n9883), .A2(n9882), .B1(n9881), .B2(n9880), .C1(n9879), .C2(n9878), .ZN(n9927) );
  XNOR2_X1 U10943 ( .A(n9885), .B(n9884), .ZN(n9925) );
  INV_X1 U10944 ( .A(n9886), .ZN(n9887) );
  AOI222_X1 U10945 ( .A1(n9925), .A2(n9888), .B1(n9887), .B2(n9905), .C1(n9924), .C2(n4350), .ZN(n9889) );
  OAI221_X1 U10946 ( .B1(n9910), .B2(n9927), .C1(n8710), .C2(n6980), .A(n9889), 
        .ZN(P2_U3229) );
  XNOR2_X1 U10947 ( .A(n9897), .B(n9890), .ZN(n9919) );
  OAI22_X1 U10948 ( .A1(n9894), .A2(n9893), .B1(n9892), .B2(n9891), .ZN(n9902)
         );
  NAND3_X1 U10949 ( .A1(n9898), .A2(n9897), .A3(n9896), .ZN(n9900) );
  AOI21_X1 U10950 ( .B1(n9895), .B2(n9900), .A(n9899), .ZN(n9901) );
  AOI211_X1 U10951 ( .C1(n9919), .C2(n9903), .A(n9902), .B(n9901), .ZN(n9916)
         );
  NOR2_X1 U10952 ( .A1(n9904), .A2(n9955), .ZN(n9918) );
  AOI22_X1 U10953 ( .A1(n9918), .A2(n9906), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n9905), .ZN(n9909) );
  AOI22_X1 U10954 ( .A1(n9919), .A2(n9907), .B1(P2_REG2_REG_2__SCAN_IN), .B2(
        n9910), .ZN(n9908) );
  OAI221_X1 U10955 ( .B1(n9910), .B2(n9916), .C1(n9910), .C2(n9909), .A(n9908), 
        .ZN(P2_U3231) );
  INV_X1 U10956 ( .A(n9911), .ZN(n9915) );
  OAI22_X1 U10957 ( .A1(n9913), .A2(n9957), .B1(n9912), .B2(n9955), .ZN(n9914)
         );
  NOR2_X1 U10958 ( .A1(n9915), .A2(n9914), .ZN(n9972) );
  AOI22_X1 U10959 ( .A1(n9970), .A2(n5858), .B1(n9972), .B2(n9968), .ZN(
        P2_U3393) );
  INV_X1 U10960 ( .A(n9916), .ZN(n9917) );
  AOI211_X1 U10961 ( .C1(n9919), .C2(n4693), .A(n9918), .B(n9917), .ZN(n9973)
         );
  AOI22_X1 U10962 ( .A1(n9970), .A2(n5877), .B1(n9973), .B2(n9968), .ZN(
        P2_U3396) );
  AOI22_X1 U10963 ( .A1(n9921), .A2(n9948), .B1(n9967), .B2(n9920), .ZN(n9922)
         );
  AND2_X1 U10964 ( .A1(n9923), .A2(n9922), .ZN(n9975) );
  AOI22_X1 U10965 ( .A1(n9970), .A2(n5889), .B1(n9975), .B2(n9968), .ZN(
        P2_U3399) );
  INV_X1 U10966 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n9928) );
  AOI22_X1 U10967 ( .A1(n9925), .A2(n9948), .B1(n9967), .B2(n9924), .ZN(n9926)
         );
  AND2_X1 U10968 ( .A1(n9927), .A2(n9926), .ZN(n9976) );
  AOI22_X1 U10969 ( .A1(n9970), .A2(n9928), .B1(n9976), .B2(n9968), .ZN(
        P2_U3402) );
  INV_X1 U10970 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9933) );
  NOR2_X1 U10971 ( .A1(n9929), .A2(n9955), .ZN(n9931) );
  AOI211_X1 U10972 ( .C1(n4693), .C2(n9932), .A(n9931), .B(n9930), .ZN(n9977)
         );
  AOI22_X1 U10973 ( .A1(n9970), .A2(n9933), .B1(n9977), .B2(n9968), .ZN(
        P2_U3405) );
  INV_X1 U10974 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9938) );
  NOR2_X1 U10975 ( .A1(n9934), .A2(n9955), .ZN(n9936) );
  AOI211_X1 U10976 ( .C1(n9937), .C2(n9948), .A(n9936), .B(n9935), .ZN(n9978)
         );
  AOI22_X1 U10977 ( .A1(n9970), .A2(n9938), .B1(n9978), .B2(n9968), .ZN(
        P2_U3408) );
  INV_X1 U10978 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9943) );
  OAI22_X1 U10979 ( .A1(n9940), .A2(n9957), .B1(n9939), .B2(n9955), .ZN(n9941)
         );
  NOR2_X1 U10980 ( .A1(n9942), .A2(n9941), .ZN(n9980) );
  AOI22_X1 U10981 ( .A1(n9970), .A2(n9943), .B1(n9980), .B2(n9968), .ZN(
        P2_U3411) );
  INV_X1 U10982 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9949) );
  NOR2_X1 U10983 ( .A1(n9944), .A2(n9955), .ZN(n9946) );
  AOI211_X1 U10984 ( .C1(n9948), .C2(n9947), .A(n9946), .B(n9945), .ZN(n9981)
         );
  AOI22_X1 U10985 ( .A1(n9970), .A2(n9949), .B1(n9981), .B2(n9968), .ZN(
        P2_U3414) );
  INV_X1 U10986 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9954) );
  OAI22_X1 U10987 ( .A1(n9951), .A2(n9957), .B1(n9950), .B2(n9955), .ZN(n9952)
         );
  NOR2_X1 U10988 ( .A1(n9953), .A2(n9952), .ZN(n9982) );
  AOI22_X1 U10989 ( .A1(n9970), .A2(n9954), .B1(n9982), .B2(n9968), .ZN(
        P2_U3417) );
  INV_X1 U10990 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9961) );
  OAI22_X1 U10991 ( .A1(n9958), .A2(n9957), .B1(n9956), .B2(n9955), .ZN(n9959)
         );
  NOR2_X1 U10992 ( .A1(n9960), .A2(n9959), .ZN(n9983) );
  AOI22_X1 U10993 ( .A1(n9970), .A2(n9961), .B1(n9983), .B2(n9968), .ZN(
        P2_U3420) );
  INV_X1 U10994 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9969) );
  NOR2_X1 U10995 ( .A1(n9963), .A2(n9962), .ZN(n9965) );
  AOI211_X1 U10996 ( .C1(n9967), .C2(n9966), .A(n9965), .B(n9964), .ZN(n9985)
         );
  AOI22_X1 U10997 ( .A1(n9970), .A2(n9969), .B1(n9985), .B2(n9968), .ZN(
        P2_U3423) );
  INV_X1 U10998 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U10999 ( .A1(n9986), .A2(n9972), .B1(n9971), .B2(n9984), .ZN(
        P2_U3460) );
  AOI22_X1 U11000 ( .A1(n9986), .A2(n9973), .B1(n6902), .B2(n9984), .ZN(
        P2_U3461) );
  INV_X1 U11001 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n9974) );
  AOI22_X1 U11002 ( .A1(n9986), .A2(n9975), .B1(n9974), .B2(n9984), .ZN(
        P2_U3462) );
  AOI22_X1 U11003 ( .A1(n9986), .A2(n9976), .B1(n6973), .B2(n9984), .ZN(
        P2_U3463) );
  AOI22_X1 U11004 ( .A1(n9986), .A2(n9977), .B1(n5913), .B2(n9984), .ZN(
        P2_U3464) );
  AOI22_X1 U11005 ( .A1(n9986), .A2(n9978), .B1(n7235), .B2(n9984), .ZN(
        P2_U3465) );
  INV_X1 U11006 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n9979) );
  AOI22_X1 U11007 ( .A1(n9986), .A2(n9980), .B1(n9979), .B2(n9984), .ZN(
        P2_U3466) );
  AOI22_X1 U11008 ( .A1(n9986), .A2(n9981), .B1(n5954), .B2(n9984), .ZN(
        P2_U3467) );
  AOI22_X1 U11009 ( .A1(n9986), .A2(n9982), .B1(n5970), .B2(n9984), .ZN(
        P2_U3468) );
  AOI22_X1 U11010 ( .A1(n9986), .A2(n9983), .B1(n8452), .B2(n9984), .ZN(
        P2_U3469) );
  AOI22_X1 U11011 ( .A1(n9986), .A2(n9985), .B1(n5998), .B2(n9984), .ZN(
        P2_U3470) );
  NAND3_X1 U11012 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n9989) );
  AND2_X1 U11013 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .ZN(n9987) );
  NOR2_X1 U11014 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n9987), .ZN(n9988) );
  INV_X1 U11015 ( .A(n9988), .ZN(n10005) );
  NAND2_X1 U11016 ( .A1(n9990), .A2(n9989), .ZN(n10004) );
  OAI222_X1 U11017 ( .A1(n9990), .A2(n9989), .B1(n9990), .B2(n10005), .C1(
        n9988), .C2(n10004), .ZN(ADD_1068_U5) );
  XOR2_X1 U11018 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  INV_X1 U11019 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10224) );
  NOR2_X1 U11020 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9991) );
  AOI21_X1 U11021 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9991), .ZN(n10012) );
  NOR2_X1 U11022 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9992) );
  AOI21_X1 U11023 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9992), .ZN(n10015) );
  NOR2_X1 U11024 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9993) );
  AOI21_X1 U11025 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9993), .ZN(n10018) );
  NOR2_X1 U11026 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9994) );
  AOI21_X1 U11027 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9994), .ZN(n10021) );
  NOR2_X1 U11028 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9995) );
  AOI21_X1 U11029 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9995), .ZN(n10024) );
  NOR2_X1 U11030 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9996) );
  AOI21_X1 U11031 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9996), .ZN(n10027) );
  NOR2_X1 U11032 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n9997) );
  AOI21_X1 U11033 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9997), .ZN(n10030) );
  NOR2_X1 U11034 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n9998) );
  AOI21_X1 U11035 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9998), .ZN(n10033) );
  NOR2_X1 U11036 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n9999) );
  AOI21_X1 U11037 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n9999), .ZN(n10236) );
  NOR2_X1 U11038 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n10000) );
  AOI21_X1 U11039 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n10000), .ZN(n10239) );
  NOR2_X1 U11040 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n10001) );
  AOI21_X1 U11041 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n10001), .ZN(n10242) );
  NOR2_X1 U11042 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n10002) );
  AOI21_X1 U11043 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n10002), .ZN(n10245) );
  NOR2_X1 U11044 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(P2_ADDR_REG_5__SCAN_IN), 
        .ZN(n10003) );
  AOI21_X1 U11045 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10003), .ZN(n10248) );
  NAND2_X1 U11046 ( .A1(n10005), .A2(n10004), .ZN(n10233) );
  NAND2_X1 U11047 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10006) );
  OAI21_X1 U11048 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n10006), .ZN(n10232) );
  NOR2_X1 U11049 ( .A1(n10233), .A2(n10232), .ZN(n10231) );
  AOI21_X1 U11050 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10231), .ZN(n10251) );
  NAND2_X1 U11051 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n10007) );
  OAI21_X1 U11052 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10007), .ZN(n10250) );
  NOR2_X1 U11053 ( .A1(n10251), .A2(n10250), .ZN(n10249) );
  AOI21_X1 U11054 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n10249), .ZN(n10254) );
  NOR2_X1 U11055 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10008) );
  AOI21_X1 U11056 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n10008), .ZN(n10253) );
  NAND2_X1 U11057 ( .A1(n10254), .A2(n10253), .ZN(n10252) );
  OAI21_X1 U11058 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10252), .ZN(n10247) );
  NAND2_X1 U11059 ( .A1(n10248), .A2(n10247), .ZN(n10246) );
  OAI21_X1 U11060 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n10246), .ZN(n10244) );
  NAND2_X1 U11061 ( .A1(n10245), .A2(n10244), .ZN(n10243) );
  OAI21_X1 U11062 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10243), .ZN(n10241) );
  NAND2_X1 U11063 ( .A1(n10242), .A2(n10241), .ZN(n10240) );
  OAI21_X1 U11064 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10240), .ZN(n10238) );
  NAND2_X1 U11065 ( .A1(n10239), .A2(n10238), .ZN(n10237) );
  OAI21_X1 U11066 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10237), .ZN(n10235) );
  NAND2_X1 U11067 ( .A1(n10236), .A2(n10235), .ZN(n10234) );
  OAI21_X1 U11068 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10234), .ZN(n10032) );
  NAND2_X1 U11069 ( .A1(n10033), .A2(n10032), .ZN(n10031) );
  OAI21_X1 U11070 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10031), .ZN(n10029) );
  NAND2_X1 U11071 ( .A1(n10030), .A2(n10029), .ZN(n10028) );
  OAI21_X1 U11072 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10028), .ZN(n10026) );
  NAND2_X1 U11073 ( .A1(n10027), .A2(n10026), .ZN(n10025) );
  OAI21_X1 U11074 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10025), .ZN(n10023) );
  NAND2_X1 U11075 ( .A1(n10024), .A2(n10023), .ZN(n10022) );
  OAI21_X1 U11076 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10022), .ZN(n10020) );
  NAND2_X1 U11077 ( .A1(n10021), .A2(n10020), .ZN(n10019) );
  OAI21_X1 U11078 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10019), .ZN(n10017) );
  NAND2_X1 U11079 ( .A1(n10018), .A2(n10017), .ZN(n10016) );
  OAI21_X1 U11080 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10016), .ZN(n10014) );
  NAND2_X1 U11081 ( .A1(n10015), .A2(n10014), .ZN(n10013) );
  OAI21_X1 U11082 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10013), .ZN(n10011) );
  NAND2_X1 U11083 ( .A1(n10012), .A2(n10011), .ZN(n10010) );
  OAI21_X1 U11084 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10010), .ZN(n10223) );
  NOR2_X1 U11085 ( .A1(n10224), .A2(n10223), .ZN(n10225) );
  AOI21_X1 U11086 ( .B1(n10224), .B2(n10223), .A(n10225), .ZN(n10009) );
  XOR2_X1 U11087 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n10009), .Z(ADD_1068_U55)
         );
  OAI21_X1 U11088 ( .B1(n10012), .B2(n10011), .A(n10010), .ZN(ADD_1068_U56) );
  OAI21_X1 U11089 ( .B1(n10015), .B2(n10014), .A(n10013), .ZN(ADD_1068_U57) );
  OAI21_X1 U11090 ( .B1(n10018), .B2(n10017), .A(n10016), .ZN(ADD_1068_U58) );
  OAI21_X1 U11091 ( .B1(n10021), .B2(n10020), .A(n10019), .ZN(ADD_1068_U59) );
  OAI21_X1 U11092 ( .B1(n10024), .B2(n10023), .A(n10022), .ZN(ADD_1068_U60) );
  OAI21_X1 U11093 ( .B1(n10027), .B2(n10026), .A(n10025), .ZN(ADD_1068_U61) );
  OAI21_X1 U11094 ( .B1(n10030), .B2(n10029), .A(n10028), .ZN(ADD_1068_U62) );
  OAI21_X1 U11095 ( .B1(n10033), .B2(n10032), .A(n10031), .ZN(ADD_1068_U63) );
  XOR2_X1 U11096 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(P2_ADDR_REG_19__SCAN_IN), 
        .Z(n10230) );
  AOI22_X1 U11097 ( .A1(SI_18_), .A2(keyinput_f14), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .ZN(n10034) );
  OAI221_X1 U11098 ( .B1(SI_18_), .B2(keyinput_f14), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_f46), .A(n10034), .ZN(n10041)
         );
  AOI22_X1 U11099 ( .A1(SI_1_), .A2(keyinput_f31), .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_f37), .ZN(n10035) );
  OAI221_X1 U11100 ( .B1(SI_1_), .B2(keyinput_f31), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_f37), .A(n10035), .ZN(n10040)
         );
  AOI22_X1 U11101 ( .A1(SI_21_), .A2(keyinput_f11), .B1(P2_RD_REG_SCAN_IN), 
        .B2(keyinput_f33), .ZN(n10036) );
  OAI221_X1 U11102 ( .B1(SI_21_), .B2(keyinput_f11), .C1(P2_RD_REG_SCAN_IN), 
        .C2(keyinput_f33), .A(n10036), .ZN(n10039) );
  AOI22_X1 U11103 ( .A1(SI_8_), .A2(keyinput_f24), .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .ZN(n10037) );
  OAI221_X1 U11104 ( .B1(SI_8_), .B2(keyinput_f24), .C1(
        P2_REG3_REG_24__SCAN_IN), .C2(keyinput_f51), .A(n10037), .ZN(n10038)
         );
  NOR4_X1 U11105 ( .A1(n10041), .A2(n10040), .A3(n10039), .A4(n10038), .ZN(
        n10069) );
  XNOR2_X1 U11106 ( .A(SI_24_), .B(keyinput_f8), .ZN(n10049) );
  AOI22_X1 U11107 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(keyinput_f58), .B1(
        n10043), .B2(keyinput_f38), .ZN(n10042) );
  OAI221_X1 U11108 ( .B1(P2_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .C1(
        n10043), .C2(keyinput_f38), .A(n10042), .ZN(n10048) );
  AOI22_X1 U11109 ( .A1(SI_6_), .A2(keyinput_f26), .B1(SI_25_), .B2(
        keyinput_f7), .ZN(n10044) );
  OAI221_X1 U11110 ( .B1(SI_6_), .B2(keyinput_f26), .C1(SI_25_), .C2(
        keyinput_f7), .A(n10044), .ZN(n10047) );
  AOI22_X1 U11111 ( .A1(SI_31_), .A2(keyinput_f1), .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .ZN(n10045) );
  OAI221_X1 U11112 ( .B1(SI_31_), .B2(keyinput_f1), .C1(
        P2_REG3_REG_10__SCAN_IN), .C2(keyinput_f39), .A(n10045), .ZN(n10046)
         );
  NOR4_X1 U11113 ( .A1(n10049), .A2(n10048), .A3(n10047), .A4(n10046), .ZN(
        n10068) );
  AOI22_X1 U11114 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_f44), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .ZN(n10050) );
  OAI221_X1 U11115 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .C1(
        P2_REG3_REG_3__SCAN_IN), .C2(keyinput_f40), .A(n10050), .ZN(n10057) );
  AOI22_X1 U11116 ( .A1(SI_0_), .A2(keyinput_f32), .B1(SI_20_), .B2(
        keyinput_f12), .ZN(n10051) );
  OAI221_X1 U11117 ( .B1(SI_0_), .B2(keyinput_f32), .C1(SI_20_), .C2(
        keyinput_f12), .A(n10051), .ZN(n10056) );
  AOI22_X1 U11118 ( .A1(SI_3_), .A2(keyinput_f29), .B1(P2_STATE_REG_SCAN_IN), 
        .B2(keyinput_f34), .ZN(n10052) );
  OAI221_X1 U11119 ( .B1(SI_3_), .B2(keyinput_f29), .C1(P2_STATE_REG_SCAN_IN), 
        .C2(keyinput_f34), .A(n10052), .ZN(n10055) );
  AOI22_X1 U11120 ( .A1(SI_23_), .A2(keyinput_f9), .B1(SI_28_), .B2(
        keyinput_f4), .ZN(n10053) );
  OAI221_X1 U11121 ( .B1(SI_23_), .B2(keyinput_f9), .C1(SI_28_), .C2(
        keyinput_f4), .A(n10053), .ZN(n10054) );
  NOR4_X1 U11122 ( .A1(n10057), .A2(n10056), .A3(n10055), .A4(n10054), .ZN(
        n10067) );
  AOI22_X1 U11123 ( .A1(SI_11_), .A2(keyinput_f21), .B1(SI_27_), .B2(
        keyinput_f5), .ZN(n10058) );
  OAI221_X1 U11124 ( .B1(SI_11_), .B2(keyinput_f21), .C1(SI_27_), .C2(
        keyinput_f5), .A(n10058), .ZN(n10065) );
  AOI22_X1 U11125 ( .A1(P2_REG3_REG_18__SCAN_IN), .A2(keyinput_f60), .B1(
        P2_REG3_REG_26__SCAN_IN), .B2(keyinput_f62), .ZN(n10059) );
  OAI221_X1 U11126 ( .B1(P2_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_f62), .A(n10059), .ZN(n10064)
         );
  AOI22_X1 U11127 ( .A1(SI_2_), .A2(keyinput_f30), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(keyinput_f61), .ZN(n10060) );
  OAI221_X1 U11128 ( .B1(SI_2_), .B2(keyinput_f30), .C1(P2_REG3_REG_6__SCAN_IN), .C2(keyinput_f61), .A(n10060), .ZN(n10063) );
  AOI22_X1 U11129 ( .A1(SI_30_), .A2(keyinput_f2), .B1(SI_16_), .B2(
        keyinput_f16), .ZN(n10061) );
  OAI221_X1 U11130 ( .B1(SI_30_), .B2(keyinput_f2), .C1(SI_16_), .C2(
        keyinput_f16), .A(n10061), .ZN(n10062) );
  NOR4_X1 U11131 ( .A1(n10065), .A2(n10064), .A3(n10063), .A4(n10062), .ZN(
        n10066) );
  NAND4_X1 U11132 ( .A1(n10069), .A2(n10068), .A3(n10067), .A4(n10066), .ZN(
        n10120) );
  INV_X1 U11133 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n10150) );
  AOI22_X1 U11134 ( .A1(n6020), .A2(keyinput_f56), .B1(n10150), .B2(
        keyinput_f41), .ZN(n10070) );
  OAI221_X1 U11135 ( .B1(n6020), .B2(keyinput_f56), .C1(n10150), .C2(
        keyinput_f41), .A(n10070), .ZN(n10079) );
  AOI22_X1 U11136 ( .A1(n10143), .A2(keyinput_f6), .B1(keyinput_f20), .B2(
        n10072), .ZN(n10071) );
  OAI221_X1 U11137 ( .B1(n10143), .B2(keyinput_f6), .C1(n10072), .C2(
        keyinput_f20), .A(n10071), .ZN(n10078) );
  AOI22_X1 U11138 ( .A1(n5900), .A2(keyinput_f52), .B1(keyinput_f15), .B2(
        n10074), .ZN(n10073) );
  OAI221_X1 U11139 ( .B1(n5900), .B2(keyinput_f52), .C1(n10074), .C2(
        keyinput_f15), .A(n10073), .ZN(n10077) );
  AOI22_X1 U11140 ( .A1(n10124), .A2(keyinput_f55), .B1(n7968), .B2(
        keyinput_f42), .ZN(n10075) );
  OAI221_X1 U11141 ( .B1(n10124), .B2(keyinput_f55), .C1(n7968), .C2(
        keyinput_f42), .A(n10075), .ZN(n10076) );
  NOR4_X1 U11142 ( .A1(n10079), .A2(n10078), .A3(n10077), .A4(n10076), .ZN(
        n10118) );
  AOI22_X1 U11143 ( .A1(n10082), .A2(keyinput_f54), .B1(n10081), .B2(
        keyinput_f18), .ZN(n10080) );
  OAI221_X1 U11144 ( .B1(n10082), .B2(keyinput_f54), .C1(n10081), .C2(
        keyinput_f18), .A(n10080), .ZN(n10091) );
  AOI22_X1 U11145 ( .A1(SI_10_), .A2(keyinput_f22), .B1(n10171), .B2(
        keyinput_f23), .ZN(n10083) );
  OAI221_X1 U11146 ( .B1(SI_10_), .B2(keyinput_f22), .C1(n10171), .C2(
        keyinput_f23), .A(n10083), .ZN(n10090) );
  INV_X1 U11147 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10085) );
  AOI22_X1 U11148 ( .A1(n10085), .A2(keyinput_f50), .B1(keyinput_f17), .B2(
        n4976), .ZN(n10084) );
  OAI221_X1 U11149 ( .B1(n10085), .B2(keyinput_f50), .C1(n4976), .C2(
        keyinput_f17), .A(n10084), .ZN(n10089) );
  AOI22_X1 U11150 ( .A1(n10149), .A2(keyinput_f63), .B1(keyinput_f10), .B2(
        n10087), .ZN(n10086) );
  OAI221_X1 U11151 ( .B1(n10149), .B2(keyinput_f63), .C1(n10087), .C2(
        keyinput_f10), .A(n10086), .ZN(n10088) );
  NOR4_X1 U11152 ( .A1(n10091), .A2(n10090), .A3(n10089), .A4(n10088), .ZN(
        n10117) );
  INV_X1 U11153 ( .A(P2_WR_REG_SCAN_IN), .ZN(n10152) );
  AOI22_X1 U11154 ( .A1(n10127), .A2(keyinput_f35), .B1(keyinput_f0), .B2(
        n10152), .ZN(n10092) );
  OAI221_X1 U11155 ( .B1(n10127), .B2(keyinput_f35), .C1(n10152), .C2(
        keyinput_f0), .A(n10092), .ZN(n10102) );
  INV_X1 U11156 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10094) );
  AOI22_X1 U11157 ( .A1(n10095), .A2(keyinput_f43), .B1(n10094), .B2(
        keyinput_f45), .ZN(n10093) );
  OAI221_X1 U11158 ( .B1(n10095), .B2(keyinput_f43), .C1(n10094), .C2(
        keyinput_f45), .A(n10093), .ZN(n10101) );
  XNOR2_X1 U11159 ( .A(SI_7_), .B(keyinput_f25), .ZN(n10099) );
  XNOR2_X1 U11160 ( .A(SI_4_), .B(keyinput_f28), .ZN(n10098) );
  XNOR2_X1 U11161 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_f59), .ZN(n10097)
         );
  XNOR2_X1 U11162 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_f47), .ZN(n10096)
         );
  NAND4_X1 U11163 ( .A1(n10099), .A2(n10098), .A3(n10097), .A4(n10096), .ZN(
        n10100) );
  NOR3_X1 U11164 ( .A1(n10102), .A2(n10101), .A3(n10100), .ZN(n10116) );
  INV_X1 U11165 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U11166 ( .A1(n10153), .A2(keyinput_f36), .B1(keyinput_f13), .B2(
        n10104), .ZN(n10103) );
  OAI221_X1 U11167 ( .B1(n10153), .B2(keyinput_f36), .C1(n10104), .C2(
        keyinput_f13), .A(n10103), .ZN(n10114) );
  AOI22_X1 U11168 ( .A1(n10168), .A2(keyinput_f49), .B1(keyinput_f3), .B2(
        n6207), .ZN(n10105) );
  OAI221_X1 U11169 ( .B1(n10168), .B2(keyinput_f49), .C1(n6207), .C2(
        keyinput_f3), .A(n10105), .ZN(n10113) );
  AOI22_X1 U11170 ( .A1(n10107), .A2(keyinput_f57), .B1(keyinput_f19), .B2(
        n10156), .ZN(n10106) );
  OAI221_X1 U11171 ( .B1(n10107), .B2(keyinput_f57), .C1(n10156), .C2(
        keyinput_f19), .A(n10106), .ZN(n10112) );
  AOI22_X1 U11172 ( .A1(n10110), .A2(keyinput_f27), .B1(n10109), .B2(
        keyinput_f48), .ZN(n10108) );
  OAI221_X1 U11173 ( .B1(n10110), .B2(keyinput_f27), .C1(n10109), .C2(
        keyinput_f48), .A(n10108), .ZN(n10111) );
  NOR4_X1 U11174 ( .A1(n10114), .A2(n10113), .A3(n10112), .A4(n10111), .ZN(
        n10115) );
  NAND4_X1 U11175 ( .A1(n10118), .A2(n10117), .A3(n10116), .A4(n10115), .ZN(
        n10119) );
  OAI22_X1 U11176 ( .A1(n10120), .A2(n10119), .B1(keyinput_f53), .B2(
        P2_REG3_REG_9__SCAN_IN), .ZN(n10121) );
  AOI21_X1 U11177 ( .B1(keyinput_f53), .B2(P2_REG3_REG_9__SCAN_IN), .A(n10121), 
        .ZN(n10221) );
  AOI22_X1 U11178 ( .A1(n10124), .A2(keyinput_g55), .B1(keyinput_g16), .B2(
        n10123), .ZN(n10122) );
  OAI221_X1 U11179 ( .B1(n10124), .B2(keyinput_g55), .C1(n10123), .C2(
        keyinput_g16), .A(n10122), .ZN(n10137) );
  AOI22_X1 U11180 ( .A1(n10127), .A2(keyinput_g35), .B1(keyinput_g12), .B2(
        n10126), .ZN(n10125) );
  OAI221_X1 U11181 ( .B1(n10127), .B2(keyinput_g35), .C1(n10126), .C2(
        keyinput_g12), .A(n10125), .ZN(n10136) );
  INV_X1 U11182 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10130) );
  AOI22_X1 U11183 ( .A1(n10130), .A2(keyinput_g51), .B1(keyinput_g37), .B2(
        n10129), .ZN(n10128) );
  OAI221_X1 U11184 ( .B1(n10130), .B2(keyinput_g51), .C1(n10129), .C2(
        keyinput_g37), .A(n10128), .ZN(n10135) );
  INV_X1 U11185 ( .A(P2_RD_REG_SCAN_IN), .ZN(n10131) );
  XOR2_X1 U11186 ( .A(n10131), .B(keyinput_g33), .Z(n10133) );
  XNOR2_X1 U11187 ( .A(SI_4_), .B(keyinput_g28), .ZN(n10132) );
  NAND2_X1 U11188 ( .A1(n10133), .A2(n10132), .ZN(n10134) );
  NOR4_X1 U11189 ( .A1(n10137), .A2(n10136), .A3(n10135), .A4(n10134), .ZN(
        n10181) );
  AOI22_X1 U11190 ( .A1(SI_0_), .A2(keyinput_g32), .B1(SI_29_), .B2(
        keyinput_g3), .ZN(n10138) );
  OAI221_X1 U11191 ( .B1(SI_0_), .B2(keyinput_g32), .C1(SI_29_), .C2(
        keyinput_g3), .A(n10138), .ZN(n10147) );
  AOI22_X1 U11192 ( .A1(P2_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(
        P2_REG3_REG_8__SCAN_IN), .B2(keyinput_g43), .ZN(n10139) );
  OAI221_X1 U11193 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(
        P2_REG3_REG_8__SCAN_IN), .C2(keyinput_g43), .A(n10139), .ZN(n10146) );
  AOI22_X1 U11194 ( .A1(n5900), .A2(keyinput_g52), .B1(n10141), .B2(
        keyinput_g46), .ZN(n10140) );
  OAI221_X1 U11195 ( .B1(n5900), .B2(keyinput_g52), .C1(n10141), .C2(
        keyinput_g46), .A(n10140), .ZN(n10145) );
  AOI22_X1 U11196 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(keyinput_g45), .B1(
        n10143), .B2(keyinput_g6), .ZN(n10142) );
  OAI221_X1 U11197 ( .B1(P2_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .C1(
        n10143), .C2(keyinput_g6), .A(n10142), .ZN(n10144) );
  NOR4_X1 U11198 ( .A1(n10147), .A2(n10146), .A3(n10145), .A4(n10144), .ZN(
        n10180) );
  AOI22_X1 U11199 ( .A1(n10150), .A2(keyinput_g41), .B1(keyinput_g63), .B2(
        n10149), .ZN(n10148) );
  OAI221_X1 U11200 ( .B1(n10150), .B2(keyinput_g41), .C1(n10149), .C2(
        keyinput_g63), .A(n10148), .ZN(n10162) );
  AOI22_X1 U11201 ( .A1(n10153), .A2(keyinput_g36), .B1(keyinput_g0), .B2(
        n10152), .ZN(n10151) );
  OAI221_X1 U11202 ( .B1(n10153), .B2(keyinput_g36), .C1(n10152), .C2(
        keyinput_g0), .A(n10151), .ZN(n10161) );
  AOI22_X1 U11203 ( .A1(n10156), .A2(keyinput_g19), .B1(n10155), .B2(
        keyinput_g14), .ZN(n10154) );
  OAI221_X1 U11204 ( .B1(n10156), .B2(keyinput_g19), .C1(n10155), .C2(
        keyinput_g14), .A(n10154), .ZN(n10160) );
  XNOR2_X1 U11205 ( .A(P2_REG3_REG_22__SCAN_IN), .B(keyinput_g57), .ZN(n10158)
         );
  XNOR2_X1 U11206 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_g44), .ZN(n10157)
         );
  NAND2_X1 U11207 ( .A1(n10158), .A2(n10157), .ZN(n10159) );
  NOR4_X1 U11208 ( .A1(n10162), .A2(n10161), .A3(n10160), .A4(n10159), .ZN(
        n10179) );
  INV_X1 U11209 ( .A(SI_6_), .ZN(n10164) );
  AOI22_X1 U11210 ( .A1(n10165), .A2(keyinput_g7), .B1(keyinput_g26), .B2(
        n10164), .ZN(n10163) );
  OAI221_X1 U11211 ( .B1(n10165), .B2(keyinput_g7), .C1(n10164), .C2(
        keyinput_g26), .A(n10163), .ZN(n10177) );
  AOI22_X1 U11212 ( .A1(n10168), .A2(keyinput_g49), .B1(keyinput_g8), .B2(
        n10167), .ZN(n10166) );
  OAI221_X1 U11213 ( .B1(n10168), .B2(keyinput_g49), .C1(n10167), .C2(
        keyinput_g8), .A(n10166), .ZN(n10176) );
  AOI22_X1 U11214 ( .A1(n10171), .A2(keyinput_g23), .B1(n10170), .B2(
        keyinput_g11), .ZN(n10169) );
  OAI221_X1 U11215 ( .B1(n10171), .B2(keyinput_g23), .C1(n10170), .C2(
        keyinput_g11), .A(n10169), .ZN(n10175) );
  XNOR2_X1 U11216 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_g48), .ZN(n10173)
         );
  XNOR2_X1 U11217 ( .A(SI_1_), .B(keyinput_g31), .ZN(n10172) );
  NAND2_X1 U11218 ( .A1(n10173), .A2(n10172), .ZN(n10174) );
  NOR4_X1 U11219 ( .A1(n10177), .A2(n10176), .A3(n10175), .A4(n10174), .ZN(
        n10178) );
  NAND4_X1 U11220 ( .A1(n10181), .A2(n10180), .A3(n10179), .A4(n10178), .ZN(
        n10219) );
  AOI22_X1 U11221 ( .A1(SI_3_), .A2(keyinput_g29), .B1(SI_10_), .B2(
        keyinput_g22), .ZN(n10182) );
  OAI221_X1 U11222 ( .B1(SI_3_), .B2(keyinput_g29), .C1(SI_10_), .C2(
        keyinput_g22), .A(n10182), .ZN(n10189) );
  AOI22_X1 U11223 ( .A1(SI_17_), .A2(keyinput_g15), .B1(SI_28_), .B2(
        keyinput_g4), .ZN(n10183) );
  OAI221_X1 U11224 ( .B1(SI_17_), .B2(keyinput_g15), .C1(SI_28_), .C2(
        keyinput_g4), .A(n10183), .ZN(n10188) );
  AOI22_X1 U11225 ( .A1(SI_11_), .A2(keyinput_g21), .B1(SI_12_), .B2(
        keyinput_g20), .ZN(n10184) );
  OAI221_X1 U11226 ( .B1(SI_11_), .B2(keyinput_g21), .C1(SI_12_), .C2(
        keyinput_g20), .A(n10184), .ZN(n10187) );
  AOI22_X1 U11227 ( .A1(SI_8_), .A2(keyinput_g24), .B1(P2_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .ZN(n10185) );
  OAI221_X1 U11228 ( .B1(SI_8_), .B2(keyinput_g24), .C1(
        P2_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n10185), .ZN(n10186)
         );
  NOR4_X1 U11229 ( .A1(n10189), .A2(n10188), .A3(n10187), .A4(n10186), .ZN(
        n10217) );
  XNOR2_X1 U11230 ( .A(SI_15_), .B(keyinput_g17), .ZN(n10197) );
  AOI22_X1 U11231 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(keyinput_g38), .B1(
        n10191), .B2(keyinput_g58), .ZN(n10190) );
  OAI221_X1 U11232 ( .B1(P2_REG3_REG_23__SCAN_IN), .B2(keyinput_g38), .C1(
        n10191), .C2(keyinput_g58), .A(n10190), .ZN(n10196) );
  AOI22_X1 U11233 ( .A1(SI_14_), .A2(keyinput_g18), .B1(SI_23_), .B2(
        keyinput_g9), .ZN(n10192) );
  OAI221_X1 U11234 ( .B1(SI_14_), .B2(keyinput_g18), .C1(SI_23_), .C2(
        keyinput_g9), .A(n10192), .ZN(n10195) );
  AOI22_X1 U11235 ( .A1(SI_5_), .A2(keyinput_g27), .B1(P2_REG3_REG_26__SCAN_IN), .B2(keyinput_g62), .ZN(n10193) );
  OAI221_X1 U11236 ( .B1(SI_5_), .B2(keyinput_g27), .C1(
        P2_REG3_REG_26__SCAN_IN), .C2(keyinput_g62), .A(n10193), .ZN(n10194)
         );
  NOR4_X1 U11237 ( .A1(n10197), .A2(n10196), .A3(n10195), .A4(n10194), .ZN(
        n10216) );
  AOI22_X1 U11238 ( .A1(SI_27_), .A2(keyinput_g5), .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_g39), .ZN(n10198) );
  OAI221_X1 U11239 ( .B1(SI_27_), .B2(keyinput_g5), .C1(
        P2_REG3_REG_10__SCAN_IN), .C2(keyinput_g39), .A(n10198), .ZN(n10205)
         );
  AOI22_X1 U11240 ( .A1(SI_22_), .A2(keyinput_g10), .B1(P2_STATE_REG_SCAN_IN), 
        .B2(keyinput_g34), .ZN(n10199) );
  OAI221_X1 U11241 ( .B1(SI_22_), .B2(keyinput_g10), .C1(P2_STATE_REG_SCAN_IN), 
        .C2(keyinput_g34), .A(n10199), .ZN(n10204) );
  AOI22_X1 U11242 ( .A1(SI_2_), .A2(keyinput_g30), .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .ZN(n10200) );
  OAI221_X1 U11243 ( .B1(SI_2_), .B2(keyinput_g30), .C1(
        P2_REG3_REG_13__SCAN_IN), .C2(keyinput_g56), .A(n10200), .ZN(n10203)
         );
  AOI22_X1 U11244 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_g40), .B1(
        P2_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .ZN(n10201) );
  OAI221_X1 U11245 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_g40), .C1(
        P2_REG3_REG_25__SCAN_IN), .C2(keyinput_g47), .A(n10201), .ZN(n10202)
         );
  NOR4_X1 U11246 ( .A1(n10205), .A2(n10204), .A3(n10203), .A4(n10202), .ZN(
        n10215) );
  AOI22_X1 U11247 ( .A1(SI_30_), .A2(keyinput_g2), .B1(SI_31_), .B2(
        keyinput_g1), .ZN(n10206) );
  OAI221_X1 U11248 ( .B1(SI_30_), .B2(keyinput_g2), .C1(SI_31_), .C2(
        keyinput_g1), .A(n10206), .ZN(n10213) );
  AOI22_X1 U11249 ( .A1(SI_7_), .A2(keyinput_g25), .B1(P2_REG3_REG_6__SCAN_IN), 
        .B2(keyinput_g61), .ZN(n10207) );
  OAI221_X1 U11250 ( .B1(SI_7_), .B2(keyinput_g25), .C1(P2_REG3_REG_6__SCAN_IN), .C2(keyinput_g61), .A(n10207), .ZN(n10212) );
  AOI22_X1 U11251 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(keyinput_g50), .B1(
        P2_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n10208) );
  OAI221_X1 U11252 ( .B1(P2_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .C1(
        P2_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n10208), .ZN(n10211)
         );
  AOI22_X1 U11253 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_g59), .B1(SI_19_), .B2(keyinput_g13), .ZN(n10209) );
  OAI221_X1 U11254 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_g59), .C1(
        SI_19_), .C2(keyinput_g13), .A(n10209), .ZN(n10210) );
  NOR4_X1 U11255 ( .A1(n10213), .A2(n10212), .A3(n10211), .A4(n10210), .ZN(
        n10214) );
  NAND4_X1 U11256 ( .A1(n10217), .A2(n10216), .A3(n10215), .A4(n10214), .ZN(
        n10218) );
  OAI22_X1 U11257 ( .A1(keyinput_g53), .A2(n10222), .B1(n10219), .B2(n10218), 
        .ZN(n10220) );
  AOI211_X1 U11258 ( .C1(keyinput_g53), .C2(n10222), .A(n10221), .B(n10220), 
        .ZN(n10228) );
  NAND2_X1 U11259 ( .A1(n10224), .A2(n10223), .ZN(n10226) );
  AOI21_X1 U11260 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(n10226), .A(n10225), 
        .ZN(n10227) );
  XOR2_X1 U11261 ( .A(n10228), .B(n10227), .Z(n10229) );
  XNOR2_X1 U11262 ( .A(n10230), .B(n10229), .ZN(ADD_1068_U4) );
  AOI21_X1 U11263 ( .B1(n10233), .B2(n10232), .A(n10231), .ZN(ADD_1068_U54) );
  OAI21_X1 U11264 ( .B1(n10236), .B2(n10235), .A(n10234), .ZN(ADD_1068_U47) );
  OAI21_X1 U11265 ( .B1(n10239), .B2(n10238), .A(n10237), .ZN(ADD_1068_U48) );
  OAI21_X1 U11266 ( .B1(n10242), .B2(n10241), .A(n10240), .ZN(ADD_1068_U49) );
  OAI21_X1 U11267 ( .B1(n10245), .B2(n10244), .A(n10243), .ZN(ADD_1068_U50) );
  OAI21_X1 U11268 ( .B1(n10248), .B2(n10247), .A(n10246), .ZN(ADD_1068_U51) );
  AOI21_X1 U11269 ( .B1(n10251), .B2(n10250), .A(n10249), .ZN(ADD_1068_U53) );
  OAI21_X1 U11270 ( .B1(n10254), .B2(n10253), .A(n10252), .ZN(ADD_1068_U52) );
  NOR2_X1 U4862 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6437) );
  INV_X1 U4903 ( .A(n5213), .ZN(n6491) );
endmodule

