

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput63, keyinput62, 
        keyinput61, keyinput60, keyinput59, keyinput58, keyinput57, keyinput56, 
        keyinput55, keyinput54, keyinput53, keyinput52, keyinput51, keyinput50, 
        keyinput49, keyinput48, keyinput47, keyinput46, keyinput45, keyinput44, 
        keyinput43, keyinput42, keyinput41, keyinput40, keyinput39, keyinput38, 
        keyinput37, keyinput36, keyinput35, keyinput34, keyinput33, keyinput32, 
        keyinput31, keyinput30, keyinput29, keyinput28, keyinput27, keyinput26, 
        keyinput25, keyinput24, keyinput23, keyinput22, keyinput21, keyinput20, 
        keyinput19, keyinput18, keyinput17, keyinput16, keyinput15, keyinput14, 
        keyinput13, keyinput12, keyinput11, keyinput10, keyinput9, keyinput8, 
        keyinput7, keyinput6, keyinput5, keyinput4, keyinput3, keyinput2, 
        keyinput1, keyinput0 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080;

  INV_X4 U4754 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NAND2_X1 U4755 ( .A1(n4371), .A2(n4983), .ZN(n8017) );
  INV_X2 U4756 ( .A(n4816), .ZN(n4260) );
  AND4_X1 U4757 ( .A1(n5541), .A2(n5540), .A3(n5539), .A4(n5538), .ZN(n7669)
         );
  INV_X2 U4758 ( .A(n5535), .ZN(n5620) );
  INV_X1 U4759 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5878) );
  AND2_X1 U4760 ( .A1(n5319), .A2(n5320), .ZN(n8027) );
  INV_X1 U4761 ( .A(n4814), .ZN(n7897) );
  INV_X1 U4762 ( .A(n6613), .ZN(n4547) );
  NAND2_X1 U4763 ( .A1(n4724), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4725) );
  INV_X1 U4764 ( .A(n5537), .ZN(n7417) );
  NOR2_X1 U4765 ( .A1(n9542), .A2(n9541), .ZN(n9540) );
  XNOR2_X1 U4766 ( .A(n7390), .B(n7389), .ZN(n7414) );
  OAI211_X1 U4767 ( .C1(n5997), .C2(n8338), .A(n4783), .B(n4782), .ZN(n9793)
         );
  OAI21_X1 U4768 ( .B1(n4425), .B2(n5878), .A(n5522), .ZN(n4424) );
  INV_X1 U4769 ( .A(n8511), .ZN(n4764) );
  AND2_X1 U4770 ( .A1(n6701), .A2(n8136), .ZN(n4249) );
  AND2_X1 U4771 ( .A1(n4946), .A2(n4928), .ZN(n4250) );
  AND2_X1 U4772 ( .A1(n6300), .A2(n5533), .ZN(n4251) );
  BUF_X4 U4773 ( .A(n5843), .Z(n4252) );
  INV_X1 U4774 ( .A(n5549), .ZN(n5843) );
  AOI21_X2 U4775 ( .B1(n6956), .B2(n6955), .A(n6954), .ZN(n7088) );
  NAND2_X2 U4776 ( .A1(n6761), .A2(n8134), .ZN(n6956) );
  AND2_X4 U4777 ( .A1(n5882), .A2(n5881), .ZN(n7663) );
  OAI21_X2 U4779 ( .B1(n4645), .B2(n4644), .A(n4266), .ZN(n4984) );
  OR2_X1 U4780 ( .A1(n9861), .A2(n8511), .ZN(n4253) );
  OR2_X1 U4781 ( .A1(n9861), .A2(n8511), .ZN(n4254) );
  NAND2_X2 U4782 ( .A1(n6528), .A2(n5628), .ZN(n9645) );
  NOR2_X2 U4783 ( .A1(n5761), .A2(n5760), .ZN(n5788) );
  NAND2_X2 U4784 ( .A1(n5775), .A2(n5774), .ZN(n9334) );
  OR2_X2 U4785 ( .A1(n4745), .A2(n4737), .ZN(n4747) );
  NAND2_X4 U4786 ( .A1(n4376), .A2(n6684), .ZN(n5410) );
  XNOR2_X2 U4787 ( .A(n5041), .B(n5040), .ZN(n6128) );
  NAND2_X2 U4788 ( .A1(n4676), .A2(n4674), .ZN(n5041) );
  XNOR2_X2 U4789 ( .A(n5532), .B(n7664), .ZN(n6302) );
  XNOR2_X2 U4791 ( .A(n7396), .B(n7395), .ZN(n8109) );
  AOI211_X2 U4792 ( .C1(n9654), .C2(n9162), .A(n9131), .B(n9130), .ZN(n9306)
         );
  OR2_X1 U4793 ( .A1(n8750), .A2(n8462), .ZN(n8264) );
  OAI21_X1 U4794 ( .B1(n8917), .B2(n6480), .A(n6479), .ZN(n6483) );
  CLKBUF_X2 U4795 ( .A(P1_U4006), .Z(n4257) );
  CLKBUF_X2 U4796 ( .A(n4802), .Z(n4259) );
  AND4_X1 U4797 ( .A1(n5556), .A2(n5555), .A3(n5554), .A4(n5553), .ZN(n6432)
         );
  AND2_X1 U4798 ( .A1(n7950), .A2(n4728), .ZN(n4802) );
  INV_X4 U4799 ( .A(n5534), .ZN(n5580) );
  NAND2_X1 U4800 ( .A1(n4424), .A2(n4423), .ZN(n9010) );
  INV_X1 U4801 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4425) );
  INV_X2 U4802 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NOR2_X1 U4803 ( .A1(n4342), .A2(n7653), .ZN(n7658) );
  INV_X1 U4804 ( .A(n4343), .ZN(n4342) );
  NOR4_X2 U4805 ( .A1(n8298), .A2(n8297), .A3(n8296), .A4(n8295), .ZN(n8299)
         );
  INV_X1 U4806 ( .A(n7517), .ZN(n7694) );
  INV_X1 U4807 ( .A(n7457), .ZN(n9280) );
  AND2_X1 U4808 ( .A1(n7413), .A2(n7412), .ZN(n7457) );
  AOI21_X1 U4809 ( .B1(n8486), .B2(n4285), .A(n4665), .ZN(n8116) );
  INV_X1 U4810 ( .A(n9287), .ZN(n9069) );
  AND2_X1 U4811 ( .A1(n7416), .A2(n7415), .ZN(n9287) );
  NAND2_X1 U4812 ( .A1(n4501), .A2(n4496), .ZN(n4499) );
  AOI21_X1 U4813 ( .B1(n4279), .B2(n7631), .A(n4333), .ZN(n4332) );
  XNOR2_X1 U4814 ( .A(n7414), .B(SI_30_), .ZN(n8107) );
  NAND2_X1 U4815 ( .A1(n7387), .A2(n7386), .ZN(n7390) );
  OR2_X1 U4816 ( .A1(n7424), .A2(n7384), .ZN(n7387) );
  NAND2_X1 U4817 ( .A1(n7744), .A2(n4291), .ZN(n8953) );
  NAND2_X1 U4818 ( .A1(n5415), .A2(n5414), .ZN(n7379) );
  NAND2_X1 U4819 ( .A1(n5413), .A2(n5412), .ZN(n5415) );
  NAND2_X1 U4820 ( .A1(n7625), .A2(n7463), .ZN(n9137) );
  OR2_X1 U4821 ( .A1(n7430), .A2(n5900), .ZN(n9185) );
  AOI21_X1 U4822 ( .B1(n5896), .B2(n5895), .A(n5894), .ZN(n9475) );
  NAND2_X1 U4823 ( .A1(n5798), .A2(n5797), .ZN(n9195) );
  NAND2_X1 U4824 ( .A1(n5304), .A2(n5303), .ZN(n5333) );
  NAND2_X1 U4825 ( .A1(n5787), .A2(n5786), .ZN(n9331) );
  NAND2_X1 U4826 ( .A1(n5298), .A2(n5297), .ZN(n5304) );
  OR2_X1 U4827 ( .A1(n6897), .A2(n6987), .ZN(n6898) );
  AND2_X1 U4828 ( .A1(n6988), .A2(n6896), .ZN(n6987) );
  XNOR2_X1 U4829 ( .A(n5211), .B(n5232), .ZN(n6563) );
  NAND2_X1 U4830 ( .A1(n5290), .A2(n5289), .ZN(n5298) );
  NAND2_X1 U4831 ( .A1(n5268), .A2(n5266), .ZN(n5290) );
  AND2_X1 U4832 ( .A1(n5206), .A2(n5233), .ZN(n5211) );
  AND2_X1 U4833 ( .A1(n5134), .A2(n5027), .ZN(n7286) );
  AND2_X1 U4834 ( .A1(n7087), .A2(n6957), .ZN(n7015) );
  NAND2_X1 U4835 ( .A1(n5087), .A2(n5086), .ZN(n7917) );
  OR2_X1 U4836 ( .A1(n7301), .A2(n7300), .ZN(n7869) );
  AND2_X1 U4837 ( .A1(n8173), .A2(n8174), .ZN(n7178) );
  AOI211_X1 U4838 ( .C1(n7919), .C2(n8101), .A(n7296), .B(n7295), .ZN(n7297)
         );
  OR2_X1 U4839 ( .A1(n7170), .A2(n7306), .ZN(n8173) );
  AOI21_X1 U4840 ( .B1(n5060), .B2(n5057), .A(n4703), .ZN(n5077) );
  NAND2_X1 U4841 ( .A1(n5676), .A2(n5675), .ZN(n7038) );
  OR2_X1 U4842 ( .A1(n6642), .A2(n6641), .ZN(n6644) );
  NAND2_X2 U4843 ( .A1(n5660), .A2(n5659), .ZN(n7114) );
  AND2_X1 U4844 ( .A1(n4368), .A2(n4366), .ZN(n8044) );
  INV_X2 U4845 ( .A(n9867), .ZN(n4255) );
  INV_X2 U4846 ( .A(n9884), .ZN(n4256) );
  XNOR2_X1 U4847 ( .A(n5003), .B(n4999), .ZN(n5657) );
  AND2_X1 U4848 ( .A1(n5592), .A2(n5591), .ZN(n9699) );
  NAND2_X1 U4849 ( .A1(n5578), .A2(n4513), .ZN(n6488) );
  OAI211_X1 U4850 ( .C1(n6298), .C2(n6195), .A(n6155), .B(n6154), .ZN(n6157)
         );
  INV_X4 U4851 ( .A(n8121), .ZN(n5409) );
  AND3_X1 U4852 ( .A1(n5575), .A2(n5574), .A3(n5573), .ZN(n9688) );
  NAND4_X1 U4853 ( .A1(n4773), .A2(n4772), .A3(n4771), .A4(n4770), .ZN(n8326)
         );
  CLKBUF_X3 U4854 ( .A(n6197), .Z(n7806) );
  CLKBUF_X1 U4855 ( .A(n4940), .Z(n7899) );
  NAND2_X1 U4856 ( .A1(n6151), .A2(n6176), .ZN(n6613) );
  AND2_X1 U4857 ( .A1(n4763), .A2(n4514), .ZN(n6714) );
  NAND2_X2 U4858 ( .A1(n6177), .A2(n6176), .ZN(n7821) );
  AND3_X1 U4859 ( .A1(n5562), .A2(n5561), .A3(n5560), .ZN(n6496) );
  XNOR2_X1 U4860 ( .A(n4533), .B(n5492), .ZN(n5944) );
  NAND4_X1 U4861 ( .A1(n5569), .A2(n5568), .A3(n5567), .A4(n5566), .ZN(n9005)
         );
  BUF_X1 U4862 ( .A(n5532), .Z(n7665) );
  MUX2_X1 U4863 ( .A(n4375), .B(n8854), .S(n5997), .Z(n9773) );
  AND2_X2 U4864 ( .A1(n4729), .A2(n4728), .ZN(n4814) );
  INV_X1 U4865 ( .A(n6299), .ZN(n6176) );
  AND2_X2 U4866 ( .A1(n7950), .A2(n4726), .ZN(n4816) );
  NAND2_X1 U4867 ( .A1(n4762), .A2(n4761), .ZN(n4952) );
  BUF_X2 U4868 ( .A(n4762), .Z(n5997) );
  XNOR2_X1 U4869 ( .A(n4723), .B(n4722), .ZN(n7950) );
  NAND2_X1 U4870 ( .A1(n5468), .A2(n7904), .ZN(n4762) );
  XNOR2_X1 U4871 ( .A(n5874), .B(n5929), .ZN(n7659) );
  NAND2_X1 U4872 ( .A1(n7397), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4723) );
  XNOR2_X1 U4873 ( .A(n4749), .B(n4748), .ZN(n7904) );
  NAND2_X1 U4874 ( .A1(n5531), .A2(n7393), .ZN(n5613) );
  XNOR2_X1 U4875 ( .A(n4848), .B(SI_4_), .ZN(n4846) );
  NAND2_X2 U4876 ( .A1(n5531), .A2(n4761), .ZN(n7426) );
  AND2_X1 U4877 ( .A1(n5745), .A2(n4569), .ZN(n5945) );
  XNOR2_X1 U4878 ( .A(n4894), .B(SI_6_), .ZN(n4892) );
  NAND2_X1 U4879 ( .A1(n4926), .A2(n4925), .ZN(n4946) );
  XNOR2_X1 U4880 ( .A(n4873), .B(SI_5_), .ZN(n4871) );
  OR2_X1 U4881 ( .A1(n7402), .A2(n5878), .ZN(n5502) );
  INV_X2 U4882 ( .A(n7407), .ZN(n7850) );
  NAND2_X1 U4883 ( .A1(n5503), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5505) );
  NAND2_X1 U4884 ( .A1(n4721), .A2(n5419), .ZN(n5424) );
  INV_X2 U4885 ( .A(n6426), .ZN(n4258) );
  NAND2_X1 U4886 ( .A1(n4301), .A2(n4798), .ZN(n6335) );
  NOR2_X1 U4887 ( .A1(n5494), .A2(n5493), .ZN(n5495) );
  AND4_X1 U4888 ( .A1(n4710), .A2(n4709), .A3(n4896), .A4(n10031), .ZN(n4711)
         );
  AND3_X1 U4889 ( .A1(n4537), .A2(n4536), .A3(n4535), .ZN(n4630) );
  AND2_X1 U4890 ( .A1(n4476), .A2(n4375), .ZN(n4750) );
  NAND3_X1 U4891 ( .A1(n4755), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n4690) );
  INV_X1 U4892 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5543) );
  NOR2_X1 U4893 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n4538) );
  INV_X1 U4894 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5671) );
  INV_X1 U4895 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4737) );
  NOR2_X1 U4896 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5487) );
  INV_X1 U4897 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n4896) );
  INV_X1 U4898 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n4602) );
  INV_X1 U4899 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5929) );
  NOR2_X1 U4900 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n4374) );
  INV_X1 U4901 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n4708) );
  INV_X1 U4902 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5696) );
  NOR2_X1 U4903 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n4536) );
  NOR2_X1 U4904 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4537) );
  NOR2_X1 U4905 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n4535) );
  AOI21_X1 U4906 ( .B1(n9135), .B2(n9137), .A(n5837), .ZN(n9117) );
  AOI21_X2 U4907 ( .B1(n7881), .B2(n7880), .A(n7879), .ZN(n8681) );
  AND2_X2 U4908 ( .A1(n7157), .A2(n8161), .ZN(n7881) );
  OAI21_X2 U4909 ( .B1(n6919), .B2(n6899), .A(n6898), .ZN(n7140) );
  INV_X4 U4910 ( .A(n4781), .ZN(n4761) );
  NAND2_X4 U4911 ( .A1(n5512), .A2(n5506), .ZN(n5535) );
  INV_X2 U4912 ( .A(n7708), .ZN(n5506) );
  OAI222_X1 U4913 ( .A1(P2_U3152), .A2(n5468), .B1(n7319), .B2(n7739), .C1(
        n7318), .C2(n7947), .ZN(P2_U3330) );
  XNOR2_X2 U4914 ( .A(n4747), .B(n4746), .ZN(n5468) );
  OR2_X1 U4915 ( .A1(n8779), .A2(n8096), .ZN(n8241) );
  INV_X1 U4916 ( .A(n5151), .ZN(n5255) );
  NAND2_X1 U4917 ( .A1(n8477), .A2(n7915), .ZN(n8465) );
  NAND2_X1 U4918 ( .A1(n7550), .A2(n7549), .ZN(n7561) );
  NAND2_X1 U4919 ( .A1(n4321), .A2(n7541), .ZN(n7542) );
  AND2_X1 U4920 ( .A1(n7564), .A2(n4327), .ZN(n4326) );
  AND2_X1 U4921 ( .A1(n7569), .A2(n7547), .ZN(n4327) );
  NAND2_X1 U4922 ( .A1(n4608), .A2(n4607), .ZN(n4606) );
  INV_X1 U4923 ( .A(n8187), .ZN(n4608) );
  NAND2_X1 U4924 ( .A1(n4328), .A2(n4332), .ZN(n7638) );
  NAND2_X1 U4925 ( .A1(n7632), .A2(n4279), .ZN(n4328) );
  OR2_X1 U4926 ( .A1(n9289), .A2(n7429), .ZN(n7640) );
  NAND3_X1 U4927 ( .A1(n9772), .A2(n4764), .A3(n5463), .ZN(n4376) );
  NAND2_X1 U4928 ( .A1(n4667), .A2(n8252), .ZN(n4666) );
  OR2_X1 U4929 ( .A1(n8773), .A2(n7954), .ZN(n8252) );
  NOR2_X1 U4930 ( .A1(n8565), .A2(n8556), .ZN(n4689) );
  INV_X1 U4931 ( .A(n8597), .ZN(n4687) );
  OR2_X1 U4932 ( .A1(n8613), .A2(n7984), .ZN(n8214) );
  NAND2_X1 U4933 ( .A1(n5019), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5049) );
  NOR2_X1 U4934 ( .A1(n5013), .A2(n4601), .ZN(n5110) );
  NAND2_X1 U4935 ( .A1(n4300), .A2(n4716), .ZN(n4601) );
  NAND2_X1 U4936 ( .A1(n8939), .A2(n4544), .ZN(n4543) );
  OR2_X1 U4937 ( .A1(n9077), .A2(n8862), .ZN(n7639) );
  OR2_X1 U4938 ( .A1(n6488), .A2(n8922), .ZN(n7535) );
  NAND2_X1 U4939 ( .A1(n8922), .A2(n6488), .ZN(n7534) );
  NAND2_X1 U4940 ( .A1(n7383), .A2(n7382), .ZN(n7424) );
  NAND2_X1 U4941 ( .A1(n7379), .A2(n7378), .ZN(n7383) );
  NAND2_X1 U4942 ( .A1(n5382), .A2(n5381), .ZN(n5413) );
  OAI21_X1 U4943 ( .B1(n5354), .B2(n5353), .A(n5352), .ZN(n5380) );
  NAND2_X1 U4944 ( .A1(n5935), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5937) );
  AND2_X1 U4945 ( .A1(n5233), .A2(n5232), .ZN(n5234) );
  NAND2_X1 U4946 ( .A1(n5108), .A2(n5107), .ZN(n5151) );
  NAND2_X1 U4947 ( .A1(n8044), .A2(n4833), .ZN(n8043) );
  AND2_X1 U4948 ( .A1(n5462), .A2(n5463), .ZN(n8269) );
  AND2_X1 U4949 ( .A1(n5395), .A2(n5394), .ZN(n8096) );
  NAND2_X1 U4950 ( .A1(n8112), .A2(n8111), .ZN(n8459) );
  AND2_X1 U4951 ( .A1(n8548), .A2(n4274), .ZN(n8477) );
  NAND2_X1 U4952 ( .A1(n8617), .A2(n7934), .ZN(n7940) );
  NOR2_X1 U4953 ( .A1(n8641), .A2(n8824), .ZN(n8631) );
  NAND2_X1 U4954 ( .A1(n7075), .A2(n4404), .ZN(n7160) );
  NOR2_X1 U4955 ( .A1(n8281), .A2(n4405), .ZN(n4404) );
  INV_X1 U4956 ( .A(n7074), .ZN(n4405) );
  INV_X1 U4957 ( .A(n9861), .ZN(n8832) );
  XNOR2_X1 U4958 ( .A(n4743), .B(P2_IR_REG_20__SCAN_IN), .ZN(n8765) );
  INV_X1 U4959 ( .A(n8997), .ZN(n7193) );
  NAND2_X1 U4960 ( .A1(n6848), .A2(n9559), .ZN(n9560) );
  NOR2_X1 U4961 ( .A1(n7835), .A2(n9289), .ZN(n9067) );
  AND2_X1 U4962 ( .A1(n9077), .A2(n9087), .ZN(n7833) );
  AND2_X1 U4963 ( .A1(n7639), .A2(n7840), .ZN(n7455) );
  NOR2_X1 U4964 ( .A1(n7455), .A2(n4498), .ZN(n4497) );
  INV_X1 U4965 ( .A(n4500), .ZN(n4498) );
  NOR2_X1 U4966 ( .A1(n9085), .A2(n7452), .ZN(n4496) );
  OR2_X1 U4967 ( .A1(n9295), .A2(n9108), .ZN(n4500) );
  OR2_X1 U4968 ( .A1(n9303), .A2(n9141), .ZN(n5850) );
  OR2_X1 U4969 ( .A1(n9303), .A2(n8908), .ZN(n9128) );
  AOI21_X1 U4970 ( .B1(n4506), .B2(n4508), .A(n7623), .ZN(n4504) );
  INV_X1 U4971 ( .A(n4506), .ZN(n4505) );
  AOI21_X1 U4972 ( .B1(n4507), .B2(n5818), .A(n4296), .ZN(n4506) );
  INV_X1 U4973 ( .A(n7447), .ZN(n7587) );
  INV_X1 U4974 ( .A(n5613), .ZN(n7425) );
  AND2_X1 U4975 ( .A1(n6448), .A2(n5588), .ZN(n4512) );
  NAND2_X1 U4976 ( .A1(n8139), .A2(n8134), .ZN(n4584) );
  INV_X1 U4977 ( .A(n7675), .ZN(n4353) );
  NAND2_X1 U4978 ( .A1(n6270), .A2(n7675), .ZN(n4352) );
  OAI21_X1 U4979 ( .B1(n4587), .B2(n8128), .A(n4586), .ZN(n4585) );
  AND2_X1 U4980 ( .A1(n8139), .A2(n8129), .ZN(n4587) );
  NAND2_X1 U4981 ( .A1(n7544), .A2(n4322), .ZN(n4321) );
  NOR2_X1 U4982 ( .A1(n4324), .A2(n4323), .ZN(n4322) );
  INV_X1 U4983 ( .A(n7545), .ZN(n4323) );
  OAI21_X1 U4984 ( .B1(n7561), .B2(n4297), .A(n4326), .ZN(n7565) );
  NAND2_X1 U4985 ( .A1(n4604), .A2(n4603), .ZN(n8210) );
  NOR2_X1 U4986 ( .A1(n8198), .A2(n8200), .ZN(n4603) );
  OAI21_X1 U4987 ( .B1(n8188), .B2(n4606), .A(n4605), .ZN(n4604) );
  NAND2_X1 U4988 ( .A1(n7601), .A2(n7547), .ZN(n4337) );
  NAND2_X1 U4989 ( .A1(n7605), .A2(n7650), .ZN(n4336) );
  NAND2_X1 U4990 ( .A1(n7606), .A2(n7650), .ZN(n4339) );
  NAND2_X1 U4991 ( .A1(n7602), .A2(n7547), .ZN(n4340) );
  NOR2_X1 U4992 ( .A1(n8522), .A2(n8231), .ZN(n4597) );
  NAND2_X1 U4993 ( .A1(n4341), .A2(n7614), .ZN(n7617) );
  OAI21_X1 U4994 ( .B1(n7613), .B2(n7612), .A(n7611), .ZN(n4341) );
  CLKBUF_X1 U4995 ( .A(n8262), .Z(n4595) );
  AND2_X1 U4996 ( .A1(n8885), .A2(n4552), .ZN(n4551) );
  NAND2_X1 U4997 ( .A1(n8931), .A2(n4553), .ZN(n4552) );
  INV_X1 U4998 ( .A(n8929), .ZN(n4553) );
  INV_X1 U4999 ( .A(n8931), .ZN(n4554) );
  INV_X1 U5000 ( .A(n7645), .ZN(n4345) );
  NAND2_X1 U5001 ( .A1(n4334), .A2(n7639), .ZN(n7643) );
  OAI21_X1 U5002 ( .B1(n7632), .B2(n4331), .A(n4329), .ZN(n4334) );
  NAND2_X1 U5003 ( .A1(n4332), .A2(n7637), .ZN(n4331) );
  AOI21_X1 U5004 ( .B1(n4332), .B2(n4330), .A(n4262), .ZN(n4329) );
  OR2_X1 U5005 ( .A1(n5712), .A2(n5711), .ZN(n5714) );
  INV_X1 U5006 ( .A(n7579), .ZN(n5894) );
  INV_X1 U5007 ( .A(n4572), .ZN(n4571) );
  INV_X1 U5008 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4755) );
  INV_X1 U5009 ( .A(n4802), .ZN(n4940) );
  NAND2_X1 U5010 ( .A1(n7000), .A2(n4474), .ZN(n7002) );
  NAND2_X1 U5011 ( .A1(n7001), .A2(n8741), .ZN(n4474) );
  NOR2_X1 U5012 ( .A1(n4529), .A2(n8779), .ZN(n4528) );
  INV_X1 U5013 ( .A(n4530), .ZN(n4529) );
  NOR2_X1 U5014 ( .A1(n8786), .A2(n8534), .ZN(n4530) );
  OR2_X1 U5015 ( .A1(n8786), .A2(n7955), .ZN(n8233) );
  NOR2_X1 U5016 ( .A1(n8577), .A2(n4685), .ZN(n4684) );
  INV_X1 U5017 ( .A(n8217), .ZN(n4685) );
  NOR2_X1 U5018 ( .A1(n8693), .A2(n7917), .ZN(n4526) );
  XNOR2_X1 U5019 ( .A(n7917), .B(n8728), .ZN(n8288) );
  AND3_X1 U5020 ( .A1(n8723), .A2(n8705), .A3(n7872), .ZN(n8704) );
  OR2_X1 U5021 ( .A1(n4972), .A2(n6405), .ZN(n4993) );
  OR2_X1 U5022 ( .A1(n7062), .A2(n9844), .ZN(n8161) );
  NOR2_X1 U5023 ( .A1(n7067), .A2(n9844), .ZN(n4518) );
  OR2_X1 U5024 ( .A1(n8765), .A2(n5463), .ZN(n6684) );
  NAND2_X1 U5025 ( .A1(n4400), .A2(n9801), .ZN(n6930) );
  NAND2_X1 U5026 ( .A1(n6930), .A2(n8124), .ZN(n8272) );
  NAND2_X1 U5027 ( .A1(n6699), .A2(n6697), .ZN(n6721) );
  NAND2_X1 U5028 ( .A1(n6691), .A2(n9778), .ZN(n6703) );
  AND2_X1 U5029 ( .A1(n8682), .A2(n8690), .ZN(n8689) );
  NAND2_X1 U5030 ( .A1(n4708), .A2(n4577), .ZN(n4576) );
  INV_X1 U5031 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n4577) );
  OR2_X1 U5032 ( .A1(n6195), .A2(n6609), .ZN(n6605) );
  NAND2_X1 U5033 ( .A1(n8982), .A2(n8980), .ZN(n4566) );
  AND2_X1 U5034 ( .A1(n4312), .A2(n8980), .ZN(n4567) );
  INV_X1 U5035 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5600) );
  AND2_X1 U5036 ( .A1(n7525), .A2(n9128), .ZN(n7465) );
  INV_X1 U5037 ( .A(n4638), .ZN(n4636) );
  NOR2_X1 U5038 ( .A1(n4640), .A2(n4639), .ZN(n4638) );
  INV_X1 U5039 ( .A(n7463), .ZN(n4640) );
  INV_X1 U5040 ( .A(n7629), .ZN(n4639) );
  NOR2_X1 U5041 ( .A1(n9303), .A2(n9309), .ZN(n4463) );
  OR2_X1 U5042 ( .A1(n9309), .A2(n8899), .ZN(n7625) );
  OR2_X1 U5043 ( .A1(n5905), .A2(n4628), .ZN(n4627) );
  INV_X1 U5044 ( .A(n7611), .ZN(n4628) );
  INV_X1 U5045 ( .A(n7616), .ZN(n4624) );
  INV_X1 U5046 ( .A(n9159), .ZN(n5907) );
  OR2_X1 U5047 ( .A1(n9251), .A2(n7343), .ZN(n7598) );
  NOR2_X1 U5048 ( .A1(n9344), .A2(n4449), .ZN(n4448) );
  INV_X1 U5049 ( .A(n4450), .ZN(n4449) );
  NOR2_X1 U5050 ( .A1(n7358), .A2(n7210), .ZN(n4450) );
  OR2_X1 U5051 ( .A1(n7358), .A2(n7267), .ZN(n7591) );
  OR2_X1 U5052 ( .A1(n7240), .A2(n7256), .ZN(n7219) );
  INV_X1 U5053 ( .A(n7552), .ZN(n4617) );
  INV_X1 U5054 ( .A(n4616), .ZN(n4615) );
  OAI21_X1 U5055 ( .B1(n7439), .B2(n4617), .A(n7551), .ZN(n4616) );
  NAND2_X1 U5056 ( .A1(n5620), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n4622) );
  OR2_X1 U5057 ( .A1(n5537), .A2(n5526), .ZN(n4618) );
  NAND2_X1 U5058 ( .A1(n5339), .A2(n5338), .ZN(n5354) );
  NAND2_X1 U5059 ( .A1(n5335), .A2(n5334), .ZN(n5339) );
  AND2_X1 U5060 ( .A1(n5267), .A2(n5265), .ZN(n5266) );
  AND2_X1 U5061 ( .A1(n5230), .A2(n5231), .ZN(n5253) );
  AND2_X1 U5062 ( .A1(n5199), .A2(n5200), .ZN(n5230) );
  OR2_X1 U5063 ( .A1(n5205), .A2(n5204), .ZN(n5233) );
  AND2_X1 U5064 ( .A1(n5107), .A2(n5072), .ZN(n5105) );
  INV_X1 U5065 ( .A(n5078), .ZN(n5065) );
  NAND2_X1 U5066 ( .A1(n4669), .A2(n4671), .ZN(n5056) );
  INV_X1 U5067 ( .A(n4672), .ZN(n4671) );
  OAI21_X1 U5068 ( .B1(n4674), .B2(n4673), .A(n5042), .ZN(n4672) );
  INV_X1 U5069 ( .A(n4647), .ZN(n4644) );
  NAND2_X1 U5070 ( .A1(n4250), .A2(n4923), .ZN(n4650) );
  AND2_X1 U5071 ( .A1(n4871), .A2(n4892), .ZN(n4651) );
  INV_X1 U5072 ( .A(n4875), .ZN(n4654) );
  NOR2_X1 U5073 ( .A1(n5399), .A2(n4363), .ZN(n4362) );
  INV_X1 U5074 ( .A(n5377), .ZN(n4363) );
  INV_X1 U5075 ( .A(n5459), .ZN(n4357) );
  NAND2_X1 U5076 ( .A1(n4361), .A2(n4365), .ZN(n4360) );
  INV_X1 U5077 ( .A(n7952), .ZN(n4361) );
  NAND2_X1 U5078 ( .A1(n8083), .A2(n4879), .ZN(n8082) );
  INV_X1 U5079 ( .A(n7990), .ZN(n4378) );
  AND2_X1 U5080 ( .A1(n7717), .A2(n7716), .ZN(n8002) );
  OAI21_X1 U5081 ( .B1(n4666), .B2(n8256), .A(n8249), .ZN(n4665) );
  AND3_X1 U5082 ( .A1(n5351), .A2(n5350), .A3(n5349), .ZN(n8095) );
  NAND2_X1 U5083 ( .A1(n4259), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n4403) );
  NAND2_X1 U5084 ( .A1(n4816), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n4402) );
  AOI21_X1 U5085 ( .B1(n6337), .B2(P2_REG2_REG_1__SCAN_IN), .A(n6336), .ZN(
        n9379) );
  AOI21_X1 U5086 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n6551), .A(n8382), .ZN(
        n6553) );
  NAND2_X1 U5087 ( .A1(n6666), .A2(n6667), .ZN(n7000) );
  NAND2_X1 U5088 ( .A1(n4486), .A2(n4485), .ZN(n4484) );
  INV_X1 U5089 ( .A(n8416), .ZN(n4485) );
  NAND2_X1 U5090 ( .A1(n4664), .A2(n4666), .ZN(n8105) );
  NAND2_X1 U5091 ( .A1(n8490), .A2(n8730), .ZN(n7907) );
  OR2_X1 U5092 ( .A1(n8779), .A2(n8473), .ZN(n7943) );
  OR2_X1 U5093 ( .A1(n8786), .A2(n8489), .ZN(n7942) );
  AND2_X1 U5094 ( .A1(n8560), .A2(n8796), .ZN(n8548) );
  AND2_X1 U5095 ( .A1(n4681), .A2(n8223), .ZN(n4679) );
  INV_X1 U5096 ( .A(n8570), .ZN(n4394) );
  NOR2_X1 U5097 ( .A1(n4594), .A2(n4395), .ZN(n4392) );
  NAND2_X1 U5098 ( .A1(n4688), .A2(n4687), .ZN(n4686) );
  INV_X1 U5099 ( .A(n8605), .ZN(n8616) );
  NAND2_X1 U5100 ( .A1(n7932), .A2(n4397), .ZN(n4396) );
  NAND2_X1 U5101 ( .A1(n8639), .A2(n8211), .ZN(n4659) );
  NAND2_X1 U5102 ( .A1(n8831), .A2(n8316), .ZN(n4399) );
  NOR2_X1 U5103 ( .A1(n8181), .A2(n4412), .ZN(n4411) );
  NAND2_X1 U5104 ( .A1(n5045), .A2(n4660), .ZN(n8705) );
  AND2_X1 U5105 ( .A1(n4663), .A2(n5044), .ZN(n4660) );
  INV_X1 U5106 ( .A(n7178), .ZN(n8284) );
  NAND2_X1 U5107 ( .A1(n7160), .A2(n7159), .ZN(n7161) );
  INV_X1 U5108 ( .A(n7299), .ZN(n8285) );
  NAND2_X1 U5109 ( .A1(n6952), .A2(n6951), .ZN(n7075) );
  INV_X1 U5110 ( .A(n8110), .ZN(n5184) );
  INV_X1 U5111 ( .A(n5997), .ZN(n5183) );
  NAND2_X1 U5112 ( .A1(n9816), .A2(n4406), .ZN(n7086) );
  NOR2_X1 U5113 ( .A1(n4269), .A2(n4407), .ZN(n4406) );
  INV_X1 U5114 ( .A(n6948), .ZN(n4407) );
  OAI21_X1 U5115 ( .B1(n5156), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n4744) );
  OR2_X1 U5116 ( .A1(n6775), .A2(n6774), .ZN(n6776) );
  INV_X1 U5117 ( .A(n8650), .ZN(n8729) );
  OR2_X1 U5118 ( .A1(n9861), .A2(n4764), .ZN(n8754) );
  OR2_X1 U5119 ( .A1(n8270), .A2(n6708), .ZN(n9748) );
  INV_X1 U5120 ( .A(n8550), .ZN(n8796) );
  INV_X1 U5121 ( .A(n8675), .ZN(n9429) );
  AND3_X1 U5122 ( .A1(n4855), .A2(n4854), .A3(n4853), .ZN(n9810) );
  INV_X1 U5123 ( .A(n9843), .ZN(n9859) );
  AND2_X1 U5124 ( .A1(n5418), .A2(n4720), .ZN(n4721) );
  NOR2_X1 U5125 ( .A1(n5156), .A2(n4578), .ZN(n4738) );
  NAND2_X1 U5126 ( .A1(n4298), .A2(n4579), .ZN(n4578) );
  INV_X1 U5127 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n4579) );
  NAND2_X1 U5128 ( .A1(n4476), .A2(n4737), .ZN(n4475) );
  OAI21_X1 U5129 ( .B1(n8982), .B2(n4312), .A(n8980), .ZN(n4563) );
  NAND2_X1 U5130 ( .A1(n4568), .A2(n4567), .ZN(n4558) );
  NAND2_X1 U5131 ( .A1(n4540), .A2(n7789), .ZN(n8869) );
  INV_X1 U5132 ( .A(n4543), .ZN(n4540) );
  NAND2_X1 U5133 ( .A1(n4543), .A2(n7788), .ZN(n8870) );
  NOR2_X1 U5134 ( .A1(n4565), .A2(n4557), .ZN(n4556) );
  INV_X1 U5135 ( .A(n8895), .ZN(n4557) );
  INV_X1 U5136 ( .A(n4567), .ZN(n4561) );
  NOR2_X1 U5137 ( .A1(n5606), .A2(n5605), .ZN(n5621) );
  NAND2_X1 U5138 ( .A1(n4547), .A2(n4546), .ZN(n4548) );
  NOR2_X1 U5139 ( .A1(n6298), .A2(n6150), .ZN(n4546) );
  OR2_X1 U5140 ( .A1(n5703), .A2(n5702), .ZN(n5705) );
  AND4_X1 U5141 ( .A1(n5654), .A2(n5653), .A3(n5652), .A4(n5651), .ZN(n6879)
         );
  OR2_X1 U5142 ( .A1(n6062), .A2(n6061), .ZN(n4470) );
  NOR2_X1 U5143 ( .A1(n9534), .A2(n4418), .ZN(n9548) );
  AND2_X1 U5144 ( .A1(n9539), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n4418) );
  OR2_X1 U5145 ( .A1(n9548), .A2(n9547), .ZN(n4417) );
  OR2_X1 U5146 ( .A1(n9554), .A2(n9553), .ZN(n4442) );
  OR2_X1 U5147 ( .A1(n9586), .A2(n9585), .ZN(n4454) );
  INV_X1 U5148 ( .A(n4436), .ZN(n4435) );
  OAI21_X1 U5149 ( .B1(n9576), .B2(n6853), .A(n6854), .ZN(n4436) );
  NAND2_X1 U5150 ( .A1(n9577), .A2(n9576), .ZN(n4432) );
  AND2_X1 U5151 ( .A1(n6856), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n9038) );
  OR2_X1 U5152 ( .A1(n9602), .A2(n4319), .ZN(n4429) );
  NAND2_X1 U5153 ( .A1(n4429), .A2(n4428), .ZN(n4427) );
  INV_X1 U5154 ( .A(n9616), .ZN(n4428) );
  NAND2_X1 U5155 ( .A1(n5910), .A2(n7637), .ZN(n5912) );
  NAND2_X1 U5156 ( .A1(n5906), .A2(n5905), .ZN(n9187) );
  NAND2_X1 U5157 ( .A1(n9251), .A2(n7343), .ZN(n9229) );
  NOR2_X1 U5158 ( .A1(n9334), .A2(n9246), .ZN(n9223) );
  NAND2_X1 U5159 ( .A1(n5753), .A2(n4264), .ZN(n4511) );
  NAND2_X1 U5160 ( .A1(n4511), .A2(n4510), .ZN(n9258) );
  AND2_X1 U5161 ( .A1(n5765), .A2(n5754), .ZN(n4510) );
  AND2_X1 U5162 ( .A1(n7598), .A2(n9229), .ZN(n9255) );
  AND2_X1 U5163 ( .A1(n5898), .A2(n9238), .ZN(n9270) );
  NAND2_X1 U5164 ( .A1(n5897), .A2(n7587), .ZN(n7349) );
  NOR2_X1 U5165 ( .A1(n5705), .A2(n5688), .ZN(n5724) );
  NOR2_X1 U5166 ( .A1(n7219), .A2(n7473), .ZN(n9471) );
  NOR2_X1 U5167 ( .A1(n5663), .A2(n5662), .ZN(n5677) );
  NOR2_X1 U5168 ( .A1(n7439), .A2(n4503), .ZN(n4502) );
  INV_X1 U5169 ( .A(n5612), .ZN(n4503) );
  NAND2_X1 U5170 ( .A1(n5890), .A2(n7679), .ZN(n4632) );
  AND4_X1 U5171 ( .A1(n5598), .A2(n5597), .A3(n5596), .A4(n5595), .ZN(n6615)
         );
  AND4_X1 U5172 ( .A1(n5586), .A2(n5585), .A3(n5584), .A4(n5583), .ZN(n8922)
         );
  OR2_X1 U5173 ( .A1(n5549), .A2(n5581), .ZN(n5584) );
  INV_X1 U5174 ( .A(n7426), .ZN(n5773) );
  NAND2_X1 U5175 ( .A1(n5587), .A2(n6310), .ZN(n6312) );
  INV_X1 U5176 ( .A(n9005), .ZN(n6486) );
  INV_X1 U5177 ( .A(n9210), .ZN(n9656) );
  XNOR2_X1 U5178 ( .A(n7669), .B(n5547), .ZN(n6252) );
  OR2_X1 U5179 ( .A1(n7654), .A2(n6199), .ZN(n9210) );
  NAND2_X1 U5180 ( .A1(n7428), .A2(n7427), .ZN(n9289) );
  NAND2_X1 U5181 ( .A1(n5861), .A2(n5860), .ZN(n9295) );
  NAND2_X1 U5182 ( .A1(n5820), .A2(n5819), .ZN(n9313) );
  AND2_X1 U5183 ( .A1(n6457), .A2(n9389), .ZN(n9349) );
  INV_X1 U5184 ( .A(n6488), .ZN(n9694) );
  OR2_X1 U5185 ( .A1(n7650), .A2(n7701), .ZN(n9389) );
  XNOR2_X1 U5186 ( .A(n7379), .B(n7378), .ZN(n7317) );
  XNOR2_X1 U5187 ( .A(n5413), .B(n5412), .ZN(n7156) );
  AOI21_X1 U5188 ( .B1(n5937), .B2(n5936), .A(n5878), .ZN(n4533) );
  XNOR2_X1 U5189 ( .A(n5380), .B(n5379), .ZN(n7081) );
  XNOR2_X1 U5190 ( .A(n5182), .B(n5201), .ZN(n6538) );
  XNOR2_X1 U5191 ( .A(n5056), .B(n5057), .ZN(n6135) );
  NAND2_X1 U5192 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(n4272), .ZN(n4423) );
  AND4_X1 U5193 ( .A1(n5023), .A2(n5022), .A3(n5021), .A4(n5020), .ZN(n7365)
         );
  NAND2_X1 U5194 ( .A1(n5045), .A2(n5044), .ZN(n7871) );
  OAI21_X1 U5195 ( .B1(n5976), .B2(n5971), .A(n5975), .ZN(n7042) );
  NAND2_X1 U5196 ( .A1(n4811), .A2(n4367), .ZN(n4366) );
  NAND2_X1 U5197 ( .A1(n4813), .A2(n6569), .ZN(n4368) );
  INV_X1 U5198 ( .A(n4812), .ZN(n4367) );
  AND4_X1 U5199 ( .A1(n4945), .A2(n4944), .A3(n4943), .A4(n4942), .ZN(n7073)
         );
  NAND2_X1 U5200 ( .A1(n4370), .A2(n4369), .ZN(n6578) );
  INV_X1 U5201 ( .A(n6576), .ZN(n4369) );
  INV_X1 U5202 ( .A(n6575), .ZN(n4370) );
  INV_X1 U5203 ( .A(n6968), .ZN(n9837) );
  AND2_X1 U5204 ( .A1(n5467), .A2(n5464), .ZN(n8085) );
  NAND2_X1 U5205 ( .A1(n5454), .A2(n8739), .ZN(n8101) );
  AND2_X1 U5206 ( .A1(n5996), .A2(n5469), .ZN(n8730) );
  AND2_X1 U5207 ( .A1(n6340), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4482) );
  NAND2_X1 U5208 ( .A1(n4481), .A2(n4277), .ZN(n6360) );
  OR2_X1 U5209 ( .A1(n8414), .A2(n4487), .ZN(n4486) );
  NOR2_X1 U5210 ( .A1(n8420), .A2(n4488), .ZN(n4487) );
  INV_X1 U5211 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n4488) );
  INV_X1 U5212 ( .A(n4484), .ZN(n8433) );
  NOR2_X1 U5213 ( .A1(n8458), .A2(n8465), .ZN(n8460) );
  AND2_X1 U5214 ( .A1(n7892), .A2(n7891), .ZN(n7915) );
  OR2_X1 U5215 ( .A1(n8633), .A2(n8632), .ZN(n8828) );
  AND3_X1 U5216 ( .A1(n4900), .A2(n4899), .A3(n4898), .ZN(n9823) );
  INV_X1 U5217 ( .A(n9750), .ZN(n8739) );
  INV_X1 U5218 ( .A(n5531), .ZN(n5969) );
  OAI211_X1 U5219 ( .C1(n7657), .C2(n9146), .A(n7661), .B(n4351), .ZN(n4350)
         );
  AOI21_X1 U5220 ( .B1(n4261), .B2(n9146), .A(n6565), .ZN(n4351) );
  OAI211_X1 U5221 ( .C1(n7702), .C2(n7701), .A(n7700), .B(n7699), .ZN(n7703)
         );
  OR2_X1 U5222 ( .A1(n7698), .A2(n7697), .ZN(n7699) );
  INV_X1 U5223 ( .A(n9123), .ZN(n9088) );
  INV_X1 U5224 ( .A(n6615), .ZN(n9003) );
  NOR2_X1 U5225 ( .A1(n6091), .A2(n4414), .ZN(n9028) );
  NOR2_X1 U5226 ( .A1(n6072), .A2(n4415), .ZN(n4414) );
  INV_X1 U5227 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n4415) );
  NAND2_X1 U5228 ( .A1(n9028), .A2(n9027), .ZN(n9026) );
  NAND2_X1 U5229 ( .A1(n9508), .A2(n9509), .ZN(n9507) );
  AND2_X1 U5230 ( .A1(n6105), .A2(n4471), .ZN(n6062) );
  NAND2_X1 U5231 ( .A1(n6059), .A2(n6060), .ZN(n4471) );
  AOI21_X1 U5232 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n9635), .A(n9629), .ZN(
        n9045) );
  AOI21_X1 U5233 ( .B1(n4610), .B2(n9651), .A(n4609), .ZN(n9290) );
  OAI22_X1 U5234 ( .A1(n8862), .A2(n9212), .B1(n7459), .B2(n7845), .ZN(n4609)
         );
  XNOR2_X1 U5235 ( .A(n4611), .B(n7642), .ZN(n4610) );
  INV_X1 U5236 ( .A(n4492), .ZN(n7834) );
  OAI21_X1 U5237 ( .B1(n9098), .B2(n4289), .A(n4493), .ZN(n4492) );
  AOI21_X1 U5238 ( .B1(n4494), .B2(n4497), .A(n7833), .ZN(n4493) );
  AOI21_X1 U5239 ( .B1(n9112), .B2(n9651), .A(n9111), .ZN(n9301) );
  NAND2_X1 U5240 ( .A1(n9110), .A2(n9109), .ZN(n9111) );
  AND2_X1 U5241 ( .A1(n9678), .A2(n6285), .ZN(n9484) );
  NOR2_X1 U5242 ( .A1(n9081), .A2(n5926), .ZN(n5927) );
  NAND2_X1 U5243 ( .A1(n9073), .A2(n9718), .ZN(n5928) );
  AND2_X1 U5244 ( .A1(n4629), .A2(n5496), .ZN(n4467) );
  NAND2_X1 U5245 ( .A1(n4582), .A2(n4581), .ZN(n4580) );
  NOR2_X1 U5246 ( .A1(n6954), .A2(n4590), .ZN(n4581) );
  NAND2_X1 U5247 ( .A1(n4584), .A2(n4583), .ZN(n4582) );
  NAND2_X1 U5248 ( .A1(n8133), .A2(n8132), .ZN(n4583) );
  NAND2_X1 U5249 ( .A1(n4589), .A2(n4588), .ZN(n8139) );
  NAND2_X1 U5250 ( .A1(n8131), .A2(n4590), .ZN(n4589) );
  NOR2_X1 U5251 ( .A1(n8670), .A2(n8193), .ZN(n4605) );
  INV_X1 U5252 ( .A(n8210), .ZN(n8207) );
  NAND2_X1 U5253 ( .A1(n4594), .A2(n4287), .ZN(n4593) );
  NAND2_X1 U5254 ( .A1(n4340), .A2(n4339), .ZN(n4338) );
  NAND2_X1 U5255 ( .A1(n4337), .A2(n4336), .ZN(n4335) );
  AND2_X1 U5256 ( .A1(n7497), .A2(n7555), .ZN(n7564) );
  AOI21_X1 U5257 ( .B1(n4600), .B2(n4599), .A(n4596), .ZN(n8240) );
  INV_X1 U5258 ( .A(n8225), .ZN(n4599) );
  NAND2_X1 U5259 ( .A1(n4598), .A2(n4597), .ZN(n4596) );
  NOR2_X1 U5260 ( .A1(n4279), .A2(n7685), .ZN(n4330) );
  INV_X1 U5261 ( .A(n7633), .ZN(n4333) );
  OR2_X1 U5262 ( .A1(n5535), .A2(n9009), .ZN(n5519) );
  OR2_X1 U5263 ( .A1(n9331), .A2(n8888), .ZN(n7604) );
  AND2_X1 U5264 ( .A1(n5040), .A2(n4677), .ZN(n4670) );
  INV_X1 U5265 ( .A(n4701), .ZN(n4648) );
  INV_X1 U5266 ( .A(n4946), .ZN(n4649) );
  XNOR2_X1 U5267 ( .A(n9793), .B(n5410), .ZN(n4784) );
  AOI21_X1 U5268 ( .B1(n8250), .B2(n8255), .A(n4595), .ZN(n4574) );
  NOR2_X1 U5269 ( .A1(n8254), .A2(n4284), .ZN(n4575) );
  AND2_X1 U5270 ( .A1(n8252), .A2(n8241), .ZN(n4668) );
  NOR2_X1 U5271 ( .A1(n8812), .A2(n8613), .ZN(n4520) );
  INV_X1 U5272 ( .A(n7931), .ZN(n4397) );
  NAND2_X1 U5273 ( .A1(n4526), .A2(n9429), .ZN(n4525) );
  INV_X1 U5274 ( .A(n7311), .ZN(n4412) );
  OR2_X1 U5275 ( .A1(n8693), .A2(n7882), .ZN(n8190) );
  AND2_X1 U5276 ( .A1(n6930), .A2(n8129), .ZN(n8125) );
  INV_X1 U5277 ( .A(n6771), .ZN(n6775) );
  AND2_X1 U5278 ( .A1(n4267), .A2(n9819), .ZN(n4521) );
  INV_X1 U5279 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5420) );
  AND4_X1 U5280 ( .A1(n4373), .A2(n4712), .A3(n4374), .A4(n4750), .ZN(n4372)
         );
  AOI21_X1 U5281 ( .B1(n4551), .B2(n4554), .A(n4292), .ZN(n4550) );
  OAI211_X1 U5282 ( .C1(n7644), .C2(n7547), .A(n4346), .B(n4344), .ZN(n4343)
         );
  NOR2_X1 U5283 ( .A1(n4700), .A2(n4347), .ZN(n4346) );
  NAND2_X1 U5284 ( .A1(n4345), .A2(n7547), .ZN(n4344) );
  AND2_X1 U5285 ( .A1(n7457), .A2(n7712), .ZN(n7517) );
  NOR2_X1 U5286 ( .A1(n9299), .A2(n4462), .ZN(n4461) );
  INV_X1 U5287 ( .A(n4463), .ZN(n4462) );
  OR2_X1 U5288 ( .A1(n9313), .A2(n8943), .ZN(n7462) );
  NOR2_X1 U5289 ( .A1(n9181), .A2(n9195), .ZN(n9167) );
  OR2_X1 U5290 ( .A1(n9195), .A2(n9209), .ZN(n7608) );
  AND2_X1 U5291 ( .A1(n7598), .A2(n9238), .ZN(n7593) );
  NAND2_X1 U5292 ( .A1(n7349), .A2(n7471), .ZN(n9239) );
  NAND2_X1 U5293 ( .A1(n5891), .A2(n7558), .ZN(n4633) );
  OR2_X1 U5294 ( .A1(n9390), .A2(n6879), .ZN(n7555) );
  NAND2_X1 U5295 ( .A1(n6520), .A2(n7439), .ZN(n9647) );
  NOR2_X1 U5296 ( .A1(n6458), .A2(n8973), .ZN(n6459) );
  OR2_X1 U5297 ( .A1(n6432), .A2(n6275), .ZN(n7486) );
  AND2_X1 U5298 ( .A1(n7584), .A2(n7585), .ZN(n9476) );
  INV_X1 U5299 ( .A(n7445), .ZN(n5895) );
  AND2_X1 U5300 ( .A1(n6305), .A2(n9688), .ZN(n4469) );
  AND3_X1 U5301 ( .A1(n4468), .A2(n6496), .A3(n6305), .ZN(n6437) );
  INV_X1 U5302 ( .A(n6289), .ZN(n6305) );
  NOR2_X1 U5303 ( .A1(n4570), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n4569) );
  NAND2_X1 U5304 ( .A1(n4571), .A2(n4295), .ZN(n4570) );
  NAND2_X1 U5305 ( .A1(n5255), .A2(n5254), .ZN(n5268) );
  AND2_X1 U5306 ( .A1(n5253), .A2(n5256), .ZN(n5254) );
  NAND2_X1 U5307 ( .A1(n4573), .A2(n5771), .ZN(n4572) );
  INV_X1 U5308 ( .A(n5769), .ZN(n4573) );
  AND2_X1 U5309 ( .A1(n5231), .A2(n5210), .ZN(n5232) );
  AND2_X1 U5310 ( .A1(n5171), .A2(n5170), .ZN(n5199) );
  AND2_X1 U5311 ( .A1(n5176), .A2(n5175), .ZN(n5203) );
  OR2_X1 U5312 ( .A1(n5173), .A2(n5172), .ZN(n5176) );
  NOR2_X1 U5313 ( .A1(n5028), .A2(n4678), .ZN(n4677) );
  INV_X1 U5314 ( .A(n5001), .ZN(n4678) );
  AOI21_X1 U5315 ( .B1(n4677), .B2(n5002), .A(n4675), .ZN(n4674) );
  INV_X1 U5316 ( .A(n5008), .ZN(n4675) );
  INV_X1 U5317 ( .A(n4999), .ZN(n5002) );
  XNOR2_X1 U5318 ( .A(n5000), .B(n10044), .ZN(n4999) );
  OAI21_X1 U5319 ( .B1(n7393), .B2(P1_DATAO_REG_4__SCAN_IN), .A(n4829), .ZN(
        n4848) );
  NAND2_X1 U5320 ( .A1(n7393), .A2(n6019), .ZN(n4829) );
  NAND2_X1 U5321 ( .A1(n5529), .A2(n4491), .ZN(n4758) );
  NAND2_X1 U5322 ( .A1(n8082), .A2(n4380), .ZN(n6828) );
  AND2_X1 U5323 ( .A1(n4905), .A2(n4883), .ZN(n4380) );
  AND2_X1 U5324 ( .A1(n5228), .A2(n5198), .ZN(n4381) );
  OR2_X1 U5325 ( .A1(n5241), .A2(n10045), .ZN(n5279) );
  NOR2_X1 U5326 ( .A1(n5475), .A2(n9764), .ZN(n5467) );
  OR3_X1 U5327 ( .A1(n5049), .A2(n5048), .A3(n5047), .ZN(n5089) );
  AND2_X1 U5328 ( .A1(n5369), .A2(n5368), .ZN(n7955) );
  AND3_X1 U5329 ( .A1(n5314), .A2(n5313), .A3(n5312), .ZN(n8031) );
  AND4_X1 U5330 ( .A1(n5223), .A2(n5222), .A3(n5221), .A4(n5220), .ZN(n7984)
         );
  NAND2_X1 U5331 ( .A1(n6401), .A2(n6366), .ZN(n8354) );
  AND2_X1 U5332 ( .A1(n6548), .A2(n4490), .ZN(n8367) );
  NAND2_X1 U5333 ( .A1(n6549), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n4490) );
  NAND2_X1 U5334 ( .A1(n8367), .A2(n8366), .ZN(n8365) );
  NAND2_X1 U5335 ( .A1(n8365), .A2(n4489), .ZN(n8384) );
  OR2_X1 U5336 ( .A1(n8370), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n4489) );
  INV_X1 U5337 ( .A(n7002), .ZN(n8405) );
  XNOR2_X1 U5338 ( .A(n8443), .B(n8439), .ZN(n8435) );
  AND2_X1 U5339 ( .A1(n4484), .A2(n4483), .ZN(n8443) );
  NAND2_X1 U5340 ( .A1(n8434), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4483) );
  INV_X1 U5341 ( .A(n8487), .ZN(n8501) );
  NAND2_X1 U5342 ( .A1(n8502), .A2(n8501), .ZN(n8500) );
  NAND2_X1 U5343 ( .A1(n8548), .A2(n4528), .ZN(n8493) );
  AND2_X1 U5344 ( .A1(n8241), .A2(n8244), .ZN(n8487) );
  AOI21_X1 U5345 ( .B1(n8526), .B2(n7888), .A(n8232), .ZN(n8488) );
  OR2_X1 U5346 ( .A1(n8534), .A2(n8544), .ZN(n7941) );
  NAND2_X1 U5347 ( .A1(n8548), .A2(n4530), .ZN(n8509) );
  OR2_X1 U5348 ( .A1(n8534), .A2(n8095), .ZN(n8505) );
  NAND2_X1 U5349 ( .A1(n8548), .A2(n8791), .ZN(n8531) );
  AND2_X1 U5350 ( .A1(n8505), .A2(n8235), .ZN(n8528) );
  INV_X1 U5351 ( .A(n8528), .ZN(n8522) );
  OAI21_X1 U5352 ( .B1(n4394), .B2(n4391), .A(n4389), .ZN(n8540) );
  INV_X1 U5353 ( .A(n4392), .ZN(n4391) );
  AOI21_X1 U5354 ( .B1(n4392), .B2(n4390), .A(n4293), .ZN(n4389) );
  AND2_X1 U5355 ( .A1(n8631), .A2(n4519), .ZN(n8560) );
  AND2_X1 U5356 ( .A1(n4268), .A2(n8563), .ZN(n4519) );
  NAND2_X1 U5357 ( .A1(n4689), .A2(n4687), .ZN(n4683) );
  NAND2_X1 U5358 ( .A1(n4682), .A2(n4689), .ZN(n4681) );
  INV_X1 U5359 ( .A(n4684), .ZN(n4682) );
  NAND2_X1 U5360 ( .A1(n8631), .A2(n4268), .ZN(n8572) );
  NAND2_X1 U5361 ( .A1(n8631), .A2(n4520), .ZN(n8589) );
  AND2_X1 U5362 ( .A1(n8214), .A2(n8212), .ZN(n8605) );
  NAND2_X1 U5363 ( .A1(n5114), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5187) );
  NAND2_X1 U5364 ( .A1(n8645), .A2(n8639), .ZN(n8653) );
  AND2_X1 U5365 ( .A1(n8623), .A2(n8209), .ZN(n8639) );
  NAND2_X1 U5366 ( .A1(n8195), .A2(n8194), .ZN(n8670) );
  OR2_X1 U5367 ( .A1(n7927), .A2(n8689), .ZN(n8665) );
  NOR2_X1 U5368 ( .A1(n8738), .A2(n4524), .ZN(n8687) );
  INV_X1 U5369 ( .A(n4526), .ZN(n4524) );
  NOR2_X1 U5370 ( .A1(n8738), .A2(n7917), .ZN(n8712) );
  NOR2_X1 U5371 ( .A1(n8706), .A2(n7876), .ZN(n8702) );
  OR2_X1 U5372 ( .A1(n7873), .A2(n8704), .ZN(n7874) );
  OR2_X1 U5373 ( .A1(n7870), .A2(n7869), .ZN(n7875) );
  INV_X1 U5374 ( .A(n8288), .ZN(n8706) );
  NAND2_X1 U5375 ( .A1(n7910), .A2(n9452), .ZN(n8736) );
  OR2_X1 U5376 ( .A1(n8736), .A2(n7871), .ZN(n8738) );
  NAND2_X1 U5377 ( .A1(n7312), .A2(n7311), .ZN(n7922) );
  OR2_X1 U5378 ( .A1(n7304), .A2(n8286), .ZN(n8724) );
  NOR2_X1 U5379 ( .A1(n7180), .A2(n7170), .ZN(n7910) );
  AND2_X1 U5380 ( .A1(n7178), .A2(n8170), .ZN(n7300) );
  AND2_X1 U5381 ( .A1(n8169), .A2(n8170), .ZN(n7299) );
  NAND2_X1 U5382 ( .A1(n4518), .A2(n4517), .ZN(n7180) );
  INV_X1 U5383 ( .A(n4518), .ZN(n7163) );
  AND2_X1 U5384 ( .A1(n8154), .A2(n8162), .ZN(n8282) );
  AND4_X1 U5385 ( .A1(n4914), .A2(n4913), .A3(n4912), .A4(n4911), .ZN(n6958)
         );
  AND2_X1 U5386 ( .A1(n8152), .A2(n8151), .ZN(n8276) );
  NOR2_X1 U5387 ( .A1(n7093), .A2(n8146), .ZN(n7094) );
  AND2_X1 U5388 ( .A1(n7094), .A2(n9830), .ZN(n7021) );
  NAND2_X1 U5389 ( .A1(n4522), .A2(n4267), .ZN(n6965) );
  INV_X1 U5390 ( .A(n6769), .ZN(n8279) );
  NOR2_X1 U5391 ( .A1(n7131), .A2(n8042), .ZN(n7132) );
  INV_X1 U5392 ( .A(n4515), .ZN(n4514) );
  AND2_X1 U5393 ( .A1(n9763), .A2(n9767), .ZN(n5444) );
  XNOR2_X1 U5394 ( .A(n4388), .B(n7894), .ZN(n8771) );
  NAND2_X1 U5395 ( .A1(n8482), .A2(n4706), .ZN(n4388) );
  INV_X1 U5396 ( .A(n8760), .ZN(n8837) );
  OR2_X1 U5397 ( .A1(n8759), .A2(n8758), .ZN(n8838) );
  NAND2_X1 U5398 ( .A1(n4736), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5430) );
  NOR2_X1 U5399 ( .A1(n4384), .A2(n4576), .ZN(n4383) );
  AND2_X1 U5400 ( .A1(n4869), .A2(n4711), .ZN(n5030) );
  OR2_X1 U5401 ( .A1(n4917), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n4965) );
  NAND2_X1 U5402 ( .A1(n5594), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5606) );
  AND2_X1 U5403 ( .A1(n7141), .A2(n7146), .ZN(n4534) );
  NAND2_X1 U5404 ( .A1(n4532), .A2(n8879), .ZN(n8878) );
  INV_X1 U5405 ( .A(n6150), .ZN(n4545) );
  AND3_X1 U5406 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U5407 ( .A1(n7340), .A2(n7341), .ZN(n7744) );
  AND2_X1 U5408 ( .A1(n7788), .A2(n4542), .ZN(n4541) );
  INV_X1 U5409 ( .A(n8868), .ZN(n4542) );
  NAND2_X1 U5410 ( .A1(n8928), .A2(n8929), .ZN(n8927) );
  OR2_X1 U5411 ( .A1(n5749), .A2(n5748), .ZN(n5761) );
  INV_X1 U5412 ( .A(n5841), .ZN(n5854) );
  NAND2_X1 U5413 ( .A1(n7192), .A2(n7191), .ZN(n7201) );
  INV_X1 U5414 ( .A(n7814), .ZN(n7820) );
  AND4_X1 U5415 ( .A1(n5709), .A2(n5708), .A3(n5707), .A4(n5706), .ZN(n6903)
         );
  OAI21_X1 U5416 ( .B1(n9010), .B2(n9723), .A(n4446), .ZN(n4445) );
  NAND2_X1 U5417 ( .A1(n9010), .A2(n9723), .ZN(n4446) );
  AND2_X1 U5418 ( .A1(n6144), .A2(n6145), .ZN(n6142) );
  AOI21_X1 U5419 ( .B1(P1_REG2_REG_2__SCAN_IN), .B2(n6071), .A(n6142), .ZN(
        n6093) );
  OAI21_X1 U5420 ( .B1(n6075), .B2(P1_REG2_REG_5__SCAN_IN), .A(n9507), .ZN(
        n6109) );
  AND2_X1 U5421 ( .A1(n9514), .A2(n6058), .ZN(n6106) );
  NOR2_X1 U5422 ( .A1(n6108), .A2(n4431), .ZN(n6076) );
  AND2_X1 U5423 ( .A1(n6114), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n4431) );
  NAND2_X1 U5424 ( .A1(n6076), .A2(n6077), .ZN(n6232) );
  NAND2_X1 U5425 ( .A1(n6232), .A2(n4430), .ZN(n9521) );
  OR2_X1 U5426 ( .A1(n6233), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4430) );
  NAND2_X1 U5427 ( .A1(n9521), .A2(n9520), .ZN(n9519) );
  OAI21_X1 U5428 ( .B1(n6234), .B2(P1_REG2_REG_8__SCAN_IN), .A(n9519), .ZN(
        n9536) );
  INV_X1 U5429 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4539) );
  OR2_X1 U5430 ( .A1(n6229), .A2(n6228), .ZN(n4440) );
  AND2_X1 U5431 ( .A1(n4417), .A2(n4416), .ZN(n6238) );
  NAND2_X1 U5432 ( .A1(n9551), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4416) );
  NAND2_X1 U5433 ( .A1(n6238), .A2(n6237), .ZN(n6846) );
  OAI21_X1 U5434 ( .B1(n6847), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6846), .ZN(
        n9562) );
  AND2_X1 U5435 ( .A1(n4440), .A2(n4439), .ZN(n9568) );
  NAND2_X1 U5436 ( .A1(n6839), .A2(n5661), .ZN(n4439) );
  OR2_X1 U5437 ( .A1(n6843), .A2(n6844), .ZN(n4452) );
  NOR2_X1 U5438 ( .A1(n9040), .A2(n9591), .ZN(n9604) );
  AND2_X1 U5439 ( .A1(n4452), .A2(n4451), .ZN(n9048) );
  NAND2_X1 U5440 ( .A1(n4434), .A2(n6835), .ZN(n4451) );
  AND2_X1 U5441 ( .A1(n4427), .A2(n4426), .ZN(n9631) );
  NAND2_X1 U5442 ( .A1(n9620), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n4426) );
  NOR2_X1 U5443 ( .A1(n9631), .A2(n9630), .ZN(n9629) );
  OAI21_X1 U5444 ( .B1(n7842), .B2(n7841), .A(n7840), .ZN(n4611) );
  INV_X1 U5445 ( .A(n4496), .ZN(n4494) );
  INV_X1 U5446 ( .A(n4497), .ZN(n4495) );
  AND2_X1 U5447 ( .A1(n9153), .A2(n4459), .ZN(n9091) );
  NOR2_X1 U5448 ( .A1(n4460), .A2(n9295), .ZN(n4459) );
  INV_X1 U5449 ( .A(n4461), .ZN(n4460) );
  AND2_X1 U5450 ( .A1(n7465), .A2(n5909), .ZN(n4637) );
  NAND2_X1 U5451 ( .A1(n4635), .A2(n7522), .ZN(n4634) );
  NAND2_X1 U5452 ( .A1(n7465), .A2(n4636), .ZN(n4635) );
  AND2_X1 U5453 ( .A1(n9086), .A2(n9085), .ZN(n7842) );
  NAND2_X1 U5454 ( .A1(n9108), .A2(n9656), .ZN(n9110) );
  NAND2_X1 U5455 ( .A1(n9153), .A2(n4461), .ZN(n9099) );
  AND4_X1 U5456 ( .A1(n5859), .A2(n5858), .A3(n5857), .A4(n5856), .ZN(n9123)
         );
  NAND2_X1 U5457 ( .A1(n9139), .A2(n4638), .ZN(n9105) );
  AND2_X1 U5458 ( .A1(n9139), .A2(n7463), .ZN(n9126) );
  NAND2_X1 U5459 ( .A1(n9153), .A2(n8913), .ZN(n9143) );
  AND2_X1 U5460 ( .A1(n9309), .A2(n9162), .ZN(n5837) );
  NAND2_X1 U5461 ( .A1(n4625), .A2(n4623), .ZN(n9158) );
  AOI21_X1 U5462 ( .B1(n4626), .B2(n4628), .A(n4624), .ZN(n4623) );
  NOR2_X1 U5463 ( .A1(n9313), .A2(n9168), .ZN(n9153) );
  AND2_X1 U5464 ( .A1(n7603), .A2(n9204), .ZN(n9227) );
  NAND2_X1 U5465 ( .A1(n9471), .A2(n4271), .ZN(n9246) );
  INV_X1 U5466 ( .A(n9255), .ZN(n5765) );
  NAND2_X1 U5467 ( .A1(n9471), .A2(n4448), .ZN(n9263) );
  NAND2_X1 U5468 ( .A1(n9471), .A2(n9490), .ZN(n9470) );
  AND4_X1 U5469 ( .A1(n5683), .A2(n5682), .A3(n5681), .A4(n5680), .ZN(n7236)
         );
  AND4_X1 U5470 ( .A1(n5694), .A2(n5693), .A3(n5692), .A4(n5691), .ZN(n7472)
         );
  NAND2_X1 U5471 ( .A1(n4633), .A2(n7577), .ZN(n7233) );
  AND3_X1 U5472 ( .A1(n6977), .A2(n4270), .A3(n6530), .ZN(n7035) );
  OR2_X1 U5473 ( .A1(n5649), .A2(n6915), .ZN(n5663) );
  NAND2_X1 U5474 ( .A1(n4614), .A2(n4612), .ZN(n6748) );
  AOI21_X1 U5475 ( .B1(n4615), .B2(n4617), .A(n4613), .ZN(n4612) );
  INV_X1 U5476 ( .A(n7557), .ZN(n4613) );
  AND4_X1 U5477 ( .A1(n5668), .A2(n5667), .A3(n5666), .A4(n5665), .ZN(n6870)
         );
  NAND2_X1 U5478 ( .A1(n6530), .A2(n4265), .ZN(n9661) );
  NAND2_X1 U5479 ( .A1(n6530), .A2(n6529), .ZN(n9660) );
  AND4_X1 U5480 ( .A1(n5640), .A2(n5639), .A3(n5638), .A4(n5637), .ZN(n6809)
         );
  AND4_X1 U5481 ( .A1(n5611), .A2(n5610), .A3(n5609), .A4(n5608), .ZN(n6609)
         );
  NAND2_X1 U5482 ( .A1(n4468), .A2(n6305), .ZN(n6274) );
  NAND2_X1 U5483 ( .A1(n6305), .A2(n9683), .ZN(n6304) );
  INV_X1 U5484 ( .A(n6252), .ZN(n7431) );
  NAND2_X1 U5485 ( .A1(n5534), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n4619) );
  OR2_X1 U5486 ( .A1(n6287), .A2(n6286), .ZN(n9713) );
  NAND2_X1 U5487 ( .A1(n4642), .A2(n5504), .ZN(n4641) );
  INV_X1 U5488 ( .A(n4643), .ZN(n4642) );
  NAND2_X1 U5489 ( .A1(n5501), .A2(n5496), .ZN(n4643) );
  XNOR2_X1 U5490 ( .A(n7424), .B(n7423), .ZN(n7889) );
  AND3_X2 U5491 ( .A1(n5542), .A2(n5487), .A3(n5543), .ZN(n4629) );
  AND2_X1 U5492 ( .A1(n4283), .A2(n4630), .ZN(n4466) );
  NOR2_X1 U5493 ( .A1(n5931), .A2(n5878), .ZN(n5879) );
  XNOR2_X1 U5494 ( .A(n5237), .B(n5256), .ZN(n6517) );
  AND2_X1 U5495 ( .A1(n5236), .A2(n5257), .ZN(n5237) );
  XNOR2_X1 U5496 ( .A(n5155), .B(n5173), .ZN(n6559) );
  OAI21_X1 U5497 ( .B1(n4645), .B2(n4650), .A(n4946), .ZN(n4959) );
  NAND2_X1 U5498 ( .A1(n4652), .A2(n4653), .ZN(n4920) );
  AOI21_X1 U5499 ( .B1(n4892), .B2(n4654), .A(n4299), .ZN(n4653) );
  XNOR2_X1 U5500 ( .A(n4921), .B(SI_7_), .ZN(n4919) );
  OR2_X1 U5501 ( .A1(n5542), .A2(n5878), .ZN(n5571) );
  NAND2_X1 U5502 ( .A1(n8082), .A2(n4883), .ZN(n6817) );
  AND4_X1 U5503 ( .A1(n4868), .A2(n4867), .A3(n4866), .A4(n4865), .ZN(n7091)
         );
  NAND2_X1 U5504 ( .A1(n5388), .A2(n5387), .ZN(n8779) );
  XNOR2_X1 U5505 ( .A(n5321), .B(n5320), .ZN(n7962) );
  NAND2_X1 U5506 ( .A1(n4355), .A2(n4360), .ZN(n5460) );
  AOI21_X1 U5507 ( .B1(n4358), .B2(n4360), .A(n4357), .ZN(n4356) );
  INV_X1 U5508 ( .A(n4360), .ZN(n4359) );
  INV_X1 U5509 ( .A(n4362), .ZN(n4358) );
  AND4_X1 U5510 ( .A1(n4998), .A2(n4997), .A3(n4996), .A4(n4995), .ZN(n7328)
         );
  NAND2_X1 U5511 ( .A1(n4861), .A2(n4860), .ZN(n8083) );
  NAND2_X1 U5512 ( .A1(n5113), .A2(n5112), .ZN(n8675) );
  NAND2_X1 U5513 ( .A1(n5306), .A2(n5305), .ZN(n8550) );
  AND4_X1 U5514 ( .A1(n4978), .A2(n4977), .A3(n4976), .A4(n4975), .ZN(n7062)
         );
  NAND2_X1 U5515 ( .A1(n7865), .A2(n5198), .ZN(n8055) );
  AND4_X1 U5516 ( .A1(n5039), .A2(n5038), .A3(n5037), .A4(n5036), .ZN(n7306)
         );
  OR2_X1 U5517 ( .A1(n7042), .A2(n7041), .ZN(n4371) );
  INV_X1 U5518 ( .A(n8069), .ZN(n8059) );
  AND2_X1 U5519 ( .A1(n4812), .A2(n4768), .ZN(n6568) );
  AND2_X1 U5520 ( .A1(n6578), .A2(n4810), .ZN(n6569) );
  AND4_X1 U5521 ( .A1(n5192), .A2(n5191), .A3(n5190), .A4(n5189), .ZN(n8651)
         );
  AND4_X1 U5522 ( .A1(n5121), .A2(n5120), .A3(n5119), .A4(n5118), .ZN(n8649)
         );
  OR2_X1 U5523 ( .A1(n7998), .A2(n8650), .ZN(n8068) );
  NAND2_X1 U5524 ( .A1(n5360), .A2(n5359), .ZN(n8786) );
  INV_X1 U5525 ( .A(n6958), .ZN(n8322) );
  AND2_X1 U5526 ( .A1(n4403), .A2(n4402), .ZN(n4401) );
  NAND2_X1 U5527 ( .A1(n4814), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4805) );
  NOR2_X1 U5528 ( .A1(n9377), .A2(n4282), .ZN(n8331) );
  NOR2_X1 U5529 ( .A1(n8331), .A2(n8330), .ZN(n8329) );
  NOR2_X1 U5530 ( .A1(n6361), .A2(n4479), .ZN(n8343) );
  NOR2_X1 U5531 ( .A1(n6359), .A2(n4480), .ZN(n4479) );
  NOR2_X1 U5532 ( .A1(n8343), .A2(n8342), .ZN(n8341) );
  NAND2_X1 U5533 ( .A1(n4478), .A2(n4320), .ZN(n6401) );
  INV_X1 U5534 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4754) );
  AOI21_X1 U5535 ( .B1(n7909), .B2(n9748), .A(n7908), .ZN(n8770) );
  NAND2_X1 U5536 ( .A1(n7907), .A2(n7906), .ZN(n7908) );
  AND2_X1 U5537 ( .A1(n7911), .A2(n8465), .ZN(n8768) );
  AND2_X1 U5538 ( .A1(n8475), .A2(n8474), .ZN(n8776) );
  NAND2_X1 U5539 ( .A1(n8471), .A2(n8470), .ZN(n8469) );
  NAND2_X1 U5540 ( .A1(n4393), .A2(n4392), .ZN(n8564) );
  AND2_X1 U5541 ( .A1(n4393), .A2(n4263), .ZN(n8566) );
  NAND2_X1 U5542 ( .A1(n4394), .A2(n8577), .ZN(n4393) );
  NAND2_X1 U5543 ( .A1(n4686), .A2(n8217), .ZN(n8578) );
  NAND2_X1 U5544 ( .A1(n4398), .A2(n4399), .ZN(n8622) );
  OR2_X1 U5545 ( .A1(n8640), .A2(n7931), .ZN(n4398) );
  NAND2_X1 U5546 ( .A1(n5186), .A2(n5185), .ZN(n8824) );
  AND2_X1 U5547 ( .A1(n7070), .A2(n8832), .ZN(n9755) );
  AND2_X1 U5548 ( .A1(n7177), .A2(n7176), .ZN(n7179) );
  NAND2_X1 U5549 ( .A1(n7075), .A2(n7074), .ZN(n7076) );
  NAND2_X1 U5550 ( .A1(n4970), .A2(n4969), .ZN(n9844) );
  NAND2_X1 U5551 ( .A1(n9816), .A2(n6948), .ZN(n7084) );
  NAND2_X1 U5552 ( .A1(n6781), .A2(n4408), .ZN(n9816) );
  NOR2_X1 U5553 ( .A1(n6955), .A2(n4409), .ZN(n4408) );
  INV_X1 U5554 ( .A(n6780), .ZN(n4409) );
  NAND2_X1 U5555 ( .A1(n6781), .A2(n6780), .ZN(n6782) );
  NAND2_X1 U5556 ( .A1(n7027), .A2(n6688), .ZN(n9753) );
  INV_X1 U5557 ( .A(n9758), .ZN(n8743) );
  AND2_X1 U5558 ( .A1(n6000), .A2(n5453), .ZN(n9750) );
  OR2_X1 U5559 ( .A1(n9762), .A2(n6696), .ZN(n9758) );
  INV_X1 U5560 ( .A(n9753), .ZN(n8722) );
  NAND2_X1 U5561 ( .A1(n8753), .A2(n8752), .ZN(n8839) );
  NAND2_X1 U5562 ( .A1(n8749), .A2(n8832), .ZN(n8753) );
  OAI21_X1 U5563 ( .B1(n8750), .B2(n9859), .A(n8762), .ZN(n8751) );
  OAI21_X1 U5564 ( .B1(n8771), .B2(n9807), .A(n4387), .ZN(n8841) );
  AND2_X1 U5565 ( .A1(n8770), .A2(n8769), .ZN(n4387) );
  AOI22_X1 U5566 ( .A1(n8768), .A2(n8832), .B1(n9843), .B2(n8767), .ZN(n8769)
         );
  OR3_X1 U5567 ( .A1(n8823), .A2(n8822), .A3(n8821), .ZN(n8850) );
  NOR2_X1 U5568 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n4413) );
  XNOR2_X1 U5569 ( .A(n5432), .B(P2_IR_REG_24__SCAN_IN), .ZN(n6789) );
  OR2_X1 U5570 ( .A1(n4738), .A2(n4737), .ZN(n4740) );
  NAND2_X1 U5571 ( .A1(n4302), .A2(P2_IR_REG_0__SCAN_IN), .ZN(n4477) );
  OAI21_X1 U5572 ( .B1(n4568), .B2(n8982), .A(n4562), .ZN(n8857) );
  NAND2_X1 U5573 ( .A1(n4558), .A2(n4564), .ZN(n8856) );
  INV_X1 U5574 ( .A(n4563), .ZN(n4562) );
  NAND2_X1 U5575 ( .A1(n8870), .A2(n8868), .ZN(n8867) );
  AOI21_X1 U5576 ( .B1(n4564), .B2(n4561), .A(n4560), .ZN(n4559) );
  INV_X1 U5577 ( .A(n7819), .ZN(n4560) );
  NAND2_X1 U5578 ( .A1(n5500), .A2(n5499), .ZN(n9077) );
  NAND2_X1 U5579 ( .A1(n8927), .A2(n8931), .ZN(n8886) );
  NAND2_X1 U5580 ( .A1(n5839), .A2(n5838), .ZN(n9303) );
  NAND2_X1 U5581 ( .A1(n5700), .A2(n5699), .ZN(n7256) );
  NAND2_X1 U5582 ( .A1(n5809), .A2(n5808), .ZN(n9318) );
  AND2_X1 U5583 ( .A1(n6200), .A2(n6199), .ZN(n8985) );
  AND2_X1 U5584 ( .A1(n6200), .A2(n5916), .ZN(n8986) );
  AND2_X1 U5585 ( .A1(n6209), .A2(n6208), .ZN(n8989) );
  INV_X1 U5586 ( .A(n8993), .ZN(n8969) );
  AND2_X1 U5587 ( .A1(n6173), .A2(n9345), .ZN(n8991) );
  OR2_X1 U5588 ( .A1(n5730), .A2(n5729), .ZN(n8997) );
  OR2_X1 U5589 ( .A1(n5537), .A2(n5564), .ZN(n5569) );
  OAI211_X1 U5590 ( .C1(n4424), .C2(n4422), .A(n4420), .B(n4419), .ZN(n9018)
         );
  NAND2_X1 U5591 ( .A1(n4421), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n4420) );
  INV_X1 U5592 ( .A(n4423), .ZN(n4421) );
  NAND2_X1 U5593 ( .A1(n9018), .A2(n9017), .ZN(n9016) );
  NAND2_X1 U5594 ( .A1(n4444), .A2(n4443), .ZN(n9015) );
  INV_X1 U5595 ( .A(n9013), .ZN(n4443) );
  INV_X1 U5596 ( .A(n4445), .ZN(n4444) );
  NAND2_X1 U5597 ( .A1(n4445), .A2(n9013), .ZN(n9014) );
  NAND2_X1 U5598 ( .A1(n9026), .A2(n4288), .ZN(n9508) );
  NAND2_X1 U5599 ( .A1(n9516), .A2(n9515), .ZN(n9514) );
  AND2_X1 U5600 ( .A1(n9029), .A2(n4458), .ZN(n9516) );
  INV_X1 U5601 ( .A(n6056), .ZN(n4458) );
  INV_X1 U5602 ( .A(n4470), .ZN(n6223) );
  AND2_X1 U5603 ( .A1(n4470), .A2(n4313), .ZN(n9530) );
  INV_X1 U5604 ( .A(n4417), .ZN(n9546) );
  INV_X1 U5605 ( .A(n4442), .ZN(n9552) );
  AND2_X1 U5606 ( .A1(n4442), .A2(n4441), .ZN(n6229) );
  NAND2_X1 U5607 ( .A1(n6227), .A2(n6226), .ZN(n4441) );
  INV_X1 U5608 ( .A(n4440), .ZN(n6838) );
  INV_X1 U5609 ( .A(n4454), .ZN(n9584) );
  INV_X1 U5610 ( .A(n4432), .ZN(n9578) );
  AND2_X1 U5611 ( .A1(n4454), .A2(n4453), .ZN(n6843) );
  NAND2_X1 U5612 ( .A1(n6852), .A2(n6841), .ZN(n4453) );
  INV_X1 U5613 ( .A(n4452), .ZN(n9046) );
  AND2_X1 U5614 ( .A1(n4433), .A2(n4438), .ZN(n6856) );
  NAND2_X1 U5615 ( .A1(n4432), .A2(n4318), .ZN(n4433) );
  INV_X1 U5616 ( .A(n6853), .ZN(n4437) );
  INV_X1 U5617 ( .A(n4429), .ZN(n9617) );
  INV_X1 U5618 ( .A(n4427), .ZN(n9615) );
  NAND2_X1 U5619 ( .A1(n4499), .A2(n4500), .ZN(n5872) );
  NAND2_X1 U5620 ( .A1(n5924), .A2(n5923), .ZN(n9081) );
  NOR2_X1 U5621 ( .A1(n5922), .A2(n4699), .ZN(n5923) );
  NAND2_X1 U5622 ( .A1(n4501), .A2(n7451), .ZN(n9084) );
  NAND2_X1 U5623 ( .A1(n9187), .A2(n7611), .ZN(n9174) );
  AND2_X1 U5624 ( .A1(n9198), .A2(n5807), .ZN(n9166) );
  NAND2_X1 U5625 ( .A1(n4511), .A2(n5754), .ZN(n9256) );
  NAND2_X1 U5626 ( .A1(n7349), .A2(n7590), .ZN(n9271) );
  NAND2_X1 U5627 ( .A1(n5735), .A2(n5734), .ZN(n7358) );
  NAND2_X1 U5628 ( .A1(n5687), .A2(n5686), .ZN(n7473) );
  INV_X1 U5629 ( .A(n9484), .ZN(n9663) );
  NAND2_X1 U5630 ( .A1(n6501), .A2(n5612), .ZN(n6526) );
  NAND2_X1 U5631 ( .A1(n4632), .A2(n7483), .ZN(n6506) );
  NAND2_X1 U5632 ( .A1(n6312), .A2(n5588), .ZN(n6451) );
  OR2_X1 U5633 ( .A1(n6023), .A2(n5613), .ZN(n4513) );
  MUX2_X1 U5634 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9374), .S(n5531), .Z(n6289) );
  INV_X1 U5635 ( .A(n9268), .ZN(n9669) );
  INV_X1 U5636 ( .A(n9731), .ZN(n9729) );
  NOR2_X1 U5637 ( .A1(n4472), .A2(n9288), .ZN(n9291) );
  NAND2_X1 U5638 ( .A1(n9290), .A2(n4473), .ZN(n4472) );
  INV_X1 U5639 ( .A(n5512), .ZN(n7849) );
  NAND2_X1 U5640 ( .A1(n4655), .A2(n4875), .ZN(n4893) );
  NAND2_X1 U5641 ( .A1(n4872), .A2(n4871), .ZN(n4655) );
  OAI21_X1 U5642 ( .B1(n5571), .B2(n5543), .A(n5557), .ZN(n6139) );
  AOI211_X1 U5643 ( .C1(n7871), .C2(n8101), .A(n7374), .B(n7373), .ZN(n7375)
         );
  INV_X1 U5644 ( .A(n4486), .ZN(n8417) );
  NAND2_X1 U5645 ( .A1(n4386), .A2(n4385), .ZN(P2_U3549) );
  NAND2_X1 U5646 ( .A1(n9884), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n4385) );
  NAND2_X1 U5647 ( .A1(n8841), .A2(n4256), .ZN(n4386) );
  NAND2_X1 U5648 ( .A1(n4349), .A2(n4348), .ZN(P1_U3240) );
  OR2_X1 U5649 ( .A1(n7706), .A2(n7705), .ZN(n4348) );
  NAND2_X1 U5650 ( .A1(n4350), .A2(n7704), .ZN(n4349) );
  INV_X1 U5651 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9066) );
  MUX2_X1 U5652 ( .A(n9063), .B(n9062), .S(n9146), .Z(n9065) );
  AOI211_X1 U5653 ( .C1(n9288), .C2(n9248), .A(n7847), .B(n7846), .ZN(n7848)
         );
  NOR2_X1 U5654 ( .A1(n9301), .A2(n9274), .ZN(n9113) );
  NAND2_X1 U5655 ( .A1(n9359), .A2(n9731), .ZN(n5966) );
  AND2_X1 U5656 ( .A1(n7520), .A2(n7519), .ZN(n4261) );
  NAND2_X1 U5657 ( .A1(n7840), .A2(n7523), .ZN(n4262) );
  NAND3_X2 U5658 ( .A1(n4807), .A2(n4806), .A3(n4805), .ZN(n6691) );
  AND2_X1 U5659 ( .A1(n6151), .A2(n6299), .ZN(n6474) );
  INV_X2 U5660 ( .A(n6474), .ZN(n6195) );
  INV_X1 U5661 ( .A(n4629), .ZN(n5576) );
  NAND2_X1 U5662 ( .A1(n8576), .A2(n7985), .ZN(n4263) );
  NAND2_X1 U5663 ( .A1(n4382), .A2(n4708), .ZN(n4821) );
  INV_X1 U5664 ( .A(n8577), .ZN(n4390) );
  NAND2_X1 U5665 ( .A1(n9344), .A2(n9242), .ZN(n4264) );
  AND2_X1 U5666 ( .A1(n6529), .A2(n4456), .ZN(n4265) );
  AND2_X1 U5667 ( .A1(n4646), .A2(n4960), .ZN(n4266) );
  NAND2_X1 U5668 ( .A1(n5159), .A2(n5158), .ZN(n8831) );
  INV_X1 U5669 ( .A(n8565), .ZN(n4594) );
  AND2_X1 U5670 ( .A1(n9801), .A2(n9810), .ZN(n4267) );
  AND2_X1 U5671 ( .A1(n4520), .A2(n8576), .ZN(n4268) );
  XOR2_X1 U5672 ( .A(n8323), .B(n9823), .Z(n4269) );
  AND3_X1 U5673 ( .A1(n5546), .A2(n5545), .A3(n5544), .ZN(n6676) );
  INV_X1 U5674 ( .A(n6676), .ZN(n5547) );
  INV_X1 U5675 ( .A(n6496), .ZN(n6275) );
  AND2_X1 U5676 ( .A1(n4265), .A2(n4455), .ZN(n4270) );
  AND2_X1 U5677 ( .A1(n4448), .A2(n4447), .ZN(n4271) );
  NAND2_X1 U5678 ( .A1(n5213), .A2(n5212), .ZN(n8613) );
  AND2_X1 U5679 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4272) );
  AND2_X1 U5680 ( .A1(n4593), .A2(n4303), .ZN(n4273) );
  OR2_X1 U5681 ( .A1(n8767), .A2(n7893), .ZN(n8255) );
  AND2_X1 U5682 ( .A1(n4527), .A2(n4528), .ZN(n4274) );
  AND2_X1 U5683 ( .A1(n4399), .A2(n4290), .ZN(n4275) );
  OR2_X1 U5684 ( .A1(n8738), .A2(n4525), .ZN(n4276) );
  INV_X1 U5685 ( .A(n9146), .ZN(n9473) );
  XNOR2_X1 U5686 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6359), .ZN(n4277) );
  NAND3_X1 U5687 ( .A1(n7616), .A2(n7469), .A3(n7611), .ZN(n4278) );
  AND2_X1 U5688 ( .A1(n9107), .A2(n7630), .ZN(n4279) );
  AND2_X1 U5689 ( .A1(n4630), .A2(n4629), .ZN(n5645) );
  INV_X1 U5690 ( .A(n4400), .ZN(n6933) );
  AND2_X1 U5691 ( .A1(n4686), .A2(n4684), .ZN(n4280) );
  NAND2_X1 U5692 ( .A1(n5033), .A2(n5032), .ZN(n7170) );
  INV_X1 U5693 ( .A(n4662), .ZN(n8726) );
  NAND2_X1 U5694 ( .A1(n7872), .A2(n8705), .ZN(n4662) );
  NOR2_X1 U5695 ( .A1(n4819), .A2(n4576), .ZN(n4869) );
  NOR2_X1 U5696 ( .A1(n6648), .A2(n6644), .ZN(n4281) );
  AND2_X1 U5697 ( .A1(n9381), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4282) );
  NAND2_X1 U5698 ( .A1(n5944), .A2(n5943), .ZN(n6151) );
  NAND4_X1 U5699 ( .A1(n4791), .A2(n4790), .A3(n4789), .A4(n4788), .ZN(n6702)
         );
  NAND2_X2 U5700 ( .A1(n5512), .A2(n7708), .ZN(n5549) );
  INV_X1 U5701 ( .A(n8682), .ZN(n4607) );
  NAND2_X1 U5702 ( .A1(n7640), .A2(n7512), .ZN(n7843) );
  AND4_X1 U5703 ( .A1(n4538), .A2(n5488), .A3(n5696), .A4(n5671), .ZN(n4283)
         );
  NOR2_X2 U5704 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5542) );
  OR2_X1 U5705 ( .A1(n8256), .A2(n4590), .ZN(n4284) );
  AND4_X1 U5706 ( .A1(n5521), .A2(n5520), .A3(n5519), .A4(n5518), .ZN(n5532)
         );
  INV_X1 U5707 ( .A(n8576), .ZN(n8807) );
  AND2_X1 U5708 ( .A1(n8255), .A2(n4668), .ZN(n4285) );
  NAND2_X1 U5709 ( .A1(n5239), .A2(n5238), .ZN(n8812) );
  INV_X1 U5710 ( .A(n4508), .ZN(n4507) );
  OAI21_X1 U5711 ( .B1(n5818), .B2(n5807), .A(n4509), .ZN(n4508) );
  INV_X1 U5712 ( .A(n7646), .ZN(n4347) );
  NAND2_X1 U5713 ( .A1(n5852), .A2(n5851), .ZN(n9299) );
  NAND2_X1 U5714 ( .A1(n5830), .A2(n5829), .ZN(n9309) );
  NAND2_X1 U5715 ( .A1(n5747), .A2(n5746), .ZN(n9344) );
  AND2_X1 U5716 ( .A1(n4585), .A2(n4580), .ZN(n4286) );
  OR2_X1 U5717 ( .A1(n9295), .A2(n7813), .ZN(n7637) );
  NAND2_X1 U5718 ( .A1(n9153), .A2(n4463), .ZN(n4464) );
  AND2_X1 U5719 ( .A1(n8220), .A2(n4595), .ZN(n4287) );
  INV_X1 U5720 ( .A(n8693), .ZN(n9436) );
  NAND2_X1 U5721 ( .A1(n5076), .A2(n5075), .ZN(n8693) );
  INV_X1 U5722 ( .A(n7210), .ZN(n9490) );
  NAND2_X1 U5723 ( .A1(n5723), .A2(n5722), .ZN(n7210) );
  OR2_X1 U5724 ( .A1(n9025), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n4288) );
  OR2_X1 U5725 ( .A1(n4495), .A2(n7453), .ZN(n4289) );
  NAND2_X1 U5726 ( .A1(n8824), .A2(n8608), .ZN(n4290) );
  INV_X1 U5727 ( .A(n8534), .ZN(n8791) );
  NAND2_X1 U5728 ( .A1(n5345), .A2(n5344), .ZN(n8534) );
  NAND2_X1 U5729 ( .A1(n8233), .A2(n8236), .ZN(n8518) );
  INV_X1 U5730 ( .A(n8518), .ZN(n4598) );
  AND2_X1 U5731 ( .A1(n7748), .A2(n7743), .ZN(n4291) );
  AND2_X1 U5732 ( .A1(n7495), .A2(n9646), .ZN(n7439) );
  AND2_X1 U5733 ( .A1(n7775), .A2(n7774), .ZN(n4292) );
  NOR2_X1 U5734 ( .A1(n7915), .A2(n8472), .ZN(n8251) );
  INV_X1 U5735 ( .A(n4565), .ZN(n4564) );
  NAND2_X1 U5736 ( .A1(n8858), .A2(n4566), .ZN(n4565) );
  AND2_X1 U5737 ( .A1(n8802), .A2(n8315), .ZN(n4293) );
  OR2_X1 U5738 ( .A1(n5770), .A2(n5769), .ZN(n4294) );
  AND3_X1 U5739 ( .A1(n5931), .A2(n5930), .A3(n5929), .ZN(n4295) );
  NOR2_X1 U5740 ( .A1(n9313), .A2(n9176), .ZN(n4296) );
  NAND2_X1 U5741 ( .A1(n4750), .A2(n4374), .ZN(n4819) );
  INV_X1 U5742 ( .A(n8723), .ZN(n4661) );
  OR2_X1 U5743 ( .A1(n7563), .A2(n7562), .ZN(n4297) );
  AND2_X1 U5744 ( .A1(n8252), .A2(n8248), .ZN(n8470) );
  INV_X1 U5745 ( .A(n8470), .ZN(n4667) );
  AND2_X1 U5746 ( .A1(n4741), .A2(n4735), .ZN(n4298) );
  AND2_X1 U5747 ( .A1(n4895), .A2(SI_6_), .ZN(n4299) );
  NAND2_X1 U5748 ( .A1(n7486), .A2(n7675), .ZN(n6270) );
  AND2_X1 U5749 ( .A1(n4693), .A2(n4602), .ZN(n4300) );
  AND2_X1 U5750 ( .A1(n4477), .A2(n4475), .ZN(n4301) );
  AND2_X1 U5751 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n4302) );
  OR2_X1 U5752 ( .A1(n8223), .A2(n4590), .ZN(n4303) );
  OR2_X1 U5753 ( .A1(n8675), .A2(n8649), .ZN(n8195) );
  AND2_X1 U5754 ( .A1(n9299), .A2(n9123), .ZN(n7521) );
  AND4_X1 U5755 ( .A1(n5054), .A2(n5053), .A3(n5052), .A4(n5051), .ZN(n8123)
         );
  INV_X1 U5756 ( .A(n8123), .ZN(n4663) );
  AND2_X1 U5757 ( .A1(n4499), .A2(n4497), .ZN(n4304) );
  AND2_X1 U5758 ( .A1(n5893), .A2(n7577), .ZN(n4305) );
  AND2_X1 U5759 ( .A1(n7438), .A2(n7483), .ZN(n4306) );
  AND2_X1 U5760 ( .A1(n4594), .A2(n8221), .ZN(n4307) );
  OR2_X1 U5761 ( .A1(n5770), .A2(n4572), .ZN(n4308) );
  AND2_X1 U5762 ( .A1(n8284), .A2(n7176), .ZN(n4309) );
  INV_X1 U5763 ( .A(n5040), .ZN(n4673) );
  AND2_X1 U5764 ( .A1(n5042), .A2(n5012), .ZN(n5040) );
  AND2_X1 U5765 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n4310) );
  INV_X1 U5766 ( .A(n7932), .ZN(n7933) );
  INV_X1 U5767 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4476) );
  INV_X1 U5768 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n4422) );
  INV_X1 U5769 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n4712) );
  INV_X1 U5770 ( .A(n9676), .ZN(n9666) );
  NAND2_X1 U5771 ( .A1(n5417), .A2(n5416), .ZN(n8773) );
  INV_X1 U5772 ( .A(n8773), .ZN(n4527) );
  AND4_X1 U5773 ( .A1(n4536), .A2(n4539), .A3(n5614), .A4(n5600), .ZN(n4311)
         );
  NAND2_X1 U5774 ( .A1(n7803), .A2(n7802), .ZN(n4312) );
  OAI211_X1 U5775 ( .C1(n5997), .C2(n6359), .A(n4831), .B(n4830), .ZN(n8042)
         );
  INV_X1 U5776 ( .A(n7590), .ZN(n4631) );
  OR2_X1 U5777 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6233), .ZN(n4313) );
  AND2_X1 U5778 ( .A1(n6363), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4314) );
  OR2_X1 U5779 ( .A1(n5013), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n4315) );
  NAND2_X1 U5780 ( .A1(n4711), .A2(n4372), .ZN(n5013) );
  NAND2_X1 U5781 ( .A1(n8606), .A2(n8605), .ZN(n8604) );
  NAND2_X1 U5782 ( .A1(n4629), .A2(n4311), .ZN(n5642) );
  NOR3_X1 U5783 ( .A1(n8738), .A2(n8831), .A3(n4525), .ZN(n4523) );
  AND4_X1 U5784 ( .A1(n5164), .A2(n5163), .A3(n5162), .A4(n5161), .ZN(n7930)
         );
  NAND2_X1 U5785 ( .A1(n7885), .A2(n8195), .ZN(n8645) );
  AND2_X1 U5786 ( .A1(n8631), .A2(n8819), .ZN(n8588) );
  INV_X1 U5787 ( .A(n5399), .ZN(n4365) );
  INV_X1 U5788 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n4375) );
  AND2_X1 U5789 ( .A1(n4680), .A2(n4681), .ZN(n4316) );
  INV_X1 U5790 ( .A(n8563), .ZN(n8802) );
  AND2_X1 U5791 ( .A1(n5301), .A2(n5300), .ZN(n8563) );
  INV_X1 U5792 ( .A(n4263), .ZN(n4395) );
  INV_X1 U5793 ( .A(n6854), .ZN(n4434) );
  INV_X1 U5794 ( .A(n9668), .ZN(n4456) );
  NAND2_X1 U5795 ( .A1(n5759), .A2(n5758), .ZN(n9251) );
  INV_X1 U5796 ( .A(n9251), .ZN(n4447) );
  NAND2_X1 U5797 ( .A1(n9471), .A2(n4450), .ZN(n4317) );
  OR2_X1 U5798 ( .A1(n9699), .A2(n9003), .ZN(n7679) );
  INV_X1 U5799 ( .A(n7679), .ZN(n4324) );
  NAND2_X1 U5800 ( .A1(n6530), .A2(n4270), .ZN(n4457) );
  AND2_X1 U5801 ( .A1(n4437), .A2(n4434), .ZN(n4318) );
  AND2_X1 U5802 ( .A1(n9683), .A2(n6676), .ZN(n4468) );
  NAND2_X1 U5803 ( .A1(n7659), .A2(n9473), .ZN(n7650) );
  INV_X1 U5804 ( .A(n7251), .ZN(n4517) );
  AND2_X1 U5805 ( .A1(n9607), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n4319) );
  NAND2_X1 U5806 ( .A1(n5648), .A2(n5647), .ZN(n9390) );
  INV_X1 U5807 ( .A(n9390), .ZN(n4455) );
  NAND2_X1 U5808 ( .A1(n6301), .A2(n6302), .ZN(n6300) );
  INV_X1 U5809 ( .A(n6691), .ZN(n6690) );
  OR2_X1 U5810 ( .A1(n6728), .A2(n9793), .ZN(n7131) );
  INV_X1 U5811 ( .A(n7131), .ZN(n4522) );
  OR2_X1 U5812 ( .A1(n8341), .A2(n4314), .ZN(n4478) );
  XNOR2_X1 U5813 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6404), .ZN(n4320) );
  NOR2_X1 U5814 ( .A1(n5497), .A2(n4641), .ZN(n7402) );
  OR2_X1 U5815 ( .A1(n8329), .A2(n4482), .ZN(n4481) );
  INV_X1 U5816 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n4480) );
  NOR2_X1 U5817 ( .A1(n8130), .A2(n8262), .ZN(n4586) );
  NAND2_X1 U5818 ( .A1(n8126), .A2(n8262), .ZN(n4588) );
  INV_X1 U5819 ( .A(n8262), .ZN(n4590) );
  NAND2_X1 U5820 ( .A1(n4325), .A2(n7540), .ZN(n7544) );
  NAND2_X1 U5821 ( .A1(n7539), .A2(n7538), .ZN(n4325) );
  AOI21_X1 U5822 ( .B1(n7607), .B2(n4338), .A(n4335), .ZN(n7613) );
  OAI211_X1 U5823 ( .C1(n7487), .C2(n4353), .A(n7671), .B(n4352), .ZN(n7527)
         );
  NAND2_X1 U5824 ( .A1(n6431), .A2(n7675), .ZN(n7526) );
  NAND2_X1 U5825 ( .A1(n7487), .A2(n7433), .ZN(n6431) );
  NAND2_X1 U5826 ( .A1(n5887), .A2(n7666), .ZN(n7487) );
  NAND2_X2 U5827 ( .A1(n5916), .A2(n6046), .ZN(n5531) );
  XNOR2_X2 U5828 ( .A(n4354), .B(n5496), .ZN(n6046) );
  NAND2_X1 U5829 ( .A1(n5497), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4354) );
  NAND2_X1 U5830 ( .A1(n5378), .A2(n4362), .ZN(n4355) );
  NAND2_X1 U5831 ( .A1(n5378), .A2(n5377), .ZN(n7951) );
  OAI21_X1 U5832 ( .B1(n5378), .B2(n4359), .A(n4356), .ZN(n4364) );
  NAND2_X1 U5833 ( .A1(n4364), .A2(n5466), .ZN(n5485) );
  NAND2_X1 U5834 ( .A1(n6830), .A2(n4935), .ZN(n5976) );
  INV_X1 U5835 ( .A(n4576), .ZN(n4373) );
  INV_X1 U5836 ( .A(n5410), .ZN(n5302) );
  NAND2_X1 U5837 ( .A1(n5331), .A2(n4377), .ZN(n8092) );
  AND2_X1 U5838 ( .A1(n5332), .A2(n4378), .ZN(n4377) );
  NAND2_X1 U5839 ( .A1(n5331), .A2(n5332), .ZN(n4379) );
  MUX2_X1 U5840 ( .A(n7995), .B(n7994), .S(n4379), .Z(n7996) );
  NAND2_X1 U5841 ( .A1(n7865), .A2(n4381), .ZN(n8053) );
  NAND2_X2 U5842 ( .A1(n7854), .A2(n5194), .ZN(n7865) );
  XNOR2_X2 U5843 ( .A(n4744), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8511) );
  NAND2_X1 U5844 ( .A1(n4712), .A2(n4602), .ZN(n4384) );
  INV_X1 U5845 ( .A(n4819), .ZN(n4382) );
  AND4_X2 U5846 ( .A1(n4711), .A2(n4383), .A3(n4693), .A4(n4382), .ZN(n5419)
         );
  OAI22_X1 U5847 ( .A1(n8640), .A2(n4396), .B1(n7933), .B2(n4275), .ZN(n8617)
         );
  NAND3_X1 U5848 ( .A1(n4817), .A2(n4818), .A3(n4401), .ZN(n4400) );
  NAND2_X1 U5849 ( .A1(n7177), .A2(n4309), .ZN(n7312) );
  NAND2_X1 U5850 ( .A1(n7312), .A2(n4411), .ZN(n4410) );
  NAND2_X1 U5851 ( .A1(n7921), .A2(n4410), .ZN(n8668) );
  NAND2_X1 U5852 ( .A1(n4745), .A2(n4746), .ZN(n4724) );
  NAND2_X1 U5853 ( .A1(n4745), .A2(n4413), .ZN(n7397) );
  NAND3_X1 U5854 ( .A1(n6773), .A2(n8124), .A3(n6930), .ZN(n6771) );
  NAND3_X1 U5855 ( .A1(n4424), .A2(n4423), .A3(n4422), .ZN(n4419) );
  OAI21_X1 U5856 ( .B1(n9577), .B2(n6853), .A(n4435), .ZN(n4438) );
  INV_X1 U5857 ( .A(n4438), .ZN(n9037) );
  XNOR2_X1 U5858 ( .A(n8326), .B(n9793), .ZN(n6769) );
  NOR2_X1 U5859 ( .A1(n9604), .A2(n9603), .ZN(n9602) );
  MUX2_X1 U5860 ( .A(n7583), .B(n7582), .S(n7650), .Z(n7588) );
  NAND2_X1 U5861 ( .A1(n7542), .A2(n7650), .ZN(n7550) );
  AND3_X2 U5862 ( .A1(n4283), .A2(n4630), .A3(n4629), .ZN(n5732) );
  OAI21_X1 U5863 ( .B1(n7597), .B2(n7596), .A(n7595), .ZN(n7607) );
  NAND2_X1 U5864 ( .A1(n7566), .A2(n7565), .ZN(n7568) );
  OR2_X2 U5865 ( .A1(n8022), .A2(n8018), .ZN(n7727) );
  NAND2_X1 U5866 ( .A1(n4647), .A2(n4649), .ZN(n4646) );
  OR2_X2 U5867 ( .A1(n5145), .A2(n7370), .ZN(n7716) );
  AND2_X1 U5868 ( .A1(n5146), .A2(n7716), .ZN(n5147) );
  NAND2_X2 U5869 ( .A1(n4986), .A2(n4985), .ZN(n5003) );
  INV_X1 U5870 ( .A(n4457), .ZN(n6976) );
  INV_X1 U5871 ( .A(n4464), .ZN(n9119) );
  NAND2_X1 U5872 ( .A1(n4465), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5498) );
  NAND3_X1 U5873 ( .A1(n4467), .A2(n5495), .A3(n4466), .ZN(n4465) );
  NAND2_X1 U5874 ( .A1(n5732), .A2(n5495), .ZN(n5497) );
  NAND3_X1 U5875 ( .A1(n4469), .A2(n4468), .A3(n6496), .ZN(n6439) );
  AOI211_X1 U5876 ( .C1(n7835), .C2(n9289), .A(n9714), .B(n9067), .ZN(n9288)
         );
  NAND2_X1 U5877 ( .A1(n9289), .A2(n9345), .ZN(n4473) );
  MUX2_X1 U5878 ( .A(n5983), .B(P2_REG2_REG_1__SCAN_IN), .S(n6335), .Z(n5984)
         );
  NAND2_X2 U5879 ( .A1(n4691), .A2(n4690), .ZN(n4781) );
  NAND3_X1 U5880 ( .A1(n4691), .A2(n4690), .A3(n4310), .ZN(n4491) );
  OR2_X2 U5881 ( .A1(n9098), .A2(n7453), .ZN(n4501) );
  NAND2_X1 U5882 ( .A1(n6501), .A2(n4502), .ZN(n6528) );
  OAI21_X1 U5883 ( .B1(n9198), .B2(n4505), .A(n4504), .ZN(n9135) );
  OAI21_X1 U5884 ( .B1(n9198), .B2(n5818), .A(n4507), .ZN(n9152) );
  OR2_X1 U5885 ( .A1(n9173), .A2(n8874), .ZN(n4509) );
  NAND2_X1 U5886 ( .A1(n6312), .A2(n4512), .ZN(n6449) );
  INV_X2 U5887 ( .A(n6714), .ZN(n9786) );
  NAND3_X1 U5888 ( .A1(n9773), .A2(n9778), .A3(n6714), .ZN(n6728) );
  OAI22_X1 U5889 ( .A1(n8110), .A2(n6009), .B1(n5997), .B2(n6010), .ZN(n4515)
         );
  AND3_X2 U5890 ( .A1(n4799), .A2(n4800), .A3(n4516), .ZN(n9778) );
  OR2_X1 U5891 ( .A1(n8110), .A2(n6011), .ZN(n4516) );
  NAND2_X1 U5892 ( .A1(n4522), .A2(n4521), .ZN(n7093) );
  INV_X1 U5893 ( .A(n4523), .ZN(n8641) );
  NAND2_X1 U5894 ( .A1(n8878), .A2(n4531), .ZN(n8880) );
  OR2_X1 U5895 ( .A1(n4532), .A2(n8879), .ZN(n4531) );
  NAND2_X1 U5896 ( .A1(n8950), .A2(n8952), .ZN(n4532) );
  NAND2_X1 U5897 ( .A1(n7142), .A2(n7141), .ZN(n7148) );
  NAND2_X1 U5898 ( .A1(n7142), .A2(n4534), .ZN(n7192) );
  OAI22_X2 U5899 ( .A1(n4543), .A2(n4541), .B1(n7788), .B2(n4542), .ZN(n8904)
         );
  NAND2_X1 U5900 ( .A1(n8938), .A2(n8941), .ZN(n4544) );
  NAND2_X1 U5901 ( .A1(n7783), .A2(n7782), .ZN(n8939) );
  NAND2_X4 U5902 ( .A1(n4547), .A2(n4545), .ZN(n7814) );
  INV_X1 U5903 ( .A(n6157), .ZN(n6178) );
  NAND2_X1 U5904 ( .A1(n6156), .A2(n6157), .ZN(n6180) );
  AND2_X1 U5905 ( .A1(n6152), .A2(n4548), .ZN(n6156) );
  NAND2_X1 U5906 ( .A1(n7744), .A2(n7743), .ZN(n7751) );
  NAND2_X1 U5907 ( .A1(n4549), .A2(n4550), .ZN(n7780) );
  NAND2_X1 U5908 ( .A1(n8928), .A2(n4551), .ZN(n4549) );
  NAND2_X1 U5909 ( .A1(n8894), .A2(n4556), .ZN(n4555) );
  NAND2_X1 U5910 ( .A1(n8894), .A2(n8895), .ZN(n4568) );
  NAND2_X1 U5911 ( .A1(n4555), .A2(n4559), .ZN(n7827) );
  AND2_X1 U5912 ( .A1(n4568), .A2(n4312), .ZN(n8984) );
  NAND2_X1 U5913 ( .A1(n5745), .A2(n5744), .ZN(n5770) );
  NOR4_X1 U5914 ( .A1(n4575), .A2(n4574), .A3(n8258), .A4(n8260), .ZN(n8267)
         );
  NAND2_X1 U5915 ( .A1(n4591), .A2(n8226), .ZN(n4600) );
  NAND2_X1 U5916 ( .A1(n4592), .A2(n4273), .ZN(n4591) );
  NAND2_X1 U5917 ( .A1(n8222), .A2(n4307), .ZN(n4592) );
  OAI21_X1 U5918 ( .B1(n6520), .B2(n4617), .A(n4615), .ZN(n6745) );
  NAND2_X1 U5919 ( .A1(n6520), .A2(n4615), .ZN(n4614) );
  AND3_X1 U5920 ( .A1(n4622), .A2(n4619), .A3(n4618), .ZN(n4621) );
  AND2_X2 U5921 ( .A1(n4621), .A2(n4620), .ZN(n6298) );
  NAND2_X1 U5922 ( .A1(n4252), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n4620) );
  NAND2_X1 U5923 ( .A1(n5906), .A2(n4626), .ZN(n4625) );
  AND2_X2 U5924 ( .A1(n4627), .A2(n4702), .ZN(n4626) );
  NAND2_X1 U5925 ( .A1(n4632), .A2(n4306), .ZN(n6504) );
  NAND2_X1 U5926 ( .A1(n4633), .A2(n4305), .ZN(n7235) );
  AOI21_X1 U5927 ( .B1(n9136), .B2(n4637), .A(n4634), .ZN(n9086) );
  NAND2_X1 U5928 ( .A1(n9136), .A2(n5909), .ZN(n9139) );
  OR2_X1 U5929 ( .A1(n5497), .A2(n4643), .ZN(n5503) );
  INV_X1 U5930 ( .A(n4924), .ZN(n4645) );
  AOI21_X2 U5931 ( .B1(n4650), .B2(n4946), .A(n4648), .ZN(n4647) );
  NAND2_X1 U5932 ( .A1(n4924), .A2(n4923), .ZN(n4947) );
  NAND2_X1 U5933 ( .A1(n4872), .A2(n4651), .ZN(n4652) );
  NAND2_X1 U5934 ( .A1(n8639), .A2(n8196), .ZN(n4657) );
  NAND2_X1 U5935 ( .A1(n4656), .A2(n8211), .ZN(n4658) );
  NAND2_X1 U5936 ( .A1(n7886), .A2(n4657), .ZN(n4656) );
  OAI21_X2 U5937 ( .B1(n7885), .B2(n4659), .A(n4658), .ZN(n8606) );
  NAND2_X1 U5938 ( .A1(n8486), .A2(n4668), .ZN(n4664) );
  NAND2_X1 U5939 ( .A1(n8486), .A2(n8241), .ZN(n8471) );
  NAND2_X1 U5940 ( .A1(n5003), .A2(n4677), .ZN(n4676) );
  NAND2_X1 U5941 ( .A1(n5003), .A2(n4670), .ZN(n4669) );
  OAI21_X1 U5942 ( .B1(n5003), .B2(n5002), .A(n5001), .ZN(n5029) );
  INV_X1 U5943 ( .A(n8596), .ZN(n4688) );
  AND2_X2 U5944 ( .A1(n4680), .A2(n4679), .ZN(n8543) );
  OR2_X2 U5945 ( .A1(n8596), .A2(n4683), .ZN(n4680) );
  NAND3_X1 U5946 ( .A1(n4754), .A2(n4753), .A3(n4752), .ZN(n4691) );
  INV_X1 U5947 ( .A(n5419), .ZN(n5073) );
  NAND2_X1 U5948 ( .A1(n7197), .A2(n7196), .ZN(n7274) );
  XNOR2_X1 U5949 ( .A(n4740), .B(n4739), .ZN(n5463) );
  CLKBUF_X1 U5950 ( .A(n7275), .Z(n7277) );
  AND2_X2 U5951 ( .A1(n5144), .A2(n7293), .ZN(n7370) );
  OR2_X2 U5952 ( .A1(n5143), .A2(n7288), .ZN(n7293) );
  OR2_X1 U5953 ( .A1(n5537), .A2(n5517), .ZN(n5520) );
  NAND2_X1 U5954 ( .A1(n4308), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5877) );
  INV_X1 U5955 ( .A(n6885), .ZN(n6889) );
  OR2_X1 U5956 ( .A1(n6885), .A2(n7051), .ZN(n6986) );
  OR2_X4 U5957 ( .A1(n9772), .A2(n8765), .ZN(n9861) );
  AND2_X2 U5958 ( .A1(n7286), .A2(n7320), .ZN(n5135) );
  NAND2_X1 U5959 ( .A1(n5169), .A2(n7729), .ZN(n7854) );
  INV_X1 U5960 ( .A(n6483), .ZN(n6619) );
  OAI22_X2 U5961 ( .A1(n9468), .A2(n5731), .B1(n9490), .B2(n7193), .ZN(n7359)
         );
  NAND2_X2 U5962 ( .A1(n8903), .A2(n7795), .ZN(n8894) );
  NAND2_X2 U5963 ( .A1(n7981), .A2(n5252), .ZN(n5287) );
  XNOR2_X2 U5964 ( .A(n8030), .B(n8029), .ZN(n8034) );
  INV_X1 U5965 ( .A(n7950), .ZN(n4729) );
  OR2_X1 U5966 ( .A1(n8838), .A2(n8760), .ZN(n9884) );
  AND3_X1 U5967 ( .A1(n8003), .A2(n8004), .A3(n8006), .ZN(n4692) );
  AND2_X1 U5968 ( .A1(n5082), .A2(n4713), .ZN(n4693) );
  OR2_X1 U5969 ( .A1(n9731), .A2(n5965), .ZN(n4694) );
  NOR2_X1 U5970 ( .A1(n7559), .A2(n7547), .ZN(n4695) );
  OR3_X1 U5971 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4696) );
  AND2_X1 U5972 ( .A1(n8143), .A2(n4269), .ZN(n4697) );
  INV_X1 U5973 ( .A(n4816), .ZN(n4769) );
  INV_X1 U5974 ( .A(n5463), .ZN(n8301) );
  AND2_X1 U5975 ( .A1(n4985), .A2(n4964), .ZN(n4698) );
  AND2_X1 U5976 ( .A1(n9656), .A2(n8996), .ZN(n4699) );
  INV_X1 U5977 ( .A(n8296), .ZN(n7894) );
  AND2_X1 U5978 ( .A1(n7516), .A2(n9280), .ZN(n4700) );
  AND2_X1 U5979 ( .A1(n4960), .A2(n4951), .ZN(n4701) );
  AND2_X1 U5980 ( .A1(n7614), .A2(n7616), .ZN(n4702) );
  AND2_X1 U5981 ( .A1(n5059), .A2(SI_14_), .ZN(n4703) );
  AND2_X1 U5982 ( .A1(n5831), .A2(n8907), .ZN(n4704) );
  NAND2_X1 U5983 ( .A1(n7052), .A2(n6888), .ZN(n4705) );
  OR2_X1 U5984 ( .A1(n8773), .A2(n8490), .ZN(n4706) );
  NOR2_X1 U5985 ( .A1(n5484), .A2(n5483), .ZN(n4707) );
  INV_X1 U5986 ( .A(n7470), .ZN(n5898) );
  INV_X1 U5987 ( .A(n7232), .ZN(n5893) );
  INV_X1 U5988 ( .A(n7650), .ZN(n7547) );
  NAND2_X1 U5989 ( .A1(n7548), .A2(n7547), .ZN(n7549) );
  NAND2_X1 U5990 ( .A1(n9270), .A2(n7592), .ZN(n7596) );
  AND2_X1 U5991 ( .A1(n7103), .A2(n6703), .ZN(n6700) );
  NOR2_X1 U5992 ( .A1(n8272), .A2(n6759), .ZN(n6760) );
  INV_X1 U5993 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n4713) );
  NAND2_X1 U5994 ( .A1(n4700), .A2(n7547), .ZN(n7651) );
  INV_X1 U5995 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n10031) );
  INV_X1 U5996 ( .A(n6644), .ZN(n6645) );
  NOR2_X1 U5997 ( .A1(n6610), .A2(n6611), .ZN(n6618) );
  NAND2_X1 U5998 ( .A1(n7652), .A2(n7651), .ZN(n7653) );
  INV_X1 U5999 ( .A(n5116), .ZN(n5114) );
  INV_X1 U6000 ( .A(n5279), .ZN(n5277) );
  INV_X1 U6001 ( .A(n5034), .ZN(n5019) );
  INV_X1 U6002 ( .A(n8142), .ZN(n6954) );
  INV_X1 U6003 ( .A(n9778), .ZN(n6689) );
  INV_X1 U6004 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n4734) );
  NAND2_X1 U6005 ( .A1(n6889), .A2(n4705), .ZN(n6988) );
  INV_X1 U6006 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5605) );
  OR2_X1 U6007 ( .A1(n5904), .A2(n5903), .ZN(n5905) );
  OR2_X1 U6008 ( .A1(n5258), .A2(n5257), .ZN(n5267) );
  AND2_X1 U6009 ( .A1(n5203), .A2(n5202), .ZN(n5204) );
  NAND2_X1 U6010 ( .A1(n4949), .A2(n4948), .ZN(n4960) );
  OR2_X1 U6011 ( .A1(n5389), .A2(n7953), .ZN(n5401) );
  INV_X1 U6012 ( .A(n6816), .ZN(n4905) );
  INV_X1 U6013 ( .A(n8056), .ZN(n5228) );
  OR2_X1 U6014 ( .A1(n4993), .A2(n4992), .ZN(n5034) );
  NAND2_X1 U6015 ( .A1(n5277), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n5326) );
  OR2_X1 U6016 ( .A1(n8550), .A2(n8031), .ZN(n8228) );
  OR3_X1 U6017 ( .A1(n5187), .A2(n7735), .A3(n7860), .ZN(n5217) );
  OR2_X1 U6018 ( .A1(n5096), .A2(n5095), .ZN(n5116) );
  AND2_X1 U6019 ( .A1(n8142), .A2(n8141), .ZN(n6955) );
  AND2_X1 U6020 ( .A1(n7302), .A2(n7869), .ZN(n7304) );
  INV_X1 U6021 ( .A(n7147), .ZN(n7146) );
  OR2_X1 U6022 ( .A1(n5635), .A2(n5634), .ZN(n5649) );
  OR2_X1 U6023 ( .A1(n5810), .A2(n8942), .ZN(n5821) );
  INV_X1 U6024 ( .A(n7750), .ZN(n7748) );
  NAND2_X1 U6025 ( .A1(n5736), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5749) );
  AND2_X1 U6026 ( .A1(n5724), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5736) );
  NAND2_X1 U6027 ( .A1(n5380), .A2(n5379), .ZN(n5382) );
  OR2_X1 U6028 ( .A1(n5235), .A2(n5234), .ZN(n5257) );
  NAND2_X1 U6029 ( .A1(n5106), .A2(n5105), .ZN(n5108) );
  NAND2_X1 U6030 ( .A1(n5005), .A2(n9942), .ZN(n5008) );
  INV_X1 U6031 ( .A(n9823), .ZN(n8146) );
  INV_X1 U6032 ( .A(n6795), .ZN(n4860) );
  OR2_X1 U6033 ( .A1(n5326), .A2(n5309), .ZN(n5347) );
  NAND2_X1 U6034 ( .A1(n6365), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6366) );
  AND2_X1 U6035 ( .A1(n6354), .A2(n6353), .ZN(n6382) );
  AND2_X1 U6036 ( .A1(n8228), .A2(n8227), .ZN(n8542) );
  INV_X1 U6037 ( .A(n8812), .ZN(n8595) );
  INV_X1 U6038 ( .A(n9755), .ZN(n8745) );
  AND2_X1 U6039 ( .A1(n8269), .A2(n5461), .ZN(n9843) );
  AND2_X1 U6040 ( .A1(n9456), .A2(n8663), .ZN(n8735) );
  INV_X1 U6041 ( .A(n8730), .ZN(n8648) );
  OR2_X1 U6042 ( .A1(n5985), .A2(n5469), .ZN(n8650) );
  NOR2_X1 U6043 ( .A1(n5478), .A2(P2_U3152), .ZN(n6000) );
  OR2_X1 U6044 ( .A1(n4915), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n4917) );
  OR2_X1 U6045 ( .A1(n5821), .A2(n9972), .ZN(n5831) );
  XNOR2_X1 U6046 ( .A(n6198), .B(n7806), .ZN(n6469) );
  OR2_X1 U6047 ( .A1(n7794), .A2(n7793), .ZN(n7795) );
  NOR2_X1 U6048 ( .A1(n5831), .A2(n8907), .ZN(n5840) );
  AND2_X1 U6049 ( .A1(n5788), .A2(n5507), .ZN(n5799) );
  NAND2_X1 U6050 ( .A1(n5915), .A2(n9651), .ZN(n5924) );
  NAND2_X1 U6051 ( .A1(n5799), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5810) );
  OR2_X1 U6052 ( .A1(n7426), .A2(n6021), .ZN(n5525) );
  NAND2_X1 U6053 ( .A1(n5481), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8099) );
  INV_X1 U6054 ( .A(n8613), .ZN(n8819) );
  INV_X1 U6055 ( .A(n8099), .ZN(n8079) );
  AND2_X1 U6056 ( .A1(n5408), .A2(n5407), .ZN(n7954) );
  AND4_X1 U6057 ( .A1(n5247), .A2(n5246), .A3(n5245), .A4(n5244), .ZN(n8580)
         );
  NAND2_X1 U6058 ( .A1(n8354), .A2(n8355), .ZN(n8353) );
  INV_X1 U6059 ( .A(n9733), .ZN(n9738) );
  INV_X2 U6060 ( .A(n4952), .ZN(n8108) );
  INV_X1 U6061 ( .A(n8272), .ZN(n7127) );
  OR2_X1 U6062 ( .A1(n9768), .A2(n5444), .ZN(n8760) );
  INV_X1 U6063 ( .A(n8751), .ZN(n8752) );
  AND2_X1 U6064 ( .A1(n9791), .A2(n9847), .ZN(n9807) );
  OR2_X1 U6065 ( .A1(n7922), .A2(n8181), .ZN(n9456) );
  INV_X1 U6066 ( .A(n9807), .ZN(n9866) );
  AND2_X1 U6067 ( .A1(n7109), .A2(n5434), .ZN(n9763) );
  INV_X1 U6068 ( .A(n4726), .ZN(n4728) );
  AND2_X1 U6069 ( .A1(n4968), .A2(n4987), .ZN(n6549) );
  INV_X1 U6070 ( .A(n9713), .ZN(n9345) );
  AND4_X1 U6071 ( .A1(n5871), .A2(n5870), .A3(n5869), .A4(n5868), .ZN(n7813)
         );
  AND2_X1 U6072 ( .A1(n7637), .A2(n7523), .ZN(n9085) );
  INV_X1 U6073 ( .A(n6448), .ZN(n7540) );
  INV_X1 U6074 ( .A(n9212), .ZN(n9654) );
  AND2_X1 U6075 ( .A1(n5940), .A2(n5939), .ZN(n6281) );
  INV_X1 U6076 ( .A(n9736), .ZN(n9376) );
  AND2_X1 U6077 ( .A1(n5276), .A2(n5275), .ZN(n8576) );
  INV_X1 U6078 ( .A(n8085), .ZN(n8103) );
  INV_X1 U6079 ( .A(n8101), .ZN(n8074) );
  OR2_X1 U6080 ( .A1(n5993), .A2(n8307), .ZN(n9740) );
  INV_X1 U6081 ( .A(n8459), .ZN(n8750) );
  AND2_X1 U6082 ( .A1(n8492), .A2(n8491), .ZN(n8782) );
  INV_X1 U6083 ( .A(n6962), .ZN(n8655) );
  AND2_X1 U6084 ( .A1(n6683), .A2(n8739), .ZN(n9762) );
  OR2_X1 U6085 ( .A1(n8838), .A2(n8837), .ZN(n9867) );
  INV_X1 U6086 ( .A(n9765), .ZN(n10021) );
  OR2_X1 U6087 ( .A1(n5741), .A2(n5740), .ZN(n9478) );
  OR2_X1 U6088 ( .A1(P1_U3083), .A2(n6160), .ZN(n9643) );
  OR2_X1 U6089 ( .A1(n9676), .A2(n9472), .ZN(n9268) );
  INV_X1 U6090 ( .A(n9666), .ZN(n9274) );
  OR2_X1 U6091 ( .A1(n9676), .A2(n9466), .ZN(n9279) );
  AND2_X1 U6092 ( .A1(n6509), .A2(n9663), .ZN(n9676) );
  INV_X1 U6093 ( .A(n9722), .ZN(n9720) );
  INV_X1 U6094 ( .A(n9679), .ZN(n9680) );
  INV_X1 U6095 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n9944) );
  NAND2_X1 U6096 ( .A1(n5966), .A2(n4694), .ZN(P1_U3551) );
  NOR2_X1 U6097 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n4710) );
  NOR2_X1 U6098 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_9__SCAN_IN), .ZN(
        n4709) );
  INV_X1 U6099 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5082) );
  NOR2_X1 U6100 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n4714) );
  INV_X1 U6101 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n4739) );
  INV_X1 U6102 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n4741) );
  INV_X1 U6103 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5429) );
  NAND4_X1 U6104 ( .A1(n4714), .A2(n4739), .A3(n4741), .A4(n5429), .ZN(n4718)
         );
  INV_X1 U6105 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n4716) );
  INV_X1 U6106 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n4735) );
  INV_X1 U6107 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n4715) );
  NAND4_X1 U6108 ( .A1(n4734), .A2(n4716), .A3(n4735), .A4(n4715), .ZN(n4717)
         );
  NOR2_X1 U6109 ( .A1(n4718), .A2(n4717), .ZN(n5418) );
  INV_X1 U6110 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n4719) );
  AND2_X1 U6111 ( .A1(n4719), .A2(n5420), .ZN(n4720) );
  NOR2_X2 U6112 ( .A1(n5424), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4745) );
  INV_X1 U6113 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4746) );
  INV_X1 U6114 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n4722) );
  INV_X1 U6115 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6328) );
  OR2_X1 U6116 ( .A1(n4769), .A2(n6328), .ZN(n4733) );
  INV_X1 U6117 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n4727) );
  OR2_X1 U6118 ( .A1(n4940), .A2(n4727), .ZN(n4732) );
  NAND2_X4 U6119 ( .A1(n4729), .A2(n4726), .ZN(n4838) );
  INV_X1 U6120 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6573) );
  OR2_X1 U6121 ( .A1(n4838), .A2(n6573), .ZN(n4731) );
  NAND2_X1 U6122 ( .A1(n4814), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n4730) );
  AND4_X2 U6123 ( .A1(n4733), .A2(n4732), .A3(n4731), .A4(n4730), .ZN(n7969)
         );
  NAND2_X1 U6124 ( .A1(n5110), .A2(n4734), .ZN(n5156) );
  NAND2_X1 U6125 ( .A1(n4738), .A2(n4739), .ZN(n4736) );
  XNOR2_X1 U6126 ( .A(n5430), .B(n5429), .ZN(n5462) );
  INV_X1 U6127 ( .A(n8269), .ZN(n9772) );
  NAND2_X1 U6128 ( .A1(n4744), .A2(n4741), .ZN(n4742) );
  NAND2_X1 U6129 ( .A1(n4742), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4743) );
  OR2_X4 U6130 ( .A1(n9861), .A2(n8511), .ZN(n8121) );
  NOR2_X1 U6131 ( .A1(n7969), .A2(n5409), .ZN(n4765) );
  NAND2_X1 U6132 ( .A1(n5424), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4749) );
  INV_X1 U6133 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n4748) );
  OR2_X1 U6134 ( .A1(n4750), .A2(n4737), .ZN(n4751) );
  XNOR2_X1 U6135 ( .A(n4751), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9381) );
  INV_X1 U6136 ( .A(n9381), .ZN(n6010) );
  INV_X1 U6137 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4753) );
  INV_X1 U6138 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4752) );
  AND2_X1 U6139 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n4756) );
  NAND2_X1 U6140 ( .A1(n4781), .A2(n4756), .ZN(n5529) );
  INV_X1 U6141 ( .A(SI_1_), .ZN(n4757) );
  XNOR2_X1 U6142 ( .A(n4758), .B(n4757), .ZN(n4797) );
  MUX2_X1 U6143 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4781), .Z(n4796) );
  NAND2_X1 U6144 ( .A1(n4797), .A2(n4796), .ZN(n4760) );
  NAND2_X1 U6145 ( .A1(n4758), .A2(SI_1_), .ZN(n4759) );
  NAND2_X1 U6146 ( .A1(n4760), .A2(n4759), .ZN(n4776) );
  INV_X1 U6147 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6017) );
  INV_X1 U6148 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6009) );
  MUX2_X1 U6149 ( .A(n6017), .B(n6009), .S(n4761), .Z(n4777) );
  XNOR2_X1 U6150 ( .A(n4777), .B(SI_2_), .ZN(n4775) );
  XNOR2_X1 U6151 ( .A(n4776), .B(n4775), .ZN(n6016) );
  OR2_X1 U6152 ( .A1(n4952), .A2(n6016), .ZN(n4763) );
  INV_X8 U6153 ( .A(n4761), .ZN(n7393) );
  NAND2_X4 U6154 ( .A1(n4762), .A2(n7393), .ZN(n8110) );
  XNOR2_X1 U6155 ( .A(n9786), .B(n5410), .ZN(n4766) );
  NAND2_X1 U6156 ( .A1(n4765), .A2(n4766), .ZN(n4812) );
  INV_X1 U6157 ( .A(n4765), .ZN(n4767) );
  INV_X1 U6158 ( .A(n4766), .ZN(n7968) );
  NAND2_X1 U6159 ( .A1(n4767), .A2(n7968), .ZN(n4768) );
  INV_X1 U6160 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6325) );
  OR2_X1 U6161 ( .A1(n4260), .A2(n6325), .ZN(n4773) );
  OR2_X1 U6162 ( .A1(n4838), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n4772) );
  NAND2_X1 U6163 ( .A1(n4814), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4771) );
  NAND2_X1 U6164 ( .A1(n4259), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n4770) );
  AND2_X1 U6165 ( .A1(n8326), .A2(n4254), .ZN(n4785) );
  NAND2_X1 U6166 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4696), .ZN(n4774) );
  XNOR2_X1 U6167 ( .A(n4774), .B(P2_IR_REG_3__SCAN_IN), .ZN(n6340) );
  INV_X1 U6168 ( .A(n6340), .ZN(n8338) );
  NAND2_X1 U6169 ( .A1(n4776), .A2(n4775), .ZN(n4780) );
  INV_X1 U6170 ( .A(n4777), .ZN(n4778) );
  NAND2_X1 U6171 ( .A1(n4778), .A2(SI_2_), .ZN(n4779) );
  NAND2_X1 U6172 ( .A1(n4780), .A2(n4779), .ZN(n4824) );
  INV_X1 U6173 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6012) );
  INV_X1 U6174 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6015) );
  MUX2_X1 U6175 ( .A(n6012), .B(n6015), .S(n4781), .Z(n4825) );
  XNOR2_X1 U6176 ( .A(n4825), .B(SI_3_), .ZN(n4823) );
  XNOR2_X1 U6177 ( .A(n4824), .B(n4823), .ZN(n6014) );
  OR2_X1 U6178 ( .A1(n4952), .A2(n6014), .ZN(n4783) );
  OR2_X1 U6179 ( .A1(n8110), .A2(n6012), .ZN(n4782) );
  NAND2_X1 U6180 ( .A1(n4785), .A2(n4784), .ZN(n4832) );
  INV_X1 U6181 ( .A(n4784), .ZN(n8039) );
  INV_X1 U6182 ( .A(n4785), .ZN(n4786) );
  NAND2_X1 U6183 ( .A1(n8039), .A2(n4786), .ZN(n4787) );
  AND2_X1 U6184 ( .A1(n4832), .A2(n4787), .ZN(n4811) );
  AND2_X1 U6185 ( .A1(n6568), .A2(n4811), .ZN(n4813) );
  NAND2_X1 U6186 ( .A1(n4802), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n4791) );
  INV_X1 U6187 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n9734) );
  OR2_X1 U6188 ( .A1(n4838), .A2(n9734), .ZN(n4790) );
  NAND2_X1 U6189 ( .A1(n4814), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n4789) );
  NAND2_X1 U6190 ( .A1(n4816), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n4788) );
  NAND2_X1 U6191 ( .A1(n4761), .A2(SI_0_), .ZN(n4793) );
  INV_X1 U6192 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n4792) );
  XNOR2_X1 U6193 ( .A(n4793), .B(n4792), .ZN(n8854) );
  INV_X1 U6194 ( .A(n9773), .ZN(n9754) );
  NAND2_X1 U6195 ( .A1(n6702), .A2(n9754), .ZN(n9751) );
  INV_X1 U6196 ( .A(n9751), .ZN(n4794) );
  NAND2_X1 U6197 ( .A1(n4794), .A2(n8121), .ZN(n6594) );
  NAND2_X1 U6198 ( .A1(n5302), .A2(n9773), .ZN(n4795) );
  NAND2_X1 U6199 ( .A1(n6594), .A2(n4795), .ZN(n6576) );
  XNOR2_X1 U6200 ( .A(n4797), .B(n4796), .ZN(n6020) );
  OR2_X1 U6201 ( .A1(n4952), .A2(n6020), .ZN(n4800) );
  INV_X1 U6202 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6011) );
  INV_X1 U6203 ( .A(n4750), .ZN(n4798) );
  OR2_X1 U6204 ( .A1(n5997), .A2(n6335), .ZN(n4799) );
  XNOR2_X1 U6205 ( .A(n9778), .B(n5410), .ZN(n4809) );
  INV_X1 U6206 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n4801) );
  OR2_X1 U6207 ( .A1(n4838), .A2(n4801), .ZN(n4804) );
  NAND2_X1 U6208 ( .A1(n4802), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n4803) );
  AND2_X1 U6209 ( .A1(n4804), .A2(n4803), .ZN(n4807) );
  NAND2_X1 U6210 ( .A1(n4816), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n4806) );
  NAND2_X1 U6211 ( .A1(n6691), .A2(n4253), .ZN(n4808) );
  XNOR2_X1 U6212 ( .A(n4809), .B(n4808), .ZN(n6575) );
  NAND2_X1 U6213 ( .A1(n4809), .A2(n4808), .ZN(n4810) );
  INV_X1 U6214 ( .A(n4811), .ZN(n7970) );
  NAND2_X1 U6215 ( .A1(n4814), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n4818) );
  INV_X1 U6216 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n4815) );
  INV_X1 U6217 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6347) );
  XNOR2_X1 U6218 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n8047) );
  OR2_X1 U6219 ( .A1(n4838), .A2(n8047), .ZN(n4817) );
  NAND2_X1 U6220 ( .A1(n4400), .A2(n8121), .ZN(n4836) );
  NAND2_X1 U6221 ( .A1(n4819), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4820) );
  MUX2_X1 U6222 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4820), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n4822) );
  NAND2_X1 U6223 ( .A1(n4822), .A2(n4821), .ZN(n6359) );
  NAND2_X1 U6224 ( .A1(n4824), .A2(n4823), .ZN(n4828) );
  INV_X1 U6225 ( .A(n4825), .ZN(n4826) );
  NAND2_X1 U6226 ( .A1(n4826), .A2(SI_3_), .ZN(n4827) );
  NAND2_X1 U6227 ( .A1(n4828), .A2(n4827), .ZN(n4847) );
  INV_X1 U6228 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6013) );
  INV_X1 U6229 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6019) );
  XNOR2_X1 U6230 ( .A(n4847), .B(n4846), .ZN(n6018) );
  OR2_X1 U6231 ( .A1(n4952), .A2(n6018), .ZN(n4831) );
  OR2_X1 U6232 ( .A1(n8110), .A2(n6013), .ZN(n4830) );
  XNOR2_X1 U6233 ( .A(n8042), .B(n5410), .ZN(n4834) );
  XNOR2_X1 U6234 ( .A(n4836), .B(n4834), .ZN(n8045) );
  AND2_X1 U6235 ( .A1(n8045), .A2(n4832), .ZN(n4833) );
  INV_X1 U6236 ( .A(n4834), .ZN(n4835) );
  NAND2_X1 U6237 ( .A1(n4836), .A2(n4835), .ZN(n4837) );
  NAND2_X1 U6238 ( .A1(n8043), .A2(n4837), .ZN(n6796) );
  INV_X1 U6239 ( .A(n6796), .ZN(n4861) );
  NAND2_X1 U6240 ( .A1(n4259), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n4845) );
  INV_X1 U6241 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6344) );
  OR2_X1 U6242 ( .A1(n4260), .A2(n6344), .ZN(n4844) );
  NAND3_X1 U6243 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .A3(P2_REG3_REG_5__SCAN_IN), .ZN(n4863) );
  INV_X1 U6244 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n4840) );
  NAND2_X1 U6245 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n4839) );
  NAND2_X1 U6246 ( .A1(n4840), .A2(n4839), .ZN(n4841) );
  NAND2_X1 U6247 ( .A1(n4863), .A2(n4841), .ZN(n6937) );
  OR2_X1 U6248 ( .A1(n4838), .A2(n6937), .ZN(n4843) );
  NAND2_X1 U6249 ( .A1(n4814), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n4842) );
  NAND4_X1 U6250 ( .A1(n4845), .A2(n4844), .A3(n4843), .A4(n4842), .ZN(n8325)
         );
  AND2_X1 U6251 ( .A1(n8325), .A2(n8121), .ZN(n4856) );
  NAND2_X1 U6252 ( .A1(n4847), .A2(n4846), .ZN(n4851) );
  INV_X1 U6253 ( .A(n4848), .ZN(n4849) );
  NAND2_X1 U6254 ( .A1(n4849), .A2(SI_4_), .ZN(n4850) );
  NAND2_X1 U6255 ( .A1(n4851), .A2(n4850), .ZN(n4872) );
  INV_X1 U6256 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6022) );
  MUX2_X1 U6257 ( .A(n6022), .B(n9944), .S(n7393), .Z(n4873) );
  XNOR2_X1 U6258 ( .A(n4872), .B(n4871), .ZN(n6023) );
  OR2_X1 U6259 ( .A1(n4952), .A2(n6023), .ZN(n4855) );
  OR2_X1 U6260 ( .A1(n8110), .A2(n6022), .ZN(n4854) );
  NAND2_X1 U6261 ( .A1(n4821), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4852) );
  XNOR2_X1 U6262 ( .A(n4852), .B(P2_IR_REG_5__SCAN_IN), .ZN(n6363) );
  INV_X1 U6263 ( .A(n6363), .ZN(n8350) );
  OR2_X1 U6264 ( .A1(n5997), .A2(n8350), .ZN(n4853) );
  XNOR2_X1 U6265 ( .A(n9810), .B(n5302), .ZN(n8075) );
  NAND2_X1 U6266 ( .A1(n4856), .A2(n8075), .ZN(n4878) );
  INV_X1 U6267 ( .A(n8075), .ZN(n4858) );
  INV_X1 U6268 ( .A(n4856), .ZN(n4857) );
  NAND2_X1 U6269 ( .A1(n4858), .A2(n4857), .ZN(n4859) );
  NAND2_X1 U6270 ( .A1(n4878), .A2(n4859), .ZN(n6795) );
  NAND2_X1 U6271 ( .A1(n4259), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n4868) );
  INV_X1 U6272 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6350) );
  OR2_X1 U6273 ( .A1(n4260), .A2(n6350), .ZN(n4867) );
  INV_X1 U6274 ( .A(n4863), .ZN(n4862) );
  NAND2_X1 U6275 ( .A1(n4862), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n4886) );
  INV_X1 U6276 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n6395) );
  NAND2_X1 U6277 ( .A1(n4863), .A2(n6395), .ZN(n4864) );
  NAND2_X1 U6278 ( .A1(n4886), .A2(n4864), .ZN(n6765) );
  OR2_X1 U6279 ( .A1(n4838), .A2(n6765), .ZN(n4866) );
  INV_X1 U6280 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n6364) );
  OR2_X1 U6281 ( .A1(n7897), .A2(n6364), .ZN(n4865) );
  INV_X1 U6282 ( .A(n7091), .ZN(n8324) );
  NAND2_X1 U6283 ( .A1(n8324), .A2(n8121), .ZN(n4882) );
  OR2_X1 U6284 ( .A1(n4869), .A2(n4737), .ZN(n4870) );
  XNOR2_X1 U6285 ( .A(n4870), .B(n4896), .ZN(n6404) );
  INV_X1 U6286 ( .A(n4873), .ZN(n4874) );
  NAND2_X1 U6287 ( .A1(n4874), .A2(SI_5_), .ZN(n4875) );
  INV_X1 U6288 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6024) );
  INV_X1 U6289 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6026) );
  MUX2_X1 U6290 ( .A(n6024), .B(n6026), .S(n7393), .Z(n4894) );
  XNOR2_X1 U6291 ( .A(n4893), .B(n4892), .ZN(n6025) );
  OR2_X1 U6292 ( .A1(n4952), .A2(n6025), .ZN(n4877) );
  OR2_X1 U6293 ( .A1(n8110), .A2(n6024), .ZN(n4876) );
  OAI211_X1 U6294 ( .C1(n5997), .C2(n6404), .A(n4877), .B(n4876), .ZN(n8080)
         );
  XNOR2_X1 U6295 ( .A(n8080), .B(n5410), .ZN(n4880) );
  XNOR2_X1 U6296 ( .A(n4882), .B(n4880), .ZN(n8084) );
  AND2_X1 U6297 ( .A1(n8084), .A2(n4878), .ZN(n4879) );
  INV_X1 U6298 ( .A(n4880), .ZN(n4881) );
  NAND2_X1 U6299 ( .A1(n4882), .A2(n4881), .ZN(n4883) );
  NAND2_X1 U6300 ( .A1(n4259), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n4891) );
  INV_X1 U6301 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6343) );
  OR2_X1 U6302 ( .A1(n4260), .A2(n6343), .ZN(n4890) );
  INV_X1 U6303 ( .A(n4886), .ZN(n4884) );
  NAND2_X1 U6304 ( .A1(n4884), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n4909) );
  INV_X1 U6305 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n4885) );
  NAND2_X1 U6306 ( .A1(n4886), .A2(n4885), .ZN(n4887) );
  NAND2_X1 U6307 ( .A1(n4909), .A2(n4887), .ZN(n6818) );
  OR2_X1 U6308 ( .A1(n4838), .A2(n6818), .ZN(n4889) );
  NAND2_X1 U6309 ( .A1(n4814), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n4888) );
  NAND4_X1 U6310 ( .A1(n4891), .A2(n4890), .A3(n4889), .A4(n4888), .ZN(n8323)
         );
  AND2_X1 U6311 ( .A1(n8323), .A2(n4253), .ZN(n4902) );
  INV_X1 U6312 ( .A(n4894), .ZN(n4895) );
  INV_X1 U6313 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6027) );
  INV_X1 U6314 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6029) );
  MUX2_X1 U6315 ( .A(n6027), .B(n6029), .S(n7393), .Z(n4921) );
  XNOR2_X1 U6316 ( .A(n4920), .B(n4919), .ZN(n6028) );
  OR2_X1 U6317 ( .A1(n4952), .A2(n6028), .ZN(n4900) );
  OR2_X1 U6318 ( .A1(n8110), .A2(n6027), .ZN(n4899) );
  NAND2_X1 U6319 ( .A1(n4869), .A2(n4896), .ZN(n4915) );
  NAND2_X1 U6320 ( .A1(n4915), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4897) );
  XNOR2_X1 U6321 ( .A(n4897), .B(P2_IR_REG_7__SCAN_IN), .ZN(n8357) );
  INV_X1 U6322 ( .A(n8357), .ZN(n6370) );
  OR2_X1 U6323 ( .A1(n5997), .A2(n6370), .ZN(n4898) );
  XNOR2_X1 U6324 ( .A(n9823), .B(n5302), .ZN(n4901) );
  NAND2_X1 U6325 ( .A1(n4902), .A2(n4901), .ZN(n4906) );
  INV_X1 U6326 ( .A(n4901), .ZN(n6829) );
  INV_X1 U6327 ( .A(n4902), .ZN(n4903) );
  NAND2_X1 U6328 ( .A1(n6829), .A2(n4903), .ZN(n4904) );
  NAND2_X1 U6329 ( .A1(n4906), .A2(n4904), .ZN(n6816) );
  NAND2_X1 U6330 ( .A1(n6828), .A2(n4906), .ZN(n4931) );
  NAND2_X1 U6331 ( .A1(n4259), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n4914) );
  INV_X1 U6332 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6352) );
  OR2_X1 U6333 ( .A1(n4260), .A2(n6352), .ZN(n4913) );
  INV_X1 U6334 ( .A(n4909), .ZN(n4907) );
  NAND2_X1 U6335 ( .A1(n4907), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n4938) );
  INV_X1 U6336 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n4908) );
  NAND2_X1 U6337 ( .A1(n4909), .A2(n4908), .ZN(n4910) );
  NAND2_X1 U6338 ( .A1(n4938), .A2(n4910), .ZN(n7022) );
  OR2_X1 U6339 ( .A1(n4838), .A2(n7022), .ZN(n4912) );
  INV_X1 U6340 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6390) );
  OR2_X1 U6341 ( .A1(n7897), .A2(n6390), .ZN(n4911) );
  NAND2_X1 U6342 ( .A1(n8322), .A2(n8121), .ZN(n4932) );
  NAND2_X1 U6343 ( .A1(n4917), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4916) );
  MUX2_X1 U6344 ( .A(P2_IR_REG_31__SCAN_IN), .B(n4916), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n4918) );
  NAND2_X1 U6345 ( .A1(n4918), .A2(n4965), .ZN(n6389) );
  NAND2_X1 U6346 ( .A1(n4920), .A2(n4919), .ZN(n4924) );
  INV_X1 U6347 ( .A(n4921), .ZN(n4922) );
  NAND2_X1 U6348 ( .A1(n4922), .A2(SI_7_), .ZN(n4923) );
  INV_X1 U6349 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6032) );
  INV_X1 U6350 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6034) );
  MUX2_X1 U6351 ( .A(n6032), .B(n6034), .S(n7393), .Z(n4926) );
  INV_X1 U6352 ( .A(SI_8_), .ZN(n4925) );
  INV_X1 U6353 ( .A(n4926), .ZN(n4927) );
  NAND2_X1 U6354 ( .A1(n4927), .A2(SI_8_), .ZN(n4928) );
  XNOR2_X1 U6355 ( .A(n4947), .B(n4250), .ZN(n6033) );
  OR2_X1 U6356 ( .A1(n6033), .A2(n4952), .ZN(n4930) );
  OR2_X1 U6357 ( .A1(n8110), .A2(n6032), .ZN(n4929) );
  OAI211_X1 U6358 ( .C1(n5997), .C2(n6389), .A(n4930), .B(n4929), .ZN(n7024)
         );
  XNOR2_X1 U6359 ( .A(n7024), .B(n5410), .ZN(n4933) );
  XNOR2_X1 U6360 ( .A(n4932), .B(n4933), .ZN(n6826) );
  NAND2_X1 U6361 ( .A1(n4931), .A2(n6826), .ZN(n6830) );
  INV_X1 U6362 ( .A(n4932), .ZN(n4934) );
  NAND2_X1 U6363 ( .A1(n4934), .A2(n4933), .ZN(n4935) );
  NAND2_X1 U6364 ( .A1(n4816), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n4945) );
  INV_X1 U6365 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6964) );
  OR2_X1 U6366 ( .A1(n7897), .A2(n6964), .ZN(n4944) );
  INV_X1 U6367 ( .A(n4938), .ZN(n4936) );
  NAND2_X1 U6368 ( .A1(n4936), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n4972) );
  INV_X1 U6369 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n4937) );
  NAND2_X1 U6370 ( .A1(n4938), .A2(n4937), .ZN(n4939) );
  NAND2_X1 U6371 ( .A1(n4972), .A2(n4939), .ZN(n6963) );
  OR2_X1 U6372 ( .A1(n4838), .A2(n6963), .ZN(n4943) );
  INV_X1 U6373 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n4941) );
  OR2_X1 U6374 ( .A1(n7899), .A2(n4941), .ZN(n4942) );
  NOR2_X1 U6375 ( .A1(n7073), .A2(n5409), .ZN(n4956) );
  INV_X1 U6376 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6037) );
  INV_X1 U6377 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6036) );
  MUX2_X1 U6378 ( .A(n6037), .B(n6036), .S(n7393), .Z(n4949) );
  INV_X1 U6379 ( .A(SI_9_), .ZN(n4948) );
  INV_X1 U6380 ( .A(n4949), .ZN(n4950) );
  NAND2_X1 U6381 ( .A1(n4950), .A2(SI_9_), .ZN(n4951) );
  XNOR2_X1 U6382 ( .A(n4959), .B(n4701), .ZN(n6035) );
  NAND2_X1 U6383 ( .A1(n6035), .A2(n8108), .ZN(n4955) );
  NAND2_X1 U6384 ( .A1(n4965), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4953) );
  XNOR2_X1 U6385 ( .A(n4953), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6406) );
  AOI22_X1 U6386 ( .A1(n5184), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5183), .B2(
        n6406), .ZN(n4954) );
  NAND2_X1 U6387 ( .A1(n4955), .A2(n4954), .ZN(n6968) );
  XNOR2_X1 U6388 ( .A(n6968), .B(n5410), .ZN(n4957) );
  AND2_X1 U6389 ( .A1(n4956), .A2(n4957), .ZN(n5971) );
  INV_X1 U6390 ( .A(n4956), .ZN(n4958) );
  INV_X1 U6391 ( .A(n4957), .ZN(n5973) );
  NAND2_X1 U6392 ( .A1(n4958), .A2(n5973), .ZN(n5975) );
  INV_X1 U6393 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6040) );
  INV_X1 U6394 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6043) );
  MUX2_X1 U6395 ( .A(n6040), .B(n6043), .S(n7393), .Z(n4962) );
  INV_X1 U6396 ( .A(SI_10_), .ZN(n4961) );
  NAND2_X1 U6397 ( .A1(n4962), .A2(n4961), .ZN(n4985) );
  INV_X1 U6398 ( .A(n4962), .ZN(n4963) );
  NAND2_X1 U6399 ( .A1(n4963), .A2(SI_10_), .ZN(n4964) );
  XNOR2_X1 U6400 ( .A(n4984), .B(n4698), .ZN(n6039) );
  NAND2_X1 U6401 ( .A1(n6039), .A2(n8108), .ZN(n4970) );
  OAI21_X1 U6402 ( .B1(n4965), .B2(P2_IR_REG_9__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n4967) );
  INV_X1 U6403 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n4966) );
  OR2_X1 U6404 ( .A1(n4967), .A2(n4966), .ZN(n4968) );
  NAND2_X1 U6405 ( .A1(n4967), .A2(n4966), .ZN(n4987) );
  AOI22_X1 U6406 ( .A1(n5184), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5183), .B2(
        n6549), .ZN(n4969) );
  XNOR2_X1 U6407 ( .A(n9844), .B(n5302), .ZN(n4979) );
  NAND2_X1 U6408 ( .A1(n4816), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n4978) );
  INV_X1 U6409 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n4971) );
  OR2_X1 U6410 ( .A1(n7899), .A2(n4971), .ZN(n4977) );
  INV_X1 U6411 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U6412 ( .A1(n4972), .A2(n6405), .ZN(n4973) );
  NAND2_X1 U6413 ( .A1(n4993), .A2(n4973), .ZN(n7043) );
  OR2_X1 U6414 ( .A1(n4838), .A2(n7043), .ZN(n4976) );
  INV_X1 U6415 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n4974) );
  OR2_X1 U6416 ( .A1(n7897), .A2(n4974), .ZN(n4975) );
  INV_X1 U6417 ( .A(n7062), .ZN(n8320) );
  NAND2_X1 U6418 ( .A1(n8320), .A2(n8121), .ZN(n4980) );
  XNOR2_X1 U6419 ( .A(n4979), .B(n4980), .ZN(n7041) );
  INV_X1 U6420 ( .A(n4979), .ZN(n4982) );
  INV_X1 U6421 ( .A(n4980), .ZN(n4981) );
  NAND2_X1 U6422 ( .A1(n4982), .A2(n4981), .ZN(n4983) );
  NAND2_X1 U6423 ( .A1(n4984), .A2(n4698), .ZN(n4986) );
  MUX2_X1 U6424 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n7393), .Z(n5000) );
  INV_X1 U6425 ( .A(SI_11_), .ZN(n10044) );
  NAND2_X1 U6426 ( .A1(n5657), .A2(n8108), .ZN(n4990) );
  NAND2_X1 U6427 ( .A1(n4987), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4988) );
  XNOR2_X1 U6428 ( .A(n4988), .B(P2_IR_REG_11__SCAN_IN), .ZN(n8370) );
  AOI22_X1 U6429 ( .A1(n5184), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5183), .B2(
        n8370), .ZN(n4989) );
  NAND2_X1 U6430 ( .A1(n4990), .A2(n4989), .ZN(n7251) );
  XNOR2_X1 U6431 ( .A(n7251), .B(n5410), .ZN(n5138) );
  NAND2_X1 U6432 ( .A1(n4816), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n4998) );
  INV_X1 U6433 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n4991) );
  OR2_X1 U6434 ( .A1(n7899), .A2(n4991), .ZN(n4997) );
  INV_X1 U6435 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U6436 ( .A1(n4993), .A2(n4992), .ZN(n4994) );
  NAND2_X1 U6437 ( .A1(n5034), .A2(n4994), .ZN(n7250) );
  OR2_X1 U6438 ( .A1(n4838), .A2(n7250), .ZN(n4996) );
  INV_X1 U6439 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7165) );
  OR2_X1 U6440 ( .A1(n7897), .A2(n7165), .ZN(n4995) );
  INV_X1 U6441 ( .A(n7328), .ZN(n8319) );
  NAND2_X1 U6442 ( .A1(n8319), .A2(n8121), .ZN(n5136) );
  XNOR2_X1 U6443 ( .A(n5138), .B(n5136), .ZN(n7322) );
  NAND2_X1 U6444 ( .A1(n5000), .A2(SI_11_), .ZN(n5001) );
  INV_X1 U6445 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6103) );
  INV_X1 U6446 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5004) );
  MUX2_X1 U6447 ( .A(n6103), .B(n5004), .S(n7393), .Z(n5005) );
  INV_X1 U6448 ( .A(SI_12_), .ZN(n9942) );
  INV_X1 U6449 ( .A(n5005), .ZN(n5006) );
  NAND2_X1 U6450 ( .A1(n5006), .A2(SI_12_), .ZN(n5007) );
  NAND2_X1 U6451 ( .A1(n5008), .A2(n5007), .ZN(n5028) );
  INV_X1 U6452 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6137) );
  INV_X1 U6453 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6129) );
  MUX2_X1 U6454 ( .A(n6137), .B(n6129), .S(n7393), .Z(n5010) );
  INV_X1 U6455 ( .A(SI_13_), .ZN(n5009) );
  NAND2_X1 U6456 ( .A1(n5010), .A2(n5009), .ZN(n5042) );
  INV_X1 U6457 ( .A(n5010), .ZN(n5011) );
  NAND2_X1 U6458 ( .A1(n5011), .A2(SI_13_), .ZN(n5012) );
  NAND2_X1 U6459 ( .A1(n6128), .A2(n8108), .ZN(n5017) );
  NAND2_X1 U6460 ( .A1(n5013), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5014) );
  MUX2_X1 U6461 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5014), .S(
        P2_IR_REG_13__SCAN_IN), .Z(n5015) );
  AND2_X1 U6462 ( .A1(n5015), .A2(n4315), .ZN(n6665) );
  AOI22_X1 U6463 ( .A1(n5184), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5183), .B2(
        n6665), .ZN(n5016) );
  NAND2_X2 U6464 ( .A1(n5017), .A2(n5016), .ZN(n7919) );
  XNOR2_X1 U6465 ( .A(n7919), .B(n5410), .ZN(n5024) );
  NAND2_X1 U6466 ( .A1(n4259), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5023) );
  INV_X1 U6467 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5018) );
  OR2_X1 U6468 ( .A1(n4260), .A2(n5018), .ZN(n5022) );
  INV_X1 U6469 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5047) );
  XNOR2_X1 U6470 ( .A(n5049), .B(n5047), .ZN(n7307) );
  OR2_X1 U6471 ( .A1(n4838), .A2(n7307), .ZN(n5021) );
  INV_X1 U6472 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7308) );
  OR2_X1 U6473 ( .A1(n7897), .A2(n7308), .ZN(n5020) );
  NOR2_X1 U6474 ( .A1(n7365), .A2(n5409), .ZN(n5025) );
  NAND2_X1 U6475 ( .A1(n5024), .A2(n5025), .ZN(n5134) );
  INV_X1 U6476 ( .A(n5024), .ZN(n7364) );
  INV_X1 U6477 ( .A(n5025), .ZN(n5026) );
  NAND2_X1 U6478 ( .A1(n7364), .A2(n5026), .ZN(n5027) );
  XNOR2_X1 U6479 ( .A(n5029), .B(n5028), .ZN(n6083) );
  NAND2_X1 U6480 ( .A1(n6083), .A2(n8108), .ZN(n5033) );
  OR2_X1 U6481 ( .A1(n5030), .A2(n4737), .ZN(n5031) );
  XNOR2_X1 U6482 ( .A(n5031), .B(P2_IR_REG_12__SCAN_IN), .ZN(n6551) );
  AOI22_X1 U6483 ( .A1(n5184), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5183), .B2(
        n6551), .ZN(n5032) );
  XNOR2_X1 U6484 ( .A(n7170), .B(n5302), .ZN(n5139) );
  NAND2_X1 U6485 ( .A1(n4259), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5039) );
  INV_X1 U6486 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6544) );
  OR2_X1 U6487 ( .A1(n4260), .A2(n6544), .ZN(n5038) );
  INV_X1 U6488 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n8385) );
  NAND2_X1 U6489 ( .A1(n5034), .A2(n8385), .ZN(n5035) );
  NAND2_X1 U6490 ( .A1(n5049), .A2(n5035), .ZN(n7327) );
  OR2_X1 U6491 ( .A1(n4838), .A2(n7327), .ZN(n5037) );
  INV_X1 U6492 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7183) );
  OR2_X1 U6493 ( .A1(n7897), .A2(n7183), .ZN(n5036) );
  INV_X1 U6494 ( .A(n7306), .ZN(n8318) );
  NAND2_X1 U6495 ( .A1(n8318), .A2(n8121), .ZN(n5140) );
  NAND2_X1 U6496 ( .A1(n5139), .A2(n5140), .ZN(n7320) );
  AND2_X1 U6497 ( .A1(n7322), .A2(n5135), .ZN(n7292) );
  INV_X1 U6498 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6163) );
  INV_X1 U6499 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n5043) );
  MUX2_X1 U6500 ( .A(n6163), .B(n5043), .S(n7393), .Z(n5058) );
  XNOR2_X1 U6501 ( .A(n5058), .B(SI_14_), .ZN(n5057) );
  NAND2_X1 U6502 ( .A1(n6135), .A2(n8108), .ZN(n5045) );
  NAND2_X1 U6503 ( .A1(n4315), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5083) );
  XNOR2_X1 U6504 ( .A(n5083), .B(P2_IR_REG_14__SCAN_IN), .ZN(n6997) );
  AOI22_X1 U6505 ( .A1(n5184), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5183), .B2(
        n6997), .ZN(n5044) );
  XNOR2_X1 U6506 ( .A(n7871), .B(n5410), .ZN(n5133) );
  INV_X1 U6507 ( .A(n5133), .ZN(n5055) );
  NAND2_X1 U6508 ( .A1(n4259), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5054) );
  INV_X1 U6509 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5046) );
  OR2_X1 U6510 ( .A1(n4260), .A2(n5046), .ZN(n5053) );
  INV_X1 U6511 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5048) );
  OAI21_X1 U6512 ( .B1(n5049), .B2(n5047), .A(n5048), .ZN(n5050) );
  NAND2_X1 U6513 ( .A1(n5050), .A2(n5089), .ZN(n8740) );
  OR2_X1 U6514 ( .A1(n4838), .A2(n8740), .ZN(n5052) );
  INV_X1 U6515 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8741) );
  OR2_X1 U6516 ( .A1(n7897), .A2(n8741), .ZN(n5051) );
  NAND2_X1 U6517 ( .A1(n4663), .A2(n8121), .ZN(n5132) );
  NAND2_X1 U6518 ( .A1(n5055), .A2(n5132), .ZN(n5131) );
  AND2_X1 U6519 ( .A1(n7292), .A2(n5131), .ZN(n7715) );
  INV_X1 U6520 ( .A(n5056), .ZN(n5060) );
  INV_X1 U6521 ( .A(n5058), .ZN(n5059) );
  INV_X1 U6522 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6263) );
  INV_X1 U6523 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6261) );
  MUX2_X1 U6524 ( .A(n6263), .B(n6261), .S(n7393), .Z(n5062) );
  INV_X1 U6525 ( .A(SI_15_), .ZN(n5061) );
  NAND2_X1 U6526 ( .A1(n5062), .A2(n5061), .ZN(n5066) );
  INV_X1 U6527 ( .A(n5062), .ZN(n5063) );
  NAND2_X1 U6528 ( .A1(n5063), .A2(SI_15_), .ZN(n5064) );
  NAND2_X1 U6529 ( .A1(n5066), .A2(n5064), .ZN(n5078) );
  NAND2_X1 U6530 ( .A1(n5077), .A2(n5065), .ZN(n5080) );
  NAND2_X1 U6531 ( .A1(n5080), .A2(n5066), .ZN(n5106) );
  INV_X1 U6532 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n5068) );
  INV_X1 U6533 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5067) );
  MUX2_X1 U6534 ( .A(n5068), .B(n5067), .S(n7393), .Z(n5070) );
  INV_X1 U6535 ( .A(SI_16_), .ZN(n5069) );
  NAND2_X1 U6536 ( .A1(n5070), .A2(n5069), .ZN(n5107) );
  INV_X1 U6537 ( .A(n5070), .ZN(n5071) );
  NAND2_X1 U6538 ( .A1(n5071), .A2(SI_16_), .ZN(n5072) );
  XNOR2_X1 U6539 ( .A(n5106), .B(n5105), .ZN(n6264) );
  NAND2_X1 U6540 ( .A1(n6264), .A2(n8108), .ZN(n5076) );
  NAND2_X1 U6541 ( .A1(n5073), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5074) );
  XNOR2_X1 U6542 ( .A(n5074), .B(P2_IR_REG_16__SCAN_IN), .ZN(n8418) );
  AOI22_X1 U6543 ( .A1(n5184), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5183), .B2(
        n8418), .ZN(n5075) );
  XNOR2_X1 U6544 ( .A(n8693), .B(n5410), .ZN(n8007) );
  INV_X1 U6545 ( .A(n8007), .ZN(n5104) );
  INV_X1 U6546 ( .A(n5077), .ZN(n5079) );
  NAND2_X1 U6547 ( .A1(n5079), .A2(n5078), .ZN(n5081) );
  NAND2_X1 U6548 ( .A1(n5081), .A2(n5080), .ZN(n6260) );
  NAND2_X1 U6549 ( .A1(n6260), .A2(n8108), .ZN(n5087) );
  NAND2_X1 U6550 ( .A1(n5083), .A2(n5082), .ZN(n5084) );
  NAND2_X1 U6551 ( .A1(n5084), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5085) );
  XNOR2_X1 U6552 ( .A(n5085), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8406) );
  AOI22_X1 U6553 ( .A1(n5184), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5183), .B2(
        n8406), .ZN(n5086) );
  XNOR2_X1 U6554 ( .A(n7917), .B(n5410), .ZN(n7718) );
  NAND2_X1 U6555 ( .A1(n4259), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5094) );
  NAND2_X1 U6556 ( .A1(n4816), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5093) );
  INV_X1 U6557 ( .A(n5089), .ZN(n5088) );
  NAND2_X1 U6558 ( .A1(n5088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5096) );
  INV_X1 U6559 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10008) );
  NAND2_X1 U6560 ( .A1(n5089), .A2(n10008), .ZN(n5090) );
  NAND2_X1 U6561 ( .A1(n5096), .A2(n5090), .ZN(n8714) );
  OR2_X1 U6562 ( .A1(n4838), .A2(n8714), .ZN(n5092) );
  NAND2_X1 U6563 ( .A1(n4814), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5091) );
  NAND4_X1 U6564 ( .A1(n5094), .A2(n5093), .A3(n5092), .A4(n5091), .ZN(n8728)
         );
  AND2_X1 U6565 ( .A1(n8728), .A2(n8121), .ZN(n5129) );
  NAND2_X1 U6566 ( .A1(n4814), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5102) );
  INV_X1 U6567 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8398) );
  OR2_X1 U6568 ( .A1(n4260), .A2(n8398), .ZN(n5101) );
  INV_X1 U6569 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6570 ( .A1(n5096), .A2(n5095), .ZN(n5097) );
  NAND2_X1 U6571 ( .A1(n5116), .A2(n5097), .ZN(n8685) );
  OR2_X1 U6572 ( .A1(n4838), .A2(n8685), .ZN(n5100) );
  INV_X1 U6573 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n5098) );
  OR2_X1 U6574 ( .A1(n7899), .A2(n5098), .ZN(n5099) );
  AND4_X1 U6575 ( .A1(n5102), .A2(n5101), .A3(n5100), .A4(n5099), .ZN(n7882)
         );
  NOR2_X1 U6576 ( .A1(n7882), .A2(n5409), .ZN(n5130) );
  OAI21_X1 U6577 ( .B1(n7718), .B2(n5129), .A(n5130), .ZN(n5103) );
  INV_X1 U6578 ( .A(n7718), .ZN(n8003) );
  INV_X1 U6579 ( .A(n5129), .ZN(n8004) );
  INV_X1 U6580 ( .A(n5130), .ZN(n8006) );
  AOI21_X1 U6581 ( .B1(n5104), .B2(n5103), .A(n4692), .ZN(n5128) );
  AND2_X1 U6582 ( .A1(n7715), .A2(n5128), .ZN(n8016) );
  INV_X1 U6583 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n6446) );
  INV_X1 U6584 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5109) );
  MUX2_X1 U6585 ( .A(n6446), .B(n5109), .S(n7393), .Z(n5152) );
  XNOR2_X1 U6586 ( .A(n5152), .B(SI_17_), .ZN(n5171) );
  XNOR2_X1 U6587 ( .A(n5151), .B(n5171), .ZN(n6425) );
  NAND2_X1 U6588 ( .A1(n6425), .A2(n8108), .ZN(n5113) );
  OR2_X1 U6589 ( .A1(n5110), .A2(n4737), .ZN(n5111) );
  XNOR2_X1 U6590 ( .A(n5111), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8434) );
  AOI22_X1 U6591 ( .A1(n5184), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5183), .B2(
        n8434), .ZN(n5112) );
  XNOR2_X1 U6592 ( .A(n8675), .B(n5410), .ZN(n5122) );
  NAND2_X1 U6593 ( .A1(n4259), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5121) );
  INV_X1 U6594 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8421) );
  OR2_X1 U6595 ( .A1(n4260), .A2(n8421), .ZN(n5120) );
  INV_X1 U6596 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5115) );
  NAND2_X1 U6597 ( .A1(n5116), .A2(n5115), .ZN(n5117) );
  NAND2_X1 U6598 ( .A1(n5187), .A2(n5117), .ZN(n8672) );
  OR2_X1 U6599 ( .A1(n4838), .A2(n8672), .ZN(n5119) );
  INV_X1 U6600 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n8673) );
  OR2_X1 U6601 ( .A1(n7897), .A2(n8673), .ZN(n5118) );
  NOR2_X1 U6602 ( .A1(n8649), .A2(n5409), .ZN(n5123) );
  NAND2_X1 U6603 ( .A1(n5122), .A2(n5123), .ZN(n5149) );
  INV_X1 U6604 ( .A(n5122), .ZN(n7731) );
  INV_X1 U6605 ( .A(n5123), .ZN(n5124) );
  NAND2_X1 U6606 ( .A1(n7731), .A2(n5124), .ZN(n5125) );
  NAND2_X1 U6607 ( .A1(n5149), .A2(n5125), .ZN(n8022) );
  INV_X1 U6608 ( .A(n8022), .ZN(n5126) );
  AND2_X1 U6609 ( .A1(n8016), .A2(n5126), .ZN(n5127) );
  NAND2_X1 U6610 ( .A1(n8017), .A2(n5127), .ZN(n7728) );
  INV_X1 U6611 ( .A(n5128), .ZN(n5148) );
  AOI22_X1 U6612 ( .A1(n8007), .A2(n5130), .B1(n5129), .B2(n7718), .ZN(n5146)
         );
  INV_X1 U6613 ( .A(n5131), .ZN(n5145) );
  XNOR2_X1 U6614 ( .A(n5133), .B(n5132), .ZN(n7376) );
  AND2_X1 U6615 ( .A1(n7376), .A2(n5134), .ZN(n5144) );
  INV_X1 U6616 ( .A(n5135), .ZN(n5143) );
  INV_X1 U6617 ( .A(n5136), .ZN(n5137) );
  NAND2_X1 U6618 ( .A1(n5138), .A2(n5137), .ZN(n7323) );
  INV_X1 U6619 ( .A(n5139), .ZN(n5142) );
  INV_X1 U6620 ( .A(n5140), .ZN(n5141) );
  NAND2_X1 U6621 ( .A1(n5142), .A2(n5141), .ZN(n7321) );
  AND2_X1 U6622 ( .A1(n7323), .A2(n7321), .ZN(n7288) );
  OR2_X1 U6623 ( .A1(n5148), .A2(n5147), .ZN(n8018) );
  AND2_X1 U6624 ( .A1(n5149), .A2(n7727), .ZN(n5150) );
  NAND2_X1 U6625 ( .A1(n7728), .A2(n5150), .ZN(n5169) );
  NAND2_X1 U6626 ( .A1(n5255), .A2(n5171), .ZN(n5154) );
  INV_X1 U6627 ( .A(n5152), .ZN(n5153) );
  NAND2_X1 U6628 ( .A1(n5153), .A2(SI_17_), .ZN(n5172) );
  NAND2_X1 U6629 ( .A1(n5154), .A2(n5172), .ZN(n5155) );
  MUX2_X1 U6630 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n7393), .Z(n5174) );
  XNOR2_X1 U6631 ( .A(n5174), .B(SI_18_), .ZN(n5173) );
  NAND2_X1 U6632 ( .A1(n6559), .A2(n8108), .ZN(n5159) );
  NAND2_X1 U6633 ( .A1(n5156), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5157) );
  XNOR2_X1 U6634 ( .A(n5157), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8439) );
  AOI22_X1 U6635 ( .A1(n5184), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5183), .B2(
        n8439), .ZN(n5158) );
  XNOR2_X1 U6636 ( .A(n8831), .B(n5410), .ZN(n7852) );
  NAND2_X1 U6637 ( .A1(n4259), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n5164) );
  INV_X1 U6638 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9932) );
  OR2_X1 U6639 ( .A1(n4260), .A2(n9932), .ZN(n5163) );
  INV_X1 U6640 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n7735) );
  XNOR2_X1 U6641 ( .A(n5187), .B(n7735), .ZN(n7734) );
  OR2_X1 U6642 ( .A1(n4838), .A2(n7734), .ZN(n5162) );
  INV_X1 U6643 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5160) );
  OR2_X1 U6644 ( .A1(n7897), .A2(n5160), .ZN(n5161) );
  NOR2_X1 U6645 ( .A1(n7930), .A2(n5409), .ZN(n5165) );
  NAND2_X1 U6646 ( .A1(n7852), .A2(n5165), .ZN(n5193) );
  INV_X1 U6647 ( .A(n7852), .ZN(n5167) );
  INV_X1 U6648 ( .A(n5165), .ZN(n5166) );
  NAND2_X1 U6649 ( .A1(n5167), .A2(n5166), .ZN(n5168) );
  AND2_X1 U6650 ( .A1(n5193), .A2(n5168), .ZN(n7729) );
  INV_X1 U6651 ( .A(n5173), .ZN(n5170) );
  NAND2_X1 U6652 ( .A1(n5255), .A2(n5199), .ZN(n5177) );
  NAND2_X1 U6653 ( .A1(n5174), .A2(SI_18_), .ZN(n5175) );
  NAND2_X1 U6654 ( .A1(n5177), .A2(n5203), .ZN(n5182) );
  INV_X1 U6655 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n6539) );
  INV_X1 U6656 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n9918) );
  MUX2_X1 U6657 ( .A(n6539), .B(n9918), .S(n7393), .Z(n5179) );
  INV_X1 U6658 ( .A(SI_19_), .ZN(n5178) );
  NAND2_X1 U6659 ( .A1(n5179), .A2(n5178), .ZN(n5200) );
  INV_X1 U6660 ( .A(n5179), .ZN(n5180) );
  NAND2_X1 U6661 ( .A1(n5180), .A2(SI_19_), .ZN(n5181) );
  NAND2_X1 U6662 ( .A1(n5200), .A2(n5181), .ZN(n5201) );
  NAND2_X1 U6663 ( .A1(n6538), .A2(n8108), .ZN(n5186) );
  AOI22_X1 U6664 ( .A1(n5184), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n8511), .B2(
        n5183), .ZN(n5185) );
  XNOR2_X1 U6665 ( .A(n8824), .B(n5410), .ZN(n5195) );
  NAND2_X1 U6666 ( .A1(n4814), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n5192) );
  INV_X1 U6667 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n9920) );
  OR2_X1 U6668 ( .A1(n7899), .A2(n9920), .ZN(n5191) );
  INV_X1 U6669 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8829) );
  OR2_X1 U6670 ( .A1(n4260), .A2(n8829), .ZN(n5190) );
  INV_X1 U6671 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n7860) );
  OAI21_X1 U6672 ( .B1(n5187), .B2(n7735), .A(n7860), .ZN(n5188) );
  NAND2_X1 U6673 ( .A1(n5188), .A2(n5217), .ZN(n8634) );
  OR2_X1 U6674 ( .A1(n4838), .A2(n8634), .ZN(n5189) );
  INV_X1 U6675 ( .A(n8651), .ZN(n8608) );
  NAND2_X1 U6676 ( .A1(n8608), .A2(n4253), .ZN(n5196) );
  XNOR2_X1 U6677 ( .A(n5195), .B(n5196), .ZN(n7855) );
  AND2_X1 U6678 ( .A1(n7855), .A2(n5193), .ZN(n5194) );
  INV_X1 U6679 ( .A(n5195), .ZN(n5197) );
  NAND2_X1 U6680 ( .A1(n5197), .A2(n5196), .ZN(n5198) );
  NAND2_X1 U6681 ( .A1(n5255), .A2(n5230), .ZN(n5206) );
  INV_X1 U6682 ( .A(n5200), .ZN(n5205) );
  INV_X1 U6683 ( .A(n5201), .ZN(n5202) );
  INV_X1 U6684 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n6582) );
  INV_X1 U6685 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n6564) );
  MUX2_X1 U6686 ( .A(n6582), .B(n6564), .S(n7393), .Z(n5208) );
  INV_X1 U6687 ( .A(SI_20_), .ZN(n5207) );
  NAND2_X1 U6688 ( .A1(n5208), .A2(n5207), .ZN(n5231) );
  INV_X1 U6689 ( .A(n5208), .ZN(n5209) );
  NAND2_X1 U6690 ( .A1(n5209), .A2(SI_20_), .ZN(n5210) );
  NAND2_X1 U6691 ( .A1(n6563), .A2(n8108), .ZN(n5213) );
  OR2_X1 U6692 ( .A1(n8110), .A2(n6582), .ZN(n5212) );
  XNOR2_X1 U6693 ( .A(n8613), .B(n5410), .ZN(n5224) );
  NAND2_X1 U6694 ( .A1(n4802), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n5223) );
  INV_X1 U6695 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n5214) );
  OR2_X1 U6696 ( .A1(n4260), .A2(n5214), .ZN(n5222) );
  INV_X1 U6697 ( .A(n5217), .ZN(n5215) );
  NAND2_X1 U6698 ( .A1(n5215), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5241) );
  INV_X1 U6699 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n5216) );
  NAND2_X1 U6700 ( .A1(n5217), .A2(n5216), .ZN(n5218) );
  NAND2_X1 U6701 ( .A1(n5241), .A2(n5218), .ZN(n8057) );
  OR2_X1 U6702 ( .A1(n4838), .A2(n8057), .ZN(n5221) );
  INV_X1 U6703 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n5219) );
  OR2_X1 U6704 ( .A1(n7897), .A2(n5219), .ZN(n5220) );
  NOR2_X1 U6705 ( .A1(n7984), .A2(n5409), .ZN(n5225) );
  NAND2_X1 U6706 ( .A1(n5224), .A2(n5225), .ZN(n5229) );
  INV_X1 U6707 ( .A(n5224), .ZN(n7980) );
  INV_X1 U6708 ( .A(n5225), .ZN(n5226) );
  NAND2_X1 U6709 ( .A1(n7980), .A2(n5226), .ZN(n5227) );
  NAND2_X1 U6710 ( .A1(n5229), .A2(n5227), .ZN(n8056) );
  NAND2_X1 U6711 ( .A1(n8053), .A2(n5229), .ZN(n5248) );
  NAND2_X1 U6712 ( .A1(n5255), .A2(n5253), .ZN(n5236) );
  INV_X1 U6713 ( .A(n5231), .ZN(n5235) );
  INV_X1 U6714 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n6599) );
  INV_X1 U6715 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n6518) );
  MUX2_X1 U6716 ( .A(n6599), .B(n6518), .S(n7393), .Z(n5259) );
  XNOR2_X1 U6717 ( .A(n5259), .B(SI_21_), .ZN(n5256) );
  NAND2_X1 U6718 ( .A1(n6517), .A2(n8108), .ZN(n5239) );
  OR2_X1 U6719 ( .A1(n8110), .A2(n6599), .ZN(n5238) );
  XNOR2_X1 U6720 ( .A(n8812), .B(n5410), .ZN(n5251) );
  NAND2_X1 U6721 ( .A1(n4802), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5247) );
  INV_X1 U6722 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n5240) );
  OR2_X1 U6723 ( .A1(n4260), .A2(n5240), .ZN(n5246) );
  INV_X1 U6724 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n10045) );
  NAND2_X1 U6725 ( .A1(n5241), .A2(n10045), .ZN(n5242) );
  NAND2_X1 U6726 ( .A1(n5279), .A2(n5242), .ZN(n8592) );
  OR2_X1 U6727 ( .A1(n4838), .A2(n8592), .ZN(n5245) );
  INV_X1 U6728 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n5243) );
  OR2_X1 U6729 ( .A1(n7897), .A2(n5243), .ZN(n5244) );
  INV_X1 U6730 ( .A(n8580), .ZN(n8607) );
  NAND2_X1 U6731 ( .A1(n8607), .A2(n8121), .ZN(n5249) );
  XNOR2_X1 U6732 ( .A(n5251), .B(n5249), .ZN(n7978) );
  NAND2_X1 U6733 ( .A1(n5248), .A2(n7978), .ZN(n7981) );
  INV_X1 U6734 ( .A(n5249), .ZN(n5250) );
  NAND2_X1 U6735 ( .A1(n5251), .A2(n5250), .ZN(n5252) );
  INV_X1 U6736 ( .A(n5256), .ZN(n5258) );
  INV_X1 U6737 ( .A(n5259), .ZN(n5260) );
  NAND2_X1 U6738 ( .A1(n5260), .A2(SI_21_), .ZN(n5269) );
  INV_X1 U6739 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n5274) );
  INV_X1 U6740 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9974) );
  MUX2_X1 U6741 ( .A(n5274), .B(n9974), .S(n7393), .Z(n5261) );
  INV_X1 U6742 ( .A(SI_22_), .ZN(n9993) );
  NAND2_X1 U6743 ( .A1(n5261), .A2(n9993), .ZN(n5289) );
  INV_X1 U6744 ( .A(n5261), .ZN(n5262) );
  NAND2_X1 U6745 ( .A1(n5262), .A2(SI_22_), .ZN(n5263) );
  NAND2_X1 U6746 ( .A1(n5289), .A2(n5263), .ZN(n5271) );
  INV_X1 U6747 ( .A(n5271), .ZN(n5264) );
  AND2_X1 U6748 ( .A1(n5269), .A2(n5264), .ZN(n5265) );
  AND2_X1 U6749 ( .A1(n5268), .A2(n5267), .ZN(n5270) );
  NAND2_X1 U6750 ( .A1(n5270), .A2(n5269), .ZN(n5272) );
  NAND2_X1 U6751 ( .A1(n5272), .A2(n5271), .ZN(n5273) );
  NAND2_X1 U6752 ( .A1(n5290), .A2(n5273), .ZN(n6584) );
  NAND2_X1 U6753 ( .A1(n6584), .A2(n8108), .ZN(n5276) );
  OR2_X1 U6754 ( .A1(n8110), .A2(n5274), .ZN(n5275) );
  XNOR2_X1 U6755 ( .A(n8576), .B(n5410), .ZN(n5285) );
  XNOR2_X2 U6756 ( .A(n5287), .B(n5285), .ZN(n8065) );
  INV_X1 U6757 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6758 ( .A1(n5279), .A2(n5278), .ZN(n5280) );
  NAND2_X1 U6759 ( .A1(n5326), .A2(n5280), .ZN(n8573) );
  OR2_X1 U6760 ( .A1(n8573), .A2(n4838), .ZN(n5284) );
  NAND2_X1 U6761 ( .A1(n4259), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n5283) );
  NAND2_X1 U6762 ( .A1(n4816), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n5282) );
  NAND2_X1 U6763 ( .A1(n4814), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n5281) );
  NAND4_X1 U6764 ( .A1(n5284), .A2(n5283), .A3(n5282), .A4(n5281), .ZN(n8599)
         );
  NAND2_X1 U6765 ( .A1(n8599), .A2(n4253), .ZN(n8064) );
  INV_X1 U6766 ( .A(n5285), .ZN(n5286) );
  NOR2_X1 U6767 ( .A1(n5287), .A2(n5286), .ZN(n5288) );
  AOI21_X2 U6768 ( .B1(n8065), .B2(n8064), .A(n5288), .ZN(n5319) );
  INV_X1 U6769 ( .A(n5298), .ZN(n5295) );
  INV_X1 U6770 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n6588) );
  INV_X1 U6771 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n6592) );
  MUX2_X1 U6772 ( .A(n6588), .B(n6592), .S(n7393), .Z(n5292) );
  INV_X1 U6773 ( .A(SI_23_), .ZN(n5291) );
  NAND2_X1 U6774 ( .A1(n5292), .A2(n5291), .ZN(n5303) );
  INV_X1 U6775 ( .A(n5292), .ZN(n5293) );
  NAND2_X1 U6776 ( .A1(n5293), .A2(SI_23_), .ZN(n5294) );
  NAND2_X1 U6777 ( .A1(n5303), .A2(n5294), .ZN(n5296) );
  NAND2_X1 U6778 ( .A1(n5295), .A2(n5296), .ZN(n5299) );
  INV_X1 U6779 ( .A(n5296), .ZN(n5297) );
  NAND2_X1 U6780 ( .A1(n5299), .A2(n5304), .ZN(n6589) );
  NAND2_X1 U6781 ( .A1(n6589), .A2(n8108), .ZN(n5301) );
  OR2_X1 U6782 ( .A1(n8110), .A2(n6588), .ZN(n5300) );
  XNOR2_X1 U6783 ( .A(n8563), .B(n5302), .ZN(n5320) );
  INV_X1 U6784 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n6790) );
  INV_X1 U6785 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n6787) );
  MUX2_X1 U6786 ( .A(n6790), .B(n6787), .S(n7393), .Z(n5336) );
  XNOR2_X1 U6787 ( .A(n5336), .B(SI_24_), .ZN(n5334) );
  XNOR2_X1 U6788 ( .A(n5333), .B(n5334), .ZN(n6786) );
  NAND2_X1 U6789 ( .A1(n6786), .A2(n8108), .ZN(n5306) );
  OR2_X1 U6790 ( .A1(n8110), .A2(n6790), .ZN(n5305) );
  XNOR2_X1 U6791 ( .A(n8550), .B(n5410), .ZN(n5316) );
  INV_X1 U6792 ( .A(n5316), .ZN(n8029) );
  INV_X1 U6793 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n5308) );
  INV_X1 U6794 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5307) );
  OAI21_X1 U6795 ( .B1(n5326), .B2(n5308), .A(n5307), .ZN(n5310) );
  NAND2_X1 U6796 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .ZN(n5309) );
  AND2_X1 U6797 ( .A1(n5310), .A2(n5347), .ZN(n8549) );
  INV_X1 U6798 ( .A(n4838), .ZN(n5327) );
  NAND2_X1 U6799 ( .A1(n8549), .A2(n5327), .ZN(n5314) );
  AOI22_X1 U6800 ( .A1(n4802), .A2(P2_REG0_REG_24__SCAN_IN), .B1(n4816), .B2(
        P2_REG1_REG_24__SCAN_IN), .ZN(n5313) );
  INV_X1 U6801 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n5311) );
  OR2_X1 U6802 ( .A1(n7897), .A2(n5311), .ZN(n5312) );
  NOR2_X1 U6803 ( .A1(n8031), .A2(n5409), .ZN(n5315) );
  INV_X1 U6804 ( .A(n5315), .ZN(n8033) );
  NAND2_X1 U6805 ( .A1(n8029), .A2(n8033), .ZN(n5318) );
  AND2_X1 U6806 ( .A1(n5316), .A2(n5315), .ZN(n5317) );
  AOI21_X1 U6807 ( .B1(n8027), .B2(n5318), .A(n5317), .ZN(n5332) );
  INV_X1 U6808 ( .A(n5319), .ZN(n5321) );
  INV_X1 U6809 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U6810 ( .A1(n4814), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6811 ( .A1(n4816), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5322) );
  OAI211_X1 U6812 ( .C1(n7899), .C2(n5324), .A(n5323), .B(n5322), .ZN(n5325)
         );
  INV_X1 U6813 ( .A(n5325), .ZN(n5329) );
  XNOR2_X1 U6814 ( .A(n5326), .B(P2_REG3_REG_23__SCAN_IN), .ZN(n8561) );
  NAND2_X1 U6815 ( .A1(n8561), .A2(n5327), .ZN(n5328) );
  NAND2_X1 U6816 ( .A1(n5329), .A2(n5328), .ZN(n8315) );
  NAND2_X1 U6817 ( .A1(n8315), .A2(n4253), .ZN(n7960) );
  AOI21_X1 U6818 ( .B1(n8029), .B2(n8031), .A(n7960), .ZN(n5330) );
  NAND2_X1 U6819 ( .A1(n7962), .A2(n5330), .ZN(n5331) );
  INV_X1 U6820 ( .A(n5333), .ZN(n5335) );
  INV_X1 U6821 ( .A(n5336), .ZN(n5337) );
  NAND2_X1 U6822 ( .A1(n5337), .A2(SI_24_), .ZN(n5338) );
  INV_X1 U6823 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n6945) );
  INV_X1 U6824 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n6944) );
  MUX2_X1 U6825 ( .A(n6945), .B(n6944), .S(n7393), .Z(n5341) );
  INV_X1 U6826 ( .A(SI_25_), .ZN(n5340) );
  NAND2_X1 U6827 ( .A1(n5341), .A2(n5340), .ZN(n5352) );
  INV_X1 U6828 ( .A(n5341), .ZN(n5342) );
  NAND2_X1 U6829 ( .A1(n5342), .A2(SI_25_), .ZN(n5343) );
  NAND2_X1 U6830 ( .A1(n5352), .A2(n5343), .ZN(n5353) );
  XNOR2_X1 U6831 ( .A(n5354), .B(n5353), .ZN(n6942) );
  NAND2_X1 U6832 ( .A1(n6942), .A2(n8108), .ZN(n5345) );
  OR2_X1 U6833 ( .A1(n8110), .A2(n6945), .ZN(n5344) );
  XNOR2_X1 U6834 ( .A(n8534), .B(n5410), .ZN(n7992) );
  INV_X1 U6835 ( .A(n5347), .ZN(n5346) );
  NAND2_X1 U6836 ( .A1(n5346), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5363) );
  INV_X1 U6837 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n10039) );
  NAND2_X1 U6838 ( .A1(n5347), .A2(n10039), .ZN(n5348) );
  NAND2_X1 U6839 ( .A1(n5363), .A2(n5348), .ZN(n7997) );
  OR2_X1 U6840 ( .A1(n7997), .A2(n4838), .ZN(n5351) );
  AOI22_X1 U6841 ( .A1(n4259), .A2(P2_REG0_REG_25__SCAN_IN), .B1(n4816), .B2(
        P2_REG1_REG_25__SCAN_IN), .ZN(n5350) );
  NAND2_X1 U6842 ( .A1(n4814), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5349) );
  NOR2_X1 U6843 ( .A1(n8095), .A2(n5409), .ZN(n5370) );
  AND2_X1 U6844 ( .A1(n7992), .A2(n5370), .ZN(n7990) );
  INV_X1 U6845 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7110) );
  INV_X1 U6846 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7082) );
  MUX2_X1 U6847 ( .A(n7110), .B(n7082), .S(n7393), .Z(n5356) );
  INV_X1 U6848 ( .A(SI_26_), .ZN(n5355) );
  NAND2_X1 U6849 ( .A1(n5356), .A2(n5355), .ZN(n5381) );
  INV_X1 U6850 ( .A(n5356), .ZN(n5357) );
  NAND2_X1 U6851 ( .A1(n5357), .A2(SI_26_), .ZN(n5358) );
  AND2_X1 U6852 ( .A1(n5381), .A2(n5358), .ZN(n5379) );
  NAND2_X1 U6853 ( .A1(n7081), .A2(n8108), .ZN(n5360) );
  OR2_X1 U6854 ( .A1(n8110), .A2(n7110), .ZN(n5359) );
  XNOR2_X1 U6855 ( .A(n8786), .B(n5410), .ZN(n5376) );
  INV_X1 U6856 ( .A(n5363), .ZN(n5361) );
  NAND2_X1 U6857 ( .A1(n5361), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5389) );
  INV_X1 U6858 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5362) );
  NAND2_X1 U6859 ( .A1(n5363), .A2(n5362), .ZN(n5364) );
  NAND2_X1 U6860 ( .A1(n5389), .A2(n5364), .ZN(n8513) );
  OR2_X1 U6861 ( .A1(n8513), .A2(n4838), .ZN(n5369) );
  INV_X1 U6862 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n10037) );
  NAND2_X1 U6863 ( .A1(n4816), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5366) );
  INV_X1 U6864 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n8514) );
  OR2_X1 U6865 ( .A1(n7897), .A2(n8514), .ZN(n5365) );
  OAI211_X1 U6866 ( .C1(n10037), .C2(n7899), .A(n5366), .B(n5365), .ZN(n5367)
         );
  INV_X1 U6867 ( .A(n5367), .ZN(n5368) );
  NOR2_X1 U6868 ( .A1(n7955), .A2(n5409), .ZN(n5375) );
  XNOR2_X1 U6869 ( .A(n5376), .B(n5375), .ZN(n8093) );
  INV_X1 U6870 ( .A(n8093), .ZN(n5373) );
  INV_X1 U6871 ( .A(n7992), .ZN(n5372) );
  INV_X1 U6872 ( .A(n5370), .ZN(n5371) );
  NAND2_X1 U6873 ( .A1(n5372), .A2(n5371), .ZN(n8091) );
  AND2_X1 U6874 ( .A1(n5373), .A2(n8091), .ZN(n5374) );
  NAND2_X1 U6875 ( .A1(n8092), .A2(n5374), .ZN(n5378) );
  NAND2_X1 U6876 ( .A1(n5376), .A2(n5375), .ZN(n5377) );
  INV_X1 U6877 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n7189) );
  INV_X1 U6878 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10040) );
  MUX2_X1 U6879 ( .A(n7189), .B(n10040), .S(n7393), .Z(n5384) );
  INV_X1 U6880 ( .A(SI_27_), .ZN(n5383) );
  NAND2_X1 U6881 ( .A1(n5384), .A2(n5383), .ZN(n5414) );
  INV_X1 U6882 ( .A(n5384), .ZN(n5385) );
  NAND2_X1 U6883 ( .A1(n5385), .A2(SI_27_), .ZN(n5386) );
  AND2_X1 U6884 ( .A1(n5414), .A2(n5386), .ZN(n5412) );
  NAND2_X1 U6885 ( .A1(n7156), .A2(n8108), .ZN(n5388) );
  OR2_X1 U6886 ( .A1(n8110), .A2(n7189), .ZN(n5387) );
  XNOR2_X1 U6887 ( .A(n8779), .B(n5410), .ZN(n5398) );
  INV_X1 U6888 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n7953) );
  NAND2_X1 U6889 ( .A1(n5389), .A2(n7953), .ZN(n5390) );
  NAND2_X1 U6890 ( .A1(n5401), .A2(n5390), .ZN(n8495) );
  OR2_X1 U6891 ( .A1(n8495), .A2(n4838), .ZN(n5395) );
  INV_X1 U6892 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n10038) );
  NAND2_X1 U6893 ( .A1(n4259), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5392) );
  NAND2_X1 U6894 ( .A1(n4814), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5391) );
  OAI211_X1 U6895 ( .C1(n4260), .C2(n10038), .A(n5392), .B(n5391), .ZN(n5393)
         );
  INV_X1 U6896 ( .A(n5393), .ZN(n5394) );
  INV_X1 U6897 ( .A(n8096), .ZN(n8473) );
  NAND2_X1 U6898 ( .A1(n8473), .A2(n8121), .ZN(n5396) );
  XNOR2_X1 U6899 ( .A(n5398), .B(n5396), .ZN(n7952) );
  INV_X1 U6900 ( .A(n5396), .ZN(n5397) );
  AND2_X1 U6901 ( .A1(n5398), .A2(n5397), .ZN(n5399) );
  INV_X1 U6902 ( .A(n5401), .ZN(n5400) );
  NAND2_X1 U6903 ( .A1(n5400), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n7912) );
  INV_X1 U6904 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U6905 ( .A1(n5401), .A2(n5482), .ZN(n5402) );
  NAND2_X1 U6906 ( .A1(n7912), .A2(n5402), .ZN(n8478) );
  OR2_X1 U6907 ( .A1(n8478), .A2(n4838), .ZN(n5408) );
  INV_X1 U6908 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n5405) );
  NAND2_X1 U6909 ( .A1(n4814), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5404) );
  NAND2_X1 U6910 ( .A1(n4816), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n5403) );
  OAI211_X1 U6911 ( .C1(n7899), .C2(n5405), .A(n5404), .B(n5403), .ZN(n5406)
         );
  INV_X1 U6912 ( .A(n5406), .ZN(n5407) );
  NOR2_X1 U6913 ( .A1(n7954), .A2(n5409), .ZN(n5411) );
  XNOR2_X1 U6914 ( .A(n5411), .B(n5410), .ZN(n5458) );
  INV_X1 U6915 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n7318) );
  INV_X1 U6916 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10046) );
  MUX2_X1 U6917 ( .A(n7318), .B(n10046), .S(n7393), .Z(n7381) );
  XNOR2_X1 U6918 ( .A(n7381), .B(SI_28_), .ZN(n7378) );
  NAND2_X1 U6919 ( .A1(n7317), .A2(n8108), .ZN(n5417) );
  OR2_X1 U6920 ( .A1(n8110), .A2(n7318), .ZN(n5416) );
  NAND2_X1 U6921 ( .A1(n5419), .A2(n5418), .ZN(n5425) );
  INV_X1 U6922 ( .A(n5425), .ZN(n5421) );
  NAND2_X1 U6923 ( .A1(n5421), .A2(n5420), .ZN(n5427) );
  NAND2_X1 U6924 ( .A1(n5427), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5422) );
  MUX2_X1 U6925 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5422), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n5423) );
  AND2_X1 U6926 ( .A1(n5424), .A2(n5423), .ZN(n7109) );
  NAND2_X1 U6927 ( .A1(n5425), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5426) );
  MUX2_X1 U6928 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5426), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5428) );
  NAND2_X1 U6929 ( .A1(n5428), .A2(n5427), .ZN(n6947) );
  NAND2_X1 U6930 ( .A1(n5430), .A2(n5429), .ZN(n5431) );
  NAND2_X1 U6931 ( .A1(n5431), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5448) );
  INV_X1 U6932 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5447) );
  NAND2_X1 U6933 ( .A1(n5448), .A2(n5447), .ZN(n5450) );
  NAND2_X1 U6934 ( .A1(n5450), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5432) );
  XOR2_X1 U6935 ( .A(n6789), .B(P2_B_REG_SCAN_IN), .Z(n5433) );
  NAND2_X1 U6936 ( .A1(n6947), .A2(n5433), .ZN(n5434) );
  INV_X1 U6937 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n9769) );
  INV_X1 U6938 ( .A(n6947), .ZN(n5445) );
  NOR2_X1 U6939 ( .A1(n5445), .A2(n7109), .ZN(n9771) );
  AOI21_X1 U6940 ( .B1(n9763), .B2(n9769), .A(n9771), .ZN(n8759) );
  NOR4_X1 U6941 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_16__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n5438) );
  NOR4_X1 U6942 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n5437) );
  NOR4_X1 U6943 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_27__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n5436) );
  NOR4_X1 U6944 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_22__SCAN_IN), .ZN(n5435) );
  NAND4_X1 U6945 ( .A1(n5438), .A2(n5437), .A3(n5436), .A4(n5435), .ZN(n5443)
         );
  NOR2_X1 U6946 ( .A1(P2_D_REG_25__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .ZN(
        n10035) );
  NOR4_X1 U6947 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n5441) );
  NOR4_X1 U6948 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n5440) );
  NOR4_X1 U6949 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n5439) );
  NAND4_X1 U6950 ( .A1(n10035), .A2(n5441), .A3(n5440), .A4(n5439), .ZN(n5442)
         );
  OAI21_X1 U6951 ( .B1(n5443), .B2(n5442), .A(n9763), .ZN(n8757) );
  AND2_X1 U6952 ( .A1(n8759), .A2(n8757), .ZN(n6713) );
  NOR2_X1 U6953 ( .A1(n6789), .A2(n7109), .ZN(n9768) );
  INV_X1 U6954 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n9767) );
  NAND2_X1 U6955 ( .A1(n6713), .A2(n8837), .ZN(n5475) );
  AND2_X1 U6956 ( .A1(n7109), .A2(n5445), .ZN(n5446) );
  NAND2_X1 U6957 ( .A1(n6789), .A2(n5446), .ZN(n5970) );
  OR2_X1 U6958 ( .A1(n5448), .A2(n5447), .ZN(n5449) );
  AND2_X1 U6959 ( .A1(n5450), .A2(n5449), .ZN(n9766) );
  INV_X1 U6960 ( .A(n9766), .ZN(n5451) );
  NAND2_X1 U6961 ( .A1(n5970), .A2(n5451), .ZN(n5478) );
  INV_X1 U6962 ( .A(n6000), .ZN(n9764) );
  NAND2_X1 U6963 ( .A1(n8269), .A2(n8765), .ZN(n6696) );
  INV_X1 U6964 ( .A(n6696), .ZN(n5452) );
  NAND2_X1 U6965 ( .A1(n5467), .A2(n5452), .ZN(n5454) );
  INV_X1 U6966 ( .A(n8754), .ZN(n5453) );
  NOR3_X1 U6967 ( .A1(n4527), .A2(n5458), .A3(n8101), .ZN(n5455) );
  AOI21_X1 U6968 ( .B1(n5458), .B2(n4527), .A(n5455), .ZN(n5456) );
  NOR2_X1 U6969 ( .A1(n5460), .A2(n5456), .ZN(n5486) );
  NAND3_X1 U6970 ( .A1(n8773), .A2(n5458), .A3(n8074), .ZN(n5457) );
  OAI21_X1 U6971 ( .B1(n8773), .B2(n5458), .A(n5457), .ZN(n5459) );
  INV_X1 U6972 ( .A(n8765), .ZN(n8268) );
  AND2_X1 U6973 ( .A1(n8268), .A2(n4764), .ZN(n5476) );
  INV_X1 U6974 ( .A(n5476), .ZN(n5461) );
  INV_X1 U6975 ( .A(n5462), .ZN(n8309) );
  NAND2_X1 U6976 ( .A1(n8309), .A2(n8301), .ZN(n5985) );
  INV_X1 U6977 ( .A(n5985), .ZN(n5996) );
  NOR2_X1 U6978 ( .A1(n9843), .A2(n5996), .ZN(n5464) );
  AOI21_X1 U6979 ( .B1(n8773), .B2(n8101), .A(n8085), .ZN(n5465) );
  INV_X1 U6980 ( .A(n5465), .ZN(n5466) );
  NAND2_X1 U6981 ( .A1(n5467), .A2(n5476), .ZN(n7998) );
  INV_X1 U6982 ( .A(n5468), .ZN(n5469) );
  OR2_X1 U6983 ( .A1(n7998), .A2(n8648), .ZN(n8069) );
  OR2_X1 U6984 ( .A1(n7912), .A2(n4838), .ZN(n5474) );
  INV_X1 U6985 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n9940) );
  NAND2_X1 U6986 ( .A1(n4816), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U6987 ( .A1(n4814), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n5470) );
  OAI211_X1 U6988 ( .C1(n7899), .C2(n9940), .A(n5471), .B(n5470), .ZN(n5472)
         );
  INV_X1 U6989 ( .A(n5472), .ZN(n5473) );
  NAND2_X1 U6990 ( .A1(n5474), .A2(n5473), .ZN(n8472) );
  INV_X1 U6991 ( .A(n8472), .ZN(n7893) );
  OAI22_X1 U6992 ( .A1(n8096), .A2(n8069), .B1(n8068), .B2(n7893), .ZN(n5484)
         );
  NAND2_X1 U6993 ( .A1(n5475), .A2(n8754), .ZN(n5480) );
  NOR2_X1 U6994 ( .A1(n5985), .A2(n5476), .ZN(n5477) );
  OR2_X1 U6995 ( .A1(n5478), .A2(n5477), .ZN(n6681) );
  INV_X1 U6996 ( .A(n6681), .ZN(n5479) );
  NAND2_X1 U6997 ( .A1(n5480), .A2(n5479), .ZN(n5481) );
  OAI22_X1 U6998 ( .A1(n8099), .A2(n8478), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5482), .ZN(n5483) );
  OAI21_X1 U6999 ( .B1(n5486), .B2(n5485), .A(n4707), .ZN(P2_U3222) );
  INV_X1 U7000 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n5488) );
  NOR2_X1 U7001 ( .A1(P1_IR_REG_25__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5491) );
  NOR2_X1 U7002 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n5490) );
  NOR2_X1 U7003 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5489) );
  INV_X1 U7004 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5767) );
  NAND4_X1 U7005 ( .A1(n5491), .A2(n5490), .A3(n5489), .A4(n5767), .ZN(n5494)
         );
  INV_X1 U7006 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5947) );
  INV_X1 U7007 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5771) );
  INV_X1 U7008 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n5492) );
  NAND4_X1 U7009 ( .A1(n5947), .A2(n5771), .A3(n5929), .A4(n5492), .ZN(n5493)
         );
  INV_X1 U7010 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5496) );
  INV_X1 U7011 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5501) );
  XNOR2_X1 U7012 ( .A(n5498), .B(n5501), .ZN(n5916) );
  NAND2_X1 U7013 ( .A1(n7317), .A2(n7425), .ZN(n5500) );
  OR2_X1 U7014 ( .A1(n7426), .A2(n10046), .ZN(n5499) );
  INV_X1 U7015 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n7403) );
  XNOR2_X2 U7016 ( .A(n5502), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5512) );
  INV_X1 U7017 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n5504) );
  XNOR2_X2 U7018 ( .A(n5505), .B(n5504), .ZN(n7708) );
  AND2_X2 U7019 ( .A1(n7849), .A2(n5506), .ZN(n5534) );
  NAND2_X1 U7020 ( .A1(n5534), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5516) );
  NAND2_X2 U7021 ( .A1(n7849), .A2(n7708), .ZN(n5537) );
  INV_X1 U7022 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n9995) );
  OR2_X1 U7023 ( .A1(n5537), .A2(n9995), .ZN(n5515) );
  NAND2_X1 U7024 ( .A1(n5621), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5635) );
  INV_X1 U7025 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5634) );
  INV_X1 U7026 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n6915) );
  INV_X1 U7027 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5662) );
  NAND2_X1 U7028 ( .A1(n5677), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5703) );
  INV_X1 U7029 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5702) );
  INV_X1 U7030 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5688) );
  INV_X1 U7031 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n5748) );
  INV_X1 U7032 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n5760) );
  AND2_X1 U7033 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(P1_REG3_REG_19__SCAN_IN), 
        .ZN(n5507) );
  INV_X1 U7034 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8942) );
  INV_X1 U7035 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n9972) );
  INV_X1 U7036 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8907) );
  NAND2_X1 U7037 ( .A1(n5840), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U7038 ( .A1(P1_REG3_REG_26__SCAN_IN), .A2(n5854), .ZN(n5863) );
  INV_X1 U7039 ( .A(n5863), .ZN(n5508) );
  NAND2_X1 U7040 ( .A1(n5508), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n5866) );
  INV_X1 U7041 ( .A(n5866), .ZN(n5509) );
  NAND2_X1 U7042 ( .A1(n5509), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n7836) );
  INV_X1 U7043 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5510) );
  NAND2_X1 U7044 ( .A1(n5866), .A2(n5510), .ZN(n5511) );
  NAND2_X1 U7045 ( .A1(n7836), .A2(n5511), .ZN(n9074) );
  OR2_X1 U7046 ( .A1(n5535), .A2(n9074), .ZN(n5514) );
  INV_X1 U7047 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9075) );
  OR2_X1 U7048 ( .A1(n5549), .A2(n9075), .ZN(n5513) );
  NAND4_X1 U7049 ( .A1(n5516), .A2(n5515), .A3(n5514), .A4(n5513), .ZN(n9087)
         );
  INV_X1 U7050 ( .A(n9087), .ZN(n8862) );
  NAND2_X1 U7051 ( .A1(n9077), .A2(n8862), .ZN(n7840) );
  NAND2_X1 U7052 ( .A1(n5534), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n5521) );
  INV_X1 U7053 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5517) );
  INV_X1 U7054 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n9009) );
  NAND2_X1 U7055 ( .A1(n5843), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n5518) );
  INV_X1 U7056 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6021) );
  INV_X1 U7057 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5522) );
  OR2_X1 U7058 ( .A1(n5531), .A2(n9010), .ZN(n5524) );
  OR2_X1 U7059 ( .A1(n5613), .A2(n6020), .ZN(n5523) );
  NAND3_X2 U7060 ( .A1(n5525), .A2(n5524), .A3(n5523), .ZN(n7664) );
  INV_X1 U7061 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6047) );
  INV_X1 U7062 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6290) );
  INV_X1 U7063 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5526) );
  INV_X1 U7064 ( .A(SI_0_), .ZN(n5528) );
  INV_X1 U7065 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5527) );
  OAI21_X1 U7066 ( .B1(n4761), .B2(n5528), .A(n5527), .ZN(n5530) );
  AND2_X1 U7067 ( .A1(n5530), .A2(n5529), .ZN(n9374) );
  NOR2_X1 U7068 ( .A1(n6298), .A2(n6305), .ZN(n6301) );
  INV_X1 U7069 ( .A(n7664), .ZN(n9683) );
  OR2_X1 U7070 ( .A1(n5532), .A2(n9683), .ZN(n5533) );
  NAND2_X1 U7071 ( .A1(n5534), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5541) );
  INV_X1 U7072 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n6246) );
  OR2_X1 U7073 ( .A1(n5535), .A2(n6246), .ZN(n5540) );
  NAND2_X1 U7074 ( .A1(n5843), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5539) );
  INV_X1 U7075 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5536) );
  OR2_X1 U7076 ( .A1(n5537), .A2(n5536), .ZN(n5538) );
  OR2_X1 U7077 ( .A1(n5613), .A2(n6016), .ZN(n5546) );
  OR2_X1 U7078 ( .A1(n7426), .A2(n6017), .ZN(n5545) );
  NAND2_X1 U7079 ( .A1(n5571), .A2(n5543), .ZN(n5557) );
  OR2_X1 U7080 ( .A1(n5531), .A2(n6139), .ZN(n5544) );
  NAND2_X1 U7081 ( .A1(n4251), .A2(n6252), .ZN(n6251) );
  NAND2_X1 U7082 ( .A1(n7669), .A2(n6676), .ZN(n5548) );
  NAND2_X1 U7083 ( .A1(n6251), .A2(n5548), .ZN(n6269) );
  NAND2_X1 U7084 ( .A1(n4252), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5556) );
  INV_X1 U7085 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U7086 ( .A1(n5620), .A2(n5550), .ZN(n5555) );
  INV_X1 U7087 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n5551) );
  OR2_X1 U7088 ( .A1(n5580), .A2(n5551), .ZN(n5554) );
  INV_X1 U7089 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5552) );
  OR2_X1 U7090 ( .A1(n5537), .A2(n5552), .ZN(n5553) );
  OR2_X1 U7091 ( .A1(n6014), .A2(n5613), .ZN(n5562) );
  OR2_X1 U7092 ( .A1(n7426), .A2(n6015), .ZN(n5561) );
  NAND2_X1 U7093 ( .A1(n5557), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5559) );
  INV_X1 U7094 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5558) );
  XNOR2_X1 U7095 ( .A(n5559), .B(n5558), .ZN(n6072) );
  OR2_X1 U7096 ( .A1(n5531), .A2(n6072), .ZN(n5560) );
  NAND2_X1 U7097 ( .A1(n6432), .A2(n6275), .ZN(n7675) );
  NAND2_X1 U7098 ( .A1(n6269), .A2(n6270), .ZN(n6268) );
  NAND2_X1 U7099 ( .A1(n6432), .A2(n6496), .ZN(n5563) );
  NAND2_X1 U7100 ( .A1(n6268), .A2(n5563), .ZN(n6428) );
  INV_X1 U7101 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5564) );
  INV_X1 U7102 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n5565) );
  OR2_X1 U7103 ( .A1(n5580), .A2(n5565), .ZN(n5568) );
  XNOR2_X1 U7104 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n8919) );
  OR2_X1 U7105 ( .A1(n5535), .A2(n8919), .ZN(n5567) );
  INV_X1 U7106 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6440) );
  OR2_X1 U7107 ( .A1(n5549), .A2(n6440), .ZN(n5566) );
  OR2_X1 U7108 ( .A1(n6018), .A2(n5613), .ZN(n5575) );
  OR2_X1 U7109 ( .A1(n7426), .A2(n6019), .ZN(n5574) );
  OAI21_X1 U7110 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(P1_IR_REG_3__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5570) );
  NAND2_X1 U7111 ( .A1(n5571), .A2(n5570), .ZN(n5572) );
  XNOR2_X1 U7112 ( .A(n5572), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6073) );
  OR2_X1 U7113 ( .A1(n5531), .A2(n6073), .ZN(n5573) );
  INV_X1 U7114 ( .A(n9688), .ZN(n8920) );
  NAND2_X1 U7115 ( .A1(n6486), .A2(n8920), .ZN(n7533) );
  NAND2_X1 U7116 ( .A1(n9005), .A2(n9688), .ZN(n7671) );
  NAND2_X1 U7117 ( .A1(n7533), .A2(n7671), .ZN(n7435) );
  NAND2_X1 U7118 ( .A1(n6428), .A2(n7435), .ZN(n6310) );
  NAND2_X1 U7119 ( .A1(n5576), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5577) );
  XNOR2_X1 U7120 ( .A(n5577), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6075) );
  AOI22_X1 U7121 ( .A1(n5773), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5969), .B2(
        n6075), .ZN(n5578) );
  AOI21_X1 U7122 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5579) );
  NOR2_X1 U7123 ( .A1(n5579), .A2(n5594), .ZN(n6489) );
  NAND2_X1 U7124 ( .A1(n5620), .A2(n6489), .ZN(n5586) );
  INV_X1 U7125 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6057) );
  OR2_X1 U7126 ( .A1(n5580), .A2(n6057), .ZN(n5585) );
  INV_X1 U7127 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n5581) );
  INV_X1 U7128 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5582) );
  OR2_X1 U7129 ( .A1(n5537), .A2(n5582), .ZN(n5583) );
  NAND2_X1 U7130 ( .A1(n7535), .A2(n7534), .ZN(n7528) );
  NAND2_X1 U7131 ( .A1(n6486), .A2(n9688), .ZN(n6311) );
  AND2_X1 U7132 ( .A1(n7528), .A2(n6311), .ZN(n5587) );
  OR2_X1 U7133 ( .A1(n9694), .A2(n8922), .ZN(n5588) );
  OR2_X1 U7134 ( .A1(n6025), .A2(n5613), .ZN(n5592) );
  NOR2_X1 U7135 ( .A1(n5576), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5601) );
  INV_X1 U7136 ( .A(n5601), .ZN(n5589) );
  NAND2_X1 U7137 ( .A1(n5589), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5590) );
  XNOR2_X1 U7138 ( .A(n5590), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6114) );
  AOI22_X1 U7139 ( .A1(n5773), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5969), .B2(
        n6114), .ZN(n5591) );
  NAND2_X1 U7140 ( .A1(n4252), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5598) );
  INV_X1 U7141 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6060) );
  OR2_X1 U7142 ( .A1(n5580), .A2(n6060), .ZN(n5597) );
  INV_X1 U7143 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5593) );
  OR2_X1 U7144 ( .A1(n5537), .A2(n5593), .ZN(n5596) );
  OAI21_X1 U7145 ( .B1(n5594), .B2(P1_REG3_REG_6__SCAN_IN), .A(n5606), .ZN(
        n8972) );
  OR2_X1 U7146 ( .A1(n5535), .A2(n8972), .ZN(n5595) );
  NAND2_X1 U7147 ( .A1(n9003), .A2(n9699), .ZN(n7483) );
  NAND2_X1 U7148 ( .A1(n7679), .A2(n7483), .ZN(n6448) );
  NAND2_X1 U7149 ( .A1(n9699), .A2(n6615), .ZN(n5599) );
  NAND2_X1 U7150 ( .A1(n6449), .A2(n5599), .ZN(n6502) );
  OR2_X1 U7151 ( .A1(n6028), .A2(n5613), .ZN(n5603) );
  NAND2_X1 U7152 ( .A1(n5601), .A2(n5600), .ZN(n5629) );
  NAND2_X1 U7153 ( .A1(n5629), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5615) );
  XNOR2_X1 U7154 ( .A(n5615), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6233) );
  AOI22_X1 U7155 ( .A1(n5773), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5969), .B2(
        n6233), .ZN(n5602) );
  NAND2_X1 U7156 ( .A1(n5603), .A2(n5602), .ZN(n6736) );
  NAND2_X1 U7157 ( .A1(n7417), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5611) );
  INV_X1 U7158 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n5604) );
  OR2_X1 U7159 ( .A1(n5580), .A2(n5604), .ZN(n5610) );
  AND2_X1 U7160 ( .A1(n5606), .A2(n5605), .ZN(n5607) );
  OR2_X1 U7161 ( .A1(n5607), .A2(n5621), .ZN(n6604) );
  OR2_X1 U7162 ( .A1(n5535), .A2(n6604), .ZN(n5609) );
  INV_X1 U7163 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n6511) );
  OR2_X1 U7164 ( .A1(n5549), .A2(n6511), .ZN(n5608) );
  OR2_X1 U7165 ( .A1(n6736), .A2(n6609), .ZN(n7541) );
  NAND2_X1 U7166 ( .A1(n6736), .A2(n6609), .ZN(n7545) );
  NAND2_X1 U7167 ( .A1(n7541), .A2(n7545), .ZN(n7437) );
  NAND2_X1 U7168 ( .A1(n6502), .A2(n7437), .ZN(n6501) );
  INV_X1 U7169 ( .A(n6609), .ZN(n9002) );
  OR2_X1 U7170 ( .A1(n6736), .A2(n9002), .ZN(n5612) );
  OR2_X1 U7171 ( .A1(n6033), .A2(n5613), .ZN(n5619) );
  INV_X1 U7172 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5614) );
  NAND2_X1 U7173 ( .A1(n5615), .A2(n5614), .ZN(n5616) );
  NAND2_X1 U7174 ( .A1(n5616), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5617) );
  XNOR2_X1 U7175 ( .A(n5617), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6234) );
  AOI22_X1 U7176 ( .A1(n5773), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5969), .B2(
        n6234), .ZN(n5618) );
  NAND2_X1 U7177 ( .A1(n5619), .A2(n5618), .ZN(n6636) );
  NAND2_X1 U7178 ( .A1(n7417), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n5627) );
  INV_X1 U7179 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6222) );
  OR2_X1 U7180 ( .A1(n5580), .A2(n6222), .ZN(n5626) );
  OR2_X1 U7181 ( .A1(n5621), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5622) );
  NAND2_X1 U7182 ( .A1(n5635), .A2(n5622), .ZN(n6655) );
  OR2_X1 U7183 ( .A1(n5535), .A2(n6655), .ZN(n5625) );
  INV_X1 U7184 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n5623) );
  OR2_X1 U7185 ( .A1(n5549), .A2(n5623), .ZN(n5624) );
  NAND4_X1 U7186 ( .A1(n5627), .A2(n5626), .A3(n5625), .A4(n5624), .ZN(n9653)
         );
  INV_X1 U7187 ( .A(n9653), .ZN(n6629) );
  OR2_X1 U7188 ( .A1(n6636), .A2(n6629), .ZN(n7495) );
  NAND2_X1 U7189 ( .A1(n6636), .A2(n6629), .ZN(n9646) );
  NAND2_X1 U7190 ( .A1(n6636), .A2(n9653), .ZN(n5628) );
  NAND2_X1 U7191 ( .A1(n6035), .A2(n7425), .ZN(n5633) );
  OR3_X1 U7192 ( .A1(n5629), .A2(P1_IR_REG_8__SCAN_IN), .A3(
        P1_IR_REG_7__SCAN_IN), .ZN(n5630) );
  NAND2_X1 U7193 ( .A1(n5630), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5631) );
  XNOR2_X1 U7194 ( .A(n5631), .B(P1_IR_REG_9__SCAN_IN), .ZN(n9539) );
  AOI22_X1 U7195 ( .A1(n5773), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5969), .B2(
        n9539), .ZN(n5632) );
  NAND2_X1 U7196 ( .A1(n5633), .A2(n5632), .ZN(n9668) );
  NAND2_X1 U7197 ( .A1(n7417), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5640) );
  NAND2_X1 U7198 ( .A1(n5635), .A2(n5634), .ZN(n5636) );
  NAND2_X1 U7199 ( .A1(n5649), .A2(n5636), .ZN(n9664) );
  OR2_X1 U7200 ( .A1(n5535), .A2(n9664), .ZN(n5639) );
  INV_X1 U7201 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6224) );
  OR2_X1 U7202 ( .A1(n5580), .A2(n6224), .ZN(n5638) );
  INV_X1 U7203 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n9665) );
  OR2_X1 U7204 ( .A1(n5549), .A2(n9665), .ZN(n5637) );
  INV_X1 U7205 ( .A(n6809), .ZN(n9001) );
  AND2_X1 U7206 ( .A1(n9668), .A2(n9001), .ZN(n5641) );
  OAI22_X1 U7207 ( .A1(n9645), .A2(n5641), .B1(n9001), .B2(n9668), .ZN(n6743)
         );
  NAND2_X1 U7208 ( .A1(n6039), .A2(n7425), .ZN(n5648) );
  NAND2_X1 U7209 ( .A1(n5642), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5643) );
  MUX2_X1 U7210 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5643), .S(
        P1_IR_REG_10__SCAN_IN), .Z(n5644) );
  INV_X1 U7211 ( .A(n5644), .ZN(n5646) );
  NOR2_X1 U7212 ( .A1(n5646), .A2(n5645), .ZN(n9551) );
  AOI22_X1 U7213 ( .A1(n5773), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5969), .B2(
        n9551), .ZN(n5647) );
  NAND2_X1 U7214 ( .A1(n7417), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n5654) );
  INV_X1 U7215 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6226) );
  OR2_X1 U7216 ( .A1(n5580), .A2(n6226), .ZN(n5653) );
  NAND2_X1 U7217 ( .A1(n5649), .A2(n6915), .ZN(n5650) );
  NAND2_X1 U7218 ( .A1(n5663), .A2(n5650), .ZN(n6918) );
  OR2_X1 U7219 ( .A1(n5535), .A2(n6918), .ZN(n5652) );
  INV_X1 U7220 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6754) );
  OR2_X1 U7221 ( .A1(n5549), .A2(n6754), .ZN(n5651) );
  NAND2_X1 U7222 ( .A1(n9390), .A2(n6879), .ZN(n7557) );
  NAND2_X1 U7223 ( .A1(n7555), .A2(n7557), .ZN(n7442) );
  NAND2_X1 U7224 ( .A1(n6743), .A2(n7442), .ZN(n5656) );
  INV_X1 U7225 ( .A(n6879), .ZN(n9655) );
  OR2_X1 U7226 ( .A1(n9390), .A2(n9655), .ZN(n5655) );
  NAND2_X1 U7227 ( .A1(n5656), .A2(n5655), .ZN(n6971) );
  NAND2_X1 U7228 ( .A1(n5657), .A2(n7425), .ZN(n5660) );
  OR2_X1 U7229 ( .A1(n5645), .A2(n5878), .ZN(n5658) );
  XNOR2_X1 U7230 ( .A(n5658), .B(P1_IR_REG_11__SCAN_IN), .ZN(n6847) );
  AOI22_X1 U7231 ( .A1(n5773), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5969), .B2(
        n6847), .ZN(n5659) );
  NAND2_X1 U7232 ( .A1(n7417), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5668) );
  INV_X1 U7233 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n5661) );
  OR2_X1 U7234 ( .A1(n5580), .A2(n5661), .ZN(n5667) );
  INV_X1 U7235 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n6978) );
  OR2_X1 U7236 ( .A1(n5549), .A2(n6978), .ZN(n5666) );
  AND2_X1 U7237 ( .A1(n5663), .A2(n5662), .ZN(n5664) );
  OR2_X1 U7238 ( .A1(n5664), .A2(n5677), .ZN(n7050) );
  OR2_X1 U7239 ( .A1(n5535), .A2(n7050), .ZN(n5665) );
  INV_X1 U7240 ( .A(n6870), .ZN(n9000) );
  NOR2_X1 U7241 ( .A1(n7114), .A2(n9000), .ZN(n5670) );
  NAND2_X1 U7242 ( .A1(n7114), .A2(n9000), .ZN(n5669) );
  OAI21_X1 U7243 ( .B1(n6971), .B2(n5670), .A(n5669), .ZN(n7032) );
  NAND2_X1 U7244 ( .A1(n6083), .A2(n7425), .ZN(n5676) );
  NAND2_X1 U7245 ( .A1(n5645), .A2(n5671), .ZN(n5673) );
  NAND2_X1 U7246 ( .A1(n5673), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5672) );
  MUX2_X1 U7247 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5672), .S(
        P1_IR_REG_12__SCAN_IN), .Z(n5674) );
  OR2_X1 U7248 ( .A1(n5673), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5695) );
  AND2_X1 U7249 ( .A1(n5674), .A2(n5695), .ZN(n9566) );
  AOI22_X1 U7250 ( .A1(n5773), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5969), .B2(
        n9566), .ZN(n5675) );
  NAND2_X1 U7251 ( .A1(n4252), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n5683) );
  INV_X1 U7252 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6837) );
  OR2_X1 U7253 ( .A1(n5580), .A2(n6837), .ZN(n5682) );
  OR2_X1 U7254 ( .A1(n5677), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U7255 ( .A1(n5703), .A2(n5678), .ZN(n7033) );
  OR2_X1 U7256 ( .A1(n5535), .A2(n7033), .ZN(n5681) );
  INV_X1 U7257 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n5679) );
  OR2_X1 U7258 ( .A1(n5537), .A2(n5679), .ZN(n5680) );
  OR2_X1 U7259 ( .A1(n7038), .A2(n7236), .ZN(n7569) );
  NAND2_X1 U7260 ( .A1(n7038), .A2(n7236), .ZN(n7558) );
  NAND2_X1 U7261 ( .A1(n7569), .A2(n7558), .ZN(n7443) );
  NAND2_X1 U7262 ( .A1(n7032), .A2(n7443), .ZN(n7224) );
  INV_X1 U7263 ( .A(n7236), .ZN(n8999) );
  NAND2_X1 U7264 ( .A1(n7038), .A2(n8999), .ZN(n7223) );
  NAND2_X1 U7265 ( .A1(n6135), .A2(n7425), .ZN(n5687) );
  INV_X1 U7266 ( .A(n5695), .ZN(n5684) );
  NAND2_X1 U7267 ( .A1(n5684), .A2(n5696), .ZN(n5720) );
  NAND2_X1 U7268 ( .A1(n5720), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5685) );
  XNOR2_X1 U7269 ( .A(n5685), .B(P1_IR_REG_14__SCAN_IN), .ZN(n6854) );
  AOI22_X1 U7270 ( .A1(n5773), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5969), .B2(
        n6854), .ZN(n5686) );
  AND2_X1 U7271 ( .A1(n5705), .A2(n5688), .ZN(n5689) );
  NOR2_X1 U7272 ( .A1(n5724), .A2(n5689), .ZN(n7216) );
  NAND2_X1 U7273 ( .A1(n5620), .A2(n7216), .ZN(n5694) );
  INV_X1 U7274 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6835) );
  OR2_X1 U7275 ( .A1(n5580), .A2(n6835), .ZN(n5693) );
  INV_X1 U7276 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7218) );
  OR2_X1 U7277 ( .A1(n5549), .A2(n7218), .ZN(n5692) );
  INV_X1 U7278 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5690) );
  OR2_X1 U7279 ( .A1(n5537), .A2(n5690), .ZN(n5691) );
  INV_X1 U7280 ( .A(n7472), .ZN(n9477) );
  OR2_X1 U7281 ( .A1(n7473), .A2(n9477), .ZN(n5715) );
  INV_X1 U7282 ( .A(n5715), .ZN(n5712) );
  NAND2_X1 U7283 ( .A1(n7473), .A2(n9477), .ZN(n5710) );
  NAND2_X1 U7284 ( .A1(n6128), .A2(n7425), .ZN(n5700) );
  NAND2_X1 U7285 ( .A1(n5695), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5697) );
  MUX2_X1 U7286 ( .A(n5697), .B(P1_IR_REG_31__SCAN_IN), .S(n5696), .Z(n5698)
         );
  NAND2_X1 U7287 ( .A1(n5698), .A2(n5720), .ZN(n6852) );
  INV_X1 U7288 ( .A(n6852), .ZN(n9583) );
  AOI22_X1 U7289 ( .A1(n5773), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n5969), .B2(
        n9583), .ZN(n5699) );
  NAND2_X1 U7290 ( .A1(n4252), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5709) );
  INV_X1 U7291 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n5701) );
  OR2_X1 U7292 ( .A1(n5537), .A2(n5701), .ZN(n5708) );
  INV_X1 U7293 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6841) );
  OR2_X1 U7294 ( .A1(n5580), .A2(n6841), .ZN(n5707) );
  NAND2_X1 U7295 ( .A1(n5703), .A2(n5702), .ZN(n5704) );
  NAND2_X1 U7296 ( .A1(n5705), .A2(n5704), .ZN(n7241) );
  OR2_X1 U7297 ( .A1(n5535), .A2(n7241), .ZN(n5706) );
  INV_X1 U7298 ( .A(n6903), .ZN(n8998) );
  NAND2_X1 U7299 ( .A1(n7256), .A2(n8998), .ZN(n7226) );
  AND2_X1 U7300 ( .A1(n5710), .A2(n7226), .ZN(n5711) );
  AND2_X1 U7301 ( .A1(n7223), .A2(n5714), .ZN(n5713) );
  NAND2_X1 U7302 ( .A1(n7224), .A2(n5713), .ZN(n5719) );
  INV_X1 U7303 ( .A(n5714), .ZN(n5717) );
  OR2_X1 U7304 ( .A1(n7256), .A2(n8998), .ZN(n7225) );
  AND2_X1 U7305 ( .A1(n7225), .A2(n5715), .ZN(n5716) );
  OR2_X1 U7306 ( .A1(n5717), .A2(n5716), .ZN(n5718) );
  NAND2_X1 U7307 ( .A1(n5719), .A2(n5718), .ZN(n9468) );
  NAND2_X1 U7308 ( .A1(n6260), .A2(n7425), .ZN(n5723) );
  OAI21_X1 U7309 ( .B1(n5720), .B2(P1_IR_REG_14__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5721) );
  XNOR2_X1 U7310 ( .A(n5721), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9596) );
  AOI22_X1 U7311 ( .A1(n5773), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n9596), .B2(
        n5969), .ZN(n5722) );
  NOR2_X1 U7312 ( .A1(n5724), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n5725) );
  OR2_X1 U7313 ( .A1(n5736), .A2(n5725), .ZN(n9483) );
  NAND2_X1 U7314 ( .A1(n4252), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n5726) );
  OAI21_X1 U7315 ( .B1(n9483), .B2(n5535), .A(n5726), .ZN(n5730) );
  INV_X1 U7316 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n5728) );
  NAND2_X1 U7317 ( .A1(n7417), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n5727) );
  OAI21_X1 U7318 ( .B1(n5728), .B2(n5580), .A(n5727), .ZN(n5729) );
  NOR2_X1 U7319 ( .A1(n7210), .A2(n8997), .ZN(n5731) );
  NAND2_X1 U7320 ( .A1(n6264), .A2(n7425), .ZN(n5735) );
  BUF_X2 U7321 ( .A(n5732), .Z(n5745) );
  OR2_X1 U7322 ( .A1(n5745), .A2(n5878), .ZN(n5733) );
  XNOR2_X1 U7323 ( .A(n5733), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9607) );
  AOI22_X1 U7324 ( .A1(n5773), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n5969), .B2(
        n9607), .ZN(n5734) );
  OR2_X1 U7325 ( .A1(n5736), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5737) );
  NAND2_X1 U7326 ( .A1(n5749), .A2(n5737), .ZN(n7351) );
  NAND2_X1 U7327 ( .A1(n4252), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n5738) );
  OAI21_X1 U7328 ( .B1(n7351), .B2(n5535), .A(n5738), .ZN(n5741) );
  INV_X1 U7329 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9050) );
  NAND2_X1 U7330 ( .A1(n7417), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n5739) );
  OAI21_X1 U7331 ( .B1(n5580), .B2(n9050), .A(n5739), .ZN(n5740) );
  INV_X1 U7332 ( .A(n9478), .ZN(n7267) );
  NAND2_X1 U7333 ( .A1(n7358), .A2(n7267), .ZN(n7590) );
  NAND2_X1 U7334 ( .A1(n7591), .A2(n7590), .ZN(n7447) );
  NAND2_X1 U7335 ( .A1(n7359), .A2(n7447), .ZN(n5743) );
  NAND2_X1 U7336 ( .A1(n7358), .A2(n9478), .ZN(n5742) );
  NAND2_X1 U7337 ( .A1(n5743), .A2(n5742), .ZN(n9262) );
  INV_X1 U7338 ( .A(n9262), .ZN(n5753) );
  NAND2_X1 U7339 ( .A1(n6425), .A2(n7425), .ZN(n5747) );
  INV_X1 U7340 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5744) );
  NAND2_X1 U7341 ( .A1(n5770), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5755) );
  XNOR2_X1 U7342 ( .A(n5755), .B(P1_IR_REG_17__SCAN_IN), .ZN(n9620) );
  AOI22_X1 U7343 ( .A1(n5773), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n5969), .B2(
        n9620), .ZN(n5746) );
  NAND2_X1 U7344 ( .A1(n5749), .A2(n5748), .ZN(n5750) );
  NAND2_X1 U7345 ( .A1(n5761), .A2(n5750), .ZN(n9265) );
  AOI22_X1 U7346 ( .A1(n5534), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n7417), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n5752) );
  NAND2_X1 U7347 ( .A1(n4252), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n5751) );
  OAI211_X1 U7348 ( .C1(n9265), .C2(n5535), .A(n5752), .B(n5751), .ZN(n9242)
         );
  OR2_X1 U7349 ( .A1(n9344), .A2(n9242), .ZN(n5754) );
  NAND2_X1 U7350 ( .A1(n6559), .A2(n7425), .ZN(n5759) );
  INV_X1 U7351 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5768) );
  NAND2_X1 U7352 ( .A1(n5755), .A2(n5768), .ZN(n5756) );
  NAND2_X1 U7353 ( .A1(n5756), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5757) );
  XNOR2_X1 U7354 ( .A(n5757), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9635) );
  AOI22_X1 U7355 ( .A1(n5773), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n5969), .B2(
        n9635), .ZN(n5758) );
  AND2_X1 U7356 ( .A1(n5761), .A2(n5760), .ZN(n5762) );
  OR2_X1 U7357 ( .A1(n5762), .A2(n5788), .ZN(n9249) );
  AOI22_X1 U7358 ( .A1(n5534), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n7417), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n5764) );
  INV_X1 U7359 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9043) );
  OR2_X1 U7360 ( .A1(n5549), .A2(n9043), .ZN(n5763) );
  OAI211_X1 U7361 ( .C1(n9249), .C2(n5535), .A(n5764), .B(n5763), .ZN(n9272)
         );
  INV_X1 U7362 ( .A(n9272), .ZN(n7343) );
  NAND2_X1 U7363 ( .A1(n9251), .A2(n9272), .ZN(n5766) );
  NAND2_X1 U7364 ( .A1(n9258), .A2(n5766), .ZN(n9222) );
  NAND2_X1 U7365 ( .A1(n6538), .A2(n7425), .ZN(n5775) );
  NAND2_X1 U7366 ( .A1(n5768), .A2(n5767), .ZN(n5769) );
  NAND2_X1 U7367 ( .A1(n4294), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5772) );
  XNOR2_X1 U7368 ( .A(n5772), .B(n5771), .ZN(n9146) );
  AOI22_X1 U7369 ( .A1(n5773), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9473), .B2(
        n5969), .ZN(n5774) );
  INV_X1 U7370 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5776) );
  XNOR2_X1 U7371 ( .A(n5788), .B(n5776), .ZN(n9224) );
  NAND2_X1 U7372 ( .A1(n9224), .A2(n5620), .ZN(n5783) );
  INV_X1 U7373 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9056) );
  INV_X1 U7374 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n5777) );
  OR2_X1 U7375 ( .A1(n5537), .A2(n5777), .ZN(n5780) );
  INV_X1 U7376 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n5778) );
  OR2_X1 U7377 ( .A1(n5549), .A2(n5778), .ZN(n5779) );
  OAI211_X1 U7378 ( .C1(n5580), .C2(n9056), .A(n5780), .B(n5779), .ZN(n5781)
         );
  INV_X1 U7379 ( .A(n5781), .ZN(n5782) );
  NAND2_X1 U7380 ( .A1(n5783), .A2(n5782), .ZN(n9243) );
  OR2_X1 U7381 ( .A1(n9334), .A2(n9243), .ZN(n5785) );
  AND2_X1 U7382 ( .A1(n9334), .A2(n9243), .ZN(n5784) );
  AOI21_X1 U7383 ( .B1(n9222), .B2(n5785), .A(n5784), .ZN(n9202) );
  NAND2_X1 U7384 ( .A1(n6563), .A2(n7425), .ZN(n5787) );
  OR2_X1 U7385 ( .A1(n7426), .A2(n6564), .ZN(n5786) );
  AOI21_X1 U7386 ( .B1(n5788), .B2(P1_REG3_REG_19__SCAN_IN), .A(
        P1_REG3_REG_20__SCAN_IN), .ZN(n5789) );
  OR2_X1 U7387 ( .A1(n5799), .A2(n5789), .ZN(n9215) );
  INV_X1 U7388 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5792) );
  NAND2_X1 U7389 ( .A1(n7417), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5791) );
  NAND2_X1 U7390 ( .A1(n4252), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5790) );
  OAI211_X1 U7391 ( .C1(n5580), .C2(n5792), .A(n5791), .B(n5790), .ZN(n5793)
         );
  INV_X1 U7392 ( .A(n5793), .ZN(n5794) );
  OAI21_X1 U7393 ( .B1(n9215), .B2(n5535), .A(n5794), .ZN(n9233) );
  NAND2_X1 U7394 ( .A1(n9331), .A2(n9233), .ZN(n5796) );
  NOR2_X1 U7395 ( .A1(n9331), .A2(n9233), .ZN(n5795) );
  AOI21_X1 U7396 ( .B1(n9202), .B2(n5796), .A(n5795), .ZN(n9197) );
  NAND2_X1 U7397 ( .A1(n6517), .A2(n7425), .ZN(n5798) );
  OR2_X1 U7398 ( .A1(n7426), .A2(n6518), .ZN(n5797) );
  OR2_X1 U7399 ( .A1(n5799), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n5800) );
  AND2_X1 U7400 ( .A1(n5810), .A2(n5800), .ZN(n9194) );
  NAND2_X1 U7401 ( .A1(n9194), .A2(n5620), .ZN(n5806) );
  INV_X1 U7402 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5803) );
  NAND2_X1 U7403 ( .A1(n7417), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5802) );
  NAND2_X1 U7404 ( .A1(n4252), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5801) );
  OAI211_X1 U7405 ( .C1(n5580), .C2(n5803), .A(n5802), .B(n5801), .ZN(n5804)
         );
  INV_X1 U7406 ( .A(n5804), .ZN(n5805) );
  NAND2_X1 U7407 ( .A1(n5806), .A2(n5805), .ZN(n9175) );
  INV_X1 U7408 ( .A(n9175), .ZN(n9209) );
  NAND2_X1 U7409 ( .A1(n9195), .A2(n9209), .ZN(n7611) );
  NAND2_X1 U7410 ( .A1(n7608), .A2(n7611), .ZN(n9196) );
  NAND2_X1 U7411 ( .A1(n9197), .A2(n9196), .ZN(n9198) );
  NAND2_X1 U7412 ( .A1(n9195), .A2(n9175), .ZN(n5807) );
  NAND2_X1 U7413 ( .A1(n6584), .A2(n7425), .ZN(n5809) );
  OR2_X1 U7414 ( .A1(n7426), .A2(n9974), .ZN(n5808) );
  NAND2_X1 U7415 ( .A1(n5810), .A2(n8942), .ZN(n5811) );
  NAND2_X1 U7416 ( .A1(n5821), .A2(n5811), .ZN(n9170) );
  OR2_X1 U7417 ( .A1(n9170), .A2(n5535), .ZN(n5817) );
  INV_X1 U7418 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5814) );
  NAND2_X1 U7419 ( .A1(n7417), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5813) );
  NAND2_X1 U7420 ( .A1(n4252), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5812) );
  OAI211_X1 U7421 ( .C1(n5580), .C2(n5814), .A(n5813), .B(n5812), .ZN(n5815)
         );
  INV_X1 U7422 ( .A(n5815), .ZN(n5816) );
  NAND2_X1 U7423 ( .A1(n5817), .A2(n5816), .ZN(n9190) );
  NOR2_X1 U7424 ( .A1(n9318), .A2(n9190), .ZN(n5818) );
  INV_X1 U7425 ( .A(n9190), .ZN(n8874) );
  INV_X1 U7426 ( .A(n9318), .ZN(n9173) );
  NAND2_X1 U7427 ( .A1(n6589), .A2(n7425), .ZN(n5820) );
  OR2_X1 U7428 ( .A1(n7426), .A2(n6592), .ZN(n5819) );
  NAND2_X1 U7429 ( .A1(n5821), .A2(n9972), .ZN(n5822) );
  AND2_X1 U7430 ( .A1(n5831), .A2(n5822), .ZN(n9154) );
  NAND2_X1 U7431 ( .A1(n9154), .A2(n5620), .ZN(n5828) );
  INV_X1 U7432 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5825) );
  NAND2_X1 U7433 ( .A1(n7417), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5824) );
  NAND2_X1 U7434 ( .A1(n4252), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5823) );
  OAI211_X1 U7435 ( .C1(n5580), .C2(n5825), .A(n5824), .B(n5823), .ZN(n5826)
         );
  INV_X1 U7436 ( .A(n5826), .ZN(n5827) );
  NAND2_X1 U7437 ( .A1(n5828), .A2(n5827), .ZN(n9176) );
  NAND2_X1 U7438 ( .A1(n9313), .A2(n9176), .ZN(n7622) );
  NAND2_X1 U7439 ( .A1(n6786), .A2(n7425), .ZN(n5830) );
  OR2_X1 U7440 ( .A1(n7426), .A2(n6787), .ZN(n5829) );
  OR2_X1 U7441 ( .A1(n4704), .A2(n5840), .ZN(n9148) );
  INV_X1 U7442 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n5834) );
  NAND2_X1 U7443 ( .A1(n7417), .A2(P1_REG0_REG_24__SCAN_IN), .ZN(n5833) );
  NAND2_X1 U7444 ( .A1(n4252), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5832) );
  OAI211_X1 U7445 ( .C1(n5580), .C2(n5834), .A(n5833), .B(n5832), .ZN(n5835)
         );
  INV_X1 U7446 ( .A(n5835), .ZN(n5836) );
  OAI21_X1 U7447 ( .B1(n9148), .B2(n5535), .A(n5836), .ZN(n9162) );
  INV_X1 U7448 ( .A(n9162), .ZN(n8899) );
  NAND2_X1 U7449 ( .A1(n9309), .A2(n8899), .ZN(n7463) );
  NAND2_X1 U7450 ( .A1(n6942), .A2(n7425), .ZN(n5839) );
  OR2_X1 U7451 ( .A1(n7426), .A2(n6944), .ZN(n5838) );
  OR2_X1 U7452 ( .A1(n5840), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5842) );
  AND2_X1 U7453 ( .A1(n5842), .A2(n5841), .ZN(n9120) );
  NAND2_X1 U7454 ( .A1(n9120), .A2(n5620), .ZN(n5849) );
  INV_X1 U7455 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n5846) );
  NAND2_X1 U7456 ( .A1(n7417), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n5845) );
  NAND2_X1 U7457 ( .A1(n4252), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5844) );
  OAI211_X1 U7458 ( .C1(n5580), .C2(n5846), .A(n5845), .B(n5844), .ZN(n5847)
         );
  INV_X1 U7459 ( .A(n5847), .ZN(n5848) );
  NAND2_X1 U7460 ( .A1(n5849), .A2(n5848), .ZN(n9141) );
  INV_X1 U7461 ( .A(n9141), .ZN(n8908) );
  NAND2_X1 U7462 ( .A1(n9303), .A2(n8908), .ZN(n7629) );
  NAND2_X1 U7463 ( .A1(n9128), .A2(n7629), .ZN(n9124) );
  NAND2_X1 U7464 ( .A1(n9117), .A2(n9124), .ZN(n9116) );
  NAND2_X1 U7465 ( .A1(n9116), .A2(n5850), .ZN(n9098) );
  NAND2_X1 U7466 ( .A1(n7081), .A2(n7425), .ZN(n5852) );
  OR2_X1 U7467 ( .A1(n7426), .A2(n7082), .ZN(n5851) );
  NAND2_X1 U7468 ( .A1(n7417), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5859) );
  INV_X1 U7469 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n5853) );
  OR2_X1 U7470 ( .A1(n5580), .A2(n5853), .ZN(n5858) );
  OAI21_X1 U7471 ( .B1(P1_REG3_REG_26__SCAN_IN), .B2(n5854), .A(n5863), .ZN(
        n9101) );
  OR2_X1 U7472 ( .A1(n5535), .A2(n9101), .ZN(n5857) );
  INV_X1 U7473 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5855) );
  OR2_X1 U7474 ( .A1(n5549), .A2(n5855), .ZN(n5856) );
  NOR2_X1 U7475 ( .A1(n9299), .A2(n9088), .ZN(n7453) );
  NAND2_X1 U7476 ( .A1(n9299), .A2(n9088), .ZN(n7451) );
  NAND2_X1 U7477 ( .A1(n7156), .A2(n7425), .ZN(n5861) );
  OR2_X1 U7478 ( .A1(n7426), .A2(n10040), .ZN(n5860) );
  NAND2_X1 U7479 ( .A1(n5534), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n5871) );
  INV_X1 U7480 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n5862) );
  OR2_X1 U7481 ( .A1(n5537), .A2(n5862), .ZN(n5870) );
  INV_X1 U7482 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n5864) );
  NAND2_X1 U7483 ( .A1(n5864), .A2(n5863), .ZN(n5865) );
  NAND2_X1 U7484 ( .A1(n5866), .A2(n5865), .ZN(n8860) );
  OR2_X1 U7485 ( .A1(n5535), .A2(n8860), .ZN(n5869) );
  INV_X1 U7486 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n5867) );
  OR2_X1 U7487 ( .A1(n5549), .A2(n5867), .ZN(n5868) );
  NAND2_X1 U7488 ( .A1(n9295), .A2(n7813), .ZN(n7523) );
  INV_X1 U7489 ( .A(n7813), .ZN(n9108) );
  AOI21_X1 U7490 ( .B1(n7455), .B2(n5872), .A(n4304), .ZN(n9073) );
  INV_X1 U7491 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5930) );
  INV_X1 U7492 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5931) );
  AND2_X1 U7493 ( .A1(n5930), .A2(n5931), .ZN(n5873) );
  NAND2_X1 U7494 ( .A1(n5877), .A2(n5873), .ZN(n5876) );
  NAND2_X1 U7495 ( .A1(n5876), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5874) );
  XNOR2_X1 U7496 ( .A(n5877), .B(n5930), .ZN(n6565) );
  AND2_X1 U7497 ( .A1(n6565), .A2(n9146), .ZN(n6286) );
  AND2_X1 U7498 ( .A1(n7659), .A2(n6286), .ZN(n6150) );
  OR2_X1 U7499 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5875) );
  NAND2_X1 U7500 ( .A1(n5877), .A2(n5930), .ZN(n5880) );
  NAND2_X1 U7501 ( .A1(n5880), .A2(n5879), .ZN(n5881) );
  NAND2_X1 U7502 ( .A1(n6150), .A2(n7663), .ZN(n5884) );
  INV_X1 U7503 ( .A(n7659), .ZN(n7411) );
  NAND2_X1 U7504 ( .A1(n7411), .A2(n9146), .ZN(n6177) );
  AND2_X2 U7505 ( .A1(n7663), .A2(n6565), .ZN(n6299) );
  OR2_X1 U7506 ( .A1(n6177), .A2(n6299), .ZN(n5883) );
  AND2_X1 U7507 ( .A1(n5884), .A2(n5883), .ZN(n6457) );
  INV_X1 U7508 ( .A(n6565), .ZN(n7701) );
  INV_X1 U7509 ( .A(n9349), .ZN(n9718) );
  INV_X1 U7510 ( .A(n6302), .ZN(n7432) );
  AND2_X1 U7511 ( .A1(n6298), .A2(n6289), .ZN(n6296) );
  NAND2_X1 U7512 ( .A1(n7432), .A2(n6296), .ZN(n5886) );
  NAND2_X1 U7513 ( .A1(n7665), .A2(n7664), .ZN(n5885) );
  NAND2_X1 U7514 ( .A1(n5886), .A2(n5885), .ZN(n6255) );
  NAND2_X1 U7515 ( .A1(n6255), .A2(n7431), .ZN(n5887) );
  NAND2_X1 U7516 ( .A1(n7669), .A2(n5547), .ZN(n7666) );
  INV_X1 U7517 ( .A(n6270), .ZN(n7433) );
  AND2_X1 U7518 ( .A1(n7533), .A2(n7675), .ZN(n5888) );
  NAND2_X1 U7519 ( .A1(n6431), .A2(n5888), .ZN(n7529) );
  NAND2_X1 U7520 ( .A1(n7529), .A2(n7671), .ZN(n6452) );
  NAND2_X1 U7521 ( .A1(n6452), .A2(n7534), .ZN(n5889) );
  NAND2_X1 U7522 ( .A1(n5889), .A2(n7535), .ZN(n5890) );
  NAND2_X1 U7523 ( .A1(n6504), .A2(n7545), .ZN(n6520) );
  NAND2_X1 U7524 ( .A1(n9668), .A2(n6809), .ZN(n7475) );
  AND2_X1 U7525 ( .A1(n7475), .A2(n9646), .ZN(n7552) );
  OR2_X1 U7526 ( .A1(n9668), .A2(n6809), .ZN(n7551) );
  NAND2_X1 U7527 ( .A1(n6748), .A2(n7555), .ZN(n6972) );
  NAND2_X1 U7528 ( .A1(n7114), .A2(n6870), .ZN(n7474) );
  NAND2_X1 U7529 ( .A1(n6972), .A2(n7474), .ZN(n7029) );
  INV_X1 U7530 ( .A(n7029), .ZN(n5891) );
  OR2_X1 U7531 ( .A1(n7114), .A2(n6870), .ZN(n7028) );
  NAND2_X1 U7532 ( .A1(n7569), .A2(n7028), .ZN(n5892) );
  NAND2_X1 U7533 ( .A1(n5892), .A2(n7558), .ZN(n7577) );
  OR2_X1 U7534 ( .A1(n7256), .A2(n6903), .ZN(n7576) );
  NAND2_X1 U7535 ( .A1(n7256), .A2(n6903), .ZN(n7572) );
  NAND2_X1 U7536 ( .A1(n7576), .A2(n7572), .ZN(n7232) );
  NAND2_X1 U7537 ( .A1(n7235), .A2(n7572), .ZN(n7214) );
  INV_X1 U7538 ( .A(n7214), .ZN(n5896) );
  XNOR2_X1 U7539 ( .A(n7473), .B(n7472), .ZN(n7445) );
  OR2_X1 U7540 ( .A1(n7473), .A2(n7472), .ZN(n7579) );
  OR2_X1 U7541 ( .A1(n7210), .A2(n7193), .ZN(n7584) );
  NAND2_X1 U7542 ( .A1(n7210), .A2(n7193), .ZN(n7585) );
  NAND2_X1 U7543 ( .A1(n9475), .A2(n9476), .ZN(n9474) );
  NAND2_X1 U7544 ( .A1(n9474), .A2(n7585), .ZN(n5897) );
  INV_X1 U7545 ( .A(n9242), .ZN(n7336) );
  AND2_X1 U7546 ( .A1(n9344), .A2(n7336), .ZN(n7470) );
  OR2_X1 U7547 ( .A1(n9344), .A2(n7336), .ZN(n9238) );
  NAND2_X1 U7548 ( .A1(n9239), .A2(n7593), .ZN(n9230) );
  INV_X1 U7549 ( .A(n9196), .ZN(n9189) );
  INV_X1 U7550 ( .A(n9233), .ZN(n8888) );
  INV_X1 U7551 ( .A(n7604), .ZN(n7430) );
  AND2_X1 U7552 ( .A1(n9331), .A2(n8888), .ZN(n7600) );
  INV_X1 U7553 ( .A(n7600), .ZN(n5899) );
  INV_X1 U7554 ( .A(n9243), .ZN(n9211) );
  NAND2_X1 U7555 ( .A1(n9334), .A2(n9211), .ZN(n9204) );
  AND2_X1 U7556 ( .A1(n5899), .A2(n9204), .ZN(n5900) );
  OR2_X2 U7557 ( .A1(n9196), .A2(n9185), .ZN(n5902) );
  AND2_X1 U7558 ( .A1(n9229), .A2(n5902), .ZN(n5901) );
  NAND2_X1 U7559 ( .A1(n9230), .A2(n5901), .ZN(n5906) );
  INV_X1 U7560 ( .A(n5902), .ZN(n5904) );
  OR2_X1 U7561 ( .A1(n9334), .A2(n9211), .ZN(n7603) );
  AND2_X1 U7562 ( .A1(n9227), .A2(n7604), .ZN(n9184) );
  AND2_X1 U7563 ( .A1(n9184), .A2(n9189), .ZN(n5903) );
  OR2_X1 U7564 ( .A1(n9318), .A2(n8874), .ZN(n7614) );
  NAND2_X1 U7565 ( .A1(n9318), .A2(n8874), .ZN(n7616) );
  INV_X1 U7566 ( .A(n9158), .ZN(n5908) );
  INV_X1 U7567 ( .A(n9176), .ZN(n8943) );
  NAND2_X1 U7568 ( .A1(n9313), .A2(n8943), .ZN(n7467) );
  NAND2_X1 U7569 ( .A1(n7462), .A2(n7467), .ZN(n9159) );
  NAND2_X1 U7570 ( .A1(n5908), .A2(n5907), .ZN(n9136) );
  INV_X1 U7571 ( .A(n7462), .ZN(n9138) );
  NOR2_X1 U7572 ( .A1(n9137), .A2(n9138), .ZN(n5909) );
  OR2_X1 U7573 ( .A1(n9299), .A2(n9123), .ZN(n7525) );
  INV_X1 U7574 ( .A(n7842), .ZN(n5910) );
  INV_X1 U7575 ( .A(n7455), .ZN(n5911) );
  XNOR2_X1 U7576 ( .A(n5912), .B(n5911), .ZN(n5915) );
  OR2_X1 U7577 ( .A1(n7659), .A2(n9146), .ZN(n5914) );
  NAND2_X1 U7578 ( .A1(n7663), .A2(n7701), .ZN(n5913) );
  NAND2_X1 U7579 ( .A1(n5914), .A2(n5913), .ZN(n9651) );
  NAND2_X1 U7580 ( .A1(n7411), .A2(n7663), .ZN(n7654) );
  OR2_X1 U7581 ( .A1(n7654), .A2(n5916), .ZN(n9212) );
  NOR2_X1 U7582 ( .A1(n7813), .A2(n9212), .ZN(n5922) );
  INV_X1 U7583 ( .A(n5916), .ZN(n6199) );
  NAND2_X1 U7584 ( .A1(n5534), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U7585 ( .A1(n7417), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5920) );
  OR2_X1 U7586 ( .A1(n5535), .A2(n7836), .ZN(n5919) );
  INV_X1 U7587 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n5917) );
  OR2_X1 U7588 ( .A1(n5549), .A2(n5917), .ZN(n5918) );
  NAND4_X1 U7589 ( .A1(n5921), .A2(n5920), .A3(n5919), .A4(n5918), .ZN(n8996)
         );
  INV_X1 U7590 ( .A(n9299), .ZN(n9104) );
  INV_X1 U7591 ( .A(n9331), .ZN(n9219) );
  INV_X1 U7592 ( .A(n9344), .ZN(n9269) );
  OR2_X1 U7593 ( .A1(n6439), .A2(n6488), .ZN(n6458) );
  INV_X1 U7594 ( .A(n9699), .ZN(n8973) );
  INV_X1 U7595 ( .A(n6736), .ZN(n6510) );
  AND2_X1 U7596 ( .A1(n6459), .A2(n6510), .ZN(n6530) );
  INV_X1 U7597 ( .A(n6636), .ZN(n6529) );
  INV_X1 U7598 ( .A(n7114), .ZN(n6977) );
  INV_X1 U7599 ( .A(n7038), .ZN(n9500) );
  NAND2_X1 U7600 ( .A1(n7035), .A2(n9500), .ZN(n7240) );
  NAND2_X1 U7601 ( .A1(n9219), .A2(n9223), .ZN(n9181) );
  NAND2_X1 U7602 ( .A1(n9173), .A2(n9167), .ZN(n9168) );
  INV_X1 U7603 ( .A(n9309), .ZN(n8913) );
  INV_X1 U7604 ( .A(n9077), .ZN(n5925) );
  NAND2_X1 U7605 ( .A1(n5925), .A2(n9091), .ZN(n7835) );
  OAI21_X1 U7606 ( .B1(n9091), .B2(n5925), .A(n7835), .ZN(n9079) );
  INV_X1 U7607 ( .A(n7663), .ZN(n6519) );
  NAND2_X1 U7608 ( .A1(n7659), .A2(n6519), .ZN(n6287) );
  OR2_X1 U7609 ( .A1(n6287), .A2(n7701), .ZN(n9714) );
  OAI22_X1 U7610 ( .A1(n9079), .A2(n9714), .B1(n5925), .B2(n9713), .ZN(n5926)
         );
  NAND2_X1 U7611 ( .A1(n5928), .A2(n5927), .ZN(n9359) );
  NAND2_X1 U7612 ( .A1(n5945), .A2(n5947), .ZN(n5932) );
  NAND2_X1 U7613 ( .A1(n5932), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5933) );
  XNOR2_X1 U7614 ( .A(n5933), .B(P1_IR_REG_24__SCAN_IN), .ZN(n5941) );
  INV_X1 U7615 ( .A(n5941), .ZN(n6788) );
  NOR2_X1 U7616 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5934) );
  NAND2_X1 U7617 ( .A1(n5945), .A2(n5934), .ZN(n5935) );
  INV_X1 U7618 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5936) );
  XNOR2_X1 U7619 ( .A(n5937), .B(P1_IR_REG_25__SCAN_IN), .ZN(n5942) );
  INV_X1 U7620 ( .A(n5942), .ZN(n6943) );
  NAND3_X1 U7621 ( .A1(n6943), .A2(P1_B_REG_SCAN_IN), .A3(n6788), .ZN(n5938)
         );
  OAI211_X1 U7622 ( .C1(P1_B_REG_SCAN_IN), .C2(n6788), .A(n5944), .B(n5938), 
        .ZN(n9677) );
  OR2_X1 U7623 ( .A1(n9677), .A2(P1_D_REG_1__SCAN_IN), .ZN(n5940) );
  INV_X1 U7624 ( .A(n5944), .ZN(n7083) );
  NAND2_X1 U7625 ( .A1(n7083), .A2(n6943), .ZN(n5939) );
  NOR2_X1 U7626 ( .A1(n9389), .A2(n7663), .ZN(n6285) );
  NOR2_X1 U7627 ( .A1(n6281), .A2(n6285), .ZN(n5951) );
  AND2_X1 U7628 ( .A1(n5942), .A2(n5941), .ZN(n5943) );
  INV_X1 U7629 ( .A(n5945), .ZN(n5946) );
  NAND2_X1 U7630 ( .A1(n5946), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5948) );
  XNOR2_X1 U7631 ( .A(n5948), .B(n5947), .ZN(n6590) );
  AND2_X1 U7632 ( .A1(n6590), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5949) );
  NAND2_X1 U7633 ( .A1(n6151), .A2(n5949), .ZN(n9372) );
  OR2_X1 U7634 ( .A1(n7654), .A2(n6286), .ZN(n6203) );
  INV_X1 U7635 ( .A(n6203), .ZN(n5950) );
  NOR2_X1 U7636 ( .A1(n9372), .A2(n5950), .ZN(n6282) );
  AND2_X1 U7637 ( .A1(n5951), .A2(n6282), .ZN(n6132) );
  OR2_X1 U7638 ( .A1(n9677), .A2(P1_D_REG_0__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U7639 ( .A1(n7083), .A2(n6788), .ZN(n5952) );
  AND2_X1 U7640 ( .A1(n5953), .A2(n5952), .ZN(n9373) );
  NOR2_X1 U7641 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n5957) );
  NOR4_X1 U7642 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n5956) );
  NOR4_X1 U7643 ( .A1(P1_D_REG_8__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n5955) );
  NOR4_X1 U7644 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n5954) );
  NAND4_X1 U7645 ( .A1(n5957), .A2(n5956), .A3(n5955), .A4(n5954), .ZN(n5963)
         );
  NOR4_X1 U7646 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_18__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n5961) );
  NOR4_X1 U7647 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_14__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n5960) );
  NOR4_X1 U7648 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n5959) );
  NOR4_X1 U7649 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n5958) );
  NAND4_X1 U7650 ( .A1(n5961), .A2(n5960), .A3(n5959), .A4(n5958), .ZN(n5962)
         );
  NOR2_X1 U7651 ( .A1(n5963), .A2(n5962), .ZN(n5964) );
  OR2_X1 U7652 ( .A1(n9677), .A2(n5964), .ZN(n6130) );
  AND2_X1 U7653 ( .A1(n9373), .A2(n6130), .ZN(n6165) );
  AND2_X2 U7654 ( .A1(n6132), .A2(n6165), .ZN(n9731) );
  INV_X1 U7655 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n5965) );
  INV_X1 U7656 ( .A(n6590), .ZN(n5967) );
  OR2_X1 U7657 ( .A1(n6151), .A2(n5967), .ZN(n6044) );
  NOR2_X1 U7658 ( .A1(n6044), .A2(P1_U3084), .ZN(P1_U4006) );
  OR2_X1 U7659 ( .A1(n7654), .A2(n5967), .ZN(n5968) );
  NAND2_X1 U7660 ( .A1(n6044), .A2(n5968), .ZN(n6045) );
  OAI21_X1 U7661 ( .B1(n6045), .B2(n5969), .A(P1_STATE_REG_SCAN_IN), .ZN(
        P1_U3083) );
  OR2_X1 U7662 ( .A1(n5970), .A2(P2_U3152), .ZN(n5986) );
  OR2_X2 U7663 ( .A1(n5986), .A2(n9766), .ZN(n8328) );
  INV_X1 U7664 ( .A(n8328), .ZN(P2_U3966) );
  INV_X1 U7665 ( .A(n5975), .ZN(n5972) );
  NOR3_X1 U7666 ( .A1(n8103), .A2(n5972), .A3(n5971), .ZN(n5978) );
  NAND2_X1 U7667 ( .A1(n8085), .A2(n8121), .ZN(n8040) );
  OR3_X1 U7668 ( .A1(n8040), .A2(n7073), .A3(n5973), .ZN(n5974) );
  OAI21_X1 U7669 ( .B1(n8103), .B2(n5975), .A(n5974), .ZN(n5977) );
  MUX2_X1 U7670 ( .A(n5978), .B(n5977), .S(n5976), .Z(n5982) );
  OAI22_X1 U7671 ( .A1(n8074), .A2(n9837), .B1(n8068), .B2(n7062), .ZN(n5981)
         );
  NAND2_X1 U7672 ( .A1(n8059), .A2(n8322), .ZN(n5979) );
  NAND2_X1 U7673 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n6375) );
  OAI211_X1 U7674 ( .C1(n8099), .C2(n6963), .A(n5979), .B(n6375), .ZN(n5980)
         );
  OR3_X1 U7675 ( .A1(n5982), .A2(n5981), .A3(n5980), .ZN(P2_U3233) );
  NAND2_X1 U7676 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .ZN(n5991) );
  INV_X1 U7677 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n5983) );
  INV_X1 U7678 ( .A(n5984), .ZN(n5990) );
  NOR2_X1 U7679 ( .A1(n5990), .A2(n5991), .ZN(n6336) );
  NAND2_X1 U7680 ( .A1(n6000), .A2(n5985), .ZN(n5987) );
  NAND2_X1 U7681 ( .A1(n9766), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8311) );
  NAND3_X1 U7682 ( .A1(n5987), .A2(n8311), .A3(n5986), .ZN(n5988) );
  NAND2_X1 U7683 ( .A1(n5988), .A2(n5997), .ZN(n5993) );
  NAND2_X1 U7684 ( .A1(n5993), .A2(n8328), .ZN(n5992) );
  INV_X1 U7685 ( .A(n5992), .ZN(n5989) );
  NOR3_X4 U7686 ( .A1(n5989), .A2(n5468), .A3(n7904), .ZN(n9733) );
  AOI211_X1 U7687 ( .C1(n5991), .C2(n5990), .A(n6336), .B(n9738), .ZN(n6007)
         );
  NAND2_X1 U7688 ( .A1(n5992), .A2(n5468), .ZN(n9739) );
  NOR2_X1 U7689 ( .A1(n9739), .A2(n6335), .ZN(n6006) );
  NAND2_X1 U7690 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n5995) );
  INV_X1 U7691 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n9870) );
  MUX2_X1 U7692 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n9870), .S(n6335), .Z(n5994)
         );
  NOR2_X1 U7693 ( .A1(n5994), .A2(n5995), .ZN(n6326) );
  INV_X1 U7694 ( .A(n7904), .ZN(n8307) );
  AOI211_X1 U7695 ( .C1(n5995), .C2(n5994), .A(n6326), .B(n9740), .ZN(n6005)
         );
  NAND2_X1 U7696 ( .A1(n6000), .A2(n5996), .ZN(n5998) );
  NAND2_X1 U7697 ( .A1(n5998), .A2(n5997), .ZN(n6002) );
  INV_X1 U7698 ( .A(n8311), .ZN(n5999) );
  OR2_X1 U7699 ( .A1(n6000), .A2(n5999), .ZN(n6001) );
  NAND2_X1 U7700 ( .A1(n6002), .A2(n6001), .ZN(n9736) );
  INV_X1 U7701 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6003) );
  OAI22_X1 U7702 ( .A1(n9736), .A2(n6003), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n4801), .ZN(n6004) );
  OR4_X1 U7703 ( .A1(n6007), .A2(n6006), .A3(n6005), .A4(n6004), .ZN(P2_U3246)
         );
  NAND2_X1 U7704 ( .A1(n4761), .A2(P2_U3152), .ZN(n7949) );
  INV_X1 U7705 ( .A(n7949), .ZN(n6586) );
  INV_X1 U7706 ( .A(n6586), .ZN(n7319) );
  NOR2_X1 U7707 ( .A1(n4761), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7399) );
  INV_X2 U7708 ( .A(n7399), .ZN(n7947) );
  OAI222_X1 U7709 ( .A1(n6010), .A2(P2_U3152), .B1(n7319), .B2(n6016), .C1(
        n6009), .C2(n7947), .ZN(P2_U3356) );
  OAI222_X1 U7710 ( .A1(n6335), .A2(P2_U3152), .B1(n7319), .B2(n6020), .C1(
        n6011), .C2(n7947), .ZN(P2_U3357) );
  OAI222_X1 U7711 ( .A1(n8338), .A2(P2_U3152), .B1(n7319), .B2(n6014), .C1(
        n6012), .C2(n7947), .ZN(P2_U3355) );
  OAI222_X1 U7712 ( .A1(n6359), .A2(P2_U3152), .B1(n7949), .B2(n6018), .C1(
        n6013), .C2(n7947), .ZN(P2_U3354) );
  AND2_X1 U7713 ( .A1(n4761), .A2(P1_U3084), .ZN(n6426) );
  NOR2_X1 U7714 ( .A1(n4761), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7407) );
  OAI222_X1 U7715 ( .A1(n4258), .A2(n6015), .B1(n7850), .B2(n6014), .C1(
        P1_U3084), .C2(n6072), .ZN(P1_U3350) );
  OAI222_X1 U7716 ( .A1(n4258), .A2(n6017), .B1(n7850), .B2(n6016), .C1(
        P1_U3084), .C2(n6139), .ZN(P1_U3351) );
  OAI222_X1 U7717 ( .A1(n4258), .A2(n6019), .B1(P1_U3084), .B2(n6073), .C1(
        n7850), .C2(n6018), .ZN(P1_U3349) );
  OAI222_X1 U7718 ( .A1(n4258), .A2(n6021), .B1(n7850), .B2(n6020), .C1(
        P1_U3084), .C2(n9010), .ZN(P1_U3352) );
  OAI222_X1 U7719 ( .A1(n8350), .A2(P2_U3152), .B1(n7319), .B2(n6023), .C1(
        n6022), .C2(n7947), .ZN(P2_U3353) );
  INV_X1 U7720 ( .A(n6075), .ZN(n9510) );
  OAI222_X1 U7721 ( .A1(n4258), .A2(n9944), .B1(n7850), .B2(n6023), .C1(
        P1_U3084), .C2(n9510), .ZN(P1_U3348) );
  OAI222_X1 U7722 ( .A1(n6404), .A2(P2_U3152), .B1(n7949), .B2(n6025), .C1(
        n6024), .C2(n7947), .ZN(P2_U3352) );
  INV_X1 U7723 ( .A(n6114), .ZN(n6059) );
  OAI222_X1 U7724 ( .A1(n4258), .A2(n6026), .B1(n7850), .B2(n6025), .C1(
        P1_U3084), .C2(n6059), .ZN(P1_U3347) );
  OAI222_X1 U7725 ( .A1(n6370), .A2(P2_U3152), .B1(n7949), .B2(n6028), .C1(
        n6027), .C2(n7947), .ZN(P2_U3351) );
  INV_X1 U7726 ( .A(n6233), .ZN(n6066) );
  OAI222_X1 U7727 ( .A1(n4258), .A2(n6029), .B1(n7850), .B2(n6028), .C1(
        P1_U3084), .C2(n6066), .ZN(P1_U3346) );
  INV_X1 U7728 ( .A(n9372), .ZN(n9678) );
  INV_X1 U7729 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6031) );
  NAND2_X1 U7730 ( .A1(n6281), .A2(n9678), .ZN(n6030) );
  OAI21_X1 U7731 ( .B1(n9678), .B2(n6031), .A(n6030), .ZN(P1_U3441) );
  OAI222_X1 U7732 ( .A1(n6389), .A2(P2_U3152), .B1(n7319), .B2(n6033), .C1(
        n6032), .C2(n7947), .ZN(P2_U3350) );
  INV_X1 U7733 ( .A(n6234), .ZN(n9522) );
  OAI222_X1 U7734 ( .A1(n4258), .A2(n6034), .B1(n7850), .B2(n6033), .C1(
        P1_U3084), .C2(n9522), .ZN(P1_U3345) );
  INV_X1 U7735 ( .A(n6035), .ZN(n6038) );
  INV_X1 U7736 ( .A(n9539), .ZN(n6225) );
  OAI222_X1 U7737 ( .A1(n7850), .A2(n6038), .B1(n6225), .B2(P1_U3084), .C1(
        n6036), .C2(n4258), .ZN(P1_U3344) );
  INV_X1 U7738 ( .A(n6406), .ZN(n6419) );
  OAI222_X1 U7739 ( .A1(P2_U3152), .A2(n6419), .B1(n7319), .B2(n6038), .C1(
        n6037), .C2(n7947), .ZN(P2_U3349) );
  INV_X1 U7740 ( .A(n6549), .ZN(n6424) );
  INV_X1 U7741 ( .A(n6039), .ZN(n6042) );
  OAI222_X1 U7742 ( .A1(P2_U3152), .A2(n6424), .B1(n7319), .B2(n6042), .C1(
        n6040), .C2(n7947), .ZN(P2_U3348) );
  INV_X1 U7743 ( .A(n5657), .ZN(n6055) );
  INV_X1 U7744 ( .A(n6847), .ZN(n6839) );
  INV_X1 U7745 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6041) );
  OAI222_X1 U7746 ( .A1(n7850), .A2(n6055), .B1(n6839), .B2(P1_U3084), .C1(
        n6041), .C2(n4258), .ZN(P1_U3342) );
  INV_X1 U7747 ( .A(n9551), .ZN(n6227) );
  OAI222_X1 U7748 ( .A1(n4258), .A2(n6043), .B1(n6227), .B2(P1_U3084), .C1(
        n7850), .C2(n6042), .ZN(P1_U3343) );
  INV_X1 U7749 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n9890) );
  INV_X1 U7750 ( .A(n6044), .ZN(n6160) );
  NOR2_X1 U7751 ( .A1(n6045), .A2(P1_U3084), .ZN(n6065) );
  NAND2_X1 U7752 ( .A1(n6065), .A2(n6199), .ZN(n6078) );
  INV_X1 U7753 ( .A(n6046), .ZN(n6063) );
  OR2_X1 U7754 ( .A1(n6078), .A2(n6063), .ZN(n9640) );
  INV_X1 U7755 ( .A(n9640), .ZN(n9622) );
  NAND3_X1 U7756 ( .A1(n9622), .A2(P1_IR_REG_0__SCAN_IN), .A3(n6047), .ZN(
        n6053) );
  AOI21_X1 U7757 ( .B1(n6046), .B2(n6047), .A(P1_IR_REG_0__SCAN_IN), .ZN(n6049) );
  OAI21_X1 U7758 ( .B1(n6046), .B2(P1_REG2_REG_0__SCAN_IN), .A(n6199), .ZN(
        n6048) );
  AOI21_X1 U7759 ( .B1(n6048), .B2(n4425), .A(P1_U3084), .ZN(n6159) );
  OAI21_X1 U7760 ( .B1(n6049), .B2(n6048), .A(n6159), .ZN(n6050) );
  OAI21_X1 U7761 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n6290), .A(n6050), .ZN(n6051) );
  NAND2_X1 U7762 ( .A1(P1_U3083), .A2(n6051), .ZN(n6052) );
  OAI211_X1 U7763 ( .C1(n9890), .C2(n9643), .A(n6053), .B(n6052), .ZN(P1_U3241) );
  INV_X1 U7764 ( .A(n8370), .ZN(n6543) );
  INV_X1 U7765 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6054) );
  OAI222_X1 U7766 ( .A1(P2_U3152), .A2(n6543), .B1(n7319), .B2(n6055), .C1(
        n6054), .C2(n7947), .ZN(P2_U3347) );
  NAND2_X1 U7767 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6075), .ZN(n6058) );
  INV_X1 U7768 ( .A(n6072), .ZN(n6099) );
  INV_X1 U7769 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9723) );
  NAND2_X1 U7770 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n9013) );
  OAI21_X1 U7771 ( .B1(n9723), .B2(n9010), .A(n9015), .ZN(n6141) );
  XNOR2_X1 U7772 ( .A(n6139), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n6140) );
  INV_X1 U7773 ( .A(n6139), .ZN(n6071) );
  AOI22_X1 U7774 ( .A1(n6141), .A2(n6140), .B1(n6071), .B2(
        P1_REG1_REG_2__SCAN_IN), .ZN(n6096) );
  MUX2_X1 U7775 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n5551), .S(n6072), .Z(n6095)
         );
  NOR2_X1 U7776 ( .A1(n6096), .A2(n6095), .ZN(n6094) );
  AOI21_X1 U7777 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n6099), .A(n6094), .ZN(
        n9031) );
  INV_X1 U7778 ( .A(n6073), .ZN(n9025) );
  NOR2_X1 U7779 ( .A1(n9025), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6056) );
  AOI21_X1 U7780 ( .B1(n9025), .B2(P1_REG1_REG_4__SCAN_IN), .A(n6056), .ZN(
        n9030) );
  NAND2_X1 U7781 ( .A1(n9031), .A2(n9030), .ZN(n9029) );
  MUX2_X1 U7782 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6057), .S(n6075), .Z(n9515)
         );
  MUX2_X1 U7783 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n6060), .S(n6114), .Z(n6107)
         );
  NAND2_X1 U7784 ( .A1(n6106), .A2(n6107), .ZN(n6105) );
  AOI22_X1 U7785 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6066), .B1(n6233), .B2(
        n5604), .ZN(n6061) );
  AOI21_X1 U7786 ( .B1(n6062), .B2(n6061), .A(n6223), .ZN(n6082) );
  INV_X1 U7787 ( .A(n9643), .ZN(n9012) );
  AND2_X1 U7788 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6601) );
  AND2_X1 U7789 ( .A1(n5916), .A2(n6063), .ZN(n6064) );
  NAND2_X1 U7790 ( .A1(n6065), .A2(n6064), .ZN(n9523) );
  NOR2_X1 U7791 ( .A1(n9523), .A2(n6066), .ZN(n6067) );
  AOI211_X1 U7792 ( .C1(n9012), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n6601), .B(
        n6067), .ZN(n6081) );
  NOR2_X1 U7793 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6233), .ZN(n6068) );
  AOI21_X1 U7794 ( .B1(n6233), .B2(P1_REG2_REG_7__SCAN_IN), .A(n6068), .ZN(
        n6077) );
  NAND2_X1 U7795 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6158) );
  INV_X1 U7796 ( .A(n6158), .ZN(n9017) );
  INV_X1 U7797 ( .A(n9010), .ZN(n6069) );
  NAND2_X1 U7798 ( .A1(n6069), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7799 ( .A1(n9016), .A2(n6070), .ZN(n6144) );
  XNOR2_X1 U7800 ( .A(n6139), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6145) );
  XOR2_X1 U7801 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n6072), .Z(n6092) );
  NOR2_X1 U7802 ( .A1(n6093), .A2(n6092), .ZN(n6091) );
  XNOR2_X1 U7803 ( .A(n6073), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n9027) );
  NOR2_X1 U7804 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6075), .ZN(n6074) );
  AOI21_X1 U7805 ( .B1(n6075), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6074), .ZN(
        n9509) );
  XNOR2_X1 U7806 ( .A(n6114), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n6110) );
  NOR2_X1 U7807 ( .A1(n6109), .A2(n6110), .ZN(n6108) );
  OAI21_X1 U7808 ( .B1(n6077), .B2(n6076), .A(n6232), .ZN(n6079) );
  NOR2_X1 U7809 ( .A1(n6078), .A2(n6046), .ZN(n9526) );
  NAND2_X1 U7810 ( .A1(n6079), .A2(n9526), .ZN(n6080) );
  OAI211_X1 U7811 ( .C1(n6082), .C2(n9640), .A(n6081), .B(n6080), .ZN(P1_U3248) );
  INV_X1 U7812 ( .A(n6083), .ZN(n6104) );
  AOI22_X1 U7813 ( .A1(n9566), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n6426), .ZN(n6084) );
  OAI21_X1 U7814 ( .B1(n6104), .B2(n7850), .A(n6084), .ZN(P1_U3341) );
  INV_X1 U7815 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6088) );
  INV_X1 U7816 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n9917) );
  NAND2_X1 U7817 ( .A1(n7417), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6086) );
  INV_X1 U7818 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n7709) );
  OR2_X1 U7819 ( .A1(n5549), .A2(n7709), .ZN(n6085) );
  OAI211_X1 U7820 ( .C1(n5580), .C2(n9917), .A(n6086), .B(n6085), .ZN(n7712)
         );
  NAND2_X1 U7821 ( .A1(n4257), .A2(n7712), .ZN(n6087) );
  OAI21_X1 U7822 ( .B1(n4257), .B2(n6088), .A(n6087), .ZN(P1_U3586) );
  INV_X1 U7823 ( .A(n6298), .ZN(n6217) );
  NAND2_X1 U7824 ( .A1(n4257), .A2(n6217), .ZN(n6089) );
  OAI21_X1 U7825 ( .B1(n4257), .B2(n4792), .A(n6089), .ZN(P1_U3555) );
  NAND2_X1 U7826 ( .A1(n9190), .A2(n4257), .ZN(n6090) );
  OAI21_X1 U7827 ( .B1(n5274), .B2(n4257), .A(n6090), .ZN(P1_U3577) );
  INV_X1 U7828 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n6102) );
  INV_X1 U7829 ( .A(n9526), .ZN(n9628) );
  AOI211_X1 U7830 ( .C1(n6093), .C2(n6092), .A(n6091), .B(n9628), .ZN(n6098)
         );
  AOI211_X1 U7831 ( .C1(n6096), .C2(n6095), .A(n6094), .B(n9640), .ZN(n6097)
         );
  NOR2_X1 U7832 ( .A1(n6098), .A2(n6097), .ZN(n6101) );
  INV_X1 U7833 ( .A(n9523), .ZN(n9634) );
  AND2_X1 U7834 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6202) );
  AOI21_X1 U7835 ( .B1(n9634), .B2(n6099), .A(n6202), .ZN(n6100) );
  OAI211_X1 U7836 ( .C1(n6102), .C2(n9643), .A(n6101), .B(n6100), .ZN(P1_U3244) );
  INV_X1 U7837 ( .A(n6551), .ZN(n8388) );
  OAI222_X1 U7838 ( .A1(n8388), .A2(P2_U3152), .B1(n7319), .B2(n6104), .C1(
        n6103), .C2(n7947), .ZN(P2_U3346) );
  INV_X1 U7839 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6117) );
  OAI21_X1 U7840 ( .B1(n6107), .B2(n6106), .A(n6105), .ZN(n6112) );
  AOI211_X1 U7841 ( .C1(n6110), .C2(n6109), .A(n6108), .B(n9628), .ZN(n6111)
         );
  AOI21_X1 U7842 ( .B1(n9622), .B2(n6112), .A(n6111), .ZN(n6116) );
  INV_X1 U7843 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n6113) );
  NOR2_X1 U7844 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6113), .ZN(n8971) );
  AOI21_X1 U7845 ( .B1(n9634), .B2(n6114), .A(n8971), .ZN(n6115) );
  OAI211_X1 U7846 ( .C1(n6117), .C2(n9643), .A(n6116), .B(n6115), .ZN(P1_U3247) );
  NOR2_X1 U7847 ( .A1(n9376), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7848 ( .A(n6287), .ZN(n6121) );
  NOR2_X1 U7849 ( .A1(n6298), .A2(n6289), .ZN(n7668) );
  NOR2_X1 U7850 ( .A1(n7668), .A2(n6296), .ZN(n7434) );
  OR2_X1 U7851 ( .A1(n6177), .A2(n6176), .ZN(n7409) );
  NAND2_X1 U7852 ( .A1(n7409), .A2(n6287), .ZN(n6118) );
  OR2_X1 U7853 ( .A1(n7434), .A2(n6118), .ZN(n6120) );
  OR2_X1 U7854 ( .A1(n7665), .A2(n9210), .ZN(n6119) );
  NAND2_X1 U7855 ( .A1(n6120), .A2(n6119), .ZN(n6291) );
  AOI21_X1 U7856 ( .B1(n6289), .B2(n6121), .A(n6291), .ZN(n6133) );
  NAND2_X1 U7857 ( .A1(n9729), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6122) );
  OAI21_X1 U7858 ( .B1(n6133), .B2(n9729), .A(n6122), .ZN(P1_U3523) );
  INV_X1 U7859 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6127) );
  INV_X1 U7860 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n6125) );
  NAND2_X1 U7861 ( .A1(n4814), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6124) );
  NAND2_X1 U7862 ( .A1(n4816), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6123) );
  OAI211_X1 U7863 ( .C1(n7899), .C2(n6125), .A(n6124), .B(n6123), .ZN(n8462)
         );
  NAND2_X1 U7864 ( .A1(P2_U3966), .A2(n8462), .ZN(n6126) );
  OAI21_X1 U7865 ( .B1(P2_U3966), .B2(n6127), .A(n6126), .ZN(P2_U3583) );
  INV_X1 U7866 ( .A(n6128), .ZN(n6138) );
  OAI222_X1 U7867 ( .A1(n7850), .A2(n6138), .B1(n6852), .B2(P1_U3084), .C1(
        n6129), .C2(n4258), .ZN(P1_U3340) );
  INV_X1 U7868 ( .A(n6130), .ZN(n6131) );
  NOR2_X1 U7869 ( .A1(n9373), .A2(n6131), .ZN(n6284) );
  AND2_X2 U7870 ( .A1(n6132), .A2(n6284), .ZN(n9722) );
  OR2_X1 U7871 ( .A1(n6133), .A2(n9720), .ZN(n6134) );
  OAI21_X1 U7872 ( .B1(n9722), .B2(n5526), .A(n6134), .ZN(P1_U3454) );
  INV_X1 U7873 ( .A(n6135), .ZN(n6164) );
  AOI22_X1 U7874 ( .A1(n6854), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n6426), .ZN(n6136) );
  OAI21_X1 U7875 ( .B1(n6164), .B2(n7850), .A(n6136), .ZN(P1_U3339) );
  INV_X1 U7876 ( .A(n6665), .ZN(n6660) );
  OAI222_X1 U7877 ( .A1(P2_U3152), .A2(n6660), .B1(n7319), .B2(n6138), .C1(
        n6137), .C2(n7947), .ZN(P2_U3345) );
  OAI22_X1 U7878 ( .A1(n9523), .A2(n6139), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n6246), .ZN(n6149) );
  XNOR2_X1 U7879 ( .A(n6141), .B(n6140), .ZN(n6147) );
  INV_X1 U7880 ( .A(n6142), .ZN(n6143) );
  OAI211_X1 U7881 ( .C1(n6145), .C2(n6144), .A(n9526), .B(n6143), .ZN(n6146)
         );
  OAI21_X1 U7882 ( .B1(n6147), .B2(n9640), .A(n6146), .ZN(n6148) );
  AOI211_X1 U7883 ( .C1(n9012), .C2(P1_ADDR_REG_2__SCAN_IN), .A(n6149), .B(
        n6148), .ZN(n6162) );
  INV_X1 U7884 ( .A(n6151), .ZN(n6153) );
  AOI22_X1 U7885 ( .A1(n6474), .A2(n6289), .B1(n6153), .B2(
        P1_IR_REG_0__SCAN_IN), .ZN(n6152) );
  OR2_X1 U7886 ( .A1(n6613), .A2(n6305), .ZN(n6155) );
  NAND2_X1 U7887 ( .A1(n6153), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6154) );
  OAI21_X1 U7888 ( .B1(n6156), .B2(n6157), .A(n6180), .ZN(n6172) );
  MUX2_X1 U7889 ( .A(n6158), .B(n6172), .S(n6046), .Z(n6161) );
  OAI211_X1 U7890 ( .C1(n6161), .C2(n5916), .A(n6160), .B(n6159), .ZN(n9036)
         );
  NAND2_X1 U7891 ( .A1(n6162), .A2(n9036), .ZN(P1_U3243) );
  INV_X1 U7892 ( .A(n6997), .ZN(n7001) );
  OAI222_X1 U7893 ( .A1(P2_U3152), .A2(n7001), .B1(n7319), .B2(n6164), .C1(
        n6163), .C2(n7947), .ZN(P2_U3344) );
  NAND2_X1 U7894 ( .A1(n6165), .A2(n6281), .ZN(n6206) );
  OR2_X1 U7895 ( .A1(n6287), .A2(n6565), .ZN(n9472) );
  AND2_X1 U7896 ( .A1(n7409), .A2(n9472), .ZN(n6166) );
  NOR2_X1 U7897 ( .A1(n9372), .A2(n6166), .ZN(n6167) );
  NAND2_X1 U7898 ( .A1(n6206), .A2(n6167), .ZN(n6208) );
  AND2_X1 U7899 ( .A1(n6208), .A2(n6282), .ZN(n6173) );
  INV_X1 U7900 ( .A(n6173), .ZN(n8889) );
  AOI21_X1 U7901 ( .B1(n6206), .B2(n9713), .A(n8889), .ZN(n6247) );
  OR2_X1 U7902 ( .A1(n9372), .A2(n7409), .ZN(n6168) );
  NOR2_X1 U7903 ( .A1(n6206), .A2(n6168), .ZN(n6200) );
  INV_X1 U7904 ( .A(n7665), .ZN(n9008) );
  INV_X1 U7905 ( .A(n6206), .ZN(n6171) );
  AND2_X1 U7906 ( .A1(n9713), .A2(n7654), .ZN(n6205) );
  INV_X1 U7907 ( .A(n6205), .ZN(n6169) );
  NOR2_X1 U7908 ( .A1(n9372), .A2(n6169), .ZN(n6170) );
  NAND2_X1 U7909 ( .A1(n6171), .A2(n6170), .ZN(n8993) );
  AOI22_X1 U7910 ( .A1(n8986), .A2(n9008), .B1(n6172), .B2(n8969), .ZN(n6175)
         );
  NAND2_X1 U7911 ( .A1(n8991), .A2(n6289), .ZN(n6174) );
  OAI211_X1 U7912 ( .C1(n6247), .C2(n6290), .A(n6175), .B(n6174), .ZN(P1_U3230) );
  NAND2_X1 U7913 ( .A1(n6178), .A2(n7821), .ZN(n6179) );
  NAND2_X1 U7914 ( .A1(n6180), .A2(n6179), .ZN(n6214) );
  OR2_X1 U7915 ( .A1(n6613), .A2(n9683), .ZN(n6181) );
  OAI21_X1 U7916 ( .B1(n6195), .B2(n7665), .A(n6181), .ZN(n6182) );
  XNOR2_X1 U7917 ( .A(n6182), .B(n7821), .ZN(n6185) );
  OAI22_X1 U7918 ( .A1(n7814), .A2(n7665), .B1(n9683), .B2(n6195), .ZN(n6184)
         );
  NAND2_X1 U7919 ( .A1(n6185), .A2(n6184), .ZN(n6183) );
  NAND2_X1 U7920 ( .A1(n6214), .A2(n6183), .ZN(n6187) );
  INV_X1 U7921 ( .A(n6184), .ZN(n6213) );
  INV_X1 U7922 ( .A(n6185), .ZN(n6216) );
  NAND2_X1 U7923 ( .A1(n6213), .A2(n6216), .ZN(n6186) );
  NAND2_X1 U7924 ( .A1(n6187), .A2(n6186), .ZN(n6243) );
  OR2_X1 U7925 ( .A1(n6195), .A2(n7669), .ZN(n6188) );
  OAI21_X1 U7926 ( .B1(n6613), .B2(n6676), .A(n6188), .ZN(n6189) );
  INV_X1 U7927 ( .A(n7821), .ZN(n6197) );
  XNOR2_X1 U7928 ( .A(n6189), .B(n6197), .ZN(n6191) );
  OAI22_X1 U7929 ( .A1(n7814), .A2(n7669), .B1(n6676), .B2(n6195), .ZN(n6190)
         );
  XNOR2_X1 U7930 ( .A(n6191), .B(n6190), .ZN(n6244) );
  NAND2_X1 U7931 ( .A1(n6243), .A2(n6244), .ZN(n6194) );
  INV_X1 U7932 ( .A(n6190), .ZN(n6192) );
  NAND2_X1 U7933 ( .A1(n6192), .A2(n6191), .ZN(n6193) );
  NAND2_X1 U7934 ( .A1(n6194), .A2(n6193), .ZN(n6467) );
  OR2_X1 U7935 ( .A1(n6195), .A2(n6432), .ZN(n6196) );
  OAI21_X1 U7936 ( .B1(n6613), .B2(n6496), .A(n6196), .ZN(n6198) );
  OAI22_X1 U7937 ( .A1(n7814), .A2(n6432), .B1(n6496), .B2(n6195), .ZN(n6468)
         );
  XNOR2_X1 U7938 ( .A(n6469), .B(n6468), .ZN(n6466) );
  XOR2_X1 U7939 ( .A(n6467), .B(n6466), .Z(n6212) );
  INV_X1 U7940 ( .A(n8985), .ZN(n8898) );
  NOR2_X1 U7941 ( .A1(n8898), .A2(n7669), .ZN(n6201) );
  AOI211_X1 U7942 ( .C1(n8986), .C2(n9005), .A(n6202), .B(n6201), .ZN(n6211)
         );
  NAND3_X1 U7943 ( .A1(n6151), .A2(n6590), .A3(n6203), .ZN(n6204) );
  AOI21_X1 U7944 ( .B1(n6206), .B2(n6205), .A(n6204), .ZN(n6207) );
  OR2_X1 U7945 ( .A1(n6207), .A2(P1_U3084), .ZN(n6209) );
  INV_X1 U7946 ( .A(n8989), .ZN(n8975) );
  AOI22_X1 U7947 ( .A1(n8975), .A2(n5550), .B1(n8991), .B2(n6275), .ZN(n6210)
         );
  OAI211_X1 U7948 ( .C1(n8993), .C2(n6212), .A(n6211), .B(n6210), .ZN(P1_U3216) );
  XNOR2_X1 U7949 ( .A(n6214), .B(n6213), .ZN(n6215) );
  XNOR2_X1 U7950 ( .A(n6216), .B(n6215), .ZN(n6221) );
  INV_X1 U7951 ( .A(n7669), .ZN(n9007) );
  AOI22_X1 U7952 ( .A1(n8986), .A2(n9007), .B1(n8985), .B2(n6217), .ZN(n6218)
         );
  OAI21_X1 U7953 ( .B1(n6247), .B2(n9009), .A(n6218), .ZN(n6219) );
  AOI21_X1 U7954 ( .B1(n8991), .B2(n7664), .A(n6219), .ZN(n6220) );
  OAI21_X1 U7955 ( .B1(n8993), .B2(n6221), .A(n6220), .ZN(P1_U3220) );
  MUX2_X1 U7956 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6222), .S(n6234), .Z(n9529)
         );
  NAND2_X1 U7957 ( .A1(n9529), .A2(n9530), .ZN(n9528) );
  OAI21_X1 U7958 ( .B1(n9522), .B2(n6222), .A(n9528), .ZN(n9542) );
  MUX2_X1 U7959 ( .A(n6224), .B(P1_REG1_REG_9__SCAN_IN), .S(n9539), .Z(n9541)
         );
  AOI21_X1 U7960 ( .B1(n6225), .B2(n6224), .A(n9540), .ZN(n9554) );
  MUX2_X1 U7961 ( .A(n6226), .B(P1_REG1_REG_10__SCAN_IN), .S(n9551), .Z(n9553)
         );
  AOI22_X1 U7962 ( .A1(n6847), .A2(n5661), .B1(P1_REG1_REG_11__SCAN_IN), .B2(
        n6839), .ZN(n6228) );
  AOI21_X1 U7963 ( .B1(n6229), .B2(n6228), .A(n6838), .ZN(n6242) );
  AND2_X1 U7964 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7047) );
  NOR2_X1 U7965 ( .A1(n9523), .A2(n6839), .ZN(n6230) );
  AOI211_X1 U7966 ( .C1(n9012), .C2(P1_ADDR_REG_11__SCAN_IN), .A(n7047), .B(
        n6230), .ZN(n6241) );
  MUX2_X1 U7967 ( .A(n5623), .B(P1_REG2_REG_8__SCAN_IN), .S(n6234), .Z(n6231)
         );
  INV_X1 U7968 ( .A(n6231), .ZN(n9520) );
  NAND2_X1 U7969 ( .A1(n9539), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6235) );
  OAI21_X1 U7970 ( .B1(n9539), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6235), .ZN(
        n9535) );
  NOR2_X1 U7971 ( .A1(n9536), .A2(n9535), .ZN(n9534) );
  XNOR2_X1 U7972 ( .A(n9551), .B(P1_REG2_REG_10__SCAN_IN), .ZN(n9547) );
  NOR2_X1 U7973 ( .A1(n6847), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n6236) );
  AOI21_X1 U7974 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n6847), .A(n6236), .ZN(
        n6237) );
  OAI21_X1 U7975 ( .B1(n6238), .B2(n6237), .A(n6846), .ZN(n6239) );
  NAND2_X1 U7976 ( .A1(n9526), .A2(n6239), .ZN(n6240) );
  OAI211_X1 U7977 ( .C1(n6242), .C2(n9640), .A(n6241), .B(n6240), .ZN(P1_U3252) );
  XOR2_X1 U7978 ( .A(n6244), .B(n6243), .Z(n6250) );
  INV_X1 U7979 ( .A(n6432), .ZN(n9006) );
  AOI22_X1 U7980 ( .A1(n8985), .A2(n9008), .B1(n8986), .B2(n9006), .ZN(n6245)
         );
  OAI21_X1 U7981 ( .B1(n6247), .B2(n6246), .A(n6245), .ZN(n6248) );
  AOI21_X1 U7982 ( .B1(n8991), .B2(n5547), .A(n6248), .ZN(n6249) );
  OAI21_X1 U7983 ( .B1(n8993), .B2(n6250), .A(n6249), .ZN(P1_U3235) );
  OAI21_X1 U7984 ( .B1(n4251), .B2(n6252), .A(n6251), .ZN(n6678) );
  INV_X1 U7985 ( .A(n6274), .ZN(n6253) );
  AOI21_X1 U7986 ( .B1(n5547), .B2(n6304), .A(n6253), .ZN(n6673) );
  INV_X1 U7987 ( .A(n6673), .ZN(n6254) );
  OAI22_X1 U7988 ( .A1(n6254), .A2(n9714), .B1(n6676), .B2(n9713), .ZN(n6258)
         );
  XNOR2_X1 U7989 ( .A(n7431), .B(n6255), .ZN(n6256) );
  AOI222_X1 U7990 ( .A1(n9651), .A2(n6256), .B1(n9006), .B2(n9656), .C1(n9008), 
        .C2(n9654), .ZN(n6680) );
  INV_X1 U7991 ( .A(n6680), .ZN(n6257) );
  AOI211_X1 U7992 ( .C1(n9718), .C2(n6678), .A(n6258), .B(n6257), .ZN(n9687)
         );
  NAND2_X1 U7993 ( .A1(n9729), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6259) );
  OAI21_X1 U7994 ( .B1(n9687), .B2(n9729), .A(n6259), .ZN(P1_U3525) );
  INV_X1 U7995 ( .A(n6260), .ZN(n6262) );
  INV_X1 U7996 ( .A(n9596), .ZN(n9047) );
  OAI222_X1 U7997 ( .A1(n4258), .A2(n6261), .B1(n7850), .B2(n6262), .C1(
        P1_U3084), .C2(n9047), .ZN(P1_U3338) );
  INV_X1 U7998 ( .A(n8406), .ZN(n8395) );
  OAI222_X1 U7999 ( .A1(n7947), .A2(n6263), .B1(n7319), .B2(n6262), .C1(n8395), 
        .C2(P2_U3152), .ZN(P2_U3343) );
  INV_X1 U8000 ( .A(n6264), .ZN(n6267) );
  AOI22_X1 U8001 ( .A1(n9607), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n6426), .ZN(n6265) );
  OAI21_X1 U8002 ( .B1(n6267), .B2(n7850), .A(n6265), .ZN(P1_U3337) );
  AOI22_X1 U8003 ( .A1(n8418), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n7399), .ZN(n6266) );
  OAI21_X1 U8004 ( .B1(n6267), .B2(n7319), .A(n6266), .ZN(P2_U3342) );
  OAI21_X1 U8005 ( .B1(n6269), .B2(n6270), .A(n6268), .ZN(n6498) );
  INV_X1 U8006 ( .A(n6498), .ZN(n6277) );
  INV_X1 U8007 ( .A(n6457), .ZN(n9659) );
  OAI22_X1 U8008 ( .A1(n7669), .A2(n9212), .B1(n6486), .B2(n9210), .ZN(n6273)
         );
  XNOR2_X1 U8009 ( .A(n7487), .B(n6270), .ZN(n6271) );
  INV_X1 U8010 ( .A(n9651), .ZN(n9207) );
  NOR2_X1 U8011 ( .A1(n6271), .A2(n9207), .ZN(n6272) );
  AOI211_X1 U8012 ( .C1(n9659), .C2(n6498), .A(n6273), .B(n6272), .ZN(n6500)
         );
  AOI21_X1 U8013 ( .B1(n6275), .B2(n6274), .A(n6437), .ZN(n6493) );
  INV_X1 U8014 ( .A(n9714), .ZN(n9469) );
  AOI22_X1 U8015 ( .A1(n6493), .A2(n9469), .B1(n9345), .B2(n6275), .ZN(n6276)
         );
  OAI211_X1 U8016 ( .C1(n6277), .C2(n9389), .A(n6500), .B(n6276), .ZN(n6279)
         );
  NAND2_X1 U8017 ( .A1(n6279), .A2(n9731), .ZN(n6278) );
  OAI21_X1 U8018 ( .B1(n9731), .B2(n5551), .A(n6278), .ZN(P1_U3526) );
  NAND2_X1 U8019 ( .A1(n6279), .A2(n9722), .ZN(n6280) );
  OAI21_X1 U8020 ( .B1(n9722), .B2(n5552), .A(n6280), .ZN(P1_U3463) );
  INV_X1 U8021 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n6295) );
  AND2_X1 U8022 ( .A1(n6282), .A2(n6281), .ZN(n6283) );
  NAND2_X1 U8023 ( .A1(n6284), .A2(n6283), .ZN(n6509) );
  INV_X1 U8024 ( .A(n6286), .ZN(n7697) );
  OR2_X1 U8025 ( .A1(n6287), .A2(n7697), .ZN(n6288) );
  OR2_X1 U8026 ( .A1(n9676), .A2(n6288), .ZN(n9671) );
  INV_X1 U8027 ( .A(n9671), .ZN(n9277) );
  OAI21_X1 U8028 ( .B1(n9669), .B2(n9277), .A(n6289), .ZN(n6294) );
  NOR2_X1 U8029 ( .A1(n9663), .A2(n6290), .ZN(n6292) );
  OAI21_X1 U8030 ( .B1(n6292), .B2(n6291), .A(n9666), .ZN(n6293) );
  OAI211_X1 U8031 ( .C1(n6295), .C2(n9666), .A(n6294), .B(n6293), .ZN(P1_U3291) );
  XNOR2_X1 U8032 ( .A(n6302), .B(n6296), .ZN(n6297) );
  OAI222_X1 U8033 ( .A1(n9212), .A2(n6298), .B1(n9210), .B2(n7669), .C1(n6297), 
        .C2(n9207), .ZN(n9684) );
  NAND2_X1 U8034 ( .A1(n6299), .A2(n9473), .ZN(n6430) );
  OR2_X1 U8035 ( .A1(n6302), .A2(n6301), .ZN(n6303) );
  NAND2_X1 U8036 ( .A1(n6300), .A2(n6303), .ZN(n9681) );
  AOI21_X1 U8037 ( .B1(n6457), .B2(n6430), .A(n9681), .ZN(n6307) );
  OAI211_X1 U8038 ( .C1(n9683), .C2(n6305), .A(n9469), .B(n6304), .ZN(n9682)
         );
  OAI22_X1 U8039 ( .A1(n9663), .A2(n9009), .B1(n9473), .B2(n9682), .ZN(n6306)
         );
  NOR3_X1 U8040 ( .A1(n9684), .A2(n6307), .A3(n6306), .ZN(n6309) );
  AOI22_X1 U8041 ( .A1(n9669), .A2(n7664), .B1(n9676), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n6308) );
  OAI21_X1 U8042 ( .B1(n9676), .B2(n6309), .A(n6308), .ZN(P1_U3290) );
  INV_X1 U8043 ( .A(n7528), .ZN(n6315) );
  NAND2_X1 U8044 ( .A1(n6310), .A2(n6311), .ZN(n6314) );
  INV_X1 U8045 ( .A(n6312), .ZN(n6313) );
  AOI21_X1 U8046 ( .B1(n6315), .B2(n6314), .A(n6313), .ZN(n9697) );
  INV_X1 U8047 ( .A(n9697), .ZN(n6324) );
  NAND2_X1 U8048 ( .A1(n7409), .A2(n7821), .ZN(n9466) );
  AOI22_X1 U8049 ( .A1(n9669), .A2(n6488), .B1(n9676), .B2(
        P1_REG2_REG_5__SCAN_IN), .ZN(n6323) );
  XNOR2_X1 U8050 ( .A(n6452), .B(n7528), .ZN(n6316) );
  NAND2_X1 U8051 ( .A1(n6316), .A2(n9651), .ZN(n6318) );
  AOI22_X1 U8052 ( .A1(n9656), .A2(n9003), .B1(n9654), .B2(n9005), .ZN(n6317)
         );
  NAND2_X1 U8053 ( .A1(n6318), .A2(n6317), .ZN(n9696) );
  INV_X1 U8054 ( .A(n6439), .ZN(n6319) );
  OAI211_X1 U8055 ( .C1(n6319), .C2(n9694), .A(n9469), .B(n6458), .ZN(n9693)
         );
  INV_X1 U8056 ( .A(n6489), .ZN(n6320) );
  OAI22_X1 U8057 ( .A1(n9693), .A2(n9473), .B1(n9663), .B2(n6320), .ZN(n6321)
         );
  OAI21_X1 U8058 ( .B1(n9696), .B2(n6321), .A(n9666), .ZN(n6322) );
  OAI211_X1 U8059 ( .C1(n6324), .C2(n9279), .A(n6323), .B(n6322), .ZN(P1_U3286) );
  AND2_X1 U8060 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6334) );
  NAND2_X1 U8061 ( .A1(n6340), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6330) );
  MUX2_X1 U8062 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6325), .S(n6340), .Z(n8334)
         );
  INV_X1 U8063 ( .A(n6326), .ZN(n6327) );
  OAI21_X1 U8064 ( .B1(n9870), .B2(n6335), .A(n6327), .ZN(n9385) );
  MUX2_X1 U8065 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6328), .S(n9381), .Z(n9384)
         );
  NAND2_X1 U8066 ( .A1(n9385), .A2(n9384), .ZN(n9383) );
  NAND2_X1 U8067 ( .A1(n9381), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6329) );
  NAND2_X1 U8068 ( .A1(n9383), .A2(n6329), .ZN(n8333) );
  NAND2_X1 U8069 ( .A1(n8334), .A2(n8333), .ZN(n8332) );
  AND2_X1 U8070 ( .A1(n6330), .A2(n8332), .ZN(n6332) );
  MUX2_X1 U8071 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6347), .S(n6359), .Z(n6331)
         );
  NOR2_X1 U8072 ( .A1(n6332), .A2(n6331), .ZN(n6345) );
  AOI211_X1 U8073 ( .C1(n6332), .C2(n6331), .A(n6345), .B(n9740), .ZN(n6333)
         );
  AOI211_X1 U8074 ( .C1(n9376), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6334), .B(
        n6333), .ZN(n6342) );
  INV_X1 U8075 ( .A(n6335), .ZN(n6337) );
  NAND2_X1 U8076 ( .A1(n9381), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6338) );
  OAI21_X1 U8077 ( .B1(n9381), .B2(P2_REG2_REG_2__SCAN_IN), .A(n6338), .ZN(
        n9378) );
  NOR2_X1 U8078 ( .A1(n9379), .A2(n9378), .ZN(n9377) );
  NAND2_X1 U8079 ( .A1(n6340), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6339) );
  OAI21_X1 U8080 ( .B1(n6340), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6339), .ZN(
        n8330) );
  OAI211_X1 U8081 ( .C1(n4277), .C2(n4481), .A(n9733), .B(n6360), .ZN(n6341)
         );
  OAI211_X1 U8082 ( .C1(n9739), .C2(n6359), .A(n6342), .B(n6341), .ZN(P2_U3249) );
  NAND2_X1 U8083 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3152), .ZN(n6823) );
  INV_X1 U8084 ( .A(n6823), .ZN(n6358) );
  NAND2_X1 U8085 ( .A1(n8357), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6351) );
  MUX2_X1 U8086 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6343), .S(n8357), .Z(n8360)
         );
  NAND2_X1 U8087 ( .A1(n6363), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6348) );
  MUX2_X1 U8088 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6344), .S(n6363), .Z(n8346)
         );
  INV_X1 U8089 ( .A(n6345), .ZN(n6346) );
  OAI21_X1 U8090 ( .B1(n6359), .B2(n6347), .A(n6346), .ZN(n8345) );
  NAND2_X1 U8091 ( .A1(n8346), .A2(n8345), .ZN(n8344) );
  AND2_X1 U8092 ( .A1(n6348), .A2(n8344), .ZN(n6398) );
  MUX2_X1 U8093 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6350), .S(n6404), .Z(n6397)
         );
  NOR2_X1 U8094 ( .A1(n6398), .A2(n6397), .ZN(n6396) );
  INV_X1 U8095 ( .A(n6396), .ZN(n6349) );
  OAI21_X1 U8096 ( .B1(n6350), .B2(n6404), .A(n6349), .ZN(n8359) );
  NAND2_X1 U8097 ( .A1(n8360), .A2(n8359), .ZN(n8358) );
  NAND2_X1 U8098 ( .A1(n6351), .A2(n8358), .ZN(n6354) );
  INV_X1 U8099 ( .A(n6354), .ZN(n6356) );
  MUX2_X1 U8100 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6352), .S(n6389), .Z(n6355)
         );
  MUX2_X1 U8101 ( .A(n6352), .B(P2_REG1_REG_8__SCAN_IN), .S(n6389), .Z(n6353)
         );
  AOI211_X1 U8102 ( .C1(n6356), .C2(n6355), .A(n6382), .B(n9740), .ZN(n6357)
         );
  AOI211_X1 U8103 ( .C1(n9376), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n6358), .B(
        n6357), .ZN(n6374) );
  MUX2_X1 U8104 ( .A(n6390), .B(P2_REG2_REG_8__SCAN_IN), .S(n6389), .Z(n6372)
         );
  INV_X1 U8105 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6369) );
  INV_X1 U8106 ( .A(n6360), .ZN(n6361) );
  NAND2_X1 U8107 ( .A1(n6363), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6362) );
  OAI21_X1 U8108 ( .B1(n6363), .B2(P2_REG2_REG_5__SCAN_IN), .A(n6362), .ZN(
        n8342) );
  INV_X1 U8109 ( .A(n6404), .ZN(n6365) );
  NAND2_X1 U8110 ( .A1(n8357), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6367) );
  OAI21_X1 U8111 ( .B1(n8357), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6367), .ZN(
        n6368) );
  INV_X1 U8112 ( .A(n6368), .ZN(n8355) );
  OAI21_X1 U8113 ( .B1(n6370), .B2(n6369), .A(n8353), .ZN(n6371) );
  NAND2_X1 U8114 ( .A1(n6371), .A2(n6372), .ZN(n6388) );
  OAI211_X1 U8115 ( .C1(n6372), .C2(n6371), .A(n9733), .B(n6388), .ZN(n6373)
         );
  OAI211_X1 U8116 ( .C1(n9739), .C2(n6389), .A(n6374), .B(n6373), .ZN(P2_U3253) );
  INV_X1 U8117 ( .A(n6375), .ZN(n6385) );
  INV_X1 U8118 ( .A(n6382), .ZN(n6378) );
  INV_X1 U8119 ( .A(n6389), .ZN(n6376) );
  NAND2_X1 U8120 ( .A1(n6376), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6379) );
  INV_X1 U8121 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n9879) );
  MUX2_X1 U8122 ( .A(n9879), .B(P2_REG1_REG_9__SCAN_IN), .S(n6406), .Z(n6377)
         );
  AOI21_X1 U8123 ( .B1(n6378), .B2(n6379), .A(n6377), .ZN(n6411) );
  INV_X1 U8124 ( .A(n6379), .ZN(n6381) );
  MUX2_X1 U8125 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n9879), .S(n6406), .Z(n6380)
         );
  NOR3_X1 U8126 ( .A1(n6382), .A2(n6381), .A3(n6380), .ZN(n6383) );
  NOR3_X1 U8127 ( .A1(n9740), .A2(n6411), .A3(n6383), .ZN(n6384) );
  AOI211_X1 U8128 ( .C1(n9376), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n6385), .B(
        n6384), .ZN(n6394) );
  NAND2_X1 U8129 ( .A1(n6406), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6386) );
  OAI21_X1 U8130 ( .B1(n6406), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6386), .ZN(
        n6387) );
  INV_X1 U8131 ( .A(n6387), .ZN(n6392) );
  OAI21_X1 U8132 ( .B1(n6390), .B2(n6389), .A(n6388), .ZN(n6391) );
  NAND2_X1 U8133 ( .A1(n6391), .A2(n6392), .ZN(n6418) );
  OAI211_X1 U8134 ( .C1(n6392), .C2(n6391), .A(n9733), .B(n6418), .ZN(n6393)
         );
  OAI211_X1 U8135 ( .C1(n9739), .C2(n6419), .A(n6394), .B(n6393), .ZN(P2_U3254) );
  NOR2_X1 U8136 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6395), .ZN(n6400) );
  AOI211_X1 U8137 ( .C1(n6398), .C2(n6397), .A(n6396), .B(n9740), .ZN(n6399)
         );
  AOI211_X1 U8138 ( .C1(n9376), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n6400), .B(
        n6399), .ZN(n6403) );
  OAI211_X1 U8139 ( .C1(n4320), .C2(n4478), .A(n9733), .B(n6401), .ZN(n6402)
         );
  OAI211_X1 U8140 ( .C1(n9739), .C2(n6404), .A(n6403), .B(n6402), .ZN(P2_U3251) );
  NOR2_X1 U8141 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6405), .ZN(n6417) );
  INV_X1 U8142 ( .A(n9740), .ZN(n9732) );
  NAND2_X1 U8143 ( .A1(n6406), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n6413) );
  INV_X1 U8144 ( .A(n6413), .ZN(n6407) );
  OR2_X1 U8145 ( .A1(n6411), .A2(n6407), .ZN(n6410) );
  INV_X1 U8146 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6408) );
  MUX2_X1 U8147 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6408), .S(n6549), .Z(n6409)
         );
  NAND2_X1 U8148 ( .A1(n6410), .A2(n6409), .ZN(n8373) );
  INV_X1 U8149 ( .A(n6411), .ZN(n6414) );
  MUX2_X1 U8150 ( .A(n6408), .B(P2_REG1_REG_10__SCAN_IN), .S(n6549), .Z(n6412)
         );
  NAND3_X1 U8151 ( .A1(n6414), .A2(n6413), .A3(n6412), .ZN(n6415) );
  AND3_X1 U8152 ( .A1(n9732), .A2(n8373), .A3(n6415), .ZN(n6416) );
  AOI211_X1 U8153 ( .C1(n9376), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n6417), .B(
        n6416), .ZN(n6423) );
  XOR2_X1 U8154 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n6549), .Z(n6421) );
  OAI21_X1 U8155 ( .B1(n6964), .B2(n6419), .A(n6418), .ZN(n6420) );
  NAND2_X1 U8156 ( .A1(n6420), .A2(n6421), .ZN(n6548) );
  OAI211_X1 U8157 ( .C1(n6421), .C2(n6420), .A(n9733), .B(n6548), .ZN(n6422)
         );
  OAI211_X1 U8158 ( .C1(n9739), .C2(n6424), .A(n6423), .B(n6422), .ZN(P2_U3255) );
  INV_X1 U8159 ( .A(n6425), .ZN(n6447) );
  AOI22_X1 U8160 ( .A1(n9620), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n6426), .ZN(n6427) );
  OAI21_X1 U8161 ( .B1(n6447), .B2(n7850), .A(n6427), .ZN(P1_U3336) );
  OR2_X1 U8162 ( .A1(n6428), .A2(n7435), .ZN(n6429) );
  NAND2_X1 U8163 ( .A1(n6310), .A2(n6429), .ZN(n9692) );
  INV_X1 U8164 ( .A(n9692), .ZN(n6445) );
  OR2_X1 U8165 ( .A1(n9676), .A2(n6430), .ZN(n7246) );
  XNOR2_X1 U8166 ( .A(n7435), .B(n7526), .ZN(n6436) );
  NOR2_X1 U8167 ( .A1(n6432), .A2(n9212), .ZN(n6434) );
  NOR2_X1 U8168 ( .A1(n8922), .A2(n9210), .ZN(n6433) );
  AOI211_X1 U8169 ( .C1(n9692), .C2(n9659), .A(n6434), .B(n6433), .ZN(n6435)
         );
  OAI21_X1 U8170 ( .B1(n9207), .B2(n6436), .A(n6435), .ZN(n9690) );
  NAND2_X1 U8171 ( .A1(n9690), .A2(n9666), .ZN(n6444) );
  OR2_X1 U8172 ( .A1(n6437), .A2(n9688), .ZN(n6438) );
  NAND2_X1 U8173 ( .A1(n6439), .A2(n6438), .ZN(n9689) );
  NOR2_X1 U8174 ( .A1(n9671), .A2(n9689), .ZN(n6442) );
  OAI22_X1 U8175 ( .A1(n9666), .A2(n6440), .B1(n8919), .B2(n9663), .ZN(n6441)
         );
  AOI211_X1 U8176 ( .C1(n9669), .C2(n8920), .A(n6442), .B(n6441), .ZN(n6443)
         );
  OAI211_X1 U8177 ( .C1(n6445), .C2(n7246), .A(n6444), .B(n6443), .ZN(P1_U3287) );
  INV_X1 U8178 ( .A(n8434), .ZN(n8430) );
  OAI222_X1 U8179 ( .A1(P2_U3152), .A2(n8430), .B1(n7319), .B2(n6447), .C1(
        n6446), .C2(n7947), .ZN(P2_U3341) );
  INV_X1 U8180 ( .A(n6449), .ZN(n6450) );
  AOI21_X1 U8181 ( .B1(n7540), .B2(n6451), .A(n6450), .ZN(n9698) );
  INV_X1 U8182 ( .A(n7535), .ZN(n7484) );
  OAI21_X1 U8183 ( .B1(n6452), .B2(n7484), .A(n7534), .ZN(n6453) );
  XNOR2_X1 U8184 ( .A(n6453), .B(n7540), .ZN(n6455) );
  OAI22_X1 U8185 ( .A1(n8922), .A2(n9212), .B1(n6609), .B2(n9210), .ZN(n6454)
         );
  AOI21_X1 U8186 ( .B1(n6455), .B2(n9651), .A(n6454), .ZN(n6456) );
  OAI21_X1 U8187 ( .B1(n9698), .B2(n6457), .A(n6456), .ZN(n9701) );
  NAND2_X1 U8188 ( .A1(n9701), .A2(n9666), .ZN(n6465) );
  INV_X1 U8189 ( .A(n6458), .ZN(n6460) );
  INV_X1 U8190 ( .A(n6459), .ZN(n6508) );
  OAI21_X1 U8191 ( .B1(n9699), .B2(n6460), .A(n6508), .ZN(n9700) );
  NOR2_X1 U8192 ( .A1(n9671), .A2(n9700), .ZN(n6463) );
  INV_X1 U8193 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6461) );
  OAI22_X1 U8194 ( .A1(n9666), .A2(n6461), .B1(n8972), .B2(n9663), .ZN(n6462)
         );
  AOI211_X1 U8195 ( .C1(n9669), .C2(n8973), .A(n6463), .B(n6462), .ZN(n6464)
         );
  OAI211_X1 U8196 ( .C1(n9698), .C2(n7246), .A(n6465), .B(n6464), .ZN(P1_U3285) );
  OAI22_X1 U8197 ( .A1(n7814), .A2(n8922), .B1(n9694), .B2(n6195), .ZN(n6610)
         );
  NAND2_X1 U8198 ( .A1(n6467), .A2(n6466), .ZN(n6472) );
  INV_X1 U8199 ( .A(n6468), .ZN(n6470) );
  NAND2_X1 U8200 ( .A1(n6470), .A2(n6469), .ZN(n6471) );
  NAND2_X1 U8201 ( .A1(n6472), .A2(n6471), .ZN(n8917) );
  NOR2_X1 U8202 ( .A1(n6195), .A2(n9688), .ZN(n6473) );
  AOI21_X1 U8203 ( .B1(n7820), .B2(n9005), .A(n6473), .ZN(n8914) );
  OR2_X1 U8204 ( .A1(n6195), .A2(n6486), .ZN(n6475) );
  OAI21_X1 U8205 ( .B1(n6613), .B2(n9688), .A(n6475), .ZN(n6476) );
  XNOR2_X1 U8206 ( .A(n6476), .B(n7806), .ZN(n6477) );
  AND2_X1 U8207 ( .A1(n8914), .A2(n6477), .ZN(n6480) );
  INV_X1 U8208 ( .A(n6477), .ZN(n8915) );
  INV_X1 U8209 ( .A(n8914), .ZN(n6478) );
  NAND2_X1 U8210 ( .A1(n8915), .A2(n6478), .ZN(n6479) );
  OR2_X1 U8211 ( .A1(n6195), .A2(n8922), .ZN(n6481) );
  OAI21_X1 U8212 ( .B1(n6613), .B2(n9694), .A(n6481), .ZN(n6482) );
  XNOR2_X1 U8213 ( .A(n6482), .B(n7821), .ZN(n6611) );
  INV_X1 U8214 ( .A(n6611), .ZN(n6484) );
  OR2_X1 U8215 ( .A1(n6483), .A2(n6611), .ZN(n8962) );
  OAI21_X1 U8216 ( .B1(n6619), .B2(n6484), .A(n8962), .ZN(n6485) );
  NOR2_X1 U8217 ( .A1(n6485), .A2(n6610), .ZN(n8964) );
  AOI21_X1 U8218 ( .B1(n6610), .B2(n6485), .A(n8964), .ZN(n6492) );
  INV_X1 U8219 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n10030) );
  NOR2_X1 U8220 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n10030), .ZN(n9512) );
  NOR2_X1 U8221 ( .A1(n8898), .A2(n6486), .ZN(n6487) );
  AOI211_X1 U8222 ( .C1(n8986), .C2(n9003), .A(n9512), .B(n6487), .ZN(n6491)
         );
  AOI22_X1 U8223 ( .A1(n8975), .A2(n6489), .B1(n8991), .B2(n6488), .ZN(n6490)
         );
  OAI211_X1 U8224 ( .C1(n6492), .C2(n8993), .A(n6491), .B(n6490), .ZN(P1_U3225) );
  INV_X1 U8225 ( .A(n7246), .ZN(n9673) );
  NAND2_X1 U8226 ( .A1(n9277), .A2(n6493), .ZN(n6495) );
  AOI22_X1 U8227 ( .A1(n9676), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9484), .B2(
        n5550), .ZN(n6494) );
  OAI211_X1 U8228 ( .C1(n6496), .C2(n9268), .A(n6495), .B(n6494), .ZN(n6497)
         );
  AOI21_X1 U8229 ( .B1(n9673), .B2(n6498), .A(n6497), .ZN(n6499) );
  OAI21_X1 U8230 ( .B1(n6500), .B2(n9274), .A(n6499), .ZN(P1_U3288) );
  OAI21_X1 U8231 ( .B1(n6502), .B2(n7437), .A(n6501), .ZN(n6503) );
  INV_X1 U8232 ( .A(n6503), .ZN(n6738) );
  INV_X1 U8233 ( .A(n6504), .ZN(n6505) );
  AOI21_X1 U8234 ( .B1(n7437), .B2(n6506), .A(n6505), .ZN(n6507) );
  OAI222_X1 U8235 ( .A1(n9210), .A2(n6629), .B1(n9212), .B2(n6615), .C1(n9207), 
        .C2(n6507), .ZN(n6734) );
  NAND2_X1 U8236 ( .A1(n6734), .A2(n9666), .ZN(n6516) );
  AOI211_X1 U8237 ( .C1(n6736), .C2(n6508), .A(n9714), .B(n6530), .ZN(n6735)
         );
  OR2_X1 U8238 ( .A1(n6509), .A2(n9473), .ZN(n7355) );
  INV_X1 U8239 ( .A(n7355), .ZN(n6514) );
  NOR2_X1 U8240 ( .A1(n9268), .A2(n6510), .ZN(n6513) );
  OAI22_X1 U8241 ( .A1(n9666), .A2(n6511), .B1(n6604), .B2(n9663), .ZN(n6512)
         );
  AOI211_X1 U8242 ( .C1(n6735), .C2(n6514), .A(n6513), .B(n6512), .ZN(n6515)
         );
  OAI211_X1 U8243 ( .C1(n6738), .C2(n9279), .A(n6516), .B(n6515), .ZN(P1_U3284) );
  INV_X1 U8244 ( .A(n6517), .ZN(n6600) );
  OAI222_X1 U8245 ( .A1(n7850), .A2(n6600), .B1(n6519), .B2(P1_U3084), .C1(
        n6518), .C2(n4258), .ZN(P1_U3332) );
  OAI21_X1 U8246 ( .B1(n7439), .B2(n6520), .A(n9647), .ZN(n6521) );
  NAND2_X1 U8247 ( .A1(n6521), .A2(n9651), .ZN(n6525) );
  OR2_X1 U8248 ( .A1(n6609), .A2(n9212), .ZN(n6522) );
  OAI21_X1 U8249 ( .B1(n6809), .B2(n9210), .A(n6522), .ZN(n6523) );
  INV_X1 U8250 ( .A(n6523), .ZN(n6524) );
  NAND2_X1 U8251 ( .A1(n6525), .A2(n6524), .ZN(n9709) );
  INV_X1 U8252 ( .A(n9709), .ZN(n6537) );
  NAND2_X1 U8253 ( .A1(n6526), .A2(n7439), .ZN(n6527) );
  AND2_X1 U8254 ( .A1(n6528), .A2(n6527), .ZN(n9705) );
  INV_X1 U8255 ( .A(n9279), .ZN(n7360) );
  OR2_X1 U8256 ( .A1(n6530), .A2(n6529), .ZN(n6531) );
  NAND2_X1 U8257 ( .A1(n9660), .A2(n6531), .ZN(n9707) );
  NAND2_X1 U8258 ( .A1(n9669), .A2(n6636), .ZN(n6534) );
  INV_X1 U8259 ( .A(n6655), .ZN(n6532) );
  AOI22_X1 U8260 ( .A1(n9676), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n6532), .B2(
        n9484), .ZN(n6533) );
  OAI211_X1 U8261 ( .C1(n9707), .C2(n9671), .A(n6534), .B(n6533), .ZN(n6535)
         );
  AOI21_X1 U8262 ( .B1(n9705), .B2(n7360), .A(n6535), .ZN(n6536) );
  OAI21_X1 U8263 ( .B1(n9676), .B2(n6537), .A(n6536), .ZN(P1_U3283) );
  INV_X1 U8264 ( .A(n6538), .ZN(n6540) );
  OAI222_X1 U8265 ( .A1(n4764), .A2(P2_U3152), .B1(n7319), .B2(n6540), .C1(
        n6539), .C2(n7947), .ZN(P2_U3339) );
  OAI222_X1 U8266 ( .A1(n4258), .A2(n9918), .B1(n7850), .B2(n6540), .C1(
        P1_U3084), .C2(n9146), .ZN(P1_U3334) );
  INV_X1 U8267 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9882) );
  NAND2_X1 U8268 ( .A1(n6549), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n8372) );
  NAND2_X1 U8269 ( .A1(n8373), .A2(n8372), .ZN(n6542) );
  MUX2_X1 U8270 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n9882), .S(n8370), .Z(n6541)
         );
  NAND2_X1 U8271 ( .A1(n6542), .A2(n6541), .ZN(n8375) );
  OAI21_X1 U8272 ( .B1(n9882), .B2(n6543), .A(n8375), .ZN(n8381) );
  MUX2_X1 U8273 ( .A(n6544), .B(P2_REG1_REG_12__SCAN_IN), .S(n6551), .Z(n8380)
         );
  NOR2_X1 U8274 ( .A1(n8381), .A2(n8380), .ZN(n8379) );
  AOI21_X1 U8275 ( .B1(n8388), .B2(n6544), .A(n8379), .ZN(n6546) );
  AOI22_X1 U8276 ( .A1(n6665), .A2(n5018), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n6660), .ZN(n6545) );
  NOR2_X1 U8277 ( .A1(n6546), .A2(n6545), .ZN(n6659) );
  AOI21_X1 U8278 ( .B1(n6546), .B2(n6545), .A(n6659), .ZN(n6558) );
  NAND2_X1 U8279 ( .A1(n6551), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6547) );
  OAI21_X1 U8280 ( .B1(n6551), .B2(P2_REG2_REG_12__SCAN_IN), .A(n6547), .ZN(
        n8383) );
  NOR2_X1 U8281 ( .A1(n8370), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n6550) );
  AOI21_X1 U8282 ( .B1(n8370), .B2(P2_REG2_REG_11__SCAN_IN), .A(n6550), .ZN(
        n8366) );
  NOR2_X1 U8283 ( .A1(n8383), .A2(n8384), .ZN(n8382) );
  AOI22_X1 U8284 ( .A1(n6665), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7308), .B2(
        n6660), .ZN(n6552) );
  NAND2_X1 U8285 ( .A1(n6553), .A2(n6552), .ZN(n6664) );
  OAI21_X1 U8286 ( .B1(n6553), .B2(n6552), .A(n6664), .ZN(n6556) );
  AOI22_X1 U8287 ( .A1(n9376), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3152), .ZN(n6554) );
  OAI21_X1 U8288 ( .B1(n9739), .B2(n6660), .A(n6554), .ZN(n6555) );
  AOI21_X1 U8289 ( .B1(n6556), .B2(n9733), .A(n6555), .ZN(n6557) );
  OAI21_X1 U8290 ( .B1(n6558), .B2(n9740), .A(n6557), .ZN(P2_U3258) );
  INV_X1 U8291 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n6560) );
  INV_X1 U8292 ( .A(n6559), .ZN(n6562) );
  INV_X1 U8293 ( .A(n9635), .ZN(n9054) );
  OAI222_X1 U8294 ( .A1(n4258), .A2(n6560), .B1(n7850), .B2(n6562), .C1(
        P1_U3084), .C2(n9054), .ZN(P1_U3335) );
  INV_X1 U8295 ( .A(n8439), .ZN(n8448) );
  INV_X1 U8296 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n6561) );
  OAI222_X1 U8297 ( .A1(n8448), .A2(P2_U3152), .B1(n7319), .B2(n6562), .C1(
        n6561), .C2(n7947), .ZN(P2_U3340) );
  INV_X1 U8298 ( .A(n6563), .ZN(n6583) );
  OAI222_X1 U8299 ( .A1(n7850), .A2(n6583), .B1(n6565), .B2(P1_U3084), .C1(
        n6564), .C2(n4258), .ZN(P1_U3333) );
  NOR2_X1 U8300 ( .A1(n8079), .A2(P2_U3152), .ZN(n6598) );
  NAND2_X1 U8301 ( .A1(n8326), .A2(n8729), .ZN(n6567) );
  NAND2_X1 U8302 ( .A1(n6691), .A2(n8730), .ZN(n6566) );
  AND2_X1 U8303 ( .A1(n6567), .A2(n6566), .ZN(n6724) );
  NAND2_X1 U8304 ( .A1(n6569), .A2(n6568), .ZN(n7971) );
  OAI211_X1 U8305 ( .C1(n6569), .C2(n6568), .A(n8085), .B(n7971), .ZN(n6570)
         );
  OAI21_X1 U8306 ( .B1(n6724), .B2(n7998), .A(n6570), .ZN(n6571) );
  AOI21_X1 U8307 ( .B1(n9786), .B2(n8101), .A(n6571), .ZN(n6572) );
  OAI21_X1 U8308 ( .B1(n6598), .B2(n6573), .A(n6572), .ZN(P2_U3239) );
  INV_X1 U8309 ( .A(n7998), .ZN(n8097) );
  NAND2_X1 U8310 ( .A1(n6702), .A2(n8730), .ZN(n6574) );
  OAI21_X1 U8311 ( .B1(n7969), .B2(n8650), .A(n6574), .ZN(n9747) );
  NAND2_X1 U8312 ( .A1(n6576), .A2(n6575), .ZN(n6577) );
  NAND2_X1 U8313 ( .A1(n6578), .A2(n6577), .ZN(n6579) );
  AOI22_X1 U8314 ( .A1(n8097), .A2(n9747), .B1(n8085), .B2(n6579), .ZN(n6581)
         );
  NAND2_X1 U8315 ( .A1(n8101), .A2(n6689), .ZN(n6580) );
  OAI211_X1 U8316 ( .C1(n6598), .C2(n4801), .A(n6581), .B(n6580), .ZN(P2_U3224) );
  OAI222_X1 U8317 ( .A1(P2_U3152), .A2(n8268), .B1(n7319), .B2(n6583), .C1(
        n6582), .C2(n7947), .ZN(P2_U3338) );
  INV_X1 U8318 ( .A(n6584), .ZN(n6585) );
  OAI222_X1 U8319 ( .A1(n4258), .A2(n9974), .B1(n7850), .B2(n6585), .C1(
        P1_U3084), .C2(n7659), .ZN(P1_U3331) );
  OAI222_X1 U8320 ( .A1(n5462), .A2(P2_U3152), .B1(n7319), .B2(n6585), .C1(
        n7947), .C2(n5274), .ZN(P2_U3336) );
  NAND2_X1 U8321 ( .A1(n6589), .A2(n6586), .ZN(n6587) );
  OAI211_X1 U8322 ( .C1(n6588), .C2(n7947), .A(n6587), .B(n8311), .ZN(P2_U3335) );
  NAND2_X1 U8323 ( .A1(n6589), .A2(n7407), .ZN(n6591) );
  NOR2_X1 U8324 ( .A1(n6590), .A2(P1_U3084), .ZN(n7700) );
  INV_X1 U8325 ( .A(n7700), .ZN(n7410) );
  OAI211_X1 U8326 ( .C1(n6592), .C2(n4258), .A(n6591), .B(n7410), .ZN(P1_U3330) );
  INV_X1 U8327 ( .A(n6702), .ZN(n6593) );
  OAI22_X1 U8328 ( .A1(n6593), .A2(n8040), .B1(n8103), .B2(n9773), .ZN(n6595)
         );
  NAND2_X1 U8329 ( .A1(n6595), .A2(n6594), .ZN(n6597) );
  INV_X1 U8330 ( .A(n8068), .ZN(n8058) );
  AOI22_X1 U8331 ( .A1(n8058), .A2(n6691), .B1(n9754), .B2(n8101), .ZN(n6596)
         );
  OAI211_X1 U8332 ( .C1(n6598), .C2(n9734), .A(n6597), .B(n6596), .ZN(P2_U3234) );
  OAI222_X1 U8333 ( .A1(P2_U3152), .A2(n5463), .B1(n7319), .B2(n6600), .C1(
        n6599), .C2(n7947), .ZN(P2_U3337) );
  AOI21_X1 U8334 ( .B1(n8985), .B2(n9003), .A(n6601), .ZN(n6603) );
  NAND2_X1 U8335 ( .A1(n8986), .A2(n9653), .ZN(n6602) );
  OAI211_X1 U8336 ( .C1(n8989), .C2(n6604), .A(n6603), .B(n6602), .ZN(n6627)
         );
  INV_X2 U8337 ( .A(n6613), .ZN(n7823) );
  NAND2_X1 U8338 ( .A1(n7823), .A2(n6736), .ZN(n6606) );
  NAND2_X1 U8339 ( .A1(n6606), .A2(n6605), .ZN(n6607) );
  XNOR2_X1 U8340 ( .A(n6607), .B(n7806), .ZN(n6634) );
  INV_X2 U8341 ( .A(n6195), .ZN(n7796) );
  NAND2_X1 U8342 ( .A1(n7796), .A2(n6736), .ZN(n6608) );
  OAI21_X1 U8343 ( .B1(n7814), .B2(n6609), .A(n6608), .ZN(n6633) );
  XNOR2_X1 U8344 ( .A(n6634), .B(n6633), .ZN(n6641) );
  NAND2_X1 U8345 ( .A1(n6611), .A2(n6610), .ZN(n6616) );
  OR2_X1 U8346 ( .A1(n6195), .A2(n6615), .ZN(n6612) );
  OAI21_X1 U8347 ( .B1(n6613), .B2(n9699), .A(n6612), .ZN(n6614) );
  XNOR2_X1 U8348 ( .A(n6614), .B(n7821), .ZN(n6621) );
  OAI22_X1 U8349 ( .A1(n7814), .A2(n6615), .B1(n9699), .B2(n6195), .ZN(n6620)
         );
  NAND2_X1 U8350 ( .A1(n6621), .A2(n6620), .ZN(n8965) );
  AND2_X1 U8351 ( .A1(n6616), .A2(n8965), .ZN(n6617) );
  OAI21_X2 U8352 ( .B1(n6619), .B2(n6618), .A(n6617), .ZN(n6647) );
  INV_X1 U8353 ( .A(n6620), .ZN(n6623) );
  INV_X1 U8354 ( .A(n6621), .ZN(n6622) );
  NAND2_X1 U8355 ( .A1(n6623), .A2(n6622), .ZN(n8966) );
  NAND2_X1 U8356 ( .A1(n6647), .A2(n8966), .ZN(n6624) );
  XOR2_X1 U8357 ( .A(n6641), .B(n6624), .Z(n6625) );
  NOR2_X1 U8358 ( .A1(n6625), .A2(n8993), .ZN(n6626) );
  AOI211_X1 U8359 ( .C1(n8991), .C2(n6736), .A(n6627), .B(n6626), .ZN(n6628)
         );
  INV_X1 U8360 ( .A(n6628), .ZN(P1_U3211) );
  NAND2_X1 U8361 ( .A1(n6636), .A2(n9345), .ZN(n9706) );
  NAND2_X1 U8362 ( .A1(n6636), .A2(n7823), .ZN(n6631) );
  OR2_X1 U8363 ( .A1(n6195), .A2(n6629), .ZN(n6630) );
  NAND2_X1 U8364 ( .A1(n6631), .A2(n6630), .ZN(n6632) );
  XNOR2_X1 U8365 ( .A(n6632), .B(n7806), .ZN(n6802) );
  INV_X1 U8366 ( .A(n6633), .ZN(n6635) );
  NAND2_X1 U8367 ( .A1(n6635), .A2(n6634), .ZN(n6640) );
  AND2_X1 U8368 ( .A1(n8966), .A2(n6640), .ZN(n6646) );
  NAND2_X1 U8369 ( .A1(n6636), .A2(n7796), .ZN(n6638) );
  NAND2_X1 U8370 ( .A1(n7820), .A2(n9653), .ZN(n6637) );
  AND2_X1 U8371 ( .A1(n6638), .A2(n6637), .ZN(n6648) );
  INV_X1 U8372 ( .A(n6648), .ZN(n6639) );
  AND2_X1 U8373 ( .A1(n6646), .A2(n6639), .ZN(n6643) );
  INV_X1 U8374 ( .A(n6640), .ZN(n6642) );
  AOI21_X2 U8375 ( .B1(n6647), .B2(n6643), .A(n4281), .ZN(n6803) );
  AOI21_X1 U8376 ( .B1(n6647), .B2(n6646), .A(n6645), .ZN(n6649) );
  NAND2_X1 U8377 ( .A1(n6649), .A2(n6648), .ZN(n6805) );
  NAND2_X1 U8378 ( .A1(n6803), .A2(n6805), .ZN(n6650) );
  XOR2_X1 U8379 ( .A(n6802), .B(n6650), .Z(n6651) );
  NAND2_X1 U8380 ( .A1(n6651), .A2(n8969), .ZN(n6658) );
  INV_X1 U8381 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6652) );
  NOR2_X1 U8382 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6652), .ZN(n9525) );
  AOI21_X1 U8383 ( .B1(n8985), .B2(n9002), .A(n9525), .ZN(n6654) );
  NAND2_X1 U8384 ( .A1(n8986), .A2(n9001), .ZN(n6653) );
  OAI211_X1 U8385 ( .C1(n8989), .C2(n6655), .A(n6654), .B(n6653), .ZN(n6656)
         );
  INV_X1 U8386 ( .A(n6656), .ZN(n6657) );
  OAI211_X1 U8387 ( .C1(n8889), .C2(n9706), .A(n6658), .B(n6657), .ZN(P1_U3219) );
  AOI21_X1 U8388 ( .B1(n6660), .B2(n5018), .A(n6659), .ZN(n6662) );
  AOI22_X1 U8389 ( .A1(n6997), .A2(n5046), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7001), .ZN(n6661) );
  NOR2_X1 U8390 ( .A1(n6662), .A2(n6661), .ZN(n6999) );
  AOI21_X1 U8391 ( .B1(n6662), .B2(n6661), .A(n6999), .ZN(n6672) );
  NOR2_X1 U8392 ( .A1(n6997), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n6663) );
  AOI21_X1 U8393 ( .B1(P2_REG2_REG_14__SCAN_IN), .B2(n6997), .A(n6663), .ZN(
        n6667) );
  OAI21_X1 U8394 ( .B1(n6665), .B2(P2_REG2_REG_13__SCAN_IN), .A(n6664), .ZN(
        n6666) );
  OAI21_X1 U8395 ( .B1(n6667), .B2(n6666), .A(n7000), .ZN(n6670) );
  NAND2_X1 U8396 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7368) );
  NAND2_X1 U8397 ( .A1(n9376), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n6668) );
  OAI211_X1 U8398 ( .C1(n9739), .C2(n7001), .A(n7368), .B(n6668), .ZN(n6669)
         );
  AOI21_X1 U8399 ( .B1(n6670), .B2(n9733), .A(n6669), .ZN(n6671) );
  OAI21_X1 U8400 ( .B1(n6672), .B2(n9740), .A(n6671), .ZN(P2_U3259) );
  NAND2_X1 U8401 ( .A1(n9277), .A2(n6673), .ZN(n6675) );
  AOI22_X1 U8402 ( .A1(n9274), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9484), .ZN(n6674) );
  OAI211_X1 U8403 ( .C1(n6676), .C2(n9268), .A(n6675), .B(n6674), .ZN(n6677)
         );
  AOI21_X1 U8404 ( .B1(n7360), .B2(n6678), .A(n6677), .ZN(n6679) );
  OAI21_X1 U8405 ( .B1(n9676), .B2(n6680), .A(n6679), .ZN(P1_U3289) );
  NOR2_X1 U8406 ( .A1(n6681), .A2(P2_U3152), .ZN(n8755) );
  AND2_X1 U8407 ( .A1(n8755), .A2(n8760), .ZN(n6682) );
  NAND2_X1 U8408 ( .A1(n6713), .A2(n6682), .ZN(n6683) );
  INV_X1 U8409 ( .A(n6684), .ZN(n6686) );
  NAND2_X1 U8410 ( .A1(n6686), .A2(n8511), .ZN(n6685) );
  OR2_X1 U8411 ( .A1(n9762), .A2(n6685), .ZN(n7027) );
  XNOR2_X1 U8412 ( .A(n6686), .B(n5462), .ZN(n6687) );
  NAND2_X1 U8413 ( .A1(n6687), .A2(n4764), .ZN(n9791) );
  OR2_X1 U8414 ( .A1(n9762), .A2(n9791), .ZN(n6688) );
  NAND2_X1 U8415 ( .A1(n6690), .A2(n6689), .ZN(n6704) );
  NAND2_X1 U8416 ( .A1(n6704), .A2(n6703), .ZN(n9752) );
  NAND2_X1 U8417 ( .A1(n9752), .A2(n9751), .ZN(n6693) );
  OR2_X1 U8418 ( .A1(n6691), .A2(n6689), .ZN(n6692) );
  NAND2_X1 U8419 ( .A1(n6693), .A2(n6692), .ZN(n6722) );
  INV_X1 U8420 ( .A(n7969), .ZN(n8327) );
  NAND2_X1 U8421 ( .A1(n8327), .A2(n6714), .ZN(n6699) );
  NAND2_X1 U8422 ( .A1(n7969), .A2(n9786), .ZN(n6697) );
  NAND2_X1 U8423 ( .A1(n6722), .A2(n6721), .ZN(n6695) );
  NAND2_X1 U8424 ( .A1(n7969), .A2(n6714), .ZN(n6694) );
  NAND2_X1 U8425 ( .A1(n6695), .A2(n6694), .ZN(n7123) );
  XNOR2_X1 U8426 ( .A(n7123), .B(n6769), .ZN(n9796) );
  NAND2_X1 U8427 ( .A1(n6704), .A2(n6697), .ZN(n6698) );
  NAND2_X1 U8428 ( .A1(n6698), .A2(n6699), .ZN(n6701) );
  NAND2_X1 U8429 ( .A1(n6702), .A2(n9773), .ZN(n7103) );
  NAND2_X1 U8430 ( .A1(n6700), .A2(n6699), .ZN(n8136) );
  NOR2_X1 U8431 ( .A1(n6702), .A2(n9773), .ZN(n7102) );
  NAND2_X1 U8432 ( .A1(n7102), .A2(n6703), .ZN(n6705) );
  NAND2_X1 U8433 ( .A1(n6705), .A2(n6704), .ZN(n6723) );
  NOR2_X1 U8434 ( .A1(n6721), .A2(n6723), .ZN(n6706) );
  NOR2_X1 U8435 ( .A1(n4249), .A2(n6706), .ZN(n6707) );
  NAND2_X1 U8436 ( .A1(n6707), .A2(n6769), .ZN(n8135) );
  OAI21_X1 U8437 ( .B1(n6707), .B2(n6769), .A(n8135), .ZN(n6711) );
  AND2_X1 U8438 ( .A1(n8309), .A2(n8511), .ZN(n8270) );
  NAND2_X1 U8439 ( .A1(n8301), .A2(n8765), .ZN(n8120) );
  INV_X1 U8440 ( .A(n8120), .ZN(n6708) );
  NOR2_X1 U8441 ( .A1(n6933), .A2(n8650), .ZN(n6710) );
  NOR2_X1 U8442 ( .A1(n7969), .A2(n8648), .ZN(n6709) );
  OR2_X1 U8443 ( .A1(n6710), .A2(n6709), .ZN(n7974) );
  AOI21_X1 U8444 ( .B1(n6711), .B2(n9748), .A(n7974), .ZN(n9795) );
  AND3_X1 U8445 ( .A1(n8755), .A2(n4764), .A3(n8760), .ZN(n6712) );
  AND2_X1 U8446 ( .A1(n6713), .A2(n6712), .ZN(n7070) );
  AOI21_X1 U8447 ( .B1(n6728), .B2(n9793), .A(n9861), .ZN(n6715) );
  AND2_X1 U8448 ( .A1(n6715), .A2(n7131), .ZN(n9792) );
  INV_X1 U8449 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6716) );
  AOI22_X1 U8450 ( .A1(n7070), .A2(n9792), .B1(n9750), .B2(n6716), .ZN(n6718)
         );
  NAND2_X1 U8451 ( .A1(n9762), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6717) );
  OAI211_X1 U8452 ( .C1(n9762), .C2(n9795), .A(n6718), .B(n6717), .ZN(n6719)
         );
  AOI21_X1 U8453 ( .B1(n8743), .B2(n9793), .A(n6719), .ZN(n6720) );
  OAI21_X1 U8454 ( .B1(n8722), .B2(n9796), .A(n6720), .ZN(P2_U3293) );
  INV_X1 U8455 ( .A(n6721), .ZN(n8274) );
  XNOR2_X1 U8456 ( .A(n6722), .B(n8274), .ZN(n9789) );
  XNOR2_X1 U8457 ( .A(n6723), .B(n8274), .ZN(n6726) );
  INV_X1 U8458 ( .A(n6724), .ZN(n6725) );
  AOI21_X1 U8459 ( .B1(n6726), .B2(n9748), .A(n6725), .ZN(n9788) );
  NAND2_X1 U8460 ( .A1(n9778), .A2(n9773), .ZN(n6727) );
  AOI21_X1 U8461 ( .B1(n6727), .B2(n9786), .A(n9861), .ZN(n6729) );
  AND2_X1 U8462 ( .A1(n6729), .A2(n6728), .ZN(n9785) );
  AOI22_X1 U8463 ( .A1(n7070), .A2(n9785), .B1(n9750), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n6731) );
  NAND2_X1 U8464 ( .A1(n9762), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6730) );
  OAI211_X1 U8465 ( .C1(n9762), .C2(n9788), .A(n6731), .B(n6730), .ZN(n6732)
         );
  AOI21_X1 U8466 ( .B1(n8743), .B2(n9786), .A(n6732), .ZN(n6733) );
  OAI21_X1 U8467 ( .B1(n8722), .B2(n9789), .A(n6733), .ZN(P2_U3294) );
  AOI211_X1 U8468 ( .C1(n9345), .C2(n6736), .A(n6735), .B(n6734), .ZN(n6737)
         );
  OAI21_X1 U8469 ( .B1(n9349), .B2(n6738), .A(n6737), .ZN(n6740) );
  NAND2_X1 U8470 ( .A1(n6740), .A2(n9731), .ZN(n6739) );
  OAI21_X1 U8471 ( .B1(n9731), .B2(n5604), .A(n6739), .ZN(P1_U3530) );
  INV_X1 U8472 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n6742) );
  NAND2_X1 U8473 ( .A1(n6740), .A2(n9722), .ZN(n6741) );
  OAI21_X1 U8474 ( .B1(n9722), .B2(n6742), .A(n6741), .ZN(P1_U3475) );
  XNOR2_X1 U8475 ( .A(n6743), .B(n7442), .ZN(n9393) );
  INV_X1 U8476 ( .A(n7555), .ZN(n6747) );
  INV_X1 U8477 ( .A(n7442), .ZN(n6744) );
  OR2_X1 U8478 ( .A1(n6745), .A2(n6744), .ZN(n6746) );
  OAI211_X1 U8479 ( .C1(n6748), .C2(n6747), .A(n6746), .B(n9651), .ZN(n6750)
         );
  OR2_X1 U8480 ( .A1(n6809), .A2(n9212), .ZN(n6749) );
  OAI211_X1 U8481 ( .C1(n6870), .C2(n9210), .A(n6750), .B(n6749), .ZN(n6751)
         );
  AOI21_X1 U8482 ( .B1(n9393), .B2(n9659), .A(n6751), .ZN(n9395) );
  NAND2_X1 U8483 ( .A1(n9661), .A2(n9390), .ZN(n6752) );
  NAND2_X1 U8484 ( .A1(n6752), .A2(n9469), .ZN(n6753) );
  OR2_X1 U8485 ( .A1(n6976), .A2(n6753), .ZN(n9391) );
  OAI22_X1 U8486 ( .A1(n9666), .A2(n6754), .B1(n6918), .B2(n9663), .ZN(n6755)
         );
  AOI21_X1 U8487 ( .B1(n9669), .B2(n9390), .A(n6755), .ZN(n6756) );
  OAI21_X1 U8488 ( .B1(n9391), .B2(n7355), .A(n6756), .ZN(n6757) );
  AOI21_X1 U8489 ( .B1(n9393), .B2(n9673), .A(n6757), .ZN(n6758) );
  OAI21_X1 U8490 ( .B1(n9395), .B2(n9274), .A(n6758), .ZN(P1_U3281) );
  INV_X1 U8491 ( .A(n8042), .ZN(n9801) );
  NAND2_X1 U8492 ( .A1(n6933), .A2(n8042), .ZN(n8124) );
  INV_X1 U8493 ( .A(n8326), .ZN(n6772) );
  NAND2_X1 U8494 ( .A1(n6772), .A2(n9793), .ZN(n8132) );
  INV_X1 U8495 ( .A(n8132), .ZN(n6759) );
  NAND2_X1 U8496 ( .A1(n8135), .A2(n6760), .ZN(n6929) );
  NAND2_X1 U8497 ( .A1(n8325), .A2(n9810), .ZN(n8129) );
  NAND2_X1 U8498 ( .A1(n6929), .A2(n8125), .ZN(n6761) );
  INV_X1 U8499 ( .A(n8325), .ZN(n6779) );
  INV_X1 U8500 ( .A(n9810), .ZN(n6939) );
  NAND2_X1 U8501 ( .A1(n6779), .A2(n6939), .ZN(n8134) );
  NAND2_X1 U8502 ( .A1(n7091), .A2(n8080), .ZN(n8142) );
  INV_X1 U8503 ( .A(n8080), .ZN(n9819) );
  NAND2_X1 U8504 ( .A1(n8324), .A2(n9819), .ZN(n8141) );
  INV_X1 U8505 ( .A(n6955), .ZN(n8278) );
  XNOR2_X1 U8506 ( .A(n6956), .B(n8278), .ZN(n6763) );
  INV_X1 U8507 ( .A(n9748), .ZN(n8661) );
  INV_X1 U8508 ( .A(n8323), .ZN(n8145) );
  OAI22_X1 U8509 ( .A1(n8145), .A2(n8650), .B1(n6779), .B2(n8648), .ZN(n8081)
         );
  INV_X1 U8510 ( .A(n8081), .ZN(n6762) );
  OAI21_X1 U8511 ( .B1(n6763), .B2(n8661), .A(n6762), .ZN(n9821) );
  XNOR2_X1 U8512 ( .A(n6965), .B(n9819), .ZN(n6764) );
  NAND2_X1 U8513 ( .A1(n6764), .A2(n8832), .ZN(n9817) );
  INV_X1 U8514 ( .A(n9817), .ZN(n6766) );
  INV_X1 U8515 ( .A(n6765), .ZN(n8078) );
  AOI22_X1 U8516 ( .A1(n7070), .A2(n6766), .B1(n8078), .B2(n9750), .ZN(n6768)
         );
  NAND2_X1 U8517 ( .A1(n9762), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6767) );
  OAI211_X1 U8518 ( .C1(n9758), .C2(n9819), .A(n6768), .B(n6767), .ZN(n6784)
         );
  NAND2_X1 U8519 ( .A1(n6933), .A2(n9801), .ZN(n6773) );
  AND2_X1 U8520 ( .A1(n8279), .A2(n6771), .ZN(n6770) );
  NAND2_X1 U8521 ( .A1(n7123), .A2(n6770), .ZN(n6777) );
  INV_X1 U8522 ( .A(n9793), .ZN(n8127) );
  NAND2_X1 U8523 ( .A1(n6772), .A2(n8127), .ZN(n7124) );
  AND2_X1 U8524 ( .A1(n7124), .A2(n6773), .ZN(n6774) );
  NAND2_X1 U8525 ( .A1(n6777), .A2(n6776), .ZN(n6928) );
  NAND2_X1 U8526 ( .A1(n8134), .A2(n6939), .ZN(n6778) );
  NAND2_X1 U8527 ( .A1(n6928), .A2(n6778), .ZN(n6781) );
  NAND2_X1 U8528 ( .A1(n6779), .A2(n9810), .ZN(n6780) );
  NAND2_X1 U8529 ( .A1(n6782), .A2(n6955), .ZN(n9815) );
  AND3_X1 U8530 ( .A1(n9753), .A2(n9816), .A3(n9815), .ZN(n6783) );
  AOI211_X1 U8531 ( .C1(n6962), .C2(n9821), .A(n6784), .B(n6783), .ZN(n6785)
         );
  INV_X1 U8532 ( .A(n6785), .ZN(P2_U3290) );
  INV_X1 U8533 ( .A(n6786), .ZN(n6791) );
  OAI222_X1 U8534 ( .A1(n7850), .A2(n6791), .B1(P1_U3084), .B2(n6788), .C1(
        n6787), .C2(n4258), .ZN(P1_U3329) );
  INV_X1 U8535 ( .A(n6789), .ZN(n6792) );
  OAI222_X1 U8536 ( .A1(P2_U3152), .A2(n6792), .B1(n7319), .B2(n6791), .C1(
        n6790), .C2(n7947), .ZN(P2_U3334) );
  OAI22_X1 U8537 ( .A1(n8099), .A2(n6937), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n4840), .ZN(n6794) );
  OAI22_X1 U8538 ( .A1(n8074), .A2(n9810), .B1(n8068), .B2(n7091), .ZN(n6793)
         );
  AOI211_X1 U8539 ( .C1(n8059), .C2(n4400), .A(n6794), .B(n6793), .ZN(n6799)
         );
  NAND2_X1 U8540 ( .A1(n6796), .A2(n6795), .ZN(n6797) );
  NAND3_X1 U8541 ( .A1(n8085), .A2(n8083), .A3(n6797), .ZN(n6798) );
  NAND2_X1 U8542 ( .A1(n6799), .A2(n6798), .ZN(P2_U3229) );
  AND2_X1 U8543 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n9538) );
  AOI21_X1 U8544 ( .B1(n8985), .B2(n9653), .A(n9538), .ZN(n6801) );
  NAND2_X1 U8545 ( .A1(n8986), .A2(n9655), .ZN(n6800) );
  OAI211_X1 U8546 ( .C1(n8989), .C2(n9664), .A(n6801), .B(n6800), .ZN(n6813)
         );
  NAND2_X1 U8547 ( .A1(n6803), .A2(n6802), .ZN(n6804) );
  NAND2_X1 U8548 ( .A1(n6805), .A2(n6804), .ZN(n6861) );
  NAND2_X1 U8549 ( .A1(n9668), .A2(n7823), .ZN(n6807) );
  OR2_X1 U8550 ( .A1(n6195), .A2(n6809), .ZN(n6806) );
  NAND2_X1 U8551 ( .A1(n6807), .A2(n6806), .ZN(n6808) );
  XNOR2_X1 U8552 ( .A(n6808), .B(n7821), .ZN(n6862) );
  NOR2_X1 U8553 ( .A1(n7814), .A2(n6809), .ZN(n6810) );
  AOI21_X1 U8554 ( .B1(n9668), .B2(n7796), .A(n6810), .ZN(n6863) );
  XNOR2_X1 U8555 ( .A(n6862), .B(n6863), .ZN(n6860) );
  XOR2_X1 U8556 ( .A(n6861), .B(n6860), .Z(n6811) );
  NOR2_X1 U8557 ( .A1(n6811), .A2(n8993), .ZN(n6812) );
  AOI211_X1 U8558 ( .C1(n8991), .C2(n9668), .A(n6813), .B(n6812), .ZN(n6814)
         );
  INV_X1 U8559 ( .A(n6814), .ZN(P1_U3229) );
  INV_X1 U8560 ( .A(n6828), .ZN(n6815) );
  AOI211_X1 U8561 ( .C1(n6817), .C2(n6816), .A(n8103), .B(n6815), .ZN(n6822)
         );
  AOI22_X1 U8562 ( .A1(n8058), .A2(n8322), .B1(n8146), .B2(n8101), .ZN(n6820)
         );
  INV_X1 U8563 ( .A(n6818), .ZN(n7092) );
  AOI22_X1 U8564 ( .A1(n8079), .A2(n7092), .B1(P2_REG3_REG_7__SCAN_IN), .B2(
        P2_U3152), .ZN(n6819) );
  OAI211_X1 U8565 ( .C1(n7091), .C2(n8069), .A(n6820), .B(n6819), .ZN(n6821)
         );
  OR2_X1 U8566 ( .A1(n6822), .A2(n6821), .ZN(P2_U3215) );
  OAI21_X1 U8567 ( .B1(n8099), .B2(n7022), .A(n6823), .ZN(n6825) );
  INV_X1 U8568 ( .A(n7024), .ZN(n9830) );
  OAI22_X1 U8569 ( .A1(n8074), .A2(n9830), .B1(n8068), .B2(n7073), .ZN(n6824)
         );
  AOI211_X1 U8570 ( .C1(n8059), .C2(n8323), .A(n6825), .B(n6824), .ZN(n6834)
         );
  INV_X1 U8571 ( .A(n6826), .ZN(n6827) );
  AOI21_X1 U8572 ( .B1(n6828), .B2(n6827), .A(n8103), .ZN(n6832) );
  NOR3_X1 U8573 ( .A1(n8040), .A2(n8145), .A3(n6829), .ZN(n6831) );
  OAI21_X1 U8574 ( .B1(n6832), .B2(n6831), .A(n6830), .ZN(n6833) );
  NAND2_X1 U8575 ( .A1(n6834), .A2(n6833), .ZN(P2_U3223) );
  NOR2_X1 U8576 ( .A1(n6854), .A2(n6835), .ZN(n6836) );
  AOI21_X1 U8577 ( .B1(n6854), .B2(n6835), .A(n6836), .ZN(n6844) );
  INV_X1 U8578 ( .A(n9566), .ZN(n6840) );
  MUX2_X1 U8579 ( .A(n6837), .B(P1_REG1_REG_12__SCAN_IN), .S(n9566), .Z(n9567)
         );
  NOR2_X1 U8580 ( .A1(n9567), .A2(n9568), .ZN(n9572) );
  AOI21_X1 U8581 ( .B1(n6837), .B2(n6840), .A(n9572), .ZN(n9586) );
  NOR2_X1 U8582 ( .A1(n9583), .A2(n6841), .ZN(n6842) );
  AOI21_X1 U8583 ( .B1(n6841), .B2(n9583), .A(n6842), .ZN(n9585) );
  AOI21_X1 U8584 ( .B1(n6844), .B2(n6843), .A(n9046), .ZN(n6859) );
  NAND2_X1 U8585 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n7150) );
  OAI21_X1 U8586 ( .B1(n9523), .B2(n4434), .A(n7150), .ZN(n6845) );
  AOI21_X1 U8587 ( .B1(n9012), .B2(P1_ADDR_REG_14__SCAN_IN), .A(n6845), .ZN(
        n6858) );
  INV_X1 U8588 ( .A(n9562), .ZN(n6848) );
  INV_X1 U8589 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7034) );
  XNOR2_X1 U8590 ( .A(n9566), .B(n7034), .ZN(n9559) );
  NAND2_X1 U8591 ( .A1(n9566), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n6849) );
  NAND2_X1 U8592 ( .A1(n9560), .A2(n6849), .ZN(n9577) );
  NAND2_X1 U8593 ( .A1(n6852), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n6850) );
  OAI21_X1 U8594 ( .B1(n6852), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6850), .ZN(
        n9576) );
  INV_X1 U8595 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n6851) );
  NOR2_X1 U8596 ( .A1(n6852), .A2(n6851), .ZN(n6853) );
  INV_X1 U8597 ( .A(n9038), .ZN(n6855) );
  OAI211_X1 U8598 ( .C1(n6856), .C2(P1_REG2_REG_14__SCAN_IN), .A(n9526), .B(
        n6855), .ZN(n6857) );
  OAI211_X1 U8599 ( .C1(n6859), .C2(n9640), .A(n6858), .B(n6857), .ZN(P1_U3255) );
  NAND2_X1 U8600 ( .A1(n6861), .A2(n6860), .ZN(n6866) );
  INV_X1 U8601 ( .A(n6862), .ZN(n6864) );
  NAND2_X1 U8602 ( .A1(n6864), .A2(n6863), .ZN(n6865) );
  NAND2_X1 U8603 ( .A1(n6866), .A2(n6865), .ZN(n6919) );
  NAND2_X1 U8604 ( .A1(n7114), .A2(n7823), .ZN(n6868) );
  OR2_X1 U8605 ( .A1(n6195), .A2(n6870), .ZN(n6867) );
  NAND2_X1 U8606 ( .A1(n6868), .A2(n6867), .ZN(n6869) );
  XNOR2_X1 U8607 ( .A(n6869), .B(n7821), .ZN(n6874) );
  NOR2_X1 U8608 ( .A1(n7814), .A2(n6870), .ZN(n6871) );
  AOI21_X1 U8609 ( .B1(n7114), .B2(n7796), .A(n6871), .ZN(n6873) );
  INV_X1 U8610 ( .A(n6873), .ZN(n6872) );
  NAND2_X1 U8611 ( .A1(n6874), .A2(n6872), .ZN(n6888) );
  INV_X1 U8612 ( .A(n6888), .ZN(n6875) );
  XNOR2_X1 U8613 ( .A(n6874), .B(n6873), .ZN(n7054) );
  NOR2_X1 U8614 ( .A1(n6875), .A2(n7054), .ZN(n6885) );
  NAND2_X1 U8615 ( .A1(n9390), .A2(n7823), .ZN(n6877) );
  OR2_X1 U8616 ( .A1(n6195), .A2(n6879), .ZN(n6876) );
  NAND2_X1 U8617 ( .A1(n6877), .A2(n6876), .ZN(n6878) );
  XNOR2_X1 U8618 ( .A(n6878), .B(n7806), .ZN(n6921) );
  NOR2_X1 U8619 ( .A1(n7814), .A2(n6879), .ZN(n6880) );
  AOI21_X1 U8620 ( .B1(n9390), .B2(n7796), .A(n6880), .ZN(n6920) );
  AND2_X1 U8621 ( .A1(n6921), .A2(n6920), .ZN(n7051) );
  NAND2_X1 U8622 ( .A1(n7038), .A2(n7823), .ZN(n6882) );
  OR2_X1 U8623 ( .A1(n6195), .A2(n7236), .ZN(n6881) );
  NAND2_X1 U8624 ( .A1(n6882), .A2(n6881), .ZN(n6883) );
  XNOR2_X1 U8625 ( .A(n6883), .B(n7806), .ZN(n6890) );
  NOR2_X1 U8626 ( .A1(n7814), .A2(n7236), .ZN(n6884) );
  AOI21_X1 U8627 ( .B1(n7038), .B2(n7796), .A(n6884), .ZN(n6891) );
  NAND2_X1 U8628 ( .A1(n6890), .A2(n6891), .ZN(n6895) );
  INV_X1 U8629 ( .A(n6895), .ZN(n6897) );
  OR2_X1 U8630 ( .A1(n6986), .A2(n6897), .ZN(n6899) );
  INV_X1 U8631 ( .A(n6921), .ZN(n6887) );
  INV_X1 U8632 ( .A(n6920), .ZN(n6886) );
  NAND2_X1 U8633 ( .A1(n6887), .A2(n6886), .ZN(n7052) );
  INV_X1 U8634 ( .A(n6890), .ZN(n6893) );
  INV_X1 U8635 ( .A(n6891), .ZN(n6892) );
  NAND2_X1 U8636 ( .A1(n6893), .A2(n6892), .ZN(n6894) );
  NAND2_X1 U8637 ( .A1(n6895), .A2(n6894), .ZN(n6990) );
  INV_X1 U8638 ( .A(n6990), .ZN(n6896) );
  NAND2_X1 U8639 ( .A1(n7256), .A2(n7823), .ZN(n6901) );
  OR2_X1 U8640 ( .A1(n6195), .A2(n6903), .ZN(n6900) );
  NAND2_X1 U8641 ( .A1(n6901), .A2(n6900), .ZN(n6902) );
  XNOR2_X1 U8642 ( .A(n6902), .B(n7806), .ZN(n6905) );
  NOR2_X1 U8643 ( .A1(n7814), .A2(n6903), .ZN(n6904) );
  AOI21_X1 U8644 ( .B1(n7256), .B2(n7796), .A(n6904), .ZN(n6906) );
  NAND2_X1 U8645 ( .A1(n6905), .A2(n6906), .ZN(n7139) );
  INV_X1 U8646 ( .A(n6905), .ZN(n6908) );
  INV_X1 U8647 ( .A(n6906), .ZN(n6907) );
  NAND2_X1 U8648 ( .A1(n6908), .A2(n6907), .ZN(n7141) );
  NAND2_X1 U8649 ( .A1(n7139), .A2(n7141), .ZN(n6909) );
  XOR2_X1 U8650 ( .A(n7140), .B(n6909), .Z(n6914) );
  AND2_X1 U8651 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9582) );
  INV_X1 U8652 ( .A(n8986), .ZN(n8956) );
  NOR2_X1 U8653 ( .A1(n8956), .A2(n7472), .ZN(n6910) );
  AOI211_X1 U8654 ( .C1(n8985), .C2(n8999), .A(n9582), .B(n6910), .ZN(n6911)
         );
  OAI21_X1 U8655 ( .B1(n8989), .B2(n7241), .A(n6911), .ZN(n6912) );
  AOI21_X1 U8656 ( .B1(n8991), .B2(n7256), .A(n6912), .ZN(n6913) );
  OAI21_X1 U8657 ( .B1(n6914), .B2(n8993), .A(n6913), .ZN(P1_U3232) );
  NOR2_X1 U8658 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6915), .ZN(n9550) );
  AOI21_X1 U8659 ( .B1(n8985), .B2(n9001), .A(n9550), .ZN(n6917) );
  NAND2_X1 U8660 ( .A1(n8986), .A2(n9000), .ZN(n6916) );
  OAI211_X1 U8661 ( .C1(n8989), .C2(n6918), .A(n6917), .B(n6916), .ZN(n6925)
         );
  XNOR2_X1 U8662 ( .A(n6921), .B(n6920), .ZN(n6922) );
  XNOR2_X1 U8663 ( .A(n6919), .B(n6922), .ZN(n6923) );
  NOR2_X1 U8664 ( .A1(n6923), .A2(n8993), .ZN(n6924) );
  AOI211_X1 U8665 ( .C1(n8991), .C2(n9390), .A(n6925), .B(n6924), .ZN(n6926)
         );
  INV_X1 U8666 ( .A(n6926), .ZN(P1_U3215) );
  NAND2_X1 U8667 ( .A1(n8134), .A2(n8129), .ZN(n8273) );
  INV_X1 U8668 ( .A(n8273), .ZN(n6927) );
  XNOR2_X1 U8669 ( .A(n6928), .B(n6927), .ZN(n9808) );
  NAND2_X1 U8670 ( .A1(n6929), .A2(n6930), .ZN(n6931) );
  XNOR2_X1 U8671 ( .A(n6931), .B(n8273), .ZN(n6932) );
  NAND2_X1 U8672 ( .A1(n6932), .A2(n9748), .ZN(n6936) );
  OAI22_X1 U8673 ( .A1(n7091), .A2(n8650), .B1(n6933), .B2(n8648), .ZN(n6934)
         );
  INV_X1 U8674 ( .A(n6934), .ZN(n6935) );
  NAND2_X1 U8675 ( .A1(n6936), .A2(n6935), .ZN(n9813) );
  OAI211_X1 U8676 ( .C1(n7132), .C2(n9810), .A(n8832), .B(n6965), .ZN(n9809)
         );
  OAI22_X1 U8677 ( .A1(n9809), .A2(n8511), .B1(n8739), .B2(n6937), .ZN(n6938)
         );
  OAI21_X1 U8678 ( .B1(n9813), .B2(n6938), .A(n6962), .ZN(n6941) );
  AOI22_X1 U8679 ( .A1(n8743), .A2(n6939), .B1(P2_REG2_REG_5__SCAN_IN), .B2(
        n8655), .ZN(n6940) );
  OAI211_X1 U8680 ( .C1(n8722), .C2(n9808), .A(n6941), .B(n6940), .ZN(P2_U3291) );
  INV_X1 U8681 ( .A(n6942), .ZN(n6946) );
  OAI222_X1 U8682 ( .A1(n4258), .A2(n6944), .B1(n7850), .B2(n6946), .C1(n6943), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  OAI222_X1 U8683 ( .A1(n6947), .A2(P2_U3152), .B1(n7319), .B2(n6946), .C1(
        n6945), .C2(n7947), .ZN(P2_U3333) );
  NAND2_X1 U8684 ( .A1(n8324), .A2(n8080), .ZN(n6948) );
  NAND2_X1 U8685 ( .A1(n6958), .A2(n7024), .ZN(n8152) );
  NAND2_X1 U8686 ( .A1(n8322), .A2(n9830), .ZN(n8151) );
  NOR2_X1 U8687 ( .A1(n8323), .A2(n8146), .ZN(n7009) );
  NOR2_X1 U8688 ( .A1(n8276), .A2(n7009), .ZN(n6949) );
  NAND2_X1 U8689 ( .A1(n7086), .A2(n6949), .ZN(n6952) );
  INV_X1 U8690 ( .A(n6952), .ZN(n7012) );
  NOR2_X1 U8691 ( .A1(n6958), .A2(n9830), .ZN(n6950) );
  NAND2_X1 U8692 ( .A1(n7073), .A2(n6968), .ZN(n8154) );
  INV_X1 U8693 ( .A(n7073), .ZN(n8321) );
  NAND2_X1 U8694 ( .A1(n9837), .A2(n8321), .ZN(n8162) );
  OAI21_X1 U8695 ( .B1(n7012), .B2(n6950), .A(n8282), .ZN(n6953) );
  NOR2_X1 U8696 ( .A1(n8282), .A2(n6950), .ZN(n6951) );
  AND2_X1 U8697 ( .A1(n6953), .A2(n7075), .ZN(n9836) );
  NAND2_X1 U8698 ( .A1(n7088), .A2(n4269), .ZN(n7087) );
  NAND2_X1 U8699 ( .A1(n8323), .A2(n9823), .ZN(n6957) );
  NAND2_X1 U8700 ( .A1(n7015), .A2(n8276), .ZN(n7014) );
  NAND2_X1 U8701 ( .A1(n7014), .A2(n8152), .ZN(n7060) );
  XNOR2_X1 U8702 ( .A(n7060), .B(n8282), .ZN(n6960) );
  OAI22_X1 U8703 ( .A1(n7062), .A2(n8650), .B1(n6958), .B2(n8648), .ZN(n6959)
         );
  AOI21_X1 U8704 ( .B1(n6960), .B2(n9748), .A(n6959), .ZN(n6961) );
  OAI21_X1 U8705 ( .B1(n9836), .B2(n9791), .A(n6961), .ZN(n9839) );
  INV_X1 U8706 ( .A(n9762), .ZN(n6962) );
  NAND2_X1 U8707 ( .A1(n9839), .A2(n6962), .ZN(n6970) );
  OAI22_X1 U8708 ( .A1(n6962), .A2(n6964), .B1(n6963), .B2(n8739), .ZN(n6967)
         );
  NAND2_X1 U8709 ( .A1(n7021), .A2(n9837), .ZN(n7067) );
  OAI21_X1 U8710 ( .B1(n7021), .B2(n9837), .A(n7067), .ZN(n9838) );
  NOR2_X1 U8711 ( .A1(n8745), .A2(n9838), .ZN(n6966) );
  AOI211_X1 U8712 ( .C1(n8743), .C2(n6968), .A(n6967), .B(n6966), .ZN(n6969)
         );
  OAI211_X1 U8713 ( .C1(n9836), .C2(n7027), .A(n6970), .B(n6969), .ZN(P2_U3287) );
  XNOR2_X1 U8714 ( .A(n7114), .B(n9000), .ZN(n7567) );
  XOR2_X1 U8715 ( .A(n6971), .B(n7567), .Z(n7113) );
  XNOR2_X1 U8716 ( .A(n6972), .B(n7567), .ZN(n6974) );
  AOI22_X1 U8717 ( .A1(n9654), .A2(n9655), .B1(n8999), .B2(n9656), .ZN(n6973)
         );
  OAI21_X1 U8718 ( .B1(n6974), .B2(n9207), .A(n6973), .ZN(n6975) );
  AOI21_X1 U8719 ( .B1(n7113), .B2(n9659), .A(n6975), .ZN(n7117) );
  AOI21_X1 U8720 ( .B1(n7114), .B2(n4457), .A(n7035), .ZN(n7115) );
  NOR2_X1 U8721 ( .A1(n6977), .A2(n9268), .ZN(n6980) );
  OAI22_X1 U8722 ( .A1(n9666), .A2(n6978), .B1(n7050), .B2(n9663), .ZN(n6979)
         );
  AOI211_X1 U8723 ( .C1(n7115), .C2(n9277), .A(n6980), .B(n6979), .ZN(n6982)
         );
  NAND2_X1 U8724 ( .A1(n7113), .A2(n9673), .ZN(n6981) );
  OAI211_X1 U8725 ( .C1(n7117), .C2(n9274), .A(n6982), .B(n6981), .ZN(P1_U3280) );
  INV_X1 U8726 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n6983) );
  NOR2_X1 U8727 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6983), .ZN(n9565) );
  AOI21_X1 U8728 ( .B1(n8985), .B2(n9000), .A(n9565), .ZN(n6985) );
  NAND2_X1 U8729 ( .A1(n8986), .A2(n8998), .ZN(n6984) );
  OAI211_X1 U8730 ( .C1(n8989), .C2(n7033), .A(n6985), .B(n6984), .ZN(n6995)
         );
  OR2_X1 U8731 ( .A1(n6919), .A2(n6986), .ZN(n6989) );
  NAND2_X1 U8732 ( .A1(n6989), .A2(n6987), .ZN(n6993) );
  NAND2_X1 U8733 ( .A1(n6989), .A2(n6988), .ZN(n6991) );
  NAND2_X1 U8734 ( .A1(n6991), .A2(n6990), .ZN(n6992) );
  AOI21_X1 U8735 ( .B1(n6993), .B2(n6992), .A(n8993), .ZN(n6994) );
  AOI211_X1 U8736 ( .C1(n8991), .C2(n7038), .A(n6995), .B(n6994), .ZN(n6996)
         );
  INV_X1 U8737 ( .A(n6996), .ZN(P1_U3222) );
  NOR2_X1 U8738 ( .A1(n6997), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6998) );
  NOR2_X1 U8739 ( .A1(n6999), .A2(n6998), .ZN(n8393) );
  XNOR2_X1 U8740 ( .A(n8393), .B(n8406), .ZN(n8397) );
  XOR2_X1 U8741 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8397), .Z(n7008) );
  XNOR2_X1 U8742 ( .A(n7002), .B(n8395), .ZN(n8404) );
  XNOR2_X1 U8743 ( .A(n8404), .B(P2_REG2_REG_15__SCAN_IN), .ZN(n7006) );
  NOR2_X1 U8744 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10008), .ZN(n7003) );
  AOI21_X1 U8745 ( .B1(n9376), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7003), .ZN(
        n7004) );
  OAI21_X1 U8746 ( .B1(n9739), .B2(n8395), .A(n7004), .ZN(n7005) );
  AOI21_X1 U8747 ( .B1(n7006), .B2(n9733), .A(n7005), .ZN(n7007) );
  OAI21_X1 U8748 ( .B1(n7008), .B2(n9740), .A(n7007), .ZN(P2_U3260) );
  INV_X1 U8749 ( .A(n7009), .ZN(n7010) );
  NAND2_X1 U8750 ( .A1(n7086), .A2(n7010), .ZN(n7011) );
  AND2_X1 U8751 ( .A1(n7011), .A2(n8276), .ZN(n7013) );
  OR2_X1 U8752 ( .A1(n7013), .A2(n7012), .ZN(n9829) );
  AOI22_X1 U8753 ( .A1(n8321), .A2(n8729), .B1(n8730), .B2(n8323), .ZN(n7018)
         );
  OAI21_X1 U8754 ( .B1(n7015), .B2(n8276), .A(n7014), .ZN(n7016) );
  NAND2_X1 U8755 ( .A1(n7016), .A2(n9748), .ZN(n7017) );
  OAI211_X1 U8756 ( .C1(n9829), .C2(n9791), .A(n7018), .B(n7017), .ZN(n9832)
         );
  MUX2_X1 U8757 ( .A(n9832), .B(P2_REG2_REG_8__SCAN_IN), .S(n9762), .Z(n7019)
         );
  INV_X1 U8758 ( .A(n7019), .ZN(n7026) );
  NOR2_X1 U8759 ( .A1(n7094), .A2(n9830), .ZN(n7020) );
  OR2_X1 U8760 ( .A1(n7021), .A2(n7020), .ZN(n9831) );
  OAI22_X1 U8761 ( .A1(n8745), .A2(n9831), .B1(n7022), .B2(n8739), .ZN(n7023)
         );
  AOI21_X1 U8762 ( .B1(n8743), .B2(n7024), .A(n7023), .ZN(n7025) );
  OAI211_X1 U8763 ( .C1(n9829), .C2(n7027), .A(n7026), .B(n7025), .ZN(P2_U3288) );
  NAND2_X1 U8764 ( .A1(n7029), .A2(n7028), .ZN(n7030) );
  XNOR2_X1 U8765 ( .A(n7030), .B(n7443), .ZN(n7031) );
  AOI222_X1 U8766 ( .A1(n9651), .A2(n7031), .B1(n8998), .B2(n9656), .C1(n9000), 
        .C2(n9654), .ZN(n9499) );
  XOR2_X1 U8767 ( .A(n7032), .B(n7443), .Z(n9502) );
  NAND2_X1 U8768 ( .A1(n9502), .A2(n7360), .ZN(n7040) );
  OAI22_X1 U8769 ( .A1(n9666), .A2(n7034), .B1(n7033), .B2(n9663), .ZN(n7037)
         );
  OAI211_X1 U8770 ( .C1(n7035), .C2(n9500), .A(n9469), .B(n7240), .ZN(n9498)
         );
  NOR2_X1 U8771 ( .A1(n9498), .A2(n7355), .ZN(n7036) );
  AOI211_X1 U8772 ( .C1(n9669), .C2(n7038), .A(n7037), .B(n7036), .ZN(n7039)
         );
  OAI211_X1 U8773 ( .C1(n9676), .C2(n9499), .A(n7040), .B(n7039), .ZN(P1_U3279) );
  XNOR2_X1 U8774 ( .A(n7042), .B(n7041), .ZN(n7046) );
  OAI22_X1 U8775 ( .A1(n7328), .A2(n8650), .B1(n7073), .B2(n8648), .ZN(n7065)
         );
  AOI22_X1 U8776 ( .A1(n8097), .A2(n7065), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n7045) );
  INV_X1 U8777 ( .A(n7043), .ZN(n7071) );
  AOI22_X1 U8778 ( .A1(n8101), .A2(n9844), .B1(n8079), .B2(n7071), .ZN(n7044)
         );
  OAI211_X1 U8779 ( .C1(n7046), .C2(n8103), .A(n7045), .B(n7044), .ZN(P2_U3219) );
  AOI21_X1 U8780 ( .B1(n8985), .B2(n9655), .A(n7047), .ZN(n7049) );
  NAND2_X1 U8781 ( .A1(n8986), .A2(n8999), .ZN(n7048) );
  OAI211_X1 U8782 ( .C1(n8989), .C2(n7050), .A(n7049), .B(n7048), .ZN(n7058)
         );
  OR2_X1 U8783 ( .A1(n6919), .A2(n7051), .ZN(n7053) );
  NAND2_X1 U8784 ( .A1(n7053), .A2(n7052), .ZN(n7055) );
  XNOR2_X1 U8785 ( .A(n7055), .B(n7054), .ZN(n7056) );
  NOR2_X1 U8786 ( .A1(n7056), .A2(n8993), .ZN(n7057) );
  AOI211_X1 U8787 ( .C1(n8991), .C2(n7114), .A(n7058), .B(n7057), .ZN(n7059)
         );
  INV_X1 U8788 ( .A(n7059), .ZN(P1_U3234) );
  NAND2_X1 U8789 ( .A1(n7060), .A2(n8282), .ZN(n7061) );
  NAND2_X1 U8790 ( .A1(n7061), .A2(n8154), .ZN(n7063) );
  NAND2_X1 U8791 ( .A1(n9844), .A2(n7062), .ZN(n8160) );
  NAND2_X1 U8792 ( .A1(n8161), .A2(n8160), .ZN(n8159) );
  AOI21_X1 U8793 ( .B1(n7063), .B2(n8159), .A(n8661), .ZN(n7066) );
  INV_X1 U8794 ( .A(n7063), .ZN(n7064) );
  NAND2_X1 U8795 ( .A1(n7064), .A2(n8281), .ZN(n7157) );
  AOI21_X1 U8796 ( .B1(n7066), .B2(n7157), .A(n7065), .ZN(n9849) );
  INV_X1 U8797 ( .A(n7067), .ZN(n7069) );
  INV_X1 U8798 ( .A(n9844), .ZN(n7068) );
  OAI211_X1 U8799 ( .C1(n7069), .C2(n7068), .A(n8832), .B(n7163), .ZN(n9845)
         );
  INV_X1 U8800 ( .A(n7070), .ZN(n8718) );
  AOI22_X1 U8801 ( .A1(n9762), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7071), .B2(
        n9750), .ZN(n7072) );
  OAI21_X1 U8802 ( .B1(n9845), .B2(n8718), .A(n7072), .ZN(n7079) );
  NAND2_X1 U8803 ( .A1(n7073), .A2(n9837), .ZN(n7074) );
  INV_X1 U8804 ( .A(n8159), .ZN(n8281) );
  NAND2_X1 U8805 ( .A1(n7076), .A2(n8281), .ZN(n7077) );
  NAND2_X1 U8806 ( .A1(n7160), .A2(n7077), .ZN(n9848) );
  NOR2_X1 U8807 ( .A1(n9848), .A2(n8722), .ZN(n7078) );
  AOI211_X1 U8808 ( .C1(n8743), .C2(n9844), .A(n7079), .B(n7078), .ZN(n7080)
         );
  OAI21_X1 U8809 ( .B1(n9762), .B2(n9849), .A(n7080), .ZN(P2_U3286) );
  INV_X1 U8810 ( .A(n7081), .ZN(n7111) );
  OAI222_X1 U8811 ( .A1(n7850), .A2(n7111), .B1(P1_U3084), .B2(n7083), .C1(
        n7082), .C2(n4258), .ZN(P1_U3327) );
  NAND2_X1 U8812 ( .A1(n7084), .A2(n4269), .ZN(n7085) );
  NAND2_X1 U8813 ( .A1(n7086), .A2(n7085), .ZN(n9827) );
  INV_X1 U8814 ( .A(n9827), .ZN(n7101) );
  OAI211_X1 U8815 ( .C1(n7088), .C2(n4269), .A(n7087), .B(n9748), .ZN(n7090)
         );
  NAND2_X1 U8816 ( .A1(n8322), .A2(n8729), .ZN(n7089) );
  OAI211_X1 U8817 ( .C1(n7091), .C2(n8648), .A(n7090), .B(n7089), .ZN(n9825)
         );
  AOI22_X1 U8818 ( .A1(n8655), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7092), .B2(
        n9750), .ZN(n7098) );
  AND2_X1 U8819 ( .A1(n7093), .A2(n8146), .ZN(n7095) );
  OR2_X1 U8820 ( .A1(n7095), .A2(n7094), .ZN(n9824) );
  INV_X1 U8821 ( .A(n9824), .ZN(n7096) );
  NAND2_X1 U8822 ( .A1(n9755), .A2(n7096), .ZN(n7097) );
  OAI211_X1 U8823 ( .C1(n9758), .C2(n9823), .A(n7098), .B(n7097), .ZN(n7099)
         );
  AOI21_X1 U8824 ( .B1(n9825), .B2(n6962), .A(n7099), .ZN(n7100) );
  OAI21_X1 U8825 ( .B1(n8722), .B2(n7101), .A(n7100), .ZN(P2_U3289) );
  INV_X1 U8826 ( .A(n7102), .ZN(n9746) );
  AND2_X1 U8827 ( .A1(n9746), .A2(n7103), .ZN(n9774) );
  OAI22_X1 U8828 ( .A1(n9774), .A2(n8661), .B1(n6690), .B2(n8650), .ZN(n9776)
         );
  AND2_X1 U8829 ( .A1(n9750), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n7104) );
  NOR2_X1 U8830 ( .A1(n9776), .A2(n7104), .ZN(n7105) );
  NOR2_X1 U8831 ( .A1(n8655), .A2(n7105), .ZN(n7107) );
  AOI21_X1 U8832 ( .B1(n8745), .B2(n9758), .A(n9773), .ZN(n7106) );
  AOI211_X1 U8833 ( .C1(n9762), .C2(P2_REG2_REG_0__SCAN_IN), .A(n7107), .B(
        n7106), .ZN(n7108) );
  OAI21_X1 U8834 ( .B1(n9774), .B2(n8722), .A(n7108), .ZN(P2_U3296) );
  INV_X1 U8835 ( .A(n7109), .ZN(n7112) );
  OAI222_X1 U8836 ( .A1(P2_U3152), .A2(n7112), .B1(n7949), .B2(n7111), .C1(
        n7110), .C2(n7947), .ZN(P2_U3332) );
  INV_X1 U8837 ( .A(n7113), .ZN(n7118) );
  AOI22_X1 U8838 ( .A1(n7115), .A2(n9469), .B1(n9345), .B2(n7114), .ZN(n7116)
         );
  OAI211_X1 U8839 ( .C1(n9389), .C2(n7118), .A(n7117), .B(n7116), .ZN(n7120)
         );
  NAND2_X1 U8840 ( .A1(n7120), .A2(n9731), .ZN(n7119) );
  OAI21_X1 U8841 ( .B1(n9731), .B2(n5661), .A(n7119), .ZN(P1_U3534) );
  INV_X1 U8842 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7122) );
  NAND2_X1 U8843 ( .A1(n7120), .A2(n9722), .ZN(n7121) );
  OAI21_X1 U8844 ( .B1(n9722), .B2(n7122), .A(n7121), .ZN(P1_U3487) );
  NAND2_X1 U8845 ( .A1(n7123), .A2(n8279), .ZN(n7125) );
  NAND2_X1 U8846 ( .A1(n7125), .A2(n7124), .ZN(n7126) );
  XNOR2_X1 U8847 ( .A(n7126), .B(n7127), .ZN(n9800) );
  AND2_X1 U8848 ( .A1(n8135), .A2(n8132), .ZN(n7128) );
  OAI211_X1 U8849 ( .C1(n7128), .C2(n7127), .A(n6929), .B(n9748), .ZN(n7130)
         );
  AOI22_X1 U8850 ( .A1(n8730), .A2(n8326), .B1(n8325), .B2(n8729), .ZN(n7129)
         );
  AND2_X1 U8851 ( .A1(n7130), .A2(n7129), .ZN(n9803) );
  OAI22_X1 U8852 ( .A1(n9803), .A2(n8655), .B1(n8047), .B2(n8739), .ZN(n7135)
         );
  INV_X1 U8853 ( .A(n7132), .ZN(n7133) );
  OAI21_X1 U8854 ( .B1(n9801), .B2(n4522), .A(n7133), .ZN(n9802) );
  OAI22_X1 U8855 ( .A1(n8745), .A2(n9802), .B1(n6962), .B2(n4480), .ZN(n7134)
         );
  AOI211_X1 U8856 ( .C1(n8743), .C2(n8042), .A(n7135), .B(n7134), .ZN(n7136)
         );
  OAI21_X1 U8857 ( .B1(n8722), .B2(n9800), .A(n7136), .ZN(P2_U3292) );
  NAND2_X1 U8858 ( .A1(n7473), .A2(n7796), .ZN(n7138) );
  NAND2_X1 U8859 ( .A1(n7820), .A2(n9477), .ZN(n7137) );
  NAND2_X1 U8860 ( .A1(n7138), .A2(n7137), .ZN(n7191) );
  NAND2_X1 U8861 ( .A1(n7140), .A2(n7139), .ZN(n7142) );
  NAND2_X1 U8862 ( .A1(n7473), .A2(n7823), .ZN(n7144) );
  OR2_X1 U8863 ( .A1(n6195), .A2(n7472), .ZN(n7143) );
  NAND2_X1 U8864 ( .A1(n7144), .A2(n7143), .ZN(n7145) );
  XNOR2_X1 U8865 ( .A(n7145), .B(n7821), .ZN(n7147) );
  NAND2_X1 U8866 ( .A1(n7148), .A2(n7147), .ZN(n7199) );
  NAND2_X1 U8867 ( .A1(n7192), .A2(n7199), .ZN(n7149) );
  XOR2_X1 U8868 ( .A(n7191), .B(n7149), .Z(n7155) );
  NAND2_X1 U8869 ( .A1(n8985), .A2(n8998), .ZN(n7151) );
  OAI211_X1 U8870 ( .C1(n8956), .C2(n7193), .A(n7151), .B(n7150), .ZN(n7152)
         );
  AOI21_X1 U8871 ( .B1(n7216), .B2(n8975), .A(n7152), .ZN(n7154) );
  NAND2_X1 U8872 ( .A1(n7473), .A2(n8991), .ZN(n7153) );
  OAI211_X1 U8873 ( .C1(n7155), .C2(n8993), .A(n7154), .B(n7153), .ZN(P1_U3213) );
  INV_X1 U8874 ( .A(n7156), .ZN(n7190) );
  OAI222_X1 U8875 ( .A1(n7850), .A2(n7190), .B1(n6046), .B2(P1_U3084), .C1(
        n10040), .C2(n4258), .ZN(P1_U3326) );
  OR2_X1 U8876 ( .A1(n7251), .A2(n7328), .ZN(n8169) );
  NAND2_X1 U8877 ( .A1(n7251), .A2(n7328), .ZN(n8170) );
  NAND2_X1 U8878 ( .A1(n7881), .A2(n7299), .ZN(n7171) );
  OAI21_X1 U8879 ( .B1(n7881), .B2(n7299), .A(n7171), .ZN(n7158) );
  AOI222_X1 U8880 ( .A1(n9748), .A2(n7158), .B1(n8318), .B2(n8729), .C1(n8320), 
        .C2(n8730), .ZN(n9855) );
  NAND2_X1 U8881 ( .A1(n8320), .A2(n9844), .ZN(n7159) );
  NAND2_X1 U8882 ( .A1(n7161), .A2(n8285), .ZN(n7177) );
  OAI21_X1 U8883 ( .B1(n7161), .B2(n8285), .A(n7177), .ZN(n7162) );
  INV_X1 U8884 ( .A(n7162), .ZN(n9858) );
  NAND2_X1 U8885 ( .A1(n7163), .A2(n7251), .ZN(n7164) );
  NAND2_X1 U8886 ( .A1(n7180), .A2(n7164), .ZN(n9854) );
  OAI22_X1 U8887 ( .A1(n6962), .A2(n7165), .B1(n7250), .B2(n8739), .ZN(n7166)
         );
  AOI21_X1 U8888 ( .B1(n8743), .B2(n7251), .A(n7166), .ZN(n7167) );
  OAI21_X1 U8889 ( .B1(n8745), .B2(n9854), .A(n7167), .ZN(n7168) );
  AOI21_X1 U8890 ( .B1(n9858), .B2(n9753), .A(n7168), .ZN(n7169) );
  OAI21_X1 U8891 ( .B1(n9855), .B2(n8655), .A(n7169), .ZN(P2_U3285) );
  AND2_X1 U8892 ( .A1(n7171), .A2(n8170), .ZN(n7173) );
  NAND2_X1 U8893 ( .A1(n7170), .A2(n7306), .ZN(n8174) );
  NAND2_X1 U8894 ( .A1(n7171), .A2(n7300), .ZN(n7172) );
  OAI211_X1 U8895 ( .C1(n7173), .C2(n7178), .A(n7172), .B(n9748), .ZN(n7175)
         );
  INV_X1 U8896 ( .A(n7365), .ZN(n8731) );
  NAND2_X1 U8897 ( .A1(n8731), .A2(n8729), .ZN(n7174) );
  OAI211_X1 U8898 ( .C1(n7328), .C2(n8648), .A(n7175), .B(n7174), .ZN(n9863)
         );
  INV_X1 U8899 ( .A(n9863), .ZN(n7188) );
  NAND2_X1 U8900 ( .A1(n7251), .A2(n8319), .ZN(n7176) );
  OAI21_X1 U8901 ( .B1(n7179), .B2(n8284), .A(n7312), .ZN(n9865) );
  INV_X1 U8902 ( .A(n7910), .ZN(n7182) );
  NAND2_X1 U8903 ( .A1(n7180), .A2(n7170), .ZN(n7181) );
  NAND2_X1 U8904 ( .A1(n7182), .A2(n7181), .ZN(n9862) );
  OAI22_X1 U8905 ( .A1(n6962), .A2(n7183), .B1(n7327), .B2(n8739), .ZN(n7184)
         );
  AOI21_X1 U8906 ( .B1(n8743), .B2(n7170), .A(n7184), .ZN(n7185) );
  OAI21_X1 U8907 ( .B1(n9862), .B2(n8745), .A(n7185), .ZN(n7186) );
  AOI21_X1 U8908 ( .B1(n9865), .B2(n9753), .A(n7186), .ZN(n7187) );
  OAI21_X1 U8909 ( .B1(n7188), .B2(n8655), .A(n7187), .ZN(P2_U3284) );
  OAI222_X1 U8910 ( .A1(P2_U3152), .A2(n7904), .B1(n7949), .B2(n7190), .C1(
        n7189), .C2(n7947), .ZN(P2_U3331) );
  NAND2_X1 U8911 ( .A1(n7201), .A2(n7199), .ZN(n7197) );
  NOR2_X1 U8912 ( .A1(n6195), .A2(n7193), .ZN(n7194) );
  AOI21_X1 U8913 ( .B1(n7210), .B2(n7823), .A(n7194), .ZN(n7195) );
  XNOR2_X1 U8914 ( .A(n7195), .B(n7821), .ZN(n7198) );
  INV_X1 U8915 ( .A(n7198), .ZN(n7196) );
  INV_X1 U8916 ( .A(n7274), .ZN(n7204) );
  AND2_X1 U8917 ( .A1(n7199), .A2(n7198), .ZN(n7200) );
  NAND2_X1 U8918 ( .A1(n7201), .A2(n7200), .ZN(n7206) );
  NAND2_X1 U8919 ( .A1(n7210), .A2(n7796), .ZN(n7203) );
  NAND2_X1 U8920 ( .A1(n7820), .A2(n8997), .ZN(n7202) );
  NAND2_X1 U8921 ( .A1(n7203), .A2(n7202), .ZN(n7205) );
  NAND2_X1 U8922 ( .A1(n7206), .A2(n7205), .ZN(n7275) );
  OAI21_X1 U8923 ( .B1(n7204), .B2(n7277), .A(n8969), .ZN(n7213) );
  AOI21_X1 U8924 ( .B1(n7274), .B2(n7206), .A(n7205), .ZN(n7212) );
  AND2_X1 U8925 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n9595) );
  NOR2_X1 U8926 ( .A1(n8898), .A2(n7472), .ZN(n7207) );
  AOI211_X1 U8927 ( .C1(n8986), .C2(n9478), .A(n9595), .B(n7207), .ZN(n7208)
         );
  OAI21_X1 U8928 ( .B1(n8989), .B2(n9483), .A(n7208), .ZN(n7209) );
  AOI21_X1 U8929 ( .B1(n8991), .B2(n7210), .A(n7209), .ZN(n7211) );
  OAI21_X1 U8930 ( .B1(n7213), .B2(n7212), .A(n7211), .ZN(P1_U3239) );
  XOR2_X1 U8931 ( .A(n7214), .B(n7445), .Z(n7215) );
  AOI222_X1 U8932 ( .A1(n9651), .A2(n7215), .B1(n8997), .B2(n9656), .C1(n8998), 
        .C2(n9654), .ZN(n9494) );
  INV_X1 U8933 ( .A(n7216), .ZN(n7217) );
  OAI22_X1 U8934 ( .A1(n9666), .A2(n7218), .B1(n7217), .B2(n9663), .ZN(n7222)
         );
  INV_X1 U8935 ( .A(n7473), .ZN(n9495) );
  INV_X1 U8936 ( .A(n7219), .ZN(n7239) );
  INV_X1 U8937 ( .A(n9471), .ZN(n7220) );
  OAI211_X1 U8938 ( .C1(n9495), .C2(n7239), .A(n7220), .B(n9469), .ZN(n9493)
         );
  NOR2_X1 U8939 ( .A1(n9493), .A2(n7355), .ZN(n7221) );
  AOI211_X1 U8940 ( .C1(n9669), .C2(n7473), .A(n7222), .B(n7221), .ZN(n7230)
         );
  NAND2_X1 U8941 ( .A1(n7224), .A2(n7223), .ZN(n7231) );
  NAND2_X1 U8942 ( .A1(n7231), .A2(n7225), .ZN(n7227) );
  NAND2_X1 U8943 ( .A1(n7227), .A2(n7226), .ZN(n7228) );
  XOR2_X1 U8944 ( .A(n7445), .B(n7228), .Z(n9497) );
  NAND2_X1 U8945 ( .A1(n9497), .A2(n7360), .ZN(n7229) );
  OAI211_X1 U8946 ( .C1(n9494), .C2(n9274), .A(n7230), .B(n7229), .ZN(P1_U3277) );
  XNOR2_X1 U8947 ( .A(n7231), .B(n5893), .ZN(n7245) );
  NAND2_X1 U8948 ( .A1(n7233), .A2(n7232), .ZN(n7234) );
  AOI21_X1 U8949 ( .B1(n7235), .B2(n7234), .A(n9207), .ZN(n7238) );
  OAI22_X1 U8950 ( .A1(n7472), .A2(n9210), .B1(n7236), .B2(n9212), .ZN(n7237)
         );
  AOI211_X1 U8951 ( .C1(n7245), .C2(n9659), .A(n7238), .B(n7237), .ZN(n7259)
         );
  AOI21_X1 U8952 ( .B1(n7256), .B2(n7240), .A(n7239), .ZN(n7257) );
  INV_X1 U8953 ( .A(n7256), .ZN(n7244) );
  INV_X1 U8954 ( .A(n7241), .ZN(n7242) );
  AOI22_X1 U8955 ( .A1(n9274), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7242), .B2(
        n9484), .ZN(n7243) );
  OAI21_X1 U8956 ( .B1(n7244), .B2(n9268), .A(n7243), .ZN(n7248) );
  INV_X1 U8957 ( .A(n7245), .ZN(n7260) );
  NOR2_X1 U8958 ( .A1(n7260), .A2(n7246), .ZN(n7247) );
  AOI211_X1 U8959 ( .C1(n7257), .C2(n9277), .A(n7248), .B(n7247), .ZN(n7249)
         );
  OAI21_X1 U8960 ( .B1(n9676), .B2(n7259), .A(n7249), .ZN(P1_U3278) );
  XNOR2_X1 U8961 ( .A(n8017), .B(n7322), .ZN(n7255) );
  OAI22_X1 U8962 ( .A1(n8099), .A2(n7250), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n4992), .ZN(n7253) );
  OAI22_X1 U8963 ( .A1(n8074), .A2(n4517), .B1(n8068), .B2(n7306), .ZN(n7252)
         );
  AOI211_X1 U8964 ( .C1(n8059), .C2(n8320), .A(n7253), .B(n7252), .ZN(n7254)
         );
  OAI21_X1 U8965 ( .B1(n7255), .B2(n8103), .A(n7254), .ZN(P2_U3238) );
  AOI22_X1 U8966 ( .A1(n7257), .A2(n9469), .B1(n9345), .B2(n7256), .ZN(n7258)
         );
  OAI211_X1 U8967 ( .C1(n9389), .C2(n7260), .A(n7259), .B(n7258), .ZN(n7262)
         );
  NAND2_X1 U8968 ( .A1(n7262), .A2(n9731), .ZN(n7261) );
  OAI21_X1 U8969 ( .B1(n9731), .B2(n6841), .A(n7261), .ZN(P1_U3536) );
  NAND2_X1 U8970 ( .A1(n7262), .A2(n9722), .ZN(n7263) );
  OAI21_X1 U8971 ( .B1(n9722), .B2(n5701), .A(n7263), .ZN(P1_U3493) );
  NAND2_X1 U8972 ( .A1(n7358), .A2(n9345), .ZN(n9353) );
  NAND2_X1 U8973 ( .A1(n7358), .A2(n7823), .ZN(n7265) );
  NAND2_X1 U8974 ( .A1(n7796), .A2(n9478), .ZN(n7264) );
  NAND2_X1 U8975 ( .A1(n7265), .A2(n7264), .ZN(n7266) );
  XNOR2_X1 U8976 ( .A(n7266), .B(n7806), .ZN(n7269) );
  NOR2_X1 U8977 ( .A1(n7814), .A2(n7267), .ZN(n7268) );
  AOI21_X1 U8978 ( .B1(n7358), .B2(n7796), .A(n7268), .ZN(n7270) );
  NAND2_X1 U8979 ( .A1(n7269), .A2(n7270), .ZN(n7338) );
  INV_X1 U8980 ( .A(n7269), .ZN(n7272) );
  INV_X1 U8981 ( .A(n7270), .ZN(n7271) );
  NAND2_X1 U8982 ( .A1(n7272), .A2(n7271), .ZN(n7273) );
  AND2_X1 U8983 ( .A1(n7338), .A2(n7273), .ZN(n7276) );
  NAND3_X1 U8984 ( .A1(n7275), .A2(n7276), .A3(n7274), .ZN(n7339) );
  INV_X1 U8985 ( .A(n7339), .ZN(n7279) );
  AOI21_X1 U8986 ( .B1(n7277), .B2(n7274), .A(n7276), .ZN(n7278) );
  OAI21_X1 U8987 ( .B1(n7279), .B2(n7278), .A(n8969), .ZN(n7285) );
  INV_X1 U8988 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n7280) );
  NOR2_X1 U8989 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7280), .ZN(n9606) );
  AOI21_X1 U8990 ( .B1(n8985), .B2(n8997), .A(n9606), .ZN(n7282) );
  NAND2_X1 U8991 ( .A1(n8986), .A2(n9242), .ZN(n7281) );
  OAI211_X1 U8992 ( .C1(n8989), .C2(n7351), .A(n7282), .B(n7281), .ZN(n7283)
         );
  INV_X1 U8993 ( .A(n7283), .ZN(n7284) );
  OAI211_X1 U8994 ( .C1(n9353), .C2(n8889), .A(n7285), .B(n7284), .ZN(P1_U3224) );
  AND2_X1 U8995 ( .A1(n7322), .A2(n7320), .ZN(n7287) );
  NAND2_X1 U8996 ( .A1(n8017), .A2(n7287), .ZN(n7291) );
  INV_X1 U8997 ( .A(n7320), .ZN(n7289) );
  OR2_X1 U8998 ( .A1(n7289), .A2(n7288), .ZN(n7290) );
  NAND2_X1 U8999 ( .A1(n7291), .A2(n7290), .ZN(n7294) );
  NAND2_X1 U9000 ( .A1(n8017), .A2(n7292), .ZN(n7371) );
  AND2_X1 U9001 ( .A1(n7371), .A2(n7293), .ZN(n7363) );
  OAI211_X1 U9002 ( .C1(n7286), .C2(n7294), .A(n7363), .B(n8085), .ZN(n7298)
         );
  OAI22_X1 U9003 ( .A1(n8099), .A2(n7307), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n5047), .ZN(n7296) );
  OAI22_X1 U9004 ( .A1(n7306), .A2(n8069), .B1(n8068), .B2(n8123), .ZN(n7295)
         );
  NAND2_X1 U9005 ( .A1(n7298), .A2(n7297), .ZN(P2_U3236) );
  AND2_X1 U9006 ( .A1(n7299), .A2(n8173), .ZN(n7868) );
  NAND2_X1 U9007 ( .A1(n7881), .A2(n7868), .ZN(n7302) );
  INV_X1 U9008 ( .A(n8173), .ZN(n7301) );
  OR2_X1 U9009 ( .A1(n7919), .A2(n7365), .ZN(n8178) );
  NAND2_X1 U9010 ( .A1(n7919), .A2(n7365), .ZN(n8723) );
  NAND2_X1 U9011 ( .A1(n8178), .A2(n8723), .ZN(n8286) );
  INV_X1 U9012 ( .A(n8724), .ZN(n7303) );
  AOI21_X1 U9013 ( .B1(n7304), .B2(n8286), .A(n7303), .ZN(n7305) );
  OAI222_X1 U9014 ( .A1(n8650), .A2(n8123), .B1(n8648), .B2(n7306), .C1(n8661), 
        .C2(n7305), .ZN(n9454) );
  INV_X1 U9015 ( .A(n9454), .ZN(n7316) );
  OAI22_X1 U9016 ( .A1(n6962), .A2(n7308), .B1(n7307), .B2(n8739), .ZN(n7310)
         );
  INV_X1 U9017 ( .A(n7919), .ZN(n9452) );
  XNOR2_X1 U9018 ( .A(n7910), .B(n9452), .ZN(n9453) );
  NOR2_X1 U9019 ( .A1(n9453), .A2(n8745), .ZN(n7309) );
  AOI211_X1 U9020 ( .C1(n8743), .C2(n7919), .A(n7310), .B(n7309), .ZN(n7315)
         );
  OR2_X1 U9021 ( .A1(n7170), .A2(n8318), .ZN(n7311) );
  INV_X1 U9022 ( .A(n8286), .ZN(n8181) );
  AND2_X1 U9023 ( .A1(n7922), .A2(n8181), .ZN(n9451) );
  INV_X1 U9024 ( .A(n9451), .ZN(n7313) );
  NAND3_X1 U9025 ( .A1(n7313), .A2(n9456), .A3(n9753), .ZN(n7314) );
  OAI211_X1 U9026 ( .C1(n7316), .C2(n8655), .A(n7315), .B(n7314), .ZN(P2_U3283) );
  INV_X1 U9027 ( .A(n7317), .ZN(n7739) );
  NAND2_X1 U9028 ( .A1(n7321), .A2(n7320), .ZN(n7326) );
  NAND2_X1 U9029 ( .A1(n8017), .A2(n7322), .ZN(n7324) );
  NAND2_X1 U9030 ( .A1(n7324), .A2(n7323), .ZN(n7325) );
  XOR2_X1 U9031 ( .A(n7326), .B(n7325), .Z(n7332) );
  OAI22_X1 U9032 ( .A1(n8099), .A2(n7327), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8385), .ZN(n7330) );
  INV_X1 U9033 ( .A(n7170), .ZN(n9860) );
  OAI22_X1 U9034 ( .A1(n8074), .A2(n9860), .B1(n8069), .B2(n7328), .ZN(n7329)
         );
  AOI211_X1 U9035 ( .C1(n8058), .C2(n8731), .A(n7330), .B(n7329), .ZN(n7331)
         );
  OAI21_X1 U9036 ( .B1(n7332), .B2(n8103), .A(n7331), .ZN(P2_U3226) );
  INV_X1 U9037 ( .A(n8991), .ZN(n8961) );
  NAND2_X1 U9038 ( .A1(n9344), .A2(n7823), .ZN(n7334) );
  NAND2_X1 U9039 ( .A1(n7796), .A2(n9242), .ZN(n7333) );
  NAND2_X1 U9040 ( .A1(n7334), .A2(n7333), .ZN(n7335) );
  XNOR2_X1 U9041 ( .A(n7335), .B(n7821), .ZN(n7740) );
  NOR2_X1 U9042 ( .A1(n7814), .A2(n7336), .ZN(n7337) );
  AOI21_X1 U9043 ( .B1(n9344), .B2(n7796), .A(n7337), .ZN(n7741) );
  XNOR2_X1 U9044 ( .A(n7740), .B(n7741), .ZN(n7341) );
  NAND2_X1 U9045 ( .A1(n7339), .A2(n7338), .ZN(n7340) );
  OAI21_X1 U9046 ( .B1(n7341), .B2(n7340), .A(n7744), .ZN(n7342) );
  NAND2_X1 U9047 ( .A1(n7342), .A2(n8969), .ZN(n7347) );
  NOR2_X1 U9048 ( .A1(n8989), .A2(n9265), .ZN(n7345) );
  NAND2_X1 U9049 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n9614) );
  OAI21_X1 U9050 ( .B1(n8956), .B2(n7343), .A(n9614), .ZN(n7344) );
  AOI211_X1 U9051 ( .C1(n8985), .C2(n9478), .A(n7345), .B(n7344), .ZN(n7346)
         );
  OAI211_X1 U9052 ( .C1(n9269), .C2(n8961), .A(n7347), .B(n7346), .ZN(P1_U3226) );
  NAND3_X1 U9053 ( .A1(n9474), .A2(n7585), .A3(n7447), .ZN(n7348) );
  NAND2_X1 U9054 ( .A1(n7349), .A2(n7348), .ZN(n7350) );
  AOI222_X1 U9055 ( .A1(n9651), .A2(n7350), .B1(n9242), .B2(n9656), .C1(n8997), 
        .C2(n9654), .ZN(n9354) );
  INV_X1 U9056 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n7352) );
  OAI22_X1 U9057 ( .A1(n9666), .A2(n7352), .B1(n7351), .B2(n9663), .ZN(n7357)
         );
  INV_X1 U9058 ( .A(n7358), .ZN(n7354) );
  INV_X1 U9059 ( .A(n9470), .ZN(n7353) );
  OAI211_X1 U9060 ( .C1(n7354), .C2(n7353), .A(n4317), .B(n9469), .ZN(n9352)
         );
  NOR2_X1 U9061 ( .A1(n9352), .A2(n7355), .ZN(n7356) );
  AOI211_X1 U9062 ( .C1(n9669), .C2(n7358), .A(n7357), .B(n7356), .ZN(n7362)
         );
  XNOR2_X1 U9063 ( .A(n7359), .B(n7587), .ZN(n9351) );
  NAND2_X1 U9064 ( .A1(n9351), .A2(n7360), .ZN(n7361) );
  OAI211_X1 U9065 ( .C1(n9354), .C2(n9274), .A(n7362), .B(n7361), .ZN(P1_U3275) );
  INV_X1 U9066 ( .A(n7363), .ZN(n7367) );
  NOR3_X1 U9067 ( .A1(n8040), .A2(n7365), .A3(n7364), .ZN(n7366) );
  AOI21_X1 U9068 ( .B1(n7367), .B2(n8085), .A(n7366), .ZN(n7377) );
  AOI22_X1 U9069 ( .A1(n8058), .A2(n8728), .B1(n8059), .B2(n8731), .ZN(n7369)
         );
  OAI211_X1 U9070 ( .C1(n8099), .C2(n8740), .A(n7369), .B(n7368), .ZN(n7374)
         );
  NAND2_X1 U9071 ( .A1(n7371), .A2(n7370), .ZN(n7372) );
  NOR2_X1 U9072 ( .A1(n7372), .A2(n8103), .ZN(n7373) );
  OAI21_X1 U9073 ( .B1(n7377), .B2(n7376), .A(n7375), .ZN(P2_U3217) );
  INV_X1 U9074 ( .A(SI_28_), .ZN(n7380) );
  NAND2_X1 U9075 ( .A1(n7381), .A2(n7380), .ZN(n7382) );
  INV_X1 U9076 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n7890) );
  INV_X1 U9077 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n7707) );
  MUX2_X1 U9078 ( .A(n7890), .B(n7707), .S(n7393), .Z(n7422) );
  INV_X1 U9079 ( .A(n7422), .ZN(n7385) );
  NOR2_X1 U9080 ( .A1(n7385), .A2(SI_29_), .ZN(n7384) );
  NAND2_X1 U9081 ( .A1(n7385), .A2(SI_29_), .ZN(n7386) );
  MUX2_X1 U9082 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n7393), .Z(n7389) );
  INV_X1 U9083 ( .A(n7414), .ZN(n7388) );
  NAND2_X1 U9084 ( .A1(n7388), .A2(SI_30_), .ZN(n7392) );
  NAND2_X1 U9085 ( .A1(n7390), .A2(n7389), .ZN(n7391) );
  NAND2_X1 U9086 ( .A1(n7392), .A2(n7391), .ZN(n7396) );
  MUX2_X1 U9087 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n7393), .Z(n7394) );
  XNOR2_X1 U9088 ( .A(n7394), .B(SI_31_), .ZN(n7395) );
  INV_X1 U9089 ( .A(n8109), .ZN(n7401) );
  NOR4_X1 U9090 ( .A1(n7397), .A2(P2_IR_REG_30__SCAN_IN), .A3(n4737), .A4(
        P2_U3152), .ZN(n7398) );
  AOI21_X1 U9091 ( .B1(n7399), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n7398), .ZN(
        n7400) );
  OAI21_X1 U9092 ( .B1(n7401), .B2(n7949), .A(n7400), .ZN(P2_U3327) );
  INV_X1 U9093 ( .A(n7402), .ZN(n7405) );
  NAND3_X1 U9094 ( .A1(n7403), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n7404) );
  OAI22_X1 U9095 ( .A1(n7405), .A2(n7404), .B1(n6127), .B2(n4258), .ZN(n7406)
         );
  AOI21_X1 U9096 ( .B1(n8109), .B2(n7407), .A(n7406), .ZN(n7408) );
  INV_X1 U9097 ( .A(n7408), .ZN(P1_U3322) );
  NOR4_X1 U9098 ( .A1(n9372), .A2(n7409), .A3(n5916), .A4(n6046), .ZN(n7706)
         );
  OAI21_X1 U9099 ( .B1(n7411), .B2(n7410), .A(P1_B_REG_SCAN_IN), .ZN(n7705) );
  NAND2_X1 U9100 ( .A1(n8109), .A2(n7425), .ZN(n7413) );
  OR2_X1 U9101 ( .A1(n7426), .A2(n6127), .ZN(n7412) );
  NAND2_X1 U9102 ( .A1(n8107), .A2(n7425), .ZN(n7416) );
  INV_X1 U9103 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n7851) );
  OR2_X1 U9104 ( .A1(n7426), .A2(n7851), .ZN(n7415) );
  INV_X1 U9105 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n7421) );
  NAND2_X1 U9106 ( .A1(n7417), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n7420) );
  INV_X1 U9107 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n7418) );
  OR2_X1 U9108 ( .A1(n5549), .A2(n7418), .ZN(n7419) );
  OAI211_X1 U9109 ( .C1(n5580), .C2(n7421), .A(n7420), .B(n7419), .ZN(n8995)
         );
  NOR2_X1 U9110 ( .A1(n9287), .A2(n8995), .ZN(n7692) );
  XNOR2_X1 U9111 ( .A(n7422), .B(SI_29_), .ZN(n7423) );
  NAND2_X1 U9112 ( .A1(n7889), .A2(n7425), .ZN(n7428) );
  OR2_X1 U9113 ( .A1(n7426), .A2(n7707), .ZN(n7427) );
  INV_X1 U9114 ( .A(n8996), .ZN(n7429) );
  NAND2_X1 U9115 ( .A1(n9289), .A2(n7429), .ZN(n7512) );
  NOR2_X1 U9116 ( .A1(n7430), .A2(n7600), .ZN(n9206) );
  NAND2_X1 U9117 ( .A1(n7551), .A2(n7475), .ZN(n9648) );
  NAND4_X1 U9118 ( .A1(n7434), .A2(n7433), .A3(n7432), .A4(n7431), .ZN(n7436)
         );
  NOR3_X1 U9119 ( .A1(n7436), .A2(n7528), .A3(n7435), .ZN(n7440) );
  INV_X1 U9120 ( .A(n7437), .ZN(n7438) );
  NAND4_X1 U9121 ( .A1(n7440), .A2(n7540), .A3(n7439), .A4(n7438), .ZN(n7441)
         );
  NOR4_X1 U9122 ( .A1(n7443), .A2(n7442), .A3(n9648), .A4(n7441), .ZN(n7444)
         );
  NAND4_X1 U9123 ( .A1(n9476), .A2(n5893), .A3(n7444), .A4(n7567), .ZN(n7446)
         );
  NOR3_X1 U9124 ( .A1(n7447), .A2(n7446), .A3(n7445), .ZN(n7448) );
  AND4_X1 U9125 ( .A1(n9227), .A2(n9270), .A3(n9255), .A4(n7448), .ZN(n7449)
         );
  NAND4_X1 U9126 ( .A1(n4702), .A2(n9189), .A3(n9206), .A4(n7449), .ZN(n7450)
         );
  NOR4_X1 U9127 ( .A1(n9124), .A2(n9137), .A3(n9159), .A4(n7450), .ZN(n7454)
         );
  INV_X1 U9128 ( .A(n7451), .ZN(n7452) );
  OR2_X1 U9129 ( .A1(n7453), .A2(n7452), .ZN(n9107) );
  NAND4_X1 U9130 ( .A1(n7455), .A2(n9085), .A3(n7454), .A4(n9107), .ZN(n7456)
         );
  NOR4_X1 U9131 ( .A1(n7517), .A2(n7692), .A3(n7843), .A4(n7456), .ZN(n7460)
         );
  INV_X1 U9132 ( .A(n7712), .ZN(n7458) );
  AND2_X1 U9133 ( .A1(n9280), .A2(n7458), .ZN(n7647) );
  INV_X1 U9134 ( .A(n8995), .ZN(n7459) );
  NOR2_X1 U9135 ( .A1(n9069), .A2(n7459), .ZN(n7514) );
  NOR2_X1 U9136 ( .A1(n7647), .A2(n7514), .ZN(n7693) );
  AOI21_X1 U9137 ( .B1(n7460), .B2(n7693), .A(n7663), .ZN(n7655) );
  INV_X1 U9138 ( .A(n7655), .ZN(n7520) );
  NAND2_X1 U9139 ( .A1(n8995), .A2(n7712), .ZN(n7461) );
  NAND2_X1 U9140 ( .A1(n9069), .A2(n7461), .ZN(n7646) );
  NAND3_X1 U9141 ( .A1(n7465), .A2(n7625), .A3(n7462), .ZN(n7509) );
  AND2_X1 U9142 ( .A1(n7629), .A2(n7463), .ZN(n7624) );
  INV_X1 U9143 ( .A(n7624), .ZN(n7464) );
  AOI21_X1 U9144 ( .B1(n7465), .B2(n7464), .A(n7521), .ZN(n7466) );
  OAI21_X1 U9145 ( .B1(n7509), .B2(n7467), .A(n7466), .ZN(n7468) );
  AOI21_X1 U9146 ( .B1(n7637), .B2(n7468), .A(n4262), .ZN(n7688) );
  NAND2_X1 U9147 ( .A1(n7608), .A2(n7600), .ZN(n7469) );
  INV_X1 U9148 ( .A(n9204), .ZN(n7599) );
  NOR2_X1 U9149 ( .A1(n4278), .A2(n7599), .ZN(n7505) );
  NOR2_X1 U9150 ( .A1(n7470), .A2(n4631), .ZN(n7471) );
  AND2_X1 U9151 ( .A1(n9229), .A2(n7471), .ZN(n7504) );
  INV_X1 U9152 ( .A(n7504), .ZN(n7481) );
  INV_X1 U9153 ( .A(n7585), .ZN(n7480) );
  AND2_X1 U9154 ( .A1(n7473), .A2(n7472), .ZN(n7573) );
  INV_X1 U9155 ( .A(n7573), .ZN(n7500) );
  AND2_X1 U9156 ( .A1(n7500), .A2(n7572), .ZN(n7580) );
  INV_X1 U9157 ( .A(n7580), .ZN(n7479) );
  NAND2_X1 U9158 ( .A1(n7558), .A2(n7474), .ZN(n7570) );
  INV_X1 U9159 ( .A(n7570), .ZN(n7477) );
  NAND2_X1 U9160 ( .A1(n7557), .A2(n7475), .ZN(n7563) );
  INV_X1 U9161 ( .A(n7563), .ZN(n7476) );
  NAND4_X1 U9162 ( .A1(n7477), .A2(n7476), .A3(n9646), .A4(n7545), .ZN(n7478)
         );
  NOR4_X1 U9163 ( .A1(n7481), .A2(n7480), .A3(n7479), .A4(n7478), .ZN(n7482)
         );
  NAND2_X1 U9164 ( .A1(n7505), .A2(n7482), .ZN(n7683) );
  AND2_X1 U9165 ( .A1(n7541), .A2(n7483), .ZN(n7543) );
  INV_X1 U9166 ( .A(n7543), .ZN(n7490) );
  AND2_X1 U9167 ( .A1(n7679), .A2(n7484), .ZN(n7485) );
  NOR2_X1 U9168 ( .A1(n7490), .A2(n7485), .ZN(n7677) );
  NAND2_X1 U9169 ( .A1(n7677), .A2(n7486), .ZN(n7672) );
  NAND2_X1 U9170 ( .A1(n7487), .A2(n7671), .ZN(n7492) );
  NAND2_X1 U9171 ( .A1(n7535), .A2(n7671), .ZN(n7532) );
  AOI21_X1 U9172 ( .B1(n7675), .B2(n7533), .A(n7532), .ZN(n7489) );
  INV_X1 U9173 ( .A(n7534), .ZN(n7488) );
  NOR3_X1 U9174 ( .A1(n7489), .A2(n4324), .A3(n7488), .ZN(n7491) );
  OAI22_X1 U9175 ( .A1(n7672), .A2(n7492), .B1(n7491), .B2(n7490), .ZN(n7510)
         );
  AND2_X1 U9176 ( .A1(n9204), .A2(n9229), .ZN(n7606) );
  INV_X1 U9177 ( .A(n7593), .ZN(n7494) );
  INV_X1 U9178 ( .A(n7603), .ZN(n7493) );
  NAND2_X1 U9179 ( .A1(n7608), .A2(n7604), .ZN(n7612) );
  AOI211_X1 U9180 ( .C1(n7606), .C2(n7494), .A(n7493), .B(n7612), .ZN(n7507)
         );
  NAND2_X1 U9181 ( .A1(n7551), .A2(n7495), .ZN(n7554) );
  INV_X1 U9182 ( .A(n7554), .ZN(n7496) );
  OR2_X1 U9183 ( .A1(n7563), .A2(n7496), .ZN(n7497) );
  OAI21_X1 U9184 ( .B1(n7570), .B2(n7564), .A(n7577), .ZN(n7499) );
  AND2_X1 U9185 ( .A1(n7579), .A2(n7576), .ZN(n7574) );
  INV_X1 U9186 ( .A(n7574), .ZN(n7498) );
  AOI21_X1 U9187 ( .B1(n7572), .B2(n7499), .A(n7498), .ZN(n7502) );
  NAND2_X1 U9188 ( .A1(n7585), .A2(n7500), .ZN(n7501) );
  OAI211_X1 U9189 ( .C1(n7502), .C2(n7501), .A(n7591), .B(n7584), .ZN(n7503)
         );
  NAND3_X1 U9190 ( .A1(n7505), .A2(n7504), .A3(n7503), .ZN(n7506) );
  OAI211_X1 U9191 ( .C1(n7507), .C2(n4278), .A(n7614), .B(n7506), .ZN(n7508)
         );
  NOR2_X1 U9192 ( .A1(n7509), .A2(n7508), .ZN(n7662) );
  OAI211_X1 U9193 ( .C1(n7683), .C2(n7510), .A(n7662), .B(n7637), .ZN(n7511)
         );
  NAND2_X1 U9194 ( .A1(n7640), .A2(n7639), .ZN(n7687) );
  AOI21_X1 U9195 ( .B1(n7688), .B2(n7511), .A(n7687), .ZN(n7513) );
  INV_X1 U9196 ( .A(n7512), .ZN(n7691) );
  NOR3_X1 U9197 ( .A1(n4347), .A2(n7513), .A3(n7691), .ZN(n7518) );
  INV_X1 U9198 ( .A(n7514), .ZN(n7515) );
  NAND2_X1 U9199 ( .A1(n7515), .A2(n7712), .ZN(n7516) );
  OAI211_X1 U9200 ( .C1(n7518), .C2(n4700), .A(n7663), .B(n7694), .ZN(n7519)
         );
  INV_X1 U9201 ( .A(n7843), .ZN(n7642) );
  INV_X1 U9202 ( .A(n7521), .ZN(n7522) );
  AND2_X1 U9203 ( .A1(n7523), .A2(n7522), .ZN(n7524) );
  MUX2_X1 U9204 ( .A(n7525), .B(n7524), .S(n7547), .Z(n7633) );
  NAND2_X1 U9205 ( .A1(n7527), .A2(n7650), .ZN(n7531) );
  AOI21_X1 U9206 ( .B1(n7529), .B2(n7547), .A(n7528), .ZN(n7530) );
  NAND2_X1 U9207 ( .A1(n7531), .A2(n7530), .ZN(n7539) );
  NAND2_X1 U9208 ( .A1(n7532), .A2(n7534), .ZN(n7537) );
  NAND2_X1 U9209 ( .A1(n7534), .A2(n7533), .ZN(n7676) );
  NAND2_X1 U9210 ( .A1(n7676), .A2(n7535), .ZN(n7536) );
  MUX2_X1 U9211 ( .A(n7537), .B(n7536), .S(n7650), .Z(n7538) );
  NAND2_X1 U9212 ( .A1(n7544), .A2(n7543), .ZN(n7546) );
  NAND2_X1 U9213 ( .A1(n7546), .A2(n7545), .ZN(n7548) );
  INV_X1 U9214 ( .A(n7551), .ZN(n7553) );
  OAI22_X1 U9215 ( .A1(n7561), .A2(n7554), .B1(n7553), .B2(n7552), .ZN(n7556)
         );
  NAND2_X1 U9216 ( .A1(n7556), .A2(n7555), .ZN(n7560) );
  NAND2_X1 U9217 ( .A1(n7558), .A2(n7557), .ZN(n7559) );
  NAND2_X1 U9218 ( .A1(n7560), .A2(n4695), .ZN(n7566) );
  INV_X1 U9219 ( .A(n9646), .ZN(n7562) );
  NAND2_X1 U9220 ( .A1(n7568), .A2(n7567), .ZN(n7578) );
  NAND2_X1 U9221 ( .A1(n7570), .A2(n7569), .ZN(n7571) );
  NAND3_X1 U9222 ( .A1(n7578), .A2(n7572), .A3(n7571), .ZN(n7575) );
  AOI21_X1 U9223 ( .B1(n7575), .B2(n7574), .A(n7573), .ZN(n7583) );
  NAND3_X1 U9224 ( .A1(n7578), .A2(n7577), .A3(n7576), .ZN(n7581) );
  AOI21_X1 U9225 ( .B1(n7581), .B2(n7580), .A(n5894), .ZN(n7582) );
  INV_X1 U9226 ( .A(n9476), .ZN(n9467) );
  MUX2_X1 U9227 ( .A(n7585), .B(n7584), .S(n7650), .Z(n7586) );
  OAI211_X1 U9228 ( .C1(n7588), .C2(n9467), .A(n7587), .B(n7586), .ZN(n7589)
         );
  INV_X1 U9229 ( .A(n7589), .ZN(n7597) );
  MUX2_X1 U9230 ( .A(n7591), .B(n7590), .S(n7650), .Z(n7592) );
  AND2_X1 U9231 ( .A1(n9229), .A2(n5898), .ZN(n7594) );
  MUX2_X1 U9232 ( .A(n7594), .B(n7593), .S(n7650), .Z(n7595) );
  AND2_X1 U9233 ( .A1(n7603), .A2(n7598), .ZN(n7602) );
  OR2_X1 U9234 ( .A1(n7600), .A2(n7599), .ZN(n7601) );
  NAND2_X1 U9235 ( .A1(n7604), .A2(n7603), .ZN(n7605) );
  AOI21_X1 U9236 ( .B1(n7613), .B2(n7608), .A(n4278), .ZN(n7609) );
  INV_X1 U9237 ( .A(n7609), .ZN(n7610) );
  AOI22_X1 U9238 ( .A1(n7610), .A2(n7614), .B1(n9313), .B2(n7622), .ZN(n7619)
         );
  AND2_X1 U9239 ( .A1(n7622), .A2(n9176), .ZN(n7615) );
  AOI21_X1 U9240 ( .B1(n7617), .B2(n7616), .A(n7615), .ZN(n7618) );
  MUX2_X1 U9241 ( .A(n7619), .B(n7618), .S(n7547), .Z(n7621) );
  INV_X1 U9242 ( .A(n9137), .ZN(n7620) );
  AND2_X1 U9243 ( .A1(n7621), .A2(n7620), .ZN(n7632) );
  INV_X1 U9244 ( .A(n9313), .ZN(n9156) );
  INV_X1 U9245 ( .A(n7622), .ZN(n7623) );
  OR2_X1 U9246 ( .A1(n9137), .A2(n7623), .ZN(n7626) );
  OAI21_X1 U9247 ( .B1(n9156), .B2(n7626), .A(n7624), .ZN(n7628) );
  OAI211_X1 U9248 ( .C1(n7626), .C2(n8943), .A(n9128), .B(n7625), .ZN(n7627)
         );
  MUX2_X1 U9249 ( .A(n7628), .B(n7627), .S(n7650), .Z(n7631) );
  MUX2_X1 U9250 ( .A(n9128), .B(n7629), .S(n7650), .Z(n7630) );
  NAND2_X1 U9251 ( .A1(n7639), .A2(n7637), .ZN(n7841) );
  INV_X1 U9252 ( .A(n7841), .ZN(n7634) );
  NAND2_X1 U9253 ( .A1(n7638), .A2(n7634), .ZN(n7635) );
  NAND2_X1 U9254 ( .A1(n7635), .A2(n7840), .ZN(n7636) );
  AOI21_X1 U9255 ( .B1(n7642), .B2(n7636), .A(n7691), .ZN(n7645) );
  INV_X1 U9256 ( .A(n7637), .ZN(n7685) );
  INV_X1 U9257 ( .A(n7640), .ZN(n7641) );
  AOI21_X1 U9258 ( .B1(n7643), .B2(n7642), .A(n7641), .ZN(n7644) );
  OAI21_X1 U9259 ( .B1(n7547), .B2(n7646), .A(n7694), .ZN(n7649) );
  INV_X1 U9260 ( .A(n7647), .ZN(n7648) );
  NAND2_X1 U9261 ( .A1(n7649), .A2(n7648), .ZN(n7652) );
  INV_X1 U9262 ( .A(n7654), .ZN(n7656) );
  AOI21_X1 U9263 ( .B1(n7658), .B2(n7656), .A(n7655), .ZN(n7657) );
  INV_X1 U9264 ( .A(n7658), .ZN(n7660) );
  NAND4_X1 U9265 ( .A1(n7660), .A2(n7663), .A3(n7694), .A4(n7659), .ZN(n7661)
         );
  INV_X1 U9266 ( .A(n7662), .ZN(n7686) );
  OAI21_X1 U9267 ( .B1(n7665), .B2(n7664), .A(n7663), .ZN(n7667) );
  OAI21_X1 U9268 ( .B1(n7668), .B2(n7667), .A(n7666), .ZN(n7670) );
  OAI22_X1 U9269 ( .A1(n6255), .A2(n7670), .B1(n7669), .B2(n5547), .ZN(n7674)
         );
  INV_X1 U9270 ( .A(n7671), .ZN(n7673) );
  AOI211_X1 U9271 ( .C1(n7675), .C2(n7674), .A(n7673), .B(n7672), .ZN(n7682)
         );
  INV_X1 U9272 ( .A(n7676), .ZN(n7680) );
  INV_X1 U9273 ( .A(n7677), .ZN(n7678) );
  AOI21_X1 U9274 ( .B1(n7680), .B2(n7679), .A(n7678), .ZN(n7681) );
  NOR3_X1 U9275 ( .A1(n7683), .A2(n7682), .A3(n7681), .ZN(n7684) );
  OR3_X1 U9276 ( .A1(n7686), .A2(n7685), .A3(n7684), .ZN(n7689) );
  AOI21_X1 U9277 ( .B1(n7689), .B2(n7688), .A(n7687), .ZN(n7690) );
  NOR3_X1 U9278 ( .A1(n7692), .A2(n7691), .A3(n7690), .ZN(n7696) );
  INV_X1 U9279 ( .A(n7693), .ZN(n7695) );
  OAI21_X1 U9280 ( .B1(n7696), .B2(n7695), .A(n7694), .ZN(n7698) );
  NAND2_X1 U9281 ( .A1(n7698), .A2(n9473), .ZN(n7702) );
  INV_X1 U9282 ( .A(n7703), .ZN(n7704) );
  INV_X1 U9283 ( .A(n7889), .ZN(n7866) );
  OAI222_X1 U9284 ( .A1(n7850), .A2(n7866), .B1(n7708), .B2(P1_U3084), .C1(
        n7707), .C2(n4258), .ZN(P1_U3324) );
  NAND2_X1 U9285 ( .A1(n9287), .A2(n9067), .ZN(n9283) );
  XNOR2_X1 U9286 ( .A(n9280), .B(n9283), .ZN(n9282) );
  NOR2_X1 U9287 ( .A1(n9666), .A2(n7709), .ZN(n7713) );
  INV_X1 U9288 ( .A(P1_B_REG_SCAN_IN), .ZN(n7710) );
  NOR2_X1 U9289 ( .A1(n6046), .A2(n7710), .ZN(n7711) );
  NOR2_X1 U9290 ( .A1(n9210), .A2(n7711), .ZN(n7844) );
  NAND2_X1 U9291 ( .A1(n7844), .A2(n7712), .ZN(n9285) );
  NOR2_X1 U9292 ( .A1(n9274), .A2(n9285), .ZN(n9070) );
  AOI211_X1 U9293 ( .C1(n9280), .C2(n9669), .A(n7713), .B(n9070), .ZN(n7714)
         );
  OAI21_X1 U9294 ( .B1(n9282), .B2(n9671), .A(n7714), .ZN(P1_U3261) );
  INV_X1 U9295 ( .A(n7917), .ZN(n9442) );
  INV_X1 U9296 ( .A(n8040), .ZN(n8077) );
  NAND2_X1 U9297 ( .A1(n8077), .A2(n8728), .ZN(n7720) );
  NAND2_X1 U9298 ( .A1(n8085), .A2(n8004), .ZN(n7719) );
  NAND2_X1 U9299 ( .A1(n8017), .A2(n7715), .ZN(n7717) );
  XNOR2_X1 U9300 ( .A(n8002), .B(n7718), .ZN(n8005) );
  MUX2_X1 U9301 ( .A(n7720), .B(n7719), .S(n8005), .Z(n7726) );
  INV_X1 U9302 ( .A(n8714), .ZN(n7724) );
  INV_X1 U9303 ( .A(n7882), .ZN(n8317) );
  NAND2_X1 U9304 ( .A1(n8317), .A2(n8729), .ZN(n7722) );
  NAND2_X1 U9305 ( .A1(n4663), .A2(n8730), .ZN(n7721) );
  AND2_X1 U9306 ( .A1(n7722), .A2(n7721), .ZN(n8709) );
  OAI22_X1 U9307 ( .A1(n7998), .A2(n8709), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10008), .ZN(n7723) );
  AOI21_X1 U9308 ( .B1(n7724), .B2(n8079), .A(n7723), .ZN(n7725) );
  OAI211_X1 U9309 ( .C1(n9442), .C2(n8074), .A(n7726), .B(n7725), .ZN(P2_U3243) );
  INV_X1 U9310 ( .A(n8831), .ZN(n8644) );
  AND2_X1 U9311 ( .A1(n7728), .A2(n7727), .ZN(n8020) );
  INV_X1 U9312 ( .A(n7729), .ZN(n7730) );
  AOI21_X1 U9313 ( .B1(n8020), .B2(n7730), .A(n8103), .ZN(n7733) );
  NOR3_X1 U9314 ( .A1(n7731), .A2(n8649), .A3(n8040), .ZN(n7732) );
  OAI21_X1 U9315 ( .B1(n7733), .B2(n7732), .A(n7854), .ZN(n7738) );
  INV_X1 U9316 ( .A(n7734), .ZN(n8642) );
  NOR2_X1 U9317 ( .A1(n7735), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8438) );
  OAI22_X1 U9318 ( .A1(n8649), .A2(n8069), .B1(n8068), .B2(n8651), .ZN(n7736)
         );
  AOI211_X1 U9319 ( .C1(n8079), .C2(n8642), .A(n8438), .B(n7736), .ZN(n7737)
         );
  OAI211_X1 U9320 ( .C1(n8644), .C2(n8074), .A(n7738), .B(n7737), .ZN(P2_U3240) );
  OAI222_X1 U9321 ( .A1(n7850), .A2(n7739), .B1(n5916), .B2(P1_U3084), .C1(
        n10046), .C2(n4258), .ZN(P1_U3325) );
  INV_X1 U9322 ( .A(n7740), .ZN(n7742) );
  NAND2_X1 U9323 ( .A1(n7742), .A2(n7741), .ZN(n7743) );
  NAND2_X1 U9324 ( .A1(n9251), .A2(n7823), .ZN(n7746) );
  NAND2_X1 U9325 ( .A1(n9272), .A2(n7796), .ZN(n7745) );
  NAND2_X1 U9326 ( .A1(n7746), .A2(n7745), .ZN(n7747) );
  XNOR2_X1 U9327 ( .A(n7747), .B(n7806), .ZN(n7750) );
  AND2_X1 U9328 ( .A1(n7820), .A2(n9272), .ZN(n7749) );
  AOI21_X1 U9329 ( .B1(n9251), .B2(n7796), .A(n7749), .ZN(n8951) );
  NAND2_X1 U9330 ( .A1(n8953), .A2(n8951), .ZN(n8950) );
  NAND2_X1 U9331 ( .A1(n7751), .A2(n7750), .ZN(n8952) );
  NAND2_X1 U9332 ( .A1(n9334), .A2(n7823), .ZN(n7753) );
  NAND2_X1 U9333 ( .A1(n9243), .A2(n7796), .ZN(n7752) );
  NAND2_X1 U9334 ( .A1(n7753), .A2(n7752), .ZN(n7754) );
  XNOR2_X1 U9335 ( .A(n7754), .B(n7821), .ZN(n7756) );
  AND2_X1 U9336 ( .A1(n9243), .A2(n7820), .ZN(n7755) );
  AOI21_X1 U9337 ( .B1(n9334), .B2(n7796), .A(n7755), .ZN(n7757) );
  XNOR2_X1 U9338 ( .A(n7756), .B(n7757), .ZN(n8879) );
  INV_X1 U9339 ( .A(n7756), .ZN(n7758) );
  NAND2_X1 U9340 ( .A1(n7758), .A2(n7757), .ZN(n7759) );
  NAND2_X1 U9341 ( .A1(n8878), .A2(n7759), .ZN(n8928) );
  NAND2_X1 U9342 ( .A1(n9331), .A2(n7823), .ZN(n7761) );
  NAND2_X1 U9343 ( .A1(n9233), .A2(n7796), .ZN(n7760) );
  NAND2_X1 U9344 ( .A1(n7761), .A2(n7760), .ZN(n7762) );
  XNOR2_X1 U9345 ( .A(n7762), .B(n7821), .ZN(n7765) );
  NAND2_X1 U9346 ( .A1(n9331), .A2(n7796), .ZN(n7764) );
  NAND2_X1 U9347 ( .A1(n9233), .A2(n7820), .ZN(n7763) );
  NAND2_X1 U9348 ( .A1(n7764), .A2(n7763), .ZN(n7766) );
  NAND2_X1 U9349 ( .A1(n7765), .A2(n7766), .ZN(n8929) );
  INV_X1 U9350 ( .A(n7765), .ZN(n7768) );
  INV_X1 U9351 ( .A(n7766), .ZN(n7767) );
  NAND2_X1 U9352 ( .A1(n7768), .A2(n7767), .ZN(n8931) );
  NAND2_X1 U9353 ( .A1(n9195), .A2(n7823), .ZN(n7770) );
  NAND2_X1 U9354 ( .A1(n9175), .A2(n7796), .ZN(n7769) );
  NAND2_X1 U9355 ( .A1(n7770), .A2(n7769), .ZN(n7771) );
  XNOR2_X1 U9356 ( .A(n7771), .B(n7821), .ZN(n7773) );
  AND2_X1 U9357 ( .A1(n9175), .A2(n7820), .ZN(n7772) );
  AOI21_X1 U9358 ( .B1(n9195), .B2(n7796), .A(n7772), .ZN(n7774) );
  XNOR2_X1 U9359 ( .A(n7773), .B(n7774), .ZN(n8885) );
  INV_X1 U9360 ( .A(n7773), .ZN(n7775) );
  AND2_X1 U9361 ( .A1(n9190), .A2(n7820), .ZN(n7776) );
  AOI21_X1 U9362 ( .B1(n9318), .B2(n7796), .A(n7776), .ZN(n7781) );
  NAND2_X1 U9363 ( .A1(n7780), .A2(n7781), .ZN(n8938) );
  NAND2_X1 U9364 ( .A1(n9318), .A2(n7823), .ZN(n7778) );
  NAND2_X1 U9365 ( .A1(n9190), .A2(n7796), .ZN(n7777) );
  NAND2_X1 U9366 ( .A1(n7778), .A2(n7777), .ZN(n7779) );
  XNOR2_X1 U9367 ( .A(n7779), .B(n7821), .ZN(n8941) );
  INV_X1 U9368 ( .A(n7780), .ZN(n7783) );
  INV_X1 U9369 ( .A(n7781), .ZN(n7782) );
  NAND2_X1 U9370 ( .A1(n9313), .A2(n7823), .ZN(n7785) );
  NAND2_X1 U9371 ( .A1(n9176), .A2(n7796), .ZN(n7784) );
  NAND2_X1 U9372 ( .A1(n7785), .A2(n7784), .ZN(n7786) );
  XNOR2_X1 U9373 ( .A(n7786), .B(n7821), .ZN(n7788) );
  AND2_X1 U9374 ( .A1(n9176), .A2(n7820), .ZN(n7787) );
  AOI21_X1 U9375 ( .B1(n9313), .B2(n7796), .A(n7787), .ZN(n8868) );
  INV_X1 U9376 ( .A(n7788), .ZN(n7789) );
  OAI22_X1 U9377 ( .A1(n8913), .A2(n6195), .B1(n8899), .B2(n7814), .ZN(n7793)
         );
  NAND2_X1 U9378 ( .A1(n9309), .A2(n7823), .ZN(n7791) );
  NAND2_X1 U9379 ( .A1(n9162), .A2(n7796), .ZN(n7790) );
  NAND2_X1 U9380 ( .A1(n7791), .A2(n7790), .ZN(n7792) );
  XNOR2_X1 U9381 ( .A(n7792), .B(n7821), .ZN(n7794) );
  XOR2_X1 U9382 ( .A(n7793), .B(n7794), .Z(n8905) );
  NAND2_X1 U9383 ( .A1(n8904), .A2(n8905), .ZN(n8903) );
  INV_X1 U9384 ( .A(n9303), .ZN(n9122) );
  OAI22_X1 U9385 ( .A1(n9122), .A2(n6195), .B1(n8908), .B2(n7814), .ZN(n7801)
         );
  NAND2_X1 U9386 ( .A1(n9303), .A2(n7823), .ZN(n7798) );
  NAND2_X1 U9387 ( .A1(n9141), .A2(n7796), .ZN(n7797) );
  NAND2_X1 U9388 ( .A1(n7798), .A2(n7797), .ZN(n7799) );
  XNOR2_X1 U9389 ( .A(n7799), .B(n7821), .ZN(n7800) );
  XOR2_X1 U9390 ( .A(n7801), .B(n7800), .Z(n8895) );
  INV_X1 U9391 ( .A(n7800), .ZN(n7803) );
  INV_X1 U9392 ( .A(n7801), .ZN(n7802) );
  NAND2_X1 U9393 ( .A1(n9299), .A2(n7823), .ZN(n7805) );
  OR2_X1 U9394 ( .A1(n6195), .A2(n9123), .ZN(n7804) );
  NAND2_X1 U9395 ( .A1(n7805), .A2(n7804), .ZN(n7807) );
  XNOR2_X1 U9396 ( .A(n7807), .B(n7806), .ZN(n7810) );
  NOR2_X1 U9397 ( .A1(n7814), .A2(n9123), .ZN(n7808) );
  AOI21_X1 U9398 ( .B1(n9299), .B2(n7796), .A(n7808), .ZN(n7809) );
  NOR2_X1 U9399 ( .A1(n7810), .A2(n7809), .ZN(n8982) );
  NAND2_X1 U9400 ( .A1(n7810), .A2(n7809), .ZN(n8980) );
  NOR2_X1 U9401 ( .A1(n6195), .A2(n7813), .ZN(n7811) );
  AOI21_X1 U9402 ( .B1(n9295), .B2(n7823), .A(n7811), .ZN(n7812) );
  XNOR2_X1 U9403 ( .A(n7812), .B(n7821), .ZN(n7817) );
  NOR2_X1 U9404 ( .A1(n7814), .A2(n7813), .ZN(n7815) );
  AOI21_X1 U9405 ( .B1(n9295), .B2(n7796), .A(n7815), .ZN(n7816) );
  NAND2_X1 U9406 ( .A1(n7817), .A2(n7816), .ZN(n7819) );
  OAI21_X1 U9407 ( .B1(n7817), .B2(n7816), .A(n7819), .ZN(n7818) );
  INV_X1 U9408 ( .A(n7818), .ZN(n8858) );
  AOI22_X1 U9409 ( .A1(n9077), .A2(n7796), .B1(n7820), .B2(n9087), .ZN(n7822)
         );
  XNOR2_X1 U9410 ( .A(n7822), .B(n7821), .ZN(n7825) );
  AOI22_X1 U9411 ( .A1(n9077), .A2(n7823), .B1(n7796), .B2(n9087), .ZN(n7824)
         );
  XNOR2_X1 U9412 ( .A(n7825), .B(n7824), .ZN(n7826) );
  XNOR2_X1 U9413 ( .A(n7827), .B(n7826), .ZN(n7832) );
  AOI22_X1 U9414 ( .A1(n8985), .A2(n9108), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n7829) );
  NAND2_X1 U9415 ( .A1(n8986), .A2(n8996), .ZN(n7828) );
  OAI211_X1 U9416 ( .C1(n8989), .C2(n9074), .A(n7829), .B(n7828), .ZN(n7830)
         );
  AOI21_X1 U9417 ( .B1(n9077), .B2(n8991), .A(n7830), .ZN(n7831) );
  OAI21_X1 U9418 ( .B1(n7832), .B2(n8993), .A(n7831), .ZN(P1_U3218) );
  XNOR2_X1 U9419 ( .A(n7834), .B(n7642), .ZN(n9292) );
  NOR2_X1 U9420 ( .A1(n9274), .A2(n9473), .ZN(n9248) );
  INV_X1 U9421 ( .A(n9289), .ZN(n7839) );
  INV_X1 U9422 ( .A(n7836), .ZN(n7837) );
  AOI22_X1 U9423 ( .A1(n9676), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n7837), .B2(
        n9484), .ZN(n7838) );
  OAI21_X1 U9424 ( .B1(n7839), .B2(n9268), .A(n7838), .ZN(n7847) );
  INV_X1 U9425 ( .A(n7844), .ZN(n7845) );
  NOR2_X1 U9426 ( .A1(n9290), .A2(n9274), .ZN(n7846) );
  OAI21_X1 U9427 ( .B1(n9292), .B2(n9279), .A(n7848), .ZN(P1_U3355) );
  INV_X1 U9428 ( .A(n8107), .ZN(n7948) );
  OAI222_X1 U9429 ( .A1(n4258), .A2(n7851), .B1(n7850), .B2(n7948), .C1(
        P1_U3084), .C2(n7849), .ZN(P1_U3323) );
  INV_X1 U9430 ( .A(n7930), .ZN(n8316) );
  NAND3_X1 U9431 ( .A1(n7852), .A2(n8077), .A3(n8316), .ZN(n7853) );
  OAI21_X1 U9432 ( .B1(n7854), .B2(n8103), .A(n7853), .ZN(n7857) );
  INV_X1 U9433 ( .A(n7855), .ZN(n7856) );
  NAND2_X1 U9434 ( .A1(n7857), .A2(n7856), .ZN(n7864) );
  NOR2_X1 U9435 ( .A1(n8099), .A2(n8634), .ZN(n7862) );
  INV_X1 U9436 ( .A(n7984), .ZN(n8600) );
  NAND2_X1 U9437 ( .A1(n8600), .A2(n8729), .ZN(n7859) );
  NAND2_X1 U9438 ( .A1(n8316), .A2(n8730), .ZN(n7858) );
  AND2_X1 U9439 ( .A1(n7859), .A2(n7858), .ZN(n8627) );
  OAI22_X1 U9440 ( .A1(n7998), .A2(n8627), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7860), .ZN(n7861) );
  AOI211_X1 U9441 ( .C1(n8824), .C2(n8101), .A(n7862), .B(n7861), .ZN(n7863)
         );
  OAI211_X1 U9442 ( .C1(n8103), .C2(n7865), .A(n7864), .B(n7863), .ZN(P2_U3221) );
  OAI222_X1 U9443 ( .A1(n7947), .A2(n7890), .B1(n7949), .B2(n7866), .C1(
        P2_U3152), .C2(n4728), .ZN(P2_U3329) );
  INV_X1 U9444 ( .A(n8705), .ZN(n7873) );
  OR2_X1 U9445 ( .A1(n8286), .A2(n7873), .ZN(n7870) );
  INV_X1 U9446 ( .A(n7870), .ZN(n7867) );
  AND2_X1 U9447 ( .A1(n7868), .A2(n7867), .ZN(n8701) );
  NAND2_X1 U9448 ( .A1(n9442), .A2(n8728), .ZN(n7877) );
  AND2_X1 U9449 ( .A1(n8701), .A2(n7877), .ZN(n7880) );
  NAND2_X1 U9450 ( .A1(n7871), .A2(n8123), .ZN(n7872) );
  NAND2_X1 U9451 ( .A1(n7875), .A2(n7874), .ZN(n7876) );
  INV_X1 U9452 ( .A(n7877), .ZN(n7878) );
  NOR2_X1 U9453 ( .A1(n8702), .A2(n7878), .ZN(n7879) );
  NAND2_X1 U9454 ( .A1(n8693), .A2(n7882), .ZN(n8189) );
  NAND2_X1 U9455 ( .A1(n8190), .A2(n8189), .ZN(n8682) );
  OAI21_X1 U9456 ( .B1(n8681), .B2(n8682), .A(n8189), .ZN(n8659) );
  INV_X1 U9457 ( .A(n8659), .ZN(n7884) );
  NAND2_X1 U9458 ( .A1(n8675), .A2(n8649), .ZN(n8194) );
  INV_X1 U9459 ( .A(n8670), .ZN(n7883) );
  NAND2_X1 U9460 ( .A1(n7884), .A2(n7883), .ZN(n7885) );
  OR2_X1 U9461 ( .A1(n8831), .A2(n7930), .ZN(n8623) );
  NAND2_X1 U9462 ( .A1(n8831), .A2(n7930), .ZN(n8209) );
  OR2_X1 U9463 ( .A1(n8824), .A2(n8651), .ZN(n8199) );
  NAND2_X1 U9464 ( .A1(n8824), .A2(n8651), .ZN(n8211) );
  NAND2_X1 U9465 ( .A1(n8199), .A2(n8211), .ZN(n8624) );
  INV_X1 U9466 ( .A(n8623), .ZN(n8200) );
  NOR2_X1 U9467 ( .A1(n8624), .A2(n8200), .ZN(n7886) );
  INV_X1 U9468 ( .A(n8211), .ZN(n8201) );
  NAND2_X1 U9469 ( .A1(n8613), .A2(n7984), .ZN(n8212) );
  NAND2_X1 U9470 ( .A1(n8604), .A2(n8214), .ZN(n8596) );
  XNOR2_X1 U9471 ( .A(n8812), .B(n8580), .ZN(n8597) );
  NAND2_X1 U9472 ( .A1(n8812), .A2(n8580), .ZN(n8217) );
  NAND2_X1 U9473 ( .A1(n8576), .A2(n8599), .ZN(n8205) );
  INV_X1 U9474 ( .A(n8599), .ZN(n7985) );
  NAND2_X1 U9475 ( .A1(n8807), .A2(n7985), .ZN(n8219) );
  NAND2_X1 U9476 ( .A1(n8205), .A2(n8219), .ZN(n8577) );
  INV_X1 U9477 ( .A(n8205), .ZN(n8556) );
  NAND2_X1 U9478 ( .A1(n8563), .A2(n8315), .ZN(n8224) );
  INV_X1 U9479 ( .A(n8315), .ZN(n8579) );
  NAND2_X1 U9480 ( .A1(n8802), .A2(n8579), .ZN(n8223) );
  NAND2_X1 U9481 ( .A1(n8224), .A2(n8223), .ZN(n8565) );
  NAND2_X1 U9482 ( .A1(n8550), .A2(n8031), .ZN(n8227) );
  NAND2_X1 U9483 ( .A1(n8543), .A2(n8542), .ZN(n8541) );
  NAND2_X1 U9484 ( .A1(n8541), .A2(n8228), .ZN(n8527) );
  NAND2_X1 U9485 ( .A1(n8534), .A2(n8095), .ZN(n8235) );
  NAND2_X1 U9486 ( .A1(n8527), .A2(n8528), .ZN(n8526) );
  NAND2_X1 U9487 ( .A1(n8786), .A2(n7955), .ZN(n8236) );
  INV_X1 U9488 ( .A(n8505), .ZN(n7887) );
  NOR2_X1 U9489 ( .A1(n8518), .A2(n7887), .ZN(n7888) );
  INV_X1 U9490 ( .A(n8236), .ZN(n8232) );
  NAND2_X1 U9491 ( .A1(n8779), .A2(n8096), .ZN(n8244) );
  NAND2_X1 U9492 ( .A1(n8488), .A2(n8487), .ZN(n8486) );
  NAND2_X1 U9493 ( .A1(n8773), .A2(n7954), .ZN(n8248) );
  NAND2_X1 U9494 ( .A1(n7889), .A2(n8108), .ZN(n7892) );
  OR2_X1 U9495 ( .A1(n8110), .A2(n7890), .ZN(n7891) );
  INV_X1 U9496 ( .A(n7915), .ZN(n8767) );
  INV_X1 U9497 ( .A(n8251), .ZN(n8249) );
  NAND2_X1 U9498 ( .A1(n8255), .A2(n8249), .ZN(n8296) );
  XNOR2_X1 U9499 ( .A(n8105), .B(n7894), .ZN(n7909) );
  INV_X1 U9500 ( .A(n7954), .ZN(n8490) );
  INV_X1 U9501 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n7895) );
  OR2_X1 U9502 ( .A1(n4260), .A2(n7895), .ZN(n7902) );
  INV_X1 U9503 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n7896) );
  OR2_X1 U9504 ( .A1(n7897), .A2(n7896), .ZN(n7901) );
  INV_X1 U9505 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n7898) );
  OR2_X1 U9506 ( .A1(n7899), .A2(n7898), .ZN(n7900) );
  AND3_X1 U9507 ( .A1(n7902), .A2(n7901), .A3(n7900), .ZN(n8114) );
  INV_X1 U9508 ( .A(n8114), .ZN(n8313) );
  INV_X1 U9509 ( .A(P2_B_REG_SCAN_IN), .ZN(n7903) );
  NOR2_X1 U9510 ( .A1(n7904), .A2(n7903), .ZN(n7905) );
  NOR2_X1 U9511 ( .A1(n8650), .A2(n7905), .ZN(n8461) );
  NAND2_X1 U9512 ( .A1(n8313), .A2(n8461), .ZN(n7906) );
  OR2_X1 U9513 ( .A1(n8477), .A2(n7915), .ZN(n7911) );
  INV_X1 U9514 ( .A(n7912), .ZN(n7913) );
  AOI22_X1 U9515 ( .A1(n8655), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n7913), .B2(
        n9750), .ZN(n7914) );
  OAI21_X1 U9516 ( .B1(n7915), .B2(n9758), .A(n7914), .ZN(n7916) );
  AOI21_X1 U9517 ( .B1(n8768), .B2(n9755), .A(n7916), .ZN(n7946) );
  OR2_X1 U9518 ( .A1(n7917), .A2(n8728), .ZN(n7924) );
  INV_X1 U9519 ( .A(n7924), .ZN(n7918) );
  OR2_X1 U9520 ( .A1(n7918), .A2(n8706), .ZN(n7926) );
  AND2_X1 U9521 ( .A1(n4662), .A2(n7926), .ZN(n8688) );
  NAND2_X1 U9522 ( .A1(n8693), .A2(n8317), .ZN(n7923) );
  AND2_X1 U9523 ( .A1(n8688), .A2(n7923), .ZN(n8664) );
  AND2_X1 U9524 ( .A1(n8664), .A2(n8670), .ZN(n7920) );
  NAND2_X1 U9525 ( .A1(n7919), .A2(n8731), .ZN(n8663) );
  AND2_X1 U9526 ( .A1(n7920), .A2(n8663), .ZN(n7921) );
  INV_X1 U9527 ( .A(n7923), .ZN(n7927) );
  OR2_X1 U9528 ( .A1(n7871), .A2(n4663), .ZN(n8699) );
  NAND2_X1 U9529 ( .A1(n8699), .A2(n7924), .ZN(n7925) );
  NAND2_X1 U9530 ( .A1(n7926), .A2(n7925), .ZN(n8690) );
  OR2_X1 U9531 ( .A1(n8665), .A2(n7883), .ZN(n8667) );
  INV_X1 U9532 ( .A(n8649), .ZN(n8683) );
  OR2_X1 U9533 ( .A1(n8675), .A2(n8683), .ZN(n7928) );
  AND2_X1 U9534 ( .A1(n8667), .A2(n7928), .ZN(n7929) );
  NAND2_X1 U9535 ( .A1(n8668), .A2(n7929), .ZN(n8640) );
  NOR2_X1 U9536 ( .A1(n8831), .A2(n8316), .ZN(n7931) );
  OR2_X1 U9537 ( .A1(n8824), .A2(n8608), .ZN(n7932) );
  OR2_X1 U9538 ( .A1(n8812), .A2(n8607), .ZN(n7935) );
  AND2_X1 U9539 ( .A1(n8616), .A2(n7935), .ZN(n7934) );
  INV_X1 U9540 ( .A(n7935), .ZN(n7936) );
  NAND2_X1 U9541 ( .A1(n8613), .A2(n8600), .ZN(n8586) );
  OR2_X1 U9542 ( .A1(n7936), .A2(n8586), .ZN(n7938) );
  NAND2_X1 U9543 ( .A1(n8812), .A2(n8607), .ZN(n7937) );
  AND2_X1 U9544 ( .A1(n7938), .A2(n7937), .ZN(n7939) );
  NAND2_X1 U9545 ( .A1(n7940), .A2(n7939), .ZN(n8570) );
  INV_X1 U9546 ( .A(n8031), .ZN(n8314) );
  OAI22_X1 U9547 ( .A1(n8540), .A2(n8542), .B1(n8314), .B2(n8550), .ZN(n8523)
         );
  NAND2_X1 U9548 ( .A1(n8523), .A2(n8522), .ZN(n8525) );
  INV_X1 U9549 ( .A(n8095), .ZN(n8544) );
  NAND2_X1 U9550 ( .A1(n8525), .A2(n7941), .ZN(n8519) );
  NAND2_X1 U9551 ( .A1(n8519), .A2(n8518), .ZN(n8517) );
  INV_X1 U9552 ( .A(n7955), .ZN(n8489) );
  NAND2_X1 U9553 ( .A1(n8517), .A2(n7942), .ZN(n8502) );
  NAND2_X1 U9554 ( .A1(n8500), .A2(n7943), .ZN(n8483) );
  NAND2_X1 U9555 ( .A1(n8483), .A2(n4667), .ZN(n8482) );
  INV_X1 U9556 ( .A(n8771), .ZN(n7944) );
  NAND2_X1 U9557 ( .A1(n7944), .A2(n9753), .ZN(n7945) );
  OAI211_X1 U9558 ( .C1(n8770), .C2(n8655), .A(n7946), .B(n7945), .ZN(P2_U3267) );
  INV_X1 U9559 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n9997) );
  OAI222_X1 U9560 ( .A1(n7950), .A2(P2_U3152), .B1(n7949), .B2(n7948), .C1(
        n9997), .C2(n7947), .ZN(P2_U3328) );
  XNOR2_X1 U9561 ( .A(n7951), .B(n7952), .ZN(n7959) );
  OAI22_X1 U9562 ( .A1(n8099), .A2(n8495), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7953), .ZN(n7957) );
  OAI22_X1 U9563 ( .A1(n7955), .A2(n8069), .B1(n8068), .B2(n7954), .ZN(n7956)
         );
  AOI211_X1 U9564 ( .C1(n8779), .C2(n8101), .A(n7957), .B(n7956), .ZN(n7958)
         );
  OAI21_X1 U9565 ( .B1(n7959), .B2(n8103), .A(n7958), .ZN(P2_U3216) );
  INV_X1 U9566 ( .A(n7962), .ZN(n7961) );
  NOR2_X1 U9567 ( .A1(n7961), .A2(n7960), .ZN(n8028) );
  AOI22_X1 U9568 ( .A1(n7962), .A2(n8085), .B1(n8077), .B2(n8315), .ZN(n7967)
         );
  INV_X1 U9569 ( .A(n8561), .ZN(n7964) );
  OAI22_X1 U9570 ( .A1(n8031), .A2(n8650), .B1(n7985), .B2(n8648), .ZN(n8558)
         );
  AOI22_X1 U9571 ( .A1(n8097), .A2(n8558), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n7963) );
  OAI21_X1 U9572 ( .B1(n7964), .B2(n8099), .A(n7963), .ZN(n7965) );
  AOI21_X1 U9573 ( .B1(n8802), .B2(n8101), .A(n7965), .ZN(n7966) );
  OAI21_X1 U9574 ( .B1(n8028), .B2(n7967), .A(n7966), .ZN(P2_U3218) );
  NOR3_X1 U9575 ( .A1(n8040), .A2(n7969), .A3(n7968), .ZN(n7973) );
  AOI21_X1 U9576 ( .B1(n7971), .B2(n7970), .A(n8103), .ZN(n7972) );
  OAI21_X1 U9577 ( .B1(n7973), .B2(n7972), .A(n8044), .ZN(n7977) );
  AOI22_X1 U9578 ( .A1(n8097), .A2(n7974), .B1(n8101), .B2(n9793), .ZN(n7976)
         );
  MUX2_X1 U9579 ( .A(n8099), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n7975) );
  NAND3_X1 U9580 ( .A1(n7977), .A2(n7976), .A3(n7975), .ZN(P2_U3220) );
  INV_X1 U9581 ( .A(n7978), .ZN(n7979) );
  AOI21_X1 U9582 ( .B1(n8053), .B2(n7979), .A(n8103), .ZN(n7983) );
  NOR3_X1 U9583 ( .A1(n7980), .A2(n7984), .A3(n8040), .ZN(n7982) );
  OAI21_X1 U9584 ( .B1(n7983), .B2(n7982), .A(n7981), .ZN(n7989) );
  OAI22_X1 U9585 ( .A1(n8099), .A2(n8592), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10045), .ZN(n7987) );
  OAI22_X1 U9586 ( .A1(n7985), .A2(n8068), .B1(n8069), .B2(n7984), .ZN(n7986)
         );
  AOI211_X1 U9587 ( .C1(n8812), .C2(n8101), .A(n7987), .B(n7986), .ZN(n7988)
         );
  NAND2_X1 U9588 ( .A1(n7989), .A2(n7988), .ZN(P2_U3225) );
  INV_X1 U9589 ( .A(n8091), .ZN(n7991) );
  NOR3_X1 U9590 ( .A1(n7991), .A2(n7990), .A3(n8103), .ZN(n7995) );
  NAND3_X1 U9591 ( .A1(n7992), .A2(n8077), .A3(n8544), .ZN(n7993) );
  OAI21_X1 U9592 ( .B1(n8091), .B2(n8103), .A(n7993), .ZN(n7994) );
  INV_X1 U9593 ( .A(n7996), .ZN(n8001) );
  INV_X1 U9594 ( .A(n7997), .ZN(n8533) );
  AOI22_X1 U9595 ( .A1(n8489), .A2(n8729), .B1(n8730), .B2(n8314), .ZN(n8529)
         );
  OAI22_X1 U9596 ( .A1(n7998), .A2(n8529), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10039), .ZN(n7999) );
  AOI21_X1 U9597 ( .B1(n8533), .B2(n8079), .A(n7999), .ZN(n8000) );
  OAI211_X1 U9598 ( .C1(n8791), .C2(n8074), .A(n8001), .B(n8000), .ZN(P2_U3227) );
  AOI22_X1 U9599 ( .A1(n8005), .A2(n8004), .B1(n8003), .B2(n8002), .ZN(n8009)
         );
  XNOR2_X1 U9600 ( .A(n8007), .B(n8006), .ZN(n8008) );
  XNOR2_X1 U9601 ( .A(n8009), .B(n8008), .ZN(n8013) );
  AOI22_X1 U9602 ( .A1(n8059), .A2(n8728), .B1(n8058), .B2(n8683), .ZN(n8010)
         );
  NAND2_X1 U9603 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n8401) );
  OAI211_X1 U9604 ( .C1(n8685), .C2(n8099), .A(n8010), .B(n8401), .ZN(n8011)
         );
  AOI21_X1 U9605 ( .B1(n8693), .B2(n8101), .A(n8011), .ZN(n8012) );
  OAI21_X1 U9606 ( .B1(n8013), .B2(n8103), .A(n8012), .ZN(P2_U3228) );
  AOI22_X1 U9607 ( .A1(n8730), .A2(n8317), .B1(n8316), .B2(n8729), .ZN(n8660)
         );
  INV_X1 U9608 ( .A(n8660), .ZN(n8014) );
  AOI22_X1 U9609 ( .A1(n8097), .A2(n8014), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n8015) );
  OAI21_X1 U9610 ( .B1(n8672), .B2(n8099), .A(n8015), .ZN(n8025) );
  NAND2_X1 U9611 ( .A1(n8017), .A2(n8016), .ZN(n8019) );
  AND2_X1 U9612 ( .A1(n8019), .A2(n8018), .ZN(n8023) );
  INV_X1 U9613 ( .A(n8020), .ZN(n8021) );
  AOI211_X1 U9614 ( .C1(n8023), .C2(n8022), .A(n8103), .B(n8021), .ZN(n8024)
         );
  AOI211_X1 U9615 ( .C1(n8675), .C2(n8101), .A(n8025), .B(n8024), .ZN(n8026)
         );
  INV_X1 U9616 ( .A(n8026), .ZN(P2_U3230) );
  NOR2_X1 U9617 ( .A1(n8028), .A2(n8027), .ZN(n8030) );
  OAI22_X1 U9618 ( .A1(n8034), .A2(n8103), .B1(n8031), .B2(n8040), .ZN(n8032)
         );
  OAI21_X1 U9619 ( .B1(n8034), .B2(n8033), .A(n8032), .ZN(n8038) );
  AOI22_X1 U9620 ( .A1(n8079), .A2(n8549), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8037) );
  AOI22_X1 U9621 ( .A1(n8058), .A2(n8544), .B1(n8059), .B2(n8315), .ZN(n8036)
         );
  NAND2_X1 U9622 ( .A1(n8550), .A2(n8101), .ZN(n8035) );
  NAND4_X1 U9623 ( .A1(n8038), .A2(n8037), .A3(n8036), .A4(n8035), .ZN(
        P2_U3231) );
  NOR3_X1 U9624 ( .A1(n8040), .A2(n8039), .A3(n8045), .ZN(n8041) );
  OAI21_X1 U9625 ( .B1(n8041), .B2(n8059), .A(n8326), .ZN(n8052) );
  AOI22_X1 U9626 ( .A1(n8058), .A2(n8325), .B1(n8042), .B2(n8101), .ZN(n8051)
         );
  OAI21_X1 U9627 ( .B1(n8045), .B2(n8044), .A(n8043), .ZN(n8049) );
  INV_X1 U9628 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8046) );
  OAI22_X1 U9629 ( .A1(n8099), .A2(n8047), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8046), .ZN(n8048) );
  AOI21_X1 U9630 ( .B1(n8085), .B2(n8049), .A(n8048), .ZN(n8050) );
  NAND3_X1 U9631 ( .A1(n8052), .A2(n8051), .A3(n8050), .ZN(P2_U3232) );
  INV_X1 U9632 ( .A(n8053), .ZN(n8054) );
  AOI211_X1 U9633 ( .C1(n8056), .C2(n8055), .A(n8103), .B(n8054), .ZN(n8063)
         );
  INV_X1 U9634 ( .A(n8057), .ZN(n8612) );
  AOI22_X1 U9635 ( .A1(n8079), .A2(n8612), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8061) );
  AOI22_X1 U9636 ( .A1(n8059), .A2(n8608), .B1(n8058), .B2(n8607), .ZN(n8060)
         );
  OAI211_X1 U9637 ( .C1(n8819), .C2(n8074), .A(n8061), .B(n8060), .ZN(n8062)
         );
  OR2_X1 U9638 ( .A1(n8063), .A2(n8062), .ZN(P2_U3235) );
  NAND2_X1 U9639 ( .A1(n8077), .A2(n8599), .ZN(n8067) );
  NAND2_X1 U9640 ( .A1(n8085), .A2(n8064), .ZN(n8066) );
  MUX2_X1 U9641 ( .A(n8067), .B(n8066), .S(n8065), .Z(n8073) );
  NOR2_X1 U9642 ( .A1(n8099), .A2(n8573), .ZN(n8071) );
  OAI22_X1 U9643 ( .A1(n8580), .A2(n8069), .B1(n8068), .B2(n8579), .ZN(n8070)
         );
  AOI211_X1 U9644 ( .C1(P2_REG3_REG_22__SCAN_IN), .C2(P2_U3152), .A(n8071), 
        .B(n8070), .ZN(n8072) );
  OAI211_X1 U9645 ( .C1(n8576), .C2(n8074), .A(n8073), .B(n8072), .ZN(P2_U3237) );
  INV_X1 U9646 ( .A(n8084), .ZN(n8076) );
  NAND4_X1 U9647 ( .A1(n8077), .A2(n8076), .A3(n8325), .A4(n8075), .ZN(n8090)
         );
  AOI22_X1 U9648 ( .A1(n8101), .A2(n8080), .B1(n8079), .B2(n8078), .ZN(n8089)
         );
  AOI22_X1 U9649 ( .A1(n8097), .A2(n8081), .B1(P2_REG3_REG_6__SCAN_IN), .B2(
        P2_U3152), .ZN(n8088) );
  OAI21_X1 U9650 ( .B1(n8084), .B2(n8083), .A(n8082), .ZN(n8086) );
  NAND2_X1 U9651 ( .A1(n8086), .A2(n8085), .ZN(n8087) );
  NAND4_X1 U9652 ( .A1(n8090), .A2(n8089), .A3(n8088), .A4(n8087), .ZN(
        P2_U3241) );
  NAND2_X1 U9653 ( .A1(n8092), .A2(n8091), .ZN(n8094) );
  XNOR2_X1 U9654 ( .A(n8094), .B(n8093), .ZN(n8104) );
  OAI22_X1 U9655 ( .A1(n8096), .A2(n8650), .B1(n8095), .B2(n8648), .ZN(n8507)
         );
  AOI22_X1 U9656 ( .A1(n8097), .A2(n8507), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3152), .ZN(n8098) );
  OAI21_X1 U9657 ( .B1(n8513), .B2(n8099), .A(n8098), .ZN(n8100) );
  AOI21_X1 U9658 ( .B1(n8786), .B2(n8101), .A(n8100), .ZN(n8102) );
  OAI21_X1 U9659 ( .B1(n8104), .B2(n8103), .A(n8102), .ZN(P2_U3242) );
  NOR2_X1 U9660 ( .A1(n8110), .A2(n9997), .ZN(n8106) );
  AOI21_X2 U9661 ( .B1(n8107), .B2(n8108), .A(n8106), .ZN(n8764) );
  AND2_X1 U9662 ( .A1(n8764), .A2(n8313), .ZN(n8260) );
  NAND2_X1 U9663 ( .A1(n8109), .A2(n8108), .ZN(n8112) );
  OR2_X1 U9664 ( .A1(n8110), .A2(n6088), .ZN(n8111) );
  INV_X1 U9665 ( .A(n8462), .ZN(n8113) );
  OR2_X2 U9666 ( .A1(n8459), .A2(n8113), .ZN(n8263) );
  INV_X1 U9667 ( .A(n8764), .ZN(n8458) );
  NAND2_X1 U9668 ( .A1(n8458), .A2(n8114), .ZN(n8257) );
  AND2_X2 U9669 ( .A1(n8263), .A2(n8257), .ZN(n8259) );
  OAI21_X1 U9670 ( .B1(n8116), .B2(n8260), .A(n8259), .ZN(n8118) );
  NAND2_X1 U9671 ( .A1(n8113), .A2(n8301), .ZN(n8115) );
  AOI21_X1 U9672 ( .B1(n8116), .B2(n8764), .A(n8115), .ZN(n8117) );
  OAI21_X1 U9673 ( .B1(n8118), .B2(n8117), .A(n8264), .ZN(n8119) );
  XNOR2_X1 U9674 ( .A(n8119), .B(n8511), .ZN(n8306) );
  NAND2_X1 U9675 ( .A1(n4253), .A2(n8120), .ZN(n8305) );
  INV_X1 U9676 ( .A(n7871), .ZN(n9446) );
  AND2_X1 U9677 ( .A1(n8301), .A2(n8511), .ZN(n8122) );
  NAND2_X1 U9678 ( .A1(n5462), .A2(n8122), .ZN(n8262) );
  MUX2_X1 U9679 ( .A(n9446), .B(n8123), .S(n8262), .Z(n8184) );
  NAND2_X1 U9680 ( .A1(n8134), .A2(n8124), .ZN(n8131) );
  INV_X1 U9681 ( .A(n8125), .ZN(n8126) );
  AOI21_X1 U9682 ( .B1(n8127), .B2(n8326), .A(n8126), .ZN(n8128) );
  INV_X1 U9683 ( .A(n8141), .ZN(n8130) );
  INV_X1 U9684 ( .A(n8131), .ZN(n8133) );
  INV_X1 U9685 ( .A(n8135), .ZN(n8138) );
  NAND2_X1 U9686 ( .A1(n5462), .A2(n8511), .ZN(n8766) );
  AOI211_X1 U9687 ( .C1(n8136), .C2(n8766), .A(n5463), .B(n8279), .ZN(n8137)
         );
  OAI22_X1 U9688 ( .A1(n8138), .A2(n8137), .B1(n4249), .B2(n8262), .ZN(n8140)
         );
  NOR2_X1 U9689 ( .A1(n8140), .A2(n8139), .ZN(n8144) );
  MUX2_X1 U9690 ( .A(n8142), .B(n8141), .S(n8262), .Z(n8143) );
  OAI21_X1 U9691 ( .B1(n4286), .B2(n8144), .A(n4697), .ZN(n8150) );
  NAND2_X1 U9692 ( .A1(n8323), .A2(n4590), .ZN(n8148) );
  NAND2_X1 U9693 ( .A1(n8145), .A2(n8262), .ZN(n8147) );
  MUX2_X1 U9694 ( .A(n8148), .B(n8147), .S(n8146), .Z(n8149) );
  NAND3_X1 U9695 ( .A1(n8150), .A2(n8276), .A3(n8149), .ZN(n8155) );
  MUX2_X1 U9696 ( .A(n8152), .B(n8151), .S(n8262), .Z(n8153) );
  NAND3_X1 U9697 ( .A1(n8155), .A2(n8154), .A3(n8153), .ZN(n8168) );
  INV_X1 U9698 ( .A(n8282), .ZN(n8158) );
  INV_X1 U9699 ( .A(n8161), .ZN(n8157) );
  NAND2_X1 U9700 ( .A1(n8162), .A2(n4590), .ZN(n8156) );
  OAI22_X1 U9701 ( .A1(n8159), .A2(n8158), .B1(n8157), .B2(n8156), .ZN(n8167)
         );
  NAND2_X1 U9702 ( .A1(n8170), .A2(n8160), .ZN(n8165) );
  INV_X1 U9703 ( .A(n8160), .ZN(n8163) );
  OAI211_X1 U9704 ( .C1(n8163), .C2(n8162), .A(n8169), .B(n8161), .ZN(n8164)
         );
  MUX2_X1 U9705 ( .A(n8165), .B(n8164), .S(n8262), .Z(n8166) );
  AOI21_X1 U9706 ( .B1(n8168), .B2(n8167), .A(n8166), .ZN(n8177) );
  NAND2_X1 U9707 ( .A1(n8173), .A2(n8169), .ZN(n8172) );
  NAND2_X1 U9708 ( .A1(n8174), .A2(n8170), .ZN(n8171) );
  MUX2_X1 U9709 ( .A(n8172), .B(n8171), .S(n8262), .Z(n8176) );
  MUX2_X1 U9710 ( .A(n8174), .B(n8173), .S(n8262), .Z(n8175) );
  OAI21_X1 U9711 ( .B1(n8177), .B2(n8176), .A(n8175), .ZN(n8182) );
  INV_X1 U9712 ( .A(n8178), .ZN(n8179) );
  MUX2_X1 U9713 ( .A(n4661), .B(n8179), .S(n8262), .Z(n8180) );
  AOI211_X1 U9714 ( .C1(n8182), .C2(n8181), .A(n8180), .B(n4662), .ZN(n8183)
         );
  AOI211_X1 U9715 ( .C1(n8699), .C2(n8184), .A(n8706), .B(n8183), .ZN(n8188)
         );
  NOR2_X1 U9716 ( .A1(n9442), .A2(n8262), .ZN(n8186) );
  NOR2_X1 U9717 ( .A1(n7917), .A2(n4590), .ZN(n8185) );
  MUX2_X1 U9718 ( .A(n8186), .B(n8185), .S(n8728), .Z(n8187) );
  INV_X1 U9719 ( .A(n8189), .ZN(n8192) );
  INV_X1 U9720 ( .A(n8190), .ZN(n8191) );
  MUX2_X1 U9721 ( .A(n8192), .B(n8191), .S(n4590), .Z(n8193) );
  NAND2_X1 U9722 ( .A1(n8209), .A2(n8194), .ZN(n8197) );
  INV_X1 U9723 ( .A(n8195), .ZN(n8196) );
  MUX2_X1 U9724 ( .A(n8197), .B(n8196), .S(n8262), .Z(n8198) );
  INV_X1 U9725 ( .A(n8199), .ZN(n8208) );
  NOR3_X1 U9726 ( .A1(n8207), .A2(n8200), .A3(n8208), .ZN(n8202) );
  NOR2_X1 U9727 ( .A1(n8202), .A2(n8201), .ZN(n8204) );
  INV_X1 U9728 ( .A(n8214), .ZN(n8203) );
  OAI211_X1 U9729 ( .C1(n8204), .C2(n8203), .A(n8217), .B(n8212), .ZN(n8206)
         );
  NAND2_X1 U9730 ( .A1(n8595), .A2(n8607), .ZN(n8213) );
  NAND4_X1 U9731 ( .A1(n8206), .A2(n4590), .A3(n8205), .A4(n8213), .ZN(n8226)
         );
  AOI21_X1 U9732 ( .B1(n8210), .B2(n8209), .A(n8208), .ZN(n8216) );
  NAND2_X1 U9733 ( .A1(n8212), .A2(n8211), .ZN(n8215) );
  OAI211_X1 U9734 ( .C1(n8216), .C2(n8215), .A(n8214), .B(n8213), .ZN(n8218)
         );
  NAND3_X1 U9735 ( .A1(n8218), .A2(n8217), .A3(n4595), .ZN(n8222) );
  OAI21_X1 U9736 ( .B1(n8807), .B2(n4595), .A(n8577), .ZN(n8221) );
  INV_X1 U9737 ( .A(n8219), .ZN(n8220) );
  AOI22_X1 U9738 ( .A1(n8542), .A2(n8224), .B1(n8227), .B2(n4595), .ZN(n8225)
         );
  INV_X1 U9739 ( .A(n8227), .ZN(n8230) );
  INV_X1 U9740 ( .A(n8228), .ZN(n8229) );
  MUX2_X1 U9741 ( .A(n8230), .B(n8229), .S(n4595), .Z(n8231) );
  AOI21_X1 U9742 ( .B1(n8505), .B2(n8233), .A(n8232), .ZN(n8238) );
  INV_X1 U9743 ( .A(n8233), .ZN(n8234) );
  AOI21_X1 U9744 ( .B1(n8236), .B2(n8235), .A(n8234), .ZN(n8237) );
  MUX2_X1 U9745 ( .A(n8238), .B(n8237), .S(n8262), .Z(n8239) );
  NOR2_X1 U9746 ( .A1(n8240), .A2(n8239), .ZN(n8247) );
  INV_X1 U9747 ( .A(n8252), .ZN(n8243) );
  INV_X1 U9748 ( .A(n8241), .ZN(n8242) );
  NOR2_X1 U9749 ( .A1(n8243), .A2(n8242), .ZN(n8245) );
  MUX2_X1 U9750 ( .A(n8245), .B(n8244), .S(n8262), .Z(n8246) );
  OAI211_X1 U9751 ( .C1(n8247), .C2(n8501), .A(n8246), .B(n8248), .ZN(n8253)
         );
  NAND3_X1 U9752 ( .A1(n8253), .A2(n8249), .A3(n8248), .ZN(n8250) );
  AOI21_X1 U9753 ( .B1(n8253), .B2(n8252), .A(n8251), .ZN(n8254) );
  INV_X1 U9754 ( .A(n8255), .ZN(n8256) );
  INV_X1 U9755 ( .A(n8257), .ZN(n8258) );
  INV_X1 U9756 ( .A(n8259), .ZN(n8297) );
  INV_X1 U9757 ( .A(n8260), .ZN(n8261) );
  NAND2_X1 U9758 ( .A1(n8264), .A2(n8261), .ZN(n8298) );
  MUX2_X1 U9759 ( .A(n8297), .B(n8298), .S(n8262), .Z(n8266) );
  MUX2_X1 U9760 ( .A(n8264), .B(n8263), .S(n8262), .Z(n8265) );
  OAI21_X1 U9761 ( .B1(n8267), .B2(n8266), .A(n8265), .ZN(n8271) );
  OAI211_X1 U9762 ( .C1(n8269), .C2(n8270), .A(n8271), .B(n8268), .ZN(n8304)
         );
  NOR2_X1 U9763 ( .A1(n8271), .A2(n8270), .ZN(n8302) );
  INV_X1 U9764 ( .A(n8542), .ZN(n8293) );
  INV_X1 U9765 ( .A(n8639), .ZN(n8646) );
  NOR3_X1 U9766 ( .A1(n8273), .A2(n8272), .A3(n9752), .ZN(n8275) );
  NAND4_X1 U9767 ( .A1(n8275), .A2(n8765), .A3(n8274), .A4(n9774), .ZN(n8280)
         );
  INV_X1 U9768 ( .A(n8276), .ZN(n8277) );
  NOR4_X1 U9769 ( .A1(n8280), .A2(n8279), .A3(n8278), .A4(n8277), .ZN(n8283)
         );
  NAND4_X1 U9770 ( .A1(n8283), .A2(n8282), .A3(n8281), .A4(n4269), .ZN(n8287)
         );
  NOR4_X1 U9771 ( .A1(n8287), .A2(n8286), .A3(n8285), .A4(n8284), .ZN(n8289)
         );
  NAND4_X1 U9772 ( .A1(n4607), .A2(n8726), .A3(n8289), .A4(n8288), .ZN(n8290)
         );
  NOR4_X1 U9773 ( .A1(n8624), .A2(n8646), .A3(n8670), .A4(n8290), .ZN(n8291)
         );
  NAND4_X1 U9774 ( .A1(n4594), .A2(n8605), .A3(n4390), .A4(n8291), .ZN(n8292)
         );
  NOR4_X1 U9775 ( .A1(n8522), .A2(n8293), .A3(n8292), .A4(n8597), .ZN(n8294)
         );
  NAND4_X1 U9776 ( .A1(n8470), .A2(n4598), .A3(n8487), .A4(n8294), .ZN(n8295)
         );
  XNOR2_X1 U9777 ( .A(n8299), .B(n8511), .ZN(n8300) );
  OAI22_X1 U9778 ( .A1(n8302), .A2(n8765), .B1(n8301), .B2(n8300), .ZN(n8303)
         );
  AOI22_X1 U9779 ( .A1(n8306), .A2(n8305), .B1(n8304), .B2(n8303), .ZN(n8312)
         );
  NAND3_X1 U9780 ( .A1(n8755), .A2(n8307), .A3(n8730), .ZN(n8308) );
  OAI211_X1 U9781 ( .C1(n8309), .C2(n8311), .A(n8308), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8310) );
  OAI21_X1 U9782 ( .B1(n8312), .B2(n8311), .A(n8310), .ZN(P2_U3244) );
  MUX2_X1 U9783 ( .A(n8313), .B(P2_DATAO_REG_30__SCAN_IN), .S(n8328), .Z(
        P2_U3582) );
  MUX2_X1 U9784 ( .A(n8472), .B(P2_DATAO_REG_29__SCAN_IN), .S(n8328), .Z(
        P2_U3581) );
  MUX2_X1 U9785 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n8490), .S(P2_U3966), .Z(
        P2_U3580) );
  MUX2_X1 U9786 ( .A(n8473), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8328), .Z(
        P2_U3579) );
  MUX2_X1 U9787 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n8489), .S(P2_U3966), .Z(
        P2_U3578) );
  MUX2_X1 U9788 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8544), .S(P2_U3966), .Z(
        P2_U3577) );
  MUX2_X1 U9789 ( .A(n8314), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8328), .Z(
        P2_U3576) );
  MUX2_X1 U9790 ( .A(n8315), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8328), .Z(
        P2_U3575) );
  MUX2_X1 U9791 ( .A(n8599), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8328), .Z(
        P2_U3574) );
  MUX2_X1 U9792 ( .A(n8607), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8328), .Z(
        P2_U3573) );
  MUX2_X1 U9793 ( .A(n8600), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8328), .Z(
        P2_U3572) );
  MUX2_X1 U9794 ( .A(n8608), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8328), .Z(
        P2_U3571) );
  MUX2_X1 U9795 ( .A(n8316), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8328), .Z(
        P2_U3570) );
  MUX2_X1 U9796 ( .A(n8683), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8328), .Z(
        P2_U3569) );
  MUX2_X1 U9797 ( .A(n8317), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8328), .Z(
        P2_U3568) );
  MUX2_X1 U9798 ( .A(n8728), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8328), .Z(
        P2_U3567) );
  MUX2_X1 U9799 ( .A(n4663), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8328), .Z(
        P2_U3566) );
  MUX2_X1 U9800 ( .A(n8731), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8328), .Z(
        P2_U3565) );
  MUX2_X1 U9801 ( .A(n8318), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8328), .Z(
        P2_U3564) );
  MUX2_X1 U9802 ( .A(n8319), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8328), .Z(
        P2_U3563) );
  MUX2_X1 U9803 ( .A(n8320), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8328), .Z(
        P2_U3562) );
  MUX2_X1 U9804 ( .A(n8321), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8328), .Z(
        P2_U3561) );
  MUX2_X1 U9805 ( .A(n8322), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8328), .Z(
        P2_U3560) );
  MUX2_X1 U9806 ( .A(n8323), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8328), .Z(
        P2_U3559) );
  MUX2_X1 U9807 ( .A(n8324), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8328), .Z(
        P2_U3558) );
  MUX2_X1 U9808 ( .A(n8325), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8328), .Z(
        P2_U3557) );
  MUX2_X1 U9809 ( .A(n4400), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8328), .Z(
        P2_U3556) );
  MUX2_X1 U9810 ( .A(n8326), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8328), .Z(
        P2_U3555) );
  MUX2_X1 U9811 ( .A(n8327), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8328), .Z(
        P2_U3554) );
  MUX2_X1 U9812 ( .A(n6691), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8328), .Z(
        P2_U3553) );
  MUX2_X1 U9813 ( .A(n6702), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8328), .Z(
        P2_U3552) );
  AOI211_X1 U9814 ( .C1(n8331), .C2(n8330), .A(n8329), .B(n9738), .ZN(n8340)
         );
  OAI211_X1 U9815 ( .C1(n8334), .C2(n8333), .A(n9732), .B(n8332), .ZN(n8337)
         );
  AND2_X1 U9816 ( .A1(P2_U3152), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n8335) );
  AOI21_X1 U9817 ( .B1(n9376), .B2(P2_ADDR_REG_3__SCAN_IN), .A(n8335), .ZN(
        n8336) );
  OAI211_X1 U9818 ( .C1(n9739), .C2(n8338), .A(n8337), .B(n8336), .ZN(n8339)
         );
  OR2_X1 U9819 ( .A1(n8340), .A2(n8339), .ZN(P2_U3248) );
  AOI211_X1 U9820 ( .C1(n8343), .C2(n8342), .A(n8341), .B(n9738), .ZN(n8352)
         );
  OAI211_X1 U9821 ( .C1(n8346), .C2(n8345), .A(n9732), .B(n8344), .ZN(n8349)
         );
  NOR2_X1 U9822 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4840), .ZN(n8347) );
  AOI21_X1 U9823 ( .B1(n9376), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n8347), .ZN(
        n8348) );
  OAI211_X1 U9824 ( .C1(n9739), .C2(n8350), .A(n8349), .B(n8348), .ZN(n8351)
         );
  OR2_X1 U9825 ( .A1(n8352), .A2(n8351), .ZN(P2_U3250) );
  OAI211_X1 U9826 ( .C1(n8355), .C2(n8354), .A(n9733), .B(n8353), .ZN(n8364)
         );
  AND2_X1 U9827 ( .A1(P2_U3152), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n8356) );
  AOI21_X1 U9828 ( .B1(n9376), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n8356), .ZN(
        n8363) );
  INV_X1 U9829 ( .A(n9739), .ZN(n9382) );
  NAND2_X1 U9830 ( .A1(n9382), .A2(n8357), .ZN(n8362) );
  OAI211_X1 U9831 ( .C1(n8360), .C2(n8359), .A(n9732), .B(n8358), .ZN(n8361)
         );
  NAND4_X1 U9832 ( .A1(n8364), .A2(n8363), .A3(n8362), .A4(n8361), .ZN(
        P2_U3252) );
  OAI21_X1 U9833 ( .B1(n8367), .B2(n8366), .A(n8365), .ZN(n8368) );
  AOI22_X1 U9834 ( .A1(n9733), .A2(n8368), .B1(n8370), .B2(n9382), .ZN(n8378)
         );
  NOR2_X1 U9835 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n4992), .ZN(n8369) );
  AOI21_X1 U9836 ( .B1(n9376), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n8369), .ZN(
        n8377) );
  MUX2_X1 U9837 ( .A(n9882), .B(P2_REG1_REG_11__SCAN_IN), .S(n8370), .Z(n8371)
         );
  NAND3_X1 U9838 ( .A1(n8373), .A2(n8372), .A3(n8371), .ZN(n8374) );
  NAND3_X1 U9839 ( .A1(n8375), .A2(n9732), .A3(n8374), .ZN(n8376) );
  NAND3_X1 U9840 ( .A1(n8378), .A2(n8377), .A3(n8376), .ZN(P2_U3256) );
  AOI21_X1 U9841 ( .B1(n8381), .B2(n8380), .A(n8379), .ZN(n8392) );
  AOI211_X1 U9842 ( .C1(n8384), .C2(n8383), .A(n8382), .B(n9738), .ZN(n8390)
         );
  NOR2_X1 U9843 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8385), .ZN(n8386) );
  AOI21_X1 U9844 ( .B1(n9376), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n8386), .ZN(
        n8387) );
  OAI21_X1 U9845 ( .B1(n9739), .B2(n8388), .A(n8387), .ZN(n8389) );
  NOR2_X1 U9846 ( .A1(n8390), .A2(n8389), .ZN(n8391) );
  OAI21_X1 U9847 ( .B1(n8392), .B2(n9740), .A(n8391), .ZN(P2_U3257) );
  INV_X1 U9848 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8396) );
  INV_X1 U9849 ( .A(n8393), .ZN(n8394) );
  OAI22_X1 U9850 ( .A1(n8397), .A2(n8396), .B1(n8395), .B2(n8394), .ZN(n8400)
         );
  MUX2_X1 U9851 ( .A(n8398), .B(P2_REG1_REG_16__SCAN_IN), .S(n8418), .Z(n8399)
         );
  NOR2_X1 U9852 ( .A1(n8399), .A2(n8400), .ZN(n8419) );
  AOI21_X1 U9853 ( .B1(n8400), .B2(n8399), .A(n8419), .ZN(n8413) );
  INV_X1 U9854 ( .A(n8401), .ZN(n8402) );
  AOI21_X1 U9855 ( .B1(n9376), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n8402), .ZN(
        n8403) );
  INV_X1 U9856 ( .A(n8403), .ZN(n8411) );
  OAI22_X1 U9857 ( .A1(n8406), .A2(n8405), .B1(n8404), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U9858 ( .A1(n8418), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n8407) );
  OAI21_X1 U9859 ( .B1(n8418), .B2(P2_REG2_REG_16__SCAN_IN), .A(n8407), .ZN(
        n8408) );
  NOR2_X1 U9860 ( .A1(n8408), .A2(n8409), .ZN(n8414) );
  AOI211_X1 U9861 ( .C1(n8409), .C2(n8408), .A(n8414), .B(n9738), .ZN(n8410)
         );
  AOI211_X1 U9862 ( .C1(n9382), .C2(n8418), .A(n8411), .B(n8410), .ZN(n8412)
         );
  OAI21_X1 U9863 ( .B1(n8413), .B2(n9740), .A(n8412), .ZN(P2_U3261) );
  NAND2_X1 U9864 ( .A1(n8434), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8415) );
  OAI21_X1 U9865 ( .B1(n8434), .B2(P2_REG2_REG_17__SCAN_IN), .A(n8415), .ZN(
        n8416) );
  AOI211_X1 U9866 ( .C1(n8417), .C2(n8416), .A(n8433), .B(n9738), .ZN(n8428)
         );
  INV_X1 U9867 ( .A(n8418), .ZN(n8420) );
  AOI21_X1 U9868 ( .B1(n8420), .B2(n8398), .A(n8419), .ZN(n8423) );
  MUX2_X1 U9869 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8421), .S(n8434), .Z(n8422)
         );
  NAND2_X1 U9870 ( .A1(n8422), .A2(n8423), .ZN(n8429) );
  OAI211_X1 U9871 ( .C1(n8423), .C2(n8422), .A(n9732), .B(n8429), .ZN(n8426)
         );
  AND2_X1 U9872 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8424) );
  AOI21_X1 U9873 ( .B1(n9376), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8424), .ZN(
        n8425) );
  OAI211_X1 U9874 ( .C1(n9739), .C2(n8430), .A(n8426), .B(n8425), .ZN(n8427)
         );
  OR2_X1 U9875 ( .A1(n8428), .A2(n8427), .ZN(P2_U3262) );
  OAI21_X1 U9876 ( .B1(n8421), .B2(n8430), .A(n8429), .ZN(n8432) );
  AOI22_X1 U9877 ( .A1(n8439), .A2(n9932), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8448), .ZN(n8431) );
  NOR2_X1 U9878 ( .A1(n8432), .A2(n8431), .ZN(n8447) );
  AOI21_X1 U9879 ( .B1(n8432), .B2(n8431), .A(n8447), .ZN(n8442) );
  NAND2_X1 U9880 ( .A1(n8435), .A2(n5160), .ZN(n8445) );
  OAI21_X1 U9881 ( .B1(n8435), .B2(n5160), .A(n8445), .ZN(n8436) );
  NAND2_X1 U9882 ( .A1(n8436), .A2(n9733), .ZN(n8441) );
  INV_X1 U9883 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10070) );
  NOR2_X1 U9884 ( .A1(n9736), .A2(n10070), .ZN(n8437) );
  AOI211_X1 U9885 ( .C1(n9382), .C2(n8439), .A(n8438), .B(n8437), .ZN(n8440)
         );
  OAI211_X1 U9886 ( .C1(n8442), .C2(n9740), .A(n8441), .B(n8440), .ZN(P2_U3263) );
  NAND2_X1 U9887 ( .A1(n8443), .A2(n8448), .ZN(n8444) );
  NAND2_X1 U9888 ( .A1(n8445), .A2(n8444), .ZN(n8446) );
  XNOR2_X1 U9889 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8446), .ZN(n8453) );
  INV_X1 U9890 ( .A(n8453), .ZN(n8451) );
  AOI21_X1 U9891 ( .B1(n8448), .B2(n9932), .A(n8447), .ZN(n8449) );
  XNOR2_X1 U9892 ( .A(n8829), .B(n8449), .ZN(n8452) );
  OAI21_X1 U9893 ( .B1(n8452), .B2(n9740), .A(n9739), .ZN(n8450) );
  AOI21_X1 U9894 ( .B1(n8451), .B2(n9733), .A(n8450), .ZN(n8455) );
  AOI22_X1 U9895 ( .A1(n8453), .A2(n9733), .B1(n9732), .B2(n8452), .ZN(n8454)
         );
  MUX2_X1 U9896 ( .A(n8455), .B(n8454), .S(n4764), .Z(n8457) );
  NAND2_X1 U9897 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_U3152), .ZN(n8456) );
  OAI211_X1 U9898 ( .C1(n4754), .C2(n9736), .A(n8457), .B(n8456), .ZN(P2_U3264) );
  XNOR2_X1 U9899 ( .A(n8460), .B(n8459), .ZN(n8749) );
  NAND2_X1 U9900 ( .A1(n8749), .A2(n9755), .ZN(n8464) );
  NAND2_X1 U9901 ( .A1(n8462), .A2(n8461), .ZN(n8762) );
  NOR2_X1 U9902 ( .A1(n8655), .A2(n8762), .ZN(n8466) );
  AOI21_X1 U9903 ( .B1(n9762), .B2(P2_REG2_REG_31__SCAN_IN), .A(n8466), .ZN(
        n8463) );
  OAI211_X1 U9904 ( .C1(n8750), .C2(n9758), .A(n8464), .B(n8463), .ZN(P2_U3265) );
  XNOR2_X1 U9905 ( .A(n8465), .B(n8764), .ZN(n8761) );
  NAND2_X1 U9906 ( .A1(n8761), .A2(n9755), .ZN(n8468) );
  AOI21_X1 U9907 ( .B1(n9762), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8466), .ZN(
        n8467) );
  OAI211_X1 U9908 ( .C1(n8764), .C2(n9758), .A(n8468), .B(n8467), .ZN(P2_U3266) );
  OAI211_X1 U9909 ( .C1(n8471), .C2(n8470), .A(n8469), .B(n9748), .ZN(n8475)
         );
  AOI22_X1 U9910 ( .A1(n8473), .A2(n8730), .B1(n8729), .B2(n8472), .ZN(n8474)
         );
  AND2_X1 U9911 ( .A1(n8493), .A2(n8773), .ZN(n8476) );
  NOR2_X1 U9912 ( .A1(n8477), .A2(n8476), .ZN(n8774) );
  INV_X1 U9913 ( .A(n8478), .ZN(n8479) );
  AOI22_X1 U9914 ( .A1(n8655), .A2(P2_REG2_REG_28__SCAN_IN), .B1(n8479), .B2(
        n9750), .ZN(n8480) );
  OAI21_X1 U9915 ( .B1(n4527), .B2(n9758), .A(n8480), .ZN(n8481) );
  AOI21_X1 U9916 ( .B1(n8774), .B2(n9755), .A(n8481), .ZN(n8485) );
  OAI21_X1 U9917 ( .B1(n8483), .B2(n4667), .A(n8482), .ZN(n8772) );
  NAND2_X1 U9918 ( .A1(n8772), .A2(n9753), .ZN(n8484) );
  OAI211_X1 U9919 ( .C1(n8776), .C2(n8655), .A(n8485), .B(n8484), .ZN(P2_U3268) );
  OAI211_X1 U9920 ( .C1(n8488), .C2(n8487), .A(n8486), .B(n9748), .ZN(n8492)
         );
  AOI22_X1 U9921 ( .A1(n8490), .A2(n8729), .B1(n8730), .B2(n8489), .ZN(n8491)
         );
  INV_X1 U9922 ( .A(n8493), .ZN(n8494) );
  AOI21_X1 U9923 ( .B1(n8779), .B2(n8509), .A(n8494), .ZN(n8780) );
  INV_X1 U9924 ( .A(n8779), .ZN(n8498) );
  INV_X1 U9925 ( .A(n8495), .ZN(n8496) );
  AOI22_X1 U9926 ( .A1(n9762), .A2(P2_REG2_REG_27__SCAN_IN), .B1(n8496), .B2(
        n9750), .ZN(n8497) );
  OAI21_X1 U9927 ( .B1(n8498), .B2(n9758), .A(n8497), .ZN(n8499) );
  AOI21_X1 U9928 ( .B1(n8780), .B2(n9755), .A(n8499), .ZN(n8504) );
  OAI21_X1 U9929 ( .B1(n8502), .B2(n8501), .A(n8500), .ZN(n8778) );
  NAND2_X1 U9930 ( .A1(n8778), .A2(n9753), .ZN(n8503) );
  OAI211_X1 U9931 ( .C1(n8782), .C2(n8655), .A(n8504), .B(n8503), .ZN(P2_U3269) );
  NAND2_X1 U9932 ( .A1(n8526), .A2(n8505), .ZN(n8506) );
  XNOR2_X1 U9933 ( .A(n8506), .B(n8518), .ZN(n8508) );
  AOI21_X1 U9934 ( .B1(n8508), .B2(n9748), .A(n8507), .ZN(n8788) );
  INV_X1 U9935 ( .A(n8509), .ZN(n8510) );
  AOI211_X1 U9936 ( .C1(n8786), .C2(n8531), .A(n9861), .B(n8510), .ZN(n8785)
         );
  NOR2_X1 U9937 ( .A1(n8655), .A2(n8511), .ZN(n8532) );
  INV_X1 U9938 ( .A(n8786), .ZN(n8512) );
  NOR2_X1 U9939 ( .A1(n8512), .A2(n9758), .ZN(n8516) );
  OAI22_X1 U9940 ( .A1(n6962), .A2(n8514), .B1(n8513), .B2(n8739), .ZN(n8515)
         );
  AOI211_X1 U9941 ( .C1(n8785), .C2(n8532), .A(n8516), .B(n8515), .ZN(n8521)
         );
  OAI21_X1 U9942 ( .B1(n8519), .B2(n8518), .A(n8517), .ZN(n8784) );
  NAND2_X1 U9943 ( .A1(n8784), .A2(n9753), .ZN(n8520) );
  OAI211_X1 U9944 ( .C1(n8788), .C2(n8655), .A(n8521), .B(n8520), .ZN(P2_U3270) );
  OR2_X1 U9945 ( .A1(n8523), .A2(n8522), .ZN(n8524) );
  NAND2_X1 U9946 ( .A1(n8525), .A2(n8524), .ZN(n8794) );
  INV_X1 U9947 ( .A(n8794), .ZN(n8539) );
  OAI211_X1 U9948 ( .C1(n8528), .C2(n8527), .A(n8526), .B(n9748), .ZN(n8530)
         );
  NAND2_X1 U9949 ( .A1(n8530), .A2(n8529), .ZN(n8792) );
  OAI211_X1 U9950 ( .C1(n8548), .C2(n8791), .A(n8832), .B(n8531), .ZN(n8790)
         );
  INV_X1 U9951 ( .A(n8532), .ZN(n8677) );
  AOI22_X1 U9952 ( .A1(n9762), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n8533), .B2(
        n9750), .ZN(n8536) );
  NAND2_X1 U9953 ( .A1(n8534), .A2(n8743), .ZN(n8535) );
  OAI211_X1 U9954 ( .C1(n8790), .C2(n8677), .A(n8536), .B(n8535), .ZN(n8537)
         );
  AOI21_X1 U9955 ( .B1(n8792), .B2(n6962), .A(n8537), .ZN(n8538) );
  OAI21_X1 U9956 ( .B1(n8722), .B2(n8539), .A(n8538), .ZN(P2_U3271) );
  XNOR2_X1 U9957 ( .A(n8540), .B(n8542), .ZN(n8800) );
  INV_X1 U9958 ( .A(n8800), .ZN(n8555) );
  OAI211_X1 U9959 ( .C1(n8543), .C2(n8542), .A(n8541), .B(n9748), .ZN(n8546)
         );
  NAND2_X1 U9960 ( .A1(n8544), .A2(n8729), .ZN(n8545) );
  OAI211_X1 U9961 ( .C1(n8579), .C2(n8648), .A(n8546), .B(n8545), .ZN(n8798)
         );
  NOR2_X1 U9962 ( .A1(n8560), .A2(n8796), .ZN(n8547) );
  OR2_X1 U9963 ( .A1(n8548), .A2(n8547), .ZN(n8797) );
  AOI22_X1 U9964 ( .A1(n8655), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n8549), .B2(
        n9750), .ZN(n8552) );
  NAND2_X1 U9965 ( .A1(n8550), .A2(n8743), .ZN(n8551) );
  OAI211_X1 U9966 ( .C1(n8797), .C2(n8745), .A(n8552), .B(n8551), .ZN(n8553)
         );
  AOI21_X1 U9967 ( .B1(n8798), .B2(n6962), .A(n8553), .ZN(n8554) );
  OAI21_X1 U9968 ( .B1(n8722), .B2(n8555), .A(n8554), .ZN(P2_U3272) );
  OAI21_X1 U9969 ( .B1(n4280), .B2(n8556), .A(n8565), .ZN(n8557) );
  NAND2_X1 U9970 ( .A1(n4316), .A2(n8557), .ZN(n8559) );
  AOI21_X1 U9971 ( .B1(n8559), .B2(n9748), .A(n8558), .ZN(n8805) );
  AOI21_X1 U9972 ( .B1(n8802), .B2(n8572), .A(n8560), .ZN(n8803) );
  AOI22_X1 U9973 ( .A1(n9762), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n8561), .B2(
        n9750), .ZN(n8562) );
  OAI21_X1 U9974 ( .B1(n8563), .B2(n9758), .A(n8562), .ZN(n8568) );
  OAI21_X1 U9975 ( .B1(n8566), .B2(n8565), .A(n8564), .ZN(n8806) );
  NOR2_X1 U9976 ( .A1(n8806), .A2(n8722), .ZN(n8567) );
  AOI211_X1 U9977 ( .C1(n8803), .C2(n9755), .A(n8568), .B(n8567), .ZN(n8569)
         );
  OAI21_X1 U9978 ( .B1(n8805), .B2(n8655), .A(n8569), .ZN(P2_U3273) );
  XNOR2_X1 U9979 ( .A(n8570), .B(n8577), .ZN(n8811) );
  NAND2_X1 U9980 ( .A1(n8589), .A2(n8807), .ZN(n8571) );
  AND2_X1 U9981 ( .A1(n8572), .A2(n8571), .ZN(n8808) );
  INV_X1 U9982 ( .A(n8573), .ZN(n8574) );
  AOI22_X1 U9983 ( .A1(n9762), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8574), .B2(
        n9750), .ZN(n8575) );
  OAI21_X1 U9984 ( .B1(n8576), .B2(n9758), .A(n8575), .ZN(n8584) );
  AOI211_X1 U9985 ( .C1(n8578), .C2(n8577), .A(n8661), .B(n4280), .ZN(n8582)
         );
  OAI22_X1 U9986 ( .A1(n8580), .A2(n8648), .B1(n8579), .B2(n8650), .ZN(n8581)
         );
  NOR2_X1 U9987 ( .A1(n8582), .A2(n8581), .ZN(n8810) );
  NOR2_X1 U9988 ( .A1(n8810), .A2(n8655), .ZN(n8583) );
  AOI211_X1 U9989 ( .C1(n8808), .C2(n9755), .A(n8584), .B(n8583), .ZN(n8585)
         );
  OAI21_X1 U9990 ( .B1(n8722), .B2(n8811), .A(n8585), .ZN(P2_U3274) );
  NAND2_X1 U9991 ( .A1(n8617), .A2(n8616), .ZN(n8618) );
  NAND2_X1 U9992 ( .A1(n8618), .A2(n8586), .ZN(n8587) );
  XNOR2_X1 U9993 ( .A(n8587), .B(n8597), .ZN(n8816) );
  INV_X1 U9994 ( .A(n8588), .ZN(n8591) );
  INV_X1 U9995 ( .A(n8589), .ZN(n8590) );
  AOI21_X1 U9996 ( .B1(n8812), .B2(n8591), .A(n8590), .ZN(n8813) );
  INV_X1 U9997 ( .A(n8592), .ZN(n8593) );
  AOI22_X1 U9998 ( .A1(n9762), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8593), .B2(
        n9750), .ZN(n8594) );
  OAI21_X1 U9999 ( .B1(n8595), .B2(n9758), .A(n8594), .ZN(n8602) );
  XNOR2_X1 U10000 ( .A(n8596), .B(n8597), .ZN(n8598) );
  AOI222_X1 U10001 ( .A1(n8600), .A2(n8730), .B1(n8599), .B2(n8729), .C1(n9748), .C2(n8598), .ZN(n8815) );
  NOR2_X1 U10002 ( .A1(n8815), .A2(n8655), .ZN(n8601) );
  AOI211_X1 U10003 ( .C1(n8813), .C2(n9755), .A(n8602), .B(n8601), .ZN(n8603)
         );
  OAI21_X1 U10004 ( .B1(n8722), .B2(n8816), .A(n8603), .ZN(P2_U3275) );
  OAI211_X1 U10005 ( .C1(n8606), .C2(n8605), .A(n8604), .B(n9748), .ZN(n8610)
         );
  AOI22_X1 U10006 ( .A1(n8730), .A2(n8608), .B1(n8607), .B2(n8729), .ZN(n8609)
         );
  NAND2_X1 U10007 ( .A1(n8610), .A2(n8609), .ZN(n8822) );
  NOR2_X1 U10008 ( .A1(n8631), .A2(n8819), .ZN(n8611) );
  OR2_X1 U10009 ( .A1(n8588), .A2(n8611), .ZN(n8820) );
  AOI22_X1 U10010 ( .A1(n8655), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8612), .B2(
        n9750), .ZN(n8615) );
  NAND2_X1 U10011 ( .A1(n8613), .A2(n8743), .ZN(n8614) );
  OAI211_X1 U10012 ( .C1(n8820), .C2(n8745), .A(n8615), .B(n8614), .ZN(n8620)
         );
  NOR2_X1 U10013 ( .A1(n8617), .A2(n8616), .ZN(n8818) );
  INV_X1 U10014 ( .A(n8618), .ZN(n8817) );
  NOR3_X1 U10015 ( .A1(n8818), .A2(n8817), .A3(n8722), .ZN(n8619) );
  AOI211_X1 U10016 ( .C1(n6962), .C2(n8822), .A(n8620), .B(n8619), .ZN(n8621)
         );
  INV_X1 U10017 ( .A(n8621), .ZN(P2_U3276) );
  XNOR2_X1 U10018 ( .A(n8622), .B(n8624), .ZN(n8826) );
  NAND2_X1 U10019 ( .A1(n8653), .A2(n8623), .ZN(n8625) );
  XNOR2_X1 U10020 ( .A(n8625), .B(n8624), .ZN(n8626) );
  NAND2_X1 U10021 ( .A1(n8626), .A2(n9748), .ZN(n8628) );
  NAND2_X1 U10022 ( .A1(n8628), .A2(n8627), .ZN(n8633) );
  NAND2_X1 U10023 ( .A1(n8641), .A2(n8824), .ZN(n8629) );
  NAND2_X1 U10024 ( .A1(n8629), .A2(n8832), .ZN(n8630) );
  NOR2_X1 U10025 ( .A1(n8631), .A2(n8630), .ZN(n8632) );
  OAI211_X1 U10026 ( .C1(n4764), .C2(n8633), .A(n8828), .B(n6962), .ZN(n8638)
         );
  INV_X1 U10027 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8635) );
  OAI22_X1 U10028 ( .A1(n6962), .A2(n8635), .B1(n8634), .B2(n8739), .ZN(n8636)
         );
  AOI21_X1 U10029 ( .B1(n8824), .B2(n8743), .A(n8636), .ZN(n8637) );
  OAI211_X1 U10030 ( .C1(n8722), .C2(n8826), .A(n8638), .B(n8637), .ZN(
        P2_U3277) );
  XNOR2_X1 U10031 ( .A(n8640), .B(n8639), .ZN(n8836) );
  AOI21_X1 U10032 ( .B1(n8831), .B2(n4276), .A(n4523), .ZN(n8833) );
  AOI22_X1 U10033 ( .A1(n8655), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8642), .B2(
        n9750), .ZN(n8643) );
  OAI21_X1 U10034 ( .B1(n8644), .B2(n9758), .A(n8643), .ZN(n8657) );
  INV_X1 U10035 ( .A(n8645), .ZN(n8647) );
  AOI21_X1 U10036 ( .B1(n8647), .B2(n8646), .A(n8661), .ZN(n8654) );
  OAI22_X1 U10037 ( .A1(n8651), .A2(n8650), .B1(n8649), .B2(n8648), .ZN(n8652)
         );
  AOI21_X1 U10038 ( .B1(n8654), .B2(n8653), .A(n8652), .ZN(n8835) );
  NOR2_X1 U10039 ( .A1(n8835), .A2(n8655), .ZN(n8656) );
  AOI211_X1 U10040 ( .C1(n8833), .C2(n9755), .A(n8657), .B(n8656), .ZN(n8658)
         );
  OAI21_X1 U10041 ( .B1(n8722), .B2(n8836), .A(n8658), .ZN(P2_U3278) );
  XNOR2_X1 U10042 ( .A(n8659), .B(n8670), .ZN(n8662) );
  OAI21_X1 U10043 ( .B1(n8662), .B2(n8661), .A(n8660), .ZN(n9430) );
  INV_X1 U10044 ( .A(n9430), .ZN(n8680) );
  NAND2_X1 U10045 ( .A1(n8735), .A2(n8664), .ZN(n8666) );
  NAND2_X1 U10046 ( .A1(n8666), .A2(n8665), .ZN(n8671) );
  AND2_X1 U10047 ( .A1(n8668), .A2(n8667), .ZN(n8669) );
  OAI21_X1 U10048 ( .B1(n8671), .B2(n8670), .A(n8669), .ZN(n9432) );
  OAI211_X1 U10049 ( .C1(n8687), .C2(n9429), .A(n8832), .B(n4276), .ZN(n9428)
         );
  OAI22_X1 U10050 ( .A1(n6962), .A2(n8673), .B1(n8672), .B2(n8739), .ZN(n8674)
         );
  AOI21_X1 U10051 ( .B1(n8675), .B2(n8743), .A(n8674), .ZN(n8676) );
  OAI21_X1 U10052 ( .B1(n9428), .B2(n8677), .A(n8676), .ZN(n8678) );
  AOI21_X1 U10053 ( .B1(n9432), .B2(n9753), .A(n8678), .ZN(n8679) );
  OAI21_X1 U10054 ( .B1(n8680), .B2(n8655), .A(n8679), .ZN(P2_U3279) );
  XNOR2_X1 U10055 ( .A(n8681), .B(n8682), .ZN(n8684) );
  AOI222_X1 U10056 ( .A1(n9748), .A2(n8684), .B1(n8683), .B2(n8729), .C1(n8728), .C2(n8730), .ZN(n9433) );
  OAI21_X1 U10057 ( .B1(n8685), .B2(n8739), .A(n9433), .ZN(n8697) );
  NOR2_X1 U10058 ( .A1(n8712), .A2(n9436), .ZN(n8686) );
  OR2_X1 U10059 ( .A1(n8687), .A2(n8686), .ZN(n9437) );
  NAND2_X1 U10060 ( .A1(n8735), .A2(n8688), .ZN(n8691) );
  NAND2_X1 U10061 ( .A1(n8691), .A2(n8689), .ZN(n9435) );
  NAND2_X1 U10062 ( .A1(n8691), .A2(n8690), .ZN(n8692) );
  NAND2_X1 U10063 ( .A1(n8692), .A2(n4607), .ZN(n9434) );
  NAND3_X1 U10064 ( .A1(n9435), .A2(n9753), .A3(n9434), .ZN(n8695) );
  AOI22_X1 U10065 ( .A1(n8743), .A2(n8693), .B1(n9762), .B2(
        P2_REG2_REG_16__SCAN_IN), .ZN(n8694) );
  OAI211_X1 U10066 ( .C1(n8745), .C2(n9437), .A(n8695), .B(n8694), .ZN(n8696)
         );
  AOI21_X1 U10067 ( .B1(n8697), .B2(n6962), .A(n8696), .ZN(n8698) );
  INV_X1 U10068 ( .A(n8698), .ZN(P2_U3280) );
  NAND2_X1 U10069 ( .A1(n8735), .A2(n4662), .ZN(n8734) );
  NAND2_X1 U10070 ( .A1(n8734), .A2(n8699), .ZN(n8700) );
  XNOR2_X1 U10071 ( .A(n8700), .B(n8706), .ZN(n9445) );
  INV_X1 U10072 ( .A(n9445), .ZN(n8721) );
  NAND2_X1 U10073 ( .A1(n7881), .A2(n8701), .ZN(n8703) );
  NAND2_X1 U10074 ( .A1(n8703), .A2(n8702), .ZN(n8708) );
  NAND2_X1 U10075 ( .A1(n8724), .A2(n8704), .ZN(n8725) );
  NAND3_X1 U10076 ( .A1(n8725), .A2(n8706), .A3(n8705), .ZN(n8707) );
  NAND3_X1 U10077 ( .A1(n8708), .A2(n9748), .A3(n8707), .ZN(n8710) );
  NAND2_X1 U10078 ( .A1(n8710), .A2(n8709), .ZN(n9443) );
  NAND2_X1 U10079 ( .A1(n8738), .A2(n7917), .ZN(n8711) );
  NAND2_X1 U10080 ( .A1(n8711), .A2(n8832), .ZN(n8713) );
  OR2_X1 U10081 ( .A1(n8713), .A2(n8712), .ZN(n9441) );
  INV_X1 U10082 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8715) );
  OAI22_X1 U10083 ( .A1(n6962), .A2(n8715), .B1(n8714), .B2(n8739), .ZN(n8716)
         );
  AOI21_X1 U10084 ( .B1(n8743), .B2(n7917), .A(n8716), .ZN(n8717) );
  OAI21_X1 U10085 ( .B1(n9441), .B2(n8718), .A(n8717), .ZN(n8719) );
  AOI21_X1 U10086 ( .B1(n9443), .B2(n6962), .A(n8719), .ZN(n8720) );
  OAI21_X1 U10087 ( .B1(n8722), .B2(n8721), .A(n8720), .ZN(P2_U3281) );
  AND2_X1 U10088 ( .A1(n8724), .A2(n8723), .ZN(n8727) );
  OAI211_X1 U10089 ( .C1(n8727), .C2(n8726), .A(n8725), .B(n9748), .ZN(n8733)
         );
  AOI22_X1 U10090 ( .A1(n8731), .A2(n8730), .B1(n8729), .B2(n8728), .ZN(n8732)
         );
  NAND2_X1 U10091 ( .A1(n8733), .A2(n8732), .ZN(n9448) );
  INV_X1 U10092 ( .A(n9448), .ZN(n8748) );
  OAI21_X1 U10093 ( .B1(n8735), .B2(n4662), .A(n8734), .ZN(n9450) );
  NAND2_X1 U10094 ( .A1(n8736), .A2(n7871), .ZN(n8737) );
  NAND2_X1 U10095 ( .A1(n8738), .A2(n8737), .ZN(n9447) );
  OAI22_X1 U10096 ( .A1(n6962), .A2(n8741), .B1(n8740), .B2(n8739), .ZN(n8742)
         );
  AOI21_X1 U10097 ( .B1(n8743), .B2(n7871), .A(n8742), .ZN(n8744) );
  OAI21_X1 U10098 ( .B1(n9447), .B2(n8745), .A(n8744), .ZN(n8746) );
  AOI21_X1 U10099 ( .B1(n9450), .B2(n9753), .A(n8746), .ZN(n8747) );
  OAI21_X1 U10100 ( .B1(n8748), .B2(n8655), .A(n8747), .ZN(P2_U3282) );
  AND2_X1 U10101 ( .A1(n8755), .A2(n8754), .ZN(n8756) );
  NAND2_X1 U10102 ( .A1(n8757), .A2(n8756), .ZN(n8758) );
  MUX2_X1 U10103 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n8839), .S(n4256), .Z(
        P2_U3551) );
  NAND2_X1 U10104 ( .A1(n8761), .A2(n8832), .ZN(n8763) );
  OAI211_X1 U10105 ( .C1(n8764), .C2(n9859), .A(n8763), .B(n8762), .ZN(n8840)
         );
  MUX2_X1 U10106 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8840), .S(n4256), .Z(
        P2_U3550) );
  OR2_X1 U10107 ( .A1(n8766), .A2(n8765), .ZN(n9847) );
  INV_X1 U10108 ( .A(n8772), .ZN(n8777) );
  AOI22_X1 U10109 ( .A1(n8774), .A2(n8832), .B1(n9843), .B2(n8773), .ZN(n8775)
         );
  OAI211_X1 U10110 ( .C1(n9807), .C2(n8777), .A(n8776), .B(n8775), .ZN(n8842)
         );
  MUX2_X1 U10111 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8842), .S(n4256), .Z(
        P2_U3548) );
  INV_X1 U10112 ( .A(n8778), .ZN(n8783) );
  AOI22_X1 U10113 ( .A1(n8780), .A2(n8832), .B1(n9843), .B2(n8779), .ZN(n8781)
         );
  OAI211_X1 U10114 ( .C1(n9807), .C2(n8783), .A(n8782), .B(n8781), .ZN(n8843)
         );
  MUX2_X1 U10115 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8843), .S(n4256), .Z(
        P2_U3547) );
  INV_X1 U10116 ( .A(n8784), .ZN(n8789) );
  AOI21_X1 U10117 ( .B1(n9843), .B2(n8786), .A(n8785), .ZN(n8787) );
  OAI211_X1 U10118 ( .C1(n9807), .C2(n8789), .A(n8788), .B(n8787), .ZN(n8844)
         );
  MUX2_X1 U10119 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8844), .S(n4256), .Z(
        P2_U3546) );
  OAI21_X1 U10120 ( .B1(n8791), .B2(n9859), .A(n8790), .ZN(n8793) );
  AOI211_X1 U10121 ( .C1(n9866), .C2(n8794), .A(n8793), .B(n8792), .ZN(n8795)
         );
  INV_X1 U10122 ( .A(n8795), .ZN(n8845) );
  MUX2_X1 U10123 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8845), .S(n4256), .Z(
        P2_U3545) );
  OAI22_X1 U10124 ( .A1(n8797), .A2(n9861), .B1(n8796), .B2(n9859), .ZN(n8799)
         );
  AOI211_X1 U10125 ( .C1(n8800), .C2(n9866), .A(n8799), .B(n8798), .ZN(n8801)
         );
  INV_X1 U10126 ( .A(n8801), .ZN(n8846) );
  MUX2_X1 U10127 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8846), .S(n4256), .Z(
        P2_U3544) );
  AOI22_X1 U10128 ( .A1(n8803), .A2(n8832), .B1(n9843), .B2(n8802), .ZN(n8804)
         );
  OAI211_X1 U10129 ( .C1(n9807), .C2(n8806), .A(n8805), .B(n8804), .ZN(n8847)
         );
  MUX2_X1 U10130 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8847), .S(n4256), .Z(
        P2_U3543) );
  AOI22_X1 U10131 ( .A1(n8808), .A2(n8832), .B1(n9843), .B2(n8807), .ZN(n8809)
         );
  OAI211_X1 U10132 ( .C1(n9807), .C2(n8811), .A(n8810), .B(n8809), .ZN(n8848)
         );
  MUX2_X1 U10133 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8848), .S(n4256), .Z(
        P2_U3542) );
  AOI22_X1 U10134 ( .A1(n8813), .A2(n8832), .B1(n9843), .B2(n8812), .ZN(n8814)
         );
  OAI211_X1 U10135 ( .C1(n9807), .C2(n8816), .A(n8815), .B(n8814), .ZN(n8849)
         );
  MUX2_X1 U10136 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8849), .S(n4256), .Z(
        P2_U3541) );
  NOR3_X1 U10137 ( .A1(n8818), .A2(n8817), .A3(n9807), .ZN(n8823) );
  OAI22_X1 U10138 ( .A1(n8820), .A2(n9861), .B1(n8819), .B2(n9859), .ZN(n8821)
         );
  MUX2_X1 U10139 ( .A(n8850), .B(P2_REG1_REG_20__SCAN_IN), .S(n9884), .Z(
        P2_U3540) );
  INV_X1 U10140 ( .A(n8824), .ZN(n8825) );
  OAI22_X1 U10141 ( .A1(n8826), .A2(n9807), .B1(n8825), .B2(n9859), .ZN(n8827)
         );
  NOR2_X1 U10142 ( .A1(n8828), .A2(n8827), .ZN(n8851) );
  MUX2_X1 U10143 ( .A(n8829), .B(n8851), .S(n4256), .Z(n8830) );
  INV_X1 U10144 ( .A(n8830), .ZN(P2_U3539) );
  AOI22_X1 U10145 ( .A1(n8833), .A2(n8832), .B1(n9843), .B2(n8831), .ZN(n8834)
         );
  OAI211_X1 U10146 ( .C1(n9807), .C2(n8836), .A(n8835), .B(n8834), .ZN(n8853)
         );
  MUX2_X1 U10147 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8853), .S(n4256), .Z(
        P2_U3538) );
  MUX2_X1 U10148 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n8839), .S(n4255), .Z(
        P2_U3519) );
  MUX2_X1 U10149 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8840), .S(n4255), .Z(
        P2_U3518) );
  MUX2_X1 U10150 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8841), .S(n4255), .Z(
        P2_U3517) );
  MUX2_X1 U10151 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8842), .S(n4255), .Z(
        P2_U3516) );
  MUX2_X1 U10152 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8843), .S(n4255), .Z(
        P2_U3515) );
  MUX2_X1 U10153 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8844), .S(n4255), .Z(
        P2_U3514) );
  MUX2_X1 U10154 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8845), .S(n4255), .Z(
        P2_U3513) );
  MUX2_X1 U10155 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8846), .S(n4255), .Z(
        P2_U3512) );
  MUX2_X1 U10156 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8847), .S(n4255), .Z(
        P2_U3511) );
  MUX2_X1 U10157 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8848), .S(n4255), .Z(
        P2_U3510) );
  MUX2_X1 U10158 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8849), .S(n4255), .Z(
        P2_U3509) );
  MUX2_X1 U10159 ( .A(n8850), .B(P2_REG0_REG_20__SCAN_IN), .S(n9867), .Z(
        P2_U3508) );
  MUX2_X1 U10160 ( .A(n9920), .B(n8851), .S(n4255), .Z(n8852) );
  INV_X1 U10161 ( .A(n8852), .ZN(P2_U3507) );
  MUX2_X1 U10162 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8853), .S(n4255), .Z(
        P2_U3505) );
  INV_X1 U10163 ( .A(n8854), .ZN(n8855) );
  MUX2_X1 U10164 ( .A(n8855), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  INV_X1 U10165 ( .A(n9295), .ZN(n9095) );
  OAI21_X1 U10166 ( .B1(n8858), .B2(n8857), .A(n8856), .ZN(n8859) );
  NAND2_X1 U10167 ( .A1(n8859), .A2(n8969), .ZN(n8865) );
  INV_X1 U10168 ( .A(n8860), .ZN(n9092) );
  AOI22_X1 U10169 ( .A1(n8985), .A2(n9088), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8861) );
  OAI21_X1 U10170 ( .B1(n8862), .B2(n8956), .A(n8861), .ZN(n8863) );
  AOI21_X1 U10171 ( .B1(n9092), .B2(n8975), .A(n8863), .ZN(n8864) );
  OAI211_X1 U10172 ( .C1(n9095), .C2(n8961), .A(n8865), .B(n8864), .ZN(
        P1_U3212) );
  INV_X1 U10173 ( .A(n8869), .ZN(n8866) );
  NOR2_X1 U10174 ( .A1(n8867), .A2(n8866), .ZN(n8872) );
  AOI21_X1 U10175 ( .B1(n8870), .B2(n8869), .A(n8868), .ZN(n8871) );
  OAI21_X1 U10176 ( .B1(n8872), .B2(n8871), .A(n8969), .ZN(n8877) );
  AOI22_X1 U10177 ( .A1(n9162), .A2(n8986), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n8873) );
  OAI21_X1 U10178 ( .B1(n8874), .B2(n8898), .A(n8873), .ZN(n8875) );
  AOI21_X1 U10179 ( .B1(n9154), .B2(n8975), .A(n8875), .ZN(n8876) );
  OAI211_X1 U10180 ( .C1(n9156), .C2(n8961), .A(n8877), .B(n8876), .ZN(
        P1_U3214) );
  INV_X1 U10181 ( .A(n9334), .ZN(n9226) );
  NAND2_X1 U10182 ( .A1(n8880), .A2(n8969), .ZN(n8884) );
  NAND2_X1 U10183 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9064) );
  NAND2_X1 U10184 ( .A1(n8985), .A2(n9272), .ZN(n8881) );
  OAI211_X1 U10185 ( .C1(n8956), .C2(n8888), .A(n9064), .B(n8881), .ZN(n8882)
         );
  AOI21_X1 U10186 ( .B1(n9224), .B2(n8975), .A(n8882), .ZN(n8883) );
  OAI211_X1 U10187 ( .C1(n9226), .C2(n8961), .A(n8884), .B(n8883), .ZN(
        P1_U3217) );
  XOR2_X1 U10188 ( .A(n8886), .B(n8885), .Z(n8893) );
  AOI22_X1 U10189 ( .A1(n8986), .A2(n9190), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n8887) );
  OAI21_X1 U10190 ( .B1(n8888), .B2(n8898), .A(n8887), .ZN(n8891) );
  NAND2_X1 U10191 ( .A1(n9195), .A2(n9345), .ZN(n9326) );
  NOR2_X1 U10192 ( .A1(n9326), .A2(n8889), .ZN(n8890) );
  AOI211_X1 U10193 ( .C1(n9194), .C2(n8975), .A(n8891), .B(n8890), .ZN(n8892)
         );
  OAI21_X1 U10194 ( .B1(n8893), .B2(n8993), .A(n8892), .ZN(P1_U3221) );
  XOR2_X1 U10195 ( .A(n8895), .B(n8894), .Z(n8902) );
  AOI22_X1 U10196 ( .A1(n8986), .A2(n9088), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n8897) );
  NAND2_X1 U10197 ( .A1(n8975), .A2(n9120), .ZN(n8896) );
  OAI211_X1 U10198 ( .C1(n8899), .C2(n8898), .A(n8897), .B(n8896), .ZN(n8900)
         );
  AOI21_X1 U10199 ( .B1(n9303), .B2(n8991), .A(n8900), .ZN(n8901) );
  OAI21_X1 U10200 ( .B1(n8902), .B2(n8993), .A(n8901), .ZN(P1_U3223) );
  OAI21_X1 U10201 ( .B1(n8905), .B2(n8904), .A(n8903), .ZN(n8906) );
  NAND2_X1 U10202 ( .A1(n8906), .A2(n8969), .ZN(n8912) );
  NOR2_X1 U10203 ( .A1(n8989), .A2(n9148), .ZN(n8910) );
  OAI22_X1 U10204 ( .A1(n8908), .A2(n8956), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8907), .ZN(n8909) );
  AOI211_X1 U10205 ( .C1(n8985), .C2(n9176), .A(n8910), .B(n8909), .ZN(n8911)
         );
  OAI211_X1 U10206 ( .C1(n8913), .C2(n8961), .A(n8912), .B(n8911), .ZN(
        P1_U3227) );
  XNOR2_X1 U10207 ( .A(n8915), .B(n8914), .ZN(n8916) );
  XNOR2_X1 U10208 ( .A(n8917), .B(n8916), .ZN(n8918) );
  NAND2_X1 U10209 ( .A1(n8918), .A2(n8969), .ZN(n8926) );
  AND2_X1 U10210 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9024) );
  AOI21_X1 U10211 ( .B1(n8985), .B2(n9006), .A(n9024), .ZN(n8925) );
  INV_X1 U10212 ( .A(n8919), .ZN(n8921) );
  AOI22_X1 U10213 ( .A1(n8975), .A2(n8921), .B1(n8991), .B2(n8920), .ZN(n8924)
         );
  INV_X1 U10214 ( .A(n8922), .ZN(n9004) );
  NAND2_X1 U10215 ( .A1(n8986), .A2(n9004), .ZN(n8923) );
  NAND4_X1 U10216 ( .A1(n8926), .A2(n8925), .A3(n8924), .A4(n8923), .ZN(
        P1_U3228) );
  INV_X1 U10217 ( .A(n8927), .ZN(n8932) );
  AOI21_X1 U10218 ( .B1(n8929), .B2(n8931), .A(n8928), .ZN(n8930) );
  AOI21_X1 U10219 ( .B1(n8932), .B2(n8931), .A(n8930), .ZN(n8937) );
  AOI22_X1 U10220 ( .A1(n8986), .A2(n9175), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n8934) );
  NAND2_X1 U10221 ( .A1(n8985), .A2(n9243), .ZN(n8933) );
  OAI211_X1 U10222 ( .C1(n8989), .C2(n9215), .A(n8934), .B(n8933), .ZN(n8935)
         );
  AOI21_X1 U10223 ( .B1(n9331), .B2(n8991), .A(n8935), .ZN(n8936) );
  OAI21_X1 U10224 ( .B1(n8937), .B2(n8993), .A(n8936), .ZN(P1_U3231) );
  NAND2_X1 U10225 ( .A1(n8939), .A2(n8938), .ZN(n8940) );
  XOR2_X1 U10226 ( .A(n8941), .B(n8940), .Z(n8948) );
  OAI22_X1 U10227 ( .A1(n8956), .A2(n8943), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n8942), .ZN(n8944) );
  AOI21_X1 U10228 ( .B1(n8985), .B2(n9175), .A(n8944), .ZN(n8945) );
  OAI21_X1 U10229 ( .B1(n8989), .B2(n9170), .A(n8945), .ZN(n8946) );
  AOI21_X1 U10230 ( .B1(n9318), .B2(n8991), .A(n8946), .ZN(n8947) );
  OAI21_X1 U10231 ( .B1(n8948), .B2(n8993), .A(n8947), .ZN(P1_U3233) );
  INV_X1 U10232 ( .A(n8952), .ZN(n8949) );
  NOR2_X1 U10233 ( .A1(n8950), .A2(n8949), .ZN(n8955) );
  AOI21_X1 U10234 ( .B1(n8953), .B2(n8952), .A(n8951), .ZN(n8954) );
  OAI21_X1 U10235 ( .B1(n8955), .B2(n8954), .A(n8969), .ZN(n8960) );
  NOR2_X1 U10236 ( .A1(n8989), .A2(n9249), .ZN(n8958) );
  NAND2_X1 U10237 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9627) );
  OAI21_X1 U10238 ( .B1(n8956), .B2(n9211), .A(n9627), .ZN(n8957) );
  AOI211_X1 U10239 ( .C1(n8985), .C2(n9242), .A(n8958), .B(n8957), .ZN(n8959)
         );
  OAI211_X1 U10240 ( .C1(n4447), .C2(n8961), .A(n8960), .B(n8959), .ZN(
        P1_U3236) );
  INV_X1 U10241 ( .A(n8962), .ZN(n8963) );
  NOR2_X1 U10242 ( .A1(n8964), .A2(n8963), .ZN(n8968) );
  NAND2_X1 U10243 ( .A1(n8966), .A2(n8965), .ZN(n8967) );
  XNOR2_X1 U10244 ( .A(n8968), .B(n8967), .ZN(n8970) );
  NAND2_X1 U10245 ( .A1(n8970), .A2(n8969), .ZN(n8979) );
  AOI21_X1 U10246 ( .B1(n8985), .B2(n9004), .A(n8971), .ZN(n8978) );
  INV_X1 U10247 ( .A(n8972), .ZN(n8974) );
  AOI22_X1 U10248 ( .A1(n8975), .A2(n8974), .B1(n8991), .B2(n8973), .ZN(n8977)
         );
  NAND2_X1 U10249 ( .A1(n8986), .A2(n9002), .ZN(n8976) );
  NAND4_X1 U10250 ( .A1(n8979), .A2(n8978), .A3(n8977), .A4(n8976), .ZN(
        P1_U3237) );
  INV_X1 U10251 ( .A(n8980), .ZN(n8981) );
  NOR2_X1 U10252 ( .A1(n8982), .A2(n8981), .ZN(n8983) );
  XNOR2_X1 U10253 ( .A(n8984), .B(n8983), .ZN(n8994) );
  AOI22_X1 U10254 ( .A1(n9141), .A2(n8985), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n8988) );
  NAND2_X1 U10255 ( .A1(n8986), .A2(n9108), .ZN(n8987) );
  OAI211_X1 U10256 ( .C1(n8989), .C2(n9101), .A(n8988), .B(n8987), .ZN(n8990)
         );
  AOI21_X1 U10257 ( .B1(n9299), .B2(n8991), .A(n8990), .ZN(n8992) );
  OAI21_X1 U10258 ( .B1(n8994), .B2(n8993), .A(n8992), .ZN(P1_U3238) );
  MUX2_X1 U10259 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n8995), .S(n4257), .Z(
        P1_U3585) );
  MUX2_X1 U10260 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n8996), .S(n4257), .Z(
        P1_U3584) );
  MUX2_X1 U10261 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9087), .S(n4257), .Z(
        P1_U3583) );
  MUX2_X1 U10262 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9108), .S(n4257), .Z(
        P1_U3582) );
  MUX2_X1 U10263 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9088), .S(n4257), .Z(
        P1_U3581) );
  MUX2_X1 U10264 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9141), .S(n4257), .Z(
        P1_U3580) );
  MUX2_X1 U10265 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9162), .S(n4257), .Z(
        P1_U3579) );
  MUX2_X1 U10266 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9176), .S(n4257), .Z(
        P1_U3578) );
  MUX2_X1 U10267 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9175), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10268 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9233), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10269 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9243), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10270 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9272), .S(n4257), .Z(
        P1_U3573) );
  MUX2_X1 U10271 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9242), .S(n4257), .Z(
        P1_U3572) );
  MUX2_X1 U10272 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9478), .S(n4257), .Z(
        P1_U3571) );
  MUX2_X1 U10273 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n8997), .S(n4257), .Z(
        P1_U3570) );
  MUX2_X1 U10274 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9477), .S(n4257), .Z(
        P1_U3569) );
  MUX2_X1 U10275 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n8998), .S(n4257), .Z(
        P1_U3568) );
  MUX2_X1 U10276 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n8999), .S(n4257), .Z(
        P1_U3567) );
  MUX2_X1 U10277 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9000), .S(n4257), .Z(
        P1_U3566) );
  MUX2_X1 U10278 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9655), .S(n4257), .Z(
        P1_U3565) );
  MUX2_X1 U10279 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9001), .S(n4257), .Z(
        P1_U3564) );
  MUX2_X1 U10280 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9653), .S(n4257), .Z(
        P1_U3563) );
  MUX2_X1 U10281 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9002), .S(n4257), .Z(
        P1_U3562) );
  MUX2_X1 U10282 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9003), .S(n4257), .Z(
        P1_U3561) );
  MUX2_X1 U10283 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9004), .S(n4257), .Z(
        P1_U3560) );
  MUX2_X1 U10284 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9005), .S(n4257), .Z(
        P1_U3559) );
  MUX2_X1 U10285 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9006), .S(n4257), .Z(
        P1_U3558) );
  MUX2_X1 U10286 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9007), .S(n4257), .Z(
        P1_U3557) );
  MUX2_X1 U10287 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9008), .S(n4257), .Z(
        P1_U3556) );
  OAI22_X1 U10288 ( .A1(n9523), .A2(n9010), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9009), .ZN(n9011) );
  AOI21_X1 U10289 ( .B1(n9012), .B2(P1_ADDR_REG_1__SCAN_IN), .A(n9011), .ZN(
        n9021) );
  NAND3_X1 U10290 ( .A1(n9622), .A2(n9015), .A3(n9014), .ZN(n9020) );
  OAI211_X1 U10291 ( .C1(n9018), .C2(n9017), .A(n9526), .B(n9016), .ZN(n9019)
         );
  NAND3_X1 U10292 ( .A1(n9021), .A2(n9020), .A3(n9019), .ZN(P1_U3242) );
  INV_X1 U10293 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9022) );
  NOR2_X1 U10294 ( .A1(n9643), .A2(n9022), .ZN(n9023) );
  AOI211_X1 U10295 ( .C1(n9634), .C2(n9025), .A(n9024), .B(n9023), .ZN(n9035)
         );
  OAI21_X1 U10296 ( .B1(n9028), .B2(n9027), .A(n9026), .ZN(n9033) );
  OAI21_X1 U10297 ( .B1(n9031), .B2(n9030), .A(n9029), .ZN(n9032) );
  AOI22_X1 U10298 ( .A1(n9526), .A2(n9033), .B1(n9622), .B2(n9032), .ZN(n9034)
         );
  NAND3_X1 U10299 ( .A1(n9036), .A2(n9035), .A3(n9034), .ZN(P1_U3245) );
  NOR2_X1 U10300 ( .A1(n9038), .A2(n9037), .ZN(n9039) );
  NOR2_X1 U10301 ( .A1(n9039), .A2(n9047), .ZN(n9040) );
  INV_X1 U10302 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9592) );
  XNOR2_X1 U10303 ( .A(n9047), .B(n9039), .ZN(n9593) );
  NOR2_X1 U10304 ( .A1(n9592), .A2(n9593), .ZN(n9591) );
  NAND2_X1 U10305 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9607), .ZN(n9041) );
  OAI21_X1 U10306 ( .B1(n9607), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9041), .ZN(
        n9603) );
  NAND2_X1 U10307 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9620), .ZN(n9042) );
  OAI21_X1 U10308 ( .B1(n9620), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9042), .ZN(
        n9616) );
  NOR2_X1 U10309 ( .A1(n9635), .A2(n9043), .ZN(n9044) );
  AOI21_X1 U10310 ( .B1(n9635), .B2(n9043), .A(n9044), .ZN(n9630) );
  XNOR2_X1 U10311 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9045), .ZN(n9061) );
  INV_X1 U10312 ( .A(n9061), .ZN(n9059) );
  INV_X1 U10313 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9055) );
  XNOR2_X1 U10314 ( .A(n9635), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n9638) );
  INV_X1 U10315 ( .A(n9620), .ZN(n9053) );
  INV_X1 U10316 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9052) );
  XNOR2_X1 U10317 ( .A(n9053), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n9624) );
  INV_X1 U10318 ( .A(n9607), .ZN(n9051) );
  XOR2_X1 U10319 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9607), .Z(n9609) );
  NAND2_X1 U10320 ( .A1(n9596), .A2(n9048), .ZN(n9049) );
  XNOR2_X1 U10321 ( .A(n9048), .B(n9047), .ZN(n9598) );
  NAND2_X1 U10322 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9598), .ZN(n9597) );
  NAND2_X1 U10323 ( .A1(n9049), .A2(n9597), .ZN(n9610) );
  NAND2_X1 U10324 ( .A1(n9609), .A2(n9610), .ZN(n9608) );
  OAI21_X1 U10325 ( .B1(n9051), .B2(n9050), .A(n9608), .ZN(n9623) );
  NAND2_X1 U10326 ( .A1(n9624), .A2(n9623), .ZN(n9621) );
  OAI21_X1 U10327 ( .B1(n9053), .B2(n9052), .A(n9621), .ZN(n9637) );
  NOR2_X1 U10328 ( .A1(n9638), .A2(n9637), .ZN(n9636) );
  AOI21_X1 U10329 ( .B1(n9055), .B2(n9054), .A(n9636), .ZN(n9057) );
  XNOR2_X1 U10330 ( .A(n9057), .B(n9056), .ZN(n9060) );
  OAI21_X1 U10331 ( .B1(n9060), .B2(n9640), .A(n9523), .ZN(n9058) );
  AOI21_X1 U10332 ( .B1(n9059), .B2(n9526), .A(n9058), .ZN(n9063) );
  AOI22_X1 U10333 ( .A1(n9061), .A2(n9526), .B1(n9622), .B2(n9060), .ZN(n9062)
         );
  OAI211_X1 U10334 ( .C1(n9066), .C2(n9643), .A(n9065), .B(n9064), .ZN(
        P1_U3260) );
  INV_X1 U10335 ( .A(n9067), .ZN(n9068) );
  NAND2_X1 U10336 ( .A1(n9069), .A2(n9068), .ZN(n9284) );
  NAND3_X1 U10337 ( .A1(n9284), .A2(n9277), .A3(n9283), .ZN(n9072) );
  AOI21_X1 U10338 ( .B1(n9676), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9070), .ZN(
        n9071) );
  OAI211_X1 U10339 ( .C1(n9287), .C2(n9268), .A(n9072), .B(n9071), .ZN(
        P1_U3262) );
  INV_X1 U10340 ( .A(n9073), .ZN(n9083) );
  OAI22_X1 U10341 ( .A1(n9666), .A2(n9075), .B1(n9074), .B2(n9663), .ZN(n9076)
         );
  AOI21_X1 U10342 ( .B1(n9077), .B2(n9669), .A(n9076), .ZN(n9078) );
  OAI21_X1 U10343 ( .B1(n9079), .B2(n9671), .A(n9078), .ZN(n9080) );
  AOI21_X1 U10344 ( .B1(n9081), .B2(n9666), .A(n9080), .ZN(n9082) );
  OAI21_X1 U10345 ( .B1(n9083), .B2(n9279), .A(n9082), .ZN(P1_U3263) );
  XOR2_X1 U10346 ( .A(n9085), .B(n9084), .Z(n9297) );
  OAI21_X1 U10347 ( .B1(n9086), .B2(n9085), .A(n9651), .ZN(n9090) );
  AOI22_X1 U10348 ( .A1(n9654), .A2(n9088), .B1(n9656), .B2(n9087), .ZN(n9089)
         );
  OAI21_X1 U10349 ( .B1(n9090), .B2(n7842), .A(n9089), .ZN(n9293) );
  AOI211_X1 U10350 ( .C1(n9295), .C2(n9099), .A(n9714), .B(n9091), .ZN(n9294)
         );
  NAND2_X1 U10351 ( .A1(n9294), .A2(n9248), .ZN(n9094) );
  AOI22_X1 U10352 ( .A1(n9274), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9092), .B2(
        n9484), .ZN(n9093) );
  OAI211_X1 U10353 ( .C1(n9095), .C2(n9268), .A(n9094), .B(n9093), .ZN(n9096)
         );
  AOI21_X1 U10354 ( .B1(n9293), .B2(n9666), .A(n9096), .ZN(n9097) );
  OAI21_X1 U10355 ( .B1(n9297), .B2(n9279), .A(n9097), .ZN(P1_U3264) );
  XNOR2_X1 U10356 ( .A(n9098), .B(n9107), .ZN(n9302) );
  INV_X1 U10357 ( .A(n9099), .ZN(n9100) );
  AOI211_X1 U10358 ( .C1(n9299), .C2(n4464), .A(n9714), .B(n9100), .ZN(n9298)
         );
  INV_X1 U10359 ( .A(n9101), .ZN(n9102) );
  AOI22_X1 U10360 ( .A1(n9274), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9102), .B2(
        n9484), .ZN(n9103) );
  OAI21_X1 U10361 ( .B1(n9104), .B2(n9268), .A(n9103), .ZN(n9114) );
  NAND2_X1 U10362 ( .A1(n9105), .A2(n9128), .ZN(n9106) );
  XOR2_X1 U10363 ( .A(n9107), .B(n9106), .Z(n9112) );
  NAND2_X1 U10364 ( .A1(n9141), .A2(n9654), .ZN(n9109) );
  AOI211_X1 U10365 ( .C1(n9298), .C2(n9248), .A(n9114), .B(n9113), .ZN(n9115)
         );
  OAI21_X1 U10366 ( .B1(n9279), .B2(n9302), .A(n9115), .ZN(P1_U3265) );
  OAI21_X1 U10367 ( .B1(n9117), .B2(n9124), .A(n9116), .ZN(n9118) );
  INV_X1 U10368 ( .A(n9118), .ZN(n9307) );
  AOI21_X1 U10369 ( .B1(n9303), .B2(n9143), .A(n9119), .ZN(n9304) );
  AOI22_X1 U10370 ( .A1(n9120), .A2(n9484), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n9274), .ZN(n9121) );
  OAI21_X1 U10371 ( .B1(n9122), .B2(n9268), .A(n9121), .ZN(n9133) );
  NOR2_X1 U10372 ( .A1(n9123), .A2(n9210), .ZN(n9131) );
  INV_X1 U10373 ( .A(n9105), .ZN(n9129) );
  INV_X1 U10374 ( .A(n9124), .ZN(n9125) );
  OAI21_X1 U10375 ( .B1(n9126), .B2(n9125), .A(n9651), .ZN(n9127) );
  AOI21_X1 U10376 ( .B1(n9129), .B2(n9128), .A(n9127), .ZN(n9130) );
  NOR2_X1 U10377 ( .A1(n9306), .A2(n9274), .ZN(n9132) );
  AOI211_X1 U10378 ( .C1(n9304), .C2(n9277), .A(n9133), .B(n9132), .ZN(n9134)
         );
  OAI21_X1 U10379 ( .B1(n9307), .B2(n9279), .A(n9134), .ZN(P1_U3266) );
  XNOR2_X1 U10380 ( .A(n9135), .B(n9137), .ZN(n9312) );
  AOI22_X1 U10381 ( .A1(n9309), .A2(n9669), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9676), .ZN(n9151) );
  INV_X1 U10382 ( .A(n9136), .ZN(n9157) );
  OAI21_X1 U10383 ( .B1(n9157), .B2(n9138), .A(n9137), .ZN(n9140) );
  NAND2_X1 U10384 ( .A1(n9140), .A2(n9139), .ZN(n9142) );
  AOI222_X1 U10385 ( .A1(n9651), .A2(n9142), .B1(n9141), .B2(n9656), .C1(n9176), .C2(n9654), .ZN(n9311) );
  INV_X1 U10386 ( .A(n9153), .ZN(n9145) );
  INV_X1 U10387 ( .A(n9143), .ZN(n9144) );
  AOI211_X1 U10388 ( .C1(n9309), .C2(n9145), .A(n9714), .B(n9144), .ZN(n9308)
         );
  NAND2_X1 U10389 ( .A1(n9308), .A2(n9146), .ZN(n9147) );
  OAI211_X1 U10390 ( .C1(n9663), .C2(n9148), .A(n9311), .B(n9147), .ZN(n9149)
         );
  NAND2_X1 U10391 ( .A1(n9149), .A2(n9666), .ZN(n9150) );
  OAI211_X1 U10392 ( .C1(n9312), .C2(n9279), .A(n9151), .B(n9150), .ZN(
        P1_U3267) );
  XNOR2_X1 U10393 ( .A(n9152), .B(n9159), .ZN(n9317) );
  AOI21_X1 U10394 ( .B1(n9313), .B2(n9168), .A(n9153), .ZN(n9314) );
  AOI22_X1 U10395 ( .A1(n9676), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9154), .B2(
        n9484), .ZN(n9155) );
  OAI21_X1 U10396 ( .B1(n9156), .B2(n9268), .A(n9155), .ZN(n9164) );
  AND2_X1 U10397 ( .A1(n9190), .A2(n9654), .ZN(n9161) );
  AOI211_X1 U10398 ( .C1(n9159), .C2(n9158), .A(n9207), .B(n9157), .ZN(n9160)
         );
  AOI211_X1 U10399 ( .C1(n9656), .C2(n9162), .A(n9161), .B(n9160), .ZN(n9316)
         );
  NOR2_X1 U10400 ( .A1(n9316), .A2(n9274), .ZN(n9163) );
  AOI211_X1 U10401 ( .C1(n9314), .C2(n9277), .A(n9164), .B(n9163), .ZN(n9165)
         );
  OAI21_X1 U10402 ( .B1(n9279), .B2(n9317), .A(n9165), .ZN(P1_U3268) );
  XNOR2_X1 U10403 ( .A(n9166), .B(n4702), .ZN(n9322) );
  INV_X1 U10404 ( .A(n9167), .ZN(n9182) );
  INV_X1 U10405 ( .A(n9168), .ZN(n9169) );
  AOI21_X1 U10406 ( .B1(n9318), .B2(n9182), .A(n9169), .ZN(n9319) );
  INV_X1 U10407 ( .A(n9170), .ZN(n9171) );
  AOI22_X1 U10408 ( .A1(n9676), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9171), .B2(
        n9484), .ZN(n9172) );
  OAI21_X1 U10409 ( .B1(n9173), .B2(n9268), .A(n9172), .ZN(n9179) );
  XNOR2_X1 U10410 ( .A(n9174), .B(n4702), .ZN(n9177) );
  AOI222_X1 U10411 ( .A1(n9651), .A2(n9177), .B1(n9176), .B2(n9656), .C1(n9175), .C2(n9654), .ZN(n9321) );
  NOR2_X1 U10412 ( .A1(n9321), .A2(n9274), .ZN(n9178) );
  AOI211_X1 U10413 ( .C1(n9319), .C2(n9277), .A(n9179), .B(n9178), .ZN(n9180)
         );
  OAI21_X1 U10414 ( .B1(n9279), .B2(n9322), .A(n9180), .ZN(P1_U3269) );
  INV_X1 U10415 ( .A(n9195), .ZN(n9183) );
  INV_X1 U10416 ( .A(n9181), .ZN(n9213) );
  OAI211_X1 U10417 ( .C1(n9183), .C2(n9213), .A(n9182), .B(n9469), .ZN(n9325)
         );
  NOR2_X1 U10418 ( .A1(n9325), .A2(n9473), .ZN(n9193) );
  NAND2_X1 U10419 ( .A1(n9230), .A2(n9229), .ZN(n9203) );
  NAND2_X1 U10420 ( .A1(n9203), .A2(n9184), .ZN(n9186) );
  NAND2_X1 U10421 ( .A1(n9186), .A2(n9185), .ZN(n9188) );
  OAI21_X1 U10422 ( .B1(n9189), .B2(n9188), .A(n9187), .ZN(n9191) );
  AOI222_X1 U10423 ( .A1(n9651), .A2(n9191), .B1(n9233), .B2(n9654), .C1(n9190), .C2(n9656), .ZN(n9327) );
  INV_X1 U10424 ( .A(n9327), .ZN(n9192) );
  AOI211_X1 U10425 ( .C1(n9484), .C2(n9194), .A(n9193), .B(n9192), .ZN(n9201)
         );
  AOI22_X1 U10426 ( .A1(n9195), .A2(n9669), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9274), .ZN(n9200) );
  NOR2_X1 U10427 ( .A1(n9197), .A2(n9196), .ZN(n9323) );
  INV_X1 U10428 ( .A(n9198), .ZN(n9324) );
  OR3_X1 U10429 ( .A1(n9323), .A2(n9324), .A3(n9279), .ZN(n9199) );
  OAI211_X1 U10430 ( .C1(n9201), .C2(n9274), .A(n9200), .B(n9199), .ZN(
        P1_U3270) );
  XNOR2_X1 U10431 ( .A(n9202), .B(n9206), .ZN(n9333) );
  NAND2_X1 U10432 ( .A1(n9203), .A2(n9227), .ZN(n9232) );
  NAND2_X1 U10433 ( .A1(n9232), .A2(n9204), .ZN(n9205) );
  XOR2_X1 U10434 ( .A(n9206), .B(n9205), .Z(n9208) );
  OAI222_X1 U10435 ( .A1(n9212), .A2(n9211), .B1(n9210), .B2(n9209), .C1(n9208), .C2(n9207), .ZN(n9329) );
  INV_X1 U10436 ( .A(n9223), .ZN(n9214) );
  AOI211_X1 U10437 ( .C1(n9331), .C2(n9214), .A(n9714), .B(n9213), .ZN(n9330)
         );
  NAND2_X1 U10438 ( .A1(n9330), .A2(n9248), .ZN(n9218) );
  INV_X1 U10439 ( .A(n9215), .ZN(n9216) );
  AOI22_X1 U10440 ( .A1(n9274), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9216), .B2(
        n9484), .ZN(n9217) );
  OAI211_X1 U10441 ( .C1(n9219), .C2(n9268), .A(n9218), .B(n9217), .ZN(n9220)
         );
  AOI21_X1 U10442 ( .B1(n9329), .B2(n9666), .A(n9220), .ZN(n9221) );
  OAI21_X1 U10443 ( .B1(n9279), .B2(n9333), .A(n9221), .ZN(P1_U3271) );
  XOR2_X1 U10444 ( .A(n9222), .B(n9227), .Z(n9338) );
  AOI21_X1 U10445 ( .B1(n9334), .B2(n9246), .A(n9223), .ZN(n9335) );
  AOI22_X1 U10446 ( .A1(n9676), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9224), .B2(
        n9484), .ZN(n9225) );
  OAI21_X1 U10447 ( .B1(n9226), .B2(n9268), .A(n9225), .ZN(n9236) );
  INV_X1 U10448 ( .A(n9227), .ZN(n9228) );
  NAND3_X1 U10449 ( .A1(n9230), .A2(n9229), .A3(n9228), .ZN(n9231) );
  NAND2_X1 U10450 ( .A1(n9232), .A2(n9231), .ZN(n9234) );
  AOI222_X1 U10451 ( .A1(n9651), .A2(n9234), .B1(n9233), .B2(n9656), .C1(n9272), .C2(n9654), .ZN(n9337) );
  NOR2_X1 U10452 ( .A1(n9337), .A2(n9274), .ZN(n9235) );
  AOI211_X1 U10453 ( .C1(n9335), .C2(n9277), .A(n9236), .B(n9235), .ZN(n9237)
         );
  OAI21_X1 U10454 ( .B1(n9279), .B2(n9338), .A(n9237), .ZN(P1_U3272) );
  NAND2_X1 U10455 ( .A1(n9239), .A2(n9238), .ZN(n9240) );
  XNOR2_X1 U10456 ( .A(n9240), .B(n5765), .ZN(n9241) );
  NAND2_X1 U10457 ( .A1(n9241), .A2(n9651), .ZN(n9245) );
  AOI22_X1 U10458 ( .A1(n9243), .A2(n9656), .B1(n9654), .B2(n9242), .ZN(n9244)
         );
  NAND2_X1 U10459 ( .A1(n9245), .A2(n9244), .ZN(n9341) );
  AOI21_X1 U10460 ( .B1(n9251), .B2(n9263), .A(n9714), .ZN(n9247) );
  NAND2_X1 U10461 ( .A1(n9247), .A2(n9246), .ZN(n9339) );
  INV_X1 U10462 ( .A(n9248), .ZN(n9254) );
  INV_X1 U10463 ( .A(n9249), .ZN(n9250) );
  AOI22_X1 U10464 ( .A1(n9676), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n9250), .B2(
        n9484), .ZN(n9253) );
  NAND2_X1 U10465 ( .A1(n9251), .A2(n9669), .ZN(n9252) );
  OAI211_X1 U10466 ( .C1(n9339), .C2(n9254), .A(n9253), .B(n9252), .ZN(n9260)
         );
  NAND2_X1 U10467 ( .A1(n9256), .A2(n9255), .ZN(n9257) );
  NAND2_X1 U10468 ( .A1(n9258), .A2(n9257), .ZN(n9343) );
  NOR2_X1 U10469 ( .A1(n9343), .A2(n9279), .ZN(n9259) );
  AOI211_X1 U10470 ( .C1(n9666), .C2(n9341), .A(n9260), .B(n9259), .ZN(n9261)
         );
  INV_X1 U10471 ( .A(n9261), .ZN(P1_U3273) );
  XOR2_X1 U10472 ( .A(n9262), .B(n9270), .Z(n9350) );
  INV_X1 U10473 ( .A(n9263), .ZN(n9264) );
  AOI21_X1 U10474 ( .B1(n9344), .B2(n4317), .A(n9264), .ZN(n9346) );
  INV_X1 U10475 ( .A(n9265), .ZN(n9266) );
  AOI22_X1 U10476 ( .A1(n9676), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9266), .B2(
        n9484), .ZN(n9267) );
  OAI21_X1 U10477 ( .B1(n9269), .B2(n9268), .A(n9267), .ZN(n9276) );
  XNOR2_X1 U10478 ( .A(n9271), .B(n9270), .ZN(n9273) );
  AOI222_X1 U10479 ( .A1(n9651), .A2(n9273), .B1(n9272), .B2(n9656), .C1(n9478), .C2(n9654), .ZN(n9348) );
  NOR2_X1 U10480 ( .A1(n9348), .A2(n9274), .ZN(n9275) );
  AOI211_X1 U10481 ( .C1(n9346), .C2(n9277), .A(n9276), .B(n9275), .ZN(n9278)
         );
  OAI21_X1 U10482 ( .B1(n9279), .B2(n9350), .A(n9278), .ZN(P1_U3274) );
  NAND2_X1 U10483 ( .A1(n9280), .A2(n9345), .ZN(n9281) );
  OAI211_X1 U10484 ( .C1(n9282), .C2(n9714), .A(n9281), .B(n9285), .ZN(n9356)
         );
  MUX2_X1 U10485 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9356), .S(n9731), .Z(
        P1_U3554) );
  NAND3_X1 U10486 ( .A1(n9284), .A2(n9469), .A3(n9283), .ZN(n9286) );
  OAI211_X1 U10487 ( .C1(n9287), .C2(n9713), .A(n9286), .B(n9285), .ZN(n9357)
         );
  MUX2_X1 U10488 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9357), .S(n9731), .Z(
        P1_U3553) );
  OAI21_X1 U10489 ( .B1(n9292), .B2(n9349), .A(n9291), .ZN(n9358) );
  MUX2_X1 U10490 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9358), .S(n9731), .Z(
        P1_U3552) );
  AOI211_X1 U10491 ( .C1(n9345), .C2(n9295), .A(n9294), .B(n9293), .ZN(n9296)
         );
  OAI21_X1 U10492 ( .B1(n9297), .B2(n9349), .A(n9296), .ZN(n9360) );
  MUX2_X1 U10493 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9360), .S(n9731), .Z(
        P1_U3550) );
  AOI21_X1 U10494 ( .B1(n9345), .B2(n9299), .A(n9298), .ZN(n9300) );
  OAI211_X1 U10495 ( .C1(n9302), .C2(n9349), .A(n9301), .B(n9300), .ZN(n9361)
         );
  MUX2_X1 U10496 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9361), .S(n9731), .Z(
        P1_U3549) );
  AOI22_X1 U10497 ( .A1(n9304), .A2(n9469), .B1(n9345), .B2(n9303), .ZN(n9305)
         );
  OAI211_X1 U10498 ( .C1(n9307), .C2(n9349), .A(n9306), .B(n9305), .ZN(n9362)
         );
  MUX2_X1 U10499 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9362), .S(n9731), .Z(
        P1_U3548) );
  AOI21_X1 U10500 ( .B1(n9345), .B2(n9309), .A(n9308), .ZN(n9310) );
  OAI211_X1 U10501 ( .C1(n9312), .C2(n9349), .A(n9311), .B(n9310), .ZN(n9363)
         );
  MUX2_X1 U10502 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9363), .S(n9731), .Z(
        P1_U3547) );
  AOI22_X1 U10503 ( .A1(n9314), .A2(n9469), .B1(n9345), .B2(n9313), .ZN(n9315)
         );
  OAI211_X1 U10504 ( .C1(n9349), .C2(n9317), .A(n9316), .B(n9315), .ZN(n9364)
         );
  MUX2_X1 U10505 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9364), .S(n9731), .Z(
        P1_U3546) );
  AOI22_X1 U10506 ( .A1(n9319), .A2(n9469), .B1(n9345), .B2(n9318), .ZN(n9320)
         );
  OAI211_X1 U10507 ( .C1(n9322), .C2(n9349), .A(n9321), .B(n9320), .ZN(n9365)
         );
  MUX2_X1 U10508 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9365), .S(n9731), .Z(
        P1_U3545) );
  OR3_X1 U10509 ( .A1(n9324), .A2(n9323), .A3(n9349), .ZN(n9328) );
  NAND4_X1 U10510 ( .A1(n9328), .A2(n9327), .A3(n9326), .A4(n9325), .ZN(n9366)
         );
  MUX2_X1 U10511 ( .A(n9366), .B(P1_REG1_REG_21__SCAN_IN), .S(n9729), .Z(
        P1_U3544) );
  AOI211_X1 U10512 ( .C1(n9345), .C2(n9331), .A(n9330), .B(n9329), .ZN(n9332)
         );
  OAI21_X1 U10513 ( .B1(n9349), .B2(n9333), .A(n9332), .ZN(n9367) );
  MUX2_X1 U10514 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9367), .S(n9731), .Z(
        P1_U3543) );
  AOI22_X1 U10515 ( .A1(n9335), .A2(n9469), .B1(n9345), .B2(n9334), .ZN(n9336)
         );
  OAI211_X1 U10516 ( .C1(n9338), .C2(n9349), .A(n9337), .B(n9336), .ZN(n9368)
         );
  MUX2_X1 U10517 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9368), .S(n9731), .Z(
        P1_U3542) );
  OAI21_X1 U10518 ( .B1(n4447), .B2(n9713), .A(n9339), .ZN(n9340) );
  NOR2_X1 U10519 ( .A1(n9341), .A2(n9340), .ZN(n9342) );
  OAI21_X1 U10520 ( .B1(n9343), .B2(n9349), .A(n9342), .ZN(n9369) );
  MUX2_X1 U10521 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n9369), .S(n9731), .Z(
        P1_U3541) );
  AOI22_X1 U10522 ( .A1(n9346), .A2(n9469), .B1(n9345), .B2(n9344), .ZN(n9347)
         );
  OAI211_X1 U10523 ( .C1(n9350), .C2(n9349), .A(n9348), .B(n9347), .ZN(n9370)
         );
  MUX2_X1 U10524 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9370), .S(n9731), .Z(
        P1_U3540) );
  NAND2_X1 U10525 ( .A1(n9351), .A2(n9718), .ZN(n9355) );
  NAND4_X1 U10526 ( .A1(n9355), .A2(n9354), .A3(n9353), .A4(n9352), .ZN(n9371)
         );
  MUX2_X1 U10527 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9371), .S(n9731), .Z(
        P1_U3539) );
  MUX2_X1 U10528 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9356), .S(n9722), .Z(
        P1_U3522) );
  MUX2_X1 U10529 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9357), .S(n9722), .Z(
        P1_U3521) );
  MUX2_X1 U10530 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9358), .S(n9722), .Z(
        P1_U3520) );
  MUX2_X1 U10531 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9359), .S(n9722), .Z(
        P1_U3519) );
  MUX2_X1 U10532 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9360), .S(n9722), .Z(
        P1_U3518) );
  MUX2_X1 U10533 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9361), .S(n9722), .Z(
        P1_U3517) );
  MUX2_X1 U10534 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9362), .S(n9722), .Z(
        P1_U3516) );
  MUX2_X1 U10535 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9363), .S(n9722), .Z(
        P1_U3515) );
  MUX2_X1 U10536 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9364), .S(n9722), .Z(
        P1_U3514) );
  MUX2_X1 U10537 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9365), .S(n9722), .Z(
        P1_U3513) );
  MUX2_X1 U10538 ( .A(n9366), .B(P1_REG0_REG_21__SCAN_IN), .S(n9720), .Z(
        P1_U3512) );
  MUX2_X1 U10539 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9367), .S(n9722), .Z(
        P1_U3511) );
  MUX2_X1 U10540 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9368), .S(n9722), .Z(
        P1_U3510) );
  MUX2_X1 U10541 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n9369), .S(n9722), .Z(
        P1_U3508) );
  MUX2_X1 U10542 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9370), .S(n9722), .Z(
        P1_U3505) );
  MUX2_X1 U10543 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9371), .S(n9722), .Z(
        P1_U3502) );
  MUX2_X1 U10544 ( .A(n9373), .B(P1_D_REG_0__SCAN_IN), .S(n9372), .Z(P1_U3440)
         );
  MUX2_X1 U10545 ( .A(n9374), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  AOI22_X1 U10546 ( .A1(n9376), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9388) );
  AOI211_X1 U10547 ( .C1(n9379), .C2(n9378), .A(n9377), .B(n9738), .ZN(n9380)
         );
  AOI21_X1 U10548 ( .B1(n9382), .B2(n9381), .A(n9380), .ZN(n9387) );
  OAI211_X1 U10549 ( .C1(n9385), .C2(n9384), .A(n9732), .B(n9383), .ZN(n9386)
         );
  NAND3_X1 U10550 ( .A1(n9388), .A2(n9387), .A3(n9386), .ZN(P2_U3247) );
  INV_X1 U10551 ( .A(n9389), .ZN(n9704) );
  OAI21_X1 U10552 ( .B1(n4455), .B2(n9713), .A(n9391), .ZN(n9392) );
  AOI21_X1 U10553 ( .B1(n9393), .B2(n9704), .A(n9392), .ZN(n9394) );
  AND2_X1 U10554 ( .A1(n9395), .A2(n9394), .ZN(n9397) );
  INV_X1 U10555 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n9396) );
  AOI22_X1 U10556 ( .A1(n9722), .A2(n9397), .B1(n9396), .B2(n9720), .ZN(
        P1_U3484) );
  AOI22_X1 U10557 ( .A1(n9731), .A2(n9397), .B1(n6226), .B2(n9729), .ZN(
        P1_U3533) );
  NOR2_X1 U10558 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9398) );
  AOI21_X1 U10559 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9398), .ZN(n9893) );
  NOR2_X1 U10560 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9399) );
  AOI21_X1 U10561 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9399), .ZN(n9896) );
  NOR2_X1 U10562 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9400) );
  AOI21_X1 U10563 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9400), .ZN(n9899) );
  NOR2_X1 U10564 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9401) );
  AOI21_X1 U10565 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9401), .ZN(n9902) );
  NOR2_X1 U10566 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9402) );
  AOI21_X1 U10567 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9402), .ZN(n9905) );
  NOR2_X1 U10568 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n9408) );
  XNOR2_X1 U10569 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10080) );
  NAND2_X1 U10570 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9406) );
  XOR2_X1 U10571 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(P2_ADDR_REG_3__SCAN_IN), .Z(
        n10078) );
  NAND2_X1 U10572 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9404) );
  XOR2_X1 U10573 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10076) );
  AOI21_X1 U10574 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9886) );
  NAND3_X1 U10575 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n9888) );
  OAI21_X1 U10576 ( .B1(n9886), .B2(n6003), .A(n9888), .ZN(n10075) );
  NAND2_X1 U10577 ( .A1(n10076), .A2(n10075), .ZN(n9403) );
  NAND2_X1 U10578 ( .A1(n9404), .A2(n9403), .ZN(n10077) );
  NAND2_X1 U10579 ( .A1(n10078), .A2(n10077), .ZN(n9405) );
  NAND2_X1 U10580 ( .A1(n9406), .A2(n9405), .ZN(n10079) );
  NOR2_X1 U10581 ( .A1(n10080), .A2(n10079), .ZN(n9407) );
  NOR2_X1 U10582 ( .A1(n9408), .A2(n9407), .ZN(n9409) );
  NOR2_X1 U10583 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9409), .ZN(n10064) );
  AND2_X1 U10584 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9409), .ZN(n10065) );
  NOR2_X1 U10585 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10065), .ZN(n9410) );
  NOR2_X1 U10586 ( .A1(n10064), .A2(n9410), .ZN(n9411) );
  NAND2_X1 U10587 ( .A1(n9411), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9413) );
  XOR2_X1 U10588 ( .A(n9411), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10062) );
  NAND2_X1 U10589 ( .A1(n10062), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9412) );
  NAND2_X1 U10590 ( .A1(n9413), .A2(n9412), .ZN(n9414) );
  NAND2_X1 U10591 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9414), .ZN(n9416) );
  XOR2_X1 U10592 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9414), .Z(n10061) );
  NAND2_X1 U10593 ( .A1(n10061), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n9415) );
  NAND2_X1 U10594 ( .A1(n9416), .A2(n9415), .ZN(n9417) );
  NAND2_X1 U10595 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9417), .ZN(n9419) );
  XOR2_X1 U10596 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n9417), .Z(n10063) );
  NAND2_X1 U10597 ( .A1(n10063), .A2(P2_ADDR_REG_8__SCAN_IN), .ZN(n9418) );
  NAND2_X1 U10598 ( .A1(n9419), .A2(n9418), .ZN(n9420) );
  AND2_X1 U10599 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9420), .ZN(n9421) );
  INV_X1 U10600 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10074) );
  XNOR2_X1 U10601 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n9420), .ZN(n10073) );
  NOR2_X1 U10602 ( .A1(n10074), .A2(n10073), .ZN(n10072) );
  NOR2_X1 U10603 ( .A1(n9421), .A2(n10072), .ZN(n9914) );
  NAND2_X1 U10604 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9422) );
  OAI21_X1 U10605 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9422), .ZN(n9913) );
  NOR2_X1 U10606 ( .A1(n9914), .A2(n9913), .ZN(n9912) );
  AOI21_X1 U10607 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n9912), .ZN(n9911) );
  NAND2_X1 U10608 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9423) );
  OAI21_X1 U10609 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9423), .ZN(n9910) );
  NOR2_X1 U10610 ( .A1(n9911), .A2(n9910), .ZN(n9909) );
  AOI21_X1 U10611 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n9909), .ZN(n9908) );
  NOR2_X1 U10612 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9424) );
  AOI21_X1 U10613 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9424), .ZN(n9907) );
  NAND2_X1 U10614 ( .A1(n9908), .A2(n9907), .ZN(n9906) );
  OAI21_X1 U10615 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n9906), .ZN(n9904) );
  NAND2_X1 U10616 ( .A1(n9905), .A2(n9904), .ZN(n9903) );
  OAI21_X1 U10617 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n9903), .ZN(n9901) );
  NAND2_X1 U10618 ( .A1(n9902), .A2(n9901), .ZN(n9900) );
  OAI21_X1 U10619 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n9900), .ZN(n9898) );
  NAND2_X1 U10620 ( .A1(n9899), .A2(n9898), .ZN(n9897) );
  OAI21_X1 U10621 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n9897), .ZN(n9895) );
  NAND2_X1 U10622 ( .A1(n9896), .A2(n9895), .ZN(n9894) );
  OAI21_X1 U10623 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n9894), .ZN(n9892) );
  NAND2_X1 U10624 ( .A1(n9893), .A2(n9892), .ZN(n9891) );
  OAI21_X1 U10625 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n9891), .ZN(n10069) );
  NOR2_X1 U10626 ( .A1(n10070), .A2(n10069), .ZN(n9425) );
  NAND2_X1 U10627 ( .A1(n10070), .A2(n10069), .ZN(n10068) );
  OAI21_X1 U10628 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9425), .A(n10068), .ZN(
        n9427) );
  XOR2_X1 U10629 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .Z(n9426) );
  XNOR2_X1 U10630 ( .A(n9427), .B(n9426), .ZN(ADD_1071_U4) );
  OAI21_X1 U10631 ( .B1(n9429), .B2(n9859), .A(n9428), .ZN(n9431) );
  AOI211_X1 U10632 ( .C1(n9866), .C2(n9432), .A(n9431), .B(n9430), .ZN(n9459)
         );
  AOI22_X1 U10633 ( .A1(n4256), .A2(n9459), .B1(n8421), .B2(n9884), .ZN(
        P2_U3537) );
  INV_X1 U10634 ( .A(n9433), .ZN(n9440) );
  AND3_X1 U10635 ( .A1(n9435), .A2(n9866), .A3(n9434), .ZN(n9439) );
  OAI22_X1 U10636 ( .A1(n9437), .A2(n9861), .B1(n9436), .B2(n9859), .ZN(n9438)
         );
  NOR3_X1 U10637 ( .A1(n9440), .A2(n9439), .A3(n9438), .ZN(n9460) );
  AOI22_X1 U10638 ( .A1(n4256), .A2(n9460), .B1(n8398), .B2(n9884), .ZN(
        P2_U3536) );
  OAI21_X1 U10639 ( .B1(n9442), .B2(n9859), .A(n9441), .ZN(n9444) );
  AOI211_X1 U10640 ( .C1(n9445), .C2(n9866), .A(n9444), .B(n9443), .ZN(n9462)
         );
  AOI22_X1 U10641 ( .A1(n4256), .A2(n9462), .B1(n8396), .B2(n9884), .ZN(
        P2_U3535) );
  OAI22_X1 U10642 ( .A1(n9447), .A2(n9861), .B1(n9446), .B2(n9859), .ZN(n9449)
         );
  AOI211_X1 U10643 ( .C1(n9866), .C2(n9450), .A(n9449), .B(n9448), .ZN(n9464)
         );
  AOI22_X1 U10644 ( .A1(n4256), .A2(n9464), .B1(n5046), .B2(n9884), .ZN(
        P2_U3534) );
  NOR2_X1 U10645 ( .A1(n9451), .A2(n9807), .ZN(n9457) );
  OAI22_X1 U10646 ( .A1(n9453), .A2(n9861), .B1(n9452), .B2(n9859), .ZN(n9455)
         );
  AOI211_X1 U10647 ( .C1(n9457), .C2(n9456), .A(n9455), .B(n9454), .ZN(n9465)
         );
  AOI22_X1 U10648 ( .A1(n4256), .A2(n9465), .B1(n5018), .B2(n9884), .ZN(
        P2_U3533) );
  INV_X1 U10649 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9458) );
  AOI22_X1 U10650 ( .A1(n4255), .A2(n9459), .B1(n9458), .B2(n9867), .ZN(
        P2_U3502) );
  AOI22_X1 U10651 ( .A1(n4255), .A2(n9460), .B1(n5098), .B2(n9867), .ZN(
        P2_U3499) );
  INV_X1 U10652 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n9461) );
  AOI22_X1 U10653 ( .A1(n4255), .A2(n9462), .B1(n9461), .B2(n9867), .ZN(
        P2_U3496) );
  INV_X1 U10654 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9463) );
  AOI22_X1 U10655 ( .A1(n4255), .A2(n9464), .B1(n9463), .B2(n9867), .ZN(
        P2_U3493) );
  INV_X1 U10656 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9930) );
  AOI22_X1 U10657 ( .A1(n4255), .A2(n9465), .B1(n9930), .B2(n9867), .ZN(
        P2_U3490) );
  INV_X1 U10658 ( .A(n9466), .ZN(n9482) );
  XNOR2_X1 U10659 ( .A(n9468), .B(n9467), .ZN(n9492) );
  OAI211_X1 U10660 ( .C1(n9471), .C2(n9490), .A(n9470), .B(n9469), .ZN(n9488)
         );
  OAI22_X1 U10661 ( .A1(n9488), .A2(n9473), .B1(n9490), .B2(n9472), .ZN(n9481)
         );
  OAI21_X1 U10662 ( .B1(n9476), .B2(n9475), .A(n9474), .ZN(n9479) );
  AOI222_X1 U10663 ( .A1(n9651), .A2(n9479), .B1(n9478), .B2(n9656), .C1(n9477), .C2(n9654), .ZN(n9489) );
  INV_X1 U10664 ( .A(n9489), .ZN(n9480) );
  AOI211_X1 U10665 ( .C1(n9482), .C2(n9492), .A(n9481), .B(n9480), .ZN(n9487)
         );
  INV_X1 U10666 ( .A(n9483), .ZN(n9485) );
  AOI22_X1 U10667 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n9676), .B1(n9485), .B2(
        n9484), .ZN(n9486) );
  OAI21_X1 U10668 ( .B1(n9676), .B2(n9487), .A(n9486), .ZN(P1_U3276) );
  OAI211_X1 U10669 ( .C1(n9490), .C2(n9713), .A(n9489), .B(n9488), .ZN(n9491)
         );
  AOI21_X1 U10670 ( .B1(n9718), .B2(n9492), .A(n9491), .ZN(n9504) );
  AOI22_X1 U10671 ( .A1(n9731), .A2(n9504), .B1(n5728), .B2(n9729), .ZN(
        P1_U3538) );
  OAI211_X1 U10672 ( .C1(n9495), .C2(n9713), .A(n9494), .B(n9493), .ZN(n9496)
         );
  AOI21_X1 U10673 ( .B1(n9718), .B2(n9497), .A(n9496), .ZN(n9505) );
  AOI22_X1 U10674 ( .A1(n9731), .A2(n9505), .B1(n6835), .B2(n9729), .ZN(
        P1_U3537) );
  OAI211_X1 U10675 ( .C1(n9500), .C2(n9713), .A(n9499), .B(n9498), .ZN(n9501)
         );
  AOI21_X1 U10676 ( .B1(n9502), .B2(n9718), .A(n9501), .ZN(n9506) );
  AOI22_X1 U10677 ( .A1(n9731), .A2(n9506), .B1(n6837), .B2(n9729), .ZN(
        P1_U3535) );
  INV_X1 U10678 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n9503) );
  AOI22_X1 U10679 ( .A1(n9722), .A2(n9504), .B1(n9503), .B2(n9720), .ZN(
        P1_U3499) );
  AOI22_X1 U10680 ( .A1(n9722), .A2(n9505), .B1(n5690), .B2(n9720), .ZN(
        P1_U3496) );
  AOI22_X1 U10681 ( .A1(n9722), .A2(n9506), .B1(n5679), .B2(n9720), .ZN(
        P1_U3490) );
  XNOR2_X1 U10682 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U10683 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U10684 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10066) );
  OAI21_X1 U10685 ( .B1(n9509), .B2(n9508), .A(n9507), .ZN(n9513) );
  NOR2_X1 U10686 ( .A1(n9523), .A2(n9510), .ZN(n9511) );
  AOI211_X1 U10687 ( .C1(n9526), .C2(n9513), .A(n9512), .B(n9511), .ZN(n9518)
         );
  OAI211_X1 U10688 ( .C1(n9516), .C2(n9515), .A(n9622), .B(n9514), .ZN(n9517)
         );
  OAI211_X1 U10689 ( .C1(n10066), .C2(n9643), .A(n9518), .B(n9517), .ZN(
        P1_U3246) );
  INV_X1 U10690 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9533) );
  OAI21_X1 U10691 ( .B1(n9521), .B2(n9520), .A(n9519), .ZN(n9527) );
  NOR2_X1 U10692 ( .A1(n9523), .A2(n9522), .ZN(n9524) );
  AOI211_X1 U10693 ( .C1(n9527), .C2(n9526), .A(n9525), .B(n9524), .ZN(n9532)
         );
  OAI211_X1 U10694 ( .C1(n9530), .C2(n9529), .A(n9622), .B(n9528), .ZN(n9531)
         );
  OAI211_X1 U10695 ( .C1(n9533), .C2(n9643), .A(n9532), .B(n9531), .ZN(
        P1_U3249) );
  AOI211_X1 U10696 ( .C1(n9536), .C2(n9535), .A(n9534), .B(n9628), .ZN(n9537)
         );
  AOI211_X1 U10697 ( .C1(n9634), .C2(n9539), .A(n9538), .B(n9537), .ZN(n9545)
         );
  AOI21_X1 U10698 ( .B1(n9542), .B2(n9541), .A(n9540), .ZN(n9543) );
  OR2_X1 U10699 ( .A1(n9640), .A2(n9543), .ZN(n9544) );
  OAI211_X1 U10700 ( .C1(n10074), .C2(n9643), .A(n9545), .B(n9544), .ZN(
        P1_U3250) );
  INV_X1 U10701 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n9558) );
  AOI211_X1 U10702 ( .C1(n9548), .C2(n9547), .A(n9546), .B(n9628), .ZN(n9549)
         );
  AOI211_X1 U10703 ( .C1(n9634), .C2(n9551), .A(n9550), .B(n9549), .ZN(n9557)
         );
  AOI21_X1 U10704 ( .B1(n9554), .B2(n9553), .A(n9552), .ZN(n9555) );
  OR2_X1 U10705 ( .A1(n9640), .A2(n9555), .ZN(n9556) );
  OAI211_X1 U10706 ( .C1(n9558), .C2(n9643), .A(n9557), .B(n9556), .ZN(
        P1_U3251) );
  INV_X1 U10707 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9575) );
  INV_X1 U10708 ( .A(n9559), .ZN(n9563) );
  INV_X1 U10709 ( .A(n9560), .ZN(n9561) );
  AOI211_X1 U10710 ( .C1(n9563), .C2(n9562), .A(n9561), .B(n9628), .ZN(n9564)
         );
  AOI211_X1 U10711 ( .C1(n9634), .C2(n9566), .A(n9565), .B(n9564), .ZN(n9574)
         );
  INV_X1 U10712 ( .A(n9567), .ZN(n9570) );
  INV_X1 U10713 ( .A(n9568), .ZN(n9569) );
  NOR2_X1 U10714 ( .A1(n9570), .A2(n9569), .ZN(n9571) );
  OAI21_X1 U10715 ( .B1(n9572), .B2(n9571), .A(n9622), .ZN(n9573) );
  OAI211_X1 U10716 ( .C1(n9575), .C2(n9643), .A(n9574), .B(n9573), .ZN(
        P1_U3253) );
  INV_X1 U10717 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9590) );
  INV_X1 U10718 ( .A(n9576), .ZN(n9580) );
  INV_X1 U10719 ( .A(n9577), .ZN(n9579) );
  AOI211_X1 U10720 ( .C1(n9580), .C2(n9579), .A(n9578), .B(n9628), .ZN(n9581)
         );
  AOI211_X1 U10721 ( .C1(n9634), .C2(n9583), .A(n9582), .B(n9581), .ZN(n9589)
         );
  AOI21_X1 U10722 ( .B1(n9586), .B2(n9585), .A(n9584), .ZN(n9587) );
  OR2_X1 U10723 ( .A1(n9640), .A2(n9587), .ZN(n9588) );
  OAI211_X1 U10724 ( .C1(n9590), .C2(n9643), .A(n9589), .B(n9588), .ZN(
        P1_U3254) );
  INV_X1 U10725 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n9601) );
  AOI211_X1 U10726 ( .C1(n9593), .C2(n9592), .A(n9591), .B(n9628), .ZN(n9594)
         );
  AOI211_X1 U10727 ( .C1(n9634), .C2(n9596), .A(n9595), .B(n9594), .ZN(n9600)
         );
  OAI211_X1 U10728 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9598), .A(n9622), .B(
        n9597), .ZN(n9599) );
  OAI211_X1 U10729 ( .C1(n9601), .C2(n9643), .A(n9600), .B(n9599), .ZN(
        P1_U3256) );
  INV_X1 U10730 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9613) );
  AOI211_X1 U10731 ( .C1(n9604), .C2(n9603), .A(n9602), .B(n9628), .ZN(n9605)
         );
  AOI211_X1 U10732 ( .C1(n9634), .C2(n9607), .A(n9606), .B(n9605), .ZN(n9612)
         );
  OAI211_X1 U10733 ( .C1(n9610), .C2(n9609), .A(n9622), .B(n9608), .ZN(n9611)
         );
  OAI211_X1 U10734 ( .C1(n9613), .C2(n9643), .A(n9612), .B(n9611), .ZN(
        P1_U3257) );
  INV_X1 U10735 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10028) );
  INV_X1 U10736 ( .A(n9614), .ZN(n9619) );
  AOI211_X1 U10737 ( .C1(n9617), .C2(n9616), .A(n9615), .B(n9628), .ZN(n9618)
         );
  AOI211_X1 U10738 ( .C1(n9620), .C2(n9634), .A(n9619), .B(n9618), .ZN(n9626)
         );
  OAI211_X1 U10739 ( .C1(n9624), .C2(n9623), .A(n9622), .B(n9621), .ZN(n9625)
         );
  OAI211_X1 U10740 ( .C1(n10028), .C2(n9643), .A(n9626), .B(n9625), .ZN(
        P1_U3258) );
  INV_X1 U10741 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9644) );
  INV_X1 U10742 ( .A(n9627), .ZN(n9633) );
  AOI211_X1 U10743 ( .C1(n9631), .C2(n9630), .A(n9629), .B(n9628), .ZN(n9632)
         );
  AOI211_X1 U10744 ( .C1(n9635), .C2(n9634), .A(n9633), .B(n9632), .ZN(n9642)
         );
  AOI21_X1 U10745 ( .B1(n9638), .B2(n9637), .A(n9636), .ZN(n9639) );
  OR2_X1 U10746 ( .A1(n9640), .A2(n9639), .ZN(n9641) );
  OAI211_X1 U10747 ( .C1(n9644), .C2(n9643), .A(n9642), .B(n9641), .ZN(
        P1_U3259) );
  XOR2_X1 U10748 ( .A(n9648), .B(n9645), .Z(n9719) );
  NAND2_X1 U10749 ( .A1(n9647), .A2(n9646), .ZN(n9650) );
  INV_X1 U10750 ( .A(n9648), .ZN(n9649) );
  XNOR2_X1 U10751 ( .A(n9650), .B(n9649), .ZN(n9652) );
  NAND2_X1 U10752 ( .A1(n9652), .A2(n9651), .ZN(n9658) );
  AOI22_X1 U10753 ( .A1(n9656), .A2(n9655), .B1(n9654), .B2(n9653), .ZN(n9657)
         );
  NAND2_X1 U10754 ( .A1(n9658), .A2(n9657), .ZN(n9717) );
  AOI21_X1 U10755 ( .B1(n9719), .B2(n9659), .A(n9717), .ZN(n9675) );
  INV_X1 U10756 ( .A(n9660), .ZN(n9662) );
  OAI21_X1 U10757 ( .B1(n9662), .B2(n4456), .A(n9661), .ZN(n9715) );
  OAI22_X1 U10758 ( .A1(n9666), .A2(n9665), .B1(n9664), .B2(n9663), .ZN(n9667)
         );
  AOI21_X1 U10759 ( .B1(n9669), .B2(n9668), .A(n9667), .ZN(n9670) );
  OAI21_X1 U10760 ( .B1(n9715), .B2(n9671), .A(n9670), .ZN(n9672) );
  AOI21_X1 U10761 ( .B1(n9719), .B2(n9673), .A(n9672), .ZN(n9674) );
  OAI21_X1 U10762 ( .B1(n9676), .B2(n9675), .A(n9674), .ZN(P1_U3282) );
  AND2_X1 U10763 ( .A1(n9678), .A2(n9677), .ZN(n9679) );
  AND2_X1 U10764 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9680), .ZN(P1_U3292) );
  AND2_X1 U10765 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9680), .ZN(P1_U3293) );
  AND2_X1 U10766 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n9680), .ZN(P1_U3294) );
  AND2_X1 U10767 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9680), .ZN(P1_U3295) );
  AND2_X1 U10768 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n9680), .ZN(P1_U3296) );
  AND2_X1 U10769 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9680), .ZN(P1_U3297) );
  AND2_X1 U10770 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9680), .ZN(P1_U3298) );
  AND2_X1 U10771 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9680), .ZN(P1_U3299) );
  AND2_X1 U10772 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9680), .ZN(P1_U3300) );
  AND2_X1 U10773 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9680), .ZN(P1_U3301) );
  AND2_X1 U10774 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9680), .ZN(P1_U3302) );
  AND2_X1 U10775 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n9680), .ZN(P1_U3303) );
  INV_X1 U10776 ( .A(P1_D_REG_19__SCAN_IN), .ZN(n9952) );
  NOR2_X1 U10777 ( .A1(n9679), .A2(n9952), .ZN(P1_U3304) );
  AND2_X1 U10778 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9680), .ZN(P1_U3305) );
  AND2_X1 U10779 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9680), .ZN(P1_U3306) );
  AND2_X1 U10780 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n9680), .ZN(P1_U3307) );
  AND2_X1 U10781 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9680), .ZN(P1_U3308) );
  AND2_X1 U10782 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9680), .ZN(P1_U3309) );
  INV_X1 U10783 ( .A(P1_D_REG_13__SCAN_IN), .ZN(n9970) );
  NOR2_X1 U10784 ( .A1(n9679), .A2(n9970), .ZN(P1_U3310) );
  AND2_X1 U10785 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9680), .ZN(P1_U3311) );
  AND2_X1 U10786 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n9680), .ZN(P1_U3312) );
  AND2_X1 U10787 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9680), .ZN(P1_U3313) );
  AND2_X1 U10788 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9680), .ZN(P1_U3314) );
  AND2_X1 U10789 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9680), .ZN(P1_U3315) );
  AND2_X1 U10790 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9680), .ZN(P1_U3316) );
  AND2_X1 U10791 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9680), .ZN(P1_U3317) );
  AND2_X1 U10792 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9680), .ZN(P1_U3318) );
  AND2_X1 U10793 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9680), .ZN(P1_U3319) );
  INV_X1 U10794 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n9960) );
  NOR2_X1 U10795 ( .A1(n9679), .A2(n9960), .ZN(P1_U3320) );
  AND2_X1 U10796 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9680), .ZN(P1_U3321) );
  INV_X1 U10797 ( .A(n9681), .ZN(n9686) );
  OAI21_X1 U10798 ( .B1(n9683), .B2(n9713), .A(n9682), .ZN(n9685) );
  AOI211_X1 U10799 ( .C1(n9686), .C2(n9718), .A(n9685), .B(n9684), .ZN(n9724)
         );
  AOI22_X1 U10800 ( .A1(n9722), .A2(n9724), .B1(n5517), .B2(n9720), .ZN(
        P1_U3457) );
  AOI22_X1 U10801 ( .A1(n9722), .A2(n9687), .B1(n5536), .B2(n9720), .ZN(
        P1_U3460) );
  OAI22_X1 U10802 ( .A1(n9689), .A2(n9714), .B1(n9688), .B2(n9713), .ZN(n9691)
         );
  AOI211_X1 U10803 ( .C1(n9704), .C2(n9692), .A(n9691), .B(n9690), .ZN(n9725)
         );
  AOI22_X1 U10804 ( .A1(n9722), .A2(n9725), .B1(n5564), .B2(n9720), .ZN(
        P1_U3466) );
  OAI21_X1 U10805 ( .B1(n9694), .B2(n9713), .A(n9693), .ZN(n9695) );
  AOI211_X1 U10806 ( .C1(n9697), .C2(n9718), .A(n9696), .B(n9695), .ZN(n9726)
         );
  AOI22_X1 U10807 ( .A1(n9722), .A2(n9726), .B1(n5582), .B2(n9720), .ZN(
        P1_U3469) );
  INV_X1 U10808 ( .A(n9698), .ZN(n9703) );
  OAI22_X1 U10809 ( .A1(n9700), .A2(n9714), .B1(n9699), .B2(n9713), .ZN(n9702)
         );
  AOI211_X1 U10810 ( .C1(n9704), .C2(n9703), .A(n9702), .B(n9701), .ZN(n9727)
         );
  AOI22_X1 U10811 ( .A1(n9722), .A2(n9727), .B1(n5593), .B2(n9720), .ZN(
        P1_U3472) );
  NAND2_X1 U10812 ( .A1(n9705), .A2(n9718), .ZN(n9711) );
  OAI21_X1 U10813 ( .B1(n9707), .B2(n9714), .A(n9706), .ZN(n9708) );
  NOR2_X1 U10814 ( .A1(n9709), .A2(n9708), .ZN(n9710) );
  AND2_X1 U10815 ( .A1(n9711), .A2(n9710), .ZN(n9728) );
  INV_X1 U10816 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n9712) );
  AOI22_X1 U10817 ( .A1(n9722), .A2(n9728), .B1(n9712), .B2(n9720), .ZN(
        P1_U3478) );
  OAI22_X1 U10818 ( .A1(n9715), .A2(n9714), .B1(n4456), .B2(n9713), .ZN(n9716)
         );
  AOI211_X1 U10819 ( .C1(n9719), .C2(n9718), .A(n9717), .B(n9716), .ZN(n9730)
         );
  INV_X1 U10820 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n9721) );
  AOI22_X1 U10821 ( .A1(n9722), .A2(n9730), .B1(n9721), .B2(n9720), .ZN(
        P1_U3481) );
  AOI22_X1 U10822 ( .A1(n9731), .A2(n9724), .B1(n9723), .B2(n9729), .ZN(
        P1_U3524) );
  AOI22_X1 U10823 ( .A1(n9731), .A2(n9725), .B1(n5565), .B2(n9729), .ZN(
        P1_U3527) );
  AOI22_X1 U10824 ( .A1(n9731), .A2(n9726), .B1(n6057), .B2(n9729), .ZN(
        P1_U3528) );
  AOI22_X1 U10825 ( .A1(n9731), .A2(n9727), .B1(n6060), .B2(n9729), .ZN(
        P1_U3529) );
  AOI22_X1 U10826 ( .A1(n9731), .A2(n9728), .B1(n6222), .B2(n9729), .ZN(
        P1_U3531) );
  AOI22_X1 U10827 ( .A1(n9731), .A2(n9730), .B1(n6224), .B2(n9729), .ZN(
        P1_U3532) );
  AOI22_X1 U10828 ( .A1(n9733), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n9732), .ZN(n9745) );
  INV_X1 U10829 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n9735) );
  OAI22_X1 U10830 ( .A1(n9736), .A2(n9735), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9734), .ZN(n9737) );
  INV_X1 U10831 ( .A(n9737), .ZN(n9744) );
  NOR2_X1 U10832 ( .A1(n9738), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n9742) );
  OAI21_X1 U10833 ( .B1(n9740), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9739), .ZN(
        n9741) );
  OAI21_X1 U10834 ( .B1(n9742), .B2(n9741), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n9743) );
  OAI211_X1 U10835 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n9745), .A(n9744), .B(
        n9743), .ZN(P2_U3245) );
  XNOR2_X1 U10836 ( .A(n9746), .B(n9752), .ZN(n9749) );
  AOI21_X1 U10837 ( .B1(n9749), .B2(n9748), .A(n9747), .ZN(n9780) );
  AOI22_X1 U10838 ( .A1(n9750), .A2(P2_REG3_REG_1__SCAN_IN), .B1(
        P2_REG2_REG_1__SCAN_IN), .B2(n9762), .ZN(n9761) );
  XNOR2_X1 U10839 ( .A(n9752), .B(n9751), .ZN(n9783) );
  NAND2_X1 U10840 ( .A1(n9753), .A2(n9783), .ZN(n9757) );
  XNOR2_X1 U10841 ( .A(n9754), .B(n9778), .ZN(n9777) );
  NAND2_X1 U10842 ( .A1(n9755), .A2(n9777), .ZN(n9756) );
  OAI211_X1 U10843 ( .C1(n9778), .C2(n9758), .A(n9757), .B(n9756), .ZN(n9759)
         );
  INV_X1 U10844 ( .A(n9759), .ZN(n9760) );
  OAI211_X1 U10845 ( .C1(n9762), .C2(n9780), .A(n9761), .B(n9760), .ZN(
        P2_U3295) );
  NOR2_X1 U10846 ( .A1(n9764), .A2(n9763), .ZN(n9765) );
  INV_X1 U10847 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n9982) );
  NOR2_X1 U10848 ( .A1(n9765), .A2(n9982), .ZN(P2_U3297) );
  AND2_X1 U10849 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10021), .ZN(P2_U3298) );
  AND2_X1 U10850 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10021), .ZN(P2_U3299) );
  AND2_X1 U10851 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10021), .ZN(P2_U3300) );
  AND2_X1 U10852 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10021), .ZN(P2_U3301) );
  AND2_X1 U10853 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10021), .ZN(P2_U3302) );
  INV_X1 U10854 ( .A(P2_D_REG_25__SCAN_IN), .ZN(n9955) );
  NOR2_X1 U10855 ( .A1(n9765), .A2(n9955), .ZN(P2_U3303) );
  AND2_X1 U10856 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10021), .ZN(P2_U3304) );
  AND2_X1 U10857 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10021), .ZN(P2_U3305) );
  AND2_X1 U10858 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10021), .ZN(P2_U3306) );
  AND2_X1 U10859 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10021), .ZN(P2_U3307) );
  AND2_X1 U10860 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10021), .ZN(P2_U3308) );
  AND2_X1 U10861 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10021), .ZN(P2_U3309) );
  AND2_X1 U10862 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10021), .ZN(P2_U3311) );
  AND2_X1 U10863 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10021), .ZN(P2_U3312) );
  AND2_X1 U10864 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10021), .ZN(P2_U3313) );
  INV_X1 U10865 ( .A(P2_D_REG_14__SCAN_IN), .ZN(n10033) );
  NOR2_X1 U10866 ( .A1(n9765), .A2(n10033), .ZN(P2_U3314) );
  AND2_X1 U10867 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10021), .ZN(P2_U3315) );
  AND2_X1 U10868 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10021), .ZN(P2_U3316) );
  AND2_X1 U10869 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10021), .ZN(P2_U3317) );
  AND2_X1 U10870 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10021), .ZN(P2_U3318) );
  AND2_X1 U10871 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10021), .ZN(P2_U3319) );
  AND2_X1 U10872 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10021), .ZN(P2_U3320) );
  AND2_X1 U10873 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10021), .ZN(P2_U3321) );
  AND2_X1 U10874 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10021), .ZN(P2_U3322) );
  AND2_X1 U10875 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10021), .ZN(P2_U3323) );
  AND2_X1 U10876 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10021), .ZN(P2_U3324) );
  AND2_X1 U10877 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10021), .ZN(P2_U3325) );
  AND2_X1 U10878 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10021), .ZN(P2_U3326) );
  NOR2_X1 U10879 ( .A1(n9766), .A2(P2_U3152), .ZN(n9770) );
  AOI22_X1 U10880 ( .A1(n9768), .A2(n9770), .B1(n9767), .B2(n10021), .ZN(
        P2_U3437) );
  AOI22_X1 U10881 ( .A1(n9771), .A2(n9770), .B1(n9769), .B2(n10021), .ZN(
        P2_U3438) );
  OAI22_X1 U10882 ( .A1(n9774), .A2(n9807), .B1(n9773), .B2(n9772), .ZN(n9775)
         );
  NOR2_X1 U10883 ( .A1(n9776), .A2(n9775), .ZN(n9869) );
  INV_X1 U10884 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n9934) );
  AOI22_X1 U10885 ( .A1(n4255), .A2(n9869), .B1(n9934), .B2(n9867), .ZN(
        P2_U3451) );
  INV_X1 U10886 ( .A(n9777), .ZN(n9779) );
  OAI22_X1 U10887 ( .A1(n9779), .A2(n9861), .B1(n9778), .B2(n9859), .ZN(n9782)
         );
  INV_X1 U10888 ( .A(n9780), .ZN(n9781) );
  AOI211_X1 U10889 ( .C1(n9866), .C2(n9783), .A(n9782), .B(n9781), .ZN(n9871)
         );
  INV_X1 U10890 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n9784) );
  AOI22_X1 U10891 ( .A1(n4255), .A2(n9871), .B1(n9784), .B2(n9867), .ZN(
        P2_U3454) );
  AOI21_X1 U10892 ( .B1(n9843), .B2(n9786), .A(n9785), .ZN(n9787) );
  OAI211_X1 U10893 ( .C1(n9807), .C2(n9789), .A(n9788), .B(n9787), .ZN(n9790)
         );
  INV_X1 U10894 ( .A(n9790), .ZN(n9872) );
  AOI22_X1 U10895 ( .A1(n4255), .A2(n9872), .B1(n4727), .B2(n9867), .ZN(
        P2_U3457) );
  INV_X1 U10896 ( .A(n9791), .ZN(n9853) );
  INV_X1 U10897 ( .A(n9796), .ZN(n9798) );
  AOI21_X1 U10898 ( .B1(n9843), .B2(n9793), .A(n9792), .ZN(n9794) );
  OAI211_X1 U10899 ( .C1(n9847), .C2(n9796), .A(n9795), .B(n9794), .ZN(n9797)
         );
  AOI21_X1 U10900 ( .B1(n9853), .B2(n9798), .A(n9797), .ZN(n9873) );
  INV_X1 U10901 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9799) );
  AOI22_X1 U10902 ( .A1(n4255), .A2(n9873), .B1(n9799), .B2(n9867), .ZN(
        P2_U3460) );
  INV_X1 U10903 ( .A(n9800), .ZN(n9806) );
  OAI22_X1 U10904 ( .A1(n9802), .A2(n9861), .B1(n9801), .B2(n9859), .ZN(n9805)
         );
  INV_X1 U10905 ( .A(n9803), .ZN(n9804) );
  AOI211_X1 U10906 ( .C1(n9866), .C2(n9806), .A(n9805), .B(n9804), .ZN(n9874)
         );
  AOI22_X1 U10907 ( .A1(n4255), .A2(n9874), .B1(n4815), .B2(n9867), .ZN(
        P2_U3463) );
  NOR2_X1 U10908 ( .A1(n9808), .A2(n9807), .ZN(n9812) );
  OAI21_X1 U10909 ( .B1(n9810), .B2(n9859), .A(n9809), .ZN(n9811) );
  NOR3_X1 U10910 ( .A1(n9813), .A2(n9812), .A3(n9811), .ZN(n9875) );
  INV_X1 U10911 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n9814) );
  AOI22_X1 U10912 ( .A1(n4255), .A2(n9875), .B1(n9814), .B2(n9867), .ZN(
        P2_U3466) );
  NAND3_X1 U10913 ( .A1(n9816), .A2(n9815), .A3(n9866), .ZN(n9818) );
  OAI211_X1 U10914 ( .C1(n9819), .C2(n9859), .A(n9818), .B(n9817), .ZN(n9820)
         );
  NOR2_X1 U10915 ( .A1(n9821), .A2(n9820), .ZN(n9876) );
  INV_X1 U10916 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9822) );
  AOI22_X1 U10917 ( .A1(n4255), .A2(n9876), .B1(n9822), .B2(n9867), .ZN(
        P2_U3469) );
  OAI22_X1 U10918 ( .A1(n9824), .A2(n9861), .B1(n9823), .B2(n9859), .ZN(n9826)
         );
  AOI211_X1 U10919 ( .C1(n9866), .C2(n9827), .A(n9826), .B(n9825), .ZN(n9877)
         );
  INV_X1 U10920 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9828) );
  AOI22_X1 U10921 ( .A1(n4255), .A2(n9877), .B1(n9828), .B2(n9867), .ZN(
        P2_U3472) );
  INV_X1 U10922 ( .A(n9847), .ZN(n9842) );
  INV_X1 U10923 ( .A(n9829), .ZN(n9834) );
  OAI22_X1 U10924 ( .A1(n9831), .A2(n9861), .B1(n9830), .B2(n9859), .ZN(n9833)
         );
  AOI211_X1 U10925 ( .C1(n9842), .C2(n9834), .A(n9833), .B(n9832), .ZN(n9878)
         );
  INV_X1 U10926 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n9835) );
  AOI22_X1 U10927 ( .A1(n4255), .A2(n9878), .B1(n9835), .B2(n9867), .ZN(
        P2_U3475) );
  INV_X1 U10928 ( .A(n9836), .ZN(n9841) );
  OAI22_X1 U10929 ( .A1(n9838), .A2(n9861), .B1(n9837), .B2(n9859), .ZN(n9840)
         );
  AOI211_X1 U10930 ( .C1(n9842), .C2(n9841), .A(n9840), .B(n9839), .ZN(n9880)
         );
  AOI22_X1 U10931 ( .A1(n4255), .A2(n9880), .B1(n4941), .B2(n9867), .ZN(
        P2_U3478) );
  INV_X1 U10932 ( .A(n9848), .ZN(n9852) );
  NAND2_X1 U10933 ( .A1(n9844), .A2(n9843), .ZN(n9846) );
  OAI211_X1 U10934 ( .C1(n9848), .C2(n9847), .A(n9846), .B(n9845), .ZN(n9851)
         );
  INV_X1 U10935 ( .A(n9849), .ZN(n9850) );
  AOI211_X1 U10936 ( .C1(n9853), .C2(n9852), .A(n9851), .B(n9850), .ZN(n9881)
         );
  AOI22_X1 U10937 ( .A1(n4255), .A2(n9881), .B1(n4971), .B2(n9867), .ZN(
        P2_U3481) );
  OAI22_X1 U10938 ( .A1(n9854), .A2(n9861), .B1(n4517), .B2(n9859), .ZN(n9857)
         );
  INV_X1 U10939 ( .A(n9855), .ZN(n9856) );
  AOI211_X1 U10940 ( .C1(n9858), .C2(n9866), .A(n9857), .B(n9856), .ZN(n9883)
         );
  AOI22_X1 U10941 ( .A1(n4255), .A2(n9883), .B1(n4991), .B2(n9867), .ZN(
        P2_U3484) );
  OAI22_X1 U10942 ( .A1(n9862), .A2(n9861), .B1(n9860), .B2(n9859), .ZN(n9864)
         );
  AOI211_X1 U10943 ( .C1(n9866), .C2(n9865), .A(n9864), .B(n9863), .ZN(n9885)
         );
  INV_X1 U10944 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10029) );
  AOI22_X1 U10945 ( .A1(n4255), .A2(n9885), .B1(n10029), .B2(n9867), .ZN(
        P2_U3487) );
  INV_X1 U10946 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n9868) );
  AOI22_X1 U10947 ( .A1(n4256), .A2(n9869), .B1(n9868), .B2(n9884), .ZN(
        P2_U3520) );
  AOI22_X1 U10948 ( .A1(n4256), .A2(n9871), .B1(n9870), .B2(n9884), .ZN(
        P2_U3521) );
  AOI22_X1 U10949 ( .A1(n4256), .A2(n9872), .B1(n6328), .B2(n9884), .ZN(
        P2_U3522) );
  AOI22_X1 U10950 ( .A1(n4256), .A2(n9873), .B1(n6325), .B2(n9884), .ZN(
        P2_U3523) );
  AOI22_X1 U10951 ( .A1(n4256), .A2(n9874), .B1(n6347), .B2(n9884), .ZN(
        P2_U3524) );
  AOI22_X1 U10952 ( .A1(n4256), .A2(n9875), .B1(n6344), .B2(n9884), .ZN(
        P2_U3525) );
  AOI22_X1 U10953 ( .A1(n4256), .A2(n9876), .B1(n6350), .B2(n9884), .ZN(
        P2_U3526) );
  AOI22_X1 U10954 ( .A1(n4256), .A2(n9877), .B1(n6343), .B2(n9884), .ZN(
        P2_U3527) );
  AOI22_X1 U10955 ( .A1(n4256), .A2(n9878), .B1(n6352), .B2(n9884), .ZN(
        P2_U3528) );
  AOI22_X1 U10956 ( .A1(n4256), .A2(n9880), .B1(n9879), .B2(n9884), .ZN(
        P2_U3529) );
  AOI22_X1 U10957 ( .A1(n4256), .A2(n9881), .B1(n6408), .B2(n9884), .ZN(
        P2_U3530) );
  AOI22_X1 U10958 ( .A1(n4256), .A2(n9883), .B1(n9882), .B2(n9884), .ZN(
        P2_U3531) );
  AOI22_X1 U10959 ( .A1(n4256), .A2(n9885), .B1(n6544), .B2(n9884), .ZN(
        P2_U3532) );
  INV_X1 U10960 ( .A(n9886), .ZN(n9887) );
  NAND2_X1 U10961 ( .A1(n9888), .A2(n9887), .ZN(n9889) );
  XNOR2_X1 U10962 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n9889), .ZN(ADD_1071_U5) );
  AOI22_X1 U10963 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .B1(n9735), .B2(n9890), .ZN(ADD_1071_U46) );
  OAI21_X1 U10964 ( .B1(n9893), .B2(n9892), .A(n9891), .ZN(ADD_1071_U56) );
  OAI21_X1 U10965 ( .B1(n9896), .B2(n9895), .A(n9894), .ZN(ADD_1071_U57) );
  OAI21_X1 U10966 ( .B1(n9899), .B2(n9898), .A(n9897), .ZN(ADD_1071_U58) );
  OAI21_X1 U10967 ( .B1(n9902), .B2(n9901), .A(n9900), .ZN(ADD_1071_U59) );
  OAI21_X1 U10968 ( .B1(n9905), .B2(n9904), .A(n9903), .ZN(ADD_1071_U60) );
  OAI21_X1 U10969 ( .B1(n9908), .B2(n9907), .A(n9906), .ZN(ADD_1071_U61) );
  AOI21_X1 U10970 ( .B1(n9911), .B2(n9910), .A(n9909), .ZN(ADD_1071_U62) );
  AOI21_X1 U10971 ( .B1(n9914), .B2(n9913), .A(n9912), .ZN(ADD_1071_U63) );
  AOI22_X1 U10972 ( .A1(n7403), .A2(keyinput43), .B1(n10030), .B2(keyinput44), 
        .ZN(n9915) );
  OAI221_X1 U10973 ( .B1(n7403), .B2(keyinput43), .C1(n10030), .C2(keyinput44), 
        .A(n9915), .ZN(n9926) );
  AOI22_X1 U10974 ( .A1(n9918), .A2(keyinput10), .B1(keyinput49), .B2(n9917), 
        .ZN(n9916) );
  OAI221_X1 U10975 ( .B1(n9918), .B2(keyinput10), .C1(n9917), .C2(keyinput49), 
        .A(n9916), .ZN(n9925) );
  AOI22_X1 U10976 ( .A1(n10037), .A2(keyinput23), .B1(keyinput14), .B2(n9920), 
        .ZN(n9919) );
  OAI221_X1 U10977 ( .B1(n10037), .B2(keyinput23), .C1(n9920), .C2(keyinput14), 
        .A(n9919), .ZN(n9924) );
  XOR2_X1 U10978 ( .A(n5701), .B(keyinput32), .Z(n9922) );
  XNOR2_X1 U10979 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput20), .ZN(n9921) );
  NAND2_X1 U10980 ( .A1(n9922), .A2(n9921), .ZN(n9923) );
  NOR4_X1 U10981 ( .A1(n9926), .A2(n9925), .A3(n9924), .A4(n9923), .ZN(n9968)
         );
  INV_X1 U10982 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n9928) );
  AOI22_X1 U10983 ( .A1(n9928), .A2(keyinput63), .B1(n10040), .B2(keyinput6), 
        .ZN(n9927) );
  OAI221_X1 U10984 ( .B1(n9928), .B2(keyinput63), .C1(n10040), .C2(keyinput6), 
        .A(n9927), .ZN(n9938) );
  AOI22_X1 U10985 ( .A1(n9930), .A2(keyinput9), .B1(keyinput19), .B2(n10029), 
        .ZN(n9929) );
  OAI221_X1 U10986 ( .B1(n9930), .B2(keyinput9), .C1(n10029), .C2(keyinput19), 
        .A(n9929), .ZN(n9937) );
  AOI22_X1 U10987 ( .A1(n4425), .A2(keyinput35), .B1(keyinput51), .B2(n9932), 
        .ZN(n9931) );
  OAI221_X1 U10988 ( .B1(n4425), .B2(keyinput35), .C1(n9932), .C2(keyinput51), 
        .A(n9931), .ZN(n9936) );
  AOI22_X1 U10989 ( .A1(n8514), .A2(keyinput42), .B1(keyinput56), .B2(n9934), 
        .ZN(n9933) );
  OAI221_X1 U10990 ( .B1(n8514), .B2(keyinput42), .C1(n9934), .C2(keyinput56), 
        .A(n9933), .ZN(n9935) );
  NOR4_X1 U10991 ( .A1(n9938), .A2(n9937), .A3(n9936), .A4(n9935), .ZN(n9967)
         );
  AOI22_X1 U10992 ( .A1(n4971), .A2(keyinput8), .B1(keyinput25), .B2(n9940), 
        .ZN(n9939) );
  OAI221_X1 U10993 ( .B1(n4971), .B2(keyinput8), .C1(n9940), .C2(keyinput25), 
        .A(n9939), .ZN(n9950) );
  AOI22_X1 U10994 ( .A1(n6461), .A2(keyinput50), .B1(n9942), .B2(keyinput29), 
        .ZN(n9941) );
  OAI221_X1 U10995 ( .B1(n6461), .B2(keyinput50), .C1(n9942), .C2(keyinput29), 
        .A(n9941), .ZN(n9949) );
  AOI22_X1 U10996 ( .A1(n5778), .A2(keyinput13), .B1(n9944), .B2(keyinput45), 
        .ZN(n9943) );
  OAI221_X1 U10997 ( .B1(n5778), .B2(keyinput13), .C1(n9944), .C2(keyinput45), 
        .A(n9943), .ZN(n9948) );
  XNOR2_X1 U10998 ( .A(P2_REG1_REG_27__SCAN_IN), .B(keyinput62), .ZN(n9946) );
  XNOR2_X1 U10999 ( .A(P2_IR_REG_14__SCAN_IN), .B(keyinput0), .ZN(n9945) );
  NAND2_X1 U11000 ( .A1(n9946), .A2(n9945), .ZN(n9947) );
  NOR4_X1 U11001 ( .A1(n9950), .A2(n9949), .A3(n9948), .A4(n9947), .ZN(n9966)
         );
  INV_X1 U11002 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9953) );
  AOI22_X1 U11003 ( .A1(n9953), .A2(keyinput11), .B1(n9952), .B2(keyinput61), 
        .ZN(n9951) );
  OAI221_X1 U11004 ( .B1(n9953), .B2(keyinput11), .C1(n9952), .C2(keyinput61), 
        .A(n9951), .ZN(n9964) );
  INV_X1 U11005 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n9956) );
  AOI22_X1 U11006 ( .A1(n9956), .A2(keyinput53), .B1(n9955), .B2(keyinput40), 
        .ZN(n9954) );
  OAI221_X1 U11007 ( .B1(n9956), .B2(keyinput53), .C1(n9955), .C2(keyinput40), 
        .A(n9954), .ZN(n9963) );
  XOR2_X1 U11008 ( .A(n5564), .B(keyinput38), .Z(n9959) );
  XNOR2_X1 U11009 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(keyinput2), .ZN(n9958) );
  XNOR2_X1 U11010 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput16), .ZN(n9957) );
  NAND3_X1 U11011 ( .A1(n9959), .A2(n9958), .A3(n9957), .ZN(n9962) );
  XNOR2_X1 U11012 ( .A(n9960), .B(keyinput48), .ZN(n9961) );
  NOR4_X1 U11013 ( .A1(n9964), .A2(n9963), .A3(n9962), .A4(n9961), .ZN(n9965)
         );
  NAND4_X1 U11014 ( .A1(n9968), .A2(n9967), .A3(n9966), .A4(n9965), .ZN(n10020) );
  AOI22_X1 U11015 ( .A1(n9970), .A2(keyinput21), .B1(keyinput34), .B2(n4815), 
        .ZN(n9969) );
  OAI221_X1 U11016 ( .B1(n9970), .B2(keyinput21), .C1(n4815), .C2(keyinput34), 
        .A(n9969), .ZN(n9980) );
  AOI22_X1 U11017 ( .A1(n10028), .A2(keyinput60), .B1(n9972), .B2(keyinput15), 
        .ZN(n9971) );
  OAI221_X1 U11018 ( .B1(n10028), .B2(keyinput60), .C1(n9972), .C2(keyinput15), 
        .A(n9971), .ZN(n9979) );
  AOI22_X1 U11019 ( .A1(n10045), .A2(keyinput36), .B1(n9974), .B2(keyinput55), 
        .ZN(n9973) );
  OAI221_X1 U11020 ( .B1(n10045), .B2(keyinput36), .C1(n9974), .C2(keyinput55), 
        .A(n9973), .ZN(n9978) );
  XNOR2_X1 U11021 ( .A(P1_ADDR_REG_19__SCAN_IN), .B(keyinput24), .ZN(n9976) );
  XNOR2_X1 U11022 ( .A(P1_REG0_REG_18__SCAN_IN), .B(keyinput39), .ZN(n9975) );
  NAND2_X1 U11023 ( .A1(n9976), .A2(n9975), .ZN(n9977) );
  NOR4_X1 U11024 ( .A1(n9980), .A2(n9979), .A3(n9978), .A4(n9977), .ZN(n10018)
         );
  AOI22_X1 U11025 ( .A1(n5593), .A2(keyinput47), .B1(keyinput17), .B2(n9982), 
        .ZN(n9981) );
  OAI221_X1 U11026 ( .B1(n5593), .B2(keyinput47), .C1(n9982), .C2(keyinput17), 
        .A(n9981), .ZN(n9991) );
  INV_X1 U11027 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n9984) );
  AOI22_X1 U11028 ( .A1(n6352), .A2(keyinput22), .B1(keyinput41), .B2(n9984), 
        .ZN(n9983) );
  OAI221_X1 U11029 ( .B1(n6352), .B2(keyinput22), .C1(n9984), .C2(keyinput41), 
        .A(n9983), .ZN(n9990) );
  XNOR2_X1 U11030 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput3), .ZN(n9988) );
  XNOR2_X1 U11031 ( .A(P1_REG0_REG_19__SCAN_IN), .B(keyinput37), .ZN(n9987) );
  XNOR2_X1 U11032 ( .A(P2_IR_REG_11__SCAN_IN), .B(keyinput57), .ZN(n9986) );
  XNOR2_X1 U11033 ( .A(P1_REG3_REG_27__SCAN_IN), .B(keyinput18), .ZN(n9985) );
  NAND4_X1 U11034 ( .A1(n9988), .A2(n9987), .A3(n9986), .A4(n9985), .ZN(n9989)
         );
  NOR3_X1 U11035 ( .A1(n9991), .A2(n9990), .A3(n9989), .ZN(n10017) );
  AOI22_X1 U11036 ( .A1(n9993), .A2(keyinput31), .B1(keyinput12), .B2(n6408), 
        .ZN(n9992) );
  OAI221_X1 U11037 ( .B1(n9993), .B2(keyinput31), .C1(n6408), .C2(keyinput12), 
        .A(n9992), .ZN(n10003) );
  AOI22_X1 U11038 ( .A1(n9995), .A2(keyinput58), .B1(keyinput26), .B2(n10033), 
        .ZN(n9994) );
  OAI221_X1 U11039 ( .B1(n9995), .B2(keyinput58), .C1(n10033), .C2(keyinput26), 
        .A(n9994), .ZN(n10002) );
  AOI22_X1 U11040 ( .A1(n10044), .A2(keyinput54), .B1(keyinput4), .B2(n9997), 
        .ZN(n9996) );
  OAI221_X1 U11041 ( .B1(n10044), .B2(keyinput54), .C1(n9997), .C2(keyinput4), 
        .A(n9996), .ZN(n10001) );
  XNOR2_X1 U11042 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput59), .ZN(n9999) );
  XNOR2_X1 U11043 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput46), .ZN(n9998) );
  NAND2_X1 U11044 ( .A1(n9999), .A2(n9998), .ZN(n10000) );
  NOR4_X1 U11045 ( .A1(n10003), .A2(n10002), .A3(n10001), .A4(n10000), .ZN(
        n10016) );
  INV_X1 U11046 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n10005) );
  AOI22_X1 U11047 ( .A1(n5311), .A2(keyinput5), .B1(keyinput52), .B2(n10005), 
        .ZN(n10004) );
  OAI221_X1 U11048 ( .B1(n5311), .B2(keyinput5), .C1(n10005), .C2(keyinput52), 
        .A(n10004), .ZN(n10014) );
  INV_X1 U11049 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10027) );
  AOI22_X1 U11050 ( .A1(n10046), .A2(keyinput30), .B1(keyinput7), .B2(n10027), 
        .ZN(n10006) );
  OAI221_X1 U11051 ( .B1(n10046), .B2(keyinput30), .C1(n10027), .C2(keyinput7), 
        .A(n10006), .ZN(n10013) );
  AOI22_X1 U11052 ( .A1(n4941), .A2(keyinput28), .B1(n10008), .B2(keyinput27), 
        .ZN(n10007) );
  OAI221_X1 U11053 ( .B1(n4941), .B2(keyinput28), .C1(n10008), .C2(keyinput27), 
        .A(n10007), .ZN(n10012) );
  XOR2_X1 U11054 ( .A(n5867), .B(keyinput1), .Z(n10010) );
  XNOR2_X1 U11055 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput33), .ZN(n10009) );
  NAND2_X1 U11056 ( .A1(n10010), .A2(n10009), .ZN(n10011) );
  NOR4_X1 U11057 ( .A1(n10014), .A2(n10013), .A3(n10012), .A4(n10011), .ZN(
        n10015) );
  NAND4_X1 U11058 ( .A1(n10018), .A2(n10017), .A3(n10016), .A4(n10015), .ZN(
        n10019) );
  NOR2_X1 U11059 ( .A1(n10020), .A2(n10019), .ZN(n10023) );
  NAND2_X1 U11060 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10021), .ZN(n10022) );
  XNOR2_X1 U11061 ( .A(n10023), .B(n10022), .ZN(n10060) );
  NOR3_X1 U11062 ( .A1(P1_ADDR_REG_19__SCAN_IN), .A2(P1_REG2_REG_27__SCAN_IN), 
        .A3(P2_REG2_REG_26__SCAN_IN), .ZN(n10058) );
  NAND4_X1 U11063 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_REG0_REG_19__SCAN_IN), 
        .A3(P1_REG0_REG_18__SCAN_IN), .A4(P1_REG2_REG_17__SCAN_IN), .ZN(n10026) );
  NAND4_X1 U11064 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(P2_REG3_REG_15__SCAN_IN), 
        .A3(P2_REG2_REG_24__SCAN_IN), .A4(P2_REG2_REG_31__SCAN_IN), .ZN(n10025) );
  NAND4_X1 U11065 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(SI_22_), .A3(
        P2_DATAO_REG_19__SCAN_IN), .A4(SI_12_), .ZN(n10024) );
  NOR3_X1 U11066 ( .A1(n10026), .A2(n10025), .A3(n10024), .ZN(n10057) );
  NAND4_X1 U11067 ( .A1(P1_ADDR_REG_14__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .A3(n10028), .A4(n10027), .ZN(n10055) );
  NOR4_X1 U11068 ( .A1(n10030), .A2(n10029), .A3(n6408), .A4(n4941), .ZN(
        n10036) );
  NAND3_X1 U11069 ( .A1(n10031), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P2_IR_REG_14__SCAN_IN), .ZN(n10032) );
  NOR4_X1 U11070 ( .A1(n10033), .A2(n10032), .A3(P1_IR_REG_30__SCAN_IN), .A4(
        P2_IR_REG_3__SCAN_IN), .ZN(n10034) );
  NAND3_X1 U11071 ( .A1(n10036), .A2(n10035), .A3(n10034), .ZN(n10054) );
  NOR4_X1 U11072 ( .A1(P2_REG0_REG_13__SCAN_IN), .A2(P2_REG0_REG_10__SCAN_IN), 
        .A3(P2_REG0_REG_4__SCAN_IN), .A4(P2_REG0_REG_0__SCAN_IN), .ZN(n10043)
         );
  NOR4_X1 U11073 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(P2_DATAO_REG_1__SCAN_IN), 
        .A3(P2_REG0_REG_19__SCAN_IN), .A4(P2_REG0_REG_29__SCAN_IN), .ZN(n10042) );
  NOR4_X1 U11074 ( .A1(n10040), .A2(n10039), .A3(n10038), .A4(n10037), .ZN(
        n10041) );
  AND4_X1 U11075 ( .A1(n10044), .A2(n10043), .A3(n10042), .A4(n10041), .ZN(
        n10047) );
  NAND4_X1 U11076 ( .A1(n10047), .A2(P2_DATAO_REG_4__SCAN_IN), .A3(n10046), 
        .A4(n10045), .ZN(n10053) );
  NOR4_X1 U11077 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_REG0_REG_28__SCAN_IN), 
        .A3(P2_REG1_REG_8__SCAN_IN), .A4(P1_REG1_REG_31__SCAN_IN), .ZN(n10051)
         );
  NOR4_X1 U11078 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_REG0_REG_6__SCAN_IN), .A4(P1_REG0_REG_4__SCAN_IN), .ZN(n10050) );
  NOR4_X1 U11079 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P2_DATAO_REG_22__SCAN_IN), 
        .A3(P1_REG2_REG_6__SCAN_IN), .A4(P1_DATAO_REG_30__SCAN_IN), .ZN(n10049) );
  NOR4_X1 U11080 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG2_REG_19__SCAN_IN), 
        .A3(P1_REG0_REG_13__SCAN_IN), .A4(P2_REG1_REG_18__SCAN_IN), .ZN(n10048) );
  NAND4_X1 U11081 ( .A1(n10051), .A2(n10050), .A3(n10049), .A4(n10048), .ZN(
        n10052) );
  NOR4_X1 U11082 ( .A1(n10055), .A2(n10054), .A3(n10053), .A4(n10052), .ZN(
        n10056) );
  NAND4_X1 U11083 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(n10058), .A3(n10057), .A4(
        n10056), .ZN(n10059) );
  XNOR2_X1 U11084 ( .A(n10060), .B(n10059), .ZN(P2_U3310) );
  XOR2_X1 U11085 ( .A(n10061), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11086 ( .A(n10062), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  XOR2_X1 U11087 ( .A(n10063), .B(P2_ADDR_REG_8__SCAN_IN), .Z(ADD_1071_U48) );
  NOR2_X1 U11088 ( .A1(n10065), .A2(n10064), .ZN(n10067) );
  XNOR2_X1 U11089 ( .A(n10067), .B(n10066), .ZN(ADD_1071_U51) );
  OAI21_X1 U11090 ( .B1(n10070), .B2(n10069), .A(n10068), .ZN(n10071) );
  XNOR2_X1 U11091 ( .A(n10071), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11092 ( .B1(n10074), .B2(n10073), .A(n10072), .ZN(ADD_1071_U47) );
  XOR2_X1 U11093 ( .A(n10076), .B(n10075), .Z(ADD_1071_U54) );
  XOR2_X1 U11094 ( .A(n10078), .B(n10077), .Z(ADD_1071_U53) );
  XNOR2_X1 U11095 ( .A(n10080), .B(n10079), .ZN(ADD_1071_U52) );
  AND2_X1 U4778 ( .A1(n5876), .A2(n5875), .ZN(n5882) );
  XNOR2_X1 U4790 ( .A(n4725), .B(P2_IR_REG_29__SCAN_IN), .ZN(n4726) );
endmodule

