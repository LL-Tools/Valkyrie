

module b21_C_AntiSAT_k_256_3 ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3, 
        keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, 
        keyinput10, keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, 
        keyinput16, keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, 
        keyinput22, keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, 
        keyinput28, keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, 
        keyinput34, keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, 
        keyinput40, keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, 
        keyinput46, keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, 
        keyinput52, keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, 
        keyinput58, keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, 
        keyinput64, keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, 
        keyinput70, keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, 
        keyinput76, keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, 
        keyinput82, keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, 
        keyinput88, keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, 
        keyinput94, keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127, keyinput128, keyinput129, 
        keyinput130, keyinput131, keyinput132, keyinput133, keyinput134, 
        keyinput135, keyinput136, keyinput137, keyinput138, keyinput139, 
        keyinput140, keyinput141, keyinput142, keyinput143, keyinput144, 
        keyinput145, keyinput146, keyinput147, keyinput148, keyinput149, 
        keyinput150, keyinput151, keyinput152, keyinput153, keyinput154, 
        keyinput155, keyinput156, keyinput157, keyinput158, keyinput159, 
        keyinput160, keyinput161, keyinput162, keyinput163, keyinput164, 
        keyinput165, keyinput166, keyinput167, keyinput168, keyinput169, 
        keyinput170, keyinput171, keyinput172, keyinput173, keyinput174, 
        keyinput175, keyinput176, keyinput177, keyinput178, keyinput179, 
        keyinput180, keyinput181, keyinput182, keyinput183, keyinput184, 
        keyinput185, keyinput186, keyinput187, keyinput188, keyinput189, 
        keyinput190, keyinput191, keyinput192, keyinput193, keyinput194, 
        keyinput195, keyinput196, keyinput197, keyinput198, keyinput199, 
        keyinput200, keyinput201, keyinput202, keyinput203, keyinput204, 
        keyinput205, keyinput206, keyinput207, keyinput208, keyinput209, 
        keyinput210, keyinput211, keyinput212, keyinput213, keyinput214, 
        keyinput215, keyinput216, keyinput217, keyinput218, keyinput219, 
        keyinput220, keyinput221, keyinput222, keyinput223, keyinput224, 
        keyinput225, keyinput226, keyinput227, keyinput228, keyinput229, 
        keyinput230, keyinput231, keyinput232, keyinput233, keyinput234, 
        keyinput235, keyinput236, keyinput237, keyinput238, keyinput239, 
        keyinput240, keyinput241, keyinput242, keyinput243, keyinput244, 
        keyinput245, keyinput246, keyinput247, keyinput248, keyinput249, 
        keyinput250, keyinput251, keyinput252, keyinput253, keyinput254, 
        keyinput255, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, 
        ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, 
        ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, 
        ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, 
        ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, 
        P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, 
        P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, 
        P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, 
        P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, 
        P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, 
        P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, 
        P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, 
        P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, 
        P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, 
        P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, 
        P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, 
        P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, 
        P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, 
        P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, 
        P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, 
        P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, 
        P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, 
        P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, 
        P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, 
        P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, 
        P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, 
        P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, 
        P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, 
        P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, 
        P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, 
        P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, 
        P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, 
        P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, 
        P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, 
        P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, 
        P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, 
        P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, 
        P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, 
        P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, 
        P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, 
        P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, 
        P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, 
        P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, 
        P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, 
        P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, 
        P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, 
        P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, 
        P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, 
        P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, 
        P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, 
        P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, 
        P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, 
        P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, 
        P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, 
        P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, 
        P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, 
        P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, 
        P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, 
        P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, 
        P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, 
        P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, 
        P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, 
        P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, 
        P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, 
        P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, 
        P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, 
        P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, 
        P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, 
        P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3152, P2_U3151, P2_U3966 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4490, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
         n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
         n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
         n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
         n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
         n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
         n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
         n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
         n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
         n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
         n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
         n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
         n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
         n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
         n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
         n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
         n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
         n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
         n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
         n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871,
         n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881,
         n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891,
         n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901,
         n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911,
         n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
         n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
         n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941,
         n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951,
         n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961,
         n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971,
         n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981,
         n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991,
         n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10523;

  CLKBUF_X3 U4995 ( .A(n6228), .Z(n6193) );
  BUF_X2 U4996 ( .A(n5981), .Z(n8017) );
  INV_X2 U4998 ( .A(n5174), .ZN(n5640) );
  NAND2_X1 U4999 ( .A1(n8353), .A2(n9377), .ZN(n5174) );
  AND4_X1 U5000 ( .A1(n4840), .A2(n5864), .A3(n5863), .A4(n5865), .ZN(n4506)
         );
  INV_X1 U5001 ( .A(n10523), .ZN(n4490) );
  INV_X2 U5002 ( .A(n4490), .ZN(P1_U3084) );
  INV_X1 U5003 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n10523) );
  NOR2_X1 U5005 ( .A1(n5861), .A2(n4838), .ZN(n4837) );
  INV_X1 U5006 ( .A(n4493), .ZN(n4496) );
  INV_X1 U5007 ( .A(n5660), .ZN(n5448) );
  INV_X1 U5008 ( .A(n5992), .ZN(n6301) );
  INV_X4 U5009 ( .A(n8314), .ZN(n8341) );
  INV_X1 U5010 ( .A(n5644), .ZN(n5606) );
  INV_X1 U5011 ( .A(n4496), .ZN(n5431) );
  AND2_X1 U5012 ( .A1(n9203), .A2(n4724), .ZN(n9137) );
  AOI21_X1 U5013 ( .B1(n6066), .B2(n5066), .A(n6065), .ZN(n6084) );
  NAND2_X1 U5014 ( .A1(n5875), .A2(n5876), .ZN(n6003) );
  NAND2_X2 U5015 ( .A1(n5104), .A2(n9377), .ZN(n5644) );
  INV_X1 U5016 ( .A(n4493), .ZN(n4495) );
  INV_X1 U5017 ( .A(n5963), .ZN(n6543) );
  NAND2_X1 U5018 ( .A1(n6084), .A2(n6085), .ZN(n7432) );
  INV_X1 U5019 ( .A(n8229), .ZN(n4695) );
  XNOR2_X1 U5020 ( .A(n5657), .B(n5656), .ZN(n9367) );
  INV_X2 U5021 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n5912) );
  INV_X1 U5022 ( .A(n5103), .ZN(n9377) );
  XNOR2_X1 U5023 ( .A(n5910), .B(n5909), .ZN(n6481) );
  OR2_X1 U5024 ( .A1(n6123), .A2(n5919), .ZN(n4492) );
  AND2_X1 U5025 ( .A1(n5104), .A2(n5103), .ZN(n4493) );
  AND2_X1 U5026 ( .A1(n4780), .A2(n4779), .ZN(n4494) );
  NAND2_X2 U5027 ( .A1(n9080), .A2(n5767), .ZN(n9063) );
  AOI21_X2 U5028 ( .B1(n7330), .B2(n7329), .A(n6586), .ZN(n7599) );
  AOI211_X1 U5029 ( .C1(n7169), .C2(n7168), .A(n10455), .B(n7322), .ZN(n7220)
         );
  AND2_X2 U5030 ( .A1(n5987), .A2(n5881), .ZN(n6196) );
  XNOR2_X2 U5031 ( .A(n5162), .B(SI_3_), .ZN(n5160) );
  NAND2_X2 U5032 ( .A1(n4586), .A2(n4585), .ZN(n5162) );
  OAI21_X2 U5033 ( .B1(n5250), .B2(n5249), .A(n5251), .ZN(n5266) );
  NAND2_X2 U5034 ( .A1(n5233), .A2(n5232), .ZN(n5250) );
  NAND3_X2 U5035 ( .A1(n5142), .A2(n5141), .A3(n4536), .ZN(n6546) );
  XNOR2_X2 U5036 ( .A(n4795), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8353) );
  OR2_X1 U5037 ( .A1(n5573), .A2(n6771), .ZN(n5132) );
  OAI21_X2 U5038 ( .B1(n10165), .B2(n7490), .A(n8128), .ZN(n7723) );
  NAND2_X2 U5039 ( .A1(n7489), .A2(n8184), .ZN(n10165) );
  XNOR2_X2 U5040 ( .A(n5221), .B(SI_6_), .ZN(n5218) );
  XNOR2_X2 U5041 ( .A(n5097), .B(P2_IR_REG_21__SCAN_IN), .ZN(n6616) );
  NAND2_X2 U5042 ( .A1(n6199), .A2(n6198), .ZN(n7917) );
  NAND2_X1 U5043 ( .A1(n4856), .A2(n8600), .ZN(n8475) );
  AOI21_X1 U5044 ( .B1(n9044), .B2(n10371), .A(n9043), .ZN(n9283) );
  AOI21_X1 U5045 ( .B1(n9039), .B2(n5802), .A(n5613), .ZN(n8460) );
  AND2_X1 U5046 ( .A1(n8318), .A2(n8317), .ZN(n8536) );
  NAND2_X1 U5047 ( .A1(n8312), .A2(n8311), .ZN(n8316) );
  NAND2_X1 U5048 ( .A1(n8495), .A2(n4887), .ZN(n8551) );
  NAND2_X2 U5049 ( .A1(n5760), .A2(n9109), .ZN(n9120) );
  NAND2_X1 U5050 ( .A1(n6761), .A2(n6762), .ZN(n6763) );
  AND2_X1 U5051 ( .A1(n5950), .A2(n5949), .ZN(n6761) );
  NAND2_X1 U5052 ( .A1(n7084), .A2(n7564), .ZN(n8243) );
  INV_X1 U5053 ( .A(n7564), .ZN(n10201) );
  NOR2_X1 U5054 ( .A1(n7314), .A2(n8341), .ZN(n6556) );
  NOR2_X1 U5055 ( .A1(n6677), .A2(n7383), .ZN(n7376) );
  AND2_X1 U5056 ( .A1(n5914), .A2(n6539), .ZN(n5917) );
  INV_X1 U5057 ( .A(n8627), .ZN(n8580) );
  BUF_X2 U5058 ( .A(n6003), .Z(n6526) );
  INV_X1 U5059 ( .A(n6546), .ZN(n4719) );
  CLKBUF_X2 U5060 ( .A(n5982), .Z(n8013) );
  CLKBUF_X2 U5061 ( .A(n7015), .Z(n7237) );
  NAND2_X1 U5062 ( .A1(n6780), .A2(n4583), .ZN(n5185) );
  NAND2_X2 U5063 ( .A1(n6797), .A2(n9385), .ZN(n6780) );
  INV_X1 U5064 ( .A(n6616), .ZN(n7520) );
  INV_X2 U5065 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n4694) );
  AOI21_X1 U5066 ( .B1(n4962), .B2(n4961), .A(n4523), .ZN(n4960) );
  NAND2_X1 U5067 ( .A1(n4706), .A2(n6430), .ZN(n9493) );
  AOI211_X1 U5068 ( .C1(n9275), .C2(n9262), .A(n8469), .B(n8468), .ZN(n8470)
         );
  NOR2_X1 U5069 ( .A1(n9397), .A2(n9399), .ZN(n9401) );
  NAND2_X1 U5070 ( .A1(n4708), .A2(n4707), .ZN(n4706) );
  AND2_X1 U5071 ( .A1(n4736), .A2(n9052), .ZN(n4670) );
  NOR2_X1 U5072 ( .A1(n6394), .A2(n6393), .ZN(n9396) );
  AOI21_X1 U5073 ( .B1(n8467), .B2(n10371), .A(n8466), .ZN(n9276) );
  OR2_X1 U5074 ( .A1(n6391), .A2(n6392), .ZN(n4710) );
  NAND2_X1 U5075 ( .A1(n8521), .A2(n8520), .ZN(n8602) );
  OR2_X1 U5076 ( .A1(n9266), .A2(n6669), .ZN(n5796) );
  AND2_X1 U5077 ( .A1(n9266), .A2(n6669), .ZN(n5799) );
  NAND2_X1 U5078 ( .A1(n4987), .A2(n4986), .ZN(n6371) );
  NAND2_X1 U5079 ( .A1(n8008), .A2(n5963), .ZN(n9921) );
  NAND2_X1 U5080 ( .A1(n9618), .A2(n4749), .ZN(n4820) );
  NAND2_X1 U5081 ( .A1(n5662), .A2(n5661), .ZN(n9266) );
  OAI21_X1 U5082 ( .B1(n9632), .B2(n8382), .A(n8381), .ZN(n9618) );
  NAND2_X1 U5083 ( .A1(n8379), .A2(n8378), .ZN(n9632) );
  INV_X1 U5084 ( .A(n9273), .ZN(n8683) );
  XNOR2_X1 U5085 ( .A(n5652), .B(n5651), .ZN(n5649) );
  AOI21_X1 U5086 ( .B1(n5035), .B2(n5038), .A(n5034), .ZN(n5033) );
  OR2_X1 U5087 ( .A1(n9280), .A2(n8342), .ZN(n5776) );
  AND2_X1 U5088 ( .A1(n4557), .A2(n5036), .ZN(n5035) );
  NAND2_X1 U5089 ( .A1(n5632), .A2(n5631), .ZN(n5652) );
  OR2_X1 U5090 ( .A1(n5629), .A2(n5628), .ZN(n5632) );
  NAND2_X1 U5091 ( .A1(n8494), .A2(n8293), .ZN(n8495) );
  NAND2_X1 U5092 ( .A1(n6464), .A2(n6463), .ZN(n9783) );
  NOR2_X1 U5093 ( .A1(n9120), .A2(n5040), .ZN(n5039) );
  OR2_X1 U5094 ( .A1(n6429), .A2(n6428), .ZN(n6430) );
  NAND2_X1 U5095 ( .A1(n6451), .A2(n6450), .ZN(n9789) );
  OAI21_X1 U5096 ( .B1(n9740), .B2(n4829), .A(n4827), .ZN(n8370) );
  NAND2_X1 U5097 ( .A1(n5600), .A2(n5599), .ZN(n5615) );
  INV_X1 U5098 ( .A(n9128), .ZN(n9305) );
  NAND2_X1 U5099 ( .A1(n5567), .A2(n5566), .ZN(n9291) );
  NAND2_X1 U5100 ( .A1(n5581), .A2(n5580), .ZN(n5598) );
  NAND2_X1 U5101 ( .A1(n7962), .A2(n4883), .ZN(n7976) );
  NAND2_X1 U5102 ( .A1(n5529), .A2(n5528), .ZN(n9300) );
  NAND2_X1 U5103 ( .A1(n6396), .A2(n6395), .ZN(n9633) );
  AND2_X1 U5104 ( .A1(n5516), .A2(n5515), .ZN(n9128) );
  AND2_X1 U5105 ( .A1(n5756), .A2(n5757), .ZN(n9143) );
  OR2_X1 U5106 ( .A1(n9310), .A2(n8567), .ZN(n5756) );
  NAND2_X1 U5107 ( .A1(n7952), .A2(n7951), .ZN(n7962) );
  NAND2_X1 U5108 ( .A1(n5496), .A2(n5495), .ZN(n9310) );
  NAND2_X1 U5109 ( .A1(n4582), .A2(n8136), .ZN(n8394) );
  NOR2_X1 U5110 ( .A1(n7855), .A2(n5058), .ZN(n7988) );
  AOI21_X1 U5111 ( .B1(n4830), .B2(n4828), .A(n4540), .ZN(n4827) );
  OR2_X1 U5112 ( .A1(n5508), .A2(n4956), .ZN(n4949) );
  AOI21_X1 U5113 ( .B1(n9961), .B2(n8052), .A(n7719), .ZN(n7720) );
  NAND2_X1 U5114 ( .A1(n5490), .A2(n5489), .ZN(n5508) );
  NAND2_X1 U5115 ( .A1(n7655), .A2(n7654), .ZN(n10265) );
  NAND2_X1 U5116 ( .A1(n5478), .A2(n5477), .ZN(n4966) );
  OR2_X1 U5117 ( .A1(n9346), .A2(n9243), .ZN(n5737) );
  AND2_X1 U5118 ( .A1(n4982), .A2(n4700), .ZN(n4699) );
  AND2_X1 U5119 ( .A1(n4983), .A2(n7639), .ZN(n4982) );
  NOR2_X1 U5120 ( .A1(n8134), .A2(n4745), .ZN(n4744) );
  NAND2_X1 U5121 ( .A1(n5374), .A2(n5373), .ZN(n9346) );
  NAND2_X1 U5122 ( .A1(n6287), .A2(n6286), .ZN(n9838) );
  NAND2_X1 U5123 ( .A1(n5430), .A2(n5429), .ZN(n9329) );
  NAND2_X1 U5124 ( .A1(n7601), .A2(n4886), .ZN(n7653) );
  NAND2_X1 U5125 ( .A1(n6268), .A2(n6267), .ZN(n9845) );
  NAND2_X1 U5126 ( .A1(n5396), .A2(n5395), .ZN(n9340) );
  NAND2_X1 U5127 ( .A1(n5412), .A2(n5411), .ZN(n9335) );
  AND2_X1 U5128 ( .A1(n9963), .A2(n9993), .ZN(n9936) );
  OR2_X1 U5129 ( .A1(n7917), .A2(n9504), .ZN(n8064) );
  AND2_X1 U5130 ( .A1(n5710), .A2(n5712), .ZN(n7849) );
  OAI21_X1 U5131 ( .B1(n5427), .B2(n5426), .A(n5425), .ZN(n5440) );
  NAND2_X1 U5132 ( .A1(n6161), .A2(n6160), .ZN(n7779) );
  NAND2_X1 U5133 ( .A1(n5313), .A2(n5312), .ZN(n10274) );
  NAND2_X1 U5134 ( .A1(n5293), .A2(n5292), .ZN(n7758) );
  NAND2_X1 U5135 ( .A1(n6138), .A2(n6137), .ZN(n9973) );
  NAND2_X1 U5136 ( .A1(n5332), .A2(n5331), .ZN(n7932) );
  OAI21_X1 U5137 ( .B1(n5363), .B2(n4970), .A(n4968), .ZN(n5407) );
  NAND2_X1 U5138 ( .A1(n5342), .A2(n5341), .ZN(n5363) );
  OR2_X1 U5139 ( .A1(n10160), .A2(n7716), .ZN(n9962) );
  OR2_X1 U5140 ( .A1(n7524), .A2(n8125), .ZN(n7583) );
  NAND2_X1 U5141 ( .A1(n6117), .A2(n6116), .ZN(n7716) );
  NAND2_X1 U5142 ( .A1(n5268), .A2(n5267), .ZN(n5287) );
  NAND2_X1 U5143 ( .A1(n4663), .A2(n8171), .ZN(n7484) );
  AND2_X2 U5144 ( .A1(n7478), .A2(n10178), .ZN(n9953) );
  INV_X2 U5145 ( .A(n7864), .ZN(n10372) );
  AND2_X1 U5146 ( .A1(n5192), .A2(n4642), .ZN(n7238) );
  OAI211_X1 U5147 ( .C1(n5963), .C2(n10027), .A(n5994), .B(n5993), .ZN(n7197)
         );
  NAND2_X1 U5148 ( .A1(n4617), .A2(n5190), .ZN(n5204) );
  OAI211_X1 U5149 ( .C1(n5963), .C2(n6831), .A(n5930), .B(n5929), .ZN(n7564)
         );
  OAI211_X1 U5150 ( .C1(n6780), .C2(n6639), .A(n5156), .B(n5155), .ZN(n7169)
         );
  NAND4_X1 U5151 ( .A1(n5986), .A2(n5985), .A3(n5984), .A4(n5983), .ZN(n9529)
         );
  OR2_X1 U5152 ( .A1(n6481), .A2(n4695), .ZN(n6964) );
  NAND4_X2 U5153 ( .A1(n5960), .A2(n5958), .A3(n5959), .A4(n5957), .ZN(n9531)
         );
  AND4_X1 U5154 ( .A1(n5146), .A2(n5145), .A3(n5144), .A4(n5143), .ZN(n7314)
         );
  NAND2_X1 U5155 ( .A1(n5908), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5910) );
  AND2_X1 U5156 ( .A1(n5908), .A2(n5887), .ZN(n6482) );
  OR2_X1 U5157 ( .A1(n5992), .A2(n6630), .ZN(n4843) );
  INV_X2 U5158 ( .A(n6013), .ZN(n8096) );
  OR2_X1 U5159 ( .A1(n5886), .A2(n5885), .ZN(n5887) );
  NAND2_X1 U5160 ( .A1(n8434), .A2(n5876), .ZN(n5981) );
  NAND2_X1 U5161 ( .A1(n5963), .A2(n4497), .ZN(n6013) );
  INV_X2 U5162 ( .A(n5185), .ZN(n5658) );
  XNOR2_X1 U5163 ( .A(n5081), .B(n5080), .ZN(n8355) );
  AOI21_X1 U5164 ( .B1(n5219), .B2(n4933), .A(n4547), .ZN(n4932) );
  XNOR2_X1 U5165 ( .A(n5873), .B(n4836), .ZN(n5874) );
  XNOR2_X1 U5167 ( .A(n5889), .B(n5888), .ZN(n8266) );
  NAND2_X1 U5168 ( .A1(n4715), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5889) );
  OAI21_X1 U5169 ( .B1(n4766), .B2(n6503), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5899) );
  CLKBUF_X3 U5170 ( .A(n5154), .Z(n8007) );
  NAND2_X2 U5171 ( .A1(n4583), .A2(P1_U3084), .ZN(n9891) );
  OAI21_X1 U5172 ( .B1(n5847), .B2(n4926), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n4738) );
  CLKBUF_X3 U5173 ( .A(n5154), .Z(n4497) );
  INV_X2 U5174 ( .A(n5112), .ZN(n5154) );
  NAND2_X1 U5175 ( .A1(n5002), .A2(n5001), .ZN(n5847) );
  NOR2_X2 U5176 ( .A1(n5988), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n5987) );
  INV_X1 U5177 ( .A(n4928), .ZN(n4926) );
  AND2_X1 U5178 ( .A1(n5121), .A2(n5068), .ZN(n5169) );
  OAI21_X1 U5179 ( .B1(P1_RD_REG_SCAN_IN), .B2(P2_ADDR_REG_19__SCAN_IN), .A(
        n4979), .ZN(n4978) );
  AND2_X1 U5180 ( .A1(n5912), .A2(n6282), .ZN(n4840) );
  NAND3_X1 U5181 ( .A1(n5904), .A2(n4694), .A3(n5962), .ZN(n5926) );
  INV_X4 U5182 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NOR2_X1 U5183 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5121) );
  INV_X1 U5184 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5888) );
  INV_X1 U5185 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6157) );
  INV_X1 U5186 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n6108) );
  NOR2_X1 U5187 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n5859) );
  INV_X1 U5188 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6177) );
  INV_X1 U5189 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5904) );
  INV_X1 U5190 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8924) );
  INV_X1 U5191 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5070) );
  AOI211_X2 U5192 ( .C1(n10163), .C2(n9779), .A(n8422), .B(n8421), .ZN(n8423)
         );
  NAND2_X2 U5193 ( .A1(n6482), .A2(n8266), .ZN(n5914) );
  XNOR2_X1 U5194 ( .A(n5915), .B(n5953), .ZN(n5975) );
  OAI21_X2 U5195 ( .B1(n6503), .B2(n4841), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5902) );
  NAND2_X1 U5196 ( .A1(n4980), .A2(n4978), .ZN(n5112) );
  XNOR2_X1 U5197 ( .A(n5899), .B(n5898), .ZN(n6524) );
  AOI21_X1 U5198 ( .B1(n4770), .B2(n4772), .A(n4769), .ZN(n4768) );
  NAND2_X1 U5199 ( .A1(n5750), .A2(n5749), .ZN(n4769) );
  AND2_X1 U5200 ( .A1(n4908), .A2(n7295), .ZN(n4905) );
  NOR2_X1 U5201 ( .A1(n4913), .A2(n7298), .ZN(n4908) );
  AND2_X1 U5202 ( .A1(n5099), .A2(n5095), .ZN(n5001) );
  NOR3_X1 U5203 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_24__SCAN_IN), .A3(
        P2_IR_REG_23__SCAN_IN), .ZN(n5099) );
  INV_X1 U5204 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5072) );
  NAND2_X1 U5205 ( .A1(n4947), .A2(n4948), .ZN(n5561) );
  AOI21_X1 U5206 ( .B1(n4956), .B2(n4500), .A(n4576), .ZN(n4948) );
  NAND2_X1 U5207 ( .A1(n5508), .A2(n4500), .ZN(n4947) );
  INV_X1 U5208 ( .A(n5699), .ZN(n4792) );
  OR2_X1 U5209 ( .A1(n5715), .A2(n5714), .ZN(n4616) );
  NAND2_X1 U5210 ( .A1(n5754), .A2(n5797), .ZN(n4778) );
  NAND2_X1 U5211 ( .A1(n5327), .A2(n5326), .ZN(n5341) );
  INV_X1 U5212 ( .A(n8353), .ZN(n5104) );
  NOR2_X1 U5213 ( .A1(n9321), .A2(n9326), .ZN(n4728) );
  OR2_X1 U5214 ( .A1(n5028), .A2(n5322), .ZN(n5027) );
  AND2_X1 U5215 ( .A1(n7849), .A2(n5029), .ZN(n5028) );
  AND2_X1 U5216 ( .A1(n7452), .A2(n5007), .ZN(n4503) );
  NAND2_X1 U5217 ( .A1(n5008), .A2(n5696), .ZN(n5007) );
  INV_X1 U5218 ( .A(n5009), .ZN(n5008) );
  NOR2_X1 U5219 ( .A1(n10343), .A2(n5010), .ZN(n5009) );
  INV_X1 U5220 ( .A(n5691), .ZN(n5010) );
  NAND2_X1 U5221 ( .A1(n7238), .A2(n10367), .ZN(n5812) );
  AND2_X1 U5222 ( .A1(n7637), .A2(n7520), .ZN(n7021) );
  INV_X1 U5223 ( .A(n9451), .ZN(n4985) );
  INV_X1 U5224 ( .A(n8434), .ZN(n5875) );
  NAND2_X1 U5225 ( .A1(n4799), .A2(n4521), .ZN(n4796) );
  INV_X1 U5226 ( .A(n4816), .ZN(n4815) );
  OAI21_X1 U5227 ( .B1(n8133), .B2(n4817), .A(n7782), .ZN(n4816) );
  NOR2_X1 U5228 ( .A1(n4823), .A2(n4822), .ZN(n4821) );
  NAND2_X1 U5229 ( .A1(n5619), .A2(n5618), .ZN(n5629) );
  NAND2_X1 U5230 ( .A1(n5615), .A2(n5614), .ZN(n5619) );
  NOR2_X1 U5231 ( .A1(n4994), .A2(n5870), .ZN(n4993) );
  NAND2_X1 U5232 ( .A1(n4995), .A2(n5901), .ZN(n4994) );
  OAI21_X1 U5233 ( .B1(n5561), .B2(n5560), .A(n5559), .ZN(n5579) );
  AOI21_X1 U5234 ( .B1(n5512), .B2(n4955), .A(n4954), .ZN(n4953) );
  INV_X1 U5235 ( .A(n5526), .ZN(n4954) );
  INV_X1 U5236 ( .A(n5506), .ZN(n4955) );
  INV_X1 U5237 ( .A(n5507), .ZN(n4957) );
  INV_X1 U5238 ( .A(n5366), .ZN(n4975) );
  AOI21_X1 U5239 ( .B1(n4502), .B2(n4946), .A(n4937), .ZN(n4936) );
  INV_X1 U5240 ( .A(n5323), .ZN(n4937) );
  AND2_X1 U5241 ( .A1(n9280), .A2(n4871), .ZN(n4870) );
  OAI21_X1 U5242 ( .B1(n4494), .B2(n5800), .A(n8355), .ZN(n5833) );
  INV_X2 U5243 ( .A(n5157), .ZN(n5573) );
  INV_X1 U5244 ( .A(n5274), .ZN(n5074) );
  OAI21_X1 U5245 ( .B1(n9283), .B2(n10372), .A(n9051), .ZN(n4737) );
  NAND2_X1 U5246 ( .A1(n4687), .A2(n4515), .ZN(n4686) );
  INV_X1 U5247 ( .A(n4690), .ZN(n4687) );
  AOI21_X1 U5248 ( .B1(n4692), .B2(n4691), .A(n4543), .ZN(n4690) );
  OR2_X1 U5249 ( .A1(n10274), .A2(n8619), .ZN(n4923) );
  NOR2_X1 U5250 ( .A1(n7849), .A2(n4922), .ZN(n4921) );
  INV_X1 U5251 ( .A(n7740), .ZN(n4922) );
  NAND2_X1 U5252 ( .A1(n10345), .A2(n4532), .ZN(n7503) );
  OAI21_X1 U5253 ( .B1(n7311), .B2(n5012), .A(n5011), .ZN(n10364) );
  INV_X1 U5254 ( .A(n5017), .ZN(n5012) );
  AOI21_X1 U5255 ( .B1(n5017), .B2(n5016), .A(n5015), .ZN(n5011) );
  INV_X1 U5256 ( .A(n5019), .ZN(n5016) );
  AND2_X1 U5257 ( .A1(n6797), .A2(n6623), .ZN(n10368) );
  XNOR2_X1 U5258 ( .A(n5102), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5103) );
  NAND2_X1 U5259 ( .A1(n5101), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5102) );
  INV_X1 U5260 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n5069) );
  NOR2_X1 U5261 ( .A1(P2_IR_REG_4__SCAN_IN), .A2(P2_IR_REG_8__SCAN_IN), .ZN(
        n5071) );
  INV_X1 U5262 ( .A(n6481), .ZN(n8273) );
  OAI21_X1 U5263 ( .B1(n4668), .B2(n4666), .A(n4664), .ZN(n8233) );
  NOR2_X1 U5264 ( .A1(n8106), .A2(n8107), .ZN(n4668) );
  AOI21_X1 U5265 ( .B1(n8146), .B2(n8090), .A(n4665), .ZN(n4664) );
  OAI21_X1 U5266 ( .B1(n8105), .B2(n8090), .A(n4667), .ZN(n4666) );
  INV_X1 U5267 ( .A(n8013), .ZN(n6433) );
  NAND2_X1 U5268 ( .A1(n5875), .A2(n5874), .ZN(n5982) );
  NOR2_X1 U5269 ( .A1(n10106), .A2(n7901), .ZN(n10105) );
  NAND2_X1 U5270 ( .A1(n9600), .A2(n8414), .ZN(n9574) );
  NOR2_X1 U5271 ( .A1(n9570), .A2(n4810), .ZN(n4809) );
  INV_X1 U5272 ( .A(n8387), .ZN(n4810) );
  NAND2_X1 U5273 ( .A1(n8376), .A2(n4517), .ZN(n4825) );
  AND2_X1 U5274 ( .A1(n6972), .A2(n6971), .ZN(n9945) );
  NAND2_X1 U5275 ( .A1(n6970), .A2(n6969), .ZN(n10172) );
  NAND2_X1 U5276 ( .A1(n6972), .A2(n4498), .ZN(n10167) );
  INV_X1 U5277 ( .A(n8392), .ZN(n9778) );
  INV_X1 U5278 ( .A(n9782), .ZN(n4762) );
  OR2_X1 U5279 ( .A1(n8107), .A2(n6968), .ZN(n9862) );
  NAND2_X1 U5280 ( .A1(n6488), .A2(n5896), .ZN(n6539) );
  CLKBUF_X1 U5281 ( .A(n6482), .Z(n6483) );
  BUF_X1 U5282 ( .A(n5112), .Z(n4583) );
  AND2_X1 U5283 ( .A1(n8268), .A2(n4965), .ZN(n4964) );
  INV_X1 U5284 ( .A(n8276), .ZN(n4965) );
  NAND2_X1 U5285 ( .A1(n8267), .A2(n8266), .ZN(n8268) );
  INV_X1 U5286 ( .A(n5706), .ZN(n4790) );
  NAND2_X1 U5287 ( .A1(n4615), .A2(n4614), .ZN(n4794) );
  OR2_X1 U5288 ( .A1(n5716), .A2(n5797), .ZN(n4793) );
  OAI21_X1 U5289 ( .B1(n4616), .B2(n7873), .A(n10274), .ZN(n4615) );
  INV_X1 U5290 ( .A(n5759), .ZN(n4777) );
  NAND2_X1 U5291 ( .A1(n4626), .A2(n4623), .ZN(n4622) );
  INV_X1 U5292 ( .A(n4625), .ZN(n4623) );
  AOI21_X1 U5293 ( .B1(n4550), .B2(n5774), .A(n9064), .ZN(n4625) );
  INV_X1 U5294 ( .A(n8204), .ZN(n4660) );
  OR2_X1 U5295 ( .A1(n8092), .A2(n8207), .ZN(n4658) );
  NOR2_X1 U5296 ( .A1(n5646), .A2(n5791), .ZN(n4781) );
  OR2_X1 U5297 ( .A1(n9296), .A2(n8604), .ZN(n5558) );
  NOR2_X1 U5298 ( .A1(n4913), .A2(n4912), .ZN(n4911) );
  INV_X1 U5299 ( .A(n4917), .ZN(n4912) );
  OR2_X1 U5300 ( .A1(n4646), .A2(n4650), .ZN(n4645) );
  NAND2_X1 U5301 ( .A1(n8415), .A2(n4647), .ZN(n4646) );
  NOR2_X1 U5302 ( .A1(n8218), .A2(n8210), .ZN(n4647) );
  NAND2_X1 U5303 ( .A1(n8149), .A2(n8415), .ZN(n4648) );
  AND2_X1 U5304 ( .A1(n4654), .A2(n4653), .ZN(n4652) );
  NAND2_X1 U5305 ( .A1(n8211), .A2(n8090), .ZN(n4653) );
  OAI21_X1 U5306 ( .B1(n8094), .B2(n8093), .A(n9605), .ZN(n8095) );
  NOR2_X1 U5307 ( .A1(n4661), .A2(n4656), .ZN(n8093) );
  INV_X1 U5308 ( .A(n5404), .ZN(n4969) );
  INV_X1 U5309 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n5269) );
  OR2_X1 U5310 ( .A1(n6048), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n6110) );
  NOR2_X1 U5311 ( .A1(n5218), .A2(n5202), .ZN(n4931) );
  NAND2_X1 U5312 ( .A1(n4859), .A2(n6555), .ZN(n4860) );
  INV_X1 U5313 ( .A(n10248), .ZN(n4859) );
  NAND2_X1 U5314 ( .A1(n8627), .A2(n8314), .ZN(n6549) );
  OR2_X1 U5315 ( .A1(n8683), .A2(n5663), .ZN(n5827) );
  OR2_X1 U5316 ( .A1(n9291), .A2(n8522), .ZN(n5769) );
  NAND2_X1 U5317 ( .A1(n5039), .A2(n5037), .ZN(n5036) );
  INV_X1 U5318 ( .A(n5505), .ZN(n5037) );
  INV_X1 U5319 ( .A(n5039), .ZN(n5038) );
  AND2_X1 U5320 ( .A1(n5558), .A2(n5768), .ZN(n8448) );
  OR2_X1 U5321 ( .A1(n9300), .A2(n8540), .ZN(n5762) );
  NOR2_X1 U5322 ( .A1(n4727), .A2(n9315), .ZN(n4726) );
  INV_X1 U5323 ( .A(n4728), .ZN(n4727) );
  NAND2_X1 U5324 ( .A1(n8443), .A2(n4925), .ZN(n4924) );
  INV_X1 U5325 ( .A(n8442), .ZN(n4925) );
  NAND2_X1 U5326 ( .A1(n5045), .A2(n5041), .ZN(n9184) );
  OAI21_X1 U5327 ( .B1(n5044), .B2(n5043), .A(n5746), .ZN(n5042) );
  NOR2_X1 U5328 ( .A1(n9245), .A2(n5051), .ZN(n5050) );
  NAND2_X1 U5329 ( .A1(n7995), .A2(n5737), .ZN(n5051) );
  AND2_X1 U5330 ( .A1(n5736), .A2(n5733), .ZN(n5803) );
  AOI21_X1 U5331 ( .B1(n5027), .B2(n5025), .A(n5024), .ZN(n5023) );
  INV_X1 U5332 ( .A(n5027), .ZN(n5026) );
  INV_X1 U5333 ( .A(n4516), .ZN(n5025) );
  INV_X1 U5334 ( .A(n4734), .ZN(n4733) );
  OR2_X1 U5335 ( .A1(n10445), .A2(n10436), .ZN(n4734) );
  NAND2_X1 U5336 ( .A1(n4786), .A2(n4785), .ZN(n5815) );
  NAND2_X1 U5337 ( .A1(n8627), .A2(n4719), .ZN(n5809) );
  NOR2_X1 U5338 ( .A1(n10377), .A2(n7458), .ZN(n10358) );
  INV_X1 U5339 ( .A(n5815), .ZN(n5667) );
  NAND2_X1 U5340 ( .A1(n8424), .A2(n8431), .ZN(n7025) );
  INV_X1 U5341 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5347) );
  NAND2_X1 U5342 ( .A1(n5079), .A2(n4882), .ZN(n4881) );
  NAND2_X1 U5343 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), 
        .ZN(n4882) );
  AOI21_X1 U5344 ( .B1(n4988), .B2(n4991), .A(n4509), .ZN(n4986) );
  NAND2_X1 U5345 ( .A1(n4713), .A2(n4711), .ZN(n4987) );
  NAND2_X1 U5346 ( .A1(n6964), .A2(n5914), .ZN(n5953) );
  NAND2_X1 U5347 ( .A1(n4718), .A2(n4534), .ZN(n6255) );
  OR2_X1 U5348 ( .A1(n10092), .A2(n4588), .ZN(n4587) );
  AND2_X1 U5349 ( .A1(n10097), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4588) );
  OR2_X1 U5350 ( .A1(n9823), .A2(n8025), .ZN(n8178) );
  AND2_X1 U5351 ( .A1(n4854), .A2(n4853), .ZN(n4852) );
  NOR2_X1 U5352 ( .A1(n9838), .A2(n9845), .ZN(n4854) );
  OR2_X1 U5353 ( .A1(n7716), .A2(n10168), .ZN(n8152) );
  OR2_X1 U5354 ( .A1(n4849), .A2(n7595), .ZN(n4848) );
  OR2_X1 U5355 ( .A1(n7532), .A2(n7466), .ZN(n4849) );
  NAND2_X1 U5356 ( .A1(n6880), .A2(n6879), .ZN(n7357) );
  AND2_X1 U5357 ( .A1(n5580), .A2(n5565), .ZN(n5578) );
  NAND2_X1 U5358 ( .A1(n5443), .A2(n5442), .ZN(n5464) );
  NOR2_X1 U5359 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_14__SCAN_IN), .ZN(
        n5882) );
  AOI21_X1 U5360 ( .B1(n5362), .B2(n4974), .A(n4972), .ZN(n4971) );
  INV_X1 U5361 ( .A(n5385), .ZN(n4972) );
  AOI21_X1 U5362 ( .B1(n4944), .B2(n5301), .A(n4548), .ZN(n4943) );
  NOR2_X1 U5363 ( .A1(n5062), .A2(n4945), .ZN(n4944) );
  INV_X1 U5364 ( .A(n5287), .ZN(n4941) );
  OR2_X1 U5365 ( .A1(n5174), .A2(n5127), .ZN(n5128) );
  NAND2_X1 U5366 ( .A1(n7824), .A2(n7823), .ZN(n7952) );
  AOI21_X1 U5367 ( .B1(n4877), .B2(n4875), .A(n4874), .ZN(n4873) );
  INV_X1 U5368 ( .A(n4877), .ZN(n4876) );
  AND4_X1 U5369 ( .A1(n5265), .A2(n5264), .A3(n5263), .A4(n5262), .ZN(n7501)
         );
  AND4_X1 U5370 ( .A1(n5217), .A2(n5216), .A3(n5215), .A4(n5214), .ZN(n7444)
         );
  NOR2_X1 U5371 ( .A1(n5573), .A2(n6777), .ZN(n4788) );
  NAND2_X1 U5372 ( .A1(n10320), .A2(n4567), .ZN(n8632) );
  NAND2_X1 U5373 ( .A1(n8632), .A2(n8631), .ZN(n8630) );
  AND2_X1 U5374 ( .A1(n5074), .A2(n4525), .ZN(n5330) );
  NOR2_X1 U5375 ( .A1(n7626), .A2(n7627), .ZN(n7628) );
  NAND2_X1 U5376 ( .A1(n7628), .A2(n7629), .ZN(n7663) );
  NAND2_X1 U5377 ( .A1(n5622), .A2(n5621), .ZN(n9274) );
  OR2_X1 U5378 ( .A1(n9285), .A2(n9083), .ZN(n8452) );
  NAND2_X1 U5379 ( .A1(n9088), .A2(n8450), .ZN(n9073) );
  NAND2_X1 U5380 ( .A1(n4904), .A2(n5064), .ZN(n4903) );
  INV_X1 U5381 ( .A(n9112), .ZN(n4904) );
  INV_X1 U5382 ( .A(n4900), .ZN(n4899) );
  OAI21_X1 U5383 ( .B1(n4901), .B2(n9112), .A(n8447), .ZN(n4900) );
  OR2_X1 U5384 ( .A1(n9300), .A2(n9131), .ZN(n8447) );
  OR2_X1 U5385 ( .A1(n9120), .A2(n4902), .ZN(n4901) );
  INV_X1 U5386 ( .A(n8448), .ZN(n9098) );
  AOI21_X1 U5387 ( .B1(n9136), .B2(n8446), .A(n8445), .ZN(n9121) );
  NAND2_X1 U5388 ( .A1(n9121), .A2(n9120), .ZN(n9119) );
  NAND2_X1 U5389 ( .A1(n4682), .A2(n4681), .ZN(n9152) );
  AOI21_X1 U5390 ( .B1(n4683), .B2(n4688), .A(n4545), .ZN(n4681) );
  NAND2_X1 U5391 ( .A1(n9203), .A2(n4728), .ZN(n9166) );
  AND2_X1 U5392 ( .A1(n5751), .A2(n5750), .ZN(n9174) );
  NAND2_X1 U5393 ( .A1(n4692), .A2(n4515), .ZN(n4688) );
  AND2_X1 U5394 ( .A1(n5747), .A2(n5749), .ZN(n9185) );
  AND2_X1 U5395 ( .A1(n4554), .A2(n9245), .ZN(n4693) );
  AOI21_X1 U5396 ( .B1(n5049), .B2(n5047), .A(n5731), .ZN(n5046) );
  INV_X1 U5397 ( .A(n5052), .ZN(n5047) );
  INV_X1 U5398 ( .A(n5049), .ZN(n5048) );
  NAND2_X1 U5399 ( .A1(n7859), .A2(n4720), .ZN(n9228) );
  AND2_X1 U5400 ( .A1(n4504), .A2(n4721), .ZN(n4720) );
  NOR2_X1 U5401 ( .A1(n9228), .A2(n9329), .ZN(n9203) );
  NAND2_X1 U5402 ( .A1(n9236), .A2(n4518), .ZN(n9221) );
  INV_X1 U5403 ( .A(n5803), .ZN(n9222) );
  NAND2_X1 U5404 ( .A1(n8439), .A2(n9245), .ZN(n9236) );
  AND4_X1 U5405 ( .A1(n5420), .A2(n5419), .A3(n5418), .A4(n5417), .ZN(n9241)
         );
  NAND2_X1 U5406 ( .A1(n4920), .A2(n4535), .ZN(n7869) );
  OR2_X1 U5407 ( .A1(n5333), .A2(n7827), .ZN(n5354) );
  NOR2_X1 U5408 ( .A1(n7878), .A2(n7932), .ZN(n7859) );
  NAND2_X1 U5409 ( .A1(n4674), .A2(n4672), .ZN(n7741) );
  INV_X1 U5410 ( .A(n4673), .ZN(n4672) );
  NAND2_X1 U5411 ( .A1(n7505), .A2(n7737), .ZN(n4674) );
  OAI21_X1 U5412 ( .B1(n5819), .B2(n4675), .A(n7739), .ZN(n4673) );
  AND2_X1 U5413 ( .A1(n5706), .A2(n5705), .ZN(n7504) );
  AND2_X1 U5414 ( .A1(n5700), .A2(n5701), .ZN(n7452) );
  AND2_X1 U5415 ( .A1(n4906), .A2(n10343), .ZN(n4669) );
  OR2_X1 U5416 ( .A1(n7299), .A2(n5688), .ZN(n5227) );
  AND4_X1 U5417 ( .A1(n5248), .A2(n5247), .A3(n5246), .A4(n5245), .ZN(n7453)
         );
  AND2_X1 U5418 ( .A1(n4919), .A2(n7296), .ZN(n4917) );
  NOR2_X1 U5419 ( .A1(n7302), .A2(n8623), .ZN(n4916) );
  INV_X1 U5420 ( .A(n5812), .ZN(n5668) );
  AND2_X1 U5421 ( .A1(n5013), .A2(n5813), .ZN(n5017) );
  NAND2_X1 U5422 ( .A1(n5019), .A2(n5667), .ZN(n5013) );
  NAND2_X1 U5423 ( .A1(n7318), .A2(n7232), .ZN(n7297) );
  AND4_X1 U5424 ( .A1(n5183), .A2(n5182), .A3(n5181), .A4(n5180), .ZN(n7313)
         );
  NAND2_X1 U5425 ( .A1(n8465), .A2(n8464), .ZN(n8466) );
  NAND2_X1 U5426 ( .A1(n5470), .A2(n5469), .ZN(n9321) );
  AND2_X1 U5427 ( .A1(n8355), .A2(n7021), .ZN(n10447) );
  INV_X1 U5428 ( .A(n10447), .ZN(n10455) );
  OR2_X1 U5429 ( .A1(n10428), .A2(n6616), .ZN(n7213) );
  AND2_X1 U5430 ( .A1(n6601), .A2(n6607), .ZN(n10384) );
  NOR2_X1 U5431 ( .A1(n5031), .A2(P2_IR_REG_26__SCAN_IN), .ZN(n5030) );
  NAND2_X1 U5432 ( .A1(n5111), .A2(n5109), .ZN(n5031) );
  OAI21_X1 U5433 ( .B1(n5847), .B2(n4927), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5110) );
  NAND2_X1 U5434 ( .A1(n4928), .A2(n5111), .ZN(n4927) );
  NAND2_X1 U5435 ( .A1(n4881), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n4880) );
  NAND2_X1 U5436 ( .A1(n5078), .A2(n5077), .ZN(n5409) );
  INV_X1 U5437 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5077) );
  XNOR2_X1 U5438 ( .A(n5082), .B(n5083), .ZN(n7015) );
  OAI21_X1 U5439 ( .B1(n5409), .B2(n4881), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5082) );
  INV_X1 U5440 ( .A(n9399), .ZN(n4984) );
  AND2_X1 U5441 ( .A1(n6922), .A2(n6921), .ZN(n5936) );
  NAND2_X1 U5442 ( .A1(n5973), .A2(n5972), .ZN(n6933) );
  OR2_X1 U5443 ( .A1(n10105), .A2(n4553), .ZN(n4591) );
  AND2_X1 U5444 ( .A1(n4591), .A2(n4590), .ZN(n10115) );
  INV_X1 U5445 ( .A(n10116), .ZN(n4590) );
  NAND2_X1 U5446 ( .A1(n4845), .A2(n4844), .ZN(n9581) );
  NAND2_X1 U5447 ( .A1(n9625), .A2(n9626), .ZN(n9624) );
  AOI21_X1 U5448 ( .B1(n4831), .B2(n8368), .A(n4522), .ZN(n4830) );
  NAND2_X1 U5449 ( .A1(n4834), .A2(n8027), .ZN(n4833) );
  AND2_X1 U5450 ( .A1(n8397), .A2(n4833), .ZN(n4831) );
  OR2_X1 U5451 ( .A1(n9740), .A2(n8368), .ZN(n4832) );
  NAND2_X1 U5452 ( .A1(n9767), .A2(n8395), .ZN(n9748) );
  INV_X1 U5453 ( .A(n4800), .ZN(n4799) );
  OAI21_X1 U5454 ( .B1(n8364), .B2(n4801), .A(n8363), .ZN(n4800) );
  NAND2_X1 U5455 ( .A1(n7889), .A2(n7892), .ZN(n4801) );
  NAND2_X1 U5456 ( .A1(n4746), .A2(n8187), .ZN(n7791) );
  NAND2_X1 U5457 ( .A1(n9943), .A2(n9934), .ZN(n4746) );
  AOI21_X1 U5458 ( .B1(n4815), .B2(n4817), .A(n4537), .ZN(n4813) );
  NAND2_X1 U5459 ( .A1(n9936), .A2(n9985), .ZN(n9938) );
  NAND2_X1 U5460 ( .A1(n7720), .A2(n8133), .ZN(n7781) );
  AND2_X1 U5461 ( .A1(n8152), .A2(n8048), .ZN(n8130) );
  NAND2_X1 U5462 ( .A1(n10159), .A2(n7472), .ZN(n4812) );
  OAI21_X1 U5463 ( .B1(n7484), .B2(n7485), .A(n7483), .ZN(n8037) );
  INV_X1 U5464 ( .A(n10167), .ZN(n9947) );
  INV_X1 U5465 ( .A(n9945), .ZN(n10170) );
  NAND2_X1 U5466 ( .A1(n6235), .A2(n6234), .ZN(n9850) );
  INV_X1 U5467 ( .A(n6503), .ZN(n4992) );
  INV_X1 U5468 ( .A(n4993), .ZN(n4766) );
  NAND2_X1 U5469 ( .A1(n5598), .A2(n5597), .ZN(n5600) );
  NAND2_X1 U5470 ( .A1(n5869), .A2(n4995), .ZN(n4841) );
  XNOR2_X1 U5471 ( .A(n5893), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6488) );
  NAND2_X1 U5472 ( .A1(n5892), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5893) );
  NAND2_X1 U5473 ( .A1(n5507), .A2(n5506), .ZN(n4951) );
  AND2_X1 U5474 ( .A1(n5526), .A2(n5511), .ZN(n5512) );
  NAND2_X1 U5475 ( .A1(n5508), .A2(n5506), .ZN(n4952) );
  NAND2_X1 U5476 ( .A1(n4966), .A2(n5479), .ZN(n5485) );
  NAND2_X1 U5477 ( .A1(n4977), .A2(n5361), .ZN(n4976) );
  INV_X1 U5478 ( .A(n5363), .ZN(n4977) );
  INV_X1 U5479 ( .A(n8626), .ZN(n10251) );
  NAND2_X1 U5480 ( .A1(n4581), .A2(n4866), .ZN(n4580) );
  NAND2_X1 U5481 ( .A1(n4870), .A2(n8345), .ZN(n4867) );
  OAI21_X1 U5482 ( .B1(n4869), .B2(n4872), .A(n4865), .ZN(n4864) );
  NAND2_X1 U5483 ( .A1(n4870), .A2(n4872), .ZN(n4865) );
  AOI22_X1 U5484 ( .A1(n4870), .A2(n10246), .B1(n8347), .B2(n10246), .ZN(n4868) );
  NAND3_X1 U5485 ( .A1(n8322), .A2(n8321), .A3(n4857), .ZN(n8521) );
  OR2_X1 U5486 ( .A1(n8538), .A2(n8542), .ZN(n4857) );
  NAND2_X1 U5487 ( .A1(n7975), .A2(n7977), .ZN(n8281) );
  INV_X1 U5488 ( .A(n7238), .ZN(n10285) );
  AND3_X1 U5489 ( .A1(n5461), .A2(n5460), .A3(n5459), .ZN(n8595) );
  NAND2_X1 U5490 ( .A1(n5833), .A2(n5832), .ZN(n5834) );
  NAND2_X1 U5491 ( .A1(n4629), .A2(n4628), .ZN(n4627) );
  INV_X1 U5492 ( .A(n8333), .ZN(n9083) );
  INV_X1 U5493 ( .A(n8531), .ZN(n9218) );
  OAI211_X1 U5494 ( .C1(n6861), .C2(n6855), .A(n4610), .B(n4609), .ZN(n6856)
         );
  NOR2_X1 U5495 ( .A1(n6849), .A2(n6790), .ZN(n4610) );
  NAND2_X1 U5496 ( .A1(n6861), .A2(n6855), .ZN(n4609) );
  AND2_X1 U5497 ( .A1(n5240), .A2(n5239), .ZN(n8634) );
  NAND2_X1 U5498 ( .A1(n10331), .A2(n6994), .ZN(n6996) );
  NOR2_X1 U5499 ( .A1(n6996), .A2(n6995), .ZN(n7062) );
  INV_X1 U5500 ( .A(n7015), .ZN(n9194) );
  NAND2_X1 U5501 ( .A1(n4608), .A2(n4607), .ZN(n4606) );
  OR2_X1 U5502 ( .A1(n8667), .A2(n10295), .ZN(n4608) );
  AOI21_X1 U5503 ( .B1(n8668), .B2(n10336), .A(n10330), .ZN(n4607) );
  OAI21_X1 U5504 ( .B1(n8461), .B2(n4894), .A(n4893), .ZN(n4892) );
  NAND2_X1 U5505 ( .A1(n8461), .A2(n8453), .ZN(n4893) );
  NOR2_X1 U5506 ( .A1(n9038), .A2(n4895), .ZN(n4894) );
  INV_X1 U5507 ( .A(n8453), .ZN(n4895) );
  OR2_X1 U5508 ( .A1(n9037), .A2(n4896), .ZN(n4891) );
  NAND2_X1 U5509 ( .A1(n8454), .A2(n8453), .ZN(n4896) );
  OR2_X1 U5510 ( .A1(n9046), .A2(n8678), .ZN(n9052) );
  INV_X1 U5511 ( .A(n4737), .ZN(n4736) );
  XNOR2_X1 U5512 ( .A(n9037), .B(n5802), .ZN(n9284) );
  NAND2_X1 U5513 ( .A1(n7738), .A2(n7737), .ZN(n7751) );
  NAND2_X1 U5514 ( .A1(n9259), .A2(n7217), .ZN(n9254) );
  NAND2_X1 U5515 ( .A1(n6377), .A2(n6376), .ZN(n9811) );
  AND2_X1 U5516 ( .A1(n6508), .A2(n9483), .ZN(n6509) );
  NAND2_X1 U5517 ( .A1(n6414), .A2(n6413), .ZN(n9799) );
  NAND2_X1 U5518 ( .A1(n7920), .A2(n8096), .ZN(n6414) );
  INV_X1 U5519 ( .A(n9522), .ZN(n10168) );
  NAND2_X1 U5520 ( .A1(n6359), .A2(n6358), .ZN(n9816) );
  NAND2_X1 U5521 ( .A1(n8269), .A2(n4964), .ZN(n4958) );
  NAND2_X1 U5522 ( .A1(n8234), .A2(n6968), .ZN(n8269) );
  OR3_X1 U5523 ( .A1(n6443), .A2(n6442), .A3(n6441), .ZN(n9627) );
  NAND2_X1 U5524 ( .A1(n4492), .A2(n5925), .ZN(n9530) );
  NOR2_X1 U5525 ( .A1(n5924), .A2(n5923), .ZN(n5925) );
  OR2_X1 U5526 ( .A1(n5981), .A2(n6689), .ZN(n5957) );
  OR2_X1 U5527 ( .A1(n6003), .A2(n7384), .ZN(n5958) );
  OR2_X1 U5528 ( .A1(n5982), .A2(n5956), .ZN(n5959) );
  NAND2_X1 U5529 ( .A1(n6733), .A2(n6734), .ZN(n6732) );
  NAND2_X1 U5530 ( .A1(n6713), .A2(n6714), .ZN(n6748) );
  NAND2_X1 U5531 ( .A1(n4552), .A2(n4805), .ZN(n4804) );
  INV_X1 U5532 ( .A(n4763), .ZN(n4584) );
  AOI21_X1 U5533 ( .B1(n9517), .B2(n9945), .A(n4764), .ZN(n4763) );
  AND2_X1 U5534 ( .A1(n8098), .A2(n8097), .ZN(n8392) );
  NAND2_X1 U5535 ( .A1(n6432), .A2(n6431), .ZN(n9796) );
  OR2_X1 U5536 ( .A1(n9862), .A2(n7358), .ZN(n10178) );
  NAND2_X1 U5537 ( .A1(n4637), .A2(n4636), .ZN(n5684) );
  NAND2_X1 U5538 ( .A1(n5670), .A2(n5797), .ZN(n4637) );
  NAND2_X1 U5539 ( .A1(n5669), .A2(n5782), .ZN(n4636) );
  NAND2_X1 U5540 ( .A1(n4635), .A2(n4633), .ZN(n5687) );
  NAND2_X1 U5541 ( .A1(n4634), .A2(n5797), .ZN(n4633) );
  OR2_X1 U5542 ( .A1(n5684), .A2(n5681), .ZN(n4635) );
  OAI21_X1 U5543 ( .B1(n5684), .B2(n4542), .A(n4510), .ZN(n4634) );
  AOI21_X1 U5544 ( .B1(n4791), .B2(n4789), .A(n5709), .ZN(n5715) );
  NOR2_X1 U5545 ( .A1(n5704), .A2(n4790), .ZN(n4789) );
  INV_X1 U5546 ( .A(n4771), .ZN(n4770) );
  NOR2_X1 U5547 ( .A1(n5741), .A2(n9245), .ZN(n4774) );
  NAND2_X1 U5548 ( .A1(n4631), .A2(n4528), .ZN(n5727) );
  NAND2_X1 U5549 ( .A1(n4640), .A2(n4638), .ZN(n4776) );
  NOR2_X1 U5550 ( .A1(n4639), .A2(n9120), .ZN(n4638) );
  INV_X1 U5551 ( .A(n5758), .ZN(n4639) );
  NOR2_X1 U5552 ( .A1(n4620), .A2(n9065), .ZN(n4619) );
  INV_X1 U5553 ( .A(n4622), .ZN(n4620) );
  AND2_X1 U5554 ( .A1(n8412), .A2(n8410), .ZN(n8150) );
  OAI21_X1 U5555 ( .B1(n4659), .B2(n4529), .A(n4657), .ZN(n4656) );
  NOR2_X1 U5556 ( .A1(n4658), .A2(n8408), .ZN(n4657) );
  AOI21_X1 U5557 ( .B1(n8088), .B2(n8178), .A(n4660), .ZN(n4659) );
  AOI21_X1 U5558 ( .B1(n4662), .B2(n8405), .A(n8107), .ZN(n4661) );
  OAI21_X1 U5559 ( .B1(n8088), .B2(n8087), .A(n8404), .ZN(n4662) );
  NAND2_X1 U5560 ( .A1(n8112), .A2(n8413), .ZN(n4655) );
  AND2_X1 U5561 ( .A1(n4988), .A2(n4712), .ZN(n4711) );
  OR2_X1 U5562 ( .A1(n9409), .A2(n4714), .ZN(n4712) );
  INV_X1 U5563 ( .A(n6320), .ZN(n4714) );
  AND2_X1 U5564 ( .A1(n9415), .A2(n4989), .ZN(n4988) );
  NAND2_X1 U5565 ( .A1(n9460), .A2(n4990), .ZN(n4989) );
  INV_X1 U5566 ( .A(n9461), .ZN(n4990) );
  INV_X1 U5567 ( .A(n7469), .ZN(n4822) );
  INV_X1 U5568 ( .A(n5324), .ZN(n4938) );
  INV_X1 U5569 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n5305) );
  INV_X1 U5570 ( .A(n5288), .ZN(n4945) );
  INV_X1 U5571 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4613) );
  INV_X1 U5572 ( .A(n8286), .ZN(n4874) );
  INV_X1 U5573 ( .A(n5795), .ZN(n4779) );
  OR2_X1 U5574 ( .A1(n9274), .A2(n8614), .ZN(n5788) );
  INV_X1 U5575 ( .A(n5762), .ZN(n5034) );
  INV_X1 U5576 ( .A(n5064), .ZN(n4902) );
  INV_X1 U5577 ( .A(n5756), .ZN(n5040) );
  AND2_X1 U5578 ( .A1(n9143), .A2(n9144), .ZN(n5505) );
  AND2_X1 U5579 ( .A1(n4686), .A2(n4684), .ZN(n4683) );
  INV_X1 U5580 ( .A(n9174), .ZN(n4684) );
  INV_X1 U5581 ( .A(n4693), .ZN(n4691) );
  OR2_X1 U5582 ( .A1(n5457), .A2(n5456), .ZN(n5472) );
  NOR2_X1 U5583 ( .A1(n9346), .A2(n7993), .ZN(n4722) );
  NOR2_X1 U5584 ( .A1(n9245), .A2(n5053), .ZN(n5052) );
  INV_X1 U5585 ( .A(n5737), .ZN(n5053) );
  NAND2_X1 U5586 ( .A1(n5055), .A2(n7987), .ZN(n5054) );
  INV_X1 U5587 ( .A(n7988), .ZN(n5055) );
  INV_X1 U5588 ( .A(n10375), .ZN(n5015) );
  INV_X1 U5589 ( .A(n5673), .ZN(n5806) );
  NAND2_X1 U5590 ( .A1(n10251), .A2(n8576), .ZN(n5807) );
  AND2_X1 U5591 ( .A1(n7014), .A2(n6616), .ZN(n6623) );
  NAND2_X1 U5592 ( .A1(n8580), .A2(n6546), .ZN(n5808) );
  INV_X1 U5593 ( .A(n4916), .ZN(n4910) );
  INV_X1 U5594 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5090) );
  INV_X1 U5595 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5109) );
  AND2_X1 U5596 ( .A1(n4999), .A2(n7765), .ZN(n4998) );
  NAND2_X1 U5597 ( .A1(n7833), .A2(n7834), .ZN(n4999) );
  NAND2_X1 U5598 ( .A1(n4558), .A2(n6135), .ZN(n4983) );
  NOR2_X1 U5599 ( .A1(n6201), .A2(n7109), .ZN(n6220) );
  NOR2_X1 U5600 ( .A1(n8146), .A2(n8019), .ZN(n4667) );
  OAI21_X1 U5601 ( .B1(n8095), .B2(n4649), .A(n4644), .ZN(n8104) );
  OR2_X1 U5602 ( .A1(n8149), .A2(n4652), .ZN(n4649) );
  NAND2_X1 U5603 ( .A1(n4648), .A2(n4645), .ZN(n4644) );
  OAI21_X1 U5604 ( .B1(n8109), .B2(n8108), .A(n8262), .ZN(n4665) );
  NAND2_X1 U5605 ( .A1(n9533), .A2(n9534), .ZN(n9535) );
  INV_X1 U5606 ( .A(n4587), .ZN(n9532) );
  AND2_X1 U5607 ( .A1(n8392), .A2(n9577), .ZN(n8219) );
  AND2_X1 U5608 ( .A1(n8099), .A2(n9778), .ZN(n8259) );
  OR2_X1 U5609 ( .A1(n9783), .A2(n9597), .ZN(n8415) );
  INV_X1 U5610 ( .A(n4831), .ZN(n4828) );
  INV_X1 U5611 ( .A(n4830), .ZN(n4829) );
  AND2_X1 U5612 ( .A1(n6288), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n6304) );
  INV_X1 U5613 ( .A(n7780), .ZN(n4817) );
  NOR2_X1 U5614 ( .A1(n6092), .A2(n7513), .ZN(n6118) );
  AND2_X1 U5615 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6004) );
  NOR2_X1 U5616 ( .A1(n6033), .A2(n8893), .ZN(n6052) );
  OR2_X1 U5617 ( .A1(n6925), .A2(n6963), .ZN(n8237) );
  INV_X1 U5618 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5901) );
  NAND2_X1 U5619 ( .A1(n5884), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5886) );
  AND2_X1 U5620 ( .A1(n5479), .A2(n5468), .ZN(n5477) );
  INV_X1 U5621 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5858) );
  INV_X1 U5622 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5860) );
  INV_X1 U5623 ( .A(n4971), .ZN(n4970) );
  AOI21_X1 U5624 ( .B1(n4971), .B2(n4973), .A(n4969), .ZN(n4968) );
  OR2_X1 U5625 ( .A1(n6110), .A2(n6109), .ZN(n6114) );
  NOR2_X1 U5626 ( .A1(n6114), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6158) );
  INV_X1 U5627 ( .A(n5206), .ZN(n4933) );
  NAND2_X1 U5628 ( .A1(n8007), .A2(n6631), .ZN(n4585) );
  OR2_X1 U5629 ( .A1(n8007), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n4586) );
  INV_X1 U5630 ( .A(n8347), .ZN(n4869) );
  NOR2_X1 U5631 ( .A1(n8527), .A2(n4878), .ZN(n4877) );
  INV_X1 U5632 ( .A(n8280), .ZN(n4878) );
  OAI211_X1 U5633 ( .C1(n6551), .C2(n4860), .A(n4861), .B(n6561), .ZN(n7125)
         );
  NAND2_X1 U5634 ( .A1(n4862), .A2(n4858), .ZN(n4861) );
  CLKBUF_X1 U5635 ( .A(n7822), .Z(n10268) );
  NAND2_X1 U5636 ( .A1(n5413), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n5457) );
  INV_X1 U5637 ( .A(n5415), .ZN(n5413) );
  NOR2_X1 U5638 ( .A1(n7963), .A2(n4884), .ZN(n4883) );
  INV_X1 U5639 ( .A(n7961), .ZN(n4884) );
  NOR2_X1 U5640 ( .A1(n5801), .A2(n7021), .ZN(n4628) );
  AND2_X1 U5641 ( .A1(n5596), .A2(n5595), .ZN(n8333) );
  AND2_X1 U5642 ( .A1(n5538), .A2(n5537), .ZN(n8540) );
  AND4_X1 U5643 ( .A1(n5437), .A2(n5436), .A3(n5435), .A4(n5434), .ZN(n8531)
         );
  NOR2_X1 U5644 ( .A1(n7418), .A2(n4574), .ZN(n7624) );
  AND2_X1 U5645 ( .A1(n4525), .A2(n5076), .ZN(n4885) );
  NOR2_X1 U5646 ( .A1(n4869), .A2(n9058), .ZN(n9045) );
  AND2_X1 U5647 ( .A1(n8458), .A2(n9045), .ZN(n8679) );
  NAND2_X1 U5648 ( .A1(n4735), .A2(n9062), .ZN(n9058) );
  OR2_X1 U5649 ( .A1(n9291), .A2(n9066), .ZN(n8451) );
  AND2_X1 U5650 ( .A1(n5769), .A2(n5767), .ZN(n9082) );
  INV_X1 U5651 ( .A(n9082), .ZN(n9072) );
  NAND2_X1 U5652 ( .A1(n9105), .A2(n8449), .ZN(n9091) );
  NAND2_X1 U5653 ( .A1(n4671), .A2(n4538), .ZN(n9088) );
  NAND2_X1 U5654 ( .A1(n9121), .A2(n4899), .ZN(n4671) );
  NAND2_X1 U5655 ( .A1(n4899), .A2(n4903), .ZN(n4898) );
  NOR2_X1 U5656 ( .A1(n9122), .A2(n9300), .ZN(n9105) );
  NAND2_X1 U5657 ( .A1(n9158), .A2(n5505), .ZN(n9142) );
  NOR2_X1 U5658 ( .A1(n9310), .A2(n4725), .ZN(n4724) );
  INV_X1 U5659 ( .A(n4726), .ZN(n4725) );
  AND2_X1 U5660 ( .A1(n5755), .A2(n9144), .ZN(n9160) );
  INV_X1 U5661 ( .A(n9160), .ZN(n9153) );
  OR2_X1 U5662 ( .A1(n5398), .A2(n5397), .ZN(n5415) );
  NAND2_X1 U5663 ( .A1(n7859), .A2(n4504), .ZN(n9252) );
  NAND2_X1 U5664 ( .A1(n5054), .A2(n5737), .ZN(n9244) );
  OAI21_X1 U5665 ( .B1(n7991), .B2(n4888), .A(n7994), .ZN(n7996) );
  NAND2_X1 U5666 ( .A1(n7996), .A2(n7995), .ZN(n8438) );
  NAND2_X1 U5667 ( .A1(n7859), .A2(n9928), .ZN(n8000) );
  AND4_X1 U5668 ( .A1(n5384), .A2(n5383), .A3(n5382), .A4(n5381), .ZN(n9243)
         );
  OR2_X1 U5669 ( .A1(n5315), .A2(n5314), .ZN(n5333) );
  INV_X1 U5670 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n7827) );
  AND4_X1 U5671 ( .A1(n5360), .A2(n5359), .A3(n5358), .A4(n5357), .ZN(n7965)
         );
  NAND2_X1 U5672 ( .A1(n5022), .A2(n5027), .ZN(n7871) );
  NAND2_X1 U5673 ( .A1(n7752), .A2(n4516), .ZN(n5022) );
  NAND2_X1 U5674 ( .A1(n4731), .A2(n4730), .ZN(n7878) );
  NOR2_X1 U5675 ( .A1(n4732), .A2(n7758), .ZN(n4730) );
  NAND2_X1 U5676 ( .A1(n10454), .A2(n4733), .ZN(n4732) );
  AND4_X1 U5677 ( .A1(n5300), .A2(n5299), .A3(n5298), .A4(n5297), .ZN(n7744)
         );
  NOR3_X1 U5678 ( .A1(n10357), .A2(n4734), .A3(n7758), .ZN(n7756) );
  NOR2_X1 U5679 ( .A1(n10357), .A2(n4734), .ZN(n7755) );
  NAND2_X1 U5680 ( .A1(n5005), .A2(n5003), .ZN(n7495) );
  INV_X1 U5681 ( .A(n5701), .ZN(n5004) );
  OAI21_X1 U5682 ( .B1(n5227), .B2(n5698), .A(n4503), .ZN(n7450) );
  NAND2_X1 U5683 ( .A1(n5006), .A2(n5696), .ZN(n7451) );
  NAND2_X1 U5684 ( .A1(n5227), .A2(n5009), .ZN(n5006) );
  NAND2_X1 U5685 ( .A1(n5244), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5280) );
  INV_X1 U5686 ( .A(n6780), .ZN(n5447) );
  AND4_X1 U5687 ( .A1(n5199), .A2(n5198), .A3(n5197), .A4(n5196), .ZN(n7301)
         );
  NAND2_X1 U5688 ( .A1(n4571), .A2(n10379), .ZN(n10377) );
  INV_X1 U5689 ( .A(n10385), .ZN(n8427) );
  NAND2_X1 U5690 ( .A1(n7322), .A2(n10414), .ZN(n7321) );
  NOR2_X1 U5691 ( .A1(n7262), .A2(n8576), .ZN(n7265) );
  AND2_X1 U5692 ( .A1(n7265), .A2(n10250), .ZN(n7322) );
  OAI21_X1 U5693 ( .B1(n5673), .B2(n7270), .A(n5807), .ZN(n7163) );
  AND2_X1 U5694 ( .A1(n5671), .A2(n5682), .ZN(n7164) );
  NAND2_X1 U5695 ( .A1(n5807), .A2(n5806), .ZN(n7269) );
  NAND2_X1 U5696 ( .A1(n7025), .A2(n5808), .ZN(n7029) );
  NAND2_X1 U5697 ( .A1(n4719), .A2(n10403), .ZN(n7262) );
  AND2_X1 U5698 ( .A1(n5634), .A2(n5633), .ZN(n9273) );
  NAND2_X1 U5699 ( .A1(n9042), .A2(n9041), .ZN(n9043) );
  NAND2_X1 U5700 ( .A1(n5548), .A2(n5547), .ZN(n9296) );
  NAND2_X1 U5701 ( .A1(n5481), .A2(n5480), .ZN(n9315) );
  NAND2_X1 U5702 ( .A1(n5021), .A2(n5814), .ZN(n7233) );
  OR2_X1 U5703 ( .A1(n7311), .A2(n5667), .ZN(n5021) );
  AND3_X1 U5704 ( .A1(n5125), .A2(n5124), .A3(n5123), .ZN(n10408) );
  INV_X1 U5705 ( .A(n10444), .ZN(n10453) );
  AND3_X1 U5706 ( .A1(n8428), .A2(n7011), .A3(n8427), .ZN(n7212) );
  INV_X1 U5707 ( .A(n7021), .ZN(n10404) );
  NAND2_X1 U5708 ( .A1(n6767), .A2(n10400), .ZN(n10385) );
  AND2_X1 U5709 ( .A1(n5100), .A2(n4679), .ZN(n4928) );
  XNOR2_X1 U5710 ( .A(n5846), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6607) );
  OAI21_X1 U5711 ( .B1(n5409), .B2(P2_IR_REG_17__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5428) );
  NOR2_X1 U5712 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_3__SCAN_IN), .ZN(
        n5068) );
  OR2_X1 U5713 ( .A1(n6454), .A2(n8883), .ZN(n6468) );
  NAND2_X1 U5714 ( .A1(n6209), .A2(n6208), .ZN(n7907) );
  NAND2_X1 U5715 ( .A1(n9479), .A2(n9481), .ZN(n9408) );
  NAND2_X1 U5716 ( .A1(n9408), .A2(n9409), .ZN(n9407) );
  NOR2_X1 U5717 ( .A1(n4702), .A2(n4698), .ZN(n4697) );
  INV_X1 U5718 ( .A(n7511), .ZN(n4698) );
  INV_X1 U5719 ( .A(n6135), .ZN(n4702) );
  NAND2_X1 U5720 ( .A1(n9459), .A2(n9461), .ZN(n9458) );
  NAND2_X1 U5721 ( .A1(n9407), .A2(n6320), .ZN(n9459) );
  OR2_X1 U5722 ( .A1(n6184), .A2(n6183), .ZN(n6201) );
  NAND2_X1 U5723 ( .A1(n9442), .A2(n4533), .ZN(n9482) );
  INV_X1 U5724 ( .A(n9423), .ZN(n4707) );
  NAND2_X1 U5725 ( .A1(n4704), .A2(n4703), .ZN(n4708) );
  AOI21_X1 U5726 ( .B1(n4499), .B2(n6392), .A(n4551), .ZN(n4703) );
  NAND2_X1 U5727 ( .A1(n6220), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n6236) );
  OR2_X1 U5728 ( .A1(n5982), .A2(n5920), .ZN(n5922) );
  AND2_X1 U5729 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6870) );
  AOI21_X1 U5730 ( .B1(n6836), .B2(n4501), .A(n4539), .ZN(n4593) );
  NAND2_X1 U5731 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6896) );
  NAND2_X1 U5732 ( .A1(n6748), .A2(n4592), .ZN(n10056) );
  OR2_X1 U5733 ( .A1(n6749), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4592) );
  NAND2_X1 U5734 ( .A1(n6910), .A2(n6911), .ZN(n7112) );
  NAND2_X1 U5735 ( .A1(n7112), .A2(n4596), .ZN(n10081) );
  OR2_X1 U5736 ( .A1(n7113), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4596) );
  NOR2_X1 U5737 ( .A1(n10081), .A2(n10080), .ZN(n10079) );
  NOR2_X1 U5738 ( .A1(n10079), .A2(n4595), .ZN(n10094) );
  AND2_X1 U5739 ( .A1(n10084), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n4595) );
  XNOR2_X1 U5740 ( .A(n4587), .B(n9541), .ZN(n7115) );
  NAND2_X1 U5741 ( .A1(n7115), .A2(n6203), .ZN(n9533) );
  NOR2_X1 U5742 ( .A1(n10115), .A2(n4589), .ZN(n10130) );
  NOR2_X1 U5743 ( .A1(n9547), .A2(n6239), .ZN(n4589) );
  NOR2_X1 U5744 ( .A1(n10128), .A2(n4599), .ZN(n10145) );
  NOR2_X1 U5745 ( .A1(n9549), .A2(n4600), .ZN(n4599) );
  NOR2_X1 U5746 ( .A1(n10145), .A2(n10144), .ZN(n10143) );
  XNOR2_X1 U5747 ( .A(n4597), .B(P1_REG2_REG_19__SCAN_IN), .ZN(n9556) );
  OR2_X1 U5748 ( .A1(n10143), .A2(n4598), .ZN(n4597) );
  AND2_X1 U5749 ( .A1(n10149), .A2(P1_REG2_REG_18__SCAN_IN), .ZN(n4598) );
  NAND2_X1 U5750 ( .A1(n8010), .A2(n8009), .ZN(n9566) );
  NOR2_X1 U5751 ( .A1(n4808), .A2(n4807), .ZN(n4806) );
  INV_X1 U5752 ( .A(n4552), .ZN(n4807) );
  INV_X1 U5753 ( .A(n9595), .ZN(n4808) );
  INV_X1 U5754 ( .A(n4809), .ZN(n4805) );
  AND2_X1 U5755 ( .A1(n8420), .A2(n9516), .ZN(n4764) );
  NOR2_X1 U5756 ( .A1(n8219), .A2(n8259), .ZN(n8418) );
  AOI21_X1 U5757 ( .B1(n9605), .B2(n4751), .A(n8147), .ZN(n4750) );
  NOR2_X1 U5758 ( .A1(n4752), .A2(n4749), .ZN(n4748) );
  NAND2_X1 U5759 ( .A1(n9619), .A2(n8356), .ZN(n9607) );
  AND2_X1 U5760 ( .A1(n5067), .A2(n8383), .ZN(n4819) );
  AND2_X1 U5761 ( .A1(n5063), .A2(n8377), .ZN(n4824) );
  OR2_X1 U5762 ( .A1(n6324), .A2(n6323), .ZN(n6344) );
  OR2_X1 U5763 ( .A1(n9826), .A2(n9718), .ZN(n9683) );
  NOR2_X1 U5764 ( .A1(n9826), .A2(n4851), .ZN(n4850) );
  INV_X1 U5765 ( .A(n4852), .ZN(n4851) );
  OAI21_X1 U5766 ( .B1(n9767), .B2(n4757), .A(n4753), .ZN(n9715) );
  AOI21_X1 U5767 ( .B1(n4756), .B2(n4755), .A(n4754), .ZN(n4753) );
  INV_X1 U5768 ( .A(n8398), .ZN(n4754) );
  INV_X1 U5769 ( .A(n8395), .ZN(n4755) );
  NAND2_X1 U5770 ( .A1(n9761), .A2(n4854), .ZN(n9731) );
  NAND2_X1 U5771 ( .A1(n9761), .A2(n4834), .ZN(n9741) );
  AND2_X1 U5772 ( .A1(n8396), .A2(n8075), .ZN(n9749) );
  AND2_X1 U5773 ( .A1(n8195), .A2(n9750), .ZN(n9769) );
  INV_X1 U5774 ( .A(n7892), .ZN(n4802) );
  INV_X1 U5775 ( .A(n9769), .ZN(n9758) );
  AOI21_X1 U5776 ( .B1(n4744), .B2(n9942), .A(n4742), .ZN(n4741) );
  INV_X1 U5777 ( .A(n8064), .ZN(n4742) );
  NAND2_X1 U5778 ( .A1(n6140), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n6162) );
  INV_X1 U5779 ( .A(n4848), .ZN(n4846) );
  NOR2_X1 U5780 ( .A1(n4848), .A2(n7400), .ZN(n10161) );
  NOR2_X1 U5781 ( .A1(n7400), .A2(n4849), .ZN(n7591) );
  NOR2_X1 U5782 ( .A1(n7400), .A2(n7466), .ZN(n7528) );
  INV_X1 U5783 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n8893) );
  NAND2_X1 U5784 ( .A1(n7565), .A2(n8169), .ZN(n4663) );
  NAND2_X1 U5785 ( .A1(n4643), .A2(n6966), .ZN(n8238) );
  NOR2_X1 U5786 ( .A1(n7357), .A2(n6882), .ZN(n6955) );
  XNOR2_X1 U5787 ( .A(n5649), .B(SI_30_), .ZN(n8351) );
  XNOR2_X1 U5788 ( .A(n5629), .B(n5620), .ZN(n8471) );
  NAND2_X1 U5789 ( .A1(n5579), .A2(n5578), .ZN(n5581) );
  AND2_X1 U5790 ( .A1(n5599), .A2(n5585), .ZN(n5597) );
  XNOR2_X1 U5791 ( .A(n5561), .B(n5560), .ZN(n7920) );
  NAND2_X1 U5792 ( .A1(n4949), .A2(n4953), .ZN(n5542) );
  NOR2_X1 U5793 ( .A1(n4531), .A2(n4717), .ZN(n4716) );
  INV_X1 U5794 ( .A(n5882), .ZN(n4717) );
  INV_X1 U5795 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U5796 ( .A1(n6196), .A2(n5882), .ZN(n6233) );
  NAND2_X1 U5797 ( .A1(n4967), .A2(n4971), .ZN(n5405) );
  NAND2_X1 U5798 ( .A1(n5363), .A2(n4974), .ZN(n4967) );
  NAND2_X1 U5799 ( .A1(n4939), .A2(n4943), .ZN(n5325) );
  NAND2_X1 U5800 ( .A1(n4941), .A2(n4940), .ZN(n4939) );
  NAND2_X1 U5801 ( .A1(n4942), .A2(n5288), .ZN(n5304) );
  NAND2_X1 U5802 ( .A1(n5287), .A2(n5062), .ZN(n4942) );
  NAND2_X1 U5803 ( .A1(n4934), .A2(n5206), .ZN(n5220) );
  NAND2_X1 U5804 ( .A1(n5204), .A2(n5203), .ZN(n4934) );
  INV_X1 U5805 ( .A(n5926), .ZN(n5867) );
  AND2_X1 U5806 ( .A1(n5577), .A2(n5576), .ZN(n8522) );
  AND2_X1 U5807 ( .A1(n7608), .A2(n7600), .ZN(n4886) );
  NAND2_X1 U5808 ( .A1(n7601), .A2(n7600), .ZN(n7606) );
  NAND2_X1 U5809 ( .A1(n8574), .A2(n6555), .ZN(n10247) );
  OAI21_X1 U5810 ( .B1(n7243), .B2(n7242), .A(n6582), .ZN(n7330) );
  AND3_X1 U5811 ( .A1(n5476), .A2(n5475), .A3(n5474), .ZN(n8615) );
  AND4_X1 U5812 ( .A1(n5339), .A2(n5338), .A3(n5337), .A4(n5336), .ZN(n10261)
         );
  NAND2_X1 U5813 ( .A1(n8281), .A2(n4877), .ZN(n8589) );
  NAND2_X1 U5814 ( .A1(n8281), .A2(n8280), .ZN(n8528) );
  AND2_X1 U5815 ( .A1(n5133), .A2(n5132), .ZN(n8424) );
  NOR2_X1 U5816 ( .A1(n4495), .A2(n5126), .ZN(n5131) );
  AND2_X1 U5817 ( .A1(n8302), .A2(n8297), .ZN(n4887) );
  INV_X1 U5818 ( .A(n8549), .ZN(n8302) );
  NAND2_X1 U5819 ( .A1(n8495), .A2(n8297), .ZN(n8550) );
  AND2_X1 U5820 ( .A1(n10279), .A2(n10366), .ZN(n10257) );
  AND4_X1 U5821 ( .A1(n5285), .A2(n5284), .A3(n5283), .A4(n5282), .ZN(n7736)
         );
  NAND2_X1 U5822 ( .A1(n8505), .A2(n8506), .ZN(n8582) );
  NAND2_X1 U5823 ( .A1(n6551), .A2(n8577), .ZN(n8574) );
  CLKBUF_X1 U5824 ( .A(n8494), .Z(n8591) );
  NAND2_X1 U5825 ( .A1(n8602), .A2(n8327), .ZN(n4856) );
  NAND2_X1 U5826 ( .A1(n6620), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10292) );
  XNOR2_X1 U5827 ( .A(n5836), .B(P2_IR_REG_22__SCAN_IN), .ZN(n7014) );
  NOR2_X1 U5828 ( .A1(n4788), .A2(n4530), .ZN(n4787) );
  NAND4_X1 U5829 ( .A1(n5108), .A2(n5107), .A3(n5106), .A4(n5105), .ZN(n8626)
         );
  AND2_X1 U5830 ( .A1(n5137), .A2(n5136), .ZN(n5000) );
  INV_X1 U5831 ( .A(n8424), .ZN(n8629) );
  NAND2_X1 U5832 ( .A1(n8630), .A2(n4568), .ZN(n6822) );
  NAND2_X1 U5833 ( .A1(n6822), .A2(n6821), .ZN(n6993) );
  NAND2_X1 U5834 ( .A1(n5074), .A2(n5056), .ZN(n5310) );
  NOR2_X1 U5835 ( .A1(n7062), .A2(n7063), .ZN(n7065) );
  NAND2_X1 U5836 ( .A1(n7065), .A2(n4601), .ZN(n7143) );
  NOR2_X1 U5837 ( .A1(n4603), .A2(n4602), .ZN(n4601) );
  NOR2_X1 U5838 ( .A1(n7075), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n4602) );
  INV_X1 U5839 ( .A(n7144), .ZN(n4603) );
  NOR2_X1 U5840 ( .A1(n7339), .A2(n7340), .ZN(n7342) );
  NOR2_X1 U5841 ( .A1(n7342), .A2(n7341), .ZN(n7418) );
  AND2_X1 U5842 ( .A1(n5349), .A2(n5371), .ZN(n7351) );
  XNOR2_X1 U5843 ( .A(n7624), .B(n7625), .ZN(n7419) );
  NAND2_X1 U5844 ( .A1(n7663), .A2(n7664), .ZN(n7665) );
  NAND2_X1 U5845 ( .A1(n7665), .A2(n7666), .ZN(n8642) );
  AND2_X1 U5846 ( .A1(n6799), .A2(n6797), .ZN(n10330) );
  INV_X1 U5847 ( .A(n9296), .ZN(n8449) );
  NAND2_X1 U5848 ( .A1(n9119), .A2(n5064), .ZN(n9104) );
  NAND2_X1 U5849 ( .A1(n9203), .A2(n9188), .ZN(n9168) );
  NAND2_X1 U5850 ( .A1(n4685), .A2(n4686), .ZN(n9165) );
  OR2_X1 U5851 ( .A1(n8439), .A2(n4688), .ZN(n4685) );
  NAND2_X1 U5852 ( .A1(n4689), .A2(n4692), .ZN(n9182) );
  NAND2_X1 U5853 ( .A1(n8439), .A2(n4693), .ZN(n4689) );
  OAI21_X1 U5854 ( .B1(n7988), .B2(n5048), .A(n5046), .ZN(n9207) );
  NAND2_X1 U5855 ( .A1(n9221), .A2(n8442), .ZN(n9202) );
  AND2_X1 U5856 ( .A1(n9236), .A2(n8441), .ZN(n9223) );
  NAND2_X1 U5857 ( .A1(n4920), .A2(n4923), .ZN(n7867) );
  INV_X1 U5858 ( .A(n7505), .ZN(n4676) );
  NAND2_X1 U5859 ( .A1(n10345), .A2(n7446), .ZN(n7448) );
  NAND2_X1 U5860 ( .A1(n5227), .A2(n5691), .ZN(n10344) );
  NAND2_X1 U5861 ( .A1(n7297), .A2(n4573), .ZN(n4918) );
  NAND2_X1 U5862 ( .A1(n5014), .A2(n5017), .ZN(n10365) );
  NAND2_X1 U5863 ( .A1(n7311), .A2(n5019), .ZN(n5014) );
  NAND2_X1 U5864 ( .A1(n4914), .A2(n7295), .ZN(n10376) );
  OR2_X1 U5865 ( .A1(n7297), .A2(n7296), .ZN(n4914) );
  AND2_X1 U5866 ( .A1(n5191), .A2(n4560), .ZN(n4642) );
  INV_X1 U5867 ( .A(n9254), .ZN(n10355) );
  BUF_X1 U5868 ( .A(n7864), .Z(n9259) );
  INV_X2 U5869 ( .A(n10471), .ZN(n10473) );
  AND2_X1 U5870 ( .A1(n4892), .A2(n10459), .ZN(n4889) );
  INV_X2 U5871 ( .A(n10461), .ZN(n10462) );
  AND2_X1 U5872 ( .A1(n6618), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10400) );
  AND2_X1 U5873 ( .A1(n5030), .A2(n4678), .ZN(n4677) );
  INV_X1 U5874 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n4678) );
  INV_X1 U5875 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7797) );
  XNOR2_X1 U5876 ( .A(n5852), .B(n5851), .ZN(n7799) );
  INV_X1 U5877 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7636) );
  INV_X1 U5878 ( .A(n7014), .ZN(n7637) );
  INV_X1 U5879 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7518) );
  INV_X1 U5880 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n8813) );
  OAI21_X1 U5881 ( .B1(n5409), .B2(n4879), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n5081) );
  NAND2_X1 U5882 ( .A1(n4880), .A2(n5083), .ZN(n4879) );
  INV_X1 U5883 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7287) );
  INV_X1 U5884 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7098) );
  INV_X1 U5885 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7048) );
  INV_X1 U5886 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7046) );
  INV_X1 U5887 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6980) );
  INV_X1 U5888 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6863) );
  INV_X1 U5889 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6686) );
  INV_X1 U5890 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6663) );
  XNOR2_X1 U5891 ( .A(n4611), .B(n5139), .ZN(n6861) );
  NAND2_X1 U5892 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n4611) );
  INV_X1 U5893 ( .A(n6214), .ZN(n7910) );
  XNOR2_X1 U5894 ( .A(n5933), .B(n6387), .ZN(n6922) );
  NAND2_X1 U5895 ( .A1(n9390), .A2(n9388), .ZN(n6512) );
  AND2_X1 U5896 ( .A1(n7429), .A2(n7430), .ZN(n7510) );
  NAND2_X1 U5897 ( .A1(n9458), .A2(n9460), .ZN(n9416) );
  NAND2_X1 U5898 ( .A1(n4705), .A2(n4709), .ZN(n9450) );
  NAND2_X1 U5899 ( .A1(n6391), .A2(n4505), .ZN(n4709) );
  NAND2_X1 U5900 ( .A1(n4710), .A2(n4499), .ZN(n4705) );
  INV_X1 U5901 ( .A(n9530), .ZN(n7084) );
  AND2_X1 U5902 ( .A1(n6532), .A2(n4498), .ZN(n9507) );
  XNOR2_X1 U5903 ( .A(n6370), .B(n7389), .ZN(n9472) );
  OR2_X1 U5904 ( .A1(n7537), .A2(n4558), .ZN(n4981) );
  XNOR2_X1 U5905 ( .A(n5975), .B(n5974), .ZN(n6942) );
  CLKBUF_X1 U5906 ( .A(n6918), .Z(n6919) );
  AND2_X1 U5907 ( .A1(n10226), .A2(n6506), .ZN(n9483) );
  OR3_X1 U5908 ( .A1(n6128), .A2(n6127), .A3(n6126), .ZN(n9522) );
  NOR2_X1 U5909 ( .A1(n5940), .A2(n5939), .ZN(n5943) );
  OR2_X1 U5910 ( .A1(n6889), .A2(n4501), .ZN(n6835) );
  AND2_X1 U5911 ( .A1(n6732), .A2(n6712), .ZN(n6713) );
  INV_X1 U5912 ( .A(n4591), .ZN(n10117) );
  INV_X1 U5913 ( .A(n9566), .ZN(n9981) );
  NAND2_X1 U5914 ( .A1(n4811), .A2(n8387), .ZN(n9571) );
  NAND2_X1 U5915 ( .A1(n9624), .A2(n8412), .ZN(n9612) );
  NAND2_X1 U5916 ( .A1(n4820), .A2(n8383), .ZN(n9606) );
  NAND2_X1 U5917 ( .A1(n4825), .A2(n8377), .ZN(n9652) );
  NAND2_X1 U5918 ( .A1(n6342), .A2(n6341), .ZN(n9823) );
  NAND2_X1 U5919 ( .A1(n4826), .A2(n4830), .ZN(n9713) );
  NAND2_X1 U5920 ( .A1(n9740), .A2(n4831), .ZN(n4826) );
  NAND2_X1 U5921 ( .A1(n4832), .A2(n4833), .ZN(n9729) );
  NAND2_X1 U5922 ( .A1(n4832), .A2(n4831), .ZN(n9837) );
  NAND2_X1 U5923 ( .A1(n9748), .A2(n4756), .ZN(n9726) );
  NAND2_X1 U5924 ( .A1(n4798), .A2(n7892), .ZN(n8365) );
  NAND2_X1 U5925 ( .A1(n7891), .A2(n7890), .ZN(n4798) );
  NAND2_X1 U5926 ( .A1(n6219), .A2(n6218), .ZN(n9856) );
  NAND2_X1 U5927 ( .A1(n4746), .A2(n4744), .ZN(n7893) );
  NAND2_X1 U5928 ( .A1(n6182), .A2(n6181), .ZN(n9956) );
  NAND2_X1 U5929 ( .A1(n7781), .A2(n7780), .ZN(n9935) );
  NAND2_X1 U5930 ( .A1(n4812), .A2(n7473), .ZN(n7476) );
  NAND2_X1 U5931 ( .A1(n7521), .A2(n7469), .ZN(n7582) );
  NAND2_X1 U5932 ( .A1(n7199), .A2(n7198), .ZN(n7391) );
  NAND2_X1 U5933 ( .A1(n10181), .A2(n6515), .ZN(n10177) );
  INV_X1 U5934 ( .A(n10177), .ZN(n9957) );
  INV_X1 U5935 ( .A(n10245), .ZN(n10243) );
  NAND2_X1 U5936 ( .A1(n9780), .A2(n4759), .ZN(n9864) );
  AND2_X1 U5937 ( .A1(n9781), .A2(n4760), .ZN(n4759) );
  NAND2_X1 U5938 ( .A1(n4762), .A2(n4761), .ZN(n4760) );
  INV_X1 U5939 ( .A(n10236), .ZN(n10234) );
  AND2_X1 U5940 ( .A1(n6539), .A2(n6505), .ZN(n8270) );
  INV_X1 U5941 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n5871) );
  NAND2_X1 U5942 ( .A1(n4835), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U5943 ( .A1(n4952), .A2(n4950), .ZN(n5527) );
  AND2_X1 U5944 ( .A1(n4951), .A2(n5512), .ZN(n4950) );
  INV_X1 U5945 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8749) );
  INV_X1 U5946 ( .A(n6483), .ZN(n8236) );
  INV_X1 U5947 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8898) );
  INV_X1 U5948 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7286) );
  INV_X1 U5949 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6954) );
  INV_X1 U5950 ( .A(n7106), .ZN(n9541) );
  INV_X1 U5951 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n6949) );
  INV_X1 U5952 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6683) );
  INV_X1 U5953 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n8761) );
  INV_X1 U5954 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6665) );
  NOR2_X1 U5955 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n5903) );
  NAND2_X1 U5956 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n5961) );
  NOR2_X1 U5957 ( .A1(n7702), .A2(n10512), .ZN(n10501) );
  AOI21_X1 U5958 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10499), .ZN(n10498) );
  NOR2_X1 U5959 ( .A1(n10498), .A2(n10497), .ZN(n10496) );
  INV_X1 U5960 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8671) );
  AND2_X1 U5961 ( .A1(n8350), .A2(n4575), .ZN(n4578) );
  OAI21_X1 U5962 ( .B1(n8669), .B2(n9194), .A(n4604), .ZN(P2_U3264) );
  AOI21_X1 U5963 ( .B1(n4606), .B2(n9194), .A(n4605), .ZN(n4604) );
  OAI21_X1 U5964 ( .B1(n10304), .B2(n8671), .A(n8670), .ZN(n4605) );
  OAI21_X1 U5965 ( .B1(n9284), .B2(n9233), .A(n4670), .ZN(n9053) );
  OR2_X1 U5966 ( .A1(n8275), .A2(n8274), .ZN(n4963) );
  INV_X1 U5967 ( .A(n4964), .ZN(n4959) );
  NAND2_X1 U5968 ( .A1(n6835), .A2(n6836), .ZN(n6834) );
  AND2_X1 U5969 ( .A1(n4985), .A2(n4984), .ZN(n4499) );
  INV_X2 U5970 ( .A(n4549), .ZN(n6228) );
  NAND2_X1 U5971 ( .A1(n4511), .A2(n4554), .ZN(n4692) );
  AND2_X1 U5972 ( .A1(n4953), .A2(n5539), .ZN(n4500) );
  AND2_X1 U5973 ( .A1(n5788), .A2(n5789), .ZN(n8461) );
  INV_X1 U5974 ( .A(n9605), .ZN(n4752) );
  AND2_X1 U5975 ( .A1(n6708), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n4501) );
  AND2_X1 U5976 ( .A1(n4943), .A2(n4938), .ZN(n4502) );
  INV_X1 U5977 ( .A(n7441), .ZN(n4913) );
  INV_X1 U5978 ( .A(n8624), .ZN(n4786) );
  AND2_X1 U5979 ( .A1(n9255), .A2(n4722), .ZN(n4504) );
  AND2_X1 U5980 ( .A1(n4985), .A2(n6392), .ZN(n4505) );
  INV_X1 U5981 ( .A(n8412), .ZN(n4751) );
  AND4_X1 U5982 ( .A1(n5071), .A2(n5070), .A3(n5069), .A4(n8924), .ZN(n4507)
         );
  AND2_X1 U5983 ( .A1(n4993), .A2(n5898), .ZN(n4508) );
  INV_X1 U5984 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9369) );
  XNOR2_X1 U5985 ( .A(n9285), .B(n8333), .ZN(n9064) );
  AND2_X1 U5986 ( .A1(n6357), .A2(n6356), .ZN(n4509) );
  NOR2_X1 U5987 ( .A1(n5672), .A2(n5018), .ZN(n4510) );
  NAND2_X1 U5988 ( .A1(n5868), .A2(n4997), .ZN(n4996) );
  INV_X1 U5989 ( .A(n4996), .ZN(n4995) );
  OR2_X1 U5990 ( .A1(n9799), .A2(n9643), .ZN(n8211) );
  NAND2_X1 U5991 ( .A1(n4518), .A2(n8443), .ZN(n4511) );
  AND2_X1 U5992 ( .A1(n7295), .A2(n4911), .ZN(n4512) );
  OR2_X1 U5993 ( .A1(n10274), .A2(n7873), .ZN(n5710) );
  INV_X1 U5994 ( .A(n8397), .ZN(n4758) );
  NAND2_X1 U5995 ( .A1(n4957), .A2(n5512), .ZN(n4956) );
  INV_X1 U5996 ( .A(n9845), .ZN(n4834) );
  NAND2_X1 U5997 ( .A1(n8355), .A2(n7237), .ZN(n5844) );
  AND2_X1 U5998 ( .A1(n8574), .A2(n4862), .ZN(n4513) );
  NAND2_X1 U5999 ( .A1(n5809), .A2(n5808), .ZN(n7017) );
  AND2_X1 U6000 ( .A1(n9142), .A2(n5039), .ZN(n4514) );
  NOR2_X1 U6001 ( .A1(n5668), .A2(n5020), .ZN(n5019) );
  NAND2_X1 U6002 ( .A1(n9326), .A2(n9210), .ZN(n4515) );
  AND2_X1 U6003 ( .A1(n5710), .A2(n5804), .ZN(n4516) );
  NAND2_X1 U6004 ( .A1(n9816), .A2(n9662), .ZN(n4517) );
  AND2_X1 U6005 ( .A1(n9222), .A2(n8441), .ZN(n4518) );
  NAND4_X1 U6006 ( .A1(n5880), .A2(n5879), .A3(n5878), .A4(n5877), .ZN(n6925)
         );
  AND2_X1 U6007 ( .A1(n5001), .A2(n4679), .ZN(n4519) );
  OR2_X1 U6008 ( .A1(n7833), .A2(n7834), .ZN(n4520) );
  OR2_X1 U6009 ( .A1(n8364), .A2(n4802), .ZN(n4521) );
  AND2_X1 U6010 ( .A1(n5776), .A2(n5781), .ZN(n5802) );
  INV_X1 U6011 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4836) );
  AND2_X1 U6012 ( .A1(n9838), .A2(n9752), .ZN(n4522) );
  AND2_X1 U6013 ( .A1(n8230), .A2(n8229), .ZN(n4523) );
  INV_X1 U6014 ( .A(n8461), .ZN(n8454) );
  NOR2_X1 U6015 ( .A1(n5862), .A2(n5861), .ZN(n5881) );
  NAND2_X1 U6016 ( .A1(n5587), .A2(n5586), .ZN(n9285) );
  NAND2_X1 U6017 ( .A1(n5351), .A2(n5350), .ZN(n7993) );
  OR3_X1 U6018 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .A3(
        P2_IR_REG_0__SCAN_IN), .ZN(n4524) );
  AND2_X1 U6019 ( .A1(n5056), .A2(n5088), .ZN(n4525) );
  AND2_X1 U6020 ( .A1(n5054), .A2(n5052), .ZN(n4526) );
  OAI211_X1 U6021 ( .C1(n4495), .C2(n4680), .A(n5000), .B(n5138), .ZN(n8627)
         );
  INV_X1 U6022 ( .A(n5813), .ZN(n5018) );
  NAND2_X1 U6023 ( .A1(n5002), .A2(n5095), .ZN(n5098) );
  NAND2_X1 U6024 ( .A1(n6196), .A2(n4716), .ZN(n5911) );
  OR2_X1 U6025 ( .A1(n6503), .A2(n4996), .ZN(n5890) );
  INV_X1 U6026 ( .A(n5002), .ZN(n5096) );
  NAND2_X1 U6027 ( .A1(n6322), .A2(n6321), .ZN(n9826) );
  NOR2_X1 U6028 ( .A1(n9401), .A2(n9396), .ZN(n4527) );
  OR2_X1 U6029 ( .A1(n5723), .A2(n5782), .ZN(n4528) );
  INV_X1 U6030 ( .A(n4735), .ZN(n9075) );
  NOR2_X1 U6031 ( .A1(n9091), .A2(n9291), .ZN(n4735) );
  OR2_X1 U6032 ( .A1(n8089), .A2(n8090), .ZN(n4529) );
  NOR2_X1 U6033 ( .A1(n4495), .A2(n7323), .ZN(n4530) );
  INV_X1 U6034 ( .A(n7737), .ZN(n4675) );
  INV_X1 U6035 ( .A(n9326), .ZN(n9188) );
  NAND2_X1 U6036 ( .A1(n5450), .A2(n5449), .ZN(n9326) );
  AND2_X1 U6037 ( .A1(n8211), .A2(n8412), .ZN(n9626) );
  INV_X1 U6038 ( .A(n9626), .ZN(n4749) );
  INV_X1 U6039 ( .A(n4946), .ZN(n4940) );
  NAND2_X1 U6040 ( .A1(n5301), .A2(n5288), .ZN(n4946) );
  NAND3_X1 U6041 ( .A1(n6282), .A2(n6264), .A3(n5883), .ZN(n4531) );
  AND2_X1 U6042 ( .A1(n7447), .A2(n7446), .ZN(n4532) );
  INV_X1 U6043 ( .A(n4845), .ZN(n9590) );
  NOR2_X1 U6044 ( .A1(n9607), .A2(n9789), .ZN(n4845) );
  AND2_X1 U6045 ( .A1(n6297), .A2(n6281), .ZN(n4533) );
  AND2_X1 U6046 ( .A1(n4520), .A2(n7907), .ZN(n4534) );
  AND2_X1 U6047 ( .A1(n5024), .A2(n4923), .ZN(n4535) );
  OR2_X1 U6048 ( .A1(n6780), .A2(n6861), .ZN(n4536) );
  INV_X1 U6049 ( .A(n8136), .ZN(n7894) );
  AND2_X1 U6050 ( .A1(n8194), .A2(n8393), .ZN(n8136) );
  INV_X1 U6051 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5111) );
  AND2_X1 U6052 ( .A1(n9956), .A2(n9520), .ZN(n4537) );
  AND2_X1 U6053 ( .A1(n4898), .A2(n9098), .ZN(n4538) );
  NOR2_X1 U6054 ( .A1(n6831), .A2(n5920), .ZN(n4539) );
  NOR2_X1 U6055 ( .A1(n9833), .A2(n9727), .ZN(n4540) );
  INV_X1 U6056 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5898) );
  OR2_X1 U6057 ( .A1(n9329), .A2(n9218), .ZN(n4541) );
  AND2_X1 U6058 ( .A1(n5815), .A2(n5671), .ZN(n4542) );
  AND2_X1 U6059 ( .A1(n9188), .A2(n8595), .ZN(n4543) );
  INV_X1 U6060 ( .A(n7298), .ZN(n4919) );
  OR2_X1 U6061 ( .A1(n6512), .A2(n6511), .ZN(n4544) );
  NOR2_X1 U6062 ( .A1(n9171), .A2(n8615), .ZN(n4545) );
  AND2_X1 U6063 ( .A1(n5718), .A2(n5720), .ZN(n7872) );
  INV_X1 U6064 ( .A(n7872), .ZN(n5024) );
  AND2_X1 U6065 ( .A1(n9142), .A2(n5756), .ZN(n4546) );
  AND2_X1 U6066 ( .A1(n5221), .A2(SI_6_), .ZN(n4547) );
  INV_X1 U6067 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5100) );
  INV_X1 U6068 ( .A(n4757), .ZN(n4756) );
  NAND2_X1 U6069 ( .A1(n4758), .A2(n8396), .ZN(n4757) );
  AND2_X1 U6070 ( .A1(n5303), .A2(SI_11_), .ZN(n4548) );
  NAND2_X1 U6071 ( .A1(n5897), .A2(n6539), .ZN(n4549) );
  NAND3_X1 U6072 ( .A1(n9082), .A2(n5764), .A3(n8448), .ZN(n4550) );
  AND2_X1 U6073 ( .A1(n6412), .A2(n6411), .ZN(n4551) );
  NAND2_X1 U6074 ( .A1(n9783), .A2(n9517), .ZN(n4552) );
  AND2_X1 U6075 ( .A1(n9536), .A2(n10109), .ZN(n4553) );
  AND2_X1 U6076 ( .A1(n4541), .A2(n4924), .ZN(n4554) );
  OR2_X1 U6077 ( .A1(n9335), .A2(n9241), .ZN(n5736) );
  AND2_X1 U6078 ( .A1(n5046), .A2(n5735), .ZN(n4555) );
  AND2_X1 U6079 ( .A1(n8461), .A2(n9038), .ZN(n4556) );
  AND2_X1 U6080 ( .A1(n9112), .A2(n9109), .ZN(n4557) );
  AND2_X1 U6081 ( .A1(n7539), .A2(n7538), .ZN(n4558) );
  AND2_X1 U6082 ( .A1(n4716), .A2(n5912), .ZN(n4559) );
  OR2_X1 U6083 ( .A1(n6780), .A2(n6647), .ZN(n4560) );
  AND2_X1 U6084 ( .A1(n4796), .A2(n9758), .ZN(n4561) );
  AND2_X1 U6085 ( .A1(n7474), .A2(n7473), .ZN(n4562) );
  OAI21_X1 U6086 ( .B1(n4913), .B2(n4910), .A(n7445), .ZN(n4909) );
  OR2_X1 U6087 ( .A1(n6503), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4563) );
  OR2_X1 U6088 ( .A1(n4499), .A2(n4505), .ZN(n4564) );
  INV_X1 U6089 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n4679) );
  INV_X1 U6090 ( .A(n4651), .ZN(n4650) );
  NAND2_X1 U6091 ( .A1(n4655), .A2(n8090), .ZN(n4651) );
  AND2_X1 U6092 ( .A1(n4811), .A2(n4809), .ZN(n4565) );
  INV_X1 U6093 ( .A(n8187), .ZN(n4745) );
  INV_X1 U6094 ( .A(n9460), .ZN(n4991) );
  NAND2_X1 U6095 ( .A1(n4814), .A2(n4813), .ZN(n7888) );
  NAND2_X1 U6096 ( .A1(n4981), .A2(n6135), .ZN(n7638) );
  NAND2_X1 U6097 ( .A1(n7741), .A2(n7740), .ZN(n7850) );
  NAND2_X1 U6098 ( .A1(n6176), .A2(n7765), .ZN(n7832) );
  AND4_X1 U6099 ( .A1(n5321), .A2(n5320), .A3(n5319), .A4(n5318), .ZN(n7873)
         );
  INV_X1 U6100 ( .A(n9783), .ZN(n4844) );
  NAND2_X1 U6101 ( .A1(n5737), .A2(n5734), .ZN(n7995) );
  NAND2_X1 U6102 ( .A1(n4907), .A2(n4669), .ZN(n10345) );
  NAND2_X1 U6103 ( .A1(n4907), .A2(n4906), .ZN(n10346) );
  AND2_X1 U6104 ( .A1(n9748), .A2(n8396), .ZN(n4566) );
  INV_X1 U6105 ( .A(n4974), .ZN(n4973) );
  NOR2_X1 U6106 ( .A1(n5386), .A2(n4975), .ZN(n4974) );
  NAND2_X1 U6107 ( .A1(n9203), .A2(n4726), .ZN(n4729) );
  NAND2_X1 U6108 ( .A1(n9761), .A2(n4852), .ZN(n4855) );
  NAND2_X1 U6109 ( .A1(n7859), .A2(n4722), .ZN(n4723) );
  OR2_X1 U6110 ( .A1(n6818), .A2(n7305), .ZN(n4567) );
  OR2_X1 U6111 ( .A1(n6820), .A2(n6819), .ZN(n4568) );
  OAI21_X1 U6112 ( .B1(n4869), .B2(n8345), .A(n4867), .ZN(n4866) );
  NAND2_X1 U6113 ( .A1(n4519), .A2(n5002), .ZN(n4569) );
  AND2_X1 U6114 ( .A1(n5486), .A2(n5479), .ZN(n4570) );
  INV_X1 U6115 ( .A(n10286), .ZN(n4871) );
  INV_X1 U6116 ( .A(n7992), .ZN(n4888) );
  INV_X1 U6117 ( .A(n7977), .ZN(n4875) );
  NAND2_X1 U6118 ( .A1(n6303), .A2(n6302), .ZN(n9833) );
  INV_X1 U6119 ( .A(n9833), .ZN(n4853) );
  INV_X1 U6120 ( .A(n4860), .ZN(n4862) );
  NAND2_X1 U6121 ( .A1(n4676), .A2(n5819), .ZN(n7738) );
  NOR2_X1 U6122 ( .A1(n7321), .A2(n10285), .ZN(n4571) );
  OR2_X1 U6123 ( .A1(n10357), .A2(n10436), .ZN(n4572) );
  NAND2_X1 U6124 ( .A1(n4918), .A2(n4915), .ZN(n7442) );
  NAND2_X1 U6125 ( .A1(n7509), .A2(n6106), .ZN(n7537) );
  INV_X1 U6126 ( .A(n9335), .ZN(n4721) );
  AND2_X1 U6127 ( .A1(n7295), .A2(n4919), .ZN(n4573) );
  AND2_X1 U6128 ( .A1(n7423), .A2(n7860), .ZN(n4574) );
  OR2_X1 U6129 ( .A1(n8614), .A2(n10260), .ZN(n4575) );
  AND2_X1 U6130 ( .A1(n5541), .A2(SI_24_), .ZN(n4576) );
  INV_X1 U6131 ( .A(n9853), .ZN(n4761) );
  INV_X1 U6132 ( .A(n8577), .ZN(n4858) );
  AND3_X1 U6133 ( .A1(n5173), .A2(n5172), .A3(n5171), .ZN(n10414) );
  INV_X1 U6134 ( .A(n10414), .ZN(n4785) );
  AND2_X1 U6135 ( .A1(n6612), .A2(n6611), .ZN(n10287) );
  AND2_X1 U6136 ( .A1(n10349), .A2(n10428), .ZN(n9926) );
  NAND2_X1 U6137 ( .A1(n6481), .A2(n4695), .ZN(n8107) );
  OR2_X1 U6138 ( .A1(n7375), .A2(n8117), .ZN(n7373) );
  NAND2_X1 U6139 ( .A1(n6935), .A2(n6937), .ZN(n6932) );
  AND2_X1 U6140 ( .A1(n6932), .A2(n6933), .ZN(n4577) );
  INV_X1 U6141 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5073) );
  INV_X1 U6142 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6264) );
  XNOR2_X1 U6143 ( .A(n5872), .B(n5871), .ZN(n8434) );
  AND3_X1 U6144 ( .A1(n4519), .A2(n5002), .A3(n4677), .ZN(n9368) );
  INV_X1 U6145 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n4680) );
  INV_X1 U6146 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n4600) );
  INV_X1 U6147 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n4979) );
  NAND2_X1 U6148 ( .A1(n4579), .A2(n4578), .ZN(P2_U3222) );
  NAND3_X1 U6149 ( .A1(n4580), .A2(n4868), .A3(n4863), .ZN(n4579) );
  INV_X1 U6150 ( .A(n8346), .ZN(n4581) );
  XNOR2_X2 U6151 ( .A(n8316), .B(n8317), .ZN(n8486) );
  AOI21_X2 U6152 ( .B1(n9097), .B2(n8448), .A(n5765), .ZN(n9081) );
  NAND2_X1 U6153 ( .A1(n4976), .A2(n5366), .ZN(n5387) );
  INV_X1 U6154 ( .A(n5046), .ZN(n5044) );
  INV_X1 U6155 ( .A(n5042), .ZN(n5041) );
  NOR2_X1 U6156 ( .A1(n5421), .A2(n5050), .ZN(n5049) );
  AND2_X4 U6157 ( .A1(n5874), .A2(n8434), .ZN(n8011) );
  NAND2_X1 U6158 ( .A1(n7790), .A2(n8154), .ZN(n9943) );
  NAND2_X1 U6159 ( .A1(n7085), .A2(n8237), .ZN(n8166) );
  OAI21_X2 U6160 ( .B1(n7723), .B2(n7722), .A(n8152), .ZN(n9967) );
  INV_X1 U6161 ( .A(n7895), .ZN(n4582) );
  NAND2_X1 U6162 ( .A1(n9706), .A2(n9705), .ZN(n9704) );
  OR2_X2 U6163 ( .A1(n9596), .A2(n9595), .ZN(n9600) );
  INV_X1 U6164 ( .A(n5393), .ZN(n5078) );
  OR2_X2 U6165 ( .A1(n9943), .A2(n4743), .ZN(n4740) );
  XNOR2_X1 U6166 ( .A(n8419), .B(n8418), .ZN(n4765) );
  MUX2_X1 U6167 ( .A(n5778), .B(n5777), .S(n5797), .Z(n5780) );
  NAND2_X1 U6168 ( .A1(n5407), .A2(n5406), .ZN(n5427) );
  NAND2_X1 U6169 ( .A1(n5186), .A2(n5187), .ZN(n4617) );
  INV_X1 U6170 ( .A(n5833), .ZN(n4629) );
  NAND2_X1 U6171 ( .A1(n5440), .A2(n5439), .ZN(n5443) );
  NAND2_X1 U6172 ( .A1(n5834), .A2(n4627), .ZN(n5842) );
  NAND2_X1 U6173 ( .A1(n4626), .A2(n5774), .ZN(n4624) );
  NAND2_X1 U6174 ( .A1(n4618), .A2(n8461), .ZN(n5783) );
  NAND2_X1 U6175 ( .A1(n5165), .A2(n5164), .ZN(n5186) );
  NAND2_X1 U6176 ( .A1(n4930), .A2(n4932), .ZN(n5230) );
  NAND2_X1 U6177 ( .A1(n4613), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n4612) );
  NAND2_X1 U6178 ( .A1(n5340), .A2(n5057), .ZN(n5342) );
  NAND2_X1 U6179 ( .A1(n5266), .A2(n5061), .ZN(n5268) );
  NAND2_X1 U6180 ( .A1(n4747), .A2(n4750), .ZN(n9596) );
  INV_X1 U6181 ( .A(n4744), .ZN(n4743) );
  AOI21_X2 U6182 ( .B1(n4765), .B2(n10172), .A(n4584), .ZN(n9780) );
  NAND2_X2 U6183 ( .A1(n9768), .A2(n9769), .ZN(n9767) );
  NAND2_X1 U6184 ( .A1(n4594), .A2(n4593), .ZN(n10022) );
  NAND2_X1 U6185 ( .A1(n6889), .A2(n6836), .ZN(n4594) );
  MUX2_X1 U6186 ( .A(n9896), .B(P1_IR_REG_0__SCAN_IN), .S(P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  MUX2_X1 U6187 ( .A(P1_IR_REG_0__SCAN_IN), .B(n9896), .S(n5963), .Z(n7369) );
  NAND3_X1 U6188 ( .A1(n10135), .A2(P1_IR_REG_0__SCAN_IN), .A3(n10019), .ZN(
        n10020) );
  NAND2_X1 U6189 ( .A1(n4612), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n4980) );
  AOI21_X1 U6190 ( .B1(n4616), .B2(n7873), .A(n5782), .ZN(n4614) );
  XNOR2_X1 U6191 ( .A(n5204), .B(n5202), .ZN(n6643) );
  NAND2_X1 U6192 ( .A1(n4621), .A2(n4619), .ZN(n4618) );
  OR2_X1 U6193 ( .A1(n4775), .A2(n4624), .ZN(n4621) );
  NAND2_X1 U6194 ( .A1(n4621), .A2(n4622), .ZN(n5787) );
  NOR2_X2 U6195 ( .A1(n5780), .A2(n5779), .ZN(n4626) );
  NAND2_X1 U6196 ( .A1(n4630), .A2(n4773), .ZN(n5748) );
  NAND2_X1 U6197 ( .A1(n5727), .A2(n4774), .ZN(n4630) );
  INV_X1 U6198 ( .A(n4632), .ZN(n4631) );
  OAI22_X1 U6199 ( .A1(n5724), .A2(n5797), .B1(n5726), .B2(n5725), .ZN(n4632)
         );
  NAND3_X1 U6200 ( .A1(n4641), .A2(n4778), .A3(n4777), .ZN(n4640) );
  NAND4_X1 U6201 ( .A1(n5745), .A2(n9144), .A3(n5782), .A4(n5750), .ZN(n4641)
         );
  OAI21_X1 U6202 ( .B1(n7376), .B2(n8117), .A(n4643), .ZN(n7379) );
  NAND2_X1 U6203 ( .A1(n7376), .A2(n8117), .ZN(n4643) );
  OAI21_X1 U6204 ( .B1(n8095), .B2(n4652), .A(n4651), .ZN(n8103) );
  OR2_X1 U6205 ( .A1(n4751), .A2(n8090), .ZN(n4654) );
  NAND3_X1 U6206 ( .A1(n4519), .A2(n5002), .A3(n5030), .ZN(n5101) );
  NAND2_X1 U6207 ( .A1(n8439), .A2(n4683), .ZN(n4682) );
  NAND2_X1 U6208 ( .A1(n5976), .A2(n6918), .ZN(n5980) );
  NAND3_X1 U6209 ( .A1(n6932), .A2(n6933), .A3(n6942), .ZN(n6918) );
  NAND2_X1 U6210 ( .A1(n4696), .A2(n4699), .ZN(n6156) );
  NAND3_X1 U6211 ( .A1(n7429), .A2(n4697), .A3(n7430), .ZN(n4696) );
  NAND3_X1 U6212 ( .A1(n7429), .A2(n7430), .A3(n7511), .ZN(n7509) );
  NAND2_X1 U6213 ( .A1(n6135), .A2(n4701), .ZN(n4700) );
  INV_X1 U6214 ( .A(n6106), .ZN(n4701) );
  NAND2_X1 U6215 ( .A1(n6391), .A2(n4564), .ZN(n4704) );
  INV_X1 U6216 ( .A(n6391), .ZN(n6394) );
  INV_X1 U6217 ( .A(n4710), .ZN(n9397) );
  INV_X1 U6218 ( .A(n4708), .ZN(n9422) );
  NAND3_X1 U6219 ( .A1(n9479), .A2(n9481), .A3(n6320), .ZN(n4713) );
  NAND2_X1 U6220 ( .A1(n6196), .A2(n4559), .ZN(n4715) );
  NAND2_X1 U6221 ( .A1(n6176), .A2(n4998), .ZN(n4718) );
  NAND2_X1 U6222 ( .A1(n4718), .A2(n4520), .ZN(n6214) );
  NAND2_X1 U6223 ( .A1(n8580), .A2(n4719), .ZN(n7157) );
  INV_X1 U6224 ( .A(n4723), .ZN(n9251) );
  INV_X1 U6225 ( .A(n4729), .ZN(n9154) );
  INV_X1 U6226 ( .A(n10357), .ZN(n4731) );
  XNOR2_X2 U6227 ( .A(n4738), .B(n5111), .ZN(n9385) );
  NAND3_X2 U6228 ( .A1(n4739), .A2(n5060), .A3(n5964), .ZN(n7386) );
  OR2_X1 U6229 ( .A1(n6013), .A2(n6632), .ZN(n4739) );
  NAND2_X2 U6230 ( .A1(n6524), .A2(n8271), .ZN(n5963) );
  NAND2_X1 U6231 ( .A1(n4740), .A2(n4741), .ZN(n7895) );
  NAND2_X1 U6232 ( .A1(n9625), .A2(n4748), .ZN(n4747) );
  AND2_X2 U6233 ( .A1(n5094), .A2(n5093), .ZN(n5002) );
  NAND2_X1 U6234 ( .A1(n5727), .A2(n4770), .ZN(n4767) );
  NAND2_X1 U6235 ( .A1(n4767), .A2(n4768), .ZN(n5752) );
  OAI21_X1 U6236 ( .B1(n4772), .B2(n4774), .A(n5747), .ZN(n4771) );
  NAND2_X1 U6237 ( .A1(n4773), .A2(n5746), .ZN(n4772) );
  OR2_X1 U6238 ( .A1(n5741), .A2(n5742), .ZN(n4773) );
  NAND3_X1 U6239 ( .A1(n4776), .A2(n5761), .A3(n9112), .ZN(n4775) );
  NAND2_X1 U6240 ( .A1(n4782), .A2(n4781), .ZN(n4780) );
  NAND2_X1 U6241 ( .A1(n4783), .A2(n5792), .ZN(n4782) );
  NAND2_X1 U6242 ( .A1(n5785), .A2(n4784), .ZN(n4783) );
  OR2_X1 U6243 ( .A1(n5787), .A2(n5786), .ZN(n4784) );
  NAND3_X1 U6244 ( .A1(n4787), .A2(n5158), .A3(n5159), .ZN(n8624) );
  NAND3_X1 U6245 ( .A1(n5695), .A2(n5701), .A3(n4792), .ZN(n4791) );
  NAND3_X1 U6246 ( .A1(n4794), .A2(n4793), .A3(n7872), .ZN(n5725) );
  NOR2_X1 U6247 ( .A1(n9368), .A2(n9369), .ZN(n4795) );
  NAND2_X1 U6248 ( .A1(n6228), .A2(n9531), .ZN(n5966) );
  OAI21_X1 U6249 ( .B1(n7891), .B2(n4521), .A(n4799), .ZN(n9759) );
  NAND2_X1 U6250 ( .A1(n4797), .A2(n4561), .ZN(n8367) );
  NAND2_X1 U6251 ( .A1(n7891), .A2(n4799), .ZN(n4797) );
  NAND2_X1 U6252 ( .A1(n8386), .A2(n4806), .ZN(n4803) );
  NAND2_X1 U6253 ( .A1(n4803), .A2(n4804), .ZN(n8388) );
  NAND2_X1 U6254 ( .A1(n8386), .A2(n9595), .ZN(n4811) );
  NAND2_X1 U6255 ( .A1(n4812), .A2(n4562), .ZN(n7718) );
  NAND2_X1 U6256 ( .A1(n7720), .A2(n4815), .ZN(n4814) );
  AND2_X1 U6257 ( .A1(n7393), .A2(n7201), .ZN(n7202) );
  NAND2_X1 U6258 ( .A1(n4818), .A2(n7199), .ZN(n7393) );
  AND2_X1 U6259 ( .A1(n7200), .A2(n7198), .ZN(n4818) );
  NAND2_X1 U6260 ( .A1(n4820), .A2(n4819), .ZN(n8385) );
  NAND2_X1 U6261 ( .A1(n7521), .A2(n4821), .ZN(n7471) );
  NAND2_X1 U6262 ( .A1(n7522), .A2(n8125), .ZN(n7521) );
  INV_X1 U6263 ( .A(n8126), .ZN(n4823) );
  NAND2_X1 U6264 ( .A1(n4825), .A2(n4824), .ZN(n8379) );
  NAND2_X1 U6265 ( .A1(n4992), .A2(n4508), .ZN(n9881) );
  NAND3_X1 U6266 ( .A1(n4992), .A2(n4508), .A3(n4836), .ZN(n4835) );
  NAND2_X1 U6267 ( .A1(n7373), .A2(n6959), .ZN(n6960) );
  NOR2_X2 U6268 ( .A1(n7899), .A2(n9856), .ZN(n9760) );
  OR2_X2 U6269 ( .A1(n9938), .A2(n7917), .ZN(n7899) );
  NAND3_X2 U6270 ( .A1(n4839), .A2(n4506), .A3(n4837), .ZN(n6503) );
  NAND3_X1 U6271 ( .A1(n5866), .A2(n5927), .A3(n5888), .ZN(n4838) );
  NOR2_X2 U6272 ( .A1(n5862), .A2(n5926), .ZN(n4839) );
  OAI211_X2 U6273 ( .C1(n6013), .C2(n6635), .A(n4843), .B(n4842), .ZN(n7553)
         );
  OR2_X1 U6274 ( .A1(n5963), .A2(n6886), .ZN(n4842) );
  NAND2_X2 U6275 ( .A1(n5963), .A2(n4583), .ZN(n5992) );
  NOR2_X2 U6276 ( .A1(n9634), .A2(n9799), .ZN(n9619) );
  INV_X1 U6277 ( .A(n7400), .ZN(n4847) );
  NAND3_X1 U6278 ( .A1(n4847), .A2(n10227), .A3(n4846), .ZN(n10160) );
  NAND2_X1 U6279 ( .A1(n9761), .A2(n4850), .ZN(n9699) );
  INV_X1 U6280 ( .A(n4855), .ZN(n9719) );
  NAND2_X1 U6281 ( .A1(n8346), .A2(n4864), .ZN(n4863) );
  INV_X1 U6282 ( .A(n8345), .ZN(n4872) );
  OAI21_X1 U6283 ( .B1(n7975), .B2(n4876), .A(n4873), .ZN(n8291) );
  NAND2_X1 U6284 ( .A1(n7962), .A2(n7961), .ZN(n7964) );
  NAND2_X1 U6285 ( .A1(n5074), .A2(n4885), .ZN(n5393) );
  NAND2_X1 U6286 ( .A1(n7653), .A2(n7652), .ZN(n7655) );
  NAND2_X1 U6287 ( .A1(n8551), .A2(n8303), .ZN(n8304) );
  OR2_X2 U6288 ( .A1(n5844), .A2(n10404), .ZN(n8314) );
  NAND2_X1 U6289 ( .A1(n9037), .A2(n4556), .ZN(n4890) );
  NAND3_X1 U6290 ( .A1(n4891), .A2(n4890), .A3(n4892), .ZN(n9279) );
  NAND3_X1 U6291 ( .A1(n4891), .A2(n4890), .A3(n4889), .ZN(n4897) );
  NAND2_X1 U6292 ( .A1(n4897), .A2(n9278), .ZN(n9352) );
  OAI21_X1 U6293 ( .B1(n9121), .B2(n4903), .A(n4899), .ZN(n9089) );
  NAND2_X1 U6294 ( .A1(n7297), .A2(n4905), .ZN(n4907) );
  NOR2_X1 U6295 ( .A1(n4512), .A2(n4909), .ZN(n4906) );
  AOI21_X1 U6296 ( .B1(n7295), .B2(n4917), .A(n4916), .ZN(n4915) );
  NAND2_X1 U6297 ( .A1(n7741), .A2(n4921), .ZN(n4920) );
  NAND2_X1 U6298 ( .A1(n4929), .A2(n5140), .ZN(n5120) );
  NAND2_X1 U6299 ( .A1(n5117), .A2(n5116), .ZN(n4929) );
  XNOR2_X1 U6300 ( .A(n4929), .B(n5140), .ZN(n6632) );
  NAND2_X1 U6301 ( .A1(n5204), .A2(n4931), .ZN(n4930) );
  NAND2_X1 U6302 ( .A1(n5287), .A2(n4502), .ZN(n4935) );
  NAND2_X1 U6303 ( .A1(n4935), .A2(n4936), .ZN(n5340) );
  OAI21_X1 U6304 ( .B1(n5508), .B2(n5507), .A(n5506), .ZN(n5513) );
  OAI211_X1 U6305 ( .C1(n4960), .C2(n4959), .A(n4958), .B(n4963), .ZN(P1_U3240) );
  AOI21_X1 U6306 ( .B1(n8145), .B2(n8144), .A(n8229), .ZN(n4961) );
  NAND2_X1 U6307 ( .A1(n8233), .A2(n8145), .ZN(n4962) );
  NAND2_X1 U6308 ( .A1(n4966), .A2(n4570), .ZN(n5490) );
  NAND3_X1 U6309 ( .A1(n6023), .A2(n6026), .A3(n6027), .ZN(n7051) );
  NAND2_X1 U6310 ( .A1(n7051), .A2(n6027), .ZN(n7132) );
  NAND2_X1 U6311 ( .A1(n6023), .A2(n6027), .ZN(n7050) );
  NAND2_X1 U6312 ( .A1(n9442), .A2(n6281), .ZN(n6300) );
  NAND2_X1 U6313 ( .A1(n9482), .A2(n9480), .ZN(n9479) );
  INV_X1 U6314 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n4997) );
  NAND2_X1 U6315 ( .A1(n5227), .A2(n4503), .ZN(n5005) );
  AOI21_X1 U6316 ( .B1(n4503), .B2(n5698), .A(n5004), .ZN(n5003) );
  INV_X1 U6317 ( .A(n5814), .ZN(n5020) );
  OAI21_X1 U6318 ( .B1(n7752), .B2(n5026), .A(n5023), .ZN(n7870) );
  OAI21_X1 U6319 ( .B1(n7752), .B2(n5714), .A(n5804), .ZN(n7742) );
  NAND2_X1 U6320 ( .A1(n5714), .A2(n5804), .ZN(n5029) );
  NAND2_X1 U6321 ( .A1(n9158), .A2(n5035), .ZN(n5032) );
  NAND2_X1 U6322 ( .A1(n5032), .A2(n5033), .ZN(n9097) );
  NAND2_X1 U6323 ( .A1(n7988), .A2(n4555), .ZN(n5045) );
  NAND2_X1 U6324 ( .A1(n5048), .A2(n5735), .ZN(n5043) );
  AND2_X1 U6325 ( .A1(n7978), .A2(n7976), .ZN(n7972) );
  CLKBUF_X1 U6326 ( .A(n7952), .Z(n7942) );
  OR2_X1 U6327 ( .A1(n9572), .A2(n4565), .ZN(n9788) );
  NAND2_X1 U6328 ( .A1(n6374), .A2(n6373), .ZN(n9470) );
  INV_X1 U6329 ( .A(n6371), .ZN(n6374) );
  NAND2_X1 U6330 ( .A1(n9881), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5873) );
  AND2_X1 U6331 ( .A1(n9277), .A2(n9276), .ZN(n9278) );
  OR2_X1 U6332 ( .A1(n5644), .A2(n6855), .ZN(n5138) );
  NAND2_X1 U6333 ( .A1(n7017), .A2(n7016), .ZN(n7158) );
  AND2_X1 U6334 ( .A1(n5089), .A2(n5073), .ZN(n5056) );
  INV_X1 U6335 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n7715) );
  AND2_X1 U6336 ( .A1(n5341), .A2(n5329), .ZN(n5057) );
  AND2_X1 U6337 ( .A1(n9928), .A2(n8617), .ZN(n5058) );
  OR2_X1 U6338 ( .A1(n6003), .A2(n5941), .ZN(n5059) );
  OR2_X1 U6339 ( .A1(n5963), .A2(n6868), .ZN(n5060) );
  INV_X1 U6340 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7711) );
  INV_X1 U6341 ( .A(n5827), .ZN(n5646) );
  AND2_X1 U6342 ( .A1(n5267), .A2(n5256), .ZN(n5061) );
  AND2_X1 U6343 ( .A1(n5288), .A2(n5273), .ZN(n5062) );
  INV_X1 U6344 ( .A(n7859), .ZN(n7880) );
  AND2_X1 U6345 ( .A1(n5612), .A2(n5611), .ZN(n8342) );
  AND3_X1 U6346 ( .A1(n5504), .A2(n5503), .A3(n5502), .ZN(n8567) );
  INV_X1 U6347 ( .A(n9280), .ZN(n8347) );
  OR2_X1 U6348 ( .A1(n9811), .A2(n9677), .ZN(n5063) );
  OR2_X1 U6349 ( .A1(n9128), .A2(n8545), .ZN(n5064) );
  OR2_X1 U6350 ( .A1(n9564), .A2(n9563), .ZN(P1_U3260) );
  INV_X1 U6351 ( .A(n8604), .ZN(n9114) );
  AND2_X1 U6352 ( .A1(n5557), .A2(n5556), .ZN(n8604) );
  NAND2_X1 U6353 ( .A1(n6064), .A2(n6063), .ZN(n5066) );
  OR2_X1 U6354 ( .A1(n9796), .A2(n9627), .ZN(n5067) );
  INV_X1 U6355 ( .A(n8266), .ZN(n6968) );
  INV_X2 U6356 ( .A(n9953), .ZN(n10181) );
  OR2_X1 U6357 ( .A1(n6962), .A2(n8266), .ZN(n7361) );
  INV_X1 U6358 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5088) );
  INV_X1 U6359 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n5866) );
  OAI21_X1 U6360 ( .B1(n9273), .B2(n5645), .A(n5789), .ZN(n5638) );
  INV_X1 U6361 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6362 ( .A1(n7386), .A2(n6478), .ZN(n5965) );
  INV_X1 U6363 ( .A(n7053), .ZN(n6026) );
  AOI21_X1 U6364 ( .B1(n6228), .B2(n7369), .A(n5948), .ZN(n5949) );
  INV_X1 U6365 ( .A(n5869), .ZN(n5870) );
  INV_X1 U6366 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n5868) );
  INV_X1 U6367 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n6111) );
  INV_X1 U6368 ( .A(n5354), .ZN(n5352) );
  INV_X1 U6369 ( .A(n5518), .ZN(n5517) );
  OR2_X1 U6370 ( .A1(n5589), .A2(n5588), .ZN(n5604) );
  INV_X1 U6371 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5835) );
  NAND2_X1 U6372 ( .A1(n5907), .A2(n5906), .ZN(n5915) );
  NOR2_X1 U6373 ( .A1(n6270), .A2(n6269), .ZN(n6288) );
  AND2_X1 U6374 ( .A1(n6118), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6140) );
  INV_X1 U6375 ( .A(n8118), .ZN(n6967) );
  INV_X1 U6376 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5885) );
  INV_X1 U6377 ( .A(n5438), .ZN(n5439) );
  INV_X1 U6378 ( .A(SI_8_), .ZN(n8922) );
  NAND2_X1 U6379 ( .A1(n5352), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n5377) );
  INV_X1 U6380 ( .A(n5472), .ZN(n5471) );
  NAND2_X1 U6381 ( .A1(n5517), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n5531) );
  OR2_X1 U6382 ( .A1(n5500), .A2(n5499), .ZN(n5518) );
  OR2_X1 U6383 ( .A1(n5569), .A2(n5568), .ZN(n5589) );
  INV_X1 U6384 ( .A(SI_19_), .ZN(n8913) );
  AND2_X1 U6385 ( .A1(n5604), .A2(n5590), .ZN(n9060) );
  INV_X1 U6386 ( .A(n8567), .ZN(n8444) );
  NOR2_X1 U6387 ( .A1(n5280), .A2(n5279), .ZN(n5295) );
  AND2_X1 U6388 ( .A1(n5209), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5244) );
  NAND2_X1 U6389 ( .A1(n7269), .A2(n7261), .ZN(n7260) );
  INV_X1 U6390 ( .A(n5802), .ZN(n9038) );
  OR2_X1 U6391 ( .A1(n5200), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5222) );
  INV_X1 U6392 ( .A(n6379), .ZN(n6398) );
  INV_X1 U6393 ( .A(n7177), .ZN(n6065) );
  OR2_X1 U6394 ( .A1(n8144), .A2(n6516), .ZN(n6517) );
  INV_X1 U6395 ( .A(n6372), .ZN(n6373) );
  INV_X1 U6396 ( .A(n6972), .ZN(n8144) );
  NAND2_X1 U6397 ( .A1(n6304), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n6324) );
  INV_X1 U6398 ( .A(n5874), .ZN(n5876) );
  AND2_X1 U6399 ( .A1(n6491), .A2(n6649), .ZN(n7354) );
  OR2_X1 U6400 ( .A1(n6162), .A2(n7768), .ZN(n6184) );
  OR2_X1 U6401 ( .A1(n6074), .A2(n7435), .ZN(n6092) );
  AND2_X1 U6402 ( .A1(n8129), .A2(n8128), .ZN(n10166) );
  NAND2_X1 U6403 ( .A1(n5307), .A2(n5306), .ZN(n5323) );
  INV_X1 U6404 ( .A(n7607), .ZN(n7608) );
  NAND2_X1 U6405 ( .A1(n5471), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5500) );
  INV_X1 U6406 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n5314) );
  AND3_X1 U6407 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_5__SCAN_IN), 
        .A3(P2_REG3_REG_3__SCAN_IN), .ZN(n5193) );
  OR2_X1 U6408 ( .A1(n5531), .A2(n5530), .ZN(n5550) );
  XNOR2_X1 U6409 ( .A(n6549), .B(n8578), .ZN(n8505) );
  NOR2_X1 U6410 ( .A1(n9310), .A2(n8444), .ZN(n8445) );
  AND2_X1 U6411 ( .A1(n5193), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5209) );
  NAND2_X1 U6412 ( .A1(n7214), .A2(n8427), .ZN(n9256) );
  INV_X1 U6413 ( .A(n8355), .ZN(n6615) );
  AND2_X1 U6414 ( .A1(n5689), .A2(n5686), .ZN(n10375) );
  INV_X1 U6415 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5083) );
  NAND2_X1 U6416 ( .A1(n9501), .A2(n9503), .ZN(n9432) );
  AND2_X1 U6417 ( .A1(n6517), .A2(n8270), .ZN(n6880) );
  INV_X1 U6418 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7513) );
  INV_X1 U6419 ( .A(n9495), .ZN(n9505) );
  AND2_X1 U6420 ( .A1(n6522), .A2(n6521), .ZN(n9510) );
  NOR2_X1 U6421 ( .A1(n6344), .A2(n6343), .ZN(n6360) );
  OR2_X1 U6422 ( .A1(n6236), .A2(n9436), .ZN(n6270) );
  INV_X1 U6423 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7435) );
  INV_X1 U6424 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7768) );
  INV_X1 U6425 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7109) );
  INV_X1 U6426 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9436) );
  AND2_X1 U6427 ( .A1(n8273), .A2(n6483), .ZN(n6972) );
  NAND2_X1 U6428 ( .A1(n7202), .A2(n8036), .ZN(n7468) );
  INV_X1 U6429 ( .A(n10226), .ZN(n9849) );
  INV_X1 U6430 ( .A(n10172), .ZN(n9949) );
  OR2_X1 U6431 ( .A1(n6962), .A2(n6968), .ZN(n10228) );
  AND2_X1 U6432 ( .A1(n7361), .A2(n6484), .ZN(n10226) );
  AND2_X1 U6433 ( .A1(n5406), .A2(n5392), .ZN(n5404) );
  NOR2_X1 U6434 ( .A1(n6622), .A2(n6621), .ZN(n10279) );
  AND2_X1 U6435 ( .A1(n6617), .A2(n8430), .ZN(n10286) );
  AND4_X1 U6436 ( .A1(n5403), .A2(n5402), .A3(n5401), .A4(n5400), .ZN(n8440)
         );
  AND2_X1 U6437 ( .A1(n6782), .A2(n6781), .ZN(n10336) );
  INV_X1 U6438 ( .A(n10295), .ZN(n10332) );
  AND2_X1 U6439 ( .A1(n9236), .A2(n9239), .ZN(n9339) );
  NAND2_X1 U6440 ( .A1(n7218), .A2(n9256), .ZN(n7864) );
  AND2_X1 U6441 ( .A1(n5845), .A2(n6623), .ZN(n10366) );
  AND2_X1 U6442 ( .A1(n7213), .A2(n7012), .ZN(n7013) );
  OR2_X1 U6443 ( .A1(n6615), .A2(n6614), .ZN(n10428) );
  AND2_X1 U6444 ( .A1(n7213), .A2(n7035), .ZN(n7036) );
  INV_X1 U6445 ( .A(n9926), .ZN(n10459) );
  AND2_X1 U6446 ( .A1(n6532), .A2(n6971), .ZN(n9495) );
  AND2_X1 U6447 ( .A1(n9455), .A2(n9849), .ZN(n9512) );
  OR2_X1 U6448 ( .A1(n6526), .A2(n9582), .ZN(n6471) );
  INV_X1 U6449 ( .A(n10142), .ZN(n10058) );
  NOR2_X1 U6450 ( .A1(n6702), .A2(n8359), .ZN(n10135) );
  AND2_X1 U6451 ( .A1(n9554), .A2(n6715), .ZN(n10148) );
  OR2_X1 U6452 ( .A1(n7357), .A2(n7356), .ZN(n7478) );
  INV_X1 U6453 ( .A(n10228), .ZN(n9984) );
  AND2_X1 U6454 ( .A1(n10175), .A2(n9862), .ZN(n9853) );
  INV_X1 U6455 ( .A(n9880), .ZN(n7355) );
  OAI211_X1 U6456 ( .C1(P1_B_REG_SCAN_IN), .C2(n7778), .A(n6488), .B(n6487), 
        .ZN(n6648) );
  AND2_X1 U6457 ( .A1(n6088), .A2(n6071), .ZN(n10051) );
  INV_X1 U6458 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n8859) );
  INV_X1 U6459 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n8810) );
  OR2_X1 U6460 ( .A1(n5853), .A2(n7799), .ZN(n6767) );
  INV_X1 U6461 ( .A(n10287), .ZN(n10246) );
  INV_X1 U6462 ( .A(n8342), .ZN(n9065) );
  INV_X1 U6463 ( .A(n8595), .ZN(n9210) );
  INV_X1 U6464 ( .A(n7873), .ZN(n8619) );
  INV_X1 U6465 ( .A(n7301), .ZN(n8623) );
  INV_X1 U6466 ( .A(n10336), .ZN(n10294) );
  AND2_X1 U6467 ( .A1(n7457), .A2(n7456), .ZN(n10443) );
  AND2_X1 U6468 ( .A1(n10360), .A2(n7229), .ZN(n9233) );
  NAND2_X1 U6469 ( .A1(n7212), .A2(n7013), .ZN(n10471) );
  AND4_X1 U6470 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .ZN(
        n10470) );
  NAND2_X1 U6471 ( .A1(n7212), .A2(n7036), .ZN(n10461) );
  NOR2_X1 U6472 ( .A1(n10385), .A2(n10384), .ZN(n10395) );
  INV_X1 U6473 ( .A(n10395), .ZN(n10398) );
  INV_X1 U6474 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6951) );
  OR2_X1 U6475 ( .A1(n6539), .A2(n7713), .ZN(n6717) );
  INV_X1 U6476 ( .A(n9512), .ZN(n9492) );
  OR3_X1 U6477 ( .A1(n6459), .A2(n6458), .A3(n6457), .ZN(n9576) );
  CLKBUF_X1 U6478 ( .A(P1_U4006), .Z(n9527) );
  INV_X1 U6479 ( .A(n10135), .ZN(n10154) );
  OR2_X1 U6480 ( .A1(P1_U3083), .A2(n6718), .ZN(n10157) );
  NAND2_X1 U6481 ( .A1(n10181), .A2(n7390), .ZN(n9777) );
  AND2_X2 U6482 ( .A1(n6955), .A2(n9880), .ZN(n10245) );
  AND2_X1 U6483 ( .A1(n9990), .A2(n9989), .ZN(n10006) );
  AND2_X2 U6484 ( .A1(n6955), .A2(n7355), .ZN(n10236) );
  NAND2_X1 U6485 ( .A1(n8270), .A2(n6648), .ZN(n10193) );
  AND2_X1 U6486 ( .A1(n6490), .A2(n6489), .ZN(n9880) );
  INV_X1 U6487 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7777) );
  INV_X1 U6488 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8474) );
  INV_X1 U6489 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7045) );
  INV_X1 U6490 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6685) );
  NOR2_X1 U6491 ( .A1(n10514), .A2(n10513), .ZN(n10512) );
  NOR2_X1 U6492 ( .A1(n10501), .A2(n10500), .ZN(n10499) );
  AND2_X2 U6493 ( .A1(n5169), .A2(n4507), .ZN(n5094) );
  NAND2_X1 U6494 ( .A1(n5094), .A2(n5072), .ZN(n5274) );
  INV_X2 U6495 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5089) );
  INV_X1 U6496 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n5075) );
  INV_X1 U6497 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5343) );
  AND3_X1 U6498 ( .A1(n5075), .A2(n5347), .A3(n5343), .ZN(n5076) );
  INV_X1 U6499 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5079) );
  INV_X1 U6500 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5080) );
  NOR2_X1 U6501 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n5087) );
  NOR2_X1 U6502 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5086) );
  NOR2_X1 U6503 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n5085) );
  NOR2_X1 U6504 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n5084) );
  NAND4_X1 U6505 ( .A1(n5087), .A2(n5086), .A3(n5085), .A4(n5084), .ZN(n5092)
         );
  NAND4_X1 U6506 ( .A1(n5090), .A2(n5089), .A3(n5347), .A4(n5088), .ZN(n5091)
         );
  NOR2_X1 U6507 ( .A1(n5092), .A2(n5091), .ZN(n5093) );
  NAND2_X1 U6508 ( .A1(n5098), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5836) );
  NAND2_X1 U6509 ( .A1(n5096), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5097) );
  NAND2_X1 U6510 ( .A1(n6615), .A2(n6616), .ZN(n7024) );
  AND2_X2 U6511 ( .A1(n8353), .A2(n5103), .ZN(n5157) );
  INV_X1 U6512 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6773) );
  OR2_X1 U6513 ( .A1(n5573), .A2(n6773), .ZN(n5108) );
  NAND2_X1 U6514 ( .A1(n5640), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5107) );
  INV_X1 U6515 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6791) );
  OR2_X1 U6516 ( .A1(n5644), .A2(n6791), .ZN(n5106) );
  NAND2_X1 U6517 ( .A1(n5431), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5105) );
  XNOR2_X2 U6518 ( .A(n5110), .B(n5109), .ZN(n6797) );
  AND2_X1 U6519 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5113) );
  NAND2_X1 U6520 ( .A1(n5154), .A2(n5113), .ZN(n5946) );
  NAND3_X1 U6521 ( .A1(n5112), .A2(SI_0_), .A3(P1_DATAO_REG_0__SCAN_IN), .ZN(
        n5114) );
  NAND2_X1 U6522 ( .A1(n5946), .A2(n5114), .ZN(n5118) );
  INV_X1 U6523 ( .A(SI_1_), .ZN(n5115) );
  XNOR2_X1 U6524 ( .A(n5118), .B(n5115), .ZN(n5140) );
  OR2_X1 U6525 ( .A1(n5154), .A2(n6633), .ZN(n5117) );
  NAND2_X1 U6526 ( .A1(n4497), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n5116) );
  NAND2_X1 U6527 ( .A1(n5118), .A2(SI_1_), .ZN(n5119) );
  NAND2_X1 U6528 ( .A1(n5120), .A2(n5119), .ZN(n5149) );
  INV_X1 U6529 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6634) );
  INV_X1 U6530 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6630) );
  MUX2_X1 U6531 ( .A(n6634), .B(n6630), .S(n5154), .Z(n5150) );
  XNOR2_X1 U6532 ( .A(n5150), .B(SI_2_), .ZN(n5148) );
  XNOR2_X1 U6533 ( .A(n5149), .B(n5148), .ZN(n6635) );
  OR2_X1 U6534 ( .A1(n5185), .A2(n6635), .ZN(n5125) );
  NAND2_X4 U6535 ( .A1(n6780), .A2(n4497), .ZN(n5660) );
  OR2_X1 U6536 ( .A1(n5660), .A2(n6634), .ZN(n5124) );
  OR2_X1 U6537 ( .A1(n5121), .A2(n9369), .ZN(n5122) );
  XNOR2_X1 U6538 ( .A(n5122), .B(P2_IR_REG_2__SCAN_IN), .ZN(n9910) );
  INV_X1 U6539 ( .A(n9910), .ZN(n6636) );
  OR2_X1 U6540 ( .A1(n6780), .A2(n6636), .ZN(n5123) );
  AND2_X1 U6541 ( .A1(n8626), .A2(n10408), .ZN(n5673) );
  INV_X1 U6542 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n5126) );
  INV_X1 U6543 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6790) );
  OR2_X1 U6544 ( .A1(n5644), .A2(n6790), .ZN(n5129) );
  INV_X1 U6545 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5127) );
  NAND2_X1 U6546 ( .A1(n5129), .A2(n5128), .ZN(n5130) );
  NOR2_X1 U6547 ( .A1(n5131), .A2(n5130), .ZN(n5133) );
  INV_X1 U6548 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6771) );
  NAND2_X1 U6549 ( .A1(n4583), .A2(SI_0_), .ZN(n5134) );
  XNOR2_X1 U6550 ( .A(n5134), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9386) );
  MUX2_X1 U6551 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9386), .S(n6780), .Z(n8431) );
  INV_X1 U6552 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6855) );
  INV_X1 U6553 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5135) );
  OR2_X1 U6554 ( .A1(n5174), .A2(n5135), .ZN(n5137) );
  NAND2_X1 U6555 ( .A1(n5157), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5136) );
  INV_X1 U6556 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5139) );
  INV_X1 U6557 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6633) );
  OR2_X1 U6558 ( .A1(n5660), .A2(n6633), .ZN(n5142) );
  OR2_X1 U6559 ( .A1(n5185), .A2(n6632), .ZN(n5141) );
  NAND2_X1 U6560 ( .A1(n7029), .A2(n5809), .ZN(n7270) );
  INV_X1 U6561 ( .A(n10408), .ZN(n8576) );
  NAND2_X1 U6562 ( .A1(n5640), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5146) );
  OR2_X1 U6563 ( .A1(n4495), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5145) );
  INV_X1 U6564 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6789) );
  OR2_X1 U6565 ( .A1(n5644), .A2(n6789), .ZN(n5144) );
  INV_X1 U6566 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6770) );
  OR2_X1 U6567 ( .A1(n5573), .A2(n6770), .ZN(n5143) );
  NAND2_X1 U6568 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n4524), .ZN(n5147) );
  XNOR2_X1 U6569 ( .A(n5147), .B(P2_IR_REG_3__SCAN_IN), .ZN(n10306) );
  INV_X1 U6570 ( .A(n10306), .ZN(n6639) );
  NAND2_X1 U6571 ( .A1(n5149), .A2(n5148), .ZN(n5153) );
  INV_X1 U6572 ( .A(n5150), .ZN(n5151) );
  NAND2_X1 U6573 ( .A1(n5151), .A2(SI_2_), .ZN(n5152) );
  NAND2_X1 U6574 ( .A1(n5153), .A2(n5152), .ZN(n5161) );
  INV_X1 U6575 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6637) );
  INV_X1 U6576 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6631) );
  XNOR2_X1 U6577 ( .A(n5161), .B(n5160), .ZN(n6638) );
  OR2_X1 U6578 ( .A1(n5185), .A2(n6638), .ZN(n5156) );
  OR2_X1 U6579 ( .A1(n5660), .A2(n6637), .ZN(n5155) );
  NAND2_X1 U6580 ( .A1(n7314), .A2(n7169), .ZN(n5671) );
  INV_X1 U6581 ( .A(n7314), .ZN(n8625) );
  INV_X1 U6582 ( .A(n7169), .ZN(n10250) );
  NAND2_X1 U6583 ( .A1(n8625), .A2(n10250), .ZN(n5682) );
  NAND2_X1 U6584 ( .A1(n7163), .A2(n7164), .ZN(n7162) );
  NAND2_X1 U6585 ( .A1(n7162), .A2(n5671), .ZN(n7311) );
  NAND2_X1 U6586 ( .A1(n5606), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5159) );
  NAND2_X1 U6587 ( .A1(n5640), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5158) );
  XNOR2_X1 U6588 ( .A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n7323) );
  INV_X1 U6589 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6777) );
  NAND2_X1 U6590 ( .A1(n5161), .A2(n5160), .ZN(n5165) );
  INV_X1 U6591 ( .A(n5162), .ZN(n5163) );
  NAND2_X1 U6592 ( .A1(n5163), .A2(SI_3_), .ZN(n5164) );
  INV_X1 U6593 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6641) );
  INV_X1 U6594 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n6640) );
  MUX2_X1 U6595 ( .A(n6641), .B(n6640), .S(n4497), .Z(n5188) );
  XNOR2_X1 U6596 ( .A(n5188), .B(SI_4_), .ZN(n5187) );
  XNOR2_X1 U6597 ( .A(n5186), .B(n5187), .ZN(n6642) );
  OR2_X1 U6598 ( .A1(n5185), .A2(n6642), .ZN(n5173) );
  OR2_X1 U6599 ( .A1(n5660), .A2(n6641), .ZN(n5172) );
  NOR2_X1 U6600 ( .A1(n5169), .A2(n9369), .ZN(n5166) );
  MUX2_X1 U6601 ( .A(n9369), .B(n5166), .S(P2_IR_REG_4__SCAN_IN), .Z(n5167) );
  INV_X1 U6602 ( .A(n5167), .ZN(n5170) );
  INV_X1 U6603 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5168) );
  NAND2_X1 U6604 ( .A1(n5169), .A2(n5168), .ZN(n5200) );
  NAND2_X1 U6605 ( .A1(n5170), .A2(n5200), .ZN(n6848) );
  OR2_X1 U6606 ( .A1(n6780), .A2(n6848), .ZN(n5171) );
  NAND2_X1 U6607 ( .A1(n8624), .A2(n10414), .ZN(n5814) );
  INV_X1 U6608 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7235) );
  OR2_X1 U6609 ( .A1(n5644), .A2(n7235), .ZN(n5183) );
  INV_X1 U6610 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6769) );
  OR2_X1 U6611 ( .A1(n5573), .A2(n6769), .ZN(n5182) );
  INV_X1 U6612 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n5175) );
  OR2_X1 U6613 ( .A1(n5174), .A2(n5175), .ZN(n5181) );
  INV_X1 U6614 ( .A(n5193), .ZN(n5179) );
  INV_X1 U6615 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6616 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n5176) );
  NAND2_X1 U6617 ( .A1(n5177), .A2(n5176), .ZN(n5178) );
  NAND2_X1 U6618 ( .A1(n5179), .A2(n5178), .ZN(n10291) );
  OR2_X1 U6619 ( .A1(n4496), .A2(n10291), .ZN(n5180) );
  INV_X1 U6620 ( .A(n7313), .ZN(n10367) );
  NAND2_X1 U6621 ( .A1(n5200), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5184) );
  XNOR2_X1 U6622 ( .A(n5184), .B(P2_IR_REG_5__SCAN_IN), .ZN(n9900) );
  INV_X1 U6623 ( .A(n9900), .ZN(n6647) );
  INV_X1 U6624 ( .A(n5188), .ZN(n5189) );
  NAND2_X1 U6625 ( .A1(n5189), .A2(SI_4_), .ZN(n5190) );
  MUX2_X1 U6626 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n8007), .Z(n5205) );
  XNOR2_X1 U6627 ( .A(n5205), .B(SI_5_), .ZN(n5202) );
  NAND2_X1 U6628 ( .A1(n5658), .A2(n6643), .ZN(n5192) );
  INV_X1 U6629 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6645) );
  OR2_X1 U6630 ( .A1(n5660), .A2(n6645), .ZN(n5191) );
  NAND2_X1 U6631 ( .A1(n7313), .A2(n10285), .ZN(n5813) );
  NAND2_X1 U6632 ( .A1(n5640), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5199) );
  NOR2_X1 U6633 ( .A1(n5193), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5194) );
  NOR2_X1 U6634 ( .A1(n5209), .A2(n5194), .ZN(n10374) );
  INV_X1 U6635 ( .A(n10374), .ZN(n7190) );
  OR2_X1 U6636 ( .A1(n4496), .A2(n7190), .ZN(n5198) );
  INV_X1 U6637 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5195) );
  OR2_X1 U6638 ( .A1(n5644), .A2(n5195), .ZN(n5197) );
  INV_X1 U6639 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6779) );
  OR2_X1 U6640 ( .A1(n5573), .A2(n6779), .ZN(n5196) );
  NAND2_X1 U6641 ( .A1(n5222), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5201) );
  XNOR2_X1 U6642 ( .A(n5201), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6815) );
  AOI22_X1 U6643 ( .A1(n5448), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n5447), .B2(
        n6815), .ZN(n5208) );
  INV_X1 U6644 ( .A(n5202), .ZN(n5203) );
  NAND2_X1 U6645 ( .A1(n5205), .A2(SI_5_), .ZN(n5206) );
  MUX2_X1 U6646 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n8007), .Z(n5221) );
  XNOR2_X1 U6647 ( .A(n5220), .B(n5218), .ZN(n6652) );
  NAND2_X1 U6648 ( .A1(n6652), .A2(n5658), .ZN(n5207) );
  NAND2_X1 U6649 ( .A1(n5208), .A2(n5207), .ZN(n7302) );
  NAND2_X1 U6650 ( .A1(n7301), .A2(n7302), .ZN(n5689) );
  INV_X1 U6651 ( .A(n7302), .ZN(n10379) );
  NAND2_X1 U6652 ( .A1(n8623), .A2(n10379), .ZN(n5686) );
  NAND2_X1 U6653 ( .A1(n10364), .A2(n5689), .ZN(n7299) );
  NAND2_X1 U6654 ( .A1(n5640), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5217) );
  INV_X1 U6655 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n7305) );
  OR2_X1 U6656 ( .A1(n5644), .A2(n7305), .ZN(n5216) );
  INV_X1 U6657 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6805) );
  OR2_X1 U6658 ( .A1(n5573), .A2(n6805), .ZN(n5215) );
  INV_X1 U6659 ( .A(n5244), .ZN(n5213) );
  INV_X1 U6660 ( .A(n5209), .ZN(n5211) );
  INV_X1 U6661 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U6662 ( .A1(n5211), .A2(n5210), .ZN(n5212) );
  NAND2_X1 U6663 ( .A1(n5213), .A2(n5212), .ZN(n7304) );
  OR2_X1 U6664 ( .A1(n4495), .A2(n7304), .ZN(n5214) );
  INV_X1 U6665 ( .A(n5218), .ZN(n5219) );
  MUX2_X1 U6666 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n4497), .Z(n5231) );
  XNOR2_X1 U6667 ( .A(n5231), .B(SI_7_), .ZN(n5228) );
  XNOR2_X1 U6668 ( .A(n5230), .B(n5228), .ZN(n6659) );
  NAND2_X1 U6669 ( .A1(n6659), .A2(n5658), .ZN(n5226) );
  INV_X1 U6670 ( .A(n5222), .ZN(n5223) );
  NAND2_X1 U6671 ( .A1(n5223), .A2(n8924), .ZN(n5237) );
  NAND2_X1 U6672 ( .A1(n5237), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5224) );
  XNOR2_X1 U6673 ( .A(n5224), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10316) );
  AOI22_X1 U6674 ( .A1(n5448), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n5447), .B2(
        n10316), .ZN(n5225) );
  NAND2_X1 U6675 ( .A1(n5226), .A2(n5225), .ZN(n7458) );
  AND2_X1 U6676 ( .A1(n7444), .A2(n7458), .ZN(n5688) );
  INV_X1 U6677 ( .A(n7458), .ZN(n7443) );
  INV_X1 U6678 ( .A(n7444), .ZN(n10369) );
  NAND2_X1 U6679 ( .A1(n7443), .A2(n10369), .ZN(n5691) );
  INV_X1 U6680 ( .A(n5228), .ZN(n5229) );
  NAND2_X1 U6681 ( .A1(n5230), .A2(n5229), .ZN(n5233) );
  NAND2_X1 U6682 ( .A1(n5231), .A2(SI_7_), .ZN(n5232) );
  MUX2_X1 U6683 ( .A(n6663), .B(n6665), .S(n8007), .Z(n5234) );
  NAND2_X1 U6684 ( .A1(n5234), .A2(n8922), .ZN(n5251) );
  INV_X1 U6685 ( .A(n5234), .ZN(n5235) );
  NAND2_X1 U6686 ( .A1(n5235), .A2(SI_8_), .ZN(n5236) );
  NAND2_X1 U6687 ( .A1(n5251), .A2(n5236), .ZN(n5249) );
  XNOR2_X1 U6688 ( .A(n5250), .B(n5249), .ZN(n6662) );
  NAND2_X1 U6689 ( .A1(n6662), .A2(n5658), .ZN(n5242) );
  OAI21_X1 U6690 ( .B1(n5237), .B2(P2_IR_REG_7__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n5238) );
  MUX2_X1 U6691 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5238), .S(
        P2_IR_REG_8__SCAN_IN), .Z(n5240) );
  INV_X1 U6692 ( .A(n5094), .ZN(n5239) );
  AOI22_X1 U6693 ( .A1(n5448), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n5447), .B2(
        n8634), .ZN(n5241) );
  NAND2_X1 U6694 ( .A1(n5242), .A2(n5241), .ZN(n10356) );
  NAND2_X1 U6695 ( .A1(n5606), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5248) );
  INV_X1 U6696 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n5243) );
  OR2_X1 U6697 ( .A1(n5174), .A2(n5243), .ZN(n5247) );
  OAI21_X1 U6698 ( .B1(n5244), .B2(P2_REG3_REG_8__SCAN_IN), .A(n5280), .ZN(
        n10353) );
  OR2_X1 U6699 ( .A1(n4496), .A2(n10353), .ZN(n5246) );
  INV_X1 U6700 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6804) );
  OR2_X1 U6701 ( .A1(n5573), .A2(n6804), .ZN(n5245) );
  XNOR2_X1 U6702 ( .A(n10356), .B(n7453), .ZN(n10343) );
  NAND2_X1 U6703 ( .A1(n10356), .A2(n7453), .ZN(n5696) );
  INV_X1 U6704 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n5252) );
  MUX2_X1 U6705 ( .A(n5252), .B(n8761), .S(n4497), .Z(n5254) );
  INV_X1 U6706 ( .A(SI_9_), .ZN(n5253) );
  NAND2_X1 U6707 ( .A1(n5254), .A2(n5253), .ZN(n5267) );
  INV_X1 U6708 ( .A(n5254), .ZN(n5255) );
  NAND2_X1 U6709 ( .A1(n5255), .A2(SI_9_), .ZN(n5256) );
  XNOR2_X1 U6710 ( .A(n5266), .B(n5061), .ZN(n6666) );
  NAND2_X1 U6711 ( .A1(n6666), .A2(n5658), .ZN(n5259) );
  OR2_X1 U6712 ( .A1(n5094), .A2(n9369), .ZN(n5257) );
  XNOR2_X1 U6713 ( .A(n5257), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6992) );
  AOI22_X1 U6714 ( .A1(n5448), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n5447), .B2(
        n6992), .ZN(n5258) );
  NAND2_X1 U6715 ( .A1(n5259), .A2(n5258), .ZN(n10436) );
  INV_X1 U6716 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n5260) );
  OR2_X1 U6717 ( .A1(n5174), .A2(n5260), .ZN(n5265) );
  INV_X1 U6718 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7461) );
  OR2_X1 U6719 ( .A1(n5644), .A2(n7461), .ZN(n5264) );
  INV_X1 U6720 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5261) );
  XNOR2_X1 U6721 ( .A(n5280), .B(n5261), .ZN(n7460) );
  OR2_X1 U6722 ( .A1(n4496), .A2(n7460), .ZN(n5263) );
  INV_X1 U6723 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6808) );
  OR2_X1 U6724 ( .A1(n5573), .A2(n6808), .ZN(n5262) );
  OR2_X1 U6725 ( .A1(n10436), .A2(n7501), .ZN(n5700) );
  NAND2_X1 U6726 ( .A1(n10436), .A2(n7501), .ZN(n5701) );
  MUX2_X1 U6727 ( .A(n5269), .B(n6685), .S(n8007), .Z(n5271) );
  INV_X1 U6728 ( .A(SI_10_), .ZN(n5270) );
  NAND2_X1 U6729 ( .A1(n5271), .A2(n5270), .ZN(n5288) );
  INV_X1 U6730 ( .A(n5271), .ZN(n5272) );
  NAND2_X1 U6731 ( .A1(n5272), .A2(SI_10_), .ZN(n5273) );
  XNOR2_X1 U6732 ( .A(n5287), .B(n5062), .ZN(n6680) );
  NAND2_X1 U6733 ( .A1(n6680), .A2(n5658), .ZN(n5276) );
  NAND2_X1 U6734 ( .A1(n5274), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5289) );
  XNOR2_X1 U6735 ( .A(n5289), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10329) );
  AOI22_X1 U6736 ( .A1(n5448), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n5447), .B2(
        n10329), .ZN(n5275) );
  NAND2_X1 U6737 ( .A1(n5276), .A2(n5275), .ZN(n10445) );
  NAND2_X1 U6738 ( .A1(n5157), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5285) );
  INV_X1 U6739 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n5277) );
  OR2_X1 U6740 ( .A1(n5174), .A2(n5277), .ZN(n5284) );
  INV_X1 U6741 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n6991) );
  OR2_X1 U6742 ( .A1(n5644), .A2(n6991), .ZN(n5283) );
  INV_X1 U6743 ( .A(n5280), .ZN(n5278) );
  AOI21_X1 U6744 ( .B1(n5278), .B2(P2_REG3_REG_9__SCAN_IN), .A(
        P2_REG3_REG_10__SCAN_IN), .ZN(n5281) );
  NAND2_X1 U6745 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_REG3_REG_9__SCAN_IN), 
        .ZN(n5279) );
  OR2_X1 U6746 ( .A1(n5281), .A2(n5295), .ZN(n7610) );
  OR2_X1 U6747 ( .A1(n4496), .A2(n7610), .ZN(n5282) );
  OR2_X1 U6748 ( .A1(n10445), .A2(n7736), .ZN(n5706) );
  NAND2_X1 U6749 ( .A1(n10445), .A2(n7736), .ZN(n5705) );
  NAND2_X1 U6750 ( .A1(n7495), .A2(n7504), .ZN(n5286) );
  NAND2_X1 U6751 ( .A1(n5286), .A2(n5705), .ZN(n7752) );
  MUX2_X1 U6752 ( .A(n6686), .B(n6683), .S(n8007), .Z(n5302) );
  XNOR2_X1 U6753 ( .A(n5302), .B(SI_11_), .ZN(n5301) );
  XNOR2_X1 U6754 ( .A(n5304), .B(n5301), .ZN(n6682) );
  NAND2_X1 U6755 ( .A1(n6682), .A2(n5658), .ZN(n5293) );
  NAND2_X1 U6756 ( .A1(n5289), .A2(n5089), .ZN(n5290) );
  NAND2_X1 U6757 ( .A1(n5290), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5291) );
  XNOR2_X1 U6758 ( .A(n5291), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7061) );
  AOI22_X1 U6759 ( .A1(n5448), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n5447), .B2(
        n7061), .ZN(n5292) );
  NAND2_X1 U6760 ( .A1(n5640), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5300) );
  INV_X1 U6761 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n5294) );
  OR2_X1 U6762 ( .A1(n5644), .A2(n5294), .ZN(n5299) );
  NAND2_X1 U6763 ( .A1(n5295), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5315) );
  OR2_X1 U6764 ( .A1(n5295), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5296) );
  NAND2_X1 U6765 ( .A1(n5315), .A2(n5296), .ZN(n7658) );
  OR2_X1 U6766 ( .A1(n4495), .A2(n7658), .ZN(n5298) );
  INV_X1 U6767 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7001) );
  OR2_X1 U6768 ( .A1(n5573), .A2(n7001), .ZN(n5297) );
  AND2_X1 U6769 ( .A1(n7758), .A2(n7744), .ZN(n5714) );
  OR2_X1 U6770 ( .A1(n7758), .A2(n7744), .ZN(n5804) );
  INV_X1 U6771 ( .A(n5302), .ZN(n5303) );
  MUX2_X1 U6772 ( .A(n6863), .B(n5305), .S(n8007), .Z(n5307) );
  INV_X1 U6773 ( .A(SI_12_), .ZN(n5306) );
  INV_X1 U6774 ( .A(n5307), .ZN(n5308) );
  NAND2_X1 U6775 ( .A1(n5308), .A2(SI_12_), .ZN(n5309) );
  NAND2_X1 U6776 ( .A1(n5323), .A2(n5309), .ZN(n5324) );
  XNOR2_X1 U6777 ( .A(n5325), .B(n5324), .ZN(n6825) );
  NAND2_X1 U6778 ( .A1(n6825), .A2(n5658), .ZN(n5313) );
  NAND2_X1 U6779 ( .A1(n5310), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5311) );
  XNOR2_X1 U6780 ( .A(n5311), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7075) );
  AOI22_X1 U6781 ( .A1(n5448), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n5447), .B2(
        n7075), .ZN(n5312) );
  NAND2_X1 U6782 ( .A1(n5606), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5321) );
  NAND2_X1 U6783 ( .A1(n5315), .A2(n5314), .ZN(n5316) );
  NAND2_X1 U6784 ( .A1(n5333), .A2(n5316), .ZN(n10276) );
  OR2_X1 U6785 ( .A1(n4495), .A2(n10276), .ZN(n5320) );
  INV_X1 U6786 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n7069) );
  OR2_X1 U6787 ( .A1(n5573), .A2(n7069), .ZN(n5319) );
  INV_X1 U6788 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n5317) );
  OR2_X1 U6789 ( .A1(n5174), .A2(n5317), .ZN(n5318) );
  NAND2_X1 U6790 ( .A1(n10274), .A2(n7873), .ZN(n5712) );
  INV_X1 U6791 ( .A(n5710), .ZN(n5322) );
  MUX2_X1 U6792 ( .A(n6951), .B(n6949), .S(n8007), .Z(n5327) );
  INV_X1 U6793 ( .A(SI_13_), .ZN(n5326) );
  INV_X1 U6794 ( .A(n5327), .ZN(n5328) );
  NAND2_X1 U6795 ( .A1(n5328), .A2(SI_13_), .ZN(n5329) );
  XNOR2_X1 U6796 ( .A(n5340), .B(n5057), .ZN(n6948) );
  NAND2_X1 U6797 ( .A1(n6948), .A2(n5658), .ZN(n5332) );
  OR2_X1 U6798 ( .A1(n5330), .A2(n9369), .ZN(n5344) );
  XNOR2_X1 U6799 ( .A(n5344), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7338) );
  AOI22_X1 U6800 ( .A1(n5448), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n5447), .B2(
        n7338), .ZN(n5331) );
  NAND2_X1 U6801 ( .A1(n5640), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5339) );
  INV_X1 U6802 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7883) );
  OR2_X1 U6803 ( .A1(n5644), .A2(n7883), .ZN(n5338) );
  NAND2_X1 U6804 ( .A1(n5333), .A2(n7827), .ZN(n5334) );
  NAND2_X1 U6805 ( .A1(n5354), .A2(n5334), .ZN(n7882) );
  OR2_X1 U6806 ( .A1(n4496), .A2(n7882), .ZN(n5337) );
  INV_X1 U6807 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n5335) );
  OR2_X1 U6808 ( .A1(n5573), .A2(n5335), .ZN(n5336) );
  OR2_X1 U6809 ( .A1(n7932), .A2(n10261), .ZN(n5718) );
  NAND2_X1 U6810 ( .A1(n7932), .A2(n10261), .ZN(n5720) );
  NAND2_X1 U6811 ( .A1(n7870), .A2(n5720), .ZN(n7852) );
  MUX2_X1 U6812 ( .A(n6980), .B(n6954), .S(n8007), .Z(n5364) );
  XNOR2_X1 U6813 ( .A(n5364), .B(SI_14_), .ZN(n5361) );
  XNOR2_X1 U6814 ( .A(n5363), .B(n5361), .ZN(n6953) );
  NAND2_X1 U6815 ( .A1(n6953), .A2(n5658), .ZN(n5351) );
  NAND2_X1 U6816 ( .A1(n5344), .A2(n5343), .ZN(n5345) );
  NAND2_X1 U6817 ( .A1(n5345), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5348) );
  INV_X1 U6818 ( .A(n5348), .ZN(n5346) );
  NAND2_X1 U6819 ( .A1(n5346), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n5349) );
  NAND2_X1 U6820 ( .A1(n5348), .A2(n5347), .ZN(n5371) );
  AOI22_X1 U6821 ( .A1(n5448), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n5447), .B2(
        n7351), .ZN(n5350) );
  NAND2_X1 U6822 ( .A1(n5640), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5360) );
  INV_X1 U6823 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7860) );
  OR2_X1 U6824 ( .A1(n5644), .A2(n7860), .ZN(n5359) );
  INV_X1 U6825 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6826 ( .A1(n5354), .A2(n5353), .ZN(n5355) );
  NAND2_X1 U6827 ( .A1(n5377), .A2(n5355), .ZN(n7949) );
  OR2_X1 U6828 ( .A1(n4496), .A2(n7949), .ZN(n5358) );
  INV_X1 U6829 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n5356) );
  OR2_X1 U6830 ( .A1(n5573), .A2(n5356), .ZN(n5357) );
  XNOR2_X1 U6831 ( .A(n7993), .B(n7965), .ZN(n7992) );
  NOR2_X1 U6832 ( .A1(n7852), .A2(n7992), .ZN(n7855) );
  INV_X1 U6833 ( .A(n7993), .ZN(n9928) );
  INV_X1 U6834 ( .A(n7965), .ZN(n8617) );
  INV_X1 U6835 ( .A(n5361), .ZN(n5362) );
  INV_X1 U6836 ( .A(n5364), .ZN(n5365) );
  NAND2_X1 U6837 ( .A1(n5365), .A2(SI_14_), .ZN(n5366) );
  MUX2_X1 U6838 ( .A(n7046), .B(n7045), .S(n8007), .Z(n5368) );
  INV_X1 U6839 ( .A(SI_15_), .ZN(n5367) );
  NAND2_X1 U6840 ( .A1(n5368), .A2(n5367), .ZN(n5385) );
  INV_X1 U6841 ( .A(n5368), .ZN(n5369) );
  NAND2_X1 U6842 ( .A1(n5369), .A2(SI_15_), .ZN(n5370) );
  NAND2_X1 U6843 ( .A1(n5385), .A2(n5370), .ZN(n5386) );
  XNOR2_X1 U6844 ( .A(n5387), .B(n5386), .ZN(n7044) );
  NAND2_X1 U6845 ( .A1(n7044), .A2(n5658), .ZN(n5374) );
  NAND2_X1 U6846 ( .A1(n5371), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5372) );
  XNOR2_X1 U6847 ( .A(n5372), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7625) );
  AOI22_X1 U6848 ( .A1(n5448), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n5447), .B2(
        n7625), .ZN(n5373) );
  NAND2_X1 U6849 ( .A1(n5640), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5384) );
  INV_X1 U6850 ( .A(n5377), .ZN(n5375) );
  NAND2_X1 U6851 ( .A1(n5375), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n5398) );
  INV_X1 U6852 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5376) );
  NAND2_X1 U6853 ( .A1(n5377), .A2(n5376), .ZN(n5378) );
  NAND2_X1 U6854 ( .A1(n5398), .A2(n5378), .ZN(n7998) );
  OR2_X1 U6855 ( .A1(n4495), .A2(n7998), .ZN(n5383) );
  INV_X1 U6856 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n5379) );
  OR2_X1 U6857 ( .A1(n5644), .A2(n5379), .ZN(n5382) );
  INV_X1 U6858 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n5380) );
  OR2_X1 U6859 ( .A1(n5573), .A2(n5380), .ZN(n5381) );
  NAND2_X1 U6860 ( .A1(n9346), .A2(n9243), .ZN(n5734) );
  INV_X1 U6861 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n5388) );
  MUX2_X1 U6862 ( .A(n7048), .B(n5388), .S(n8007), .Z(n5390) );
  INV_X1 U6863 ( .A(SI_16_), .ZN(n5389) );
  NAND2_X1 U6864 ( .A1(n5390), .A2(n5389), .ZN(n5406) );
  INV_X1 U6865 ( .A(n5390), .ZN(n5391) );
  NAND2_X1 U6866 ( .A1(n5391), .A2(SI_16_), .ZN(n5392) );
  XNOR2_X1 U6867 ( .A(n5405), .B(n5404), .ZN(n7042) );
  NAND2_X1 U6868 ( .A1(n7042), .A2(n5658), .ZN(n5396) );
  NAND2_X1 U6869 ( .A1(n5393), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5394) );
  XNOR2_X1 U6870 ( .A(n5394), .B(P2_IR_REG_16__SCAN_IN), .ZN(n7667) );
  AOI22_X1 U6871 ( .A1(n5448), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n5447), .B2(
        n7667), .ZN(n5395) );
  NAND2_X1 U6872 ( .A1(n5640), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5403) );
  INV_X1 U6873 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n9258) );
  OR2_X1 U6874 ( .A1(n5644), .A2(n9258), .ZN(n5402) );
  INV_X1 U6875 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n5397) );
  NAND2_X1 U6876 ( .A1(n5398), .A2(n5397), .ZN(n5399) );
  NAND2_X1 U6877 ( .A1(n5415), .A2(n5399), .ZN(n9257) );
  OR2_X1 U6878 ( .A1(n4496), .A2(n9257), .ZN(n5401) );
  INV_X1 U6879 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7616) );
  OR2_X1 U6880 ( .A1(n5573), .A2(n7616), .ZN(n5400) );
  OR2_X1 U6881 ( .A1(n9340), .A2(n8440), .ZN(n5728) );
  NAND2_X1 U6882 ( .A1(n9340), .A2(n8440), .ZN(n9215) );
  NAND2_X1 U6883 ( .A1(n5728), .A2(n9215), .ZN(n9245) );
  INV_X1 U6884 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n5408) );
  MUX2_X1 U6885 ( .A(n7098), .B(n5408), .S(n4497), .Z(n5423) );
  XNOR2_X1 U6886 ( .A(n5423), .B(SI_17_), .ZN(n5422) );
  XNOR2_X1 U6887 ( .A(n5427), .B(n5422), .ZN(n7078) );
  NAND2_X1 U6888 ( .A1(n7078), .A2(n5658), .ZN(n5412) );
  NAND2_X1 U6889 ( .A1(n5409), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5410) );
  XNOR2_X1 U6890 ( .A(n5410), .B(P2_IR_REG_17__SCAN_IN), .ZN(n7673) );
  AOI22_X1 U6891 ( .A1(n5448), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n5447), .B2(
        n7673), .ZN(n5411) );
  INV_X1 U6892 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n8985) );
  OR2_X1 U6893 ( .A1(n5174), .A2(n8985), .ZN(n5420) );
  INV_X1 U6894 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9226) );
  OR2_X1 U6895 ( .A1(n5644), .A2(n9226), .ZN(n5419) );
  INV_X1 U6896 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5414) );
  NAND2_X1 U6897 ( .A1(n5415), .A2(n5414), .ZN(n5416) );
  NAND2_X1 U6898 ( .A1(n5457), .A2(n5416), .ZN(n9225) );
  OR2_X1 U6899 ( .A1(n4496), .A2(n9225), .ZN(n5418) );
  INV_X1 U6900 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8647) );
  OR2_X1 U6901 ( .A1(n5573), .A2(n8647), .ZN(n5417) );
  NAND2_X1 U6902 ( .A1(n9335), .A2(n9241), .ZN(n5733) );
  NAND2_X1 U6903 ( .A1(n5803), .A2(n9215), .ZN(n5421) );
  INV_X1 U6904 ( .A(n5422), .ZN(n5426) );
  INV_X1 U6905 ( .A(n5423), .ZN(n5424) );
  NAND2_X1 U6906 ( .A1(n5424), .A2(SI_17_), .ZN(n5425) );
  MUX2_X1 U6907 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n8007), .Z(n5441) );
  XNOR2_X1 U6908 ( .A(n5441), .B(SI_18_), .ZN(n5438) );
  XNOR2_X1 U6909 ( .A(n5440), .B(n5438), .ZN(n7257) );
  NAND2_X1 U6910 ( .A1(n7257), .A2(n5658), .ZN(n5430) );
  XNOR2_X1 U6911 ( .A(n5428), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8657) );
  AOI22_X1 U6912 ( .A1(n5448), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n5447), .B2(
        n8657), .ZN(n5429) );
  XNOR2_X1 U6913 ( .A(n5457), .B(P2_REG3_REG_18__SCAN_IN), .ZN(n9204) );
  NAND2_X1 U6914 ( .A1(n9204), .A2(n5431), .ZN(n5437) );
  INV_X1 U6915 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n5432) );
  OR2_X1 U6916 ( .A1(n5174), .A2(n5432), .ZN(n5436) );
  INV_X1 U6917 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n5433) );
  OR2_X1 U6918 ( .A1(n5644), .A2(n5433), .ZN(n5435) );
  INV_X1 U6919 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n8648) );
  OR2_X1 U6920 ( .A1(n5573), .A2(n8648), .ZN(n5434) );
  NOR2_X1 U6921 ( .A1(n9329), .A2(n8531), .ZN(n5743) );
  NAND2_X1 U6922 ( .A1(n9329), .A2(n8531), .ZN(n5746) );
  NAND2_X1 U6923 ( .A1(n5441), .A2(SI_18_), .ZN(n5442) );
  MUX2_X1 U6924 ( .A(n7287), .B(n7286), .S(n4497), .Z(n5444) );
  NAND2_X1 U6925 ( .A1(n5444), .A2(n8913), .ZN(n5462) );
  INV_X1 U6926 ( .A(n5444), .ZN(n5445) );
  NAND2_X1 U6927 ( .A1(n5445), .A2(SI_19_), .ZN(n5446) );
  NAND2_X1 U6928 ( .A1(n5462), .A2(n5446), .ZN(n5463) );
  XNOR2_X1 U6929 ( .A(n5464), .B(n5463), .ZN(n7285) );
  NAND2_X1 U6930 ( .A1(n7285), .A2(n5658), .ZN(n5450) );
  AOI22_X1 U6931 ( .A1(n5448), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9194), .B2(
        n5447), .ZN(n5449) );
  INV_X1 U6932 ( .A(P2_REG0_REG_19__SCAN_IN), .ZN(n5451) );
  OR2_X1 U6933 ( .A1(n5174), .A2(n5451), .ZN(n5453) );
  INV_X1 U6934 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9198) );
  OR2_X1 U6935 ( .A1(n5644), .A2(n9198), .ZN(n5452) );
  AND2_X1 U6936 ( .A1(n5453), .A2(n5452), .ZN(n5461) );
  INV_X1 U6937 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n5455) );
  INV_X1 U6938 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5454) );
  OAI21_X1 U6939 ( .B1(n5457), .B2(n5455), .A(n5454), .ZN(n5458) );
  NAND2_X1 U6940 ( .A1(P2_REG3_REG_19__SCAN_IN), .A2(P2_REG3_REG_18__SCAN_IN), 
        .ZN(n5456) );
  AND2_X1 U6941 ( .A1(n5458), .A2(n5472), .ZN(n9196) );
  NAND2_X1 U6942 ( .A1(n9196), .A2(n5431), .ZN(n5460) );
  NAND2_X1 U6943 ( .A1(n5157), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5459) );
  OR2_X1 U6944 ( .A1(n9326), .A2(n8595), .ZN(n5747) );
  NAND2_X1 U6945 ( .A1(n9326), .A2(n8595), .ZN(n5749) );
  NAND2_X1 U6946 ( .A1(n9184), .A2(n9185), .ZN(n9183) );
  NAND2_X1 U6947 ( .A1(n9183), .A2(n5749), .ZN(n9173) );
  OAI21_X2 U6948 ( .B1(n5464), .B2(n5463), .A(n5462), .ZN(n5478) );
  MUX2_X1 U6949 ( .A(n8813), .B(n8898), .S(n4497), .Z(n5466) );
  INV_X1 U6950 ( .A(SI_20_), .ZN(n5465) );
  NAND2_X1 U6951 ( .A1(n5466), .A2(n5465), .ZN(n5479) );
  INV_X1 U6952 ( .A(n5466), .ZN(n5467) );
  NAND2_X1 U6953 ( .A1(n5467), .A2(SI_20_), .ZN(n5468) );
  XNOR2_X1 U6954 ( .A(n5478), .B(n5477), .ZN(n7408) );
  NAND2_X1 U6955 ( .A1(n7408), .A2(n5658), .ZN(n5470) );
  OR2_X1 U6956 ( .A1(n5660), .A2(n8813), .ZN(n5469) );
  INV_X1 U6957 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8811) );
  NAND2_X1 U6958 ( .A1(n5472), .A2(n8811), .ZN(n5473) );
  NAND2_X1 U6959 ( .A1(n5500), .A2(n5473), .ZN(n8553) );
  OR2_X1 U6960 ( .A1(n8553), .A2(n4496), .ZN(n5476) );
  AOI22_X1 U6961 ( .A1(n5606), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n5640), .B2(
        P2_REG0_REG_20__SCAN_IN), .ZN(n5475) );
  INV_X1 U6962 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n8933) );
  OR2_X1 U6963 ( .A1(n5573), .A2(n8933), .ZN(n5474) );
  OR2_X1 U6964 ( .A1(n9321), .A2(n8615), .ZN(n5751) );
  NAND2_X1 U6965 ( .A1(n9321), .A2(n8615), .ZN(n5750) );
  NAND2_X1 U6966 ( .A1(n9173), .A2(n9174), .ZN(n9172) );
  NAND2_X1 U6967 ( .A1(n9172), .A2(n5750), .ZN(n9159) );
  MUX2_X1 U6968 ( .A(n7518), .B(n8749), .S(n4497), .Z(n5487) );
  XNOR2_X1 U6969 ( .A(n5487), .B(SI_21_), .ZN(n5486) );
  XNOR2_X1 U6970 ( .A(n5485), .B(n5486), .ZN(n7508) );
  NAND2_X1 U6971 ( .A1(n7508), .A2(n5658), .ZN(n5481) );
  OR2_X1 U6972 ( .A1(n5660), .A2(n7518), .ZN(n5480) );
  XNOR2_X1 U6973 ( .A(n5500), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n9155) );
  INV_X1 U6974 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n8894) );
  NAND2_X1 U6975 ( .A1(n5640), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U6976 ( .A1(n5606), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5482) );
  OAI211_X1 U6977 ( .C1(n8894), .C2(n5573), .A(n5483), .B(n5482), .ZN(n5484)
         );
  AOI21_X1 U6978 ( .B1(n9155), .B2(n5431), .A(n5484), .ZN(n8558) );
  OR2_X1 U6979 ( .A1(n9315), .A2(n8558), .ZN(n5755) );
  NAND2_X1 U6980 ( .A1(n9315), .A2(n8558), .ZN(n9144) );
  NAND2_X1 U6981 ( .A1(n9159), .A2(n9160), .ZN(n9158) );
  INV_X1 U6982 ( .A(n5487), .ZN(n5488) );
  NAND2_X1 U6983 ( .A1(n5488), .A2(SI_21_), .ZN(n5489) );
  MUX2_X1 U6984 ( .A(n7636), .B(n8474), .S(n8007), .Z(n5492) );
  INV_X1 U6985 ( .A(SI_22_), .ZN(n5491) );
  NAND2_X1 U6986 ( .A1(n5492), .A2(n5491), .ZN(n5506) );
  INV_X1 U6987 ( .A(n5492), .ZN(n5493) );
  NAND2_X1 U6988 ( .A1(n5493), .A2(SI_22_), .ZN(n5494) );
  NAND2_X1 U6989 ( .A1(n5506), .A2(n5494), .ZN(n5507) );
  XNOR2_X1 U6990 ( .A(n5508), .B(n5507), .ZN(n7635) );
  NAND2_X1 U6991 ( .A1(n7635), .A2(n5658), .ZN(n5496) );
  OR2_X1 U6992 ( .A1(n5660), .A2(n7636), .ZN(n5495) );
  INV_X1 U6993 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5498) );
  INV_X1 U6994 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n5497) );
  OAI21_X1 U6995 ( .B1(n5500), .B2(n5498), .A(n5497), .ZN(n5501) );
  NAND2_X1 U6996 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n5499) );
  NAND2_X1 U6997 ( .A1(n5501), .A2(n5518), .ZN(n9138) );
  OR2_X1 U6998 ( .A1(n9138), .A2(n4495), .ZN(n5504) );
  AOI22_X1 U6999 ( .A1(n5606), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n5640), .B2(
        P2_REG0_REG_22__SCAN_IN), .ZN(n5503) );
  INV_X1 U7000 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n8873) );
  OR2_X1 U7001 ( .A1(n5573), .A2(n8873), .ZN(n5502) );
  NAND2_X1 U7002 ( .A1(n9310), .A2(n8567), .ZN(n5757) );
  MUX2_X1 U7003 ( .A(n7711), .B(n7715), .S(n8007), .Z(n5509) );
  INV_X1 U7004 ( .A(SI_23_), .ZN(n8833) );
  NAND2_X1 U7005 ( .A1(n5509), .A2(n8833), .ZN(n5526) );
  INV_X1 U7006 ( .A(n5509), .ZN(n5510) );
  NAND2_X1 U7007 ( .A1(n5510), .A2(SI_23_), .ZN(n5511) );
  OR2_X1 U7008 ( .A1(n5513), .A2(n5512), .ZN(n5514) );
  NAND2_X1 U7009 ( .A1(n5527), .A2(n5514), .ZN(n7712) );
  NAND2_X1 U7010 ( .A1(n7712), .A2(n5658), .ZN(n5516) );
  OR2_X1 U7011 ( .A1(n5660), .A2(n7711), .ZN(n5515) );
  INV_X1 U7012 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n8871) );
  NAND2_X1 U7013 ( .A1(n5518), .A2(n8871), .ZN(n5519) );
  NAND2_X1 U7014 ( .A1(n5531), .A2(n5519), .ZN(n9125) );
  OR2_X1 U7015 ( .A1(n9125), .A2(n4495), .ZN(n5525) );
  INV_X1 U7016 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n5522) );
  NAND2_X1 U7017 ( .A1(n5640), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n5521) );
  NAND2_X1 U7018 ( .A1(n5157), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n5520) );
  OAI211_X1 U7019 ( .C1(n5644), .C2(n5522), .A(n5521), .B(n5520), .ZN(n5523)
         );
  INV_X1 U7020 ( .A(n5523), .ZN(n5524) );
  NAND2_X1 U7021 ( .A1(n5525), .A2(n5524), .ZN(n9113) );
  NAND2_X1 U7022 ( .A1(n9128), .A2(n9113), .ZN(n5760) );
  INV_X1 U7023 ( .A(n9113), .ZN(n8545) );
  NAND2_X1 U7024 ( .A1(n9305), .A2(n8545), .ZN(n9109) );
  MUX2_X1 U7025 ( .A(n7797), .B(n7777), .S(n4497), .Z(n5540) );
  XNOR2_X1 U7026 ( .A(n5540), .B(SI_24_), .ZN(n5539) );
  XNOR2_X1 U7027 ( .A(n5542), .B(n5539), .ZN(n7776) );
  NAND2_X1 U7028 ( .A1(n7776), .A2(n5658), .ZN(n5529) );
  OR2_X1 U7029 ( .A1(n5660), .A2(n7797), .ZN(n5528) );
  INV_X1 U7030 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U7031 ( .A1(n5531), .A2(n5530), .ZN(n5532) );
  AND2_X1 U7032 ( .A1(n5550), .A2(n5532), .ZN(n9106) );
  NAND2_X1 U7033 ( .A1(n9106), .A2(n5431), .ZN(n5538) );
  INV_X1 U7034 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n5535) );
  NAND2_X1 U7035 ( .A1(n5640), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U7036 ( .A1(n5606), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n5533) );
  OAI211_X1 U7037 ( .C1(n5535), .C2(n5573), .A(n5534), .B(n5533), .ZN(n5536)
         );
  INV_X1 U7038 ( .A(n5536), .ZN(n5537) );
  NAND2_X1 U7039 ( .A1(n9300), .A2(n8540), .ZN(n5763) );
  AND2_X2 U7040 ( .A1(n5762), .A2(n5763), .ZN(n9112) );
  INV_X1 U7041 ( .A(n5540), .ZN(n5541) );
  INV_X1 U7042 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7921) );
  INV_X1 U7043 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n7925) );
  MUX2_X1 U7044 ( .A(n7921), .B(n7925), .S(n8007), .Z(n5544) );
  INV_X1 U7045 ( .A(SI_25_), .ZN(n5543) );
  NAND2_X1 U7046 ( .A1(n5544), .A2(n5543), .ZN(n5559) );
  INV_X1 U7047 ( .A(n5544), .ZN(n5545) );
  NAND2_X1 U7048 ( .A1(n5545), .A2(SI_25_), .ZN(n5546) );
  NAND2_X1 U7049 ( .A1(n5559), .A2(n5546), .ZN(n5560) );
  NAND2_X1 U7050 ( .A1(n7920), .A2(n5658), .ZN(n5548) );
  OR2_X1 U7051 ( .A1(n5660), .A2(n7921), .ZN(n5547) );
  INV_X1 U7052 ( .A(n5550), .ZN(n5549) );
  NAND2_X1 U7053 ( .A1(n5549), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n5569) );
  INV_X1 U7054 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8523) );
  NAND2_X1 U7055 ( .A1(n5550), .A2(n8523), .ZN(n5551) );
  NAND2_X1 U7056 ( .A1(n5569), .A2(n5551), .ZN(n9094) );
  OR2_X1 U7057 ( .A1(n9094), .A2(n4495), .ZN(n5557) );
  INV_X1 U7058 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n5554) );
  NAND2_X1 U7059 ( .A1(n5640), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U7060 ( .A1(n5606), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n5552) );
  OAI211_X1 U7061 ( .C1(n5554), .C2(n5573), .A(n5553), .B(n5552), .ZN(n5555)
         );
  INV_X1 U7062 ( .A(n5555), .ZN(n5556) );
  NAND2_X1 U7063 ( .A1(n9296), .A2(n8604), .ZN(n5768) );
  INV_X1 U7064 ( .A(n5558), .ZN(n5765) );
  INV_X1 U7065 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n7929) );
  INV_X1 U7066 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n7927) );
  MUX2_X1 U7067 ( .A(n7929), .B(n7927), .S(n8007), .Z(n5563) );
  INV_X1 U7068 ( .A(SI_26_), .ZN(n5562) );
  NAND2_X1 U7069 ( .A1(n5563), .A2(n5562), .ZN(n5580) );
  INV_X1 U7070 ( .A(n5563), .ZN(n5564) );
  NAND2_X1 U7071 ( .A1(n5564), .A2(SI_26_), .ZN(n5565) );
  XNOR2_X1 U7072 ( .A(n5579), .B(n5578), .ZN(n7926) );
  NAND2_X1 U7073 ( .A1(n7926), .A2(n5658), .ZN(n5567) );
  OR2_X1 U7074 ( .A1(n5660), .A2(n7929), .ZN(n5566) );
  INV_X1 U7075 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n5568) );
  NAND2_X1 U7076 ( .A1(n5569), .A2(n5568), .ZN(n5570) );
  NAND2_X1 U7077 ( .A1(n5589), .A2(n5570), .ZN(n9076) );
  OR2_X1 U7078 ( .A1(n9076), .A2(n4496), .ZN(n5577) );
  INV_X1 U7079 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n5574) );
  NAND2_X1 U7080 ( .A1(n5640), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5572) );
  NAND2_X1 U7081 ( .A1(n5606), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n5571) );
  OAI211_X1 U7082 ( .C1(n5574), .C2(n5573), .A(n5572), .B(n5571), .ZN(n5575)
         );
  INV_X1 U7083 ( .A(n5575), .ZN(n5576) );
  NAND2_X1 U7084 ( .A1(n9291), .A2(n8522), .ZN(n5767) );
  NAND2_X1 U7085 ( .A1(n9081), .A2(n9082), .ZN(n9080) );
  INV_X1 U7086 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9383) );
  INV_X1 U7087 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n9895) );
  MUX2_X1 U7088 ( .A(n9383), .B(n9895), .S(n4497), .Z(n5583) );
  INV_X1 U7089 ( .A(SI_27_), .ZN(n5582) );
  NAND2_X1 U7090 ( .A1(n5583), .A2(n5582), .ZN(n5599) );
  INV_X1 U7091 ( .A(n5583), .ZN(n5584) );
  NAND2_X1 U7092 ( .A1(n5584), .A2(SI_27_), .ZN(n5585) );
  XNOR2_X2 U7093 ( .A(n5598), .B(n5597), .ZN(n9893) );
  NAND2_X1 U7094 ( .A1(n9893), .A2(n5658), .ZN(n5587) );
  OR2_X1 U7095 ( .A1(n5660), .A2(n9383), .ZN(n5586) );
  INV_X1 U7096 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7097 ( .A1(n5589), .A2(n5588), .ZN(n5590) );
  NAND2_X1 U7098 ( .A1(n9060), .A2(n5431), .ZN(n5596) );
  INV_X1 U7099 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U7100 ( .A1(n5606), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n5592) );
  NAND2_X1 U7101 ( .A1(n5640), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n5591) );
  OAI211_X1 U7102 ( .C1(n5593), .C2(n5573), .A(n5592), .B(n5591), .ZN(n5594)
         );
  INV_X1 U7103 ( .A(n5594), .ZN(n5595) );
  INV_X1 U7104 ( .A(n9285), .ZN(n9062) );
  NAND2_X1 U7105 ( .A1(n9062), .A2(n9083), .ZN(n5775) );
  OAI21_X1 U7106 ( .B1(n9063), .B2(n9064), .A(n5775), .ZN(n9039) );
  INV_X1 U7107 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9381) );
  INV_X1 U7108 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9890) );
  MUX2_X1 U7109 ( .A(n9381), .B(n9890), .S(n8007), .Z(n5617) );
  XNOR2_X1 U7110 ( .A(n5617), .B(SI_28_), .ZN(n5614) );
  XNOR2_X2 U7111 ( .A(n5615), .B(n5614), .ZN(n9888) );
  NAND2_X1 U7112 ( .A1(n9888), .A2(n5658), .ZN(n5602) );
  OR2_X1 U7113 ( .A1(n5660), .A2(n9381), .ZN(n5601) );
  NAND2_X2 U7114 ( .A1(n5602), .A2(n5601), .ZN(n9280) );
  INV_X1 U7115 ( .A(n5604), .ZN(n5603) );
  NAND2_X1 U7116 ( .A1(n5603), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n5623) );
  INV_X1 U7117 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U7118 ( .A1(n5604), .A2(n8348), .ZN(n5605) );
  NAND2_X1 U7119 ( .A1(n5623), .A2(n5605), .ZN(n9047) );
  OR2_X1 U7120 ( .A1(n9047), .A2(n4495), .ZN(n5612) );
  INV_X1 U7121 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n5609) );
  NAND2_X1 U7122 ( .A1(n5640), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n5608) );
  NAND2_X1 U7123 ( .A1(n5606), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n5607) );
  OAI211_X1 U7124 ( .C1(n5609), .C2(n5573), .A(n5608), .B(n5607), .ZN(n5610)
         );
  INV_X1 U7125 ( .A(n5610), .ZN(n5611) );
  NAND2_X1 U7126 ( .A1(n9280), .A2(n8342), .ZN(n5781) );
  INV_X1 U7127 ( .A(n5776), .ZN(n5613) );
  INV_X1 U7128 ( .A(SI_28_), .ZN(n5616) );
  NAND2_X1 U7129 ( .A1(n5617), .A2(n5616), .ZN(n5618) );
  INV_X1 U7130 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n8472) );
  INV_X1 U7131 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9374) );
  MUX2_X1 U7132 ( .A(n8472), .B(n9374), .S(n4583), .Z(n5627) );
  XNOR2_X1 U7133 ( .A(n5627), .B(SI_29_), .ZN(n5620) );
  NAND2_X1 U7134 ( .A1(n8471), .A2(n5658), .ZN(n5622) );
  OR2_X1 U7135 ( .A1(n5660), .A2(n9374), .ZN(n5621) );
  INV_X1 U7136 ( .A(n5623), .ZN(n8456) );
  NAND2_X1 U7137 ( .A1(n5157), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U7138 ( .A1(n5640), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n5624) );
  OAI211_X1 U7139 ( .C1(n5644), .C2(n8896), .A(n5625), .B(n5624), .ZN(n5626)
         );
  AOI21_X1 U7140 ( .B1(n8456), .B2(n5431), .A(n5626), .ZN(n8614) );
  NAND2_X1 U7141 ( .A1(n9274), .A2(n8614), .ZN(n5789) );
  NAND2_X1 U7142 ( .A1(n8460), .A2(n8461), .ZN(n8459) );
  INV_X1 U7143 ( .A(n5627), .ZN(n5630) );
  NOR2_X1 U7144 ( .A1(n5630), .A2(SI_29_), .ZN(n5628) );
  NAND2_X1 U7145 ( .A1(n5630), .A2(SI_29_), .ZN(n5631) );
  MUX2_X1 U7146 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n4583), .Z(n5651) );
  NAND2_X1 U7147 ( .A1(n8351), .A2(n5658), .ZN(n5634) );
  INV_X1 U7148 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8352) );
  OR2_X1 U7149 ( .A1(n5660), .A2(n8352), .ZN(n5633) );
  NAND2_X1 U7150 ( .A1(n5157), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n5637) );
  INV_X1 U7151 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8675) );
  OR2_X1 U7152 ( .A1(n5644), .A2(n8675), .ZN(n5636) );
  INV_X1 U7153 ( .A(P2_REG0_REG_31__SCAN_IN), .ZN(n8934) );
  OR2_X1 U7154 ( .A1(n5174), .A2(n8934), .ZN(n5635) );
  AND3_X1 U7155 ( .A1(n5637), .A2(n5636), .A3(n5635), .ZN(n6669) );
  NAND2_X1 U7156 ( .A1(n6669), .A2(n6616), .ZN(n5645) );
  INV_X1 U7157 ( .A(n5638), .ZN(n5639) );
  NAND2_X1 U7158 ( .A1(n8459), .A2(n5639), .ZN(n5648) );
  INV_X1 U7159 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n5643) );
  NAND2_X1 U7160 ( .A1(n5157), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n5642) );
  NAND2_X1 U7161 ( .A1(n5640), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n5641) );
  OAI211_X1 U7162 ( .C1(n5644), .C2(n5643), .A(n5642), .B(n5641), .ZN(n8613)
         );
  INV_X1 U7163 ( .A(n8613), .ZN(n5663) );
  NAND2_X1 U7164 ( .A1(n5646), .A2(n5645), .ZN(n5647) );
  NAND2_X1 U7165 ( .A1(n5648), .A2(n5647), .ZN(n5664) );
  INV_X1 U7166 ( .A(n5649), .ZN(n5650) );
  NAND2_X1 U7167 ( .A1(n5650), .A2(SI_30_), .ZN(n5654) );
  NAND2_X1 U7168 ( .A1(n5652), .A2(n5651), .ZN(n5653) );
  NAND2_X1 U7169 ( .A1(n5654), .A2(n5653), .ZN(n5657) );
  MUX2_X1 U7170 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n4583), .Z(n5655) );
  XNOR2_X1 U7171 ( .A(n5655), .B(SI_31_), .ZN(n5656) );
  NAND2_X1 U7172 ( .A1(n9367), .A2(n5658), .ZN(n5662) );
  INV_X1 U7173 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5659) );
  OR2_X1 U7174 ( .A1(n5660), .A2(n5659), .ZN(n5661) );
  NAND2_X1 U7175 ( .A1(n8683), .A2(n5663), .ZN(n5790) );
  AND2_X2 U7176 ( .A1(n5796), .A2(n5790), .ZN(n5829) );
  AOI21_X1 U7177 ( .B1(n5664), .B2(n5829), .A(n5799), .ZN(n5665) );
  XNOR2_X1 U7178 ( .A(n5665), .B(n9194), .ZN(n5666) );
  AOI21_X1 U7179 ( .B1(n8314), .B2(n7024), .A(n5666), .ZN(n5843) );
  NAND2_X1 U7180 ( .A1(n9194), .A2(n7637), .ZN(n6614) );
  OR2_X2 U7181 ( .A1(n6614), .A2(n7520), .ZN(n5797) );
  INV_X1 U7182 ( .A(n5797), .ZN(n5782) );
  MUX2_X1 U7183 ( .A(n8617), .B(n7993), .S(n5782), .Z(n5726) );
  NAND2_X1 U7184 ( .A1(n5812), .A2(n5814), .ZN(n5670) );
  NAND2_X1 U7185 ( .A1(n5815), .A2(n5813), .ZN(n5669) );
  INV_X1 U7186 ( .A(n5689), .ZN(n5672) );
  OR2_X1 U7187 ( .A1(n8424), .A2(n8431), .ZN(n5810) );
  NAND2_X1 U7188 ( .A1(n5810), .A2(n6616), .ZN(n5675) );
  INV_X1 U7189 ( .A(n5809), .ZN(n7028) );
  OAI211_X1 U7190 ( .C1(n5675), .C2(n7028), .A(n5807), .B(n5808), .ZN(n5674)
         );
  NAND2_X1 U7191 ( .A1(n5674), .A2(n5806), .ZN(n5679) );
  INV_X1 U7192 ( .A(n5675), .ZN(n5676) );
  OAI211_X1 U7193 ( .C1(n5676), .C2(n7029), .A(n5806), .B(n5809), .ZN(n5677)
         );
  NAND2_X1 U7194 ( .A1(n5677), .A2(n5807), .ZN(n5678) );
  MUX2_X1 U7195 ( .A(n5679), .B(n5678), .S(n5797), .Z(n5680) );
  NAND2_X1 U7196 ( .A1(n5680), .A2(n7164), .ZN(n5681) );
  AND2_X1 U7197 ( .A1(n5814), .A2(n5682), .ZN(n5683) );
  OAI211_X1 U7198 ( .C1(n5684), .C2(n5683), .A(n5686), .B(n5812), .ZN(n5685)
         );
  AOI22_X1 U7199 ( .A1(n5687), .A2(n5686), .B1(n5782), .B2(n5685), .ZN(n5694)
         );
  INV_X1 U7200 ( .A(n5688), .ZN(n5690) );
  NAND2_X1 U7201 ( .A1(n5690), .A2(n5691), .ZN(n7441) );
  OAI21_X1 U7202 ( .B1(n5797), .B2(n5689), .A(n4913), .ZN(n5693) );
  MUX2_X1 U7203 ( .A(n5691), .B(n5690), .S(n5797), .Z(n5692) );
  INV_X1 U7204 ( .A(n10343), .ZN(n10347) );
  OAI211_X1 U7205 ( .C1(n5694), .C2(n5693), .A(n5692), .B(n10347), .ZN(n5695)
         );
  INV_X1 U7206 ( .A(n5696), .ZN(n5698) );
  OAI21_X1 U7207 ( .B1(n7453), .B2(n10356), .A(n5700), .ZN(n5697) );
  MUX2_X1 U7208 ( .A(n5698), .B(n5697), .S(n5797), .Z(n5699) );
  INV_X1 U7209 ( .A(n5700), .ZN(n5703) );
  NAND2_X1 U7210 ( .A1(n5705), .A2(n5701), .ZN(n5702) );
  MUX2_X1 U7211 ( .A(n5703), .B(n5702), .S(n5797), .Z(n5704) );
  INV_X1 U7212 ( .A(n5714), .ZN(n5805) );
  NAND2_X1 U7213 ( .A1(n5805), .A2(n5705), .ZN(n5708) );
  NAND2_X1 U7214 ( .A1(n5804), .A2(n5706), .ZN(n5707) );
  MUX2_X1 U7215 ( .A(n5708), .B(n5707), .S(n5797), .Z(n5709) );
  INV_X1 U7216 ( .A(n5715), .ZN(n5711) );
  NAND3_X1 U7217 ( .A1(n5711), .A2(n5804), .A3(n5710), .ZN(n5713) );
  AND2_X1 U7218 ( .A1(n5713), .A2(n5712), .ZN(n5716) );
  MUX2_X1 U7219 ( .A(n5718), .B(n5720), .S(n5797), .Z(n5717) );
  NAND3_X1 U7220 ( .A1(n5725), .A2(n5726), .A3(n5717), .ZN(n5722) );
  OAI21_X1 U7221 ( .B1(n7993), .B2(n5718), .A(n5737), .ZN(n5719) );
  AOI21_X1 U7222 ( .B1(n5722), .B2(n8617), .A(n5719), .ZN(n5724) );
  OAI21_X1 U7223 ( .B1(n8617), .B2(n5720), .A(n5734), .ZN(n5721) );
  AOI21_X1 U7224 ( .B1(n5722), .B2(n7993), .A(n5721), .ZN(n5723) );
  INV_X1 U7225 ( .A(n9245), .ZN(n9237) );
  INV_X1 U7226 ( .A(n5728), .ZN(n5730) );
  NAND2_X1 U7227 ( .A1(n5733), .A2(n9215), .ZN(n5729) );
  MUX2_X1 U7228 ( .A(n5730), .B(n5729), .S(n5797), .Z(n5732) );
  INV_X1 U7229 ( .A(n5736), .ZN(n5731) );
  OR2_X1 U7230 ( .A1(n5732), .A2(n5731), .ZN(n5738) );
  INV_X1 U7231 ( .A(n5738), .ZN(n5742) );
  OAI211_X1 U7232 ( .C1(n5738), .C2(n5734), .A(n5746), .B(n5733), .ZN(n5740)
         );
  INV_X1 U7233 ( .A(n5743), .ZN(n5735) );
  OAI211_X1 U7234 ( .C1(n5738), .C2(n5737), .A(n5736), .B(n5735), .ZN(n5739)
         );
  MUX2_X1 U7235 ( .A(n5740), .B(n5739), .S(n5797), .Z(n5741) );
  OAI21_X1 U7236 ( .B1(n5748), .B2(n5743), .A(n5749), .ZN(n5744) );
  NAND3_X1 U7237 ( .A1(n5744), .A2(n5747), .A3(n5751), .ZN(n5745) );
  NAND3_X1 U7238 ( .A1(n5752), .A2(n5755), .A3(n5751), .ZN(n5753) );
  NAND3_X1 U7239 ( .A1(n5753), .A2(n9144), .A3(n5757), .ZN(n5754) );
  AOI21_X1 U7240 ( .B1(n5756), .B2(n5755), .A(n5797), .ZN(n5759) );
  INV_X1 U7241 ( .A(n9120), .ZN(n9130) );
  MUX2_X1 U7242 ( .A(n5757), .B(n5756), .S(n5797), .Z(n5758) );
  MUX2_X1 U7243 ( .A(n5760), .B(n9109), .S(n5797), .Z(n5761) );
  MUX2_X1 U7244 ( .A(n5763), .B(n5762), .S(n5797), .Z(n5764) );
  INV_X1 U7245 ( .A(n5769), .ZN(n5766) );
  OAI21_X1 U7246 ( .B1(n5766), .B2(n5765), .A(n5767), .ZN(n5773) );
  INV_X1 U7247 ( .A(n5767), .ZN(n5771) );
  INV_X1 U7248 ( .A(n5768), .ZN(n5770) );
  OAI21_X1 U7249 ( .B1(n5771), .B2(n5770), .A(n5769), .ZN(n5772) );
  MUX2_X1 U7250 ( .A(n5773), .B(n5772), .S(n5797), .Z(n5774) );
  NAND2_X1 U7251 ( .A1(n5776), .A2(n5775), .ZN(n5778) );
  NOR2_X1 U7252 ( .A1(n9062), .A2(n9083), .ZN(n5777) );
  INV_X1 U7253 ( .A(n5781), .ZN(n5779) );
  OAI21_X1 U7254 ( .B1(n5782), .B2(n9280), .A(n5781), .ZN(n5786) );
  INV_X1 U7255 ( .A(n5788), .ZN(n5784) );
  OAI21_X1 U7256 ( .B1(n5784), .B2(n5797), .A(n5783), .ZN(n5785) );
  MUX2_X1 U7257 ( .A(n5789), .B(n5788), .S(n5797), .Z(n5792) );
  INV_X1 U7258 ( .A(n5790), .ZN(n5791) );
  INV_X1 U7259 ( .A(n5829), .ZN(n5794) );
  INV_X1 U7260 ( .A(n5799), .ZN(n5826) );
  NAND2_X1 U7261 ( .A1(n5826), .A2(n5827), .ZN(n5793) );
  MUX2_X1 U7262 ( .A(n5794), .B(n5793), .S(n5797), .Z(n5795) );
  INV_X1 U7263 ( .A(n5796), .ZN(n5798) );
  MUX2_X1 U7264 ( .A(n5799), .B(n5798), .S(n5797), .Z(n5800) );
  NAND2_X1 U7265 ( .A1(n9194), .A2(n7014), .ZN(n7023) );
  INV_X1 U7266 ( .A(n7023), .ZN(n5801) );
  INV_X1 U7267 ( .A(n9143), .ZN(n8446) );
  INV_X1 U7268 ( .A(n7995), .ZN(n7987) );
  NAND2_X1 U7269 ( .A1(n5805), .A2(n5804), .ZN(n7753) );
  INV_X1 U7270 ( .A(n7504), .ZN(n5819) );
  NOR2_X1 U7271 ( .A1(n7269), .A2(n7017), .ZN(n5811) );
  NAND2_X1 U7272 ( .A1(n5810), .A2(n7025), .ZN(n10406) );
  INV_X1 U7273 ( .A(n10406), .ZN(n7293) );
  NAND4_X1 U7274 ( .A1(n5811), .A2(n6615), .A3(n7164), .A4(n7293), .ZN(n5816)
         );
  NAND2_X1 U7275 ( .A1(n5813), .A2(n5812), .ZN(n7294) );
  NAND2_X1 U7276 ( .A1(n5815), .A2(n5814), .ZN(n7319) );
  NOR3_X1 U7277 ( .A1(n5816), .A2(n7294), .A3(n7319), .ZN(n5817) );
  NAND4_X1 U7278 ( .A1(n5817), .A2(n4913), .A3(n10375), .A4(n7452), .ZN(n5818)
         );
  NOR4_X1 U7279 ( .A1(n7753), .A2(n5819), .A3(n5818), .A4(n10343), .ZN(n5820)
         );
  NAND4_X1 U7280 ( .A1(n7987), .A2(n7872), .A3(n7849), .A4(n5820), .ZN(n5821)
         );
  NOR4_X1 U7281 ( .A1(n9222), .A2(n7992), .A3(n9245), .A4(n5821), .ZN(n5822)
         );
  XNOR2_X1 U7282 ( .A(n9329), .B(n9218), .ZN(n9208) );
  NAND4_X1 U7283 ( .A1(n9174), .A2(n9185), .A3(n5822), .A4(n9208), .ZN(n5823)
         );
  NOR4_X1 U7284 ( .A1(n9120), .A2(n8446), .A3(n9153), .A4(n5823), .ZN(n5824)
         );
  NAND4_X1 U7285 ( .A1(n9082), .A2(n9112), .A3(n8448), .A4(n5824), .ZN(n5825)
         );
  NOR4_X1 U7286 ( .A1(n8454), .A2(n9038), .A3(n9064), .A4(n5825), .ZN(n5828)
         );
  NAND4_X1 U7287 ( .A1(n5829), .A2(n5828), .A3(n5827), .A4(n5826), .ZN(n5830)
         );
  XNOR2_X1 U7288 ( .A(n5830), .B(n7237), .ZN(n5831) );
  OAI22_X1 U7289 ( .A1(n5831), .A2(n6616), .B1(n6615), .B2(n7023), .ZN(n5832)
         );
  AOI21_X1 U7290 ( .B1(n5836), .B2(n5835), .A(n9369), .ZN(n5837) );
  NAND2_X1 U7291 ( .A1(n5837), .A2(P2_IR_REG_23__SCAN_IN), .ZN(n5840) );
  INV_X1 U7292 ( .A(n5837), .ZN(n5839) );
  INV_X1 U7293 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5838) );
  NAND2_X1 U7294 ( .A1(n5839), .A2(n5838), .ZN(n5850) );
  NAND2_X1 U7295 ( .A1(n5840), .A2(n5850), .ZN(n6618) );
  OR2_X1 U7296 ( .A1(n6618), .A2(P2_U3152), .ZN(n7709) );
  INV_X1 U7297 ( .A(n7709), .ZN(n5841) );
  OAI21_X1 U7298 ( .B1(n5843), .B2(n5842), .A(n5841), .ZN(n5857) );
  INV_X1 U7299 ( .A(n6797), .ZN(n5845) );
  INV_X1 U7300 ( .A(n10366), .ZN(n9242) );
  NAND2_X1 U7301 ( .A1(n4569), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5846) );
  NAND2_X1 U7302 ( .A1(n5847), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5848) );
  MUX2_X1 U7303 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5848), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n5849) );
  AND2_X1 U7304 ( .A1(n5849), .A2(n4569), .ZN(n6606) );
  NAND2_X1 U7305 ( .A1(n6607), .A2(n6606), .ZN(n5853) );
  NAND2_X1 U7306 ( .A1(n5850), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5852) );
  INV_X1 U7307 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n5851) );
  NOR4_X1 U7308 ( .A1(n5844), .A2(n9242), .A3(n10385), .A4(n9385), .ZN(n5855)
         );
  OAI21_X1 U7309 ( .B1(n7709), .B2(n7014), .A(P2_B_REG_SCAN_IN), .ZN(n5854) );
  OR2_X1 U7310 ( .A1(n5855), .A2(n5854), .ZN(n5856) );
  NAND2_X1 U7311 ( .A1(n5857), .A2(n5856), .ZN(P2_U3244) );
  NAND4_X1 U7312 ( .A1(n5859), .A2(n5858), .A3(n6157), .A4(n6108), .ZN(n5862)
         );
  INV_X2 U7313 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6069) );
  NAND4_X1 U7314 ( .A1(n6111), .A2(n6177), .A3(n6069), .A4(n5860), .ZN(n5861)
         );
  NOR2_X1 U7315 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_16__SCAN_IN), .ZN(
        n5865) );
  NOR2_X1 U7316 ( .A1(P1_IR_REG_15__SCAN_IN), .A2(P1_IR_REG_21__SCAN_IN), .ZN(
        n5864) );
  NOR2_X1 U7317 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n5863) );
  INV_X2 U7318 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n5927) );
  INV_X2 U7319 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6282) );
  NOR2_X1 U7320 ( .A1(P1_IR_REG_26__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n5869) );
  NAND2_X1 U7321 ( .A1(n8011), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n5880) );
  INV_X1 U7322 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7549) );
  OR2_X1 U7323 ( .A1(n5982), .A2(n7549), .ZN(n5879) );
  INV_X1 U7324 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7548) );
  OR2_X1 U7325 ( .A1(n6003), .A2(n7548), .ZN(n5878) );
  INV_X1 U7326 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n8774) );
  OR2_X1 U7327 ( .A1(n5981), .A2(n8774), .ZN(n5877) );
  NAND2_X1 U7328 ( .A1(n5867), .A2(n5927), .ZN(n5988) );
  NAND2_X1 U7329 ( .A1(n5889), .A2(n5888), .ZN(n5884) );
  NAND2_X1 U7330 ( .A1(n5886), .A2(n5885), .ZN(n5908) );
  INV_X1 U7331 ( .A(n5914), .ZN(n5897) );
  NAND2_X1 U7332 ( .A1(n5890), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5894) );
  INV_X1 U7333 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n5891) );
  NAND2_X1 U7334 ( .A1(n5894), .A2(n5891), .ZN(n5892) );
  XNOR2_X1 U7335 ( .A(n5894), .B(P1_IR_REG_25__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U7336 ( .A1(n4563), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5895) );
  XNOR2_X1 U7337 ( .A(n5895), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6485) );
  AND2_X1 U7338 ( .A1(n6486), .A2(n6485), .ZN(n5896) );
  NAND2_X1 U7339 ( .A1(n6925), .A2(n6228), .ZN(n5907) );
  BUF_X8 U7340 ( .A(n5917), .Z(n6478) );
  INV_X1 U7341 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n5900) );
  XNOR2_X2 U7342 ( .A(n5902), .B(n5901), .ZN(n8271) );
  OR2_X1 U7343 ( .A1(n5903), .A2(n5900), .ZN(n5905) );
  XNOR2_X1 U7344 ( .A(n5905), .B(n5904), .ZN(n6886) );
  NAND2_X1 U7345 ( .A1(n6478), .A2(n7553), .ZN(n5906) );
  INV_X1 U7346 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n5909) );
  NAND2_X1 U7347 ( .A1(n5911), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5913) );
  XNOR2_X2 U7348 ( .A(n5913), .B(n5912), .ZN(n8229) );
  INV_X1 U7349 ( .A(n5975), .ZN(n5918) );
  NAND2_X1 U7350 ( .A1(n6481), .A2(n8266), .ZN(n5916) );
  AND2_X4 U7351 ( .A1(n5917), .A2(n5916), .ZN(n6474) );
  AOI22_X1 U7352 ( .A1(n6474), .A2(n6925), .B1(n6228), .B2(n7553), .ZN(n5974)
         );
  NAND2_X1 U7353 ( .A1(n5918), .A2(n5974), .ZN(n6920) );
  INV_X1 U7354 ( .A(n6920), .ZN(n5937) );
  INV_X1 U7355 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n5919) );
  INV_X1 U7356 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n5920) );
  OR2_X1 U7357 ( .A1(n6003), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5921) );
  NAND2_X1 U7358 ( .A1(n5922), .A2(n5921), .ZN(n5924) );
  INV_X1 U7359 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6694) );
  NOR2_X1 U7360 ( .A1(n5981), .A2(n6694), .ZN(n5923) );
  NAND2_X1 U7361 ( .A1(n9530), .A2(n6228), .ZN(n5932) );
  NAND2_X1 U7362 ( .A1(n5926), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5928) );
  XNOR2_X1 U7363 ( .A(n5928), .B(n5927), .ZN(n6831) );
  OR2_X1 U7364 ( .A1(n5992), .A2(n6631), .ZN(n5930) );
  OR2_X1 U7365 ( .A1(n6013), .A2(n6638), .ZN(n5929) );
  NAND2_X1 U7366 ( .A1(n6478), .A2(n7564), .ZN(n5931) );
  NAND2_X1 U7367 ( .A1(n5932), .A2(n5931), .ZN(n5933) );
  INV_X4 U7368 ( .A(n5953), .ZN(n6387) );
  NAND2_X1 U7369 ( .A1(n6474), .A2(n9530), .ZN(n5935) );
  NAND2_X1 U7370 ( .A1(n6228), .A2(n7564), .ZN(n5934) );
  AND2_X1 U7371 ( .A1(n5935), .A2(n5934), .ZN(n6921) );
  NOR2_X1 U7372 ( .A1(n5937), .A2(n5936), .ZN(n5976) );
  INV_X1 U7373 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n5938) );
  NOR2_X1 U7374 ( .A1(n5982), .A2(n5938), .ZN(n5940) );
  INV_X1 U7375 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10019) );
  NOR2_X1 U7376 ( .A1(n5981), .A2(n10019), .ZN(n5939) );
  NAND2_X1 U7377 ( .A1(n8011), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n5942) );
  INV_X1 U7378 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n5941) );
  NAND3_X1 U7379 ( .A1(n5943), .A2(n5942), .A3(n5059), .ZN(n6677) );
  NAND2_X1 U7380 ( .A1(n6677), .A2(n6474), .ZN(n5950) );
  INV_X1 U7381 ( .A(SI_0_), .ZN(n5945) );
  INV_X1 U7382 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5944) );
  OAI21_X1 U7383 ( .B1(n4583), .B2(n5945), .A(n5944), .ZN(n5947) );
  AND2_X1 U7384 ( .A1(n5947), .A2(n5946), .ZN(n9896) );
  NOR2_X1 U7385 ( .A1(n6539), .A2(n4694), .ZN(n5948) );
  NAND2_X1 U7386 ( .A1(n6677), .A2(n6228), .ZN(n5954) );
  NOR2_X1 U7387 ( .A1(n6539), .A2(n10019), .ZN(n5951) );
  AOI21_X1 U7388 ( .B1(n6478), .B2(n7369), .A(n5951), .ZN(n5952) );
  NAND2_X1 U7389 ( .A1(n5954), .A2(n5952), .ZN(n6762) );
  NAND3_X1 U7390 ( .A1(n5954), .A2(n5953), .A3(n5952), .ZN(n5955) );
  NAND2_X1 U7391 ( .A1(n6763), .A2(n5955), .ZN(n5970) );
  NAND2_X1 U7392 ( .A1(n8011), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n5960) );
  INV_X1 U7393 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5956) );
  INV_X1 U7394 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n7384) );
  INV_X1 U7395 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n6689) );
  INV_X1 U7396 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6629) );
  OR2_X1 U7397 ( .A1(n5992), .A2(n6629), .ZN(n5964) );
  INV_X1 U7398 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5962) );
  XNOR2_X1 U7399 ( .A(n5962), .B(n5961), .ZN(n6868) );
  NAND2_X1 U7400 ( .A1(n5966), .A2(n5965), .ZN(n5967) );
  XNOR2_X1 U7401 ( .A(n5967), .B(n6387), .ZN(n5971) );
  NAND2_X1 U7402 ( .A1(n5970), .A2(n5971), .ZN(n6935) );
  NAND2_X1 U7403 ( .A1(n6474), .A2(n9531), .ZN(n5969) );
  NAND2_X1 U7404 ( .A1(n6228), .A2(n7386), .ZN(n5968) );
  NAND2_X1 U7405 ( .A1(n5969), .A2(n5968), .ZN(n6937) );
  INV_X1 U7406 ( .A(n5970), .ZN(n5973) );
  INV_X1 U7407 ( .A(n5971), .ZN(n5972) );
  INV_X1 U7408 ( .A(n6922), .ZN(n5978) );
  INV_X1 U7409 ( .A(n6921), .ZN(n5977) );
  NAND2_X1 U7410 ( .A1(n5978), .A2(n5977), .ZN(n5979) );
  NAND2_X1 U7411 ( .A1(n5980), .A2(n5979), .ZN(n6982) );
  NAND2_X1 U7412 ( .A1(n8011), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n5986) );
  INV_X1 U7413 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6695) );
  OR2_X1 U7414 ( .A1(n8017), .A2(n6695), .ZN(n5985) );
  INV_X1 U7415 ( .A(n6004), .ZN(n6006) );
  OAI21_X1 U7416 ( .B1(P1_REG3_REG_3__SCAN_IN), .B2(P1_REG3_REG_4__SCAN_IN), 
        .A(n6006), .ZN(n6984) );
  OR2_X1 U7417 ( .A1(n6003), .A2(n6984), .ZN(n5984) );
  INV_X1 U7418 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6709) );
  OR2_X1 U7419 ( .A1(n5982), .A2(n6709), .ZN(n5983) );
  NAND2_X1 U7420 ( .A1(n9529), .A2(n6228), .ZN(n5996) );
  INV_X1 U7421 ( .A(n5987), .ZN(n5991) );
  NAND2_X1 U7422 ( .A1(n5988), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5989) );
  MUX2_X1 U7423 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5989), .S(
        P1_IR_REG_4__SCAN_IN), .Z(n5990) );
  NAND2_X1 U7424 ( .A1(n5991), .A2(n5990), .ZN(n10027) );
  OR2_X1 U7425 ( .A1(n6642), .A2(n6013), .ZN(n5994) );
  OR2_X1 U7426 ( .A1(n5992), .A2(n6640), .ZN(n5993) );
  NAND2_X1 U7427 ( .A1(n6478), .A2(n7197), .ZN(n5995) );
  NAND2_X1 U7428 ( .A1(n5996), .A2(n5995), .ZN(n5997) );
  INV_X4 U7429 ( .A(n6387), .ZN(n7389) );
  XNOR2_X1 U7430 ( .A(n5997), .B(n7389), .ZN(n5998) );
  AOI22_X1 U7431 ( .A1(n6474), .A2(n9529), .B1(n6228), .B2(n7197), .ZN(n5999)
         );
  XNOR2_X1 U7432 ( .A(n5998), .B(n5999), .ZN(n6983) );
  INV_X1 U7433 ( .A(n5998), .ZN(n6000) );
  NOR2_X1 U7434 ( .A1(n6000), .A2(n5999), .ZN(n6001) );
  AOI21_X2 U7435 ( .B1(n6982), .B2(n6983), .A(n6001), .ZN(n6022) );
  INV_X1 U7436 ( .A(n6022), .ZN(n6020) );
  NAND2_X1 U7437 ( .A1(n8011), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6011) );
  INV_X1 U7438 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n6002) );
  OR2_X1 U7439 ( .A1(n8013), .A2(n6002), .ZN(n6010) );
  NAND2_X1 U7440 ( .A1(n6004), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n6033) );
  INV_X1 U7441 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6005) );
  NAND2_X1 U7442 ( .A1(n6006), .A2(n6005), .ZN(n6007) );
  NAND2_X1 U7443 ( .A1(n6033), .A2(n6007), .ZN(n7054) );
  OR2_X1 U7444 ( .A1(n6526), .A2(n7054), .ZN(n6009) );
  INV_X1 U7445 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n6688) );
  OR2_X1 U7446 ( .A1(n8017), .A2(n6688), .ZN(n6008) );
  NAND4_X1 U7447 ( .A1(n6011), .A2(n6010), .A3(n6009), .A4(n6008), .ZN(n9528)
         );
  NAND2_X1 U7448 ( .A1(n9528), .A2(n6193), .ZN(n6017) );
  OR2_X1 U7449 ( .A1(n5987), .A2(n5900), .ZN(n6012) );
  XNOR2_X1 U7450 ( .A(n6012), .B(P1_IR_REG_5__SCAN_IN), .ZN(n10039) );
  AOI22_X1 U7451 ( .A1(n6301), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n6543), .B2(
        n10039), .ZN(n6015) );
  NAND2_X1 U7452 ( .A1(n6643), .A2(n8096), .ZN(n6014) );
  NAND2_X1 U7453 ( .A1(n6015), .A2(n6014), .ZN(n7398) );
  NAND2_X1 U7454 ( .A1(n6478), .A2(n7398), .ZN(n6016) );
  NAND2_X1 U7455 ( .A1(n6017), .A2(n6016), .ZN(n6018) );
  XNOR2_X1 U7456 ( .A(n6018), .B(n6387), .ZN(n6021) );
  INV_X1 U7457 ( .A(n6021), .ZN(n6019) );
  NAND2_X1 U7458 ( .A1(n6020), .A2(n6019), .ZN(n6023) );
  NAND2_X1 U7459 ( .A1(n6022), .A2(n6021), .ZN(n6027) );
  NAND2_X1 U7460 ( .A1(n6474), .A2(n9528), .ZN(n6025) );
  NAND2_X1 U7461 ( .A1(n6193), .A2(n7398), .ZN(n6024) );
  NAND2_X1 U7462 ( .A1(n6025), .A2(n6024), .ZN(n7053) );
  NAND2_X1 U7463 ( .A1(n6652), .A2(n8096), .ZN(n6031) );
  INV_X1 U7464 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7465 ( .A1(n5987), .A2(n6028), .ZN(n6048) );
  NAND2_X1 U7466 ( .A1(n6048), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6029) );
  XNOR2_X1 U7467 ( .A(n6029), .B(P1_IR_REG_6__SCAN_IN), .ZN(n6727) );
  AOI22_X1 U7468 ( .A1(n6301), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n6543), .B2(
        n6727), .ZN(n6030) );
  NAND2_X1 U7469 ( .A1(n6031), .A2(n6030), .ZN(n7466) );
  NAND2_X1 U7470 ( .A1(n7466), .A2(n6478), .ZN(n6040) );
  NAND2_X1 U7471 ( .A1(n8011), .A2(P1_REG0_REG_6__SCAN_IN), .ZN(n6038) );
  INV_X1 U7472 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6032) );
  OR2_X1 U7473 ( .A1(n8017), .A2(n6032), .ZN(n6037) );
  INV_X1 U7474 ( .A(n6052), .ZN(n6054) );
  NAND2_X1 U7475 ( .A1(n6033), .A2(n8893), .ZN(n6034) );
  NAND2_X1 U7476 ( .A1(n6054), .A2(n6034), .ZN(n7362) );
  OR2_X1 U7477 ( .A1(n6526), .A2(n7362), .ZN(n6036) );
  INV_X1 U7478 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7359) );
  OR2_X1 U7479 ( .A1(n8013), .A2(n7359), .ZN(n6035) );
  NAND4_X1 U7480 ( .A1(n6038), .A2(n6037), .A3(n6036), .A4(n6035), .ZN(n9526)
         );
  NAND2_X1 U7481 ( .A1(n9526), .A2(n6193), .ZN(n6039) );
  NAND2_X1 U7482 ( .A1(n6040), .A2(n6039), .ZN(n6041) );
  XNOR2_X1 U7483 ( .A(n6041), .B(n6387), .ZN(n6046) );
  NAND2_X1 U7484 ( .A1(n6474), .A2(n9526), .ZN(n6043) );
  NAND2_X1 U7485 ( .A1(n7466), .A2(n6193), .ZN(n6042) );
  NAND2_X1 U7486 ( .A1(n6043), .A2(n6042), .ZN(n6044) );
  XNOR2_X1 U7487 ( .A(n6046), .B(n6044), .ZN(n7134) );
  NAND2_X1 U7488 ( .A1(n7132), .A2(n7134), .ZN(n7133) );
  INV_X1 U7489 ( .A(n6044), .ZN(n6045) );
  NAND2_X1 U7490 ( .A1(n6046), .A2(n6045), .ZN(n6047) );
  NAND2_X1 U7491 ( .A1(n7133), .A2(n6047), .ZN(n7176) );
  INV_X1 U7492 ( .A(n7176), .ZN(n6066) );
  NAND2_X1 U7493 ( .A1(n6659), .A2(n8096), .ZN(n6050) );
  NAND2_X1 U7494 ( .A1(n6110), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6067) );
  XNOR2_X1 U7495 ( .A(n6067), .B(P1_IR_REG_7__SCAN_IN), .ZN(n6749) );
  AOI22_X1 U7496 ( .A1(n6301), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n6543), .B2(
        n6749), .ZN(n6049) );
  NAND2_X1 U7497 ( .A1(n6050), .A2(n6049), .ZN(n7532) );
  NAND2_X1 U7498 ( .A1(n7532), .A2(n6478), .ZN(n6061) );
  NAND2_X1 U7499 ( .A1(n8011), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n6059) );
  INV_X1 U7500 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6051) );
  OR2_X1 U7501 ( .A1(n8017), .A2(n6051), .ZN(n6058) );
  NAND2_X1 U7502 ( .A1(n6052), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n6074) );
  INV_X1 U7503 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n6053) );
  NAND2_X1 U7504 ( .A1(n6054), .A2(n6053), .ZN(n6055) );
  NAND2_X1 U7505 ( .A1(n6074), .A2(n6055), .ZN(n7529) );
  OR2_X1 U7506 ( .A1(n6526), .A2(n7529), .ZN(n6057) );
  INV_X1 U7507 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7530) );
  OR2_X1 U7508 ( .A1(n8013), .A2(n7530), .ZN(n6056) );
  NAND4_X1 U7509 ( .A1(n6059), .A2(n6058), .A3(n6057), .A4(n6056), .ZN(n9525)
         );
  NAND2_X1 U7510 ( .A1(n9525), .A2(n6193), .ZN(n6060) );
  NAND2_X1 U7511 ( .A1(n6061), .A2(n6060), .ZN(n6062) );
  XNOR2_X1 U7512 ( .A(n6062), .B(n6387), .ZN(n6064) );
  AOI22_X1 U7513 ( .A1(n7532), .A2(n6228), .B1(n6474), .B2(n9525), .ZN(n6063)
         );
  OR2_X1 U7514 ( .A1(n6064), .A2(n6063), .ZN(n7177) );
  NAND2_X1 U7515 ( .A1(n6662), .A2(n8096), .ZN(n6073) );
  NAND2_X1 U7516 ( .A1(n6067), .A2(n6108), .ZN(n6068) );
  NAND2_X1 U7517 ( .A1(n6068), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6070) );
  NAND2_X1 U7518 ( .A1(n6070), .A2(n6069), .ZN(n6088) );
  OR2_X1 U7519 ( .A1(n6070), .A2(n6069), .ZN(n6071) );
  AOI22_X1 U7520 ( .A1(n6301), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n6543), .B2(
        n10051), .ZN(n6072) );
  NAND2_X1 U7521 ( .A1(n6073), .A2(n6072), .ZN(n7595) );
  NAND2_X1 U7522 ( .A1(n8011), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n6079) );
  OR2_X1 U7523 ( .A1(n8017), .A2(n10241), .ZN(n6078) );
  NAND2_X1 U7524 ( .A1(n6074), .A2(n7435), .ZN(n6075) );
  NAND2_X1 U7525 ( .A1(n6092), .A2(n6075), .ZN(n7590) );
  OR2_X1 U7526 ( .A1(n6526), .A2(n7590), .ZN(n6077) );
  OR2_X1 U7527 ( .A1(n8013), .A2(n8772), .ZN(n6076) );
  NAND4_X1 U7528 ( .A1(n6079), .A2(n6078), .A3(n6077), .A4(n6076), .ZN(n9524)
         );
  AND2_X1 U7529 ( .A1(n6474), .A2(n9524), .ZN(n6080) );
  AOI21_X1 U7530 ( .B1(n7595), .B2(n6193), .A(n6080), .ZN(n6085) );
  NAND2_X1 U7531 ( .A1(n7595), .A2(n6478), .ZN(n6082) );
  NAND2_X1 U7532 ( .A1(n9524), .A2(n6193), .ZN(n6081) );
  NAND2_X1 U7533 ( .A1(n6082), .A2(n6081), .ZN(n6083) );
  XNOR2_X1 U7534 ( .A(n6083), .B(n7389), .ZN(n7434) );
  NAND2_X1 U7535 ( .A1(n7432), .A2(n7434), .ZN(n7429) );
  INV_X1 U7536 ( .A(n6084), .ZN(n6087) );
  INV_X1 U7537 ( .A(n6085), .ZN(n6086) );
  NAND2_X1 U7538 ( .A1(n6087), .A2(n6086), .ZN(n7430) );
  NAND2_X1 U7539 ( .A1(n6666), .A2(n8096), .ZN(n6091) );
  NAND2_X1 U7540 ( .A1(n6088), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6089) );
  XNOR2_X1 U7541 ( .A(n6089), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6746) );
  AOI22_X1 U7542 ( .A1(n6301), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n6543), .B2(
        n6746), .ZN(n6090) );
  NAND2_X1 U7543 ( .A1(n6091), .A2(n6090), .ZN(n7491) );
  NAND2_X1 U7544 ( .A1(n7491), .A2(n6478), .ZN(n6100) );
  NAND2_X1 U7545 ( .A1(n8011), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n6098) );
  INV_X1 U7546 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10180) );
  OR2_X1 U7547 ( .A1(n8013), .A2(n10180), .ZN(n6097) );
  INV_X1 U7548 ( .A(n6118), .ZN(n6119) );
  NAND2_X1 U7549 ( .A1(n6092), .A2(n7513), .ZN(n6093) );
  NAND2_X1 U7550 ( .A1(n6119), .A2(n6093), .ZN(n10179) );
  OR2_X1 U7551 ( .A1(n6526), .A2(n10179), .ZN(n6096) );
  INV_X1 U7552 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6094) );
  OR2_X1 U7553 ( .A1(n8017), .A2(n6094), .ZN(n6095) );
  NAND4_X1 U7554 ( .A1(n6098), .A2(n6097), .A3(n6096), .A4(n6095), .ZN(n9523)
         );
  NAND2_X1 U7555 ( .A1(n9523), .A2(n6228), .ZN(n6099) );
  NAND2_X1 U7556 ( .A1(n6100), .A2(n6099), .ZN(n6101) );
  XNOR2_X1 U7557 ( .A(n6101), .B(n7389), .ZN(n6103) );
  AND2_X1 U7558 ( .A1(n6474), .A2(n9523), .ZN(n6102) );
  AOI21_X1 U7559 ( .B1(n7491), .B2(n6193), .A(n6102), .ZN(n6104) );
  XNOR2_X1 U7560 ( .A(n6103), .B(n6104), .ZN(n7511) );
  INV_X1 U7561 ( .A(n6103), .ZN(n6105) );
  NAND2_X1 U7562 ( .A1(n6105), .A2(n6104), .ZN(n6106) );
  NAND2_X1 U7563 ( .A1(n6680), .A2(n8096), .ZN(n6117) );
  INV_X1 U7564 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n6107) );
  NAND3_X1 U7565 ( .A1(n6069), .A2(n6108), .A3(n6107), .ZN(n6109) );
  NAND2_X1 U7566 ( .A1(n6114), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6112) );
  MUX2_X1 U7567 ( .A(n6112), .B(P1_IR_REG_31__SCAN_IN), .S(n6111), .Z(n6113)
         );
  INV_X1 U7568 ( .A(n6113), .ZN(n6115) );
  NOR2_X1 U7569 ( .A1(n6115), .A2(n6158), .ZN(n6907) );
  AOI22_X1 U7570 ( .A1(n6301), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n6543), .B2(
        n6907), .ZN(n6116) );
  NAND2_X1 U7571 ( .A1(n7716), .A2(n6478), .ZN(n6130) );
  NAND2_X1 U7572 ( .A1(n6433), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6122) );
  INV_X1 U7573 ( .A(n6140), .ZN(n6142) );
  INV_X1 U7574 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n8792) );
  NAND2_X1 U7575 ( .A1(n6119), .A2(n8792), .ZN(n6120) );
  NAND2_X1 U7576 ( .A1(n6142), .A2(n6120), .ZN(n7544) );
  OR2_X1 U7577 ( .A1(n6526), .A2(n7544), .ZN(n6121) );
  NAND2_X1 U7578 ( .A1(n6122), .A2(n6121), .ZN(n6128) );
  INV_X1 U7579 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6124) );
  NOR2_X1 U7580 ( .A1(n6123), .A2(n6124), .ZN(n6127) );
  INV_X1 U7581 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6125) );
  NOR2_X1 U7582 ( .A1(n8017), .A2(n6125), .ZN(n6126) );
  NAND2_X1 U7583 ( .A1(n9522), .A2(n6193), .ZN(n6129) );
  NAND2_X1 U7584 ( .A1(n6130), .A2(n6129), .ZN(n6131) );
  XNOR2_X1 U7585 ( .A(n6131), .B(n6387), .ZN(n7539) );
  AND2_X1 U7586 ( .A1(n6474), .A2(n9522), .ZN(n6132) );
  AOI21_X1 U7587 ( .B1(n7716), .B2(n6193), .A(n6132), .ZN(n7538) );
  INV_X1 U7588 ( .A(n7539), .ZN(n6134) );
  INV_X1 U7589 ( .A(n7538), .ZN(n6133) );
  NAND2_X1 U7590 ( .A1(n6134), .A2(n6133), .ZN(n6135) );
  NAND2_X1 U7591 ( .A1(n6682), .A2(n8096), .ZN(n6138) );
  OR2_X1 U7592 ( .A1(n6158), .A2(n5900), .ZN(n6136) );
  XNOR2_X1 U7593 ( .A(n6136), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7113) );
  AOI22_X1 U7594 ( .A1(n6301), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n6543), .B2(
        n7113), .ZN(n6137) );
  NAND2_X1 U7595 ( .A1(n9973), .A2(n6478), .ZN(n6149) );
  INV_X1 U7596 ( .A(n8017), .ZN(n6525) );
  NAND2_X1 U7597 ( .A1(n6525), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6147) );
  INV_X1 U7598 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n6139) );
  OR2_X1 U7599 ( .A1(n6123), .A2(n6139), .ZN(n6146) );
  INV_X1 U7600 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7601 ( .A1(n6142), .A2(n6141), .ZN(n6143) );
  NAND2_X1 U7602 ( .A1(n6162), .A2(n6143), .ZN(n9974) );
  OR2_X1 U7603 ( .A1(n6526), .A2(n9974), .ZN(n6145) );
  INV_X1 U7604 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n9975) );
  OR2_X1 U7605 ( .A1(n8013), .A2(n9975), .ZN(n6144) );
  NAND4_X1 U7606 ( .A1(n6147), .A2(n6146), .A3(n6145), .A4(n6144), .ZN(n9521)
         );
  NAND2_X1 U7607 ( .A1(n9521), .A2(n6228), .ZN(n6148) );
  NAND2_X1 U7608 ( .A1(n6149), .A2(n6148), .ZN(n6150) );
  XNOR2_X1 U7609 ( .A(n6150), .B(n7389), .ZN(n6154) );
  AND2_X1 U7610 ( .A1(n6474), .A2(n9521), .ZN(n6151) );
  AOI21_X1 U7611 ( .B1(n9973), .B2(n6193), .A(n6151), .ZN(n6152) );
  XNOR2_X1 U7612 ( .A(n6154), .B(n6152), .ZN(n7639) );
  INV_X1 U7613 ( .A(n6152), .ZN(n6153) );
  NAND2_X1 U7614 ( .A1(n6154), .A2(n6153), .ZN(n6155) );
  NAND2_X1 U7615 ( .A1(n6156), .A2(n6155), .ZN(n7766) );
  NAND2_X1 U7616 ( .A1(n6825), .A2(n8096), .ZN(n6161) );
  NAND2_X1 U7617 ( .A1(n6158), .A2(n6157), .ZN(n6159) );
  NAND2_X1 U7618 ( .A1(n6159), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6178) );
  XNOR2_X1 U7619 ( .A(n6178), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10084) );
  AOI22_X1 U7620 ( .A1(n6301), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n10084), 
        .B2(n6543), .ZN(n6160) );
  NAND2_X1 U7621 ( .A1(n7779), .A2(n6478), .ZN(n6169) );
  NAND2_X1 U7622 ( .A1(n8011), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n6167) );
  INV_X1 U7623 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7728) );
  OR2_X1 U7624 ( .A1(n8013), .A2(n7728), .ZN(n6166) );
  NAND2_X1 U7625 ( .A1(n6162), .A2(n7768), .ZN(n6163) );
  NAND2_X1 U7626 ( .A1(n6184), .A2(n6163), .ZN(n7772) );
  OR2_X1 U7627 ( .A1(n6526), .A2(n7772), .ZN(n6165) );
  INV_X1 U7628 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n7102) );
  OR2_X1 U7629 ( .A1(n8017), .A2(n7102), .ZN(n6164) );
  NAND4_X1 U7630 ( .A1(n6167), .A2(n6166), .A3(n6165), .A4(n6164), .ZN(n9944)
         );
  NAND2_X1 U7631 ( .A1(n9944), .A2(n6193), .ZN(n6168) );
  NAND2_X1 U7632 ( .A1(n6169), .A2(n6168), .ZN(n6170) );
  XNOR2_X1 U7633 ( .A(n6170), .B(n6387), .ZN(n6172) );
  AND2_X1 U7634 ( .A1(n6474), .A2(n9944), .ZN(n6171) );
  AOI21_X1 U7635 ( .B1(n7779), .B2(n6193), .A(n6171), .ZN(n6173) );
  NAND2_X1 U7636 ( .A1(n6172), .A2(n6173), .ZN(n7764) );
  NAND2_X1 U7637 ( .A1(n7766), .A2(n7764), .ZN(n6176) );
  INV_X1 U7638 ( .A(n6172), .ZN(n6175) );
  INV_X1 U7639 ( .A(n6173), .ZN(n6174) );
  NAND2_X1 U7640 ( .A1(n6175), .A2(n6174), .ZN(n7765) );
  NAND2_X1 U7641 ( .A1(n6948), .A2(n8096), .ZN(n6182) );
  NAND2_X1 U7642 ( .A1(n6178), .A2(n6177), .ZN(n6179) );
  NAND2_X1 U7643 ( .A1(n6179), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6180) );
  XNOR2_X1 U7644 ( .A(n6180), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10097) );
  AOI22_X1 U7645 ( .A1(n10097), .A2(n6543), .B1(n6301), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n6181) );
  NAND2_X1 U7646 ( .A1(n9956), .A2(n6478), .ZN(n6191) );
  NAND2_X1 U7647 ( .A1(n8011), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n6189) );
  INV_X1 U7648 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n7104) );
  OR2_X1 U7649 ( .A1(n8017), .A2(n7104), .ZN(n6188) );
  INV_X1 U7650 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7651 ( .A1(n6184), .A2(n6183), .ZN(n6185) );
  NAND2_X1 U7652 ( .A1(n6201), .A2(n6185), .ZN(n9940) );
  OR2_X1 U7653 ( .A1(n6526), .A2(n9940), .ZN(n6187) );
  INV_X1 U7654 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9941) );
  OR2_X1 U7655 ( .A1(n8013), .A2(n9941), .ZN(n6186) );
  NAND4_X1 U7656 ( .A1(n6189), .A2(n6188), .A3(n6187), .A4(n6186), .ZN(n9520)
         );
  NAND2_X1 U7657 ( .A1(n9520), .A2(n6193), .ZN(n6190) );
  NAND2_X1 U7658 ( .A1(n6191), .A2(n6190), .ZN(n6192) );
  XNOR2_X1 U7659 ( .A(n6192), .B(n7389), .ZN(n7833) );
  NAND2_X1 U7660 ( .A1(n9956), .A2(n6193), .ZN(n6195) );
  NAND2_X1 U7661 ( .A1(n6474), .A2(n9520), .ZN(n6194) );
  NAND2_X1 U7662 ( .A1(n6195), .A2(n6194), .ZN(n7834) );
  NAND2_X1 U7663 ( .A1(n6953), .A2(n8096), .ZN(n6199) );
  OR2_X1 U7664 ( .A1(n6196), .A2(n5900), .ZN(n6197) );
  XNOR2_X1 U7665 ( .A(n6197), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7106) );
  AOI22_X1 U7666 ( .A1(n6301), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n6543), .B2(
        n7106), .ZN(n6198) );
  NAND2_X1 U7667 ( .A1(n7917), .A2(n6193), .ZN(n6209) );
  NAND2_X1 U7668 ( .A1(n8011), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n6207) );
  INV_X1 U7669 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6200) );
  OR2_X1 U7670 ( .A1(n8017), .A2(n6200), .ZN(n6206) );
  INV_X1 U7671 ( .A(n6220), .ZN(n6222) );
  NAND2_X1 U7672 ( .A1(n6201), .A2(n7109), .ZN(n6202) );
  NAND2_X1 U7673 ( .A1(n6222), .A2(n6202), .ZN(n7915) );
  OR2_X1 U7674 ( .A1(n6526), .A2(n7915), .ZN(n6205) );
  INV_X1 U7675 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n6203) );
  OR2_X1 U7676 ( .A1(n8013), .A2(n6203), .ZN(n6204) );
  NAND4_X1 U7677 ( .A1(n6207), .A2(n6206), .A3(n6205), .A4(n6204), .ZN(n9946)
         );
  NAND2_X1 U7678 ( .A1(n6474), .A2(n9946), .ZN(n6208) );
  NAND2_X1 U7679 ( .A1(n7917), .A2(n6478), .ZN(n6211) );
  NAND2_X1 U7680 ( .A1(n9946), .A2(n6193), .ZN(n6210) );
  NAND2_X1 U7681 ( .A1(n6211), .A2(n6210), .ZN(n6212) );
  XNOR2_X1 U7682 ( .A(n6212), .B(n6387), .ZN(n7908) );
  NAND2_X1 U7683 ( .A1(n6255), .A2(n7908), .ZN(n6232) );
  INV_X1 U7684 ( .A(n7907), .ZN(n6213) );
  NAND2_X1 U7685 ( .A1(n6214), .A2(n6213), .ZN(n6257) );
  NAND2_X1 U7686 ( .A1(n7044), .A2(n8096), .ZN(n6219) );
  INV_X1 U7687 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6215) );
  NAND2_X1 U7688 ( .A1(n6196), .A2(n6215), .ZN(n6216) );
  NAND2_X1 U7689 ( .A1(n6216), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6217) );
  XNOR2_X1 U7690 ( .A(n6217), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10109) );
  AOI22_X1 U7691 ( .A1(n6301), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n6543), .B2(
        n10109), .ZN(n6218) );
  NAND2_X1 U7692 ( .A1(n9856), .A2(n6478), .ZN(n6230) );
  NAND2_X1 U7693 ( .A1(n8011), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n6227) );
  INV_X1 U7694 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n9545) );
  OR2_X1 U7695 ( .A1(n8017), .A2(n9545), .ZN(n6226) );
  INV_X1 U7696 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n6221) );
  NAND2_X1 U7697 ( .A1(n6222), .A2(n6221), .ZN(n6223) );
  NAND2_X1 U7698 ( .A1(n6236), .A2(n6223), .ZN(n9509) );
  OR2_X1 U7699 ( .A1(n6526), .A2(n9509), .ZN(n6225) );
  INV_X1 U7700 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7901) );
  OR2_X1 U7701 ( .A1(n8013), .A2(n7901), .ZN(n6224) );
  NAND4_X1 U7702 ( .A1(n6227), .A2(n6226), .A3(n6225), .A4(n6224), .ZN(n9770)
         );
  NAND2_X1 U7703 ( .A1(n9770), .A2(n6228), .ZN(n6229) );
  NAND2_X1 U7704 ( .A1(n6230), .A2(n6229), .ZN(n6231) );
  XNOR2_X1 U7705 ( .A(n6231), .B(n7389), .ZN(n6253) );
  NAND3_X1 U7706 ( .A1(n6232), .A2(n6257), .A3(n6253), .ZN(n9430) );
  NAND2_X1 U7707 ( .A1(n7042), .A2(n8096), .ZN(n6235) );
  NAND2_X1 U7708 ( .A1(n6233), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6265) );
  XNOR2_X1 U7709 ( .A(n6265), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10120) );
  AOI22_X1 U7710 ( .A1(n6301), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n6543), .B2(
        n10120), .ZN(n6234) );
  NAND2_X1 U7711 ( .A1(n9850), .A2(n6478), .ZN(n6245) );
  NAND2_X1 U7712 ( .A1(n6236), .A2(n9436), .ZN(n6237) );
  NAND2_X1 U7713 ( .A1(n6270), .A2(n6237), .ZN(n9435) );
  INV_X1 U7714 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n6238) );
  OR2_X1 U7715 ( .A1(n6123), .A2(n6238), .ZN(n6241) );
  INV_X1 U7716 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n6239) );
  OR2_X1 U7717 ( .A1(n8013), .A2(n6239), .ZN(n6240) );
  AND2_X1 U7718 ( .A1(n6241), .A2(n6240), .ZN(n6243) );
  INV_X1 U7719 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9546) );
  OR2_X1 U7720 ( .A1(n8017), .A2(n9546), .ZN(n6242) );
  OAI211_X1 U7721 ( .C1(n9435), .C2(n6526), .A(n6243), .B(n6242), .ZN(n9751)
         );
  NAND2_X1 U7722 ( .A1(n9751), .A2(n6193), .ZN(n6244) );
  NAND2_X1 U7723 ( .A1(n6245), .A2(n6244), .ZN(n6246) );
  XNOR2_X1 U7724 ( .A(n6246), .B(n6387), .ZN(n6248) );
  AND2_X1 U7725 ( .A1(n6474), .A2(n9751), .ZN(n6247) );
  AOI21_X1 U7726 ( .B1(n9850), .B2(n6193), .A(n6247), .ZN(n6249) );
  NAND2_X1 U7727 ( .A1(n6248), .A2(n6249), .ZN(n6263) );
  INV_X1 U7728 ( .A(n6248), .ZN(n6251) );
  INV_X1 U7729 ( .A(n6249), .ZN(n6250) );
  NAND2_X1 U7730 ( .A1(n6251), .A2(n6250), .ZN(n6252) );
  AND2_X1 U7731 ( .A1(n6263), .A2(n6252), .ZN(n9431) );
  AND2_X1 U7732 ( .A1(n9430), .A2(n9431), .ZN(n6262) );
  INV_X1 U7733 ( .A(n6253), .ZN(n6254) );
  AND2_X1 U7734 ( .A1(n6255), .A2(n6254), .ZN(n6259) );
  INV_X1 U7735 ( .A(n7908), .ZN(n6256) );
  NAND2_X1 U7736 ( .A1(n6257), .A2(n6256), .ZN(n6258) );
  NAND2_X1 U7737 ( .A1(n6259), .A2(n6258), .ZN(n9501) );
  NAND2_X1 U7738 ( .A1(n9856), .A2(n6193), .ZN(n6261) );
  NAND2_X1 U7739 ( .A1(n6474), .A2(n9770), .ZN(n6260) );
  NAND2_X1 U7740 ( .A1(n6261), .A2(n6260), .ZN(n9503) );
  NAND2_X1 U7741 ( .A1(n6262), .A2(n9432), .ZN(n9429) );
  NAND2_X1 U7742 ( .A1(n9429), .A2(n6263), .ZN(n9443) );
  NAND2_X1 U7743 ( .A1(n7078), .A2(n8096), .ZN(n6268) );
  NAND2_X1 U7744 ( .A1(n6265), .A2(n6264), .ZN(n6266) );
  NAND2_X1 U7745 ( .A1(n6266), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6283) );
  XNOR2_X1 U7746 ( .A(n6283), .B(P1_IR_REG_17__SCAN_IN), .ZN(n10133) );
  AOI22_X1 U7747 ( .A1(n6301), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n6543), .B2(
        n10133), .ZN(n6267) );
  NAND2_X1 U7748 ( .A1(n9845), .A2(n6478), .ZN(n6275) );
  INV_X1 U7749 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9548) );
  INV_X1 U7750 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n6269) );
  INV_X1 U7751 ( .A(n6288), .ZN(n6290) );
  NAND2_X1 U7752 ( .A1(n6270), .A2(n6269), .ZN(n6271) );
  NAND2_X1 U7753 ( .A1(n6290), .A2(n6271), .ZN(n9744) );
  OR2_X1 U7754 ( .A1(n9744), .A2(n6526), .ZN(n6273) );
  AOI22_X1 U7755 ( .A1(n8011), .A2(P1_REG0_REG_17__SCAN_IN), .B1(n6433), .B2(
        P1_REG2_REG_17__SCAN_IN), .ZN(n6272) );
  OAI211_X1 U7756 ( .C1(n8017), .C2(n9548), .A(n6273), .B(n6272), .ZN(n9771)
         );
  NAND2_X1 U7757 ( .A1(n9771), .A2(n6193), .ZN(n6274) );
  NAND2_X1 U7758 ( .A1(n6275), .A2(n6274), .ZN(n6276) );
  XNOR2_X1 U7759 ( .A(n6276), .B(n7389), .ZN(n6278) );
  AND2_X1 U7760 ( .A1(n9771), .A2(n6474), .ZN(n6277) );
  AOI21_X1 U7761 ( .B1(n9845), .B2(n6193), .A(n6277), .ZN(n6279) );
  XNOR2_X1 U7762 ( .A(n6278), .B(n6279), .ZN(n9444) );
  NAND2_X1 U7763 ( .A1(n9443), .A2(n9444), .ZN(n9442) );
  INV_X1 U7764 ( .A(n6278), .ZN(n6280) );
  NAND2_X1 U7765 ( .A1(n6280), .A2(n6279), .ZN(n6281) );
  NAND2_X1 U7766 ( .A1(n7257), .A2(n8096), .ZN(n6287) );
  NAND2_X1 U7767 ( .A1(n6283), .A2(n6282), .ZN(n6284) );
  NAND2_X1 U7768 ( .A1(n6284), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6285) );
  XNOR2_X1 U7769 ( .A(n6285), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U7770 ( .A1(n6301), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n10149), 
        .B2(n6543), .ZN(n6286) );
  NAND2_X1 U7771 ( .A1(n9838), .A2(n6478), .ZN(n6295) );
  INV_X1 U7772 ( .A(n6304), .ZN(n6306) );
  INV_X1 U7773 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n6289) );
  NAND2_X1 U7774 ( .A1(n6290), .A2(n6289), .ZN(n6291) );
  NAND2_X1 U7775 ( .A1(n6306), .A2(n6291), .ZN(n9734) );
  AOI22_X1 U7776 ( .A1(n6525), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n8011), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n6293) );
  INV_X1 U7777 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9735) );
  OR2_X1 U7778 ( .A1(n8013), .A2(n9735), .ZN(n6292) );
  OAI211_X1 U7779 ( .C1(n9734), .C2(n6526), .A(n6293), .B(n6292), .ZN(n9752)
         );
  NAND2_X1 U7780 ( .A1(n9752), .A2(n6193), .ZN(n6294) );
  NAND2_X1 U7781 ( .A1(n6295), .A2(n6294), .ZN(n6296) );
  XNOR2_X1 U7782 ( .A(n6296), .B(n6387), .ZN(n6299) );
  INV_X1 U7783 ( .A(n6299), .ZN(n6297) );
  AND2_X1 U7784 ( .A1(n9752), .A2(n6474), .ZN(n6298) );
  AOI21_X1 U7785 ( .B1(n9838), .B2(n6193), .A(n6298), .ZN(n9480) );
  NAND2_X1 U7786 ( .A1(n6300), .A2(n6299), .ZN(n9481) );
  NAND2_X1 U7787 ( .A1(n7285), .A2(n8096), .ZN(n6303) );
  AOI22_X1 U7788 ( .A1(n6301), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n4695), .B2(
        n6543), .ZN(n6302) );
  NAND2_X1 U7789 ( .A1(n9833), .A2(n6478), .ZN(n6314) );
  INV_X1 U7790 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n6305) );
  NAND2_X1 U7791 ( .A1(n6306), .A2(n6305), .ZN(n6307) );
  NAND2_X1 U7792 ( .A1(n6324), .A2(n6307), .ZN(n9720) );
  OR2_X1 U7793 ( .A1(n9720), .A2(n6526), .ZN(n6312) );
  INV_X1 U7794 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n9552) );
  NAND2_X1 U7795 ( .A1(n6433), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n6309) );
  INV_X1 U7796 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n8885) );
  OR2_X1 U7797 ( .A1(n6123), .A2(n8885), .ZN(n6308) );
  OAI211_X1 U7798 ( .C1(n9552), .C2(n8017), .A(n6309), .B(n6308), .ZN(n6310)
         );
  INV_X1 U7799 ( .A(n6310), .ZN(n6311) );
  NAND2_X1 U7800 ( .A1(n6312), .A2(n6311), .ZN(n9727) );
  NAND2_X1 U7801 ( .A1(n9727), .A2(n6193), .ZN(n6313) );
  NAND2_X1 U7802 ( .A1(n6314), .A2(n6313), .ZN(n6315) );
  XNOR2_X1 U7803 ( .A(n6315), .B(n7389), .ZN(n6317) );
  AND2_X1 U7804 ( .A1(n9727), .A2(n6474), .ZN(n6316) );
  AOI21_X1 U7805 ( .B1(n9833), .B2(n6193), .A(n6316), .ZN(n6318) );
  XNOR2_X1 U7806 ( .A(n6317), .B(n6318), .ZN(n9409) );
  INV_X1 U7807 ( .A(n6317), .ZN(n6319) );
  NAND2_X1 U7808 ( .A1(n6319), .A2(n6318), .ZN(n6320) );
  NAND2_X1 U7809 ( .A1(n7408), .A2(n8096), .ZN(n6322) );
  OR2_X1 U7810 ( .A1(n5992), .A2(n8898), .ZN(n6321) );
  NAND2_X1 U7811 ( .A1(n9826), .A2(n6478), .ZN(n6333) );
  INV_X1 U7812 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n6323) );
  NAND2_X1 U7813 ( .A1(n6324), .A2(n6323), .ZN(n6325) );
  AND2_X1 U7814 ( .A1(n6344), .A2(n6325), .ZN(n9701) );
  INV_X1 U7815 ( .A(n6526), .ZN(n6326) );
  NAND2_X1 U7816 ( .A1(n9701), .A2(n6326), .ZN(n6331) );
  INV_X1 U7817 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8870) );
  NAND2_X1 U7818 ( .A1(n8011), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U7819 ( .A1(n6433), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n6327) );
  OAI211_X1 U7820 ( .C1(n8017), .C2(n8870), .A(n6328), .B(n6327), .ZN(n6329)
         );
  INV_X1 U7821 ( .A(n6329), .ZN(n6330) );
  NAND2_X1 U7822 ( .A1(n6331), .A2(n6330), .ZN(n9519) );
  NAND2_X1 U7823 ( .A1(n9519), .A2(n6193), .ZN(n6332) );
  NAND2_X1 U7824 ( .A1(n6333), .A2(n6332), .ZN(n6334) );
  XNOR2_X1 U7825 ( .A(n6334), .B(n7389), .ZN(n6337) );
  NAND2_X1 U7826 ( .A1(n9826), .A2(n6193), .ZN(n6336) );
  NAND2_X1 U7827 ( .A1(n9519), .A2(n6474), .ZN(n6335) );
  NAND2_X1 U7828 ( .A1(n6336), .A2(n6335), .ZN(n6338) );
  NAND2_X1 U7829 ( .A1(n6337), .A2(n6338), .ZN(n9461) );
  INV_X1 U7830 ( .A(n6337), .ZN(n6340) );
  INV_X1 U7831 ( .A(n6338), .ZN(n6339) );
  NAND2_X1 U7832 ( .A1(n6340), .A2(n6339), .ZN(n9460) );
  NAND2_X1 U7833 ( .A1(n7508), .A2(n8096), .ZN(n6342) );
  OR2_X1 U7834 ( .A1(n5992), .A2(n8749), .ZN(n6341) );
  NAND2_X1 U7835 ( .A1(n9823), .A2(n6478), .ZN(n6352) );
  INV_X1 U7836 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n6343) );
  AND2_X1 U7837 ( .A1(n6344), .A2(n6343), .ZN(n6345) );
  OR2_X1 U7838 ( .A1(n6345), .A2(n6360), .ZN(n9692) );
  INV_X1 U7839 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n6348) );
  NAND2_X1 U7840 ( .A1(n6433), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n6347) );
  NAND2_X1 U7841 ( .A1(n8011), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n6346) );
  OAI211_X1 U7842 ( .C1(n8017), .C2(n6348), .A(n6347), .B(n6346), .ZN(n6349)
         );
  INV_X1 U7843 ( .A(n6349), .ZN(n6350) );
  OAI21_X1 U7844 ( .B1(n9692), .B2(n6526), .A(n6350), .ZN(n9707) );
  NAND2_X1 U7845 ( .A1(n9707), .A2(n6193), .ZN(n6351) );
  NAND2_X1 U7846 ( .A1(n6352), .A2(n6351), .ZN(n6353) );
  XNOR2_X1 U7847 ( .A(n6353), .B(n7389), .ZN(n6355) );
  AND2_X1 U7848 ( .A1(n9707), .A2(n6474), .ZN(n6354) );
  AOI21_X1 U7849 ( .B1(n9823), .B2(n6193), .A(n6354), .ZN(n6356) );
  XNOR2_X1 U7850 ( .A(n6355), .B(n6356), .ZN(n9415) );
  INV_X1 U7851 ( .A(n6355), .ZN(n6357) );
  NAND2_X1 U7852 ( .A1(n7635), .A2(n8096), .ZN(n6359) );
  OR2_X1 U7853 ( .A1(n5992), .A2(n8474), .ZN(n6358) );
  OR2_X1 U7854 ( .A1(n6360), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6361) );
  NAND2_X1 U7855 ( .A1(n6360), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U7856 ( .A1(n6361), .A2(n6379), .ZN(n9670) );
  OR2_X1 U7857 ( .A1(n9670), .A2(n6526), .ZN(n6366) );
  INV_X1 U7858 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8764) );
  NAND2_X1 U7859 ( .A1(n6433), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n6363) );
  INV_X1 U7860 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8856) );
  OR2_X1 U7861 ( .A1(n6123), .A2(n8856), .ZN(n6362) );
  OAI211_X1 U7862 ( .C1(n8017), .C2(n8764), .A(n6363), .B(n6362), .ZN(n6364)
         );
  INV_X1 U7863 ( .A(n6364), .ZN(n6365) );
  NAND2_X1 U7864 ( .A1(n6366), .A2(n6365), .ZN(n9662) );
  AND2_X1 U7865 ( .A1(n9662), .A2(n6474), .ZN(n6367) );
  AOI21_X1 U7866 ( .B1(n9816), .B2(n6193), .A(n6367), .ZN(n6372) );
  NAND2_X1 U7867 ( .A1(n6371), .A2(n6372), .ZN(n9469) );
  NAND2_X1 U7868 ( .A1(n9816), .A2(n6478), .ZN(n6369) );
  NAND2_X1 U7869 ( .A1(n9662), .A2(n6193), .ZN(n6368) );
  NAND2_X1 U7870 ( .A1(n6369), .A2(n6368), .ZN(n6370) );
  NAND2_X1 U7871 ( .A1(n9469), .A2(n9472), .ZN(n6375) );
  AND2_X2 U7872 ( .A1(n6375), .A2(n9470), .ZN(n6391) );
  NAND2_X1 U7873 ( .A1(n7712), .A2(n8096), .ZN(n6377) );
  OR2_X1 U7874 ( .A1(n5992), .A2(n7715), .ZN(n6376) );
  NAND2_X1 U7875 ( .A1(n9811), .A2(n6478), .ZN(n6386) );
  NAND2_X1 U7876 ( .A1(n8011), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n6384) );
  INV_X1 U7877 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6378) );
  OR2_X1 U7878 ( .A1(n8013), .A2(n6378), .ZN(n6383) );
  XNOR2_X1 U7879 ( .A(P1_REG3_REG_23__SCAN_IN), .B(n6398), .ZN(n9656) );
  OR2_X1 U7880 ( .A1(n6526), .A2(n9656), .ZN(n6382) );
  INV_X1 U7881 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n6380) );
  OR2_X1 U7882 ( .A1(n8017), .A2(n6380), .ZN(n6381) );
  NAND4_X1 U7883 ( .A1(n6384), .A2(n6383), .A3(n6382), .A4(n6381), .ZN(n9677)
         );
  NAND2_X1 U7884 ( .A1(n9677), .A2(n6193), .ZN(n6385) );
  NAND2_X1 U7885 ( .A1(n6386), .A2(n6385), .ZN(n6388) );
  XNOR2_X1 U7886 ( .A(n6388), .B(n6387), .ZN(n6392) );
  NAND2_X1 U7887 ( .A1(n9811), .A2(n6193), .ZN(n6390) );
  NAND2_X1 U7888 ( .A1(n6474), .A2(n9677), .ZN(n6389) );
  NAND2_X1 U7889 ( .A1(n6390), .A2(n6389), .ZN(n9399) );
  INV_X1 U7890 ( .A(n6392), .ZN(n6393) );
  NAND2_X1 U7891 ( .A1(n7776), .A2(n8096), .ZN(n6396) );
  OR2_X1 U7892 ( .A1(n5992), .A2(n7777), .ZN(n6395) );
  NAND2_X1 U7893 ( .A1(n6525), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n6406) );
  INV_X1 U7894 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n6397) );
  OR2_X1 U7895 ( .A1(n6123), .A2(n6397), .ZN(n6405) );
  NAND3_X1 U7896 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(P1_REG3_REG_24__SCAN_IN), 
        .A3(n6398), .ZN(n6417) );
  INV_X1 U7897 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n6400) );
  NAND2_X1 U7898 ( .A1(P1_REG3_REG_23__SCAN_IN), .A2(n6398), .ZN(n6399) );
  NAND2_X1 U7899 ( .A1(n6400), .A2(n6399), .ZN(n6401) );
  NAND2_X1 U7900 ( .A1(n6417), .A2(n6401), .ZN(n9642) );
  OR2_X1 U7901 ( .A1(n6526), .A2(n9642), .ZN(n6404) );
  INV_X1 U7902 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n6402) );
  OR2_X1 U7903 ( .A1(n8013), .A2(n6402), .ZN(n6403) );
  NAND4_X1 U7904 ( .A1(n6406), .A2(n6405), .A3(n6404), .A4(n6403), .ZN(n9663)
         );
  AOI22_X1 U7905 ( .A1(n9633), .A2(n6193), .B1(n6474), .B2(n9663), .ZN(n6411)
         );
  NAND2_X1 U7906 ( .A1(n9633), .A2(n6478), .ZN(n6408) );
  NAND2_X1 U7907 ( .A1(n9663), .A2(n6193), .ZN(n6407) );
  NAND2_X1 U7908 ( .A1(n6408), .A2(n6407), .ZN(n6409) );
  XNOR2_X1 U7909 ( .A(n6409), .B(n7389), .ZN(n6410) );
  XOR2_X1 U7910 ( .A(n6411), .B(n6410), .Z(n9451) );
  INV_X1 U7911 ( .A(n6410), .ZN(n6412) );
  OR2_X1 U7912 ( .A1(n5992), .A2(n7925), .ZN(n6413) );
  NAND2_X1 U7913 ( .A1(n8011), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n6423) );
  INV_X1 U7914 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n6415) );
  OR2_X1 U7915 ( .A1(n8017), .A2(n6415), .ZN(n6422) );
  INV_X1 U7916 ( .A(n6417), .ZN(n6416) );
  NAND2_X1 U7917 ( .A1(n6416), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n6436) );
  INV_X1 U7918 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8931) );
  NAND2_X1 U7919 ( .A1(n6417), .A2(n8931), .ZN(n6418) );
  NAND2_X1 U7920 ( .A1(n6436), .A2(n6418), .ZN(n9620) );
  OR2_X1 U7921 ( .A1(n6526), .A2(n9620), .ZN(n6421) );
  INV_X1 U7922 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n6419) );
  OR2_X1 U7923 ( .A1(n8013), .A2(n6419), .ZN(n6420) );
  NAND4_X1 U7924 ( .A1(n6423), .A2(n6422), .A3(n6421), .A4(n6420), .ZN(n9518)
         );
  AOI22_X1 U7925 ( .A1(n9799), .A2(n6193), .B1(n6474), .B2(n9518), .ZN(n6427)
         );
  NAND2_X1 U7926 ( .A1(n9799), .A2(n6478), .ZN(n6425) );
  NAND2_X1 U7927 ( .A1(n9518), .A2(n6228), .ZN(n6424) );
  NAND2_X1 U7928 ( .A1(n6425), .A2(n6424), .ZN(n6426) );
  XNOR2_X1 U7929 ( .A(n6426), .B(n7389), .ZN(n6429) );
  XOR2_X1 U7930 ( .A(n6427), .B(n6429), .Z(n9423) );
  INV_X1 U7931 ( .A(n6427), .ZN(n6428) );
  NAND2_X1 U7932 ( .A1(n7926), .A2(n8096), .ZN(n6432) );
  OR2_X1 U7933 ( .A1(n5992), .A2(n7927), .ZN(n6431) );
  NAND2_X1 U7934 ( .A1(n9796), .A2(n6478), .ZN(n6445) );
  NAND2_X1 U7935 ( .A1(n6433), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n6439) );
  INV_X1 U7936 ( .A(n6436), .ZN(n6434) );
  NAND2_X1 U7937 ( .A1(n6434), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n6454) );
  INV_X1 U7938 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n6435) );
  NAND2_X1 U7939 ( .A1(n6436), .A2(n6435), .ZN(n6437) );
  NAND2_X1 U7940 ( .A1(n6454), .A2(n6437), .ZN(n9610) );
  OR2_X1 U7941 ( .A1(n6526), .A2(n9610), .ZN(n6438) );
  NAND2_X1 U7942 ( .A1(n6439), .A2(n6438), .ZN(n6443) );
  INV_X1 U7943 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8862) );
  NOR2_X1 U7944 ( .A1(n8017), .A2(n8862), .ZN(n6442) );
  INV_X1 U7945 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n6440) );
  NOR2_X1 U7946 ( .A1(n6123), .A2(n6440), .ZN(n6441) );
  NAND2_X1 U7947 ( .A1(n9627), .A2(n6193), .ZN(n6444) );
  NAND2_X1 U7948 ( .A1(n6445), .A2(n6444), .ZN(n6446) );
  XNOR2_X1 U7949 ( .A(n6446), .B(n7389), .ZN(n6447) );
  AOI22_X1 U7950 ( .A1(n9796), .A2(n6193), .B1(n6474), .B2(n9627), .ZN(n6448)
         );
  XNOR2_X1 U7951 ( .A(n6447), .B(n6448), .ZN(n9494) );
  INV_X1 U7952 ( .A(n6447), .ZN(n6449) );
  AOI22_X2 U7953 ( .A1(n9493), .A2(n9494), .B1(n6449), .B2(n6448), .ZN(n9390)
         );
  NAND2_X1 U7954 ( .A1(n9893), .A2(n8096), .ZN(n6451) );
  OR2_X1 U7955 ( .A1(n5992), .A2(n9895), .ZN(n6450) );
  NAND2_X1 U7956 ( .A1(n8011), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n6453) );
  INV_X1 U7957 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n8795) );
  OR2_X1 U7958 ( .A1(n8017), .A2(n8795), .ZN(n6452) );
  NAND2_X1 U7959 ( .A1(n6453), .A2(n6452), .ZN(n6459) );
  INV_X1 U7960 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8883) );
  NAND2_X1 U7961 ( .A1(n6454), .A2(n8883), .ZN(n6455) );
  NAND2_X1 U7962 ( .A1(n6468), .A2(n6455), .ZN(n9591) );
  NOR2_X1 U7963 ( .A1(n6526), .A2(n9591), .ZN(n6458) );
  INV_X1 U7964 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n6456) );
  NOR2_X1 U7965 ( .A1(n8013), .A2(n6456), .ZN(n6457) );
  AOI22_X1 U7966 ( .A1(n9789), .A2(n6478), .B1(n6193), .B2(n9576), .ZN(n6460)
         );
  XOR2_X1 U7967 ( .A(n7389), .B(n6460), .Z(n9388) );
  AND2_X1 U7968 ( .A1(n6474), .A2(n9576), .ZN(n6461) );
  AOI21_X1 U7969 ( .B1(n9789), .B2(n6193), .A(n6461), .ZN(n9387) );
  INV_X1 U7970 ( .A(n9387), .ZN(n6462) );
  OAI21_X1 U7971 ( .B1(n9390), .B2(n9388), .A(n6462), .ZN(n6510) );
  NAND2_X1 U7972 ( .A1(n9888), .A2(n8096), .ZN(n6464) );
  OR2_X1 U7973 ( .A1(n5992), .A2(n9890), .ZN(n6463) );
  NAND2_X1 U7974 ( .A1(n9783), .A2(n6228), .ZN(n6476) );
  NAND2_X1 U7975 ( .A1(n8011), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n6473) );
  INV_X1 U7976 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n6465) );
  OR2_X1 U7977 ( .A1(n8017), .A2(n6465), .ZN(n6472) );
  INV_X1 U7978 ( .A(n6468), .ZN(n6466) );
  NAND2_X1 U7979 ( .A1(n6466), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8389) );
  INV_X1 U7980 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U7981 ( .A1(n6468), .A2(n6467), .ZN(n6469) );
  NAND2_X1 U7982 ( .A1(n8389), .A2(n6469), .ZN(n9582) );
  INV_X1 U7983 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9583) );
  OR2_X1 U7984 ( .A1(n8013), .A2(n9583), .ZN(n6470) );
  NAND4_X1 U7985 ( .A1(n6473), .A2(n6472), .A3(n6471), .A4(n6470), .ZN(n9517)
         );
  NAND2_X1 U7986 ( .A1(n6474), .A2(n9517), .ZN(n6475) );
  NAND2_X1 U7987 ( .A1(n6476), .A2(n6475), .ZN(n6477) );
  XNOR2_X1 U7988 ( .A(n6477), .B(n7389), .ZN(n6480) );
  AOI22_X1 U7989 ( .A1(n9783), .A2(n6478), .B1(n6193), .B2(n9517), .ZN(n6479)
         );
  XNOR2_X1 U7990 ( .A(n6480), .B(n6479), .ZN(n6508) );
  INV_X1 U7991 ( .A(n6508), .ZN(n6507) );
  NAND2_X1 U7992 ( .A1(n6481), .A2(n8236), .ZN(n6962) );
  OR2_X1 U7993 ( .A1(n6962), .A2(n8229), .ZN(n6484) );
  INV_X1 U7994 ( .A(n6485), .ZN(n7778) );
  INV_X1 U7995 ( .A(n6486), .ZN(n7923) );
  NAND3_X1 U7996 ( .A1(n7923), .A2(P1_B_REG_SCAN_IN), .A3(n7778), .ZN(n6487)
         );
  OR2_X1 U7997 ( .A1(n6648), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6490) );
  INV_X1 U7998 ( .A(n6488), .ZN(n7928) );
  NAND2_X1 U7999 ( .A1(n7928), .A2(n7778), .ZN(n6489) );
  OR2_X1 U8000 ( .A1(n6648), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6491) );
  NAND2_X1 U8001 ( .A1(n7928), .A2(n7923), .ZN(n6649) );
  NOR2_X1 U8002 ( .A1(P1_D_REG_3__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .ZN(
        n6495) );
  NOR4_X1 U8003 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_16__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n6494) );
  NOR4_X1 U8004 ( .A1(P1_D_REG_5__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6493) );
  NOR4_X1 U8005 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_4__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6492) );
  NAND4_X1 U8006 ( .A1(n6495), .A2(n6494), .A3(n6493), .A4(n6492), .ZN(n6501)
         );
  NOR4_X1 U8007 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_19__SCAN_IN), .ZN(n6499) );
  NOR4_X1 U8008 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_13__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_11__SCAN_IN), .ZN(n6498) );
  NOR4_X1 U8009 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6497) );
  NOR4_X1 U8010 ( .A1(P1_D_REG_20__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6496) );
  NAND4_X1 U8011 ( .A1(n6499), .A2(n6498), .A3(n6497), .A4(n6496), .ZN(n6500)
         );
  NOR2_X1 U8012 ( .A1(n6501), .A2(n6500), .ZN(n6502) );
  OR2_X1 U8013 ( .A1(n6648), .A2(n6502), .ZN(n6879) );
  AND3_X1 U8014 ( .A1(n9880), .A2(n7354), .A3(n6879), .ZN(n6518) );
  NAND2_X1 U8015 ( .A1(n6503), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6504) );
  XNOR2_X1 U8016 ( .A(n6504), .B(n4997), .ZN(n6541) );
  AND2_X1 U8017 ( .A1(n6541), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6505) );
  NAND2_X1 U8018 ( .A1(n6518), .A2(n8270), .ZN(n6523) );
  NOR2_X1 U8019 ( .A1(n6972), .A2(n6523), .ZN(n6506) );
  NAND2_X1 U8020 ( .A1(n6507), .A2(n9483), .ZN(n6511) );
  OR2_X1 U8021 ( .A1(n6510), .A2(n6511), .ZN(n6538) );
  NAND3_X1 U8022 ( .A1(n6510), .A2(n6509), .A3(n6512), .ZN(n6537) );
  INV_X1 U8023 ( .A(n7361), .ZN(n6515) );
  INV_X1 U8024 ( .A(n6518), .ZN(n6513) );
  AND2_X1 U8025 ( .A1(n6513), .A2(n8270), .ZN(n6514) );
  NAND2_X1 U8026 ( .A1(n6515), .A2(n6514), .ZN(n6521) );
  AND2_X1 U8027 ( .A1(n8266), .A2(n8229), .ZN(n6516) );
  AND2_X1 U8028 ( .A1(n6521), .A2(n6880), .ZN(n9455) );
  AND3_X1 U8029 ( .A1(n6517), .A2(n6539), .A3(n6541), .ZN(n6519) );
  OR2_X1 U8030 ( .A1(n9849), .A2(n6518), .ZN(n6760) );
  NAND2_X1 U8031 ( .A1(n6519), .A2(n6760), .ZN(n6520) );
  NAND2_X1 U8032 ( .A1(n6520), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6522) );
  OR2_X1 U8033 ( .A1(n6964), .A2(n5914), .ZN(n8272) );
  NOR2_X1 U8034 ( .A1(n8272), .A2(n6523), .ZN(n6532) );
  NAND2_X1 U8035 ( .A1(n6525), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6531) );
  NAND2_X1 U8036 ( .A1(n8011), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n6530) );
  OR2_X1 U8037 ( .A1(n6526), .A2(n8389), .ZN(n6529) );
  INV_X1 U8038 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n6527) );
  OR2_X1 U8039 ( .A1(n8013), .A2(n6527), .ZN(n6528) );
  NAND4_X1 U8040 ( .A1(n6531), .A2(n6530), .A3(n6529), .A4(n6528), .ZN(n9577)
         );
  AOI22_X1 U8041 ( .A1(n9507), .A2(n9577), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6534) );
  INV_X1 U8042 ( .A(n4498), .ZN(n6971) );
  NAND2_X1 U8043 ( .A1(n9495), .A2(n9576), .ZN(n6533) );
  OAI211_X1 U8044 ( .C1(n9510), .C2(n9582), .A(n6534), .B(n6533), .ZN(n6535)
         );
  AOI21_X1 U8045 ( .B1(n9783), .B2(n9512), .A(n6535), .ZN(n6536) );
  NAND4_X1 U8046 ( .A1(n6538), .A2(n6537), .A3(n4544), .A4(n6536), .ZN(
        P1_U3218) );
  INV_X1 U8047 ( .A(n6541), .ZN(n7713) );
  NOR2_X2 U8048 ( .A1(n6717), .A2(P1_U3084), .ZN(P1_U4006) );
  INV_X1 U8049 ( .A(n10400), .ZN(n6540) );
  NOR2_X2 U8050 ( .A1(n6767), .A2(n6540), .ZN(P2_U3966) );
  NAND2_X1 U8051 ( .A1(n6972), .A2(n6541), .ZN(n6542) );
  NAND2_X1 U8052 ( .A1(n6542), .A2(n6717), .ZN(n10016) );
  OR2_X1 U8053 ( .A1(n10016), .A2(n6543), .ZN(n6544) );
  NAND2_X1 U8054 ( .A1(n6544), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NAND2_X1 U8055 ( .A1(n8355), .A2(n6616), .ZN(n7215) );
  NAND3_X1 U8056 ( .A1(n7023), .A2(n7520), .A3(n10404), .ZN(n6545) );
  NAND2_X1 U8057 ( .A1(n7215), .A2(n6545), .ZN(n6566) );
  XNOR2_X1 U8058 ( .A(n6566), .B(n6546), .ZN(n8578) );
  NAND2_X1 U8059 ( .A1(n8629), .A2(n8431), .ZN(n7016) );
  INV_X1 U8060 ( .A(n7016), .ZN(n7019) );
  NAND2_X1 U8061 ( .A1(n7019), .A2(n8314), .ZN(n8425) );
  OR2_X1 U8062 ( .A1(n6566), .A2(n8431), .ZN(n6547) );
  AND2_X1 U8063 ( .A1(n8425), .A2(n6547), .ZN(n8506) );
  INV_X1 U8064 ( .A(n8578), .ZN(n6548) );
  NAND2_X1 U8065 ( .A1(n6549), .A2(n6548), .ZN(n6550) );
  NAND2_X1 U8066 ( .A1(n8582), .A2(n6550), .ZN(n6551) );
  INV_X2 U8067 ( .A(n6566), .ZN(n8313) );
  XNOR2_X1 U8068 ( .A(n8313), .B(n10408), .ZN(n6552) );
  NAND2_X1 U8069 ( .A1(n8626), .A2(n8314), .ZN(n6553) );
  XNOR2_X1 U8070 ( .A(n6552), .B(n6553), .ZN(n8577) );
  INV_X1 U8071 ( .A(n6552), .ZN(n6554) );
  NAND2_X1 U8072 ( .A1(n6554), .A2(n6553), .ZN(n6555) );
  XNOR2_X1 U8073 ( .A(n6566), .B(n7169), .ZN(n6557) );
  NAND2_X1 U8074 ( .A1(n6556), .A2(n6557), .ZN(n6560) );
  INV_X1 U8075 ( .A(n6556), .ZN(n6558) );
  INV_X1 U8076 ( .A(n6557), .ZN(n7120) );
  NAND2_X1 U8077 ( .A1(n6558), .A2(n7120), .ZN(n6559) );
  NAND2_X1 U8078 ( .A1(n6560), .A2(n6559), .ZN(n10248) );
  XNOR2_X1 U8079 ( .A(n8313), .B(n10414), .ZN(n6562) );
  NAND2_X1 U8080 ( .A1(n8624), .A2(n8314), .ZN(n6563) );
  XNOR2_X1 U8081 ( .A(n6562), .B(n6563), .ZN(n7130) );
  AND2_X1 U8082 ( .A1(n7130), .A2(n6560), .ZN(n6561) );
  INV_X1 U8083 ( .A(n6562), .ZN(n6564) );
  NAND2_X1 U8084 ( .A1(n6564), .A2(n6563), .ZN(n6565) );
  NAND2_X1 U8085 ( .A1(n7125), .A2(n6565), .ZN(n10283) );
  NOR2_X1 U8086 ( .A1(n7313), .A2(n8341), .ZN(n6567) );
  XNOR2_X1 U8087 ( .A(n8343), .B(n10285), .ZN(n6568) );
  NAND2_X1 U8088 ( .A1(n6567), .A2(n6568), .ZN(n10282) );
  NAND2_X1 U8089 ( .A1(n10283), .A2(n10282), .ZN(n6571) );
  INV_X1 U8090 ( .A(n6567), .ZN(n6570) );
  INV_X1 U8091 ( .A(n6568), .ZN(n6569) );
  NAND2_X1 U8092 ( .A1(n6570), .A2(n6569), .ZN(n10281) );
  NAND2_X1 U8093 ( .A1(n6571), .A2(n10281), .ZN(n7187) );
  NOR2_X1 U8094 ( .A1(n7301), .A2(n8341), .ZN(n6572) );
  XNOR2_X1 U8095 ( .A(n7302), .B(n8343), .ZN(n6573) );
  NAND2_X1 U8096 ( .A1(n6572), .A2(n6573), .ZN(n6576) );
  INV_X1 U8097 ( .A(n6572), .ZN(n6575) );
  INV_X1 U8098 ( .A(n6573), .ZN(n6574) );
  NAND2_X1 U8099 ( .A1(n6575), .A2(n6574), .ZN(n6577) );
  AND2_X1 U8100 ( .A1(n6576), .A2(n6577), .ZN(n7188) );
  NAND2_X1 U8101 ( .A1(n7187), .A2(n7188), .ZN(n7186) );
  NAND2_X1 U8102 ( .A1(n7186), .A2(n6577), .ZN(n7243) );
  XNOR2_X1 U8103 ( .A(n7458), .B(n8313), .ZN(n6579) );
  OR2_X1 U8104 ( .A1(n7444), .A2(n8341), .ZN(n6578) );
  XNOR2_X1 U8105 ( .A(n6579), .B(n6578), .ZN(n7242) );
  INV_X1 U8106 ( .A(n6578), .ZN(n6581) );
  INV_X1 U8107 ( .A(n6579), .ZN(n6580) );
  NAND2_X1 U8108 ( .A1(n6581), .A2(n6580), .ZN(n6582) );
  XNOR2_X1 U8109 ( .A(n10356), .B(n8313), .ZN(n6583) );
  NOR2_X1 U8110 ( .A1(n7453), .A2(n8341), .ZN(n6584) );
  XNOR2_X1 U8111 ( .A(n6583), .B(n6584), .ZN(n7329) );
  INV_X1 U8112 ( .A(n6583), .ZN(n6585) );
  AND2_X1 U8113 ( .A1(n6585), .A2(n6584), .ZN(n6586) );
  XNOR2_X1 U8114 ( .A(n10436), .B(n8343), .ZN(n6590) );
  INV_X1 U8115 ( .A(n6590), .ZN(n6588) );
  NOR2_X1 U8116 ( .A1(n7501), .A2(n8341), .ZN(n6589) );
  INV_X1 U8117 ( .A(n6589), .ZN(n6587) );
  NAND2_X1 U8118 ( .A1(n6588), .A2(n6587), .ZN(n7600) );
  NAND2_X1 U8119 ( .A1(n6590), .A2(n6589), .ZN(n7598) );
  NAND2_X1 U8120 ( .A1(n7600), .A2(n7598), .ZN(n6591) );
  XNOR2_X1 U8121 ( .A(n7599), .B(n6591), .ZN(n6613) );
  AND2_X2 U8122 ( .A1(n5844), .A2(n7021), .ZN(n10444) );
  INV_X1 U8123 ( .A(n6623), .ZN(n6656) );
  NAND2_X1 U8124 ( .A1(n8427), .A2(n6656), .ZN(n6766) );
  NOR2_X1 U8125 ( .A1(n10444), .A2(n6766), .ZN(n6612) );
  NOR4_X1 U8126 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_12__SCAN_IN), .A3(
        P2_D_REG_14__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6595) );
  NOR4_X1 U8127 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_5__SCAN_IN), .A3(
        P2_D_REG_6__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6594) );
  NOR4_X1 U8128 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_24__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_29__SCAN_IN), .ZN(n6593) );
  NOR4_X1 U8129 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n6592) );
  NAND4_X1 U8130 ( .A1(n6595), .A2(n6594), .A3(n6593), .A4(n6592), .ZN(n6603)
         );
  NOR2_X1 U8131 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_15__SCAN_IN), .ZN(
        n6599) );
  NOR4_X1 U8132 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), .A3(
        P2_D_REG_17__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6598) );
  NOR4_X1 U8133 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n6597) );
  NOR4_X1 U8134 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_31__SCAN_IN), .A3(
        P2_D_REG_30__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6596) );
  NAND4_X1 U8135 ( .A1(n6599), .A2(n6598), .A3(n6597), .A4(n6596), .ZN(n6602)
         );
  INV_X1 U8136 ( .A(n6606), .ZN(n7922) );
  XNOR2_X1 U8137 ( .A(n7799), .B(P2_B_REG_SCAN_IN), .ZN(n6600) );
  NAND2_X1 U8138 ( .A1(n7922), .A2(n6600), .ZN(n6601) );
  OAI21_X1 U8139 ( .B1(n6603), .B2(n6602), .A(n10384), .ZN(n7011) );
  INV_X1 U8140 ( .A(n6607), .ZN(n7931) );
  AND2_X1 U8141 ( .A1(n7799), .A2(n7931), .ZN(n10397) );
  INV_X1 U8142 ( .A(n10397), .ZN(n6605) );
  INV_X1 U8143 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10396) );
  NAND2_X1 U8144 ( .A1(n10384), .A2(n10396), .ZN(n6604) );
  NAND2_X1 U8145 ( .A1(n6605), .A2(n6604), .ZN(n7209) );
  INV_X1 U8146 ( .A(n7209), .ZN(n7034) );
  INV_X1 U8147 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10399) );
  NAND2_X1 U8148 ( .A1(n10384), .A2(n10399), .ZN(n6609) );
  NOR2_X1 U8149 ( .A1(n6607), .A2(n6606), .ZN(n10401) );
  INV_X1 U8150 ( .A(n10401), .ZN(n6608) );
  AND2_X1 U8151 ( .A1(n6609), .A2(n6608), .ZN(n7210) );
  AND2_X1 U8152 ( .A1(n7034), .A2(n7210), .ZN(n6610) );
  NAND2_X1 U8153 ( .A1(n7011), .A2(n6610), .ZN(n6622) );
  INV_X1 U8154 ( .A(n6622), .ZN(n6611) );
  NOR2_X1 U8155 ( .A1(n6613), .A2(n10246), .ZN(n6628) );
  AND2_X1 U8156 ( .A1(n10444), .A2(n8427), .ZN(n6617) );
  NAND2_X1 U8157 ( .A1(n6622), .A2(n7213), .ZN(n8430) );
  AND2_X1 U8158 ( .A1(n10436), .A2(n10286), .ZN(n6627) );
  NAND2_X1 U8159 ( .A1(n5844), .A2(n6623), .ZN(n8428) );
  AND3_X1 U8160 ( .A1(n8428), .A2(n6618), .A3(n6767), .ZN(n6619) );
  NAND2_X1 U8161 ( .A1(n8430), .A2(n6619), .ZN(n6620) );
  NOR2_X1 U8162 ( .A1(n10292), .A2(n7460), .ZN(n6626) );
  OR2_X1 U8163 ( .A1(n5844), .A2(n10385), .ZN(n6621) );
  NAND2_X1 U8164 ( .A1(n10279), .A2(n10368), .ZN(n10260) );
  INV_X1 U8165 ( .A(n7453), .ZN(n8622) );
  NAND2_X1 U8166 ( .A1(n10257), .A2(n8622), .ZN(n6624) );
  NAND2_X1 U8167 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n6811) );
  OAI211_X1 U8168 ( .C1(n7736), .C2(n10260), .A(n6624), .B(n6811), .ZN(n6625)
         );
  OR4_X1 U8169 ( .A1(n6628), .A2(n6627), .A3(n6626), .A4(n6625), .ZN(P2_U3233)
         );
  AND2_X1 U8170 ( .A1(n4497), .A2(P1_U3084), .ZN(n9892) );
  INV_X2 U8171 ( .A(n9892), .ZN(n9886) );
  OAI222_X1 U8172 ( .A1(n9891), .A2(n6629), .B1(n9886), .B2(n6632), .C1(
        P1_U3084), .C2(n6868), .ZN(P1_U3352) );
  OAI222_X1 U8173 ( .A1(n9891), .A2(n6630), .B1(n9886), .B2(n6635), .C1(
        P1_U3084), .C2(n6886), .ZN(P1_U3351) );
  OAI222_X1 U8174 ( .A1(n9891), .A2(n6631), .B1(n9886), .B2(n6638), .C1(
        P1_U3084), .C2(n6831), .ZN(P1_U3350) );
  NOR2_X1 U8175 ( .A1(n4583), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9372) );
  INV_X2 U8176 ( .A(n9372), .ZN(n9382) );
  AND2_X1 U8177 ( .A1(n4583), .A2(P2_U3152), .ZN(n9378) );
  INV_X2 U8178 ( .A(n9378), .ZN(n9376) );
  OAI222_X1 U8179 ( .A1(n9382), .A2(n6633), .B1(n9376), .B2(n6632), .C1(n6861), 
        .C2(P2_U3152), .ZN(P2_U3357) );
  OAI222_X1 U8180 ( .A1(n6636), .A2(P2_U3152), .B1(n9376), .B2(n6635), .C1(
        n6634), .C2(n9382), .ZN(P2_U3356) );
  OAI222_X1 U8181 ( .A1(n6639), .A2(P2_U3152), .B1(n9376), .B2(n6638), .C1(
        n6637), .C2(n9382), .ZN(P2_U3355) );
  OAI222_X1 U8182 ( .A1(n9891), .A2(n6640), .B1(n9886), .B2(n6642), .C1(
        P1_U3084), .C2(n10027), .ZN(P1_U3349) );
  OAI222_X1 U8183 ( .A1(n6848), .A2(P2_U3152), .B1(n9376), .B2(n6642), .C1(
        n6641), .C2(n9382), .ZN(P2_U3354) );
  INV_X1 U8184 ( .A(n6643), .ZN(n6646) );
  INV_X1 U8185 ( .A(n9891), .ZN(n9882) );
  AOI22_X1 U8186 ( .A1(n10039), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n9882), .ZN(n6644) );
  OAI21_X1 U8187 ( .B1(n6646), .B2(n9886), .A(n6644), .ZN(P1_U3348) );
  OAI222_X1 U8188 ( .A1(n6647), .A2(P2_U3152), .B1(n9376), .B2(n6646), .C1(
        n6645), .C2(n9382), .ZN(P2_U3353) );
  INV_X1 U8189 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6651) );
  INV_X1 U8190 ( .A(n10193), .ZN(n10192) );
  OAI21_X1 U8191 ( .B1(n10192), .B2(P1_D_REG_1__SCAN_IN), .A(n6649), .ZN(n6650) );
  OAI21_X1 U8192 ( .B1(n8270), .B2(n6651), .A(n6650), .ZN(P1_U3441) );
  INV_X1 U8193 ( .A(n6652), .ZN(n6654) );
  AOI22_X1 U8194 ( .A1(n6815), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n9372), .ZN(n6653) );
  OAI21_X1 U8195 ( .B1(n6654), .B2(n9376), .A(n6653), .ZN(P2_U3352) );
  INV_X1 U8196 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6655) );
  INV_X1 U8197 ( .A(n6727), .ZN(n6698) );
  OAI222_X1 U8198 ( .A1(n9891), .A2(n6655), .B1(n9886), .B2(n6654), .C1(
        P1_U3084), .C2(n6698), .ZN(P1_U3347) );
  OAI21_X1 U8199 ( .B1(n10385), .B2(n6656), .A(n6780), .ZN(n6658) );
  NAND2_X1 U8200 ( .A1(n10385), .A2(n7709), .ZN(n6657) );
  NAND2_X1 U8201 ( .A1(n6658), .A2(n6657), .ZN(n10304) );
  INV_X1 U8202 ( .A(n10304), .ZN(n10328) );
  NOR2_X1 U8203 ( .A1(n10328), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U8204 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6660) );
  INV_X1 U8205 ( .A(n6659), .ZN(n6661) );
  INV_X1 U8206 ( .A(n6749), .ZN(n6704) );
  OAI222_X1 U8207 ( .A1(n9891), .A2(n6660), .B1(n9886), .B2(n6661), .C1(
        P1_U3084), .C2(n6704), .ZN(P1_U3346) );
  INV_X1 U8208 ( .A(n10316), .ZN(n6818) );
  INV_X1 U8209 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n8786) );
  OAI222_X1 U8210 ( .A1(n6818), .A2(P2_U3152), .B1(n9376), .B2(n6661), .C1(
        n8786), .C2(n9382), .ZN(P2_U3351) );
  INV_X1 U8211 ( .A(n8634), .ZN(n6820) );
  INV_X1 U8212 ( .A(n6662), .ZN(n6664) );
  OAI222_X1 U8213 ( .A1(n6820), .A2(P2_U3152), .B1(n9376), .B2(n6664), .C1(
        n6663), .C2(n9382), .ZN(P2_U3350) );
  INV_X1 U8214 ( .A(n10051), .ZN(n6747) );
  OAI222_X1 U8215 ( .A1(n9891), .A2(n6665), .B1(n9886), .B2(n6664), .C1(
        P1_U3084), .C2(n6747), .ZN(P1_U3345) );
  INV_X1 U8216 ( .A(n6666), .ZN(n6668) );
  AOI22_X1 U8217 ( .A1(n6992), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n9372), .ZN(n6667) );
  OAI21_X1 U8218 ( .B1(n6668), .B2(n9376), .A(n6667), .ZN(P2_U3349) );
  INV_X1 U8219 ( .A(n6746), .ZN(n10073) );
  OAI222_X1 U8220 ( .A1(n9886), .A2(n6668), .B1(n10073), .B2(P1_U3084), .C1(
        n8761), .C2(n9891), .ZN(P1_U3344) );
  INV_X1 U8221 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6671) );
  INV_X1 U8222 ( .A(n6669), .ZN(n8673) );
  NAND2_X1 U8223 ( .A1(n8673), .A2(P2_U3966), .ZN(n6670) );
  OAI21_X1 U8224 ( .B1(P2_U3966), .B2(n6671), .A(n6670), .ZN(P2_U3583) );
  INV_X1 U8225 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6675) );
  NAND2_X1 U8226 ( .A1(n8011), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6674) );
  INV_X1 U8227 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n6672) );
  OR2_X1 U8228 ( .A1(n8013), .A2(n6672), .ZN(n6673) );
  OAI211_X1 U8229 ( .C1(n8017), .C2(n6675), .A(n6674), .B(n6673), .ZN(n8360)
         );
  NAND2_X1 U8230 ( .A1(n8360), .A2(P1_U4006), .ZN(n6676) );
  OAI21_X1 U8231 ( .B1(P1_U4006), .B2(n5659), .A(n6676), .ZN(P1_U3586) );
  INV_X1 U8232 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6679) );
  NAND2_X1 U8233 ( .A1(n6677), .A2(P1_U4006), .ZN(n6678) );
  OAI21_X1 U8234 ( .B1(P1_U4006), .B2(n6679), .A(n6678), .ZN(P1_U3555) );
  INV_X1 U8235 ( .A(n6680), .ZN(n6684) );
  AOI22_X1 U8236 ( .A1(n10329), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n9372), .ZN(n6681) );
  OAI21_X1 U8237 ( .B1(n6684), .B2(n9376), .A(n6681), .ZN(P2_U3348) );
  INV_X1 U8238 ( .A(n6682), .ZN(n6687) );
  INV_X1 U8239 ( .A(n7113), .ZN(n6903) );
  OAI222_X1 U8240 ( .A1(n9886), .A2(n6687), .B1(n6903), .B2(P1_U3084), .C1(
        n6683), .C2(n9891), .ZN(P1_U3342) );
  INV_X1 U8241 ( .A(n6907), .ZN(n6743) );
  OAI222_X1 U8242 ( .A1(n9891), .A2(n6685), .B1(n6743), .B2(P1_U3084), .C1(
        n9886), .C2(n6684), .ZN(P1_U3343) );
  INV_X1 U8243 ( .A(n7061), .ZN(n7068) );
  OAI222_X1 U8244 ( .A1(P2_U3152), .A2(n7068), .B1(n9376), .B2(n6687), .C1(
        n6686), .C2(n9382), .ZN(P2_U3347) );
  NOR2_X1 U8245 ( .A1(n6727), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6699) );
  NAND2_X1 U8246 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n10039), .ZN(n6696) );
  MUX2_X1 U8247 ( .A(P1_REG1_REG_5__SCAN_IN), .B(n6688), .S(n10039), .Z(n10045) );
  MUX2_X1 U8248 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6695), .S(n10027), .Z(n10031) );
  OR2_X1 U8249 ( .A1(n6868), .A2(n6689), .ZN(n6691) );
  NAND2_X1 U8250 ( .A1(n6868), .A2(n6689), .ZN(n6690) );
  AND2_X1 U8251 ( .A1(n6691), .A2(n6690), .ZN(n6871) );
  NAND2_X1 U8252 ( .A1(n6871), .A2(n6870), .ZN(n6869) );
  NAND2_X1 U8253 ( .A1(n6869), .A2(n6691), .ZN(n6884) );
  XNOR2_X1 U8254 ( .A(n6886), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n6885) );
  NOR2_X1 U8255 ( .A1(n6886), .A2(n8774), .ZN(n6692) );
  AOI21_X1 U8256 ( .B1(n6884), .B2(n6885), .A(n6692), .ZN(n6829) );
  MUX2_X1 U8257 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n6694), .S(n6831), .Z(n6828)
         );
  NOR2_X1 U8258 ( .A1(n6829), .A2(n6828), .ZN(n6827) );
  INV_X1 U8259 ( .A(n6827), .ZN(n6693) );
  OAI21_X1 U8260 ( .B1(n6831), .B2(n6694), .A(n6693), .ZN(n10032) );
  NOR2_X1 U8261 ( .A1(n10031), .A2(n10032), .ZN(n10030) );
  AOI21_X1 U8262 ( .B1(n10027), .B2(n6695), .A(n10030), .ZN(n10046) );
  NAND2_X1 U8263 ( .A1(n10045), .A2(n10046), .ZN(n10044) );
  NAND2_X1 U8264 ( .A1(n6696), .A2(n10044), .ZN(n6726) );
  INV_X1 U8265 ( .A(n6699), .ZN(n6697) );
  OAI21_X1 U8266 ( .B1(n6032), .B2(n6698), .A(n6697), .ZN(n6725) );
  NOR2_X1 U8267 ( .A1(n6726), .A2(n6725), .ZN(n6724) );
  NOR2_X1 U8268 ( .A1(n6699), .A2(n6724), .ZN(n6701) );
  AOI22_X1 U8269 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n6704), .B1(n6749), .B2(
        n6051), .ZN(n6700) );
  NOR2_X1 U8270 ( .A1(n6701), .A2(n6700), .ZN(n6740) );
  AOI21_X1 U8271 ( .B1(n6701), .B2(n6700), .A(n6740), .ZN(n6723) );
  OR2_X1 U8272 ( .A1(n4498), .A2(P1_U3084), .ZN(n10011) );
  OR2_X1 U8273 ( .A1(n10016), .A2(n10011), .ZN(n6702) );
  INV_X1 U8274 ( .A(n8271), .ZN(n8359) );
  INV_X1 U8275 ( .A(n6702), .ZN(n6703) );
  NAND2_X1 U8276 ( .A1(n6703), .A2(n8359), .ZN(n10142) );
  AOI22_X1 U8277 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n6749), .B1(n6704), .B2(
        n7530), .ZN(n6714) );
  MUX2_X1 U8278 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n7359), .S(n6727), .Z(n6734)
         );
  OR2_X1 U8279 ( .A1(n10039), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n6711) );
  NOR2_X1 U8280 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n10039), .ZN(n6705) );
  AOI21_X1 U8281 ( .B1(n10039), .B2(P1_REG2_REG_5__SCAN_IN), .A(n6705), .ZN(
        n10042) );
  XNOR2_X1 U8282 ( .A(n6868), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n6866) );
  INV_X1 U8283 ( .A(n6896), .ZN(n6865) );
  NAND2_X1 U8284 ( .A1(n6866), .A2(n6865), .ZN(n6864) );
  INV_X1 U8285 ( .A(n6868), .ZN(n6706) );
  NAND2_X1 U8286 ( .A1(n6706), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6707) );
  NAND2_X1 U8287 ( .A1(n6864), .A2(n6707), .ZN(n6887) );
  XNOR2_X1 U8288 ( .A(n6886), .B(P1_REG2_REG_2__SCAN_IN), .ZN(n6888) );
  AND2_X1 U8289 ( .A1(n6887), .A2(n6888), .ZN(n6889) );
  INV_X1 U8290 ( .A(n6886), .ZN(n6708) );
  MUX2_X1 U8291 ( .A(n5920), .B(P1_REG2_REG_3__SCAN_IN), .S(n6831), .Z(n6836)
         );
  XNOR2_X1 U8292 ( .A(n10027), .B(n6709), .ZN(n10023) );
  OR2_X1 U8293 ( .A1(n10022), .A2(n10023), .ZN(n10024) );
  NAND2_X1 U8294 ( .A1(n10027), .A2(n6709), .ZN(n6710) );
  NAND2_X1 U8295 ( .A1(n10024), .A2(n6710), .ZN(n10041) );
  NAND2_X1 U8296 ( .A1(n10042), .A2(n10041), .ZN(n10040) );
  AND2_X1 U8297 ( .A1(n6711), .A2(n10040), .ZN(n6733) );
  NAND2_X1 U8298 ( .A1(n6727), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6712) );
  OAI21_X1 U8299 ( .B1(n6714), .B2(n6713), .A(n6748), .ZN(n6721) );
  INV_X1 U8300 ( .A(n10016), .ZN(n9554) );
  OR2_X1 U8301 ( .A1(n8271), .A2(P1_U3084), .ZN(n10010) );
  INV_X1 U8302 ( .A(n10010), .ZN(n9555) );
  AND2_X1 U8303 ( .A1(n9555), .A2(n4498), .ZN(n6715) );
  NAND2_X1 U8304 ( .A1(n10148), .A2(n6749), .ZN(n6716) );
  NAND2_X1 U8305 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7179) );
  NAND2_X1 U8306 ( .A1(n6716), .A2(n7179), .ZN(n6720) );
  INV_X1 U8307 ( .A(n6717), .ZN(n6718) );
  INV_X1 U8308 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n8831) );
  NOR2_X1 U8309 ( .A1(n10157), .A2(n8831), .ZN(n6719) );
  AOI211_X1 U8310 ( .C1(n10058), .C2(n6721), .A(n6720), .B(n6719), .ZN(n6722)
         );
  OAI21_X1 U8311 ( .B1(n6723), .B2(n10154), .A(n6722), .ZN(P1_U3248) );
  INV_X1 U8312 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n6737) );
  AOI21_X1 U8313 ( .B1(n6726), .B2(n6725), .A(n6724), .ZN(n6730) );
  NOR2_X1 U8314 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8893), .ZN(n7136) );
  INV_X1 U8315 ( .A(n7136), .ZN(n6729) );
  NAND2_X1 U8316 ( .A1(n10148), .A2(n6727), .ZN(n6728) );
  OAI211_X1 U8317 ( .C1(n10154), .C2(n6730), .A(n6729), .B(n6728), .ZN(n6731)
         );
  INV_X1 U8318 ( .A(n6731), .ZN(n6736) );
  OAI211_X1 U8319 ( .C1(n6734), .C2(n6733), .A(n10058), .B(n6732), .ZN(n6735)
         );
  OAI211_X1 U8320 ( .C1(n6737), .C2(n10157), .A(n6736), .B(n6735), .ZN(
        P1_U3247) );
  NAND2_X1 U8321 ( .A1(n9113), .A2(P2_U3966), .ZN(n6738) );
  OAI21_X1 U8322 ( .B1(P2_U3966), .B2(n7715), .A(n6738), .ZN(P2_U3575) );
  NOR2_X1 U8323 ( .A1(n6746), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6741) );
  INV_X1 U8324 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10241) );
  MUX2_X1 U8325 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10241), .S(n10051), .Z(
        n10060) );
  NOR2_X1 U8326 ( .A1(n6749), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6739) );
  NOR2_X1 U8327 ( .A1(n6740), .A2(n6739), .ZN(n10061) );
  NAND2_X1 U8328 ( .A1(n10060), .A2(n10061), .ZN(n10059) );
  OAI21_X1 U8329 ( .B1(n10241), .B2(n6747), .A(n10059), .ZN(n10068) );
  AOI22_X1 U8330 ( .A1(n6746), .A2(n6094), .B1(P1_REG1_REG_9__SCAN_IN), .B2(
        n10073), .ZN(n10067) );
  NOR2_X1 U8331 ( .A1(n10068), .A2(n10067), .ZN(n10066) );
  NOR2_X1 U8332 ( .A1(n6741), .A2(n10066), .ZN(n6745) );
  NOR2_X1 U8333 ( .A1(n6907), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6902) );
  INV_X1 U8334 ( .A(n6902), .ZN(n6742) );
  OAI21_X1 U8335 ( .B1(n6125), .B2(n6743), .A(n6742), .ZN(n6744) );
  NOR2_X1 U8336 ( .A1(n6745), .A2(n6744), .ZN(n6901) );
  AOI21_X1 U8337 ( .B1(n6745), .B2(n6744), .A(n6901), .ZN(n6759) );
  INV_X1 U8338 ( .A(n10157), .ZN(n10052) );
  INV_X1 U8339 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7480) );
  XNOR2_X1 U8340 ( .A(n6907), .B(n7480), .ZN(n6753) );
  NAND2_X1 U8341 ( .A1(n6746), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6751) );
  OAI21_X1 U8342 ( .B1(n6746), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6751), .ZN(
        n10071) );
  INV_X1 U8343 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n8772) );
  AOI22_X1 U8344 ( .A1(n10051), .A2(P1_REG2_REG_8__SCAN_IN), .B1(n8772), .B2(
        n6747), .ZN(n10055) );
  NAND2_X1 U8345 ( .A1(n10055), .A2(n10056), .ZN(n10054) );
  OAI21_X1 U8346 ( .B1(n10051), .B2(P1_REG2_REG_8__SCAN_IN), .A(n10054), .ZN(
        n10072) );
  NOR2_X1 U8347 ( .A1(n10071), .A2(n10072), .ZN(n10070) );
  INV_X1 U8348 ( .A(n10070), .ZN(n6750) );
  NAND2_X1 U8349 ( .A1(n6751), .A2(n6750), .ZN(n6752) );
  NAND2_X1 U8350 ( .A1(n6753), .A2(n6752), .ZN(n6909) );
  OAI21_X1 U8351 ( .B1(n6753), .B2(n6752), .A(n6909), .ZN(n6756) );
  NOR2_X1 U8352 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8792), .ZN(n7542) );
  INV_X1 U8353 ( .A(n7542), .ZN(n6755) );
  NAND2_X1 U8354 ( .A1(n10148), .A2(n6907), .ZN(n6754) );
  OAI211_X1 U8355 ( .C1(n10142), .C2(n6756), .A(n6755), .B(n6754), .ZN(n6757)
         );
  AOI21_X1 U8356 ( .B1(n10052), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n6757), .ZN(
        n6758) );
  OAI21_X1 U8357 ( .B1(n6759), .B2(n10154), .A(n6758), .ZN(P1_U3251) );
  NAND2_X1 U8358 ( .A1(n9455), .A2(n6760), .ZN(n6945) );
  AOI22_X1 U8359 ( .A1(n9512), .A2(n7369), .B1(n6945), .B2(
        P1_REG3_REG_0__SCAN_IN), .ZN(n6765) );
  OAI21_X1 U8360 ( .B1(n6761), .B2(n6762), .A(n6763), .ZN(n6895) );
  AOI22_X1 U8361 ( .A1(n6895), .A2(n9483), .B1(n9507), .B2(n9531), .ZN(n6764)
         );
  NAND2_X1 U8362 ( .A1(n6765), .A2(n6764), .ZN(P1_U3230) );
  OR2_X1 U8363 ( .A1(n6797), .A2(P2_U3152), .ZN(n9379) );
  OAI211_X1 U8364 ( .C1(n6767), .C2(n9379), .A(n6766), .B(n7709), .ZN(n6782)
         );
  NAND2_X1 U8365 ( .A1(n6782), .A2(n6780), .ZN(n6768) );
  INV_X2 U8366 ( .A(P2_U3966), .ZN(n8628) );
  NAND2_X1 U8367 ( .A1(n6768), .A2(n8628), .ZN(n6799) );
  INV_X1 U8368 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U8369 ( .A1(n9900), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6778) );
  MUX2_X1 U8370 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6769), .S(n9900), .Z(n9902)
         );
  NAND2_X1 U8371 ( .A1(n10306), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6775) );
  MUX2_X1 U8372 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6770), .S(n10306), .Z(n10308) );
  INV_X1 U8373 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n8857) );
  MUX2_X1 U8374 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n8857), .S(n6861), .Z(n6851)
         );
  INV_X1 U8375 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n6849) );
  NOR3_X1 U8376 ( .A1(n6851), .A2(n6771), .A3(n6849), .ZN(n6850) );
  INV_X1 U8377 ( .A(n6850), .ZN(n6772) );
  OAI21_X1 U8378 ( .B1(n8857), .B2(n6861), .A(n6772), .ZN(n9913) );
  MUX2_X1 U8379 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6773), .S(n9910), .Z(n9912)
         );
  NAND2_X1 U8380 ( .A1(n9913), .A2(n9912), .ZN(n9911) );
  NAND2_X1 U8381 ( .A1(n9910), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6774) );
  NAND2_X1 U8382 ( .A1(n9911), .A2(n6774), .ZN(n10309) );
  NAND2_X1 U8383 ( .A1(n10308), .A2(n10309), .ZN(n10307) );
  AND2_X1 U8384 ( .A1(n6775), .A2(n10307), .ZN(n6841) );
  MUX2_X1 U8385 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6777), .S(n6848), .Z(n6840)
         );
  NOR2_X1 U8386 ( .A1(n6841), .A2(n6840), .ZN(n6839) );
  INV_X1 U8387 ( .A(n6839), .ZN(n6776) );
  OAI21_X1 U8388 ( .B1(n6777), .B2(n6848), .A(n6776), .ZN(n9903) );
  NAND2_X1 U8389 ( .A1(n9902), .A2(n9903), .ZN(n9901) );
  NAND2_X1 U8390 ( .A1(n6778), .A2(n9901), .ZN(n6784) );
  MUX2_X1 U8391 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6779), .S(n6815), .Z(n6783)
         );
  AND2_X1 U8392 ( .A1(n6780), .A2(n9385), .ZN(n6781) );
  NAND2_X1 U8393 ( .A1(n6783), .A2(n6784), .ZN(n6806) );
  OAI211_X1 U8394 ( .C1(n6784), .C2(n6783), .A(n10336), .B(n6806), .ZN(n6785)
         );
  NAND2_X1 U8395 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n7191) );
  OAI211_X1 U8396 ( .C1(n10304), .C2(n6786), .A(n6785), .B(n7191), .ZN(n6787)
         );
  AOI21_X1 U8397 ( .B1(n6815), .B2(n10330), .A(n6787), .ZN(n6803) );
  NAND2_X1 U8398 ( .A1(n9900), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6795) );
  MUX2_X1 U8399 ( .A(n7235), .B(P2_REG2_REG_5__SCAN_IN), .S(n9900), .Z(n6788)
         );
  INV_X1 U8400 ( .A(n6788), .ZN(n9905) );
  INV_X1 U8401 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n6794) );
  NAND2_X1 U8402 ( .A1(n10306), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n6793) );
  MUX2_X1 U8403 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6789), .S(n10306), .Z(n10311) );
  NAND2_X1 U8404 ( .A1(n9910), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6792) );
  OAI21_X1 U8405 ( .B1(n6861), .B2(n6855), .A(n6856), .ZN(n9916) );
  MUX2_X1 U8406 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n6791), .S(n9910), .Z(n9915)
         );
  NAND2_X1 U8407 ( .A1(n9916), .A2(n9915), .ZN(n9914) );
  NAND2_X1 U8408 ( .A1(n6792), .A2(n9914), .ZN(n10312) );
  NAND2_X1 U8409 ( .A1(n10311), .A2(n10312), .ZN(n10310) );
  NAND2_X1 U8410 ( .A1(n6793), .A2(n10310), .ZN(n6845) );
  MUX2_X1 U8411 ( .A(n6794), .B(P2_REG2_REG_4__SCAN_IN), .S(n6848), .Z(n6844)
         );
  NAND2_X1 U8412 ( .A1(n6845), .A2(n6844), .ZN(n6843) );
  OAI21_X1 U8413 ( .B1(n6794), .B2(n6848), .A(n6843), .ZN(n9906) );
  NAND2_X1 U8414 ( .A1(n9905), .A2(n9906), .ZN(n9904) );
  NAND2_X1 U8415 ( .A1(n6795), .A2(n9904), .ZN(n6801) );
  MUX2_X1 U8416 ( .A(n5195), .B(P2_REG2_REG_6__SCAN_IN), .S(n6815), .Z(n6796)
         );
  INV_X1 U8417 ( .A(n6796), .ZN(n6800) );
  NOR2_X1 U8418 ( .A1(n6797), .A2(n9385), .ZN(n6798) );
  NAND2_X1 U8419 ( .A1(n6799), .A2(n6798), .ZN(n10295) );
  NAND2_X1 U8420 ( .A1(n6800), .A2(n6801), .ZN(n6816) );
  OAI211_X1 U8421 ( .C1(n6801), .C2(n6800), .A(n10332), .B(n6816), .ZN(n6802)
         );
  NAND2_X1 U8422 ( .A1(n6803), .A2(n6802), .ZN(P2_U3251) );
  INV_X1 U8423 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n6813) );
  MUX2_X1 U8424 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6804), .S(n8634), .Z(n8636)
         );
  MUX2_X1 U8425 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6805), .S(n10316), .Z(n10318) );
  NAND2_X1 U8426 ( .A1(n6815), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6807) );
  NAND2_X1 U8427 ( .A1(n6807), .A2(n6806), .ZN(n10319) );
  NAND2_X1 U8428 ( .A1(n10318), .A2(n10319), .ZN(n10317) );
  OAI21_X1 U8429 ( .B1(n6818), .B2(n6805), .A(n10317), .ZN(n8637) );
  NAND2_X1 U8430 ( .A1(n8636), .A2(n8637), .ZN(n8635) );
  OAI21_X1 U8431 ( .B1(n6820), .B2(n6804), .A(n8635), .ZN(n6810) );
  MUX2_X1 U8432 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n6808), .S(n6992), .Z(n6809)
         );
  NAND2_X1 U8433 ( .A1(n6809), .A2(n6810), .ZN(n6998) );
  OAI211_X1 U8434 ( .C1(n6810), .C2(n6809), .A(n10336), .B(n6998), .ZN(n6812)
         );
  OAI211_X1 U8435 ( .C1(n10304), .C2(n6813), .A(n6812), .B(n6811), .ZN(n6814)
         );
  AOI21_X1 U8436 ( .B1(n6992), .B2(n10330), .A(n6814), .ZN(n6824) );
  INV_X1 U8437 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6819) );
  MUX2_X1 U8438 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6819), .S(n8634), .Z(n8631)
         );
  MUX2_X1 U8439 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n7305), .S(n10316), .Z(n10321) );
  NAND2_X1 U8440 ( .A1(n6815), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n6817) );
  NAND2_X1 U8441 ( .A1(n6817), .A2(n6816), .ZN(n10322) );
  NAND2_X1 U8442 ( .A1(n10321), .A2(n10322), .ZN(n10320) );
  MUX2_X1 U8443 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7461), .S(n6992), .Z(n6821)
         );
  OAI211_X1 U8444 ( .C1(n6822), .C2(n6821), .A(n10332), .B(n6993), .ZN(n6823)
         );
  NAND2_X1 U8445 ( .A1(n6824), .A2(n6823), .ZN(P2_U3254) );
  INV_X1 U8446 ( .A(n6825), .ZN(n6862) );
  AOI22_X1 U8447 ( .A1(n10084), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9882), .ZN(n6826) );
  OAI21_X1 U8448 ( .B1(n6862), .B2(n9886), .A(n6826), .ZN(P1_U3341) );
  AOI211_X1 U8449 ( .C1(n6829), .C2(n6828), .A(n6827), .B(n10154), .ZN(n6833)
         );
  INV_X1 U8450 ( .A(n10148), .ZN(n10074) );
  INV_X1 U8451 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8923) );
  NOR2_X1 U8452 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n8923), .ZN(n6926) );
  INV_X1 U8453 ( .A(n6926), .ZN(n6830) );
  OAI21_X1 U8454 ( .B1(n10074), .B2(n6831), .A(n6830), .ZN(n6832) );
  NOR2_X1 U8455 ( .A1(n6833), .A2(n6832), .ZN(n6838) );
  OAI211_X1 U8456 ( .C1(n6836), .C2(n6835), .A(n10058), .B(n6834), .ZN(n6837)
         );
  OAI211_X1 U8457 ( .C1(n8859), .C2(n10157), .A(n6838), .B(n6837), .ZN(
        P1_U3244) );
  INV_X1 U8458 ( .A(n10330), .ZN(n10293) );
  AND2_X1 U8459 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7122) );
  AOI211_X1 U8460 ( .C1(n6841), .C2(n6840), .A(n6839), .B(n10294), .ZN(n6842)
         );
  AOI211_X1 U8461 ( .C1(n10328), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n7122), .B(
        n6842), .ZN(n6847) );
  OAI211_X1 U8462 ( .C1(n6845), .C2(n6844), .A(n10332), .B(n6843), .ZN(n6846)
         );
  OAI211_X1 U8463 ( .C1(n10293), .C2(n6848), .A(n6847), .B(n6846), .ZN(
        P2_U3249) );
  NOR2_X1 U8464 ( .A1(n4680), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6854) );
  OR2_X1 U8465 ( .A1(n6849), .A2(n6771), .ZN(n6852) );
  AOI211_X1 U8466 ( .C1(n6852), .C2(n6851), .A(n6850), .B(n10294), .ZN(n6853)
         );
  AOI211_X1 U8467 ( .C1(n10328), .C2(P2_ADDR_REG_1__SCAN_IN), .A(n6854), .B(
        n6853), .ZN(n6860) );
  AND2_X1 U8468 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(
        n6858) );
  MUX2_X1 U8469 ( .A(n6855), .B(P2_REG2_REG_1__SCAN_IN), .S(n6861), .Z(n6857)
         );
  OAI211_X1 U8470 ( .C1(n6858), .C2(n6857), .A(n10332), .B(n6856), .ZN(n6859)
         );
  OAI211_X1 U8471 ( .C1(n10293), .C2(n6861), .A(n6860), .B(n6859), .ZN(
        P2_U3246) );
  INV_X1 U8472 ( .A(n7075), .ZN(n7148) );
  OAI222_X1 U8473 ( .A1(n9382), .A2(n6863), .B1(n9376), .B2(n6862), .C1(n7148), 
        .C2(P2_U3152), .ZN(P2_U3346) );
  OAI211_X1 U8474 ( .C1(n6866), .C2(n6865), .A(n10058), .B(n6864), .ZN(n6867)
         );
  OAI21_X1 U8475 ( .B1(n10074), .B2(n6868), .A(n6867), .ZN(n6874) );
  OAI211_X1 U8476 ( .C1(n6871), .C2(n6870), .A(n10135), .B(n6869), .ZN(n6872)
         );
  OAI21_X1 U8477 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n7384), .A(n6872), .ZN(n6873) );
  AOI211_X1 U8478 ( .C1(n10052), .C2(P1_ADDR_REG_1__SCAN_IN), .A(n6874), .B(
        n6873), .ZN(n6875) );
  INV_X1 U8479 ( .A(n6875), .ZN(P1_U3242) );
  INV_X1 U8480 ( .A(n6962), .ZN(n6878) );
  INV_X1 U8481 ( .A(n9531), .ZN(n6973) );
  INV_X1 U8482 ( .A(n7369), .ZN(n7383) );
  INV_X1 U8483 ( .A(n7376), .ZN(n6876) );
  NAND2_X1 U8484 ( .A1(n6677), .A2(n7383), .ZN(n8240) );
  NAND2_X1 U8485 ( .A1(n6876), .A2(n8240), .ZN(n8119) );
  NAND3_X1 U8486 ( .A1(n8119), .A2(n8272), .A3(n6962), .ZN(n6877) );
  OAI21_X1 U8487 ( .B1(n6973), .B2(n10167), .A(n6877), .ZN(n7370) );
  AOI21_X1 U8488 ( .B1(n7369), .B2(n6878), .A(n7370), .ZN(n6958) );
  INV_X1 U8489 ( .A(n7354), .ZN(n6881) );
  OAI21_X1 U8490 ( .B1(n9862), .B2(n6483), .A(n6881), .ZN(n6882) );
  NAND2_X1 U8491 ( .A1(n10243), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6883) );
  OAI21_X1 U8492 ( .B1(n6958), .B2(n10243), .A(n6883), .ZN(P1_U3523) );
  INV_X1 U8493 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6900) );
  XOR2_X1 U8494 ( .A(n6885), .B(n6884), .Z(n6894) );
  OAI22_X1 U8495 ( .A1(n10074), .A2(n6886), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7548), .ZN(n6893) );
  INV_X1 U8496 ( .A(n6887), .ZN(n6891) );
  INV_X1 U8497 ( .A(n6888), .ZN(n6890) );
  AOI211_X1 U8498 ( .C1(n6891), .C2(n6890), .A(n6889), .B(n10142), .ZN(n6892)
         );
  AOI211_X1 U8499 ( .C1(n10135), .C2(n6894), .A(n6893), .B(n6892), .ZN(n6899)
         );
  MUX2_X1 U8500 ( .A(n6896), .B(n6895), .S(n8271), .Z(n6898) );
  NOR2_X1 U8501 ( .A1(n8271), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6897) );
  OR2_X1 U8502 ( .A1(n4498), .A2(n6897), .ZN(n10014) );
  NAND2_X1 U8503 ( .A1(n10014), .A2(n4694), .ZN(n10012) );
  OAI211_X1 U8504 ( .C1(n6898), .C2(n4498), .A(P1_U4006), .B(n10012), .ZN(
        n10036) );
  OAI211_X1 U8505 ( .C1(n6900), .C2(n10157), .A(n6899), .B(n10036), .ZN(
        P1_U3243) );
  NOR2_X1 U8506 ( .A1(n6902), .A2(n6901), .ZN(n6905) );
  INV_X1 U8507 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n10002) );
  AOI22_X1 U8508 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n6903), .B1(n7113), .B2(
        n10002), .ZN(n6904) );
  NOR2_X1 U8509 ( .A1(n6905), .A2(n6904), .ZN(n7101) );
  AOI21_X1 U8510 ( .B1(n6905), .B2(n6904), .A(n7101), .ZN(n6917) );
  NOR2_X1 U8511 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n7113), .ZN(n6906) );
  AOI21_X1 U8512 ( .B1(n7113), .B2(P1_REG2_REG_11__SCAN_IN), .A(n6906), .ZN(
        n6911) );
  NAND2_X1 U8513 ( .A1(n6907), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n6908) );
  AND2_X1 U8514 ( .A1(n6909), .A2(n6908), .ZN(n6910) );
  OAI21_X1 U8515 ( .B1(n6911), .B2(n6910), .A(n7112), .ZN(n6912) );
  INV_X1 U8516 ( .A(n6912), .ZN(n6914) );
  NOR2_X1 U8517 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6141), .ZN(n7641) );
  AOI21_X1 U8518 ( .B1(n10148), .B2(n7113), .A(n7641), .ZN(n6913) );
  OAI21_X1 U8519 ( .B1(n10142), .B2(n6914), .A(n6913), .ZN(n6915) );
  AOI21_X1 U8520 ( .B1(n10052), .B2(P1_ADDR_REG_11__SCAN_IN), .A(n6915), .ZN(
        n6916) );
  OAI21_X1 U8521 ( .B1(n6917), .B2(n10154), .A(n6916), .ZN(P1_U3252) );
  NAND2_X1 U8522 ( .A1(n6919), .A2(n6920), .ZN(n6924) );
  XNOR2_X1 U8523 ( .A(n6922), .B(n6921), .ZN(n6923) );
  XNOR2_X1 U8524 ( .A(n6924), .B(n6923), .ZN(n6931) );
  INV_X1 U8525 ( .A(n9483), .ZN(n9514) );
  INV_X1 U8526 ( .A(n9510), .ZN(n9466) );
  INV_X1 U8527 ( .A(n6925), .ZN(n7568) );
  NAND2_X1 U8528 ( .A1(n9512), .A2(n7564), .ZN(n6928) );
  AOI21_X1 U8529 ( .B1(n9507), .B2(n9529), .A(n6926), .ZN(n6927) );
  OAI211_X1 U8530 ( .C1(n7568), .C2(n9505), .A(n6928), .B(n6927), .ZN(n6929)
         );
  AOI21_X1 U8531 ( .B1(n8923), .B2(n9466), .A(n6929), .ZN(n6930) );
  OAI21_X1 U8532 ( .B1(n6931), .B2(n9514), .A(n6930), .ZN(P1_U3216) );
  INV_X1 U8533 ( .A(n6932), .ZN(n6934) );
  NAND2_X1 U8534 ( .A1(n6934), .A2(n6933), .ZN(n6936) );
  AOI22_X1 U8535 ( .A1(n6937), .A2(n6936), .B1(n4577), .B2(n6935), .ZN(n6941)
         );
  INV_X1 U8536 ( .A(n6677), .ZN(n7377) );
  INV_X1 U8537 ( .A(n9507), .ZN(n9486) );
  OAI22_X1 U8538 ( .A1(n7377), .A2(n9505), .B1(n9486), .B2(n7568), .ZN(n6939)
         );
  INV_X1 U8539 ( .A(n7386), .ZN(n10196) );
  NOR2_X1 U8540 ( .A1(n9492), .A2(n10196), .ZN(n6938) );
  AOI211_X1 U8541 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(n6945), .A(n6939), .B(
        n6938), .ZN(n6940) );
  OAI21_X1 U8542 ( .B1(n6941), .B2(n9514), .A(n6940), .ZN(P1_U3220) );
  INV_X1 U8543 ( .A(n7553), .ZN(n6963) );
  OAI21_X1 U8544 ( .B1(n6942), .B2(n4577), .A(n6919), .ZN(n6943) );
  NAND2_X1 U8545 ( .A1(n6943), .A2(n9483), .ZN(n6947) );
  OAI22_X1 U8546 ( .A1(n6973), .A2(n9505), .B1(n9486), .B2(n7084), .ZN(n6944)
         );
  AOI21_X1 U8547 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n6945), .A(n6944), .ZN(
        n6946) );
  OAI211_X1 U8548 ( .C1(n6963), .C2(n9492), .A(n6947), .B(n6946), .ZN(P1_U3235) );
  INV_X1 U8549 ( .A(n6948), .ZN(n6952) );
  INV_X1 U8550 ( .A(n10097), .ZN(n7105) );
  OAI222_X1 U8551 ( .A1(n9886), .A2(n6952), .B1(n7105), .B2(P1_U3084), .C1(
        n6949), .C2(n9891), .ZN(P1_U3340) );
  NAND2_X1 U8552 ( .A1(n9677), .A2(P1_U4006), .ZN(n6950) );
  OAI21_X1 U8553 ( .B1(n9527), .B2(n7711), .A(n6950), .ZN(P1_U3578) );
  INV_X1 U8554 ( .A(n7338), .ZN(n7345) );
  OAI222_X1 U8555 ( .A1(P2_U3152), .A2(n7345), .B1(n9376), .B2(n6952), .C1(
        n6951), .C2(n9382), .ZN(P2_U3345) );
  INV_X1 U8556 ( .A(n6953), .ZN(n6981) );
  OAI222_X1 U8557 ( .A1(n9886), .A2(n6981), .B1(n9541), .B2(P1_U3084), .C1(
        n6954), .C2(n9891), .ZN(P1_U3339) );
  INV_X1 U8558 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6956) );
  OR2_X1 U8559 ( .A1(n10236), .A2(n6956), .ZN(n6957) );
  OAI21_X1 U8560 ( .B1(n6958), .B2(n10234), .A(n6957), .ZN(P1_U3454) );
  INV_X1 U8561 ( .A(n9862), .ZN(n10233) );
  AND2_X1 U8562 ( .A1(n6677), .A2(n7369), .ZN(n7375) );
  XNOR2_X2 U8563 ( .A(n9531), .B(n7386), .ZN(n8117) );
  OR2_X1 U8564 ( .A1(n9531), .A2(n7386), .ZN(n6959) );
  NAND2_X1 U8565 ( .A1(n6925), .A2(n6963), .ZN(n8242) );
  NAND2_X2 U8566 ( .A1(n8237), .A2(n8242), .ZN(n8118) );
  NAND2_X1 U8567 ( .A1(n6960), .A2(n8118), .ZN(n7081) );
  OAI21_X1 U8568 ( .B1(n6960), .B2(n8118), .A(n7081), .ZN(n6978) );
  NOR2_X1 U8569 ( .A1(n7386), .A2(n7369), .ZN(n7381) );
  AND2_X1 U8570 ( .A1(n7381), .A2(n6963), .ZN(n7561) );
  INV_X1 U8571 ( .A(n7561), .ZN(n6961) );
  OAI21_X1 U8572 ( .B1(n6963), .B2(n7381), .A(n6961), .ZN(n7550) );
  OAI22_X1 U8573 ( .A1(n7550), .A2(n10228), .B1(n6963), .B2(n10226), .ZN(n6977) );
  INV_X1 U8574 ( .A(n6978), .ZN(n7557) );
  NAND2_X1 U8575 ( .A1(n6481), .A2(n8229), .ZN(n6965) );
  MUX2_X1 U8576 ( .A(n6965), .B(n6964), .S(n5914), .Z(n10175) );
  OR2_X1 U8577 ( .A1(n9531), .A2(n10196), .ZN(n6966) );
  NAND2_X1 U8578 ( .A1(n8238), .A2(n6967), .ZN(n7085) );
  OAI21_X1 U8579 ( .B1(n6967), .B2(n8238), .A(n7085), .ZN(n6975) );
  OR2_X1 U8580 ( .A1(n6481), .A2(n8229), .ZN(n6970) );
  NAND2_X1 U8581 ( .A1(n6483), .A2(n6968), .ZN(n6969) );
  OAI22_X1 U8582 ( .A1(n10170), .A2(n6973), .B1(n7084), .B2(n10167), .ZN(n6974) );
  AOI21_X1 U8583 ( .B1(n6975), .B2(n10172), .A(n6974), .ZN(n6976) );
  OAI21_X1 U8584 ( .B1(n7557), .B2(n10175), .A(n6976), .ZN(n7554) );
  AOI211_X1 U8585 ( .C1(n10233), .C2(n6978), .A(n6977), .B(n7554), .ZN(n7039)
         );
  NAND2_X1 U8586 ( .A1(n10243), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6979) );
  OAI21_X1 U8587 ( .B1(n7039), .B2(n10243), .A(n6979), .ZN(P1_U3525) );
  INV_X1 U8588 ( .A(n7351), .ZN(n7423) );
  OAI222_X1 U8589 ( .A1(P2_U3152), .A2(n7423), .B1(n9376), .B2(n6981), .C1(
        n6980), .C2(n9382), .ZN(P2_U3344) );
  XNOR2_X1 U8590 ( .A(n6983), .B(n6982), .ZN(n6990) );
  INV_X1 U8591 ( .A(n6984), .ZN(n7410) );
  NAND2_X1 U8592 ( .A1(n9512), .A2(n7197), .ZN(n6987) );
  INV_X1 U8593 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6985) );
  NOR2_X1 U8594 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6985), .ZN(n10035) );
  AOI21_X1 U8595 ( .B1(n9507), .B2(n9528), .A(n10035), .ZN(n6986) );
  OAI211_X1 U8596 ( .C1(n7084), .C2(n9505), .A(n6987), .B(n6986), .ZN(n6988)
         );
  AOI21_X1 U8597 ( .B1(n7410), .B2(n9466), .A(n6988), .ZN(n6989) );
  OAI21_X1 U8598 ( .B1(n6990), .B2(n9514), .A(n6989), .ZN(P1_U3228) );
  NAND2_X1 U8599 ( .A1(n10329), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6994) );
  MUX2_X1 U8600 ( .A(P2_REG2_REG_10__SCAN_IN), .B(n6991), .S(n10329), .Z(
        n10333) );
  INV_X1 U8601 ( .A(n6992), .ZN(n6999) );
  OAI21_X1 U8602 ( .B1(n6999), .B2(n7461), .A(n6993), .ZN(n10334) );
  NAND2_X1 U8603 ( .A1(n10333), .A2(n10334), .ZN(n10331) );
  AOI22_X1 U8604 ( .A1(n7061), .A2(n5294), .B1(P2_REG2_REG_11__SCAN_IN), .B2(
        n7068), .ZN(n6995) );
  AOI21_X1 U8605 ( .B1(n6996), .B2(n6995), .A(n7062), .ZN(n7010) );
  NAND2_X1 U8606 ( .A1(n10329), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7000) );
  INV_X1 U8607 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6997) );
  MUX2_X1 U8608 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6997), .S(n10329), .Z(
        n10337) );
  OAI21_X1 U8609 ( .B1(n6999), .B2(n6808), .A(n6998), .ZN(n10338) );
  NAND2_X1 U8610 ( .A1(n10337), .A2(n10338), .ZN(n10335) );
  NAND2_X1 U8611 ( .A1(n7000), .A2(n10335), .ZN(n7003) );
  MUX2_X1 U8612 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n7001), .S(n7061), .Z(n7002)
         );
  NAND2_X1 U8613 ( .A1(n7002), .A2(n7003), .ZN(n7067) );
  OAI211_X1 U8614 ( .C1(n7003), .C2(n7002), .A(n10336), .B(n7067), .ZN(n7007)
         );
  INV_X1 U8615 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7004) );
  NOR2_X1 U8616 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7004), .ZN(n7005) );
  AOI21_X1 U8617 ( .B1(n10328), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7005), .ZN(
        n7006) );
  NAND2_X1 U8618 ( .A1(n7007), .A2(n7006), .ZN(n7008) );
  AOI21_X1 U8619 ( .B1(n7061), .B2(n10330), .A(n7008), .ZN(n7009) );
  OAI21_X1 U8620 ( .B1(n7010), .B2(n10295), .A(n7009), .ZN(P2_U3256) );
  NOR2_X1 U8621 ( .A1(n7210), .A2(n7209), .ZN(n7012) );
  XNOR2_X1 U8622 ( .A(n7215), .B(n7014), .ZN(n9191) );
  NAND2_X1 U8623 ( .A1(n9191), .A2(n7237), .ZN(n10349) );
  INV_X1 U8624 ( .A(n7017), .ZN(n7020) );
  INV_X1 U8625 ( .A(n7158), .ZN(n7018) );
  AOI21_X1 U8626 ( .B1(n7020), .B2(n7019), .A(n7018), .ZN(n7281) );
  INV_X1 U8627 ( .A(n8431), .ZN(n10403) );
  INV_X1 U8628 ( .A(n7262), .ZN(n7022) );
  AOI211_X1 U8629 ( .C1(n8431), .C2(n6546), .A(n10455), .B(n7022), .ZN(n7278)
         );
  NAND2_X2 U8630 ( .A1(n7024), .A2(n7023), .ZN(n10371) );
  INV_X1 U8631 ( .A(n7025), .ZN(n7026) );
  NAND2_X1 U8632 ( .A1(n7017), .A2(n7026), .ZN(n7027) );
  OAI211_X1 U8633 ( .C1(n7029), .C2(n7028), .A(n10371), .B(n7027), .ZN(n7031)
         );
  AOI22_X1 U8634 ( .A1(n8629), .A2(n10366), .B1(n10368), .B2(n8626), .ZN(n7030) );
  NAND2_X1 U8635 ( .A1(n7031), .A2(n7030), .ZN(n7282) );
  AOI211_X1 U8636 ( .C1(n10444), .C2(n6546), .A(n7278), .B(n7282), .ZN(n7032)
         );
  OAI21_X1 U8637 ( .B1(n9926), .B2(n7281), .A(n7032), .ZN(n7037) );
  NAND2_X1 U8638 ( .A1(n7037), .A2(n10473), .ZN(n7033) );
  OAI21_X1 U8639 ( .B1(n10473), .B2(n8857), .A(n7033), .ZN(P2_U3521) );
  NOR2_X1 U8640 ( .A1(n7034), .A2(n7210), .ZN(n7035) );
  NAND2_X1 U8641 ( .A1(n7037), .A2(n10462), .ZN(n7038) );
  OAI21_X1 U8642 ( .B1(n10462), .B2(n5135), .A(n7038), .ZN(P2_U3454) );
  INV_X1 U8643 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n7041) );
  OR2_X1 U8644 ( .A1(n7039), .A2(n10234), .ZN(n7040) );
  OAI21_X1 U8645 ( .B1(n10236), .B2(n7041), .A(n7040), .ZN(P1_U3460) );
  INV_X1 U8646 ( .A(n7042), .ZN(n7049) );
  AOI22_X1 U8647 ( .A1(n10120), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n9882), .ZN(n7043) );
  OAI21_X1 U8648 ( .B1(n7049), .B2(n9886), .A(n7043), .ZN(P1_U3337) );
  INV_X1 U8649 ( .A(n7044), .ZN(n7047) );
  INV_X1 U8650 ( .A(n10109), .ZN(n9544) );
  OAI222_X1 U8651 ( .A1(n9891), .A2(n7045), .B1(n9886), .B2(n7047), .C1(
        P1_U3084), .C2(n9544), .ZN(P1_U3338) );
  INV_X1 U8652 ( .A(n7625), .ZN(n7424) );
  OAI222_X1 U8653 ( .A1(n7424), .A2(P2_U3152), .B1(n9376), .B2(n7047), .C1(
        n7046), .C2(n9382), .ZN(P2_U3343) );
  INV_X1 U8654 ( .A(n7667), .ZN(n7623) );
  OAI222_X1 U8655 ( .A1(P2_U3152), .A2(n7623), .B1(n9376), .B2(n7049), .C1(
        n7048), .C2(n9382), .ZN(P2_U3342) );
  INV_X1 U8656 ( .A(n7051), .ZN(n7052) );
  AOI21_X1 U8657 ( .B1(n7053), .B2(n7050), .A(n7052), .ZN(n7060) );
  INV_X1 U8658 ( .A(n7054), .ZN(n7402) );
  INV_X1 U8659 ( .A(n9529), .ZN(n7567) );
  NAND2_X1 U8660 ( .A1(n9512), .A2(n7398), .ZN(n7057) );
  NAND2_X1 U8661 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10049) );
  INV_X1 U8662 ( .A(n10049), .ZN(n7055) );
  AOI21_X1 U8663 ( .B1(n9507), .B2(n9526), .A(n7055), .ZN(n7056) );
  OAI211_X1 U8664 ( .C1(n7567), .C2(n9505), .A(n7057), .B(n7056), .ZN(n7058)
         );
  AOI21_X1 U8665 ( .B1(n7402), .B2(n9466), .A(n7058), .ZN(n7059) );
  OAI21_X1 U8666 ( .B1(n7060), .B2(n9514), .A(n7059), .ZN(P1_U3225) );
  NOR2_X1 U8667 ( .A1(n7061), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n7063) );
  INV_X1 U8668 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7745) );
  MUX2_X1 U8669 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7745), .S(n7075), .Z(n7064)
         );
  NAND2_X1 U8670 ( .A1(n7075), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7144) );
  OAI211_X1 U8671 ( .C1(n7065), .C2(n7064), .A(n7143), .B(n10332), .ZN(n7077)
         );
  INV_X1 U8672 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n7066) );
  NAND2_X1 U8673 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n10258) );
  OAI21_X1 U8674 ( .B1(n10304), .B2(n7066), .A(n10258), .ZN(n7074) );
  OAI21_X1 U8675 ( .B1(n7001), .B2(n7068), .A(n7067), .ZN(n7071) );
  MUX2_X1 U8676 ( .A(n7069), .B(P2_REG1_REG_12__SCAN_IN), .S(n7075), .Z(n7070)
         );
  NOR2_X1 U8677 ( .A1(n7070), .A2(n7071), .ZN(n7147) );
  AOI21_X1 U8678 ( .B1(n7071), .B2(n7070), .A(n7147), .ZN(n7072) );
  NOR2_X1 U8679 ( .A1(n10294), .A2(n7072), .ZN(n7073) );
  AOI211_X1 U8680 ( .C1(n10330), .C2(n7075), .A(n7074), .B(n7073), .ZN(n7076)
         );
  NAND2_X1 U8681 ( .A1(n7077), .A2(n7076), .ZN(P2_U3257) );
  INV_X1 U8682 ( .A(n7078), .ZN(n7099) );
  AOI22_X1 U8683 ( .A1(n10133), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n9882), .ZN(n7079) );
  OAI21_X1 U8684 ( .B1(n7099), .B2(n9886), .A(n7079), .ZN(P1_U3336) );
  OR2_X1 U8685 ( .A1(n6925), .A2(n7553), .ZN(n7080) );
  NAND2_X1 U8686 ( .A1(n7081), .A2(n7080), .ZN(n7559) );
  NAND2_X1 U8687 ( .A1(n9530), .A2(n10201), .ZN(n8246) );
  AND2_X1 U8688 ( .A1(n8243), .A2(n8246), .ZN(n7566) );
  INV_X1 U8689 ( .A(n7566), .ZN(n8120) );
  NAND2_X1 U8690 ( .A1(n7559), .A2(n8120), .ZN(n7558) );
  NAND2_X1 U8691 ( .A1(n7084), .A2(n10201), .ZN(n7082) );
  NAND2_X1 U8692 ( .A1(n7558), .A2(n7082), .ZN(n7083) );
  INV_X1 U8693 ( .A(n7197), .ZN(n7413) );
  OR2_X1 U8694 ( .A1(n7413), .A2(n9529), .ZN(n8249) );
  NAND2_X1 U8695 ( .A1(n9529), .A2(n7413), .ZN(n8171) );
  AND2_X1 U8696 ( .A1(n8249), .A2(n8171), .ZN(n8123) );
  INV_X1 U8697 ( .A(n8123), .ZN(n7086) );
  NAND2_X1 U8698 ( .A1(n7083), .A2(n7086), .ZN(n7199) );
  OAI21_X1 U8699 ( .B1(n7083), .B2(n7086), .A(n7199), .ZN(n7415) );
  INV_X1 U8700 ( .A(n7415), .ZN(n7093) );
  INV_X1 U8701 ( .A(n10175), .ZN(n9952) );
  INV_X1 U8702 ( .A(n9528), .ZN(n7138) );
  OAI22_X1 U8703 ( .A1(n10170), .A2(n7084), .B1(n7138), .B2(n10167), .ZN(n7090) );
  NAND2_X1 U8704 ( .A1(n8166), .A2(n7566), .ZN(n7565) );
  NAND2_X1 U8705 ( .A1(n7565), .A2(n8243), .ZN(n7087) );
  XNOR2_X1 U8706 ( .A(n7087), .B(n7086), .ZN(n7088) );
  NOR2_X1 U8707 ( .A1(n7088), .A2(n9949), .ZN(n7089) );
  AOI211_X1 U8708 ( .C1(n9952), .C2(n7415), .A(n7090), .B(n7089), .ZN(n7417)
         );
  NAND2_X1 U8709 ( .A1(n7561), .A2(n10201), .ZN(n7560) );
  OR2_X1 U8710 ( .A1(n7560), .A2(n7197), .ZN(n7399) );
  NAND2_X1 U8711 ( .A1(n7560), .A2(n7197), .ZN(n7091) );
  AND2_X1 U8712 ( .A1(n7399), .A2(n7091), .ZN(n7409) );
  AOI22_X1 U8713 ( .A1(n7409), .A2(n9984), .B1(n7197), .B2(n9849), .ZN(n7092)
         );
  OAI211_X1 U8714 ( .C1(n7093), .C2(n9862), .A(n7417), .B(n7092), .ZN(n7095)
         );
  NAND2_X1 U8715 ( .A1(n7095), .A2(n10245), .ZN(n7094) );
  OAI21_X1 U8716 ( .B1(n10245), .B2(n6695), .A(n7094), .ZN(P1_U3527) );
  INV_X1 U8717 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n7097) );
  NAND2_X1 U8718 ( .A1(n7095), .A2(n10236), .ZN(n7096) );
  OAI21_X1 U8719 ( .B1(n10236), .B2(n7097), .A(n7096), .ZN(P1_U3466) );
  INV_X1 U8720 ( .A(n7673), .ZN(n8646) );
  OAI222_X1 U8721 ( .A1(P2_U3152), .A2(n8646), .B1(n9376), .B2(n7099), .C1(
        n7098), .C2(n9382), .ZN(P2_U3341) );
  INV_X1 U8722 ( .A(n10084), .ZN(n7103) );
  NOR2_X1 U8723 ( .A1(n7113), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7100) );
  NOR2_X1 U8724 ( .A1(n7101), .A2(n7100), .ZN(n10087) );
  MUX2_X1 U8725 ( .A(n7102), .B(P1_REG1_REG_12__SCAN_IN), .S(n10084), .Z(
        n10086) );
  NOR2_X1 U8726 ( .A1(n10087), .A2(n10086), .ZN(n10085) );
  AOI21_X1 U8727 ( .B1(n7103), .B2(n7102), .A(n10085), .ZN(n10099) );
  MUX2_X1 U8728 ( .A(n7104), .B(P1_REG1_REG_13__SCAN_IN), .S(n10097), .Z(
        n10100) );
  NOR2_X1 U8729 ( .A1(n10099), .A2(n10100), .ZN(n10098) );
  AOI21_X1 U8730 ( .B1(n7104), .B2(n7105), .A(n10098), .ZN(n7108) );
  AOI22_X1 U8731 ( .A1(n7106), .A2(n6200), .B1(P1_REG1_REG_14__SCAN_IN), .B2(
        n9541), .ZN(n7107) );
  NOR2_X1 U8732 ( .A1(n7108), .A2(n7107), .ZN(n9540) );
  AOI21_X1 U8733 ( .B1(n7108), .B2(n7107), .A(n9540), .ZN(n7119) );
  NOR2_X1 U8734 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7109), .ZN(n7913) );
  NOR2_X1 U8735 ( .A1(n10074), .A2(n9541), .ZN(n7110) );
  AOI211_X1 U8736 ( .C1(n10052), .C2(P1_ADDR_REG_14__SCAN_IN), .A(n7913), .B(
        n7110), .ZN(n7118) );
  NAND2_X1 U8737 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(n10084), .ZN(n7111) );
  OAI21_X1 U8738 ( .B1(n10084), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7111), .ZN(
        n10080) );
  NAND2_X1 U8739 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n10097), .ZN(n7114) );
  OAI21_X1 U8740 ( .B1(n10097), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7114), .ZN(
        n10093) );
  NOR2_X1 U8741 ( .A1(n10094), .A2(n10093), .ZN(n10092) );
  OAI21_X1 U8742 ( .B1(n7115), .B2(n6203), .A(n9533), .ZN(n7116) );
  NAND2_X1 U8743 ( .A1(n7116), .A2(n10058), .ZN(n7117) );
  OAI211_X1 U8744 ( .C1(n7119), .C2(n10154), .A(n7118), .B(n7117), .ZN(
        P1_U3255) );
  NAND2_X1 U8745 ( .A1(n10287), .A2(n8314), .ZN(n8603) );
  NOR3_X1 U8746 ( .A1(n8603), .A2(n7120), .A3(n7314), .ZN(n7121) );
  AOI21_X1 U8747 ( .B1(n4513), .B2(n10287), .A(n7121), .ZN(n7131) );
  INV_X1 U8748 ( .A(n10292), .ZN(n8597) );
  INV_X1 U8749 ( .A(n7323), .ZN(n7128) );
  NAND2_X1 U8750 ( .A1(n10257), .A2(n8625), .ZN(n7124) );
  AOI21_X1 U8751 ( .B1(n10286), .B2(n4785), .A(n7122), .ZN(n7123) );
  OAI211_X1 U8752 ( .C1(n7313), .C2(n10260), .A(n7124), .B(n7123), .ZN(n7127)
         );
  NOR2_X1 U8753 ( .A1(n7125), .A2(n10246), .ZN(n7126) );
  AOI211_X1 U8754 ( .C1(n8597), .C2(n7128), .A(n7127), .B(n7126), .ZN(n7129)
         );
  OAI21_X1 U8755 ( .B1(n7131), .B2(n7130), .A(n7129), .ZN(P2_U3232) );
  INV_X1 U8756 ( .A(n7466), .ZN(n7363) );
  OAI21_X1 U8757 ( .B1(n7134), .B2(n7132), .A(n7133), .ZN(n7135) );
  NAND2_X1 U8758 ( .A1(n7135), .A2(n9483), .ZN(n7142) );
  INV_X1 U8759 ( .A(n7362), .ZN(n7140) );
  AOI21_X1 U8760 ( .B1(n9507), .B2(n9525), .A(n7136), .ZN(n7137) );
  OAI21_X1 U8761 ( .B1(n9505), .B2(n7138), .A(n7137), .ZN(n7139) );
  AOI21_X1 U8762 ( .B1(n9466), .B2(n7140), .A(n7139), .ZN(n7141) );
  OAI211_X1 U8763 ( .C1(n7363), .C2(n9492), .A(n7142), .B(n7141), .ZN(P1_U3237) );
  NAND2_X1 U8764 ( .A1(n7144), .A2(n7143), .ZN(n7146) );
  AOI22_X1 U8765 ( .A1(n7338), .A2(n7883), .B1(P2_REG2_REG_13__SCAN_IN), .B2(
        n7345), .ZN(n7145) );
  NOR2_X1 U8766 ( .A1(n7146), .A2(n7145), .ZN(n7339) );
  AOI21_X1 U8767 ( .B1(n7146), .B2(n7145), .A(n7339), .ZN(n7156) );
  AOI21_X1 U8768 ( .B1(n7069), .B2(n7148), .A(n7147), .ZN(n7150) );
  AOI22_X1 U8769 ( .A1(n7338), .A2(n5335), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7345), .ZN(n7149) );
  NOR2_X1 U8770 ( .A1(n7150), .A2(n7149), .ZN(n7344) );
  AOI21_X1 U8771 ( .B1(n7150), .B2(n7149), .A(n7344), .ZN(n7153) );
  NOR2_X1 U8772 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7827), .ZN(n7151) );
  AOI21_X1 U8773 ( .B1(n10328), .B2(P2_ADDR_REG_13__SCAN_IN), .A(n7151), .ZN(
        n7152) );
  OAI21_X1 U8774 ( .B1(n10294), .B2(n7153), .A(n7152), .ZN(n7154) );
  AOI21_X1 U8775 ( .B1(n7338), .B2(n10330), .A(n7154), .ZN(n7155) );
  OAI21_X1 U8776 ( .B1(n7156), .B2(n10295), .A(n7155), .ZN(P2_U3258) );
  NAND2_X1 U8777 ( .A1(n7158), .A2(n7157), .ZN(n7261) );
  NAND2_X1 U8778 ( .A1(n10251), .A2(n10408), .ZN(n7159) );
  NAND2_X1 U8779 ( .A1(n7260), .A2(n7159), .ZN(n7161) );
  INV_X1 U8780 ( .A(n7164), .ZN(n7160) );
  NAND2_X1 U8781 ( .A1(n7161), .A2(n7160), .ZN(n7231) );
  OAI21_X1 U8782 ( .B1(n7161), .B2(n7160), .A(n7231), .ZN(n7223) );
  INV_X1 U8783 ( .A(n7223), .ZN(n7171) );
  OAI21_X1 U8784 ( .B1(n7164), .B2(n7163), .A(n7162), .ZN(n7167) );
  INV_X1 U8785 ( .A(n10368), .ZN(n9240) );
  OAI22_X1 U8786 ( .A1(n10251), .A2(n9242), .B1(n4786), .B2(n9240), .ZN(n7166)
         );
  NOR2_X1 U8787 ( .A1(n7171), .A2(n10349), .ZN(n7165) );
  AOI211_X1 U8788 ( .C1(n10371), .C2(n7167), .A(n7166), .B(n7165), .ZN(n7225)
         );
  INV_X1 U8789 ( .A(n7265), .ZN(n7168) );
  AOI21_X1 U8790 ( .B1(n10444), .B2(n7169), .A(n7220), .ZN(n7170) );
  OAI211_X1 U8791 ( .C1(n7171), .C2(n10428), .A(n7225), .B(n7170), .ZN(n7173)
         );
  NAND2_X1 U8792 ( .A1(n7173), .A2(n10473), .ZN(n7172) );
  OAI21_X1 U8793 ( .B1(n10473), .B2(n6770), .A(n7172), .ZN(P2_U3523) );
  INV_X1 U8794 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n7175) );
  NAND2_X1 U8795 ( .A1(n7173), .A2(n10462), .ZN(n7174) );
  OAI21_X1 U8796 ( .B1(n10462), .B2(n7175), .A(n7174), .ZN(P2_U3460) );
  NAND2_X1 U8797 ( .A1(n5066), .A2(n7177), .ZN(n7178) );
  XNOR2_X1 U8798 ( .A(n7176), .B(n7178), .ZN(n7185) );
  INV_X1 U8799 ( .A(n7179), .ZN(n7181) );
  INV_X1 U8800 ( .A(n9526), .ZN(n7526) );
  NOR2_X1 U8801 ( .A1(n9505), .A2(n7526), .ZN(n7180) );
  AOI211_X1 U8802 ( .C1(n9507), .C2(n9524), .A(n7181), .B(n7180), .ZN(n7182)
         );
  OAI21_X1 U8803 ( .B1(n9510), .B2(n7529), .A(n7182), .ZN(n7183) );
  AOI21_X1 U8804 ( .B1(n9512), .B2(n7532), .A(n7183), .ZN(n7184) );
  OAI21_X1 U8805 ( .B1(n7185), .B2(n9514), .A(n7184), .ZN(P1_U3211) );
  OAI21_X1 U8806 ( .B1(n7188), .B2(n7187), .A(n7186), .ZN(n7189) );
  NAND2_X1 U8807 ( .A1(n7189), .A2(n10287), .ZN(n7196) );
  NOR2_X1 U8808 ( .A1(n10292), .A2(n7190), .ZN(n7194) );
  NAND2_X1 U8809 ( .A1(n10257), .A2(n10367), .ZN(n7192) );
  OAI211_X1 U8810 ( .C1(n7444), .C2(n10260), .A(n7192), .B(n7191), .ZN(n7193)
         );
  AOI211_X1 U8811 ( .C1(n10286), .C2(n7302), .A(n7194), .B(n7193), .ZN(n7195)
         );
  NAND2_X1 U8812 ( .A1(n7196), .A2(n7195), .ZN(P2_U3241) );
  OR2_X1 U8813 ( .A1(n9529), .A2(n7197), .ZN(n7198) );
  INV_X1 U8814 ( .A(n7398), .ZN(n10207) );
  AND2_X1 U8815 ( .A1(n9528), .A2(n10207), .ZN(n7485) );
  INV_X1 U8816 ( .A(n7485), .ZN(n8170) );
  OR2_X1 U8817 ( .A1(n9528), .A2(n10207), .ZN(n7483) );
  AND2_X1 U8818 ( .A1(n8170), .A2(n7483), .ZN(n7394) );
  INV_X1 U8819 ( .A(n7394), .ZN(n7200) );
  NAND2_X1 U8820 ( .A1(n9528), .A2(n7398), .ZN(n7201) );
  OR2_X1 U8821 ( .A1(n7526), .A2(n7466), .ZN(n8122) );
  NAND2_X1 U8822 ( .A1(n7526), .A2(n7466), .ZN(n8031) );
  NAND2_X1 U8823 ( .A1(n8122), .A2(n8031), .ZN(n8036) );
  OAI21_X1 U8824 ( .B1(n7202), .B2(n8036), .A(n7468), .ZN(n7206) );
  INV_X1 U8825 ( .A(n7206), .ZN(n7368) );
  AND2_X1 U8826 ( .A1(n8243), .A2(n8249), .ZN(n8169) );
  XNOR2_X1 U8827 ( .A(n8037), .B(n8036), .ZN(n7204) );
  AOI22_X1 U8828 ( .A1(n9947), .A2(n9525), .B1(n9945), .B2(n9528), .ZN(n7203)
         );
  OAI21_X1 U8829 ( .B1(n7204), .B2(n9949), .A(n7203), .ZN(n7205) );
  AOI21_X1 U8830 ( .B1(n7206), .B2(n9952), .A(n7205), .ZN(n7360) );
  OR2_X1 U8831 ( .A1(n7399), .A2(n7398), .ZN(n7400) );
  AOI211_X1 U8832 ( .C1(n7466), .C2(n7400), .A(n10228), .B(n7528), .ZN(n7365)
         );
  AOI21_X1 U8833 ( .B1(n7466), .B2(n9849), .A(n7365), .ZN(n7207) );
  OAI211_X1 U8834 ( .C1(n7368), .C2(n9862), .A(n7360), .B(n7207), .ZN(n7226)
         );
  NAND2_X1 U8835 ( .A1(n7226), .A2(n10245), .ZN(n7208) );
  OAI21_X1 U8836 ( .B1(n10245), .B2(n6032), .A(n7208), .ZN(P1_U3529) );
  AND2_X1 U8837 ( .A1(n7210), .A2(n7209), .ZN(n7211) );
  NAND2_X1 U8838 ( .A1(n7212), .A2(n7211), .ZN(n7218) );
  INV_X1 U8839 ( .A(n7213), .ZN(n7214) );
  NOR2_X1 U8840 ( .A1(n7215), .A2(n7237), .ZN(n7216) );
  NAND2_X1 U8841 ( .A1(n9259), .A2(n7216), .ZN(n10360) );
  INV_X1 U8842 ( .A(n10360), .ZN(n9263) );
  NOR2_X1 U8843 ( .A1(n8355), .A2(n10404), .ZN(n7217) );
  OR2_X1 U8844 ( .A1(n7218), .A2(n9194), .ZN(n10359) );
  INV_X1 U8845 ( .A(n10359), .ZN(n9179) );
  OAI22_X1 U8846 ( .A1(n9259), .A2(n6789), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9256), .ZN(n7219) );
  AOI21_X1 U8847 ( .B1(n7220), .B2(n9179), .A(n7219), .ZN(n7221) );
  OAI21_X1 U8848 ( .B1(n10250), .B2(n9254), .A(n7221), .ZN(n7222) );
  AOI21_X1 U8849 ( .B1(n9263), .B2(n7223), .A(n7222), .ZN(n7224) );
  OAI21_X1 U8850 ( .B1(n7225), .B2(n10372), .A(n7224), .ZN(P2_U3293) );
  INV_X1 U8851 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7228) );
  NAND2_X1 U8852 ( .A1(n7226), .A2(n10236), .ZN(n7227) );
  OAI21_X1 U8853 ( .B1(n10236), .B2(n7228), .A(n7227), .ZN(P1_U3472) );
  INV_X1 U8854 ( .A(n10349), .ZN(n9250) );
  NAND2_X1 U8855 ( .A1(n9259), .A2(n9250), .ZN(n7229) );
  NAND2_X1 U8856 ( .A1(n7314), .A2(n10250), .ZN(n7230) );
  NAND2_X1 U8857 ( .A1(n7231), .A2(n7230), .ZN(n7320) );
  NAND2_X1 U8858 ( .A1(n7320), .A2(n7319), .ZN(n7318) );
  NAND2_X1 U8859 ( .A1(n4786), .A2(n10414), .ZN(n7232) );
  XOR2_X1 U8860 ( .A(n7294), .B(n7297), .Z(n7253) );
  XOR2_X1 U8861 ( .A(n7233), .B(n7294), .Z(n7234) );
  INV_X1 U8862 ( .A(n10371), .ZN(n9246) );
  AOI22_X1 U8863 ( .A1(n8623), .A2(n10368), .B1(n10366), .B2(n8624), .ZN(
        n10277) );
  OAI21_X1 U8864 ( .B1(n7234), .B2(n9246), .A(n10277), .ZN(n7250) );
  INV_X1 U8865 ( .A(n7250), .ZN(n7236) );
  MUX2_X1 U8866 ( .A(n7236), .B(n7235), .S(n10372), .Z(n7241) );
  AOI211_X1 U8867 ( .C1(n10285), .C2(n7321), .A(n10455), .B(n4571), .ZN(n7251)
         );
  AND2_X1 U8868 ( .A1(n9259), .A2(n7237), .ZN(n9230) );
  OAI22_X1 U8869 ( .A1(n9254), .A2(n7238), .B1(n9256), .B2(n10291), .ZN(n7239)
         );
  AOI21_X1 U8870 ( .B1(n7251), .B2(n9230), .A(n7239), .ZN(n7240) );
  OAI211_X1 U8871 ( .C1(n9233), .C2(n7253), .A(n7241), .B(n7240), .ZN(P2_U3291) );
  XNOR2_X1 U8872 ( .A(n7243), .B(n7242), .ZN(n7249) );
  NOR2_X1 U8873 ( .A1(n10292), .A2(n7304), .ZN(n7247) );
  NAND2_X1 U8874 ( .A1(n10257), .A2(n8623), .ZN(n7245) );
  OR2_X1 U8875 ( .A1(n10260), .A2(n7453), .ZN(n7244) );
  OAI211_X1 U8876 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n5210), .A(n7245), .B(n7244), .ZN(n7246) );
  AOI211_X1 U8877 ( .C1(n10286), .C2(n7458), .A(n7247), .B(n7246), .ZN(n7248)
         );
  OAI21_X1 U8878 ( .B1(n7249), .B2(n10246), .A(n7248), .ZN(P2_U3215) );
  AOI211_X1 U8879 ( .C1(n10444), .C2(n10285), .A(n7251), .B(n7250), .ZN(n7252)
         );
  OAI21_X1 U8880 ( .B1(n9926), .B2(n7253), .A(n7252), .ZN(n7255) );
  NAND2_X1 U8881 ( .A1(n7255), .A2(n10473), .ZN(n7254) );
  OAI21_X1 U8882 ( .B1(n10473), .B2(n6769), .A(n7254), .ZN(P2_U3525) );
  NAND2_X1 U8883 ( .A1(n7255), .A2(n10462), .ZN(n7256) );
  OAI21_X1 U8884 ( .B1(n10462), .B2(n5175), .A(n7256), .ZN(P2_U3466) );
  INV_X1 U8885 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n8880) );
  INV_X1 U8886 ( .A(n7257), .ZN(n7258) );
  INV_X1 U8887 ( .A(n10149), .ZN(n9551) );
  OAI222_X1 U8888 ( .A1(n9891), .A2(n8880), .B1(n9886), .B2(n7258), .C1(
        P1_U3084), .C2(n9551), .ZN(P1_U3335) );
  INV_X1 U8889 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7259) );
  INV_X1 U8890 ( .A(n8657), .ZN(n8656) );
  OAI222_X1 U8891 ( .A1(n9382), .A2(n7259), .B1(n9376), .B2(n7258), .C1(n8656), 
        .C2(P2_U3152), .ZN(P2_U3340) );
  OAI21_X1 U8892 ( .B1(n7261), .B2(n7269), .A(n7260), .ZN(n10411) );
  INV_X1 U8893 ( .A(n10411), .ZN(n7277) );
  NOR2_X1 U8894 ( .A1(n9259), .A2(n6791), .ZN(n7268) );
  NAND2_X1 U8895 ( .A1(n7262), .A2(n8576), .ZN(n7263) );
  NAND2_X1 U8896 ( .A1(n7263), .A2(n10447), .ZN(n7264) );
  OR2_X1 U8897 ( .A1(n7265), .A2(n7264), .ZN(n10407) );
  INV_X1 U8898 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7266) );
  OAI22_X1 U8899 ( .A1(n10359), .A2(n10407), .B1(n7266), .B2(n9256), .ZN(n7267) );
  AOI211_X1 U8900 ( .C1(n10355), .C2(n8576), .A(n7268), .B(n7267), .ZN(n7276)
         );
  XNOR2_X1 U8901 ( .A(n7270), .B(n7269), .ZN(n7271) );
  NAND2_X1 U8902 ( .A1(n7271), .A2(n10371), .ZN(n7274) );
  OAI22_X1 U8903 ( .A1(n8580), .A2(n9242), .B1(n7314), .B2(n9240), .ZN(n7272)
         );
  INV_X1 U8904 ( .A(n7272), .ZN(n7273) );
  NAND2_X1 U8905 ( .A1(n7274), .A2(n7273), .ZN(n10409) );
  NAND2_X1 U8906 ( .A1(n10409), .A2(n9259), .ZN(n7275) );
  OAI211_X1 U8907 ( .C1(n7277), .C2(n9233), .A(n7276), .B(n7275), .ZN(P2_U3294) );
  INV_X1 U8908 ( .A(n9256), .ZN(n10373) );
  AOI22_X1 U8909 ( .A1(n7278), .A2(n9179), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n10373), .ZN(n7280) );
  NAND2_X1 U8910 ( .A1(n10355), .A2(n6546), .ZN(n7279) );
  OAI211_X1 U8911 ( .C1(n7281), .C2(n9233), .A(n7280), .B(n7279), .ZN(n7284)
         );
  MUX2_X1 U8912 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n7282), .S(n9259), .Z(n7283)
         );
  OR2_X1 U8913 ( .A1(n7284), .A2(n7283), .ZN(P2_U3295) );
  INV_X1 U8914 ( .A(n7285), .ZN(n7288) );
  OAI222_X1 U8915 ( .A1(n9891), .A2(n7286), .B1(n9886), .B2(n7288), .C1(n8229), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OAI222_X1 U8916 ( .A1(P2_U3152), .A2(n7237), .B1(n9376), .B2(n7288), .C1(
        n7287), .C2(n9382), .ZN(P2_U3339) );
  NOR2_X2 U8917 ( .A1(n10359), .A2(n10455), .ZN(n9262) );
  OR2_X1 U8918 ( .A1(n9262), .A2(n10355), .ZN(n10380) );
  NOR2_X1 U8919 ( .A1(n8580), .A2(n9240), .ZN(n7289) );
  AOI21_X1 U8920 ( .B1(n10406), .B2(n10371), .A(n7289), .ZN(n10402) );
  AOI22_X1 U8921 ( .A1(n10372), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(n10373), .ZN(n7290) );
  OAI21_X1 U8922 ( .B1(n10402), .B2(n10372), .A(n7290), .ZN(n7291) );
  AOI21_X1 U8923 ( .B1(n8431), .B2(n10380), .A(n7291), .ZN(n7292) );
  OAI21_X1 U8924 ( .B1(n7293), .B2(n9233), .A(n7292), .ZN(P2_U3296) );
  NOR2_X1 U8925 ( .A1(n10367), .A2(n10285), .ZN(n7296) );
  OR2_X1 U8926 ( .A1(n7294), .A2(n7313), .ZN(n7295) );
  AND2_X1 U8927 ( .A1(n8623), .A2(n7302), .ZN(n7298) );
  XNOR2_X1 U8928 ( .A(n7442), .B(n7441), .ZN(n10426) );
  INV_X1 U8929 ( .A(n10426), .ZN(n7309) );
  XNOR2_X1 U8930 ( .A(n7299), .B(n7441), .ZN(n7300) );
  OAI222_X1 U8931 ( .A1(n9240), .A2(n7453), .B1(n9242), .B2(n7301), .C1(n7300), 
        .C2(n9246), .ZN(n10424) );
  NAND2_X1 U8932 ( .A1(n10424), .A2(n7864), .ZN(n7308) );
  XNOR2_X1 U8933 ( .A(n10377), .B(n7458), .ZN(n7303) );
  OAI22_X1 U8934 ( .A1(n7303), .A2(n10455), .B1(n7443), .B2(n10453), .ZN(
        n10425) );
  OAI22_X1 U8935 ( .A1(n9259), .A2(n7305), .B1(n7304), .B2(n9256), .ZN(n7306)
         );
  AOI21_X1 U8936 ( .B1(n10425), .B2(n10380), .A(n7306), .ZN(n7307) );
  OAI211_X1 U8937 ( .C1(n9233), .C2(n7309), .A(n7308), .B(n7307), .ZN(P2_U3289) );
  INV_X1 U8938 ( .A(n7319), .ZN(n7310) );
  XNOR2_X1 U8939 ( .A(n7311), .B(n7310), .ZN(n7312) );
  NAND2_X1 U8940 ( .A1(n7312), .A2(n10371), .ZN(n7317) );
  OAI22_X1 U8941 ( .A1(n7314), .A2(n9242), .B1(n7313), .B2(n9240), .ZN(n7315)
         );
  INV_X1 U8942 ( .A(n7315), .ZN(n7316) );
  NAND2_X1 U8943 ( .A1(n7317), .A2(n7316), .ZN(n10415) );
  INV_X1 U8944 ( .A(n10415), .ZN(n7328) );
  OAI21_X1 U8945 ( .B1(n7320), .B2(n7319), .A(n7318), .ZN(n10417) );
  INV_X1 U8946 ( .A(n9233), .ZN(n10381) );
  OAI211_X1 U8947 ( .C1(n7322), .C2(n10414), .A(n10447), .B(n7321), .ZN(n10413) );
  OAI22_X1 U8948 ( .A1(n6794), .A2(n9259), .B1(n7323), .B2(n9256), .ZN(n7324)
         );
  AOI21_X1 U8949 ( .B1(n10355), .B2(n4785), .A(n7324), .ZN(n7325) );
  OAI21_X1 U8950 ( .B1(n10413), .B2(n10359), .A(n7325), .ZN(n7326) );
  AOI21_X1 U8951 ( .B1(n10417), .B2(n10381), .A(n7326), .ZN(n7327) );
  OAI21_X1 U8952 ( .B1(n7328), .B2(n10372), .A(n7327), .ZN(P2_U3292) );
  XNOR2_X1 U8953 ( .A(n7330), .B(n7329), .ZN(n7337) );
  OR2_X1 U8954 ( .A1(n7444), .A2(n9242), .ZN(n7331) );
  OAI21_X1 U8955 ( .B1(n7501), .B2(n9240), .A(n7331), .ZN(n10351) );
  NAND2_X1 U8956 ( .A1(n10351), .A2(n10279), .ZN(n7334) );
  INV_X1 U8957 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7332) );
  NOR2_X1 U8958 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7332), .ZN(n8633) );
  INV_X1 U8959 ( .A(n8633), .ZN(n7333) );
  OAI211_X1 U8960 ( .C1(n10292), .C2(n10353), .A(n7334), .B(n7333), .ZN(n7335)
         );
  AOI21_X1 U8961 ( .B1(n10286), .B2(n10356), .A(n7335), .ZN(n7336) );
  OAI21_X1 U8962 ( .B1(n7337), .B2(n10246), .A(n7336), .ZN(P2_U3223) );
  NOR2_X1 U8963 ( .A1(n7338), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7340) );
  AOI22_X1 U8964 ( .A1(n7351), .A2(n7860), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n7423), .ZN(n7341) );
  AOI21_X1 U8965 ( .B1(n7342), .B2(n7341), .A(n7418), .ZN(n7353) );
  INV_X1 U8966 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n7343) );
  NAND2_X1 U8967 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3152), .ZN(n7946) );
  OAI21_X1 U8968 ( .B1(n10304), .B2(n7343), .A(n7946), .ZN(n7350) );
  AOI21_X1 U8969 ( .B1(n7345), .B2(n5335), .A(n7344), .ZN(n7347) );
  AOI22_X1 U8970 ( .A1(n7351), .A2(n5356), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7423), .ZN(n7346) );
  NOR2_X1 U8971 ( .A1(n7347), .A2(n7346), .ZN(n7422) );
  AOI21_X1 U8972 ( .B1(n7347), .B2(n7346), .A(n7422), .ZN(n7348) );
  NOR2_X1 U8973 ( .A1(n7348), .A2(n10294), .ZN(n7349) );
  AOI211_X1 U8974 ( .C1(n10330), .C2(n7351), .A(n7350), .B(n7349), .ZN(n7352)
         );
  OAI21_X1 U8975 ( .B1(n7353), .B2(n10295), .A(n7352), .ZN(P2_U3259) );
  NAND2_X1 U8976 ( .A1(n7355), .A2(n7354), .ZN(n7356) );
  NAND2_X1 U8977 ( .A1(n8236), .A2(n8270), .ZN(n7358) );
  NOR3_X1 U8978 ( .A1(n9953), .A2(n8229), .A3(n5914), .ZN(n10164) );
  INV_X1 U8979 ( .A(n10164), .ZN(n7735) );
  MUX2_X1 U8980 ( .A(n7360), .B(n7359), .S(n9953), .Z(n7367) );
  NAND2_X1 U8981 ( .A1(n10181), .A2(n8229), .ZN(n9586) );
  INV_X1 U8982 ( .A(n9586), .ZN(n9747) );
  OAI22_X1 U8983 ( .A1(n10177), .A2(n7363), .B1(n10178), .B2(n7362), .ZN(n7364) );
  AOI21_X1 U8984 ( .B1(n7365), .B2(n9747), .A(n7364), .ZN(n7366) );
  OAI211_X1 U8985 ( .C1(n7368), .C2(n7735), .A(n7367), .B(n7366), .ZN(P1_U3285) );
  NOR2_X2 U8986 ( .A1(n9586), .A2(n10228), .ZN(n10163) );
  OAI21_X1 U8987 ( .B1(n10163), .B2(n9957), .A(n7369), .ZN(n7372) );
  INV_X1 U8988 ( .A(n10178), .ZN(n9763) );
  AOI22_X1 U8989 ( .A1(n10181), .A2(n7370), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        n9763), .ZN(n7371) );
  OAI211_X1 U8990 ( .C1(n5938), .C2(n10181), .A(n7372), .B(n7371), .ZN(
        P1_U3291) );
  INV_X1 U8991 ( .A(n7373), .ZN(n7374) );
  AOI21_X1 U8992 ( .B1(n7375), .B2(n8117), .A(n7374), .ZN(n10194) );
  OAI22_X1 U8993 ( .A1(n10170), .A2(n7377), .B1(n7568), .B2(n10167), .ZN(n7378) );
  AOI21_X1 U8994 ( .B1(n7379), .B2(n10172), .A(n7378), .ZN(n7380) );
  OAI21_X1 U8995 ( .B1(n10194), .B2(n10175), .A(n7380), .ZN(n10197) );
  INV_X1 U8996 ( .A(n7381), .ZN(n7382) );
  OAI211_X1 U8997 ( .C1(n10196), .C2(n7383), .A(n9984), .B(n7382), .ZN(n10195)
         );
  OAI22_X1 U8998 ( .A1(n10195), .A2(n4695), .B1(n10178), .B2(n7384), .ZN(n7385) );
  OAI21_X1 U8999 ( .B1(n10197), .B2(n7385), .A(n10181), .ZN(n7388) );
  AOI22_X1 U9000 ( .A1(n9957), .A2(n7386), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n9953), .ZN(n7387) );
  OAI211_X1 U9001 ( .C1(n7735), .C2(n10194), .A(n7388), .B(n7387), .ZN(
        P1_U3290) );
  AND2_X1 U9002 ( .A1(n8272), .A2(n7389), .ZN(n7390) );
  INV_X1 U9003 ( .A(n9777), .ZN(n9730) );
  NAND2_X1 U9004 ( .A1(n7391), .A2(n7394), .ZN(n7392) );
  AND2_X1 U9005 ( .A1(n7393), .A2(n7392), .ZN(n10209) );
  OAI22_X1 U9006 ( .A1(n10177), .A2(n10207), .B1(n6002), .B2(n10181), .ZN(
        n7406) );
  XNOR2_X1 U9007 ( .A(n7484), .B(n7200), .ZN(n7397) );
  NAND2_X1 U9008 ( .A1(n9945), .A2(n9529), .ZN(n7395) );
  OAI21_X1 U9009 ( .B1(n7526), .B2(n10167), .A(n7395), .ZN(n7396) );
  AOI21_X1 U9010 ( .B1(n7397), .B2(n10172), .A(n7396), .ZN(n10210) );
  AOI21_X1 U9011 ( .B1(n7399), .B2(n7398), .A(n10228), .ZN(n7401) );
  NAND2_X1 U9012 ( .A1(n7401), .A2(n7400), .ZN(n10206) );
  INV_X1 U9013 ( .A(n10206), .ZN(n7403) );
  AOI22_X1 U9014 ( .A1(n7403), .A2(n8229), .B1(n9763), .B2(n7402), .ZN(n7404)
         );
  AOI21_X1 U9015 ( .B1(n10210), .B2(n7404), .A(n9953), .ZN(n7405) );
  AOI211_X1 U9016 ( .C1(n9730), .C2(n10209), .A(n7406), .B(n7405), .ZN(n7407)
         );
  INV_X1 U9017 ( .A(n7407), .ZN(P1_U3286) );
  INV_X1 U9018 ( .A(n7408), .ZN(n8354) );
  OAI222_X1 U9019 ( .A1(n9886), .A2(n8354), .B1(P1_U3084), .B2(n8266), .C1(
        n8898), .C2(n9891), .ZN(P1_U3333) );
  NAND2_X1 U9020 ( .A1(n10163), .A2(n7409), .ZN(n7412) );
  AOI22_X1 U9021 ( .A1(n9953), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7410), .B2(
        n9763), .ZN(n7411) );
  OAI211_X1 U9022 ( .C1(n7413), .C2(n10177), .A(n7412), .B(n7411), .ZN(n7414)
         );
  AOI21_X1 U9023 ( .B1(n7415), .B2(n10164), .A(n7414), .ZN(n7416) );
  OAI21_X1 U9024 ( .B1(n7417), .B2(n9953), .A(n7416), .ZN(P1_U3287) );
  NOR2_X1 U9025 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n7419), .ZN(n7626) );
  AOI21_X1 U9026 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n7419), .A(n7626), .ZN(
        n7428) );
  INV_X1 U9027 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n7420) );
  NAND2_X1 U9028 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7966) );
  OAI21_X1 U9029 ( .B1(n10304), .B2(n7420), .A(n7966), .ZN(n7421) );
  AOI21_X1 U9030 ( .B1(n10330), .B2(n7625), .A(n7421), .ZN(n7427) );
  AOI21_X1 U9031 ( .B1(n7423), .B2(n5356), .A(n7422), .ZN(n7617) );
  XNOR2_X1 U9032 ( .A(n7617), .B(n7424), .ZN(n7425) );
  NAND2_X1 U9033 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7425), .ZN(n7618) );
  OAI211_X1 U9034 ( .C1(n7425), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10336), .B(
        n7618), .ZN(n7426) );
  OAI211_X1 U9035 ( .C1(n7428), .C2(n10295), .A(n7427), .B(n7426), .ZN(
        P2_U3260) );
  INV_X1 U9036 ( .A(n7429), .ZN(n7431) );
  NAND2_X1 U9037 ( .A1(n7431), .A2(n7430), .ZN(n7433) );
  AOI22_X1 U9038 ( .A1(n7434), .A2(n7433), .B1(n7510), .B2(n7432), .ZN(n7440)
         );
  NOR2_X1 U9039 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7435), .ZN(n10053) );
  INV_X1 U9040 ( .A(n9523), .ZN(n7585) );
  NOR2_X1 U9041 ( .A1(n9486), .A2(n7585), .ZN(n7436) );
  AOI211_X1 U9042 ( .C1(n9495), .C2(n9525), .A(n10053), .B(n7436), .ZN(n7437)
         );
  OAI21_X1 U9043 ( .B1(n9510), .B2(n7590), .A(n7437), .ZN(n7438) );
  AOI21_X1 U9044 ( .B1(n9512), .B2(n7595), .A(n7438), .ZN(n7439) );
  OAI21_X1 U9045 ( .B1(n7440), .B2(n9514), .A(n7439), .ZN(P1_U3219) );
  NAND2_X1 U9046 ( .A1(n7444), .A2(n7443), .ZN(n7445) );
  NAND2_X1 U9047 ( .A1(n10356), .A2(n8622), .ZN(n7446) );
  INV_X1 U9048 ( .A(n7452), .ZN(n7447) );
  NAND2_X1 U9049 ( .A1(n7448), .A2(n7452), .ZN(n7449) );
  NAND2_X1 U9050 ( .A1(n7503), .A2(n7449), .ZN(n10441) );
  NAND2_X1 U9051 ( .A1(n10441), .A2(n9250), .ZN(n7457) );
  OAI21_X1 U9052 ( .B1(n7452), .B2(n7451), .A(n7450), .ZN(n7455) );
  OAI22_X1 U9053 ( .A1(n7453), .A2(n9242), .B1(n7736), .B2(n9240), .ZN(n7454)
         );
  AOI21_X1 U9054 ( .B1(n7455), .B2(n10371), .A(n7454), .ZN(n7456) );
  INV_X1 U9055 ( .A(n10356), .ZN(n10431) );
  NAND2_X1 U9056 ( .A1(n10358), .A2(n10431), .ZN(n10357) );
  NAND2_X1 U9057 ( .A1(n10357), .A2(n10436), .ZN(n7459) );
  NAND2_X1 U9058 ( .A1(n4572), .A2(n7459), .ZN(n10438) );
  INV_X1 U9059 ( .A(n9262), .ZN(n8678) );
  OAI22_X1 U9060 ( .A1(n9259), .A2(n7461), .B1(n7460), .B2(n9256), .ZN(n7462)
         );
  AOI21_X1 U9061 ( .B1(n10355), .B2(n10436), .A(n7462), .ZN(n7463) );
  OAI21_X1 U9062 ( .B1(n10438), .B2(n8678), .A(n7463), .ZN(n7464) );
  AOI21_X1 U9063 ( .B1(n10441), .B2(n9263), .A(n7464), .ZN(n7465) );
  OAI21_X1 U9064 ( .B1(n10443), .B2(n10372), .A(n7465), .ZN(P2_U3287) );
  NAND2_X1 U9065 ( .A1(n7716), .A2(n10168), .ZN(n8048) );
  OR2_X1 U9066 ( .A1(n7466), .A2(n9526), .ZN(n7467) );
  NAND2_X1 U9067 ( .A1(n7468), .A2(n7467), .ZN(n7522) );
  INV_X1 U9068 ( .A(n9525), .ZN(n7586) );
  OR2_X1 U9069 ( .A1(n7532), .A2(n7586), .ZN(n8038) );
  NAND2_X1 U9070 ( .A1(n7532), .A2(n7586), .ZN(n8032) );
  NAND2_X1 U9071 ( .A1(n8038), .A2(n8032), .ZN(n8125) );
  OR2_X1 U9072 ( .A1(n7532), .A2(n9525), .ZN(n7469) );
  INV_X1 U9073 ( .A(n9524), .ZN(n10169) );
  OR2_X1 U9074 ( .A1(n7595), .A2(n10169), .ZN(n8184) );
  NAND2_X1 U9075 ( .A1(n7595), .A2(n10169), .ZN(n8045) );
  NAND2_X1 U9076 ( .A1(n8184), .A2(n8045), .ZN(n8126) );
  NAND2_X1 U9077 ( .A1(n7595), .A2(n9524), .ZN(n7470) );
  NAND2_X1 U9078 ( .A1(n7471), .A2(n7470), .ZN(n10159) );
  OR2_X1 U9079 ( .A1(n7491), .A2(n9523), .ZN(n7472) );
  NAND2_X1 U9080 ( .A1(n7491), .A2(n9523), .ZN(n7473) );
  INV_X1 U9081 ( .A(n8130), .ZN(n7474) );
  INV_X1 U9082 ( .A(n7718), .ZN(n7475) );
  AOI21_X1 U9083 ( .B1(n8130), .B2(n7476), .A(n7475), .ZN(n7578) );
  INV_X1 U9084 ( .A(n7532), .ZN(n10214) );
  INV_X1 U9085 ( .A(n7595), .ZN(n10220) );
  INV_X1 U9086 ( .A(n7491), .ZN(n10227) );
  INV_X1 U9087 ( .A(n9962), .ZN(n7477) );
  AOI211_X1 U9088 ( .C1(n7716), .C2(n10160), .A(n10228), .B(n7477), .ZN(n7576)
         );
  NOR2_X1 U9089 ( .A1(n7478), .A2(n4695), .ZN(n9775) );
  INV_X1 U9090 ( .A(n7716), .ZN(n7479) );
  NOR2_X1 U9091 ( .A1(n7479), .A2(n10177), .ZN(n7482) );
  OAI22_X1 U9092 ( .A1(n10181), .A2(n7480), .B1(n7544), .B2(n10178), .ZN(n7481) );
  AOI211_X1 U9093 ( .C1(n7576), .C2(n9775), .A(n7482), .B(n7481), .ZN(n7494)
         );
  INV_X1 U9094 ( .A(n9521), .ZN(n7769) );
  NAND2_X1 U9095 ( .A1(n8031), .A2(n7483), .ZN(n8251) );
  INV_X1 U9096 ( .A(n8251), .ZN(n8175) );
  NAND2_X1 U9097 ( .A1(n7484), .A2(n8175), .ZN(n7488) );
  AND2_X1 U9098 ( .A1(n8031), .A2(n7485), .ZN(n8165) );
  INV_X1 U9099 ( .A(n8122), .ZN(n7486) );
  NOR2_X1 U9100 ( .A1(n8165), .A2(n7486), .ZN(n7487) );
  NAND2_X1 U9101 ( .A1(n7488), .A2(n7487), .ZN(n7524) );
  NAND2_X1 U9102 ( .A1(n8045), .A2(n8032), .ZN(n8039) );
  INV_X1 U9103 ( .A(n8039), .ZN(n8159) );
  NAND2_X1 U9104 ( .A1(n7583), .A2(n8159), .ZN(n7489) );
  OR2_X1 U9105 ( .A1(n7491), .A2(n7585), .ZN(n8129) );
  INV_X1 U9106 ( .A(n8129), .ZN(n7490) );
  NAND2_X1 U9107 ( .A1(n7491), .A2(n7585), .ZN(n8128) );
  XOR2_X1 U9108 ( .A(n8130), .B(n7723), .Z(n7492) );
  OAI222_X1 U9109 ( .A1(n10167), .A2(n7769), .B1(n10170), .B2(n7585), .C1(
        n7492), .C2(n9949), .ZN(n7575) );
  NAND2_X1 U9110 ( .A1(n7575), .A2(n10181), .ZN(n7493) );
  OAI211_X1 U9111 ( .C1(n7578), .C2(n9777), .A(n7494), .B(n7493), .ZN(P1_U3281) );
  XNOR2_X1 U9112 ( .A(n7495), .B(n7504), .ZN(n7497) );
  OR2_X1 U9113 ( .A1(n7501), .A2(n9242), .ZN(n7496) );
  OAI21_X1 U9114 ( .B1(n7744), .B2(n9240), .A(n7496), .ZN(n7612) );
  AOI21_X1 U9115 ( .B1(n7497), .B2(n10371), .A(n7612), .ZN(n10452) );
  AND2_X1 U9116 ( .A1(n4572), .A2(n10445), .ZN(n7498) );
  NOR2_X1 U9117 ( .A1(n7755), .A2(n7498), .ZN(n10448) );
  INV_X1 U9118 ( .A(n10445), .ZN(n7615) );
  NOR2_X1 U9119 ( .A1(n7615), .A2(n9254), .ZN(n7500) );
  OAI22_X1 U9120 ( .A1(n9259), .A2(n6991), .B1(n7610), .B2(n9256), .ZN(n7499)
         );
  AOI211_X1 U9121 ( .C1(n10448), .C2(n9262), .A(n7500), .B(n7499), .ZN(n7507)
         );
  INV_X1 U9122 ( .A(n7501), .ZN(n8621) );
  OR2_X1 U9123 ( .A1(n10436), .A2(n8621), .ZN(n7502) );
  NAND2_X1 U9124 ( .A1(n7503), .A2(n7502), .ZN(n7505) );
  NAND2_X1 U9125 ( .A1(n7505), .A2(n7504), .ZN(n10446) );
  NAND3_X1 U9126 ( .A1(n7738), .A2(n10446), .A3(n10381), .ZN(n7506) );
  OAI211_X1 U9127 ( .C1(n10452), .C2(n10372), .A(n7507), .B(n7506), .ZN(
        P2_U3286) );
  INV_X1 U9128 ( .A(n7508), .ZN(n7519) );
  OAI222_X1 U9129 ( .A1(n9886), .A2(n7519), .B1(P1_U3084), .B2(n8236), .C1(
        n8749), .C2(n9891), .ZN(P1_U3332) );
  OAI21_X1 U9130 ( .B1(n7511), .B2(n7510), .A(n7509), .ZN(n7512) );
  NAND2_X1 U9131 ( .A1(n7512), .A2(n9483), .ZN(n7517) );
  OAI22_X1 U9132 ( .A1(n9486), .A2(n10168), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7513), .ZN(n7515) );
  NOR2_X1 U9133 ( .A1(n9510), .A2(n10179), .ZN(n7514) );
  AOI211_X1 U9134 ( .C1(n9495), .C2(n9524), .A(n7515), .B(n7514), .ZN(n7516)
         );
  OAI211_X1 U9135 ( .C1(n10227), .C2(n9492), .A(n7517), .B(n7516), .ZN(
        P1_U3229) );
  OAI222_X1 U9136 ( .A1(n7520), .A2(P2_U3152), .B1(n9376), .B2(n7519), .C1(
        n7518), .C2(n9382), .ZN(P2_U3337) );
  OAI21_X1 U9137 ( .B1(n7522), .B2(n8125), .A(n7521), .ZN(n10217) );
  INV_X1 U9138 ( .A(n10217), .ZN(n7536) );
  INV_X1 U9139 ( .A(n7583), .ZN(n7523) );
  AOI21_X1 U9140 ( .B1(n8125), .B2(n7524), .A(n7523), .ZN(n7525) );
  OAI222_X1 U9141 ( .A1(n10167), .A2(n10169), .B1(n10170), .B2(n7526), .C1(
        n9949), .C2(n7525), .ZN(n10215) );
  INV_X1 U9142 ( .A(n7591), .ZN(n7527) );
  OAI211_X1 U9143 ( .C1(n10214), .C2(n7528), .A(n7527), .B(n9984), .ZN(n10213)
         );
  INV_X1 U9144 ( .A(n9775), .ZN(n7730) );
  OAI22_X1 U9145 ( .A1(n10181), .A2(n7530), .B1(n7529), .B2(n10178), .ZN(n7531) );
  AOI21_X1 U9146 ( .B1(n9957), .B2(n7532), .A(n7531), .ZN(n7533) );
  OAI21_X1 U9147 ( .B1(n10213), .B2(n7730), .A(n7533), .ZN(n7534) );
  AOI21_X1 U9148 ( .B1(n10215), .B2(n10181), .A(n7534), .ZN(n7535) );
  OAI21_X1 U9149 ( .B1(n7536), .B2(n9777), .A(n7535), .ZN(P1_U3284) );
  XNOR2_X1 U9150 ( .A(n7539), .B(n7538), .ZN(n7540) );
  XNOR2_X1 U9151 ( .A(n7537), .B(n7540), .ZN(n7547) );
  NOR2_X1 U9152 ( .A1(n9505), .A2(n7585), .ZN(n7541) );
  AOI211_X1 U9153 ( .C1(n9507), .C2(n9521), .A(n7542), .B(n7541), .ZN(n7543)
         );
  OAI21_X1 U9154 ( .B1(n9510), .B2(n7544), .A(n7543), .ZN(n7545) );
  AOI21_X1 U9155 ( .B1(n9512), .B2(n7716), .A(n7545), .ZN(n7546) );
  OAI21_X1 U9156 ( .B1(n7547), .B2(n9514), .A(n7546), .ZN(P1_U3215) );
  OAI22_X1 U9157 ( .A1(n10181), .A2(n7549), .B1(n7548), .B2(n10178), .ZN(n7552) );
  INV_X1 U9158 ( .A(n10163), .ZN(n7904) );
  NOR2_X1 U9159 ( .A1(n7904), .A2(n7550), .ZN(n7551) );
  AOI211_X1 U9160 ( .C1(n9957), .C2(n7553), .A(n7552), .B(n7551), .ZN(n7556)
         );
  NAND2_X1 U9161 ( .A1(n7554), .A2(n10181), .ZN(n7555) );
  OAI211_X1 U9162 ( .C1(n7557), .C2(n7735), .A(n7556), .B(n7555), .ZN(P1_U3289) );
  OAI21_X1 U9163 ( .B1(n7559), .B2(n8120), .A(n7558), .ZN(n10205) );
  INV_X1 U9164 ( .A(n10205), .ZN(n7574) );
  OAI22_X1 U9165 ( .A1(n10181), .A2(n5920), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10178), .ZN(n7563) );
  OAI21_X1 U9166 ( .B1(n7561), .B2(n10201), .A(n7560), .ZN(n10202) );
  NOR2_X1 U9167 ( .A1(n7904), .A2(n10202), .ZN(n7562) );
  AOI211_X1 U9168 ( .C1(n9957), .C2(n7564), .A(n7563), .B(n7562), .ZN(n7573)
         );
  OAI21_X1 U9169 ( .B1(n7566), .B2(n8166), .A(n7565), .ZN(n7570) );
  OAI22_X1 U9170 ( .A1(n10170), .A2(n7568), .B1(n7567), .B2(n10167), .ZN(n7569) );
  AOI21_X1 U9171 ( .B1(n7570), .B2(n10172), .A(n7569), .ZN(n7571) );
  OAI21_X1 U9172 ( .B1(n7574), .B2(n10175), .A(n7571), .ZN(n10203) );
  NAND2_X1 U9173 ( .A1(n10203), .A2(n10181), .ZN(n7572) );
  OAI211_X1 U9174 ( .C1(n7574), .C2(n7735), .A(n7573), .B(n7572), .ZN(P1_U3288) );
  AOI211_X1 U9175 ( .C1(n7716), .C2(n9849), .A(n7576), .B(n7575), .ZN(n7577)
         );
  OAI21_X1 U9176 ( .B1(n7578), .B2(n9853), .A(n7577), .ZN(n7580) );
  NAND2_X1 U9177 ( .A1(n7580), .A2(n10245), .ZN(n7579) );
  OAI21_X1 U9178 ( .B1(n10245), .B2(n6125), .A(n7579), .ZN(P1_U3533) );
  NAND2_X1 U9179 ( .A1(n7580), .A2(n10236), .ZN(n7581) );
  OAI21_X1 U9180 ( .B1(n10236), .B2(n6124), .A(n7581), .ZN(P1_U3484) );
  XNOR2_X1 U9181 ( .A(n7582), .B(n4823), .ZN(n10219) );
  NAND2_X1 U9182 ( .A1(n7583), .A2(n8032), .ZN(n7584) );
  XNOR2_X1 U9183 ( .A(n7584), .B(n4823), .ZN(n7588) );
  OAI22_X1 U9184 ( .A1(n10170), .A2(n7586), .B1(n7585), .B2(n10167), .ZN(n7587) );
  AOI21_X1 U9185 ( .B1(n7588), .B2(n10172), .A(n7587), .ZN(n7589) );
  OAI21_X1 U9186 ( .B1(n10219), .B2(n10175), .A(n7589), .ZN(n10222) );
  NAND2_X1 U9187 ( .A1(n10222), .A2(n10181), .ZN(n7597) );
  OAI22_X1 U9188 ( .A1(n10181), .A2(n8772), .B1(n7590), .B2(n10178), .ZN(n7594) );
  NOR2_X1 U9189 ( .A1(n7591), .A2(n10220), .ZN(n7592) );
  OR2_X1 U9190 ( .A1(n10161), .A2(n7592), .ZN(n10221) );
  NOR2_X1 U9191 ( .A1(n10221), .A2(n7904), .ZN(n7593) );
  AOI211_X1 U9192 ( .C1(n9957), .C2(n7595), .A(n7594), .B(n7593), .ZN(n7596)
         );
  OAI211_X1 U9193 ( .C1(n10219), .C2(n7735), .A(n7597), .B(n7596), .ZN(
        P1_U3283) );
  NAND2_X1 U9194 ( .A1(n7599), .A2(n7598), .ZN(n7601) );
  XNOR2_X1 U9195 ( .A(n10445), .B(n8343), .ZN(n7602) );
  NOR2_X1 U9196 ( .A1(n7736), .A2(n8341), .ZN(n7603) );
  NAND2_X1 U9197 ( .A1(n7602), .A2(n7603), .ZN(n7652) );
  INV_X1 U9198 ( .A(n7602), .ZN(n7651) );
  INV_X1 U9199 ( .A(n7603), .ZN(n7604) );
  NAND2_X1 U9200 ( .A1(n7651), .A2(n7604), .ZN(n7605) );
  NAND2_X1 U9201 ( .A1(n7652), .A2(n7605), .ZN(n7607) );
  AOI21_X1 U9202 ( .B1(n7606), .B2(n7607), .A(n10246), .ZN(n7609) );
  NAND2_X1 U9203 ( .A1(n7609), .A2(n7653), .ZN(n7614) );
  AND2_X1 U9204 ( .A1(P2_U3152), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n10327) );
  NOR2_X1 U9205 ( .A1(n10292), .A2(n7610), .ZN(n7611) );
  AOI211_X1 U9206 ( .C1(n10279), .C2(n7612), .A(n10327), .B(n7611), .ZN(n7613)
         );
  OAI211_X1 U9207 ( .C1(n7615), .C2(n4871), .A(n7614), .B(n7613), .ZN(P2_U3219) );
  AOI22_X1 U9208 ( .A1(n7667), .A2(n7616), .B1(P2_REG1_REG_16__SCAN_IN), .B2(
        n7623), .ZN(n7621) );
  NAND2_X1 U9209 ( .A1(n7625), .A2(n7617), .ZN(n7619) );
  NAND2_X1 U9210 ( .A1(n7619), .A2(n7618), .ZN(n7620) );
  NOR2_X1 U9211 ( .A1(n7621), .A2(n7620), .ZN(n7669) );
  AOI21_X1 U9212 ( .B1(n7621), .B2(n7620), .A(n7669), .ZN(n7634) );
  INV_X1 U9213 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n7622) );
  NAND2_X1 U9214 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3152), .ZN(n7981) );
  OAI21_X1 U9215 ( .B1(n10304), .B2(n7622), .A(n7981), .ZN(n7632) );
  AOI22_X1 U9216 ( .A1(n7667), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n9258), .B2(
        n7623), .ZN(n7629) );
  NOR2_X1 U9217 ( .A1(n7625), .A2(n7624), .ZN(n7627) );
  OAI21_X1 U9218 ( .B1(n7629), .B2(n7628), .A(n7663), .ZN(n7630) );
  NOR2_X1 U9219 ( .A1(n7630), .A2(n10295), .ZN(n7631) );
  AOI211_X1 U9220 ( .C1(n10330), .C2(n7667), .A(n7632), .B(n7631), .ZN(n7633)
         );
  OAI21_X1 U9221 ( .B1(n7634), .B2(n10294), .A(n7633), .ZN(P2_U3261) );
  INV_X1 U9222 ( .A(n7635), .ZN(n8473) );
  OAI222_X1 U9223 ( .A1(P2_U3152), .A2(n7637), .B1(n9376), .B2(n8473), .C1(
        n7636), .C2(n9382), .ZN(P2_U3336) );
  XNOR2_X1 U9224 ( .A(n7638), .B(n7639), .ZN(n7645) );
  NOR2_X1 U9225 ( .A1(n9505), .A2(n10168), .ZN(n7640) );
  AOI211_X1 U9226 ( .C1(n9507), .C2(n9944), .A(n7641), .B(n7640), .ZN(n7642)
         );
  OAI21_X1 U9227 ( .B1(n9510), .B2(n9974), .A(n7642), .ZN(n7643) );
  AOI21_X1 U9228 ( .B1(n9512), .B2(n9973), .A(n7643), .ZN(n7644) );
  OAI21_X1 U9229 ( .B1(n7645), .B2(n9514), .A(n7644), .ZN(P1_U3234) );
  INV_X1 U9230 ( .A(n7758), .ZN(n7802) );
  XNOR2_X1 U9231 ( .A(n7758), .B(n8343), .ZN(n10264) );
  NOR2_X1 U9232 ( .A1(n7744), .A2(n8341), .ZN(n7646) );
  NAND2_X1 U9233 ( .A1(n10264), .A2(n7646), .ZN(n7809) );
  INV_X1 U9234 ( .A(n10264), .ZN(n7648) );
  INV_X1 U9235 ( .A(n7646), .ZN(n7647) );
  NAND2_X1 U9236 ( .A1(n7648), .A2(n7647), .ZN(n7649) );
  AND2_X1 U9237 ( .A1(n7809), .A2(n7649), .ZN(n7654) );
  INV_X1 U9238 ( .A(n7654), .ZN(n7650) );
  AOI21_X1 U9239 ( .B1(n7653), .B2(n7650), .A(n10246), .ZN(n7657) );
  NOR3_X1 U9240 ( .A1(n7651), .A2(n7736), .A3(n8603), .ZN(n7656) );
  OAI21_X1 U9241 ( .B1(n7657), .B2(n7656), .A(n10265), .ZN(n7662) );
  INV_X1 U9242 ( .A(n7658), .ZN(n7800) );
  INV_X1 U9243 ( .A(n10257), .ZN(n10252) );
  INV_X1 U9244 ( .A(n10260), .ZN(n8610) );
  AOI22_X1 U9245 ( .A1(n8610), .A2(n8619), .B1(P2_REG3_REG_11__SCAN_IN), .B2(
        P2_U3152), .ZN(n7659) );
  OAI21_X1 U9246 ( .B1(n7736), .B2(n10252), .A(n7659), .ZN(n7660) );
  AOI21_X1 U9247 ( .B1(n7800), .B2(n8597), .A(n7660), .ZN(n7661) );
  OAI211_X1 U9248 ( .C1(n7802), .C2(n4871), .A(n7662), .B(n7661), .ZN(P2_U3238) );
  AOI22_X1 U9249 ( .A1(n7673), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n9226), .B2(
        n8646), .ZN(n7666) );
  NAND2_X1 U9250 ( .A1(n7667), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n7664) );
  OAI21_X1 U9251 ( .B1(n7666), .B2(n7665), .A(n8642), .ZN(n7676) );
  NOR2_X1 U9252 ( .A1(n7667), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n7668) );
  NOR2_X1 U9253 ( .A1(n7669), .A2(n7668), .ZN(n7671) );
  XNOR2_X1 U9254 ( .A(n7673), .B(n8647), .ZN(n7670) );
  NAND2_X1 U9255 ( .A1(n7670), .A2(n7671), .ZN(n8645) );
  OAI211_X1 U9256 ( .C1(n7671), .C2(n7670), .A(n10336), .B(n8645), .ZN(n7675)
         );
  INV_X1 U9257 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n8915) );
  NAND2_X1 U9258 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8530) );
  OAI21_X1 U9259 ( .B1(n10304), .B2(n8915), .A(n8530), .ZN(n7672) );
  AOI21_X1 U9260 ( .B1(n10330), .B2(n7673), .A(n7672), .ZN(n7674) );
  OAI211_X1 U9261 ( .C1(n7676), .C2(n10295), .A(n7675), .B(n7674), .ZN(
        P2_U3262) );
  INV_X1 U9262 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10510) );
  NOR2_X1 U9263 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7677) );
  AOI21_X1 U9264 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7677), .ZN(n10480) );
  NOR2_X1 U9265 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7678) );
  AOI21_X1 U9266 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7678), .ZN(n10483) );
  NOR2_X1 U9267 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7679) );
  AOI21_X1 U9268 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7679), .ZN(n10486) );
  NOR2_X1 U9269 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7680) );
  AOI21_X1 U9270 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7680), .ZN(n10489) );
  NOR2_X1 U9271 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7681) );
  AOI21_X1 U9272 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7681), .ZN(n10492) );
  NOR2_X1 U9273 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7689) );
  INV_X1 U9274 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n7682) );
  AOI22_X1 U9275 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n7682), .B1(
        P2_ADDR_REG_4__SCAN_IN), .B2(n8810), .ZN(n10520) );
  NAND2_X1 U9276 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n7687) );
  INV_X1 U9277 ( .A(P2_ADDR_REG_3__SCAN_IN), .ZN(n10303) );
  AOI22_X1 U9278 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .B1(n10303), .B2(n8859), .ZN(n10518) );
  NAND2_X1 U9279 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n7685) );
  XOR2_X1 U9280 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Z(
        n10504) );
  AOI21_X1 U9281 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10474) );
  INV_X1 U9282 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7683) );
  NAND3_X1 U9283 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_1__SCAN_IN), .ZN(n10476) );
  OAI21_X1 U9284 ( .B1(n10474), .B2(n7683), .A(n10476), .ZN(n10503) );
  NAND2_X1 U9285 ( .A1(n10504), .A2(n10503), .ZN(n7684) );
  NAND2_X1 U9286 ( .A1(n7685), .A2(n7684), .ZN(n10517) );
  NAND2_X1 U9287 ( .A1(n10518), .A2(n10517), .ZN(n7686) );
  NAND2_X1 U9288 ( .A1(n7687), .A2(n7686), .ZN(n10519) );
  NOR2_X1 U9289 ( .A1(n10520), .A2(n10519), .ZN(n7688) );
  NOR2_X1 U9290 ( .A1(n7689), .A2(n7688), .ZN(n7690) );
  NOR2_X1 U9291 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7690), .ZN(n10506) );
  AND2_X1 U9292 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n7690), .ZN(n10505) );
  NOR2_X1 U9293 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10505), .ZN(n7691) );
  NOR2_X1 U9294 ( .A1(n10506), .A2(n7691), .ZN(n7692) );
  NAND2_X1 U9295 ( .A1(n7692), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7694) );
  XOR2_X1 U9296 ( .A(n7692), .B(P1_ADDR_REG_6__SCAN_IN), .Z(n10502) );
  NAND2_X1 U9297 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10502), .ZN(n7693) );
  NAND2_X1 U9298 ( .A1(n7694), .A2(n7693), .ZN(n7695) );
  NAND2_X1 U9299 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n7695), .ZN(n7697) );
  XNOR2_X1 U9300 ( .A(n8831), .B(n7695), .ZN(n10515) );
  NAND2_X1 U9301 ( .A1(n10515), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7696) );
  NAND2_X1 U9302 ( .A1(n7697), .A2(n7696), .ZN(n7698) );
  NAND2_X1 U9303 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n7698), .ZN(n7700) );
  XOR2_X1 U9304 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n7698), .Z(n10516) );
  NAND2_X1 U9305 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10516), .ZN(n7699) );
  NAND2_X1 U9306 ( .A1(n7700), .A2(n7699), .ZN(n7701) );
  AND2_X1 U9307 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n7701), .ZN(n7702) );
  INV_X1 U9308 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10514) );
  XNOR2_X1 U9309 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n7701), .ZN(n10513) );
  NAND2_X1 U9310 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7703) );
  OAI21_X1 U9311 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n7703), .ZN(n10500) );
  NAND2_X1 U9312 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n7704) );
  OAI21_X1 U9313 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7704), .ZN(n10497) );
  AOI21_X1 U9314 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10496), .ZN(n10495) );
  NOR2_X1 U9315 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7705) );
  AOI21_X1 U9316 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7705), .ZN(n10494) );
  NAND2_X1 U9317 ( .A1(n10495), .A2(n10494), .ZN(n10493) );
  OAI21_X1 U9318 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10493), .ZN(n10491) );
  NAND2_X1 U9319 ( .A1(n10492), .A2(n10491), .ZN(n10490) );
  OAI21_X1 U9320 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10490), .ZN(n10488) );
  NAND2_X1 U9321 ( .A1(n10489), .A2(n10488), .ZN(n10487) );
  OAI21_X1 U9322 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10487), .ZN(n10485) );
  NAND2_X1 U9323 ( .A1(n10486), .A2(n10485), .ZN(n10484) );
  OAI21_X1 U9324 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10484), .ZN(n10482) );
  NAND2_X1 U9325 ( .A1(n10483), .A2(n10482), .ZN(n10481) );
  OAI21_X1 U9326 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10481), .ZN(n10479) );
  NAND2_X1 U9327 ( .A1(n10480), .A2(n10479), .ZN(n10478) );
  OAI21_X1 U9328 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10478), .ZN(n10509) );
  NOR2_X1 U9329 ( .A1(n10510), .A2(n10509), .ZN(n7706) );
  NAND2_X1 U9330 ( .A1(n10510), .A2(n10509), .ZN(n10508) );
  OAI21_X1 U9331 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n7706), .A(n10508), .ZN(
        n7708) );
  XNOR2_X1 U9332 ( .A(n8671), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7707) );
  XNOR2_X1 U9333 ( .A(n7708), .B(n7707), .ZN(ADD_1071_U4) );
  NAND2_X1 U9334 ( .A1(n7712), .A2(n9378), .ZN(n7710) );
  OAI211_X1 U9335 ( .C1(n7711), .C2(n9382), .A(n7710), .B(n7709), .ZN(P2_U3335) );
  NAND2_X1 U9336 ( .A1(n7712), .A2(n9892), .ZN(n7714) );
  NAND2_X1 U9337 ( .A1(n7713), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8276) );
  OAI211_X1 U9338 ( .C1(n7715), .C2(n9891), .A(n7714), .B(n8276), .ZN(P1_U3330) );
  OR2_X1 U9339 ( .A1(n7716), .A2(n9522), .ZN(n7717) );
  NAND2_X1 U9340 ( .A1(n7718), .A2(n7717), .ZN(n9961) );
  NAND2_X1 U9341 ( .A1(n9973), .A2(n9521), .ZN(n8052) );
  OR2_X1 U9342 ( .A1(n9973), .A2(n9521), .ZN(n8053) );
  INV_X1 U9343 ( .A(n8053), .ZN(n7719) );
  INV_X1 U9344 ( .A(n9944), .ZN(n9968) );
  OR2_X1 U9345 ( .A1(n7779), .A2(n9968), .ZN(n8056) );
  NAND2_X1 U9346 ( .A1(n7779), .A2(n9968), .ZN(n8154) );
  NAND2_X1 U9347 ( .A1(n8056), .A2(n8154), .ZN(n8133) );
  OR2_X1 U9348 ( .A1(n7720), .A2(n8133), .ZN(n7721) );
  NAND2_X1 U9349 ( .A1(n7781), .A2(n7721), .ZN(n9991) );
  INV_X1 U9350 ( .A(n8048), .ZN(n7722) );
  NAND2_X1 U9351 ( .A1(n9973), .A2(n7769), .ZN(n8153) );
  NAND2_X1 U9352 ( .A1(n9967), .A2(n8153), .ZN(n7789) );
  OR2_X1 U9353 ( .A1(n9973), .A2(n7769), .ZN(n7787) );
  NAND2_X1 U9354 ( .A1(n7789), .A2(n7787), .ZN(n7724) );
  XNOR2_X1 U9355 ( .A(n7724), .B(n8133), .ZN(n7726) );
  INV_X1 U9356 ( .A(n9520), .ZN(n7911) );
  OAI22_X1 U9357 ( .A1(n10170), .A2(n7769), .B1(n7911), .B2(n10167), .ZN(n7725) );
  AOI21_X1 U9358 ( .B1(n7726), .B2(n10172), .A(n7725), .ZN(n7727) );
  OAI21_X1 U9359 ( .B1(n9991), .B2(n10175), .A(n7727), .ZN(n9994) );
  NAND2_X1 U9360 ( .A1(n9994), .A2(n10181), .ZN(n7734) );
  OAI22_X1 U9361 ( .A1(n10181), .A2(n7728), .B1(n7772), .B2(n10178), .ZN(n7732) );
  INV_X1 U9362 ( .A(n7779), .ZN(n9993) );
  NOR2_X1 U9363 ( .A1(n9962), .A2(n9973), .ZN(n9963) );
  INV_X1 U9364 ( .A(n9936), .ZN(n7729) );
  OAI211_X1 U9365 ( .C1(n9993), .C2(n9963), .A(n7729), .B(n9984), .ZN(n9992)
         );
  NOR2_X1 U9366 ( .A1(n9992), .A2(n7730), .ZN(n7731) );
  AOI211_X1 U9367 ( .C1(n9957), .C2(n7779), .A(n7732), .B(n7731), .ZN(n7733)
         );
  OAI211_X1 U9368 ( .C1(n9991), .C2(n7735), .A(n7734), .B(n7733), .ZN(P1_U3279) );
  INV_X1 U9369 ( .A(n7736), .ZN(n8620) );
  NAND2_X1 U9370 ( .A1(n10445), .A2(n8620), .ZN(n7737) );
  INV_X1 U9371 ( .A(n7744), .ZN(n10262) );
  OR2_X1 U9372 ( .A1(n7758), .A2(n10262), .ZN(n7739) );
  NAND2_X1 U9373 ( .A1(n7758), .A2(n10262), .ZN(n7740) );
  XNOR2_X1 U9374 ( .A(n7850), .B(n7849), .ZN(n10460) );
  INV_X1 U9375 ( .A(n10460), .ZN(n7750) );
  XNOR2_X1 U9376 ( .A(n7742), .B(n7849), .ZN(n7743) );
  OAI222_X1 U9377 ( .A1(n9242), .A2(n7744), .B1(n9240), .B2(n10261), .C1(n9246), .C2(n7743), .ZN(n10457) );
  INV_X1 U9378 ( .A(n10274), .ZN(n10454) );
  OAI21_X1 U9379 ( .B1(n7756), .B2(n10454), .A(n7878), .ZN(n10456) );
  OAI22_X1 U9380 ( .A1(n9259), .A2(n7745), .B1(n10276), .B2(n9256), .ZN(n7746)
         );
  AOI21_X1 U9381 ( .B1(n10274), .B2(n10355), .A(n7746), .ZN(n7747) );
  OAI21_X1 U9382 ( .B1(n10456), .B2(n8678), .A(n7747), .ZN(n7748) );
  AOI21_X1 U9383 ( .B1(n10457), .B2(n7864), .A(n7748), .ZN(n7749) );
  OAI21_X1 U9384 ( .B1(n9233), .B2(n7750), .A(n7749), .ZN(P2_U3284) );
  INV_X1 U9385 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n7761) );
  XNOR2_X1 U9386 ( .A(n7751), .B(n7753), .ZN(n7808) );
  XOR2_X1 U9387 ( .A(n7752), .B(n7753), .Z(n7754) );
  AOI222_X1 U9388 ( .A1(n10371), .A2(n7754), .B1(n8619), .B2(n10368), .C1(
        n8620), .C2(n10366), .ZN(n7803) );
  INV_X1 U9389 ( .A(n7755), .ZN(n7757) );
  AOI21_X1 U9390 ( .B1(n7758), .B2(n7757), .A(n7756), .ZN(n7806) );
  AOI22_X1 U9391 ( .A1(n7806), .A2(n10447), .B1(n10444), .B2(n7758), .ZN(n7759) );
  OAI211_X1 U9392 ( .C1(n9926), .C2(n7808), .A(n7803), .B(n7759), .ZN(n7762)
         );
  NAND2_X1 U9393 ( .A1(n7762), .A2(n10462), .ZN(n7760) );
  OAI21_X1 U9394 ( .B1(n10462), .B2(n7761), .A(n7760), .ZN(P2_U3484) );
  NAND2_X1 U9395 ( .A1(n7762), .A2(n10473), .ZN(n7763) );
  OAI21_X1 U9396 ( .B1(n10473), .B2(n7001), .A(n7763), .ZN(P2_U3531) );
  NAND2_X1 U9397 ( .A1(n7765), .A2(n7764), .ZN(n7767) );
  XOR2_X1 U9398 ( .A(n7767), .B(n7766), .Z(n7775) );
  NOR2_X1 U9399 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7768), .ZN(n10083) );
  NOR2_X1 U9400 ( .A1(n9505), .A2(n7769), .ZN(n7770) );
  AOI211_X1 U9401 ( .C1(n9507), .C2(n9520), .A(n10083), .B(n7770), .ZN(n7771)
         );
  OAI21_X1 U9402 ( .B1(n9510), .B2(n7772), .A(n7771), .ZN(n7773) );
  AOI21_X1 U9403 ( .B1(n9512), .B2(n7779), .A(n7773), .ZN(n7774) );
  OAI21_X1 U9404 ( .B1(n7775), .B2(n9514), .A(n7774), .ZN(P1_U3222) );
  INV_X1 U9405 ( .A(n7776), .ZN(n7798) );
  OAI222_X1 U9406 ( .A1(n9886), .A2(n7798), .B1(P1_U3084), .B2(n7778), .C1(
        n7777), .C2(n9891), .ZN(P1_U3329) );
  NAND2_X1 U9407 ( .A1(n7779), .A2(n9944), .ZN(n7780) );
  OR2_X1 U9408 ( .A1(n9956), .A2(n9520), .ZN(n7782) );
  INV_X1 U9409 ( .A(n9946), .ZN(n9504) );
  NAND2_X1 U9410 ( .A1(n7917), .A2(n9504), .ZN(n8151) );
  NAND2_X1 U9411 ( .A1(n8064), .A2(n8151), .ZN(n8134) );
  XNOR2_X1 U9412 ( .A(n7888), .B(n8134), .ZN(n7844) );
  INV_X1 U9413 ( .A(n9956), .ZN(n9985) );
  INV_X1 U9414 ( .A(n7899), .ZN(n7783) );
  AOI211_X1 U9415 ( .C1(n7917), .C2(n9938), .A(n10228), .B(n7783), .ZN(n7841)
         );
  INV_X1 U9416 ( .A(n7917), .ZN(n7786) );
  INV_X1 U9417 ( .A(n7915), .ZN(n7784) );
  AOI22_X1 U9418 ( .A1(n9953), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n7784), .B2(
        n9763), .ZN(n7785) );
  OAI21_X1 U9419 ( .B1(n7786), .B2(n10177), .A(n7785), .ZN(n7795) );
  NAND2_X1 U9420 ( .A1(n8056), .A2(n7787), .ZN(n8055) );
  INV_X1 U9421 ( .A(n8055), .ZN(n7788) );
  NAND2_X1 U9422 ( .A1(n7789), .A2(n7788), .ZN(n7790) );
  OR2_X1 U9423 ( .A1(n9956), .A2(n7911), .ZN(n8054) );
  NAND2_X1 U9424 ( .A1(n9956), .A2(n7911), .ZN(n8187) );
  NAND2_X1 U9425 ( .A1(n8054), .A2(n8187), .ZN(n9942) );
  INV_X1 U9426 ( .A(n9942), .ZN(n9934) );
  AOI21_X1 U9427 ( .B1(n7791), .B2(n8134), .A(n9949), .ZN(n7793) );
  INV_X1 U9428 ( .A(n9770), .ZN(n9438) );
  OAI22_X1 U9429 ( .A1(n10170), .A2(n7911), .B1(n9438), .B2(n10167), .ZN(n7792) );
  AOI21_X1 U9430 ( .B1(n7793), .B2(n7893), .A(n7792), .ZN(n7843) );
  NOR2_X1 U9431 ( .A1(n7843), .A2(n9953), .ZN(n7794) );
  AOI211_X1 U9432 ( .C1(n7841), .C2(n9775), .A(n7795), .B(n7794), .ZN(n7796)
         );
  OAI21_X1 U9433 ( .B1(n7844), .B2(n9777), .A(n7796), .ZN(P1_U3277) );
  OAI222_X1 U9434 ( .A1(n7799), .A2(P2_U3152), .B1(n9376), .B2(n7798), .C1(
        n7797), .C2(n9382), .ZN(P2_U3334) );
  AOI22_X1 U9435 ( .A1(n10372), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n7800), .B2(
        n10373), .ZN(n7801) );
  OAI21_X1 U9436 ( .B1(n7802), .B2(n9254), .A(n7801), .ZN(n7805) );
  NOR2_X1 U9437 ( .A1(n7803), .A2(n10372), .ZN(n7804) );
  AOI211_X1 U9438 ( .C1(n7806), .C2(n9262), .A(n7805), .B(n7804), .ZN(n7807)
         );
  OAI21_X1 U9439 ( .B1(n9233), .B2(n7808), .A(n7807), .ZN(P2_U3285) );
  INV_X1 U9440 ( .A(n7932), .ZN(n7881) );
  NAND2_X1 U9441 ( .A1(n10265), .A2(n7809), .ZN(n7814) );
  XNOR2_X1 U9442 ( .A(n10274), .B(n8343), .ZN(n7810) );
  NOR2_X1 U9443 ( .A1(n7873), .A2(n8341), .ZN(n7811) );
  NAND2_X1 U9444 ( .A1(n7810), .A2(n7811), .ZN(n7821) );
  INV_X1 U9445 ( .A(n7810), .ZN(n7820) );
  INV_X1 U9446 ( .A(n7811), .ZN(n7812) );
  NAND2_X1 U9447 ( .A1(n7820), .A2(n7812), .ZN(n7813) );
  AND2_X1 U9448 ( .A1(n7821), .A2(n7813), .ZN(n10266) );
  NAND2_X1 U9449 ( .A1(n7814), .A2(n10266), .ZN(n7822) );
  XNOR2_X1 U9450 ( .A(n7932), .B(n8343), .ZN(n7815) );
  NOR2_X1 U9451 ( .A1(n10261), .A2(n8341), .ZN(n7816) );
  NAND2_X1 U9452 ( .A1(n7815), .A2(n7816), .ZN(n7950) );
  INV_X1 U9453 ( .A(n7815), .ZN(n7943) );
  INV_X1 U9454 ( .A(n7816), .ZN(n7817) );
  NAND2_X1 U9455 ( .A1(n7943), .A2(n7817), .ZN(n7818) );
  AND2_X1 U9456 ( .A1(n7950), .A2(n7818), .ZN(n7823) );
  INV_X1 U9457 ( .A(n7823), .ZN(n7819) );
  AOI21_X1 U9458 ( .B1(n10268), .B2(n7819), .A(n10246), .ZN(n7826) );
  NOR3_X1 U9459 ( .A1(n7820), .A2(n7873), .A3(n8603), .ZN(n7825) );
  NAND2_X1 U9460 ( .A1(n7822), .A2(n7821), .ZN(n7824) );
  OAI21_X1 U9461 ( .B1(n7826), .B2(n7825), .A(n7942), .ZN(n7831) );
  NOR2_X1 U9462 ( .A1(n10292), .A2(n7882), .ZN(n7829) );
  OAI22_X1 U9463 ( .A1(n10260), .A2(n7965), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7827), .ZN(n7828) );
  AOI211_X1 U9464 ( .C1(n10257), .C2(n8619), .A(n7829), .B(n7828), .ZN(n7830)
         );
  OAI211_X1 U9465 ( .C1(n7881), .C2(n4871), .A(n7831), .B(n7830), .ZN(P2_U3236) );
  XOR2_X1 U9466 ( .A(n7834), .B(n7833), .Z(n7835) );
  XNOR2_X1 U9467 ( .A(n7832), .B(n7835), .ZN(n7840) );
  AND2_X1 U9468 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n10096) );
  NOR2_X1 U9469 ( .A1(n9505), .A2(n9968), .ZN(n7836) );
  AOI211_X1 U9470 ( .C1(n9507), .C2(n9946), .A(n10096), .B(n7836), .ZN(n7837)
         );
  OAI21_X1 U9471 ( .B1(n9510), .B2(n9940), .A(n7837), .ZN(n7838) );
  AOI21_X1 U9472 ( .B1(n9956), .B2(n9512), .A(n7838), .ZN(n7839) );
  OAI21_X1 U9473 ( .B1(n7840), .B2(n9514), .A(n7839), .ZN(P1_U3232) );
  AOI21_X1 U9474 ( .B1(n7917), .B2(n9849), .A(n7841), .ZN(n7842) );
  OAI211_X1 U9475 ( .C1(n7844), .C2(n9853), .A(n7843), .B(n7842), .ZN(n7846)
         );
  NAND2_X1 U9476 ( .A1(n7846), .A2(n10245), .ZN(n7845) );
  OAI21_X1 U9477 ( .B1(n10245), .B2(n6200), .A(n7845), .ZN(P1_U3537) );
  INV_X1 U9478 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7848) );
  NAND2_X1 U9479 ( .A1(n7846), .A2(n10236), .ZN(n7847) );
  OAI21_X1 U9480 ( .B1(n10236), .B2(n7848), .A(n7847), .ZN(P1_U3496) );
  INV_X1 U9481 ( .A(n10261), .ZN(n8618) );
  NAND2_X1 U9482 ( .A1(n7932), .A2(n8618), .ZN(n7851) );
  NAND2_X1 U9483 ( .A1(n7869), .A2(n7851), .ZN(n7991) );
  XNOR2_X1 U9484 ( .A(n7991), .B(n4888), .ZN(n9931) );
  INV_X1 U9485 ( .A(n9931), .ZN(n7866) );
  NAND2_X1 U9486 ( .A1(n7852), .A2(n7992), .ZN(n7853) );
  NAND2_X1 U9487 ( .A1(n7853), .A2(n10371), .ZN(n7854) );
  OR2_X1 U9488 ( .A1(n7855), .A2(n7854), .ZN(n7858) );
  OAI22_X1 U9489 ( .A1(n9243), .A2(n9240), .B1(n10261), .B2(n9242), .ZN(n7856)
         );
  INV_X1 U9490 ( .A(n7856), .ZN(n7857) );
  NAND2_X1 U9491 ( .A1(n7858), .A2(n7857), .ZN(n9929) );
  OAI211_X1 U9492 ( .C1(n7859), .C2(n9928), .A(n10447), .B(n8000), .ZN(n9927)
         );
  OAI22_X1 U9493 ( .A1(n9259), .A2(n7860), .B1(n7949), .B2(n9256), .ZN(n7861)
         );
  AOI21_X1 U9494 ( .B1(n7993), .B2(n10355), .A(n7861), .ZN(n7862) );
  OAI21_X1 U9495 ( .B1(n9927), .B2(n10359), .A(n7862), .ZN(n7863) );
  AOI21_X1 U9496 ( .B1(n9929), .B2(n7864), .A(n7863), .ZN(n7865) );
  OAI21_X1 U9497 ( .B1(n7866), .B2(n9233), .A(n7865), .ZN(P2_U3282) );
  NAND2_X1 U9498 ( .A1(n7867), .A2(n7872), .ZN(n7868) );
  NAND2_X1 U9499 ( .A1(n7869), .A2(n7868), .ZN(n7935) );
  OR2_X1 U9500 ( .A1(n7935), .A2(n10349), .ZN(n7877) );
  OAI21_X1 U9501 ( .B1(n7872), .B2(n7871), .A(n7870), .ZN(n7875) );
  OAI22_X1 U9502 ( .A1(n7965), .A2(n9240), .B1(n7873), .B2(n9242), .ZN(n7874)
         );
  AOI21_X1 U9503 ( .B1(n7875), .B2(n10371), .A(n7874), .ZN(n7876) );
  NAND2_X1 U9504 ( .A1(n7877), .A2(n7876), .ZN(n7937) );
  NAND2_X1 U9505 ( .A1(n7937), .A2(n9259), .ZN(n7887) );
  NAND2_X1 U9506 ( .A1(n7878), .A2(n7932), .ZN(n7879) );
  AND2_X1 U9507 ( .A1(n7880), .A2(n7879), .ZN(n7933) );
  NOR2_X1 U9508 ( .A1(n7881), .A2(n9254), .ZN(n7885) );
  OAI22_X1 U9509 ( .A1(n9259), .A2(n7883), .B1(n7882), .B2(n9256), .ZN(n7884)
         );
  AOI211_X1 U9510 ( .C1(n7933), .C2(n9262), .A(n7885), .B(n7884), .ZN(n7886)
         );
  OAI211_X1 U9511 ( .C1(n7935), .C2(n10360), .A(n7887), .B(n7886), .ZN(
        P2_U3283) );
  INV_X1 U9512 ( .A(n7888), .ZN(n7891) );
  AND2_X1 U9513 ( .A1(n7917), .A2(n9946), .ZN(n7889) );
  INV_X1 U9514 ( .A(n7889), .ZN(n7890) );
  OR2_X1 U9515 ( .A1(n7917), .A2(n9946), .ZN(n7892) );
  OR2_X1 U9516 ( .A1(n9856), .A2(n9438), .ZN(n8194) );
  NAND2_X1 U9517 ( .A1(n9856), .A2(n9438), .ZN(n8393) );
  XNOR2_X1 U9518 ( .A(n8365), .B(n7894), .ZN(n9855) );
  NAND2_X1 U9519 ( .A1(n7895), .A2(n7894), .ZN(n7896) );
  AOI21_X1 U9520 ( .B1(n8394), .B2(n7896), .A(n9949), .ZN(n7898) );
  INV_X1 U9521 ( .A(n9751), .ZN(n8029) );
  OAI22_X1 U9522 ( .A1(n10170), .A2(n9504), .B1(n8029), .B2(n10167), .ZN(n7897) );
  AOI211_X1 U9523 ( .C1(n9855), .C2(n9952), .A(n7898), .B(n7897), .ZN(n9861)
         );
  AND2_X1 U9524 ( .A1(n7899), .A2(n9856), .ZN(n7900) );
  OR2_X1 U9525 ( .A1(n7900), .A2(n9760), .ZN(n9858) );
  OAI22_X1 U9526 ( .A1(n10181), .A2(n7901), .B1(n9509), .B2(n10178), .ZN(n7902) );
  AOI21_X1 U9527 ( .B1(n9856), .B2(n9957), .A(n7902), .ZN(n7903) );
  OAI21_X1 U9528 ( .B1(n9858), .B2(n7904), .A(n7903), .ZN(n7905) );
  AOI21_X1 U9529 ( .B1(n9855), .B2(n10164), .A(n7905), .ZN(n7906) );
  OAI21_X1 U9530 ( .B1(n9861), .B2(n9953), .A(n7906), .ZN(P1_U3276) );
  XNOR2_X1 U9531 ( .A(n7908), .B(n7907), .ZN(n7909) );
  XNOR2_X1 U9532 ( .A(n7910), .B(n7909), .ZN(n7919) );
  NOR2_X1 U9533 ( .A1(n9505), .A2(n7911), .ZN(n7912) );
  AOI211_X1 U9534 ( .C1(n9507), .C2(n9770), .A(n7913), .B(n7912), .ZN(n7914)
         );
  OAI21_X1 U9535 ( .B1(n9510), .B2(n7915), .A(n7914), .ZN(n7916) );
  AOI21_X1 U9536 ( .B1(n7917), .B2(n9512), .A(n7916), .ZN(n7918) );
  OAI21_X1 U9537 ( .B1(n7919), .B2(n9514), .A(n7918), .ZN(P1_U3213) );
  INV_X1 U9538 ( .A(n7920), .ZN(n7924) );
  OAI222_X1 U9539 ( .A1(P2_U3152), .A2(n7922), .B1(n9376), .B2(n7924), .C1(
        n7921), .C2(n9382), .ZN(P2_U3333) );
  OAI222_X1 U9540 ( .A1(n9891), .A2(n7925), .B1(n9886), .B2(n7924), .C1(n7923), 
        .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9541 ( .A(n7926), .ZN(n7930) );
  OAI222_X1 U9542 ( .A1(n9886), .A2(n7930), .B1(P1_U3084), .B2(n7928), .C1(
        n7927), .C2(n9891), .ZN(P1_U3327) );
  OAI222_X1 U9543 ( .A1(n7931), .A2(P2_U3152), .B1(n9376), .B2(n7930), .C1(
        n7929), .C2(n9382), .ZN(P2_U3332) );
  INV_X1 U9544 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n7938) );
  AOI22_X1 U9545 ( .A1(n7933), .A2(n10447), .B1(n10444), .B2(n7932), .ZN(n7934) );
  OAI21_X1 U9546 ( .B1(n7935), .B2(n10428), .A(n7934), .ZN(n7936) );
  NOR2_X1 U9547 ( .A1(n7937), .A2(n7936), .ZN(n7940) );
  MUX2_X1 U9548 ( .A(n7938), .B(n7940), .S(n10462), .Z(n7939) );
  INV_X1 U9549 ( .A(n7939), .ZN(P2_U3490) );
  MUX2_X1 U9550 ( .A(n5335), .B(n7940), .S(n10473), .Z(n7941) );
  INV_X1 U9551 ( .A(n7941), .ZN(P2_U3533) );
  INV_X1 U9552 ( .A(n7942), .ZN(n7945) );
  NOR3_X1 U9553 ( .A1(n7943), .A2(n10261), .A3(n8603), .ZN(n7944) );
  AOI21_X1 U9554 ( .B1(n7945), .B2(n10287), .A(n7944), .ZN(n7957) );
  XNOR2_X1 U9555 ( .A(n7993), .B(n8313), .ZN(n7960) );
  NOR2_X1 U9556 ( .A1(n7965), .A2(n8341), .ZN(n7958) );
  XNOR2_X1 U9557 ( .A(n7960), .B(n7958), .ZN(n7956) );
  INV_X1 U9558 ( .A(n9243), .ZN(n8616) );
  OAI21_X1 U9559 ( .B1(n10252), .B2(n10261), .A(n7946), .ZN(n7947) );
  AOI21_X1 U9560 ( .B1(n8610), .B2(n8616), .A(n7947), .ZN(n7948) );
  OAI21_X1 U9561 ( .B1(n7949), .B2(n10292), .A(n7948), .ZN(n7954) );
  AND2_X1 U9562 ( .A1(n7956), .A2(n7950), .ZN(n7951) );
  NOR2_X1 U9563 ( .A1(n7962), .A2(n10246), .ZN(n7953) );
  AOI211_X1 U9564 ( .C1(n10286), .C2(n7993), .A(n7954), .B(n7953), .ZN(n7955)
         );
  OAI21_X1 U9565 ( .B1(n7957), .B2(n7956), .A(n7955), .ZN(P2_U3217) );
  INV_X1 U9566 ( .A(n7958), .ZN(n7959) );
  NAND2_X1 U9567 ( .A1(n7960), .A2(n7959), .ZN(n7961) );
  XNOR2_X1 U9568 ( .A(n9346), .B(n8313), .ZN(n7963) );
  NAND2_X1 U9569 ( .A1(n7964), .A2(n7963), .ZN(n7978) );
  NOR2_X1 U9570 ( .A1(n8603), .A2(n9243), .ZN(n7979) );
  INV_X1 U9571 ( .A(n7979), .ZN(n7971) );
  OR2_X1 U9572 ( .A1(n9243), .A2(n8341), .ZN(n7973) );
  NAND3_X1 U9573 ( .A1(n7972), .A2(n10287), .A3(n7973), .ZN(n7970) );
  OAI22_X1 U9574 ( .A1(n7965), .A2(n9242), .B1(n8440), .B2(n9240), .ZN(n7989)
         );
  NAND2_X1 U9575 ( .A1(n7989), .A2(n10279), .ZN(n7967) );
  OAI211_X1 U9576 ( .C1(n10292), .C2(n7998), .A(n7967), .B(n7966), .ZN(n7968)
         );
  AOI21_X1 U9577 ( .B1(n9346), .B2(n10286), .A(n7968), .ZN(n7969) );
  OAI211_X1 U9578 ( .C1(n7972), .C2(n7971), .A(n7970), .B(n7969), .ZN(P2_U3243) );
  NAND2_X1 U9579 ( .A1(n7976), .A2(n7973), .ZN(n7974) );
  NAND2_X1 U9580 ( .A1(n7974), .A2(n7978), .ZN(n7975) );
  XNOR2_X1 U9581 ( .A(n9340), .B(n8313), .ZN(n8279) );
  NOR2_X1 U9582 ( .A1(n8440), .A2(n8341), .ZN(n8277) );
  XNOR2_X1 U9583 ( .A(n8279), .B(n8277), .ZN(n7977) );
  NOR2_X1 U9584 ( .A1(n7976), .A2(n10246), .ZN(n7980) );
  OAI211_X1 U9585 ( .C1(n7980), .C2(n7979), .A(n4875), .B(n7978), .ZN(n7986)
         );
  INV_X1 U9586 ( .A(n9241), .ZN(n9209) );
  OAI21_X1 U9587 ( .B1(n10252), .B2(n9243), .A(n7981), .ZN(n7982) );
  AOI21_X1 U9588 ( .B1(n8610), .B2(n9209), .A(n7982), .ZN(n7983) );
  OAI21_X1 U9589 ( .B1(n9257), .B2(n10292), .A(n7983), .ZN(n7984) );
  AOI21_X1 U9590 ( .B1(n9340), .B2(n10286), .A(n7984), .ZN(n7985) );
  OAI211_X1 U9591 ( .C1(n8281), .C2(n10246), .A(n7986), .B(n7985), .ZN(
        P2_U3228) );
  XNOR2_X1 U9592 ( .A(n7988), .B(n7987), .ZN(n7990) );
  AOI21_X1 U9593 ( .B1(n7990), .B2(n10371), .A(n7989), .ZN(n9348) );
  OR2_X1 U9594 ( .A1(n7993), .A2(n8617), .ZN(n7994) );
  OAI21_X1 U9595 ( .B1(n7996), .B2(n7995), .A(n8438), .ZN(n7997) );
  INV_X1 U9596 ( .A(n7997), .ZN(n9349) );
  OAI22_X1 U9597 ( .A1(n9259), .A2(n5379), .B1(n7998), .B2(n9256), .ZN(n7999)
         );
  AOI21_X1 U9598 ( .B1(n9346), .B2(n10355), .A(n7999), .ZN(n8004) );
  NAND2_X1 U9599 ( .A1(n8000), .A2(n9346), .ZN(n8001) );
  NAND2_X1 U9600 ( .A1(n8001), .A2(n10447), .ZN(n8002) );
  NOR2_X1 U9601 ( .A1(n9251), .A2(n8002), .ZN(n9345) );
  NAND2_X1 U9602 ( .A1(n9345), .A2(n9179), .ZN(n8003) );
  OAI211_X1 U9603 ( .C1(n9349), .C2(n9233), .A(n8004), .B(n8003), .ZN(n8005)
         );
  INV_X1 U9604 ( .A(n8005), .ZN(n8006) );
  OAI21_X1 U9605 ( .B1(n9348), .B2(n10372), .A(n8006), .ZN(P2_U3281) );
  MUX2_X1 U9606 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n9367), .S(n8007), .Z(n8008) );
  NOR2_X1 U9607 ( .A1(n9921), .A2(n8360), .ZN(n8109) );
  NAND2_X1 U9608 ( .A1(n8351), .A2(n8096), .ZN(n8010) );
  INV_X1 U9609 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8797) );
  OR2_X1 U9610 ( .A1(n5992), .A2(n8797), .ZN(n8009) );
  INV_X1 U9611 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8016) );
  NAND2_X1 U9612 ( .A1(n8011), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8015) );
  INV_X1 U9613 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n8012) );
  OR2_X1 U9614 ( .A1(n8013), .A2(n8012), .ZN(n8014) );
  OAI211_X1 U9615 ( .C1(n8017), .C2(n8016), .A(n8015), .B(n8014), .ZN(n9516)
         );
  NAND2_X1 U9616 ( .A1(n8360), .A2(n9516), .ZN(n8018) );
  NAND2_X1 U9617 ( .A1(n9566), .A2(n8018), .ZN(n8222) );
  INV_X1 U9618 ( .A(n8222), .ZN(n8019) );
  NAND2_X1 U9619 ( .A1(n8019), .A2(n8107), .ZN(n8108) );
  INV_X1 U9620 ( .A(n9663), .ZN(n8020) );
  NOR2_X1 U9621 ( .A1(n9633), .A2(n8020), .ZN(n8022) );
  INV_X1 U9622 ( .A(n9677), .ZN(n8021) );
  NAND2_X1 U9623 ( .A1(n9811), .A2(n8021), .ZN(n8407) );
  INV_X1 U9624 ( .A(n9518), .ZN(n9643) );
  NAND2_X1 U9625 ( .A1(n9799), .A2(n9643), .ZN(n8412) );
  NAND2_X1 U9626 ( .A1(n9633), .A2(n8020), .ZN(n8410) );
  OAI21_X1 U9627 ( .B1(n8022), .B2(n8407), .A(n8150), .ZN(n8024) );
  INV_X1 U9628 ( .A(n8410), .ZN(n8092) );
  OR2_X1 U9629 ( .A1(n9811), .A2(n8021), .ZN(n9636) );
  INV_X1 U9630 ( .A(n8022), .ZN(n8091) );
  OAI211_X1 U9631 ( .C1(n8092), .C2(n9636), .A(n8211), .B(n8091), .ZN(n8023)
         );
  MUX2_X1 U9632 ( .A(n8024), .B(n8023), .S(n8107), .Z(n8094) );
  INV_X1 U9633 ( .A(n9662), .ZN(n9689) );
  NAND2_X1 U9634 ( .A1(n9816), .A2(n9689), .ZN(n8113) );
  INV_X1 U9635 ( .A(n9707), .ZN(n8025) );
  NAND2_X1 U9636 ( .A1(n9823), .A2(n8025), .ZN(n9674) );
  NAND2_X1 U9637 ( .A1(n8113), .A2(n9674), .ZN(n8086) );
  INV_X1 U9638 ( .A(n9519), .ZN(n9718) );
  AND2_X1 U9639 ( .A1(n9826), .A2(n9718), .ZN(n8080) );
  AND2_X1 U9640 ( .A1(n8178), .A2(n8080), .ZN(n8026) );
  NOR2_X1 U9641 ( .A1(n8086), .A2(n8026), .ZN(n8204) );
  INV_X1 U9642 ( .A(n9727), .ZN(n9487) );
  NAND2_X1 U9643 ( .A1(n9833), .A2(n9487), .ZN(n8399) );
  INV_X1 U9644 ( .A(n9752), .ZN(n9717) );
  NAND2_X1 U9645 ( .A1(n9838), .A2(n9717), .ZN(n8398) );
  AND2_X1 U9646 ( .A1(n8399), .A2(n8398), .ZN(n8180) );
  OR2_X1 U9647 ( .A1(n9838), .A2(n9717), .ZN(n8116) );
  INV_X1 U9648 ( .A(n9771), .ZN(n8027) );
  OR2_X1 U9649 ( .A1(n9845), .A2(n8027), .ZN(n8396) );
  NAND2_X1 U9650 ( .A1(n8116), .A2(n8396), .ZN(n8179) );
  NAND2_X1 U9651 ( .A1(n9845), .A2(n8027), .ZN(n8075) );
  NAND2_X1 U9652 ( .A1(n8398), .A2(n8075), .ZN(n8182) );
  INV_X1 U9653 ( .A(n8107), .ZN(n8090) );
  MUX2_X1 U9654 ( .A(n8179), .B(n8182), .S(n8090), .Z(n8028) );
  INV_X1 U9655 ( .A(n8028), .ZN(n8079) );
  OR2_X1 U9656 ( .A1(n9850), .A2(n8029), .ZN(n8195) );
  NAND2_X1 U9657 ( .A1(n9850), .A2(n8029), .ZN(n9750) );
  MUX2_X1 U9658 ( .A(n9751), .B(n9850), .S(n8090), .Z(n8077) );
  INV_X1 U9659 ( .A(n8036), .ZN(n8030) );
  NAND2_X1 U9660 ( .A1(n8037), .A2(n8030), .ZN(n8035) );
  AND2_X1 U9661 ( .A1(n8032), .A2(n8031), .ZN(n8034) );
  INV_X1 U9662 ( .A(n8038), .ZN(n8033) );
  AOI21_X1 U9663 ( .B1(n8035), .B2(n8034), .A(n8033), .ZN(n8042) );
  OR2_X1 U9664 ( .A1(n8037), .A2(n8036), .ZN(n8040) );
  AND2_X1 U9665 ( .A1(n8038), .A2(n8122), .ZN(n8164) );
  AOI21_X1 U9666 ( .B1(n8040), .B2(n8164), .A(n8039), .ZN(n8041) );
  MUX2_X1 U9667 ( .A(n8042), .B(n8041), .S(n8090), .Z(n8047) );
  NAND2_X1 U9668 ( .A1(n8129), .A2(n8184), .ZN(n8043) );
  AND2_X1 U9669 ( .A1(n8048), .A2(n8128), .ZN(n8155) );
  OAI21_X1 U9670 ( .B1(n8047), .B2(n8043), .A(n8155), .ZN(n8044) );
  NAND3_X1 U9671 ( .A1(n8044), .A2(n8152), .A3(n8056), .ZN(n8051) );
  NAND2_X1 U9672 ( .A1(n8128), .A2(n8045), .ZN(n8046) );
  AOI21_X1 U9673 ( .B1(n8047), .B2(n8184), .A(n8046), .ZN(n8049) );
  NAND2_X1 U9674 ( .A1(n8152), .A2(n8129), .ZN(n8186) );
  OAI211_X1 U9675 ( .C1(n8049), .C2(n8186), .A(n8154), .B(n8048), .ZN(n8050)
         );
  MUX2_X1 U9676 ( .A(n8051), .B(n8050), .S(n8107), .Z(n8061) );
  AND2_X1 U9677 ( .A1(n8053), .A2(n8052), .ZN(n9966) );
  NAND2_X1 U9678 ( .A1(n8064), .A2(n8054), .ZN(n8191) );
  NAND2_X1 U9679 ( .A1(n8055), .A2(n8154), .ZN(n8188) );
  NAND2_X1 U9680 ( .A1(n8188), .A2(n8107), .ZN(n8059) );
  NAND2_X1 U9681 ( .A1(n8151), .A2(n8090), .ZN(n8062) );
  INV_X1 U9682 ( .A(n8056), .ZN(n8057) );
  OAI211_X1 U9683 ( .C1(n8057), .C2(n8153), .A(n8187), .B(n8154), .ZN(n8058)
         );
  OAI22_X1 U9684 ( .A1(n8191), .A2(n8059), .B1(n8062), .B2(n8058), .ZN(n8060)
         );
  OAI21_X1 U9685 ( .B1(n8061), .B2(n9966), .A(n8060), .ZN(n8068) );
  INV_X1 U9686 ( .A(n8062), .ZN(n8063) );
  NAND2_X1 U9687 ( .A1(n8063), .A2(n8191), .ZN(n8067) );
  NAND2_X1 U9688 ( .A1(n8151), .A2(n8187), .ZN(n8065) );
  NAND3_X1 U9689 ( .A1(n8065), .A2(n8064), .A3(n8107), .ZN(n8066) );
  NAND4_X1 U9690 ( .A1(n8068), .A2(n8136), .A3(n8067), .A4(n8066), .ZN(n8074)
         );
  NAND2_X1 U9691 ( .A1(n9850), .A2(n9751), .ZN(n8366) );
  NAND2_X1 U9692 ( .A1(n8077), .A2(n8366), .ZN(n8073) );
  INV_X1 U9693 ( .A(n8393), .ZN(n8070) );
  INV_X1 U9694 ( .A(n8194), .ZN(n8069) );
  MUX2_X1 U9695 ( .A(n8070), .B(n8069), .S(n8107), .Z(n8071) );
  INV_X1 U9696 ( .A(n8071), .ZN(n8072) );
  NAND3_X1 U9697 ( .A1(n8074), .A2(n8073), .A3(n8072), .ZN(n8076) );
  OAI211_X1 U9698 ( .C1(n9769), .C2(n8077), .A(n8076), .B(n9749), .ZN(n8078)
         );
  NAND2_X1 U9699 ( .A1(n8079), .A2(n8078), .ZN(n8082) );
  OR2_X1 U9700 ( .A1(n9833), .A2(n9487), .ZN(n8115) );
  NAND2_X1 U9701 ( .A1(n9683), .A2(n8115), .ZN(n8181) );
  AOI21_X1 U9702 ( .B1(n8180), .B2(n8082), .A(n8181), .ZN(n8085) );
  AND2_X1 U9703 ( .A1(n8115), .A2(n8116), .ZN(n8083) );
  INV_X1 U9704 ( .A(n8080), .ZN(n8114) );
  NAND2_X1 U9705 ( .A1(n8114), .A2(n8399), .ZN(n8081) );
  AOI21_X1 U9706 ( .B1(n8083), .B2(n8082), .A(n8081), .ZN(n8084) );
  MUX2_X1 U9707 ( .A(n8085), .B(n8084), .S(n8090), .Z(n8088) );
  NOR2_X1 U9708 ( .A1(n9816), .A2(n9689), .ZN(n8089) );
  NAND2_X1 U9709 ( .A1(n8178), .A2(n9683), .ZN(n8087) );
  INV_X1 U9710 ( .A(n8086), .ZN(n8404) );
  INV_X1 U9711 ( .A(n8089), .ZN(n8405) );
  NAND2_X1 U9712 ( .A1(n8091), .A2(n9636), .ZN(n8408) );
  INV_X1 U9713 ( .A(n8407), .ZN(n8207) );
  XNOR2_X1 U9714 ( .A(n9796), .B(n9627), .ZN(n9605) );
  INV_X1 U9715 ( .A(n9627), .ZN(n9598) );
  NAND2_X1 U9716 ( .A1(n9796), .A2(n9598), .ZN(n8413) );
  INV_X1 U9717 ( .A(n9576), .ZN(n9614) );
  NAND2_X1 U9718 ( .A1(n9789), .A2(n9614), .ZN(n8112) );
  NOR2_X1 U9719 ( .A1(n9789), .A2(n9614), .ZN(n8218) );
  INV_X1 U9720 ( .A(n8218), .ZN(n8414) );
  INV_X1 U9721 ( .A(n9517), .ZN(n9597) );
  NAND3_X1 U9722 ( .A1(n8103), .A2(n8414), .A3(n8415), .ZN(n8101) );
  NAND2_X1 U9723 ( .A1(n9783), .A2(n9597), .ZN(n8416) );
  NAND2_X1 U9724 ( .A1(n8471), .A2(n8096), .ZN(n8098) );
  OR2_X1 U9725 ( .A1(n5992), .A2(n8472), .ZN(n8097) );
  INV_X1 U9726 ( .A(n9577), .ZN(n8099) );
  INV_X1 U9727 ( .A(n8418), .ZN(n8100) );
  AOI21_X1 U9728 ( .B1(n8101), .B2(n8416), .A(n8100), .ZN(n8102) );
  NOR2_X1 U9729 ( .A1(n8102), .A2(n8259), .ZN(n8106) );
  NOR2_X1 U9730 ( .A1(n9796), .A2(n9598), .ZN(n8210) );
  NAND2_X1 U9731 ( .A1(n8416), .A2(n8112), .ZN(n8149) );
  AOI21_X1 U9732 ( .B1(n8104), .B2(n8418), .A(n8219), .ZN(n8105) );
  NAND2_X1 U9733 ( .A1(n9981), .A2(n9516), .ZN(n8110) );
  AOI21_X1 U9734 ( .B1(n8360), .B2(n8110), .A(n9921), .ZN(n8146) );
  NAND2_X1 U9735 ( .A1(n9921), .A2(n8360), .ZN(n8262) );
  INV_X1 U9736 ( .A(n8109), .ZN(n8111) );
  NAND2_X1 U9737 ( .A1(n8111), .A2(n8110), .ZN(n8263) );
  NAND2_X1 U9738 ( .A1(n8415), .A2(n8416), .ZN(n9573) );
  NAND2_X1 U9739 ( .A1(n8414), .A2(n8112), .ZN(n9595) );
  NAND2_X1 U9740 ( .A1(n9636), .A2(n8407), .ZN(n9660) );
  NAND2_X1 U9741 ( .A1(n8405), .A2(n8113), .ZN(n9676) );
  NAND2_X1 U9742 ( .A1(n8178), .A2(n9674), .ZN(n9687) );
  NAND2_X1 U9743 ( .A1(n9683), .A2(n8114), .ZN(n9697) );
  NAND2_X1 U9744 ( .A1(n8115), .A2(n8399), .ZN(n9714) );
  NAND2_X1 U9745 ( .A1(n8116), .A2(n8398), .ZN(n8397) );
  INV_X1 U9746 ( .A(n8117), .ZN(n8121) );
  NOR4_X1 U9747 ( .A1(n8121), .A2(n8120), .A3(n8119), .A4(n8118), .ZN(n8124)
         );
  NAND4_X1 U9748 ( .A1(n8124), .A2(n8123), .A3(n8170), .A4(n8122), .ZN(n8127)
         );
  NOR4_X1 U9749 ( .A1(n8127), .A2(n8251), .A3(n8126), .A4(n8125), .ZN(n8131)
         );
  INV_X1 U9750 ( .A(n9966), .ZN(n9960) );
  NAND4_X1 U9751 ( .A1(n8131), .A2(n9960), .A3(n8130), .A4(n10166), .ZN(n8132)
         );
  NOR4_X1 U9752 ( .A1(n8134), .A2(n9942), .A3(n8133), .A4(n8132), .ZN(n8135)
         );
  NAND4_X1 U9753 ( .A1(n9749), .A2(n8136), .A3(n9769), .A4(n8135), .ZN(n8137)
         );
  OR4_X1 U9754 ( .A1(n9697), .A2(n9714), .A3(n8397), .A4(n8137), .ZN(n8138) );
  NOR4_X1 U9755 ( .A1(n9660), .A2(n9676), .A3(n9687), .A4(n8138), .ZN(n8139)
         );
  OR2_X1 U9756 ( .A1(n9633), .A2(n9663), .ZN(n8381) );
  NAND2_X1 U9757 ( .A1(n9633), .A2(n9663), .ZN(n8380) );
  NAND2_X1 U9758 ( .A1(n8381), .A2(n8380), .ZN(n9638) );
  NAND3_X1 U9759 ( .A1(n9626), .A2(n8139), .A3(n9638), .ZN(n8140) );
  NOR4_X1 U9760 ( .A1(n9573), .A2(n9595), .A3(n4752), .A4(n8140), .ZN(n8142)
         );
  INV_X1 U9761 ( .A(n9516), .ZN(n8141) );
  NAND2_X1 U9762 ( .A1(n9566), .A2(n8141), .ZN(n8257) );
  NAND4_X1 U9763 ( .A1(n8262), .A2(n8418), .A3(n8142), .A4(n8257), .ZN(n8143)
         );
  OAI21_X1 U9764 ( .B1(n8263), .B2(n8143), .A(n8236), .ZN(n8145) );
  INV_X1 U9765 ( .A(n8145), .ZN(n8228) );
  INV_X1 U9766 ( .A(n8146), .ZN(n8226) );
  INV_X1 U9767 ( .A(n8413), .ZN(n8147) );
  AND2_X1 U9768 ( .A1(n8414), .A2(n8147), .ZN(n8148) );
  OR2_X1 U9769 ( .A1(n8149), .A2(n8148), .ZN(n8215) );
  INV_X1 U9770 ( .A(n8150), .ZN(n8213) );
  AND2_X1 U9771 ( .A1(n8393), .A2(n8151), .ZN(n8193) );
  INV_X1 U9772 ( .A(n8152), .ZN(n8156) );
  OAI211_X1 U9773 ( .C1(n8156), .C2(n8155), .A(n8154), .B(n8153), .ZN(n8157)
         );
  INV_X1 U9774 ( .A(n8157), .ZN(n8158) );
  AND2_X1 U9775 ( .A1(n8187), .A2(n8158), .ZN(n8183) );
  NAND4_X1 U9776 ( .A1(n9750), .A2(n8193), .A3(n8159), .A4(n8183), .ZN(n8160)
         );
  NOR2_X1 U9777 ( .A1(n8182), .A2(n8160), .ZN(n8161) );
  NAND4_X1 U9778 ( .A1(n8204), .A2(n8161), .A3(n8399), .A4(n8407), .ZN(n8162)
         );
  OR2_X1 U9779 ( .A1(n8213), .A2(n8162), .ZN(n8163) );
  OR2_X1 U9780 ( .A1(n8215), .A2(n8163), .ZN(n8248) );
  INV_X1 U9781 ( .A(n8164), .ZN(n8173) );
  NOR2_X1 U9782 ( .A1(n8173), .A2(n8165), .ZN(n8250) );
  NAND2_X1 U9783 ( .A1(n8250), .A2(n8171), .ZN(n8256) );
  INV_X1 U9784 ( .A(n8166), .ZN(n8168) );
  INV_X1 U9785 ( .A(n8246), .ZN(n8167) );
  NOR3_X1 U9786 ( .A1(n8256), .A2(n8168), .A3(n8167), .ZN(n8177) );
  INV_X1 U9787 ( .A(n8169), .ZN(n8172) );
  NAND3_X1 U9788 ( .A1(n8172), .A2(n8171), .A3(n8170), .ZN(n8174) );
  AOI21_X1 U9789 ( .B1(n8175), .B2(n8174), .A(n8173), .ZN(n8176) );
  NOR3_X1 U9790 ( .A1(n8248), .A2(n8177), .A3(n8176), .ZN(n8224) );
  INV_X1 U9791 ( .A(n8178), .ZN(n8206) );
  INV_X1 U9792 ( .A(n8179), .ZN(n8203) );
  INV_X1 U9793 ( .A(n8180), .ZN(n8202) );
  INV_X1 U9794 ( .A(n8181), .ZN(n8201) );
  INV_X1 U9795 ( .A(n8182), .ZN(n8199) );
  INV_X1 U9796 ( .A(n8183), .ZN(n8190) );
  INV_X1 U9797 ( .A(n8184), .ZN(n8185) );
  NOR2_X1 U9798 ( .A1(n8186), .A2(n8185), .ZN(n8189) );
  OAI22_X1 U9799 ( .A1(n8190), .A2(n8189), .B1(n4745), .B2(n8188), .ZN(n8192)
         );
  NOR2_X1 U9800 ( .A1(n8192), .A2(n8191), .ZN(n8197) );
  INV_X1 U9801 ( .A(n8193), .ZN(n8196) );
  OAI211_X1 U9802 ( .C1(n8197), .C2(n8196), .A(n8195), .B(n8194), .ZN(n8198)
         );
  NAND4_X1 U9803 ( .A1(n8399), .A2(n8199), .A3(n9750), .A4(n8198), .ZN(n8200)
         );
  OAI211_X1 U9804 ( .C1(n8203), .C2(n8202), .A(n8201), .B(n8200), .ZN(n8205)
         );
  OAI21_X1 U9805 ( .B1(n8206), .B2(n8205), .A(n8204), .ZN(n8208) );
  AOI21_X1 U9806 ( .B1(n8208), .B2(n8405), .A(n8207), .ZN(n8209) );
  NOR2_X1 U9807 ( .A1(n8209), .A2(n8408), .ZN(n8214) );
  INV_X1 U9808 ( .A(n8210), .ZN(n8212) );
  OAI211_X1 U9809 ( .C1(n8214), .C2(n8213), .A(n8212), .B(n8211), .ZN(n8217)
         );
  INV_X1 U9810 ( .A(n8215), .ZN(n8216) );
  OAI21_X1 U9811 ( .B1(n8218), .B2(n8217), .A(n8216), .ZN(n8221) );
  INV_X1 U9812 ( .A(n8219), .ZN(n8220) );
  NAND3_X1 U9813 ( .A1(n8221), .A2(n8220), .A3(n8415), .ZN(n8235) );
  INV_X1 U9814 ( .A(n8259), .ZN(n8223) );
  OAI211_X1 U9815 ( .C1(n8224), .C2(n8235), .A(n8223), .B(n8222), .ZN(n8225)
         );
  INV_X1 U9816 ( .A(n8262), .ZN(n8231) );
  AOI211_X1 U9817 ( .C1(n8226), .C2(n8225), .A(n8236), .B(n8231), .ZN(n8227)
         );
  NOR2_X1 U9818 ( .A1(n8228), .A2(n8227), .ZN(n8230) );
  NOR3_X1 U9819 ( .A1(n8231), .A2(n8273), .A3(n8236), .ZN(n8232) );
  NAND2_X1 U9820 ( .A1(n8233), .A2(n8232), .ZN(n8234) );
  INV_X1 U9821 ( .A(n8235), .ZN(n8261) );
  AOI21_X1 U9822 ( .B1(n9531), .B2(n10196), .A(n8236), .ZN(n8241) );
  INV_X1 U9823 ( .A(n8237), .ZN(n8239) );
  AOI211_X1 U9824 ( .C1(n8241), .C2(n8240), .A(n8239), .B(n8238), .ZN(n8245)
         );
  INV_X1 U9825 ( .A(n8242), .ZN(n8244) );
  OAI21_X1 U9826 ( .B1(n8245), .B2(n8244), .A(n8243), .ZN(n8247) );
  NAND2_X1 U9827 ( .A1(n8247), .A2(n8246), .ZN(n8255) );
  INV_X1 U9828 ( .A(n8248), .ZN(n8254) );
  INV_X1 U9829 ( .A(n8249), .ZN(n8252) );
  OAI21_X1 U9830 ( .B1(n8252), .B2(n8251), .A(n8250), .ZN(n8253) );
  OAI211_X1 U9831 ( .C1(n8256), .C2(n8255), .A(n8254), .B(n8253), .ZN(n8260)
         );
  INV_X1 U9832 ( .A(n8257), .ZN(n8258) );
  AOI211_X1 U9833 ( .C1(n8261), .C2(n8260), .A(n8259), .B(n8258), .ZN(n8264)
         );
  OAI21_X1 U9834 ( .B1(n8264), .B2(n8263), .A(n8262), .ZN(n8265) );
  XNOR2_X1 U9835 ( .A(n8265), .B(n4695), .ZN(n8267) );
  INV_X1 U9836 ( .A(n8270), .ZN(n9879) );
  NOR4_X1 U9837 ( .A1(n8272), .A2(n9879), .A3(n8271), .A4(n4498), .ZN(n8275)
         );
  OAI21_X1 U9838 ( .B1(n8273), .B2(n8276), .A(P1_B_REG_SCAN_IN), .ZN(n8274) );
  XNOR2_X1 U9839 ( .A(n9300), .B(n8313), .ZN(n8538) );
  NOR2_X1 U9840 ( .A1(n8540), .A2(n8341), .ZN(n8320) );
  INV_X1 U9841 ( .A(n8320), .ZN(n8542) );
  INV_X1 U9842 ( .A(n8277), .ZN(n8278) );
  NAND2_X1 U9843 ( .A1(n8279), .A2(n8278), .ZN(n8280) );
  XNOR2_X1 U9844 ( .A(n9335), .B(n8343), .ZN(n8282) );
  NOR2_X1 U9845 ( .A1(n9241), .A2(n8341), .ZN(n8283) );
  NAND2_X1 U9846 ( .A1(n8282), .A2(n8283), .ZN(n8286) );
  INV_X1 U9847 ( .A(n8282), .ZN(n8590) );
  INV_X1 U9848 ( .A(n8283), .ZN(n8284) );
  NAND2_X1 U9849 ( .A1(n8590), .A2(n8284), .ZN(n8285) );
  NAND2_X1 U9850 ( .A1(n8286), .A2(n8285), .ZN(n8527) );
  XNOR2_X1 U9851 ( .A(n9329), .B(n8343), .ZN(n8287) );
  NOR2_X1 U9852 ( .A1(n8531), .A2(n8341), .ZN(n8288) );
  NAND2_X1 U9853 ( .A1(n8287), .A2(n8288), .ZN(n8292) );
  INV_X1 U9854 ( .A(n8287), .ZN(n8496) );
  INV_X1 U9855 ( .A(n8288), .ZN(n8289) );
  NAND2_X1 U9856 ( .A1(n8496), .A2(n8289), .ZN(n8290) );
  AND2_X1 U9857 ( .A1(n8292), .A2(n8290), .ZN(n8587) );
  NAND2_X1 U9858 ( .A1(n8291), .A2(n8587), .ZN(n8494) );
  XNOR2_X1 U9859 ( .A(n9326), .B(n8343), .ZN(n8294) );
  NAND2_X1 U9860 ( .A1(n9210), .A2(n8314), .ZN(n8295) );
  XNOR2_X1 U9861 ( .A(n8294), .B(n8295), .ZN(n8497) );
  AND2_X1 U9862 ( .A1(n8497), .A2(n8292), .ZN(n8293) );
  INV_X1 U9863 ( .A(n8294), .ZN(n8296) );
  NAND2_X1 U9864 ( .A1(n8296), .A2(n8295), .ZN(n8297) );
  XNOR2_X1 U9865 ( .A(n9321), .B(n8343), .ZN(n8298) );
  NOR2_X1 U9866 ( .A1(n8615), .A2(n8341), .ZN(n8299) );
  NAND2_X1 U9867 ( .A1(n8298), .A2(n8299), .ZN(n8303) );
  INV_X1 U9868 ( .A(n8298), .ZN(n8513) );
  INV_X1 U9869 ( .A(n8299), .ZN(n8300) );
  NAND2_X1 U9870 ( .A1(n8513), .A2(n8300), .ZN(n8301) );
  NAND2_X1 U9871 ( .A1(n8303), .A2(n8301), .ZN(n8549) );
  XNOR2_X1 U9872 ( .A(n9315), .B(n8313), .ZN(n8305) );
  NOR2_X1 U9873 ( .A1(n8558), .A2(n8341), .ZN(n8306) );
  XNOR2_X1 U9874 ( .A(n8305), .B(n8306), .ZN(n8511) );
  NAND2_X1 U9875 ( .A1(n8304), .A2(n8511), .ZN(n8564) );
  XNOR2_X1 U9876 ( .A(n9310), .B(n8343), .ZN(n8309) );
  NOR2_X1 U9877 ( .A1(n8567), .A2(n8341), .ZN(n8310) );
  INV_X1 U9878 ( .A(n8305), .ZN(n8307) );
  AND2_X1 U9879 ( .A1(n8307), .A2(n8306), .ZN(n8562) );
  AOI21_X1 U9880 ( .B1(n8309), .B2(n8310), .A(n8562), .ZN(n8308) );
  NAND2_X1 U9881 ( .A1(n8564), .A2(n8308), .ZN(n8312) );
  INV_X1 U9882 ( .A(n8309), .ZN(n8565) );
  INV_X1 U9883 ( .A(n8310), .ZN(n8570) );
  NAND2_X1 U9884 ( .A1(n8565), .A2(n8570), .ZN(n8311) );
  XNOR2_X1 U9885 ( .A(n9128), .B(n8313), .ZN(n8317) );
  NAND2_X1 U9886 ( .A1(n9113), .A2(n8314), .ZN(n8487) );
  AOI21_X1 U9887 ( .B1(n8538), .B2(n8540), .A(n8487), .ZN(n8315) );
  NAND2_X1 U9888 ( .A1(n8486), .A2(n8315), .ZN(n8322) );
  INV_X1 U9889 ( .A(n8538), .ZN(n8319) );
  INV_X1 U9890 ( .A(n8316), .ZN(n8318) );
  OAI21_X1 U9891 ( .B1(n8320), .B2(n8319), .A(n8536), .ZN(n8321) );
  XNOR2_X1 U9892 ( .A(n9296), .B(n8343), .ZN(n8323) );
  NOR2_X1 U9893 ( .A1(n8604), .A2(n8341), .ZN(n8324) );
  NAND2_X1 U9894 ( .A1(n8323), .A2(n8324), .ZN(n8327) );
  INV_X1 U9895 ( .A(n8323), .ZN(n8605) );
  INV_X1 U9896 ( .A(n8324), .ZN(n8325) );
  NAND2_X1 U9897 ( .A1(n8605), .A2(n8325), .ZN(n8326) );
  AND2_X1 U9898 ( .A1(n8327), .A2(n8326), .ZN(n8520) );
  XNOR2_X1 U9899 ( .A(n9291), .B(n8343), .ZN(n8328) );
  NOR2_X1 U9900 ( .A1(n8522), .A2(n8341), .ZN(n8329) );
  NAND2_X1 U9901 ( .A1(n8328), .A2(n8329), .ZN(n8332) );
  INV_X1 U9902 ( .A(n8328), .ZN(n8478) );
  INV_X1 U9903 ( .A(n8329), .ZN(n8330) );
  NAND2_X1 U9904 ( .A1(n8478), .A2(n8330), .ZN(n8331) );
  AND2_X1 U9905 ( .A1(n8332), .A2(n8331), .ZN(n8600) );
  NAND2_X1 U9906 ( .A1(n8475), .A2(n8332), .ZN(n8339) );
  XNOR2_X1 U9907 ( .A(n9285), .B(n8343), .ZN(n8334) );
  NOR2_X1 U9908 ( .A1(n8333), .A2(n8341), .ZN(n8335) );
  NAND2_X1 U9909 ( .A1(n8334), .A2(n8335), .ZN(n8340) );
  INV_X1 U9910 ( .A(n8334), .ZN(n8337) );
  INV_X1 U9911 ( .A(n8335), .ZN(n8336) );
  NAND2_X1 U9912 ( .A1(n8337), .A2(n8336), .ZN(n8338) );
  AND2_X1 U9913 ( .A1(n8340), .A2(n8338), .ZN(n8476) );
  NAND2_X1 U9914 ( .A1(n8339), .A2(n8476), .ZN(n8479) );
  NAND2_X1 U9915 ( .A1(n8479), .A2(n8340), .ZN(n8346) );
  NOR2_X1 U9916 ( .A1(n8342), .A2(n8341), .ZN(n8344) );
  XNOR2_X1 U9917 ( .A(n8344), .B(n8343), .ZN(n8345) );
  OAI22_X1 U9918 ( .A1(n9047), .A2(n10292), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8348), .ZN(n8349) );
  AOI21_X1 U9919 ( .B1(n10257), .B2(n9083), .A(n8349), .ZN(n8350) );
  INV_X1 U9920 ( .A(n8351), .ZN(n8435) );
  OAI222_X1 U9921 ( .A1(n8353), .A2(P2_U3152), .B1(n9376), .B2(n8435), .C1(
        n8352), .C2(n9382), .ZN(P2_U3328) );
  OAI222_X1 U9922 ( .A1(n8355), .A2(P2_U3152), .B1(n9376), .B2(n8354), .C1(
        n8813), .C2(n9382), .ZN(P2_U3338) );
  INV_X1 U9923 ( .A(n9796), .ZN(n8356) );
  INV_X1 U9924 ( .A(n9811), .ZN(n9659) );
  INV_X1 U9925 ( .A(n9826), .ZN(n9703) );
  INV_X1 U9926 ( .A(n9850), .ZN(n9766) );
  AND2_X2 U9927 ( .A1(n9760), .A2(n9766), .ZN(n9761) );
  OR2_X2 U9928 ( .A1(n9699), .A2(n9823), .ZN(n9690) );
  NOR2_X1 U9929 ( .A1(n9816), .A2(n9690), .ZN(n9669) );
  NAND2_X1 U9930 ( .A1(n9659), .A2(n9669), .ZN(n9653) );
  OR2_X2 U9931 ( .A1(n9633), .A2(n9653), .ZN(n9634) );
  INV_X1 U9932 ( .A(n9581), .ZN(n8357) );
  AND2_X2 U9933 ( .A1(n8392), .A2(n8357), .ZN(n9565) );
  NAND2_X1 U9934 ( .A1(n9981), .A2(n9565), .ZN(n8358) );
  XNOR2_X1 U9935 ( .A(n9921), .B(n8358), .ZN(n9923) );
  NAND2_X1 U9936 ( .A1(n9923), .A2(n10163), .ZN(n8362) );
  AOI21_X1 U9937 ( .B1(n8359), .B2(P1_B_REG_SCAN_IN), .A(n10167), .ZN(n8420)
         );
  NAND2_X1 U9938 ( .A1(n8420), .A2(n8360), .ZN(n9980) );
  NOR2_X1 U9939 ( .A1(n9953), .A2(n9980), .ZN(n9567) );
  AOI21_X1 U9940 ( .B1(n9953), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9567), .ZN(
        n8361) );
  OAI211_X1 U9941 ( .C1(n9921), .C2(n10177), .A(n8362), .B(n8361), .ZN(
        P1_U3261) );
  NOR2_X1 U9942 ( .A1(n9856), .A2(n9770), .ZN(n8364) );
  NAND2_X1 U9943 ( .A1(n9856), .A2(n9770), .ZN(n8363) );
  NAND2_X1 U9944 ( .A1(n8367), .A2(n8366), .ZN(n9740) );
  AND2_X1 U9945 ( .A1(n9845), .A2(n9771), .ZN(n8368) );
  NAND2_X1 U9946 ( .A1(n9833), .A2(n9727), .ZN(n8369) );
  NAND2_X1 U9947 ( .A1(n8370), .A2(n8369), .ZN(n9698) );
  OR2_X1 U9948 ( .A1(n9826), .A2(n9519), .ZN(n8371) );
  NAND2_X1 U9949 ( .A1(n9698), .A2(n8371), .ZN(n8373) );
  NAND2_X1 U9950 ( .A1(n9826), .A2(n9519), .ZN(n8372) );
  NAND2_X1 U9951 ( .A1(n8373), .A2(n8372), .ZN(n9682) );
  NAND2_X1 U9952 ( .A1(n9682), .A2(n9687), .ZN(n8375) );
  NAND2_X1 U9953 ( .A1(n9823), .A2(n9707), .ZN(n8374) );
  NAND2_X1 U9954 ( .A1(n8375), .A2(n8374), .ZN(n9668) );
  INV_X1 U9955 ( .A(n9668), .ZN(n8376) );
  OR2_X1 U9956 ( .A1(n9816), .A2(n9662), .ZN(n8377) );
  NAND2_X1 U9957 ( .A1(n9811), .A2(n9677), .ZN(n8378) );
  INV_X1 U9958 ( .A(n8380), .ZN(n8382) );
  OR2_X1 U9959 ( .A1(n9799), .A2(n9518), .ZN(n8383) );
  NAND2_X1 U9960 ( .A1(n9796), .A2(n9627), .ZN(n8384) );
  NAND2_X1 U9961 ( .A1(n8385), .A2(n8384), .ZN(n9589) );
  INV_X1 U9962 ( .A(n9589), .ZN(n8386) );
  OR2_X1 U9963 ( .A1(n9789), .A2(n9576), .ZN(n8387) );
  INV_X1 U9964 ( .A(n9573), .ZN(n9570) );
  XNOR2_X1 U9965 ( .A(n8388), .B(n8418), .ZN(n9782) );
  AOI21_X1 U9966 ( .B1(n9778), .B2(n9581), .A(n9565), .ZN(n9779) );
  INV_X1 U9967 ( .A(n8389), .ZN(n8390) );
  AOI22_X1 U9968 ( .A1(n9953), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8390), .B2(
        n9763), .ZN(n8391) );
  OAI21_X1 U9969 ( .B1(n8392), .B2(n10177), .A(n8391), .ZN(n8422) );
  NAND2_X1 U9970 ( .A1(n8394), .A2(n8393), .ZN(n9768) );
  AND2_X1 U9971 ( .A1(n9749), .A2(n9750), .ZN(n8395) );
  INV_X1 U9972 ( .A(n9714), .ZN(n8401) );
  INV_X1 U9973 ( .A(n8399), .ZN(n8400) );
  AOI21_X1 U9974 ( .B1(n9715), .B2(n8401), .A(n8400), .ZN(n9706) );
  INV_X1 U9975 ( .A(n9697), .ZN(n9705) );
  INV_X1 U9976 ( .A(n9683), .ZN(n8402) );
  NOR2_X1 U9977 ( .A1(n9687), .A2(n8402), .ZN(n8403) );
  NAND2_X1 U9978 ( .A1(n9704), .A2(n8403), .ZN(n9684) );
  NAND2_X1 U9979 ( .A1(n9684), .A2(n8404), .ZN(n8406) );
  NAND2_X1 U9980 ( .A1(n8406), .A2(n8405), .ZN(n9661) );
  NAND2_X1 U9981 ( .A1(n9661), .A2(n8407), .ZN(n9637) );
  INV_X1 U9982 ( .A(n8408), .ZN(n8409) );
  NAND2_X1 U9983 ( .A1(n9637), .A2(n8409), .ZN(n8411) );
  NAND2_X1 U9984 ( .A1(n8411), .A2(n8410), .ZN(n9625) );
  INV_X1 U9985 ( .A(n8415), .ZN(n8417) );
  OAI21_X1 U9986 ( .B1(n9574), .B2(n8417), .A(n8416), .ZN(n8419) );
  NOR2_X1 U9987 ( .A1(n9780), .A2(n9953), .ZN(n8421) );
  OAI21_X1 U9988 ( .B1(n9782), .B2(n9777), .A(n8423), .ZN(P1_U3355) );
  OAI22_X1 U9989 ( .A1(n8424), .A2(n8603), .B1(n10246), .B2(n10403), .ZN(n8426) );
  NAND2_X1 U9990 ( .A1(n8426), .A2(n8425), .ZN(n8433) );
  AND2_X1 U9991 ( .A1(n8428), .A2(n8427), .ZN(n8429) );
  NAND2_X1 U9992 ( .A1(n8430), .A2(n8429), .ZN(n8575) );
  AOI22_X1 U9993 ( .A1(n10286), .A2(n8431), .B1(n8575), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n8432) );
  OAI211_X1 U9994 ( .C1(n8580), .C2(n10260), .A(n8433), .B(n8432), .ZN(
        P2_U3234) );
  OAI222_X1 U9995 ( .A1(n9891), .A2(n8797), .B1(n9886), .B2(n8435), .C1(
        P1_U3084), .C2(n8434), .ZN(P1_U3323) );
  INV_X1 U9996 ( .A(n9346), .ZN(n8436) );
  NAND2_X1 U9997 ( .A1(n8436), .A2(n9243), .ZN(n8437) );
  NAND2_X1 U9998 ( .A1(n8438), .A2(n8437), .ZN(n9238) );
  INV_X1 U9999 ( .A(n9238), .ZN(n8439) );
  INV_X1 U10000 ( .A(n8440), .ZN(n9219) );
  NAND2_X1 U10001 ( .A1(n9340), .A2(n9219), .ZN(n8441) );
  OR2_X1 U10002 ( .A1(n9335), .A2(n9209), .ZN(n8442) );
  NAND2_X1 U10003 ( .A1(n9329), .A2(n9218), .ZN(n8443) );
  INV_X1 U10004 ( .A(n9321), .ZN(n9171) );
  INV_X1 U10005 ( .A(n8558), .ZN(n9175) );
  AOI22_X1 U10006 ( .A1(n9152), .A2(n9153), .B1(n9175), .B2(n9315), .ZN(n9136)
         );
  INV_X1 U10007 ( .A(n9310), .ZN(n9141) );
  INV_X1 U10008 ( .A(n8540), .ZN(n9131) );
  NAND2_X1 U10009 ( .A1(n8449), .A2(n8604), .ZN(n8450) );
  NAND2_X1 U10010 ( .A1(n9073), .A2(n9072), .ZN(n9071) );
  INV_X1 U10011 ( .A(n8522), .ZN(n9066) );
  NAND2_X1 U10012 ( .A1(n9071), .A2(n8451), .ZN(n9056) );
  NAND2_X1 U10013 ( .A1(n9056), .A2(n9064), .ZN(n9055) );
  NAND2_X1 U10014 ( .A1(n9055), .A2(n8452), .ZN(n9037) );
  NAND2_X1 U10015 ( .A1(n8347), .A2(n8342), .ZN(n8453) );
  INV_X1 U10016 ( .A(n9340), .ZN(n9255) );
  NAND2_X1 U10017 ( .A1(n9137), .A2(n9128), .ZN(n9122) );
  INV_X1 U10018 ( .A(n9045), .ZN(n8455) );
  INV_X1 U10019 ( .A(n9274), .ZN(n8458) );
  AOI21_X1 U10020 ( .B1(n9274), .B2(n8455), .A(n8679), .ZN(n9275) );
  AOI22_X1 U10021 ( .A1(n8456), .A2(n10373), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n10372), .ZN(n8457) );
  OAI21_X1 U10022 ( .B1(n8458), .B2(n9254), .A(n8457), .ZN(n8469) );
  OAI21_X1 U10023 ( .B1(n8461), .B2(n8460), .A(n8459), .ZN(n8467) );
  NAND2_X1 U10024 ( .A1(n9065), .A2(n10366), .ZN(n8465) );
  INV_X1 U10025 ( .A(n9385), .ZN(n8462) );
  NAND2_X1 U10026 ( .A1(n8462), .A2(P2_B_REG_SCAN_IN), .ZN(n8463) );
  AND2_X1 U10027 ( .A1(n10368), .A2(n8463), .ZN(n8672) );
  NAND2_X1 U10028 ( .A1(n8613), .A2(n8672), .ZN(n8464) );
  NOR2_X1 U10029 ( .A1(n9276), .A2(n10372), .ZN(n8468) );
  OAI21_X1 U10030 ( .B1(n9279), .B2(n9233), .A(n8470), .ZN(P2_U3267) );
  INV_X1 U10031 ( .A(n8471), .ZN(n9375) );
  OAI222_X1 U10032 ( .A1(n9886), .A2(n9375), .B1(n5874), .B2(P1_U3084), .C1(
        n8472), .C2(n9891), .ZN(P1_U3324) );
  OAI222_X1 U10033 ( .A1(n9891), .A2(n8474), .B1(n9886), .B2(n8473), .C1(n6481), .C2(P1_U3084), .ZN(P1_U3331) );
  INV_X1 U10034 ( .A(n8476), .ZN(n8477) );
  AOI21_X1 U10035 ( .B1(n8475), .B2(n8477), .A(n10246), .ZN(n8481) );
  NOR3_X1 U10036 ( .A1(n8478), .A2(n8522), .A3(n8603), .ZN(n8480) );
  OAI21_X1 U10037 ( .B1(n8481), .B2(n8480), .A(n8479), .ZN(n8485) );
  AOI22_X1 U10038 ( .A1(n9060), .A2(n8597), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3152), .ZN(n8482) );
  OAI21_X1 U10039 ( .B1(n8522), .B2(n10252), .A(n8482), .ZN(n8483) );
  AOI21_X1 U10040 ( .B1(n9065), .B2(n8610), .A(n8483), .ZN(n8484) );
  OAI211_X1 U10041 ( .C1(n9062), .C2(n4871), .A(n8485), .B(n8484), .ZN(
        P2_U3216) );
  INV_X1 U10042 ( .A(n8486), .ZN(n8488) );
  NOR2_X1 U10043 ( .A1(n8488), .A2(n8487), .ZN(n8537) );
  INV_X1 U10044 ( .A(n8603), .ZN(n10263) );
  AOI22_X1 U10045 ( .A1(n8486), .A2(n10287), .B1(n10263), .B2(n9113), .ZN(
        n8493) );
  OAI22_X1 U10046 ( .A1(n8540), .A2(n10260), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8871), .ZN(n8489) );
  AOI21_X1 U10047 ( .B1(n10257), .B2(n8444), .A(n8489), .ZN(n8490) );
  OAI21_X1 U10048 ( .B1(n9125), .B2(n10292), .A(n8490), .ZN(n8491) );
  AOI21_X1 U10049 ( .B1(n9305), .B2(n10286), .A(n8491), .ZN(n8492) );
  OAI21_X1 U10050 ( .B1(n8537), .B2(n8493), .A(n8492), .ZN(P2_U3218) );
  OAI21_X1 U10051 ( .B1(n8497), .B2(n8591), .A(n8495), .ZN(n8503) );
  NOR3_X1 U10052 ( .A1(n8497), .A2(n8496), .A3(n8603), .ZN(n8498) );
  OAI21_X1 U10053 ( .B1(n8498), .B2(n10257), .A(n9218), .ZN(n8501) );
  NAND2_X1 U10054 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8670) );
  OAI21_X1 U10055 ( .B1(n10260), .B2(n8615), .A(n8670), .ZN(n8499) );
  AOI21_X1 U10056 ( .B1(n9196), .B2(n8597), .A(n8499), .ZN(n8500) );
  OAI211_X1 U10057 ( .C1(n9188), .C2(n4871), .A(n8501), .B(n8500), .ZN(n8502)
         );
  AOI21_X1 U10058 ( .B1(n8503), .B2(n10287), .A(n8502), .ZN(n8504) );
  INV_X1 U10059 ( .A(n8504), .ZN(P2_U3221) );
  OAI21_X1 U10060 ( .B1(n8506), .B2(n8505), .A(n8582), .ZN(n8507) );
  NAND2_X1 U10061 ( .A1(n8507), .A2(n10287), .ZN(n8510) );
  AOI22_X1 U10062 ( .A1(n10286), .A2(n6546), .B1(n8575), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n8509) );
  AOI22_X1 U10063 ( .A1(n8610), .A2(n8626), .B1(n10257), .B2(n8629), .ZN(n8508) );
  NAND3_X1 U10064 ( .A1(n8510), .A2(n8509), .A3(n8508), .ZN(P2_U3224) );
  INV_X1 U10065 ( .A(n9315), .ZN(n9157) );
  INV_X1 U10066 ( .A(n8511), .ZN(n8512) );
  AOI21_X1 U10067 ( .B1(n8551), .B2(n8512), .A(n10246), .ZN(n8515) );
  NOR3_X1 U10068 ( .A1(n8513), .A2(n8615), .A3(n8603), .ZN(n8514) );
  OAI21_X1 U10069 ( .B1(n8515), .B2(n8514), .A(n8564), .ZN(n8519) );
  AOI22_X1 U10070 ( .A1(n8444), .A2(n8610), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8516) );
  OAI21_X1 U10071 ( .B1(n8615), .B2(n10252), .A(n8516), .ZN(n8517) );
  AOI21_X1 U10072 ( .B1(n9155), .B2(n8597), .A(n8517), .ZN(n8518) );
  OAI211_X1 U10073 ( .C1(n9157), .C2(n4871), .A(n8519), .B(n8518), .ZN(
        P2_U3225) );
  OAI211_X1 U10074 ( .C1(n8521), .C2(n8520), .A(n8602), .B(n10287), .ZN(n8526)
         );
  OAI22_X1 U10075 ( .A1(n8522), .A2(n9240), .B1(n8540), .B2(n9242), .ZN(n9099)
         );
  OAI22_X1 U10076 ( .A1(n9094), .A2(n10292), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8523), .ZN(n8524) );
  AOI21_X1 U10077 ( .B1(n9099), .B2(n10279), .A(n8524), .ZN(n8525) );
  OAI211_X1 U10078 ( .C1(n8449), .C2(n4871), .A(n8526), .B(n8525), .ZN(
        P2_U3227) );
  AOI21_X1 U10079 ( .B1(n8528), .B2(n8527), .A(n10246), .ZN(n8529) );
  NAND2_X1 U10080 ( .A1(n8529), .A2(n8589), .ZN(n8535) );
  NOR2_X1 U10081 ( .A1(n10292), .A2(n9225), .ZN(n8533) );
  OAI21_X1 U10082 ( .B1(n10260), .B2(n8531), .A(n8530), .ZN(n8532) );
  AOI211_X1 U10083 ( .C1(n10257), .C2(n9219), .A(n8533), .B(n8532), .ZN(n8534)
         );
  OAI211_X1 U10084 ( .C1(n4721), .C2(n4871), .A(n8535), .B(n8534), .ZN(
        P2_U3230) );
  INV_X1 U10085 ( .A(n9300), .ZN(n9108) );
  NOR2_X1 U10086 ( .A1(n8537), .A2(n8536), .ZN(n8539) );
  XNOR2_X1 U10087 ( .A(n8539), .B(n8538), .ZN(n8543) );
  OAI22_X1 U10088 ( .A1(n8543), .A2(n10246), .B1(n8540), .B2(n8603), .ZN(n8541) );
  OAI21_X1 U10089 ( .B1(n8543), .B2(n8542), .A(n8541), .ZN(n8548) );
  AOI22_X1 U10090 ( .A1(n9114), .A2(n8610), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n8544) );
  OAI21_X1 U10091 ( .B1(n8545), .B2(n10252), .A(n8544), .ZN(n8546) );
  AOI21_X1 U10092 ( .B1(n9106), .B2(n8597), .A(n8546), .ZN(n8547) );
  OAI211_X1 U10093 ( .C1(n9108), .C2(n4871), .A(n8548), .B(n8547), .ZN(
        P2_U3231) );
  AOI21_X1 U10094 ( .B1(n8550), .B2(n8549), .A(n10246), .ZN(n8552) );
  NAND2_X1 U10095 ( .A1(n8552), .A2(n8551), .ZN(n8557) );
  INV_X1 U10096 ( .A(n8553), .ZN(n9169) );
  AOI22_X1 U10097 ( .A1(n9175), .A2(n8610), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3152), .ZN(n8554) );
  OAI21_X1 U10098 ( .B1(n8595), .B2(n10252), .A(n8554), .ZN(n8555) );
  AOI21_X1 U10099 ( .B1(n9169), .B2(n8597), .A(n8555), .ZN(n8556) );
  OAI211_X1 U10100 ( .C1(n9171), .C2(n4871), .A(n8557), .B(n8556), .ZN(
        P2_U3235) );
  NAND2_X1 U10101 ( .A1(n9113), .A2(n10368), .ZN(n8560) );
  OR2_X1 U10102 ( .A1(n8558), .A2(n9242), .ZN(n8559) );
  NAND2_X1 U10103 ( .A1(n8560), .A2(n8559), .ZN(n9147) );
  AOI22_X1 U10104 ( .A1(n9147), .A2(n10279), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3152), .ZN(n8561) );
  OAI21_X1 U10105 ( .B1(n9138), .B2(n10292), .A(n8561), .ZN(n8569) );
  INV_X1 U10106 ( .A(n8562), .ZN(n8563) );
  NAND2_X1 U10107 ( .A1(n8564), .A2(n8563), .ZN(n8566) );
  XNOR2_X1 U10108 ( .A(n8566), .B(n8565), .ZN(n8571) );
  NOR3_X1 U10109 ( .A1(n8571), .A2(n8567), .A3(n8603), .ZN(n8568) );
  AOI211_X1 U10110 ( .C1(n10286), .C2(n9310), .A(n8569), .B(n8568), .ZN(n8573)
         );
  NAND3_X1 U10111 ( .A1(n8571), .A2(n10287), .A3(n8570), .ZN(n8572) );
  NAND2_X1 U10112 ( .A1(n8573), .A2(n8572), .ZN(P2_U3237) );
  OR2_X1 U10113 ( .A1(n8574), .A2(n10246), .ZN(n8586) );
  AOI22_X1 U10114 ( .A1(n10286), .A2(n8576), .B1(n8575), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n8585) );
  AOI22_X1 U10115 ( .A1(n8610), .A2(n8625), .B1(n10257), .B2(n8627), .ZN(n8584) );
  NAND2_X1 U10116 ( .A1(n10287), .A2(n8578), .ZN(n8579) );
  OAI21_X1 U10117 ( .B1(n8603), .B2(n8580), .A(n8579), .ZN(n8581) );
  NAND3_X1 U10118 ( .A1(n8582), .A2(n4858), .A3(n8581), .ZN(n8583) );
  NAND4_X1 U10119 ( .A1(n8586), .A2(n8585), .A3(n8584), .A4(n8583), .ZN(
        P2_U3239) );
  INV_X1 U10120 ( .A(n9329), .ZN(n9206) );
  INV_X1 U10121 ( .A(n8587), .ZN(n8588) );
  AOI21_X1 U10122 ( .B1(n8589), .B2(n8588), .A(n10246), .ZN(n8593) );
  NOR3_X1 U10123 ( .A1(n8590), .A2(n9241), .A3(n8603), .ZN(n8592) );
  OAI21_X1 U10124 ( .B1(n8593), .B2(n8592), .A(n8591), .ZN(n8599) );
  NAND2_X1 U10125 ( .A1(n10257), .A2(n9209), .ZN(n8594) );
  NAND2_X1 U10126 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8644) );
  OAI211_X1 U10127 ( .C1(n8595), .C2(n10260), .A(n8594), .B(n8644), .ZN(n8596)
         );
  AOI21_X1 U10128 ( .B1(n9204), .B2(n8597), .A(n8596), .ZN(n8598) );
  OAI211_X1 U10129 ( .C1(n9206), .C2(n4871), .A(n8599), .B(n8598), .ZN(
        P2_U3240) );
  INV_X1 U10130 ( .A(n9291), .ZN(n9079) );
  INV_X1 U10131 ( .A(n8600), .ZN(n8601) );
  AOI21_X1 U10132 ( .B1(n8602), .B2(n8601), .A(n10246), .ZN(n8607) );
  NOR3_X1 U10133 ( .A1(n8605), .A2(n8604), .A3(n8603), .ZN(n8606) );
  OAI21_X1 U10134 ( .B1(n8607), .B2(n8606), .A(n8475), .ZN(n8612) );
  AOI22_X1 U10135 ( .A1(n9114), .A2(n10257), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3152), .ZN(n8608) );
  OAI21_X1 U10136 ( .B1(n9076), .B2(n10292), .A(n8608), .ZN(n8609) );
  AOI21_X1 U10137 ( .B1(n8610), .B2(n9083), .A(n8609), .ZN(n8611) );
  OAI211_X1 U10138 ( .C1(n9079), .C2(n4871), .A(n8612), .B(n8611), .ZN(
        P2_U3242) );
  MUX2_X1 U10139 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8613), .S(P2_U3966), .Z(
        P2_U3582) );
  INV_X1 U10140 ( .A(n8614), .ZN(n9040) );
  MUX2_X1 U10141 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n9040), .S(P2_U3966), .Z(
        P2_U3581) );
  MUX2_X1 U10142 ( .A(n9065), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8628), .Z(
        P2_U3580) );
  MUX2_X1 U10143 ( .A(n9083), .B(P2_DATAO_REG_27__SCAN_IN), .S(n8628), .Z(
        P2_U3579) );
  MUX2_X1 U10144 ( .A(n9066), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8628), .Z(
        P2_U3578) );
  MUX2_X1 U10145 ( .A(n9114), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8628), .Z(
        P2_U3577) );
  MUX2_X1 U10146 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9131), .S(P2_U3966), .Z(
        P2_U3576) );
  MUX2_X1 U10147 ( .A(n8444), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8628), .Z(
        P2_U3574) );
  MUX2_X1 U10148 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9175), .S(P2_U3966), .Z(
        P2_U3573) );
  INV_X1 U10149 ( .A(n8615), .ZN(n9186) );
  MUX2_X1 U10150 ( .A(n9186), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8628), .Z(
        P2_U3572) );
  MUX2_X1 U10151 ( .A(n9210), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8628), .Z(
        P2_U3571) );
  MUX2_X1 U10152 ( .A(n9218), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8628), .Z(
        P2_U3570) );
  MUX2_X1 U10153 ( .A(n9209), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8628), .Z(
        P2_U3569) );
  MUX2_X1 U10154 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9219), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10155 ( .A(n8616), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8628), .Z(
        P2_U3567) );
  MUX2_X1 U10156 ( .A(n8617), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8628), .Z(
        P2_U3566) );
  MUX2_X1 U10157 ( .A(n8618), .B(P2_DATAO_REG_13__SCAN_IN), .S(n8628), .Z(
        P2_U3565) );
  MUX2_X1 U10158 ( .A(n8619), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8628), .Z(
        P2_U3564) );
  MUX2_X1 U10159 ( .A(n10262), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8628), .Z(
        P2_U3563) );
  MUX2_X1 U10160 ( .A(n8620), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8628), .Z(
        P2_U3562) );
  MUX2_X1 U10161 ( .A(n8621), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8628), .Z(
        P2_U3561) );
  MUX2_X1 U10162 ( .A(n8622), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8628), .Z(
        P2_U3560) );
  MUX2_X1 U10163 ( .A(n10369), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8628), .Z(
        P2_U3559) );
  MUX2_X1 U10164 ( .A(n8623), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8628), .Z(
        P2_U3558) );
  MUX2_X1 U10165 ( .A(n10367), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8628), .Z(
        P2_U3557) );
  MUX2_X1 U10166 ( .A(n8624), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8628), .Z(
        P2_U3556) );
  MUX2_X1 U10167 ( .A(n8625), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8628), .Z(
        P2_U3555) );
  MUX2_X1 U10168 ( .A(n8626), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8628), .Z(
        P2_U3554) );
  MUX2_X1 U10169 ( .A(n8627), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8628), .Z(
        P2_U3553) );
  MUX2_X1 U10170 ( .A(n8629), .B(P2_DATAO_REG_0__SCAN_IN), .S(n8628), .Z(
        P2_U3552) );
  OAI211_X1 U10171 ( .C1(n8632), .C2(n8631), .A(n10332), .B(n8630), .ZN(n8641)
         );
  AOI21_X1 U10172 ( .B1(n10328), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n8633), .ZN(
        n8640) );
  NAND2_X1 U10173 ( .A1(n10330), .A2(n8634), .ZN(n8639) );
  OAI211_X1 U10174 ( .C1(n8637), .C2(n8636), .A(n10336), .B(n8635), .ZN(n8638)
         );
  NAND4_X1 U10175 ( .A1(n8641), .A2(n8640), .A3(n8639), .A4(n8638), .ZN(
        P2_U3253) );
  OAI21_X1 U10176 ( .B1(n8646), .B2(n9226), .A(n8642), .ZN(n8658) );
  XNOR2_X1 U10177 ( .A(n8658), .B(n8656), .ZN(n8643) );
  NAND2_X1 U10178 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n8643), .ZN(n8660) );
  OAI211_X1 U10179 ( .C1(n8643), .C2(P2_REG2_REG_18__SCAN_IN), .A(n10332), .B(
        n8660), .ZN(n8655) );
  INV_X1 U10180 ( .A(n8644), .ZN(n8653) );
  OAI21_X1 U10181 ( .B1(n8647), .B2(n8646), .A(n8645), .ZN(n8650) );
  NAND2_X1 U10182 ( .A1(n8656), .A2(n8648), .ZN(n8662) );
  OAI21_X1 U10183 ( .B1(n8656), .B2(n8648), .A(n8662), .ZN(n8649) );
  NOR2_X1 U10184 ( .A1(n8649), .A2(n8650), .ZN(n8664) );
  AOI21_X1 U10185 ( .B1(n8650), .B2(n8649), .A(n8664), .ZN(n8651) );
  NOR2_X1 U10186 ( .A1(n8651), .A2(n10294), .ZN(n8652) );
  AOI211_X1 U10187 ( .C1(n10328), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n8653), .B(
        n8652), .ZN(n8654) );
  OAI211_X1 U10188 ( .C1(n10293), .C2(n8656), .A(n8655), .B(n8654), .ZN(
        P2_U3263) );
  NAND2_X1 U10189 ( .A1(n8658), .A2(n8657), .ZN(n8659) );
  NAND2_X1 U10190 ( .A1(n8660), .A2(n8659), .ZN(n8661) );
  XOR2_X1 U10191 ( .A(n8661), .B(P2_REG2_REG_19__SCAN_IN), .Z(n8667) );
  INV_X1 U10192 ( .A(n8662), .ZN(n8663) );
  NOR2_X1 U10193 ( .A1(n8664), .A2(n8663), .ZN(n8665) );
  XNOR2_X1 U10194 ( .A(n8665), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8668) );
  INV_X1 U10195 ( .A(n8668), .ZN(n8666) );
  AOI22_X1 U10196 ( .A1(n8667), .A2(n10332), .B1(n8666), .B2(n10336), .ZN(
        n8669) );
  NAND2_X1 U10197 ( .A1(n9273), .A2(n8679), .ZN(n9269) );
  XNOR2_X1 U10198 ( .A(n9269), .B(n9266), .ZN(n9268) );
  NAND2_X1 U10199 ( .A1(n8673), .A2(n8672), .ZN(n9271) );
  INV_X1 U10200 ( .A(n9271), .ZN(n8674) );
  NAND2_X1 U10201 ( .A1(n8674), .A2(n9259), .ZN(n8681) );
  OAI21_X1 U10202 ( .B1(n9259), .B2(n8675), .A(n8681), .ZN(n8676) );
  AOI21_X1 U10203 ( .B1(n9266), .B2(n10355), .A(n8676), .ZN(n8677) );
  OAI21_X1 U10204 ( .B1(n9268), .B2(n8678), .A(n8677), .ZN(P2_U3265) );
  INV_X1 U10205 ( .A(n8679), .ZN(n8680) );
  NAND2_X1 U10206 ( .A1(n8683), .A2(n8680), .ZN(n9270) );
  NAND3_X1 U10207 ( .A1(n9270), .A2(n9262), .A3(n9269), .ZN(n8685) );
  OAI21_X1 U10208 ( .B1(n5643), .B2(n9259), .A(n8681), .ZN(n8682) );
  AOI21_X1 U10209 ( .B1(n8683), .B2(n10355), .A(n8682), .ZN(n8684) );
  NAND2_X1 U10210 ( .A1(n8685), .A2(n8684), .ZN(P2_U3266) );
  AOI22_X1 U10211 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(keyinput179), .B1(SI_4_), 
        .B2(keyinput135), .ZN(n8686) );
  OAI221_X1 U10212 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(keyinput179), .C1(SI_4_), 
        .C2(keyinput135), .A(n8686), .ZN(n8693) );
  AOI22_X1 U10213 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(keyinput229), .B1(
        P2_D_REG_1__SCAN_IN), .B2(keyinput163), .ZN(n8687) );
  OAI221_X1 U10214 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput229), .C1(
        P2_D_REG_1__SCAN_IN), .C2(keyinput163), .A(n8687), .ZN(n8692) );
  AOI22_X1 U10215 ( .A1(P2_REG1_REG_5__SCAN_IN), .A2(keyinput212), .B1(
        P1_REG2_REG_12__SCAN_IN), .B2(keyinput128), .ZN(n8688) );
  OAI221_X1 U10216 ( .B1(P2_REG1_REG_5__SCAN_IN), .B2(keyinput212), .C1(
        P1_REG2_REG_12__SCAN_IN), .C2(keyinput128), .A(n8688), .ZN(n8691) );
  AOI22_X1 U10217 ( .A1(P2_REG0_REG_31__SCAN_IN), .A2(keyinput148), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(keyinput162), .ZN(n8689) );
  OAI221_X1 U10218 ( .B1(P2_REG0_REG_31__SCAN_IN), .B2(keyinput148), .C1(
        P1_REG2_REG_1__SCAN_IN), .C2(keyinput162), .A(n8689), .ZN(n8690) );
  NOR4_X1 U10219 ( .A1(n8693), .A2(n8692), .A3(n8691), .A4(n8690), .ZN(n8721)
         );
  AOI22_X1 U10220 ( .A1(P2_REG0_REG_10__SCAN_IN), .A2(keyinput134), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput168), .ZN(n8694) );
  OAI221_X1 U10221 ( .B1(P2_REG0_REG_10__SCAN_IN), .B2(keyinput134), .C1(
        P1_IR_REG_19__SCAN_IN), .C2(keyinput168), .A(n8694), .ZN(n8701) );
  AOI22_X1 U10222 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(keyinput223), .B1(
        P1_D_REG_16__SCAN_IN), .B2(keyinput172), .ZN(n8695) );
  OAI221_X1 U10223 ( .B1(P1_REG2_REG_10__SCAN_IN), .B2(keyinput223), .C1(
        P1_D_REG_16__SCAN_IN), .C2(keyinput172), .A(n8695), .ZN(n8700) );
  AOI22_X1 U10224 ( .A1(P2_REG2_REG_30__SCAN_IN), .A2(keyinput199), .B1(
        P2_D_REG_15__SCAN_IN), .B2(keyinput200), .ZN(n8696) );
  OAI221_X1 U10225 ( .B1(P2_REG2_REG_30__SCAN_IN), .B2(keyinput199), .C1(
        P2_D_REG_15__SCAN_IN), .C2(keyinput200), .A(n8696), .ZN(n8699) );
  AOI22_X1 U10226 ( .A1(P2_REG2_REG_23__SCAN_IN), .A2(keyinput146), .B1(
        P2_REG0_REG_8__SCAN_IN), .B2(keyinput240), .ZN(n8697) );
  OAI221_X1 U10227 ( .B1(P2_REG2_REG_23__SCAN_IN), .B2(keyinput146), .C1(
        P2_REG0_REG_8__SCAN_IN), .C2(keyinput240), .A(n8697), .ZN(n8698) );
  NOR4_X1 U10228 ( .A1(n8701), .A2(n8700), .A3(n8699), .A4(n8698), .ZN(n8720)
         );
  AOI22_X1 U10229 ( .A1(P1_REG2_REG_3__SCAN_IN), .A2(keyinput204), .B1(
        P1_REG3_REG_9__SCAN_IN), .B2(keyinput252), .ZN(n8702) );
  OAI221_X1 U10230 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(keyinput204), .C1(
        P1_REG3_REG_9__SCAN_IN), .C2(keyinput252), .A(n8702), .ZN(n8709) );
  AOI22_X1 U10231 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput242), .B1(
        P2_REG1_REG_9__SCAN_IN), .B2(keyinput196), .ZN(n8703) );
  OAI221_X1 U10232 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput242), .C1(
        P2_REG1_REG_9__SCAN_IN), .C2(keyinput196), .A(n8703), .ZN(n8708) );
  AOI22_X1 U10233 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(keyinput177), .B1(
        P1_B_REG_SCAN_IN), .B2(keyinput203), .ZN(n8704) );
  OAI221_X1 U10234 ( .B1(P1_REG3_REG_11__SCAN_IN), .B2(keyinput177), .C1(
        P1_B_REG_SCAN_IN), .C2(keyinput203), .A(n8704), .ZN(n8707) );
  AOI22_X1 U10235 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(keyinput192), .B1(
        P1_REG1_REG_20__SCAN_IN), .B2(keyinput166), .ZN(n8705) );
  OAI221_X1 U10236 ( .B1(P2_REG3_REG_27__SCAN_IN), .B2(keyinput192), .C1(
        P1_REG1_REG_20__SCAN_IN), .C2(keyinput166), .A(n8705), .ZN(n8706) );
  NOR4_X1 U10237 ( .A1(n8709), .A2(n8708), .A3(n8707), .A4(n8706), .ZN(n8719)
         );
  AOI22_X1 U10238 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(keyinput178), .B1(
        P1_REG3_REG_6__SCAN_IN), .B2(keyinput175), .ZN(n8710) );
  OAI221_X1 U10239 ( .B1(P1_DATAO_REG_29__SCAN_IN), .B2(keyinput178), .C1(
        P1_REG3_REG_6__SCAN_IN), .C2(keyinput175), .A(n8710), .ZN(n8717) );
  AOI22_X1 U10240 ( .A1(P2_REG1_REG_1__SCAN_IN), .A2(keyinput149), .B1(
        P1_D_REG_4__SCAN_IN), .B2(keyinput187), .ZN(n8711) );
  OAI221_X1 U10241 ( .B1(P2_REG1_REG_1__SCAN_IN), .B2(keyinput149), .C1(
        P1_D_REG_4__SCAN_IN), .C2(keyinput187), .A(n8711), .ZN(n8716) );
  AOI22_X1 U10242 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(keyinput137), .B1(
        P1_IR_REG_2__SCAN_IN), .B2(keyinput197), .ZN(n8712) );
  OAI221_X1 U10243 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(keyinput137), .C1(
        P1_IR_REG_2__SCAN_IN), .C2(keyinput197), .A(n8712), .ZN(n8715) );
  AOI22_X1 U10244 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(keyinput191), .B1(
        P1_REG3_REG_27__SCAN_IN), .B2(keyinput157), .ZN(n8713) );
  OAI221_X1 U10245 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(keyinput191), .C1(
        P1_REG3_REG_27__SCAN_IN), .C2(keyinput157), .A(n8713), .ZN(n8714) );
  NOR4_X1 U10246 ( .A1(n8717), .A2(n8716), .A3(n8715), .A4(n8714), .ZN(n8718)
         );
  NAND4_X1 U10247 ( .A1(n8721), .A2(n8720), .A3(n8719), .A4(n8718), .ZN(n8854)
         );
  AOI22_X1 U10248 ( .A1(P2_REG2_REG_8__SCAN_IN), .A2(keyinput184), .B1(
        P1_D_REG_29__SCAN_IN), .B2(keyinput164), .ZN(n8722) );
  OAI221_X1 U10249 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(keyinput184), .C1(
        P1_D_REG_29__SCAN_IN), .C2(keyinput164), .A(n8722), .ZN(n8729) );
  AOI22_X1 U10250 ( .A1(P2_D_REG_17__SCAN_IN), .A2(keyinput152), .B1(
        P1_IR_REG_3__SCAN_IN), .B2(keyinput201), .ZN(n8723) );
  OAI221_X1 U10251 ( .B1(P2_D_REG_17__SCAN_IN), .B2(keyinput152), .C1(
        P1_IR_REG_3__SCAN_IN), .C2(keyinput201), .A(n8723), .ZN(n8728) );
  AOI22_X1 U10252 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(keyinput159), .B1(
        P1_REG0_REG_16__SCAN_IN), .B2(keyinput185), .ZN(n8724) );
  OAI221_X1 U10253 ( .B1(P2_IR_REG_15__SCAN_IN), .B2(keyinput159), .C1(
        P1_REG0_REG_16__SCAN_IN), .C2(keyinput185), .A(n8724), .ZN(n8727) );
  AOI22_X1 U10254 ( .A1(SI_1_), .A2(keyinput140), .B1(P1_DATAO_REG_4__SCAN_IN), 
        .B2(keyinput170), .ZN(n8725) );
  OAI221_X1 U10255 ( .B1(SI_1_), .B2(keyinput140), .C1(P1_DATAO_REG_4__SCAN_IN), .C2(keyinput170), .A(n8725), .ZN(n8726) );
  NOR4_X1 U10256 ( .A1(n8729), .A2(n8728), .A3(n8727), .A4(n8726), .ZN(n8758)
         );
  AOI22_X1 U10257 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput129), .B1(
        P1_D_REG_12__SCAN_IN), .B2(keyinput233), .ZN(n8730) );
  OAI221_X1 U10258 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput129), .C1(
        P1_D_REG_12__SCAN_IN), .C2(keyinput233), .A(n8730), .ZN(n8737) );
  AOI22_X1 U10259 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(keyinput153), .B1(
        P1_REG3_REG_25__SCAN_IN), .B2(keyinput132), .ZN(n8731) );
  OAI221_X1 U10260 ( .B1(P2_IR_REG_11__SCAN_IN), .B2(keyinput153), .C1(
        P1_REG3_REG_25__SCAN_IN), .C2(keyinput132), .A(n8731), .ZN(n8736) );
  AOI22_X1 U10261 ( .A1(P2_D_REG_8__SCAN_IN), .A2(keyinput202), .B1(SI_26_), 
        .B2(keyinput193), .ZN(n8732) );
  OAI221_X1 U10262 ( .B1(P2_D_REG_8__SCAN_IN), .B2(keyinput202), .C1(SI_26_), 
        .C2(keyinput193), .A(n8732), .ZN(n8735) );
  AOI22_X1 U10263 ( .A1(P2_REG2_REG_17__SCAN_IN), .A2(keyinput222), .B1(
        P2_IR_REG_7__SCAN_IN), .B2(keyinput189), .ZN(n8733) );
  OAI221_X1 U10264 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(keyinput222), .C1(
        P2_IR_REG_7__SCAN_IN), .C2(keyinput189), .A(n8733), .ZN(n8734) );
  NOR4_X1 U10265 ( .A1(n8737), .A2(n8736), .A3(n8735), .A4(n8734), .ZN(n8757)
         );
  INV_X1 U10266 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10393) );
  AOI22_X1 U10267 ( .A1(P1_REG1_REG_26__SCAN_IN), .A2(keyinput165), .B1(n10393), .B2(keyinput167), .ZN(n8738) );
  OAI221_X1 U10268 ( .B1(P1_REG1_REG_26__SCAN_IN), .B2(keyinput165), .C1(
        n10393), .C2(keyinput167), .A(n8738), .ZN(n8745) );
  INV_X1 U10269 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n8882) );
  AOI22_X1 U10270 ( .A1(n8915), .A2(keyinput224), .B1(n8882), .B2(keyinput144), 
        .ZN(n8739) );
  OAI221_X1 U10271 ( .B1(n8915), .B2(keyinput224), .C1(n8882), .C2(keyinput144), .A(n8739), .ZN(n8744) );
  INV_X1 U10272 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n8909) );
  AOI22_X1 U10273 ( .A1(n8909), .A2(keyinput176), .B1(n8923), .B2(keyinput158), 
        .ZN(n8740) );
  OAI221_X1 U10274 ( .B1(n8909), .B2(keyinput176), .C1(n8923), .C2(keyinput158), .A(n8740), .ZN(n8743) );
  AOI22_X1 U10275 ( .A1(n6051), .A2(keyinput243), .B1(keyinput147), .B2(n8859), 
        .ZN(n8741) );
  OAI221_X1 U10276 ( .B1(n6051), .B2(keyinput243), .C1(n8859), .C2(keyinput147), .A(n8741), .ZN(n8742) );
  NOR4_X1 U10277 ( .A1(n8745), .A2(n8744), .A3(n8743), .A4(n8742), .ZN(n8756)
         );
  INV_X1 U10278 ( .A(P2_D_REG_30__SCAN_IN), .ZN(n10387) );
  AOI22_X1 U10279 ( .A1(n9546), .A2(keyinput238), .B1(keyinput174), .B2(n10387), .ZN(n8746) );
  OAI221_X1 U10280 ( .B1(n9546), .B2(keyinput238), .C1(n10387), .C2(
        keyinput174), .A(n8746), .ZN(n8754) );
  AOI22_X1 U10281 ( .A1(n7530), .A2(keyinput246), .B1(keyinput241), .B2(n8873), 
        .ZN(n8747) );
  OAI221_X1 U10282 ( .B1(n7530), .B2(keyinput246), .C1(n8873), .C2(keyinput241), .A(n8747), .ZN(n8753) );
  AOI22_X1 U10283 ( .A1(n8749), .A2(keyinput215), .B1(keyinput156), .B2(n9436), 
        .ZN(n8748) );
  OAI221_X1 U10284 ( .B1(n8749), .B2(keyinput215), .C1(n9436), .C2(keyinput156), .A(n8748), .ZN(n8752) );
  AOI22_X1 U10285 ( .A1(n5175), .A2(keyinput247), .B1(keyinput155), .B2(n10514), .ZN(n8750) );
  OAI221_X1 U10286 ( .B1(n5175), .B2(keyinput247), .C1(n10514), .C2(
        keyinput155), .A(n8750), .ZN(n8751) );
  NOR4_X1 U10287 ( .A1(n8754), .A2(n8753), .A3(n8752), .A4(n8751), .ZN(n8755)
         );
  NAND4_X1 U10288 ( .A1(n8758), .A2(n8757), .A3(n8756), .A4(n8755), .ZN(n8853)
         );
  INV_X1 U10289 ( .A(SI_6_), .ZN(n8911) );
  AOI22_X1 U10290 ( .A1(n6139), .A2(keyinput205), .B1(n8911), .B2(keyinput221), 
        .ZN(n8759) );
  OAI221_X1 U10291 ( .B1(n6139), .B2(keyinput205), .C1(n8911), .C2(keyinput221), .A(n8759), .ZN(n8770) );
  INV_X1 U10292 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9550) );
  AOI22_X1 U10293 ( .A1(n8761), .A2(keyinput253), .B1(keyinput219), .B2(n9550), 
        .ZN(n8760) );
  OAI221_X1 U10294 ( .B1(n8761), .B2(keyinput253), .C1(n9550), .C2(keyinput219), .A(n8760), .ZN(n8769) );
  INV_X1 U10295 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n8763) );
  AOI22_X1 U10296 ( .A1(n8764), .A2(keyinput250), .B1(n8763), .B2(keyinput136), 
        .ZN(n8762) );
  OAI221_X1 U10297 ( .B1(n8764), .B2(keyinput250), .C1(n8763), .C2(keyinput136), .A(n8762), .ZN(n8768) );
  XOR2_X1 U10298 ( .A(n5838), .B(keyinput239), .Z(n8766) );
  XNOR2_X1 U10299 ( .A(P2_IR_REG_9__SCAN_IN), .B(keyinput131), .ZN(n8765) );
  NAND2_X1 U10300 ( .A1(n8766), .A2(n8765), .ZN(n8767) );
  NOR4_X1 U10301 ( .A1(n8770), .A2(n8769), .A3(n8768), .A4(n8767), .ZN(n8806)
         );
  AOI22_X1 U10302 ( .A1(n6282), .A2(keyinput231), .B1(keyinput183), .B2(n8772), 
        .ZN(n8771) );
  OAI221_X1 U10303 ( .B1(n6282), .B2(keyinput231), .C1(n8772), .C2(keyinput183), .A(n8771), .ZN(n8781) );
  AOI22_X1 U10304 ( .A1(n8774), .A2(keyinput225), .B1(keyinput216), .B2(n5379), 
        .ZN(n8773) );
  OAI221_X1 U10305 ( .B1(n8774), .B2(keyinput225), .C1(n5379), .C2(keyinput216), .A(n8773), .ZN(n8780) );
  INV_X1 U10306 ( .A(P1_D_REG_23__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U10307 ( .A1(n6804), .A2(keyinput154), .B1(n10187), .B2(keyinput195), .ZN(n8775) );
  OAI221_X1 U10308 ( .B1(n6804), .B2(keyinput154), .C1(n10187), .C2(
        keyinput195), .A(n8775), .ZN(n8779) );
  XOR2_X1 U10309 ( .A(n5083), .B(keyinput234), .Z(n8777) );
  XNOR2_X1 U10310 ( .A(P1_IR_REG_29__SCAN_IN), .B(keyinput188), .ZN(n8776) );
  NAND2_X1 U10311 ( .A1(n8777), .A2(n8776), .ZN(n8778) );
  NOR4_X1 U10312 ( .A1(n8781), .A2(n8780), .A3(n8779), .A4(n8778), .ZN(n8805)
         );
  AOI22_X1 U10313 ( .A1(n5335), .A2(keyinput180), .B1(n8913), .B2(keyinput244), 
        .ZN(n8782) );
  OAI221_X1 U10314 ( .B1(n5335), .B2(keyinput180), .C1(n8913), .C2(keyinput244), .A(n8782), .ZN(n8790) );
  INV_X1 U10315 ( .A(P2_D_REG_31__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U10316 ( .A1(n10386), .A2(keyinput227), .B1(n8898), .B2(keyinput237), .ZN(n8783) );
  OAI221_X1 U10317 ( .B1(n10386), .B2(keyinput227), .C1(n8898), .C2(
        keyinput237), .A(n8783), .ZN(n8789) );
  INV_X1 U10318 ( .A(P2_D_REG_13__SCAN_IN), .ZN(n10392) );
  AOI22_X1 U10319 ( .A1(n10392), .A2(keyinput190), .B1(P1_U3084), .B2(
        keyinput210), .ZN(n8784) );
  OAI221_X1 U10320 ( .B1(n10392), .B2(keyinput190), .C1(P1_U3084), .C2(
        keyinput210), .A(n8784), .ZN(n8788) );
  AOI22_X1 U10321 ( .A1(n8894), .A2(keyinput251), .B1(n8786), .B2(keyinput206), 
        .ZN(n8785) );
  OAI221_X1 U10322 ( .B1(n8894), .B2(keyinput251), .C1(n8786), .C2(keyinput206), .A(n8785), .ZN(n8787) );
  NOR4_X1 U10323 ( .A1(n8790), .A2(n8789), .A3(n8788), .A4(n8787), .ZN(n8804)
         );
  INV_X1 U10324 ( .A(SI_31_), .ZN(n8793) );
  AOI22_X1 U10325 ( .A1(n8793), .A2(keyinput194), .B1(n8792), .B2(keyinput173), 
        .ZN(n8791) );
  OAI221_X1 U10326 ( .B1(n8793), .B2(keyinput194), .C1(n8792), .C2(keyinput173), .A(n8791), .ZN(n8802) );
  AOI22_X1 U10327 ( .A1(n7384), .A2(keyinput171), .B1(n8795), .B2(keyinput169), 
        .ZN(n8794) );
  OAI221_X1 U10328 ( .B1(n7384), .B2(keyinput171), .C1(n8795), .C2(keyinput169), .A(n8794), .ZN(n8801) );
  AOI22_X1 U10329 ( .A1(n8797), .A2(keyinput186), .B1(n7461), .B2(keyinput160), 
        .ZN(n8796) );
  OAI221_X1 U10330 ( .B1(n8797), .B2(keyinput186), .C1(n7461), .C2(keyinput160), .A(n8796), .ZN(n8800) );
  AOI22_X1 U10331 ( .A1(n6467), .A2(keyinput138), .B1(keyinput208), .B2(n8985), 
        .ZN(n8798) );
  OAI221_X1 U10332 ( .B1(n6467), .B2(keyinput138), .C1(n8985), .C2(keyinput208), .A(n8798), .ZN(n8799) );
  NOR4_X1 U10333 ( .A1(n8802), .A2(n8801), .A3(n8800), .A4(n8799), .ZN(n8803)
         );
  NAND4_X1 U10334 ( .A1(n8806), .A2(n8805), .A3(n8804), .A4(n8803), .ZN(n8852)
         );
  INV_X1 U10335 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n8896) );
  AOI22_X1 U10336 ( .A1(n7715), .A2(keyinput226), .B1(keyinput232), .B2(n8896), 
        .ZN(n8807) );
  OAI221_X1 U10337 ( .B1(n7715), .B2(keyinput226), .C1(n8896), .C2(keyinput232), .A(n8807), .ZN(n8817) );
  AOI22_X1 U10338 ( .A1(n5260), .A2(keyinput217), .B1(n8933), .B2(keyinput213), 
        .ZN(n8808) );
  OAI221_X1 U10339 ( .B1(n5260), .B2(keyinput217), .C1(n8933), .C2(keyinput213), .A(n8808), .ZN(n8816) );
  AOI22_X1 U10340 ( .A1(n8811), .A2(keyinput230), .B1(keyinput235), .B2(n8810), 
        .ZN(n8809) );
  OAI221_X1 U10341 ( .B1(n8811), .B2(keyinput230), .C1(n8810), .C2(keyinput235), .A(n8809), .ZN(n8815) );
  AOI22_X1 U10342 ( .A1(n5127), .A2(keyinput150), .B1(n8813), .B2(keyinput248), 
        .ZN(n8812) );
  OAI221_X1 U10343 ( .B1(n5127), .B2(keyinput150), .C1(n8813), .C2(keyinput248), .A(n8812), .ZN(n8814) );
  NOR4_X1 U10344 ( .A1(n8817), .A2(n8816), .A3(n8815), .A4(n8814), .ZN(n8850)
         );
  AOI22_X1 U10345 ( .A1(n8885), .A2(keyinput207), .B1(keyinput161), .B2(n7001), 
        .ZN(n8818) );
  OAI221_X1 U10346 ( .B1(n8885), .B2(keyinput207), .C1(n7001), .C2(keyinput161), .A(n8818), .ZN(n8827) );
  AOI22_X1 U10347 ( .A1(n5089), .A2(keyinput141), .B1(n7102), .B2(keyinput182), 
        .ZN(n8819) );
  OAI221_X1 U10348 ( .B1(n5089), .B2(keyinput141), .C1(n7102), .C2(keyinput182), .A(n8819), .ZN(n8826) );
  INV_X1 U10349 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10388) );
  INV_X1 U10350 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n8821) );
  AOI22_X1 U10351 ( .A1(n10388), .A2(keyinput249), .B1(keyinput133), .B2(n8821), .ZN(n8820) );
  OAI221_X1 U10352 ( .B1(n10388), .B2(keyinput249), .C1(n8821), .C2(
        keyinput133), .A(n8820), .ZN(n8825) );
  XNOR2_X1 U10353 ( .A(P2_IR_REG_6__SCAN_IN), .B(keyinput236), .ZN(n8823) );
  XNOR2_X1 U10354 ( .A(SI_8_), .B(keyinput181), .ZN(n8822) );
  NAND2_X1 U10355 ( .A1(n8823), .A2(n8822), .ZN(n8824) );
  NOR4_X1 U10356 ( .A1(n8827), .A2(n8826), .A3(n8825), .A4(n8824), .ZN(n8849)
         );
  INV_X1 U10357 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n9924) );
  AOI22_X1 U10358 ( .A1(n9924), .A2(keyinput143), .B1(n6456), .B2(keyinput211), 
        .ZN(n8828) );
  OAI221_X1 U10359 ( .B1(n9924), .B2(keyinput143), .C1(n6456), .C2(keyinput211), .A(n8828), .ZN(n8837) );
  AOI22_X1 U10360 ( .A1(n6378), .A2(keyinput254), .B1(n8880), .B2(keyinput139), 
        .ZN(n8829) );
  OAI221_X1 U10361 ( .B1(n6378), .B2(keyinput254), .C1(n8880), .C2(keyinput139), .A(n8829), .ZN(n8836) );
  INV_X1 U10362 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n8899) );
  AOI22_X1 U10363 ( .A1(n8899), .A2(keyinput245), .B1(keyinput209), .B2(n8831), 
        .ZN(n8830) );
  OAI221_X1 U10364 ( .B1(n8899), .B2(keyinput245), .C1(n8831), .C2(keyinput209), .A(n8830), .ZN(n8835) );
  INV_X1 U10365 ( .A(P2_D_REG_23__SCAN_IN), .ZN(n10389) );
  AOI22_X1 U10366 ( .A1(n10389), .A2(keyinput198), .B1(n8833), .B2(keyinput218), .ZN(n8832) );
  OAI221_X1 U10367 ( .B1(n10389), .B2(keyinput198), .C1(n8833), .C2(
        keyinput218), .A(n8832), .ZN(n8834) );
  NOR4_X1 U10368 ( .A1(n8837), .A2(n8836), .A3(n8835), .A4(n8834), .ZN(n8848)
         );
  INV_X1 U10369 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9932) );
  INV_X1 U10370 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10191) );
  AOI22_X1 U10371 ( .A1(n9932), .A2(keyinput151), .B1(n10191), .B2(keyinput228), .ZN(n8838) );
  OAI221_X1 U10372 ( .B1(n9932), .B2(keyinput151), .C1(n10191), .C2(
        keyinput228), .A(n8838), .ZN(n8846) );
  INV_X1 U10373 ( .A(P1_D_REG_17__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U10374 ( .A1(n8856), .A2(keyinput145), .B1(n10188), .B2(keyinput220), .ZN(n8839) );
  OAI221_X1 U10375 ( .B1(n8856), .B2(keyinput145), .C1(n10188), .C2(
        keyinput220), .A(n8839), .ZN(n8845) );
  AOI22_X1 U10376 ( .A1(n7359), .A2(keyinput214), .B1(n6264), .B2(keyinput255), 
        .ZN(n8840) );
  OAI221_X1 U10377 ( .B1(n7359), .B2(keyinput214), .C1(n6264), .C2(keyinput255), .A(n8840), .ZN(n8844) );
  XNOR2_X1 U10378 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput130), .ZN(n8842) );
  XNOR2_X1 U10379 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput142), .ZN(n8841)
         );
  NAND2_X1 U10380 ( .A1(n8842), .A2(n8841), .ZN(n8843) );
  NOR4_X1 U10381 ( .A1(n8846), .A2(n8845), .A3(n8844), .A4(n8843), .ZN(n8847)
         );
  NAND4_X1 U10382 ( .A1(n8850), .A2(n8849), .A3(n8848), .A4(n8847), .ZN(n8851)
         );
  NOR4_X1 U10383 ( .A1(n8854), .A2(n8853), .A3(n8852), .A4(n8851), .ZN(n9036)
         );
  AOI22_X1 U10384 ( .A1(n8857), .A2(keyinput21), .B1(n8856), .B2(keyinput17), 
        .ZN(n8855) );
  OAI221_X1 U10385 ( .B1(n8857), .B2(keyinput21), .C1(n8856), .C2(keyinput17), 
        .A(n8855), .ZN(n8866) );
  AOI22_X1 U10386 ( .A1(n5083), .A2(keyinput106), .B1(keyinput19), .B2(n8859), 
        .ZN(n8858) );
  OAI221_X1 U10387 ( .B1(n5083), .B2(keyinput106), .C1(n8859), .C2(keyinput19), 
        .A(n8858), .ZN(n8865) );
  AOI22_X1 U10388 ( .A1(n5075), .A2(keyinput31), .B1(keyinput88), .B2(n5379), 
        .ZN(n8860) );
  OAI221_X1 U10389 ( .B1(n5075), .B2(keyinput31), .C1(n5379), .C2(keyinput88), 
        .A(n8860), .ZN(n8864) );
  AOI22_X1 U10390 ( .A1(n8862), .A2(keyinput37), .B1(keyinput68), .B2(n6808), 
        .ZN(n8861) );
  OAI221_X1 U10391 ( .B1(n8862), .B2(keyinput37), .C1(n6808), .C2(keyinput68), 
        .A(n8861), .ZN(n8863) );
  NOR4_X1 U10392 ( .A1(n8866), .A2(n8865), .A3(n8864), .A4(n8863), .ZN(n8907)
         );
  AOI22_X1 U10393 ( .A1(n7461), .A2(keyinput32), .B1(n5070), .B2(keyinput61), 
        .ZN(n8867) );
  OAI221_X1 U10394 ( .B1(n7461), .B2(keyinput32), .C1(n5070), .C2(keyinput61), 
        .A(n8867), .ZN(n8877) );
  AOI22_X1 U10395 ( .A1(n5089), .A2(keyinput13), .B1(keyinput26), .B2(n6804), 
        .ZN(n8868) );
  OAI221_X1 U10396 ( .B1(n5089), .B2(keyinput13), .C1(n6804), .C2(keyinput26), 
        .A(n8868), .ZN(n8876) );
  AOI22_X1 U10397 ( .A1(n8871), .A2(keyinput14), .B1(n8870), .B2(keyinput38), 
        .ZN(n8869) );
  OAI221_X1 U10398 ( .B1(n8871), .B2(keyinput14), .C1(n8870), .C2(keyinput38), 
        .A(n8869), .ZN(n8875) );
  INV_X1 U10399 ( .A(P1_D_REG_12__SCAN_IN), .ZN(n10189) );
  AOI22_X1 U10400 ( .A1(n10189), .A2(keyinput105), .B1(keyinput113), .B2(n8873), .ZN(n8872) );
  OAI221_X1 U10401 ( .B1(n10189), .B2(keyinput105), .C1(n8873), .C2(
        keyinput113), .A(n8872), .ZN(n8874) );
  NOR4_X1 U10402 ( .A1(n8877), .A2(n8876), .A3(n8875), .A4(n8874), .ZN(n8906)
         );
  INV_X1 U10403 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10391) );
  INV_X1 U10404 ( .A(P2_D_REG_8__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U10405 ( .A1(n10391), .A2(keyinput72), .B1(keyinput74), .B2(n10394), 
        .ZN(n8878) );
  OAI221_X1 U10406 ( .B1(n10391), .B2(keyinput72), .C1(n10394), .C2(keyinput74), .A(n8878), .ZN(n8889) );
  AOI22_X1 U10407 ( .A1(n6378), .A2(keyinput126), .B1(n8880), .B2(keyinput11), 
        .ZN(n8879) );
  OAI221_X1 U10408 ( .B1(n6378), .B2(keyinput126), .C1(n8880), .C2(keyinput11), 
        .A(n8879), .ZN(n8888) );
  AOI22_X1 U10409 ( .A1(n8883), .A2(keyinput29), .B1(keyinput16), .B2(n8882), 
        .ZN(n8881) );
  OAI221_X1 U10410 ( .B1(n8883), .B2(keyinput29), .C1(n8882), .C2(keyinput16), 
        .A(n8881), .ZN(n8887) );
  AOI22_X1 U10411 ( .A1(n8885), .A2(keyinput79), .B1(keyinput76), .B2(n5920), 
        .ZN(n8884) );
  OAI221_X1 U10412 ( .B1(n8885), .B2(keyinput79), .C1(n5920), .C2(keyinput76), 
        .A(n8884), .ZN(n8886) );
  NOR4_X1 U10413 ( .A1(n8889), .A2(n8888), .A3(n8887), .A4(n8886), .ZN(n8905)
         );
  INV_X1 U10414 ( .A(SI_4_), .ZN(n8891) );
  AOI22_X1 U10415 ( .A1(n5838), .A2(keyinput111), .B1(n8891), .B2(keyinput7), 
        .ZN(n8890) );
  OAI221_X1 U10416 ( .B1(n5838), .B2(keyinput111), .C1(n8891), .C2(keyinput7), 
        .A(n8890), .ZN(n8903) );
  AOI22_X1 U10417 ( .A1(n8894), .A2(keyinput123), .B1(n8893), .B2(keyinput47), 
        .ZN(n8892) );
  OAI221_X1 U10418 ( .B1(n8894), .B2(keyinput123), .C1(n8893), .C2(keyinput47), 
        .A(n8892), .ZN(n8902) );
  AOI22_X1 U10419 ( .A1(n8896), .A2(keyinput104), .B1(n5927), .B2(keyinput73), 
        .ZN(n8895) );
  OAI221_X1 U10420 ( .B1(n8896), .B2(keyinput104), .C1(n5927), .C2(keyinput73), 
        .A(n8895), .ZN(n8901) );
  AOI22_X1 U10421 ( .A1(n8899), .A2(keyinput117), .B1(n8898), .B2(keyinput109), 
        .ZN(n8897) );
  OAI221_X1 U10422 ( .B1(n8899), .B2(keyinput117), .C1(n8898), .C2(keyinput109), .A(n8897), .ZN(n8900) );
  NOR4_X1 U10423 ( .A1(n8903), .A2(n8902), .A3(n8901), .A4(n8900), .ZN(n8904)
         );
  NAND4_X1 U10424 ( .A1(n8907), .A2(n8906), .A3(n8905), .A4(n8904), .ZN(n9035)
         );
  AOI22_X1 U10425 ( .A1(n8909), .A2(keyinput48), .B1(keyinput22), .B2(n5127), 
        .ZN(n8908) );
  OAI221_X1 U10426 ( .B1(n8909), .B2(keyinput48), .C1(n5127), .C2(keyinput22), 
        .A(n8908), .ZN(n8919) );
  AOI22_X1 U10427 ( .A1(n8911), .A2(keyinput93), .B1(keyinput71), .B2(n5643), 
        .ZN(n8910) );
  OAI221_X1 U10428 ( .B1(n8911), .B2(keyinput93), .C1(n5643), .C2(keyinput71), 
        .A(n8910), .ZN(n8918) );
  AOI22_X1 U10429 ( .A1(n10386), .A2(keyinput99), .B1(n8913), .B2(keyinput116), 
        .ZN(n8912) );
  OAI221_X1 U10430 ( .B1(n10386), .B2(keyinput99), .C1(n8913), .C2(keyinput116), .A(n8912), .ZN(n8917) );
  AOI22_X1 U10431 ( .A1(n8915), .A2(keyinput96), .B1(n10188), .B2(keyinput92), 
        .ZN(n8914) );
  OAI221_X1 U10432 ( .B1(n8915), .B2(keyinput96), .C1(n10188), .C2(keyinput92), 
        .A(n8914), .ZN(n8916) );
  OR4_X1 U10433 ( .A1(n8919), .A2(n8918), .A3(n8917), .A4(n8916), .ZN(n9034)
         );
  AOI22_X1 U10434 ( .A1(n9374), .A2(keyinput50), .B1(n6141), .B2(keyinput49), 
        .ZN(n8920) );
  OAI221_X1 U10435 ( .B1(n9374), .B2(keyinput50), .C1(n6141), .C2(keyinput49), 
        .A(n8920), .ZN(n8928) );
  AOI22_X1 U10436 ( .A1(n8923), .A2(keyinput30), .B1(n8922), .B2(keyinput53), 
        .ZN(n8921) );
  OAI221_X1 U10437 ( .B1(n8923), .B2(keyinput30), .C1(n8922), .C2(keyinput53), 
        .A(n8921), .ZN(n8927) );
  XOR2_X1 U10438 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput8), .Z(n8926) );
  XNOR2_X1 U10439 ( .A(n8924), .B(keyinput108), .ZN(n8925) );
  NOR4_X1 U10440 ( .A1(n8928), .A2(n8927), .A3(n8926), .A4(n8925), .ZN(n8958)
         );
  INV_X1 U10441 ( .A(P1_D_REG_4__SCAN_IN), .ZN(n10190) );
  INV_X1 U10442 ( .A(P2_D_REG_17__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U10443 ( .A1(n10190), .A2(keyinput59), .B1(keyinput24), .B2(n10390), 
        .ZN(n8929) );
  OAI221_X1 U10444 ( .B1(n10190), .B2(keyinput59), .C1(n10390), .C2(keyinput24), .A(n8929), .ZN(n8937) );
  AOI22_X1 U10445 ( .A1(n8931), .A2(keyinput4), .B1(keyinput94), .B2(n9226), 
        .ZN(n8930) );
  OAI221_X1 U10446 ( .B1(n8931), .B2(keyinput4), .C1(n9226), .C2(keyinput94), 
        .A(n8930), .ZN(n8936) );
  AOI22_X1 U10447 ( .A1(n8934), .A2(keyinput20), .B1(n8933), .B2(keyinput85), 
        .ZN(n8932) );
  OAI221_X1 U10448 ( .B1(n8934), .B2(keyinput20), .C1(n8933), .C2(keyinput85), 
        .A(n8932), .ZN(n8935) );
  NOR3_X1 U10449 ( .A1(n8937), .A2(n8936), .A3(n8935), .ZN(n8957) );
  OAI22_X1 U10450 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(keyinput3), .B1(
        P2_REG3_REG_6__SCAN_IN), .B2(keyinput5), .ZN(n8938) );
  AOI221_X1 U10451 ( .B1(P2_IR_REG_9__SCAN_IN), .B2(keyinput3), .C1(keyinput5), 
        .C2(P2_REG3_REG_6__SCAN_IN), .A(n8938), .ZN(n8945) );
  OAI22_X1 U10452 ( .A1(P1_REG1_REG_22__SCAN_IN), .A2(keyinput122), .B1(
        P1_ADDR_REG_7__SCAN_IN), .B2(keyinput81), .ZN(n8939) );
  AOI221_X1 U10453 ( .B1(P1_REG1_REG_22__SCAN_IN), .B2(keyinput122), .C1(
        keyinput81), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n8939), .ZN(n8944) );
  OAI22_X1 U10454 ( .A1(P1_REG0_REG_11__SCAN_IN), .A2(keyinput77), .B1(
        P1_REG2_REG_8__SCAN_IN), .B2(keyinput55), .ZN(n8940) );
  AOI221_X1 U10455 ( .B1(P1_REG0_REG_11__SCAN_IN), .B2(keyinput77), .C1(
        keyinput55), .C2(P1_REG2_REG_8__SCAN_IN), .A(n8940), .ZN(n8943) );
  OAI22_X1 U10456 ( .A1(P2_REG0_REG_5__SCAN_IN), .A2(keyinput119), .B1(
        P2_ADDR_REG_2__SCAN_IN), .B2(keyinput9), .ZN(n8941) );
  AOI221_X1 U10457 ( .B1(P2_REG0_REG_5__SCAN_IN), .B2(keyinput119), .C1(
        keyinput9), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n8941), .ZN(n8942) );
  NAND4_X1 U10458 ( .A1(n8945), .A2(n8944), .A3(n8943), .A4(n8942), .ZN(n8955)
         );
  OAI22_X1 U10459 ( .A1(P1_STATE_REG_SCAN_IN), .A2(keyinput82), .B1(
        P1_REG1_REG_2__SCAN_IN), .B2(keyinput97), .ZN(n8946) );
  AOI221_X1 U10460 ( .B1(P1_STATE_REG_SCAN_IN), .B2(keyinput82), .C1(
        keyinput97), .C2(P1_REG1_REG_2__SCAN_IN), .A(n8946), .ZN(n8953) );
  OAI22_X1 U10461 ( .A1(P1_REG3_REG_28__SCAN_IN), .A2(keyinput10), .B1(
        keyinput86), .B2(P1_REG2_REG_6__SCAN_IN), .ZN(n8947) );
  AOI221_X1 U10462 ( .B1(P1_REG3_REG_28__SCAN_IN), .B2(keyinput10), .C1(
        P1_REG2_REG_6__SCAN_IN), .C2(keyinput86), .A(n8947), .ZN(n8952) );
  OAI22_X1 U10463 ( .A1(P2_D_REG_10__SCAN_IN), .A2(keyinput39), .B1(keyinput52), .B2(P2_REG1_REG_13__SCAN_IN), .ZN(n8948) );
  AOI221_X1 U10464 ( .B1(P2_D_REG_10__SCAN_IN), .B2(keyinput39), .C1(
        P2_REG1_REG_13__SCAN_IN), .C2(keyinput52), .A(n8948), .ZN(n8951) );
  OAI22_X1 U10465 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(keyinput110), .B1(
        P1_REG2_REG_7__SCAN_IN), .B2(keyinput118), .ZN(n8949) );
  AOI221_X1 U10466 ( .B1(P1_REG1_REG_16__SCAN_IN), .B2(keyinput110), .C1(
        keyinput118), .C2(P1_REG2_REG_7__SCAN_IN), .A(n8949), .ZN(n8950) );
  NAND4_X1 U10467 ( .A1(n8953), .A2(n8952), .A3(n8951), .A4(n8950), .ZN(n8954)
         );
  NOR2_X1 U10468 ( .A1(n8955), .A2(n8954), .ZN(n8956) );
  NAND3_X1 U10469 ( .A1(n8958), .A2(n8957), .A3(n8956), .ZN(n8997) );
  OAI22_X1 U10470 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(keyinput40), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(keyinput120), .ZN(n8959) );
  AOI221_X1 U10471 ( .B1(P1_IR_REG_19__SCAN_IN), .B2(keyinput40), .C1(
        keyinput120), .C2(P1_DATAO_REG_20__SCAN_IN), .A(n8959), .ZN(n8966) );
  OAI22_X1 U10472 ( .A1(P1_D_REG_3__SCAN_IN), .A2(keyinput100), .B1(
        P1_D_REG_23__SCAN_IN), .B2(keyinput67), .ZN(n8960) );
  AOI221_X1 U10473 ( .B1(P1_D_REG_3__SCAN_IN), .B2(keyinput100), .C1(
        keyinput67), .C2(P1_D_REG_23__SCAN_IN), .A(n8960), .ZN(n8965) );
  OAI22_X1 U10474 ( .A1(P1_D_REG_16__SCAN_IN), .A2(keyinput44), .B1(
        P2_REG3_REG_25__SCAN_IN), .B2(keyinput101), .ZN(n8961) );
  AOI221_X1 U10475 ( .B1(P1_D_REG_16__SCAN_IN), .B2(keyinput44), .C1(
        keyinput101), .C2(P2_REG3_REG_25__SCAN_IN), .A(n8961), .ZN(n8964) );
  OAI22_X1 U10476 ( .A1(SI_23_), .A2(keyinput90), .B1(keyinput121), .B2(
        P2_D_REG_27__SCAN_IN), .ZN(n8962) );
  AOI221_X1 U10477 ( .B1(SI_23_), .B2(keyinput90), .C1(P2_D_REG_27__SCAN_IN), 
        .C2(keyinput121), .A(n8962), .ZN(n8963) );
  NAND4_X1 U10478 ( .A1(n8966), .A2(n8965), .A3(n8964), .A4(n8963), .ZN(n8996)
         );
  OAI22_X1 U10479 ( .A1(P1_REG3_REG_16__SCAN_IN), .A2(keyinput28), .B1(
        P2_REG0_REG_10__SCAN_IN), .B2(keyinput6), .ZN(n8967) );
  AOI221_X1 U10480 ( .B1(P1_REG3_REG_16__SCAN_IN), .B2(keyinput28), .C1(
        keyinput6), .C2(P2_REG0_REG_10__SCAN_IN), .A(n8967), .ZN(n8974) );
  OAI22_X1 U10481 ( .A1(P2_REG0_REG_8__SCAN_IN), .A2(keyinput112), .B1(
        P1_REG0_REG_31__SCAN_IN), .B2(keyinput15), .ZN(n8968) );
  AOI221_X1 U10482 ( .B1(P2_REG0_REG_8__SCAN_IN), .B2(keyinput112), .C1(
        keyinput15), .C2(P1_REG0_REG_31__SCAN_IN), .A(n8968), .ZN(n8973) );
  OAI22_X1 U10483 ( .A1(P2_D_REG_30__SCAN_IN), .A2(keyinput46), .B1(
        keyinput102), .B2(P2_REG3_REG_20__SCAN_IN), .ZN(n8969) );
  AOI221_X1 U10484 ( .B1(P2_D_REG_30__SCAN_IN), .B2(keyinput46), .C1(
        P2_REG3_REG_20__SCAN_IN), .C2(keyinput102), .A(n8969), .ZN(n8972) );
  OAI22_X1 U10485 ( .A1(P1_IR_REG_29__SCAN_IN), .A2(keyinput60), .B1(
        P2_REG1_REG_5__SCAN_IN), .B2(keyinput84), .ZN(n8970) );
  AOI221_X1 U10486 ( .B1(P1_IR_REG_29__SCAN_IN), .B2(keyinput60), .C1(
        keyinput84), .C2(P2_REG1_REG_5__SCAN_IN), .A(n8970), .ZN(n8971) );
  NAND4_X1 U10487 ( .A1(n8974), .A2(n8973), .A3(n8972), .A4(n8971), .ZN(n8995)
         );
  OAI22_X1 U10488 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput127), .B1(
        keyinput124), .B2(P1_REG3_REG_9__SCAN_IN), .ZN(n8975) );
  AOI221_X1 U10489 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput127), .C1(
        P1_REG3_REG_9__SCAN_IN), .C2(keyinput124), .A(n8975), .ZN(n8982) );
  OAI22_X1 U10490 ( .A1(SI_26_), .A2(keyinput65), .B1(P2_D_REG_1__SCAN_IN), 
        .B2(keyinput35), .ZN(n8976) );
  AOI221_X1 U10491 ( .B1(SI_26_), .B2(keyinput65), .C1(keyinput35), .C2(
        P2_D_REG_1__SCAN_IN), .A(n8976), .ZN(n8981) );
  OAI22_X1 U10492 ( .A1(SI_31_), .A2(keyinput66), .B1(keyinput107), .B2(
        P1_ADDR_REG_4__SCAN_IN), .ZN(n8977) );
  AOI221_X1 U10493 ( .B1(SI_31_), .B2(keyinput66), .C1(P1_ADDR_REG_4__SCAN_IN), 
        .C2(keyinput107), .A(n8977), .ZN(n8980) );
  OAI22_X1 U10494 ( .A1(P2_D_REG_13__SCAN_IN), .A2(keyinput62), .B1(
        P2_ADDR_REG_6__SCAN_IN), .B2(keyinput51), .ZN(n8978) );
  AOI221_X1 U10495 ( .B1(P2_D_REG_13__SCAN_IN), .B2(keyinput62), .C1(
        keyinput51), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n8978), .ZN(n8979) );
  NAND4_X1 U10496 ( .A1(n8982), .A2(n8981), .A3(n8980), .A4(n8979), .ZN(n8993)
         );
  AOI22_X1 U10497 ( .A1(n7384), .A2(keyinput43), .B1(keyinput33), .B2(n7001), 
        .ZN(n8983) );
  OAI221_X1 U10498 ( .B1(n7384), .B2(keyinput43), .C1(n7001), .C2(keyinput33), 
        .A(n8983), .ZN(n8992) );
  AOI22_X1 U10499 ( .A1(n5073), .A2(keyinput25), .B1(keyinput80), .B2(n8985), 
        .ZN(n8984) );
  OAI221_X1 U10500 ( .B1(n5073), .B2(keyinput25), .C1(n8985), .C2(keyinput80), 
        .A(n8984), .ZN(n8991) );
  XNOR2_X1 U10501 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput87), .ZN(n8989)
         );
  XNOR2_X1 U10502 ( .A(SI_1_), .B(keyinput12), .ZN(n8988) );
  XNOR2_X1 U10503 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput2), .ZN(n8987) );
  XNOR2_X1 U10504 ( .A(P1_REG2_REG_1__SCAN_IN), .B(keyinput34), .ZN(n8986) );
  NAND4_X1 U10505 ( .A1(n8989), .A2(n8988), .A3(n8987), .A4(n8986), .ZN(n8990)
         );
  OR4_X1 U10506 ( .A1(n8993), .A2(n8992), .A3(n8991), .A4(n8990), .ZN(n8994)
         );
  NOR4_X1 U10507 ( .A1(n8997), .A2(n8996), .A3(n8995), .A4(n8994), .ZN(n9032)
         );
  OAI22_X1 U10508 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(keyinput69), .B1(keyinput89), .B2(P2_REG0_REG_9__SCAN_IN), .ZN(n8998) );
  AOI221_X1 U10509 ( .B1(P1_IR_REG_2__SCAN_IN), .B2(keyinput69), .C1(
        P2_REG0_REG_9__SCAN_IN), .C2(keyinput89), .A(n8998), .ZN(n9005) );
  OAI22_X1 U10510 ( .A1(P2_DATAO_REG_9__SCAN_IN), .A2(keyinput125), .B1(
        keyinput95), .B2(P1_REG2_REG_10__SCAN_IN), .ZN(n8999) );
  AOI221_X1 U10511 ( .B1(P2_DATAO_REG_9__SCAN_IN), .B2(keyinput125), .C1(
        P1_REG2_REG_10__SCAN_IN), .C2(keyinput95), .A(n8999), .ZN(n9004) );
  OAI22_X1 U10512 ( .A1(P1_REG2_REG_12__SCAN_IN), .A2(keyinput0), .B1(
        keyinput56), .B2(P2_REG2_REG_8__SCAN_IN), .ZN(n9000) );
  AOI221_X1 U10513 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(keyinput0), .C1(
        P2_REG2_REG_8__SCAN_IN), .C2(keyinput56), .A(n9000), .ZN(n9003) );
  OAI22_X1 U10514 ( .A1(P1_B_REG_SCAN_IN), .A2(keyinput75), .B1(keyinput45), 
        .B2(P1_REG3_REG_10__SCAN_IN), .ZN(n9001) );
  AOI221_X1 U10515 ( .B1(P1_B_REG_SCAN_IN), .B2(keyinput75), .C1(
        P1_REG3_REG_10__SCAN_IN), .C2(keyinput45), .A(n9001), .ZN(n9002) );
  NAND4_X1 U10516 ( .A1(n9005), .A2(n9004), .A3(n9003), .A4(n9002), .ZN(n9015)
         );
  OAI22_X1 U10517 ( .A1(P1_REG1_REG_12__SCAN_IN), .A2(keyinput54), .B1(
        P2_D_REG_23__SCAN_IN), .B2(keyinput70), .ZN(n9006) );
  AOI221_X1 U10518 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(keyinput54), .C1(
        keyinput70), .C2(P2_D_REG_23__SCAN_IN), .A(n9006), .ZN(n9013) );
  OAI22_X1 U10519 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(keyinput42), .B1(
        keyinput18), .B2(P2_REG2_REG_23__SCAN_IN), .ZN(n9007) );
  AOI221_X1 U10520 ( .B1(P1_DATAO_REG_4__SCAN_IN), .B2(keyinput42), .C1(
        P2_REG2_REG_23__SCAN_IN), .C2(keyinput18), .A(n9007), .ZN(n9012) );
  OAI22_X1 U10521 ( .A1(P1_REG2_REG_27__SCAN_IN), .A2(keyinput83), .B1(
        keyinput27), .B2(P1_ADDR_REG_9__SCAN_IN), .ZN(n9008) );
  AOI221_X1 U10522 ( .B1(P1_REG2_REG_27__SCAN_IN), .B2(keyinput83), .C1(
        P1_ADDR_REG_9__SCAN_IN), .C2(keyinput27), .A(n9008), .ZN(n9011) );
  OAI22_X1 U10523 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(keyinput98), .B1(
        keyinput57), .B2(P1_REG0_REG_16__SCAN_IN), .ZN(n9009) );
  AOI221_X1 U10524 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(keyinput98), .C1(
        P1_REG0_REG_16__SCAN_IN), .C2(keyinput57), .A(n9009), .ZN(n9010) );
  NAND4_X1 U10525 ( .A1(n9013), .A2(n9012), .A3(n9011), .A4(n9010), .ZN(n9014)
         );
  NOR2_X1 U10526 ( .A1(n9015), .A2(n9014), .ZN(n9031) );
  AOI22_X1 U10527 ( .A1(n9932), .A2(keyinput23), .B1(n9550), .B2(keyinput91), 
        .ZN(n9016) );
  OAI221_X1 U10528 ( .B1(n9932), .B2(keyinput23), .C1(n9550), .C2(keyinput91), 
        .A(n9016), .ZN(n9020) );
  INV_X1 U10529 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n10186) );
  XNOR2_X1 U10530 ( .A(n10186), .B(keyinput36), .ZN(n9019) );
  INV_X1 U10531 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9017) );
  XNOR2_X1 U10532 ( .A(n9017), .B(keyinput114), .ZN(n9018) );
  NOR3_X1 U10533 ( .A1(n9020), .A2(n9019), .A3(n9018), .ZN(n9030) );
  OAI22_X1 U10534 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(keyinput115), .B1(
        keyinput63), .B2(P1_REG2_REG_5__SCAN_IN), .ZN(n9021) );
  AOI221_X1 U10535 ( .B1(P1_REG1_REG_7__SCAN_IN), .B2(keyinput115), .C1(
        P1_REG2_REG_5__SCAN_IN), .C2(keyinput63), .A(n9021), .ZN(n9028) );
  OAI22_X1 U10536 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput103), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(keyinput58), .ZN(n9022) );
  AOI221_X1 U10537 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput103), .C1(
        keyinput58), .C2(P2_DATAO_REG_30__SCAN_IN), .A(n9022), .ZN(n9027) );
  OAI22_X1 U10538 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput1), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(keyinput78), .ZN(n9023) );
  AOI221_X1 U10539 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput1), .C1(
        keyinput78), .C2(P1_DATAO_REG_7__SCAN_IN), .A(n9023), .ZN(n9026) );
  OAI22_X1 U10540 ( .A1(P1_REG1_REG_27__SCAN_IN), .A2(keyinput41), .B1(
        keyinput64), .B2(P2_REG3_REG_27__SCAN_IN), .ZN(n9024) );
  AOI221_X1 U10541 ( .B1(P1_REG1_REG_27__SCAN_IN), .B2(keyinput41), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput64), .A(n9024), .ZN(n9025) );
  AND4_X1 U10542 ( .A1(n9028), .A2(n9027), .A3(n9026), .A4(n9025), .ZN(n9029)
         );
  NAND4_X1 U10543 ( .A1(n9032), .A2(n9031), .A3(n9030), .A4(n9029), .ZN(n9033)
         );
  NOR4_X1 U10544 ( .A1(n9036), .A2(n9035), .A3(n9034), .A4(n9033), .ZN(n9054)
         );
  XNOR2_X1 U10545 ( .A(n9039), .B(n9038), .ZN(n9044) );
  NAND2_X1 U10546 ( .A1(n9040), .A2(n10368), .ZN(n9042) );
  NAND2_X1 U10547 ( .A1(n9083), .A2(n10366), .ZN(n9041) );
  AOI21_X1 U10548 ( .B1(n9280), .B2(n9058), .A(n9045), .ZN(n9281) );
  INV_X1 U10549 ( .A(n9281), .ZN(n9046) );
  INV_X1 U10550 ( .A(n9047), .ZN(n9048) );
  AOI22_X1 U10551 ( .A1(n9048), .A2(n10373), .B1(P2_REG2_REG_28__SCAN_IN), 
        .B2(n10372), .ZN(n9049) );
  OAI21_X1 U10552 ( .B1(n8347), .B2(n9254), .A(n9049), .ZN(n9050) );
  INV_X1 U10553 ( .A(n9050), .ZN(n9051) );
  XOR2_X1 U10554 ( .A(n9054), .B(n9053), .Z(P2_U3268) );
  OAI21_X1 U10555 ( .B1(n9056), .B2(n9064), .A(n9055), .ZN(n9057) );
  INV_X1 U10556 ( .A(n9057), .ZN(n9289) );
  INV_X1 U10557 ( .A(n9058), .ZN(n9059) );
  AOI21_X1 U10558 ( .B1(n9285), .B2(n9075), .A(n9059), .ZN(n9286) );
  AOI22_X1 U10559 ( .A1(n9060), .A2(n10373), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n10372), .ZN(n9061) );
  OAI21_X1 U10560 ( .B1(n9062), .B2(n9254), .A(n9061), .ZN(n9069) );
  XOR2_X1 U10561 ( .A(n9064), .B(n9063), .Z(n9067) );
  AOI222_X1 U10562 ( .A1(n10371), .A2(n9067), .B1(n9066), .B2(n10366), .C1(
        n9065), .C2(n10368), .ZN(n9288) );
  NOR2_X1 U10563 ( .A1(n9288), .A2(n10372), .ZN(n9068) );
  AOI211_X1 U10564 ( .C1(n9286), .C2(n9262), .A(n9069), .B(n9068), .ZN(n9070)
         );
  OAI21_X1 U10565 ( .B1(n9233), .B2(n9289), .A(n9070), .ZN(P2_U3269) );
  OAI21_X1 U10566 ( .B1(n9073), .B2(n9072), .A(n9071), .ZN(n9074) );
  INV_X1 U10567 ( .A(n9074), .ZN(n9294) );
  AOI211_X1 U10568 ( .C1(n9291), .C2(n9091), .A(n10455), .B(n4735), .ZN(n9290)
         );
  INV_X1 U10569 ( .A(n9076), .ZN(n9077) );
  AOI22_X1 U10570 ( .A1(n9077), .A2(n10373), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n10372), .ZN(n9078) );
  OAI21_X1 U10571 ( .B1(n9079), .B2(n9254), .A(n9078), .ZN(n9086) );
  OAI21_X1 U10572 ( .B1(n9082), .B2(n9081), .A(n9080), .ZN(n9084) );
  AOI222_X1 U10573 ( .A1(n10371), .A2(n9084), .B1(n9083), .B2(n10368), .C1(
        n9114), .C2(n10366), .ZN(n9293) );
  NOR2_X1 U10574 ( .A1(n9293), .A2(n10372), .ZN(n9085) );
  AOI211_X1 U10575 ( .C1(n9290), .C2(n9230), .A(n9086), .B(n9085), .ZN(n9087)
         );
  OAI21_X1 U10576 ( .B1(n9233), .B2(n9294), .A(n9087), .ZN(P2_U3270) );
  OAI21_X1 U10577 ( .B1(n9089), .B2(n9098), .A(n9088), .ZN(n9090) );
  INV_X1 U10578 ( .A(n9090), .ZN(n9299) );
  INV_X1 U10579 ( .A(n9105), .ZN(n9093) );
  INV_X1 U10580 ( .A(n9091), .ZN(n9092) );
  AOI211_X1 U10581 ( .C1(n9296), .C2(n9093), .A(n10455), .B(n9092), .ZN(n9295)
         );
  INV_X1 U10582 ( .A(n9094), .ZN(n9095) );
  AOI22_X1 U10583 ( .A1(n9095), .A2(n10373), .B1(P2_REG2_REG_25__SCAN_IN), 
        .B2(n10372), .ZN(n9096) );
  OAI21_X1 U10584 ( .B1(n8449), .B2(n9254), .A(n9096), .ZN(n9102) );
  XNOR2_X1 U10585 ( .A(n9097), .B(n9098), .ZN(n9100) );
  AOI21_X1 U10586 ( .B1(n9100), .B2(n10371), .A(n9099), .ZN(n9298) );
  NOR2_X1 U10587 ( .A1(n9298), .A2(n10372), .ZN(n9101) );
  AOI211_X1 U10588 ( .C1(n9230), .C2(n9295), .A(n9102), .B(n9101), .ZN(n9103)
         );
  OAI21_X1 U10589 ( .B1(n9233), .B2(n9299), .A(n9103), .ZN(P2_U3271) );
  XOR2_X1 U10590 ( .A(n9112), .B(n9104), .Z(n9304) );
  AOI21_X1 U10591 ( .B1(n9300), .B2(n9122), .A(n9105), .ZN(n9301) );
  AOI22_X1 U10592 ( .A1(P2_REG2_REG_24__SCAN_IN), .A2(n10372), .B1(n9106), 
        .B2(n10373), .ZN(n9107) );
  OAI21_X1 U10593 ( .B1(n9108), .B2(n9254), .A(n9107), .ZN(n9117) );
  INV_X1 U10594 ( .A(n9109), .ZN(n9110) );
  NOR2_X1 U10595 ( .A1(n4514), .A2(n9110), .ZN(n9111) );
  XOR2_X1 U10596 ( .A(n9112), .B(n9111), .Z(n9115) );
  AOI222_X1 U10597 ( .A1(n10371), .A2(n9115), .B1(n9114), .B2(n10368), .C1(
        n9113), .C2(n10366), .ZN(n9303) );
  NOR2_X1 U10598 ( .A1(n9303), .A2(n10372), .ZN(n9116) );
  AOI211_X1 U10599 ( .C1(n9301), .C2(n9262), .A(n9117), .B(n9116), .ZN(n9118)
         );
  OAI21_X1 U10600 ( .B1(n9233), .B2(n9304), .A(n9118), .ZN(P2_U3272) );
  OAI21_X1 U10601 ( .B1(n9121), .B2(n9120), .A(n9119), .ZN(n9309) );
  INV_X1 U10602 ( .A(n9137), .ZN(n9124) );
  INV_X1 U10603 ( .A(n9122), .ZN(n9123) );
  AOI21_X1 U10604 ( .B1(n9305), .B2(n9124), .A(n9123), .ZN(n9306) );
  INV_X1 U10605 ( .A(n9125), .ZN(n9126) );
  AOI22_X1 U10606 ( .A1(n10372), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9126), 
        .B2(n10373), .ZN(n9127) );
  OAI21_X1 U10607 ( .B1(n9128), .B2(n9254), .A(n9127), .ZN(n9134) );
  INV_X1 U10608 ( .A(n4514), .ZN(n9129) );
  OAI21_X1 U10609 ( .B1(n9130), .B2(n4546), .A(n9129), .ZN(n9132) );
  AOI222_X1 U10610 ( .A1(n10371), .A2(n9132), .B1(n8444), .B2(n10366), .C1(
        n9131), .C2(n10368), .ZN(n9308) );
  NOR2_X1 U10611 ( .A1(n9308), .A2(n10372), .ZN(n9133) );
  AOI211_X1 U10612 ( .C1(n9306), .C2(n9262), .A(n9134), .B(n9133), .ZN(n9135)
         );
  OAI21_X1 U10613 ( .B1(n9233), .B2(n9309), .A(n9135), .ZN(P2_U3273) );
  XNOR2_X1 U10614 ( .A(n9136), .B(n9143), .ZN(n9314) );
  AOI21_X1 U10615 ( .B1(n9310), .B2(n4729), .A(n9137), .ZN(n9311) );
  INV_X1 U10616 ( .A(n9138), .ZN(n9139) );
  AOI22_X1 U10617 ( .A1(n10372), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9139), 
        .B2(n10373), .ZN(n9140) );
  OAI21_X1 U10618 ( .B1(n9141), .B2(n9254), .A(n9140), .ZN(n9150) );
  INV_X1 U10619 ( .A(n9142), .ZN(n9146) );
  AOI21_X1 U10620 ( .B1(n9158), .B2(n9144), .A(n9143), .ZN(n9145) );
  NOR3_X1 U10621 ( .A1(n9146), .A2(n9145), .A3(n9246), .ZN(n9148) );
  NOR2_X1 U10622 ( .A1(n9148), .A2(n9147), .ZN(n9313) );
  NOR2_X1 U10623 ( .A1(n9313), .A2(n10372), .ZN(n9149) );
  AOI211_X1 U10624 ( .C1(n9311), .C2(n9262), .A(n9150), .B(n9149), .ZN(n9151)
         );
  OAI21_X1 U10625 ( .B1(n9233), .B2(n9314), .A(n9151), .ZN(P2_U3274) );
  XNOR2_X1 U10626 ( .A(n9152), .B(n9153), .ZN(n9319) );
  AOI21_X1 U10627 ( .B1(n9315), .B2(n9166), .A(n9154), .ZN(n9316) );
  AOI22_X1 U10628 ( .A1(n10372), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9155), 
        .B2(n10373), .ZN(n9156) );
  OAI21_X1 U10629 ( .B1(n9157), .B2(n9254), .A(n9156), .ZN(n9163) );
  OAI21_X1 U10630 ( .B1(n9160), .B2(n9159), .A(n9158), .ZN(n9161) );
  AOI222_X1 U10631 ( .A1(n10371), .A2(n9161), .B1(n8444), .B2(n10368), .C1(
        n9186), .C2(n10366), .ZN(n9318) );
  NOR2_X1 U10632 ( .A1(n9318), .A2(n10372), .ZN(n9162) );
  AOI211_X1 U10633 ( .C1(n9316), .C2(n9262), .A(n9163), .B(n9162), .ZN(n9164)
         );
  OAI21_X1 U10634 ( .B1(n9233), .B2(n9319), .A(n9164), .ZN(P2_U3275) );
  XNOR2_X1 U10635 ( .A(n9165), .B(n9174), .ZN(n9324) );
  INV_X1 U10636 ( .A(n9166), .ZN(n9167) );
  AOI211_X1 U10637 ( .C1(n9321), .C2(n9168), .A(n10455), .B(n9167), .ZN(n9320)
         );
  AOI22_X1 U10638 ( .A1(n10372), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n9169), 
        .B2(n10373), .ZN(n9170) );
  OAI21_X1 U10639 ( .B1(n9171), .B2(n9254), .A(n9170), .ZN(n9178) );
  OAI21_X1 U10640 ( .B1(n9174), .B2(n9173), .A(n9172), .ZN(n9176) );
  AOI222_X1 U10641 ( .A1(n10371), .A2(n9176), .B1(n9210), .B2(n10366), .C1(
        n9175), .C2(n10368), .ZN(n9323) );
  NOR2_X1 U10642 ( .A1(n9323), .A2(n10372), .ZN(n9177) );
  AOI211_X1 U10643 ( .C1(n9320), .C2(n9179), .A(n9178), .B(n9177), .ZN(n9180)
         );
  OAI21_X1 U10644 ( .B1(n9233), .B2(n9324), .A(n9180), .ZN(P2_U3276) );
  INV_X1 U10645 ( .A(n9185), .ZN(n9181) );
  XNOR2_X1 U10646 ( .A(n9182), .B(n9181), .ZN(n9328) );
  OAI21_X1 U10647 ( .B1(n9185), .B2(n9184), .A(n9183), .ZN(n9187) );
  AOI222_X1 U10648 ( .A1(n10371), .A2(n9187), .B1(n9186), .B2(n10368), .C1(
        n9218), .C2(n10366), .ZN(n9193) );
  INV_X1 U10649 ( .A(n9328), .ZN(n9190) );
  XNOR2_X1 U10650 ( .A(n9203), .B(n9188), .ZN(n9189) );
  OAI21_X1 U10651 ( .B1(n10455), .B2(n9189), .A(n9193), .ZN(n9325) );
  AOI21_X1 U10652 ( .B1(n9191), .B2(n9190), .A(n9325), .ZN(n9192) );
  AOI211_X1 U10653 ( .C1(n9194), .C2(n9193), .A(n10372), .B(n9192), .ZN(n9195)
         );
  INV_X1 U10654 ( .A(n9195), .ZN(n9201) );
  INV_X1 U10655 ( .A(n9196), .ZN(n9197) );
  OAI22_X1 U10656 ( .A1(n9259), .A2(n9198), .B1(n9197), .B2(n9256), .ZN(n9199)
         );
  AOI21_X1 U10657 ( .B1(n9326), .B2(n10355), .A(n9199), .ZN(n9200) );
  OAI211_X1 U10658 ( .C1(n9328), .C2(n10360), .A(n9201), .B(n9200), .ZN(
        P2_U3277) );
  XNOR2_X1 U10659 ( .A(n9202), .B(n9208), .ZN(n9333) );
  AOI21_X1 U10660 ( .B1(n9329), .B2(n9228), .A(n9203), .ZN(n9330) );
  AOI22_X1 U10661 ( .A1(n10372), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9204), 
        .B2(n10373), .ZN(n9205) );
  OAI21_X1 U10662 ( .B1(n9206), .B2(n9254), .A(n9205), .ZN(n9213) );
  XOR2_X1 U10663 ( .A(n9208), .B(n9207), .Z(n9211) );
  AOI222_X1 U10664 ( .A1(n10371), .A2(n9211), .B1(n9210), .B2(n10368), .C1(
        n9209), .C2(n10366), .ZN(n9332) );
  NOR2_X1 U10665 ( .A1(n9332), .A2(n10372), .ZN(n9212) );
  AOI211_X1 U10666 ( .C1(n9330), .C2(n9262), .A(n9213), .B(n9212), .ZN(n9214)
         );
  OAI21_X1 U10667 ( .B1(n9233), .B2(n9333), .A(n9214), .ZN(P2_U3278) );
  INV_X1 U10668 ( .A(n9215), .ZN(n9216) );
  NOR2_X1 U10669 ( .A1(n4526), .A2(n9216), .ZN(n9217) );
  XNOR2_X1 U10670 ( .A(n9217), .B(n9222), .ZN(n9220) );
  AOI222_X1 U10671 ( .A1(n10371), .A2(n9220), .B1(n9219), .B2(n10366), .C1(
        n9218), .C2(n10368), .ZN(n9337) );
  OAI21_X1 U10672 ( .B1(n9223), .B2(n9222), .A(n9221), .ZN(n9224) );
  INV_X1 U10673 ( .A(n9224), .ZN(n9338) );
  OAI22_X1 U10674 ( .A1(n9259), .A2(n9226), .B1(n9225), .B2(n9256), .ZN(n9227)
         );
  AOI21_X1 U10675 ( .B1(n9335), .B2(n10355), .A(n9227), .ZN(n9232) );
  AOI21_X1 U10676 ( .B1(n9252), .B2(n9335), .A(n10455), .ZN(n9229) );
  AND2_X1 U10677 ( .A1(n9229), .A2(n9228), .ZN(n9334) );
  NAND2_X1 U10678 ( .A1(n9334), .A2(n9230), .ZN(n9231) );
  OAI211_X1 U10679 ( .C1(n9338), .C2(n9233), .A(n9232), .B(n9231), .ZN(n9234)
         );
  INV_X1 U10680 ( .A(n9234), .ZN(n9235) );
  OAI21_X1 U10681 ( .B1(n9337), .B2(n10372), .A(n9235), .ZN(P2_U3279) );
  NAND2_X1 U10682 ( .A1(n9238), .A2(n9237), .ZN(n9239) );
  OAI22_X1 U10683 ( .A1(n9243), .A2(n9242), .B1(n9241), .B2(n9240), .ZN(n9249)
         );
  AOI21_X1 U10684 ( .B1(n9245), .B2(n9244), .A(n4526), .ZN(n9247) );
  NOR2_X1 U10685 ( .A1(n9247), .A2(n9246), .ZN(n9248) );
  AOI211_X1 U10686 ( .C1(n9339), .C2(n9250), .A(n9249), .B(n9248), .ZN(n9343)
         );
  INV_X1 U10687 ( .A(n9252), .ZN(n9253) );
  AOI21_X1 U10688 ( .B1(n9340), .B2(n4723), .A(n9253), .ZN(n9341) );
  NOR2_X1 U10689 ( .A1(n9255), .A2(n9254), .ZN(n9261) );
  OAI22_X1 U10690 ( .A1(n9259), .A2(n9258), .B1(n9257), .B2(n9256), .ZN(n9260)
         );
  AOI211_X1 U10691 ( .C1(n9341), .C2(n9262), .A(n9261), .B(n9260), .ZN(n9265)
         );
  NAND2_X1 U10692 ( .A1(n9339), .A2(n9263), .ZN(n9264) );
  OAI211_X1 U10693 ( .C1(n9343), .C2(n10372), .A(n9265), .B(n9264), .ZN(
        P2_U3280) );
  NAND2_X1 U10694 ( .A1(n9266), .A2(n10444), .ZN(n9267) );
  OAI211_X1 U10695 ( .C1(n9268), .C2(n10455), .A(n9267), .B(n9271), .ZN(n9350)
         );
  MUX2_X1 U10696 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9350), .S(n10473), .Z(
        P2_U3551) );
  NAND3_X1 U10697 ( .A1(n9270), .A2(n10447), .A3(n9269), .ZN(n9272) );
  OAI211_X1 U10698 ( .C1(n9273), .C2(n10453), .A(n9272), .B(n9271), .ZN(n9351)
         );
  MUX2_X1 U10699 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9351), .S(n10473), .Z(
        P2_U3550) );
  AOI22_X1 U10700 ( .A1(n9275), .A2(n10447), .B1(n10444), .B2(n9274), .ZN(
        n9277) );
  MUX2_X1 U10701 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n9352), .S(n10473), .Z(
        P2_U3549) );
  AOI22_X1 U10702 ( .A1(n9281), .A2(n10447), .B1(n10444), .B2(n9280), .ZN(
        n9282) );
  OAI211_X1 U10703 ( .C1(n9926), .C2(n9284), .A(n9283), .B(n9282), .ZN(n9353)
         );
  MUX2_X1 U10704 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9353), .S(n10473), .Z(
        P2_U3548) );
  AOI22_X1 U10705 ( .A1(n9286), .A2(n10447), .B1(n10444), .B2(n9285), .ZN(
        n9287) );
  OAI211_X1 U10706 ( .C1(n9926), .C2(n9289), .A(n9288), .B(n9287), .ZN(n9354)
         );
  MUX2_X1 U10707 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9354), .S(n10473), .Z(
        P2_U3547) );
  AOI21_X1 U10708 ( .B1(n10444), .B2(n9291), .A(n9290), .ZN(n9292) );
  OAI211_X1 U10709 ( .C1(n9926), .C2(n9294), .A(n9293), .B(n9292), .ZN(n9355)
         );
  MUX2_X1 U10710 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9355), .S(n10473), .Z(
        P2_U3546) );
  AOI21_X1 U10711 ( .B1(n10444), .B2(n9296), .A(n9295), .ZN(n9297) );
  OAI211_X1 U10712 ( .C1(n9299), .C2(n9926), .A(n9298), .B(n9297), .ZN(n9356)
         );
  MUX2_X1 U10713 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9356), .S(n10473), .Z(
        P2_U3545) );
  AOI22_X1 U10714 ( .A1(n9301), .A2(n10447), .B1(n10444), .B2(n9300), .ZN(
        n9302) );
  OAI211_X1 U10715 ( .C1(n9926), .C2(n9304), .A(n9303), .B(n9302), .ZN(n9357)
         );
  MUX2_X1 U10716 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9357), .S(n10473), .Z(
        P2_U3544) );
  AOI22_X1 U10717 ( .A1(n9306), .A2(n10447), .B1(n10444), .B2(n9305), .ZN(
        n9307) );
  OAI211_X1 U10718 ( .C1(n9926), .C2(n9309), .A(n9308), .B(n9307), .ZN(n9358)
         );
  MUX2_X1 U10719 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9358), .S(n10473), .Z(
        P2_U3543) );
  AOI22_X1 U10720 ( .A1(n9311), .A2(n10447), .B1(n10444), .B2(n9310), .ZN(
        n9312) );
  OAI211_X1 U10721 ( .C1(n9926), .C2(n9314), .A(n9313), .B(n9312), .ZN(n9359)
         );
  MUX2_X1 U10722 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9359), .S(n10473), .Z(
        P2_U3542) );
  AOI22_X1 U10723 ( .A1(n9316), .A2(n10447), .B1(n10444), .B2(n9315), .ZN(
        n9317) );
  OAI211_X1 U10724 ( .C1(n9926), .C2(n9319), .A(n9318), .B(n9317), .ZN(n9360)
         );
  MUX2_X1 U10725 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9360), .S(n10473), .Z(
        P2_U3541) );
  AOI21_X1 U10726 ( .B1(n10444), .B2(n9321), .A(n9320), .ZN(n9322) );
  OAI211_X1 U10727 ( .C1(n9926), .C2(n9324), .A(n9323), .B(n9322), .ZN(n9361)
         );
  MUX2_X1 U10728 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9361), .S(n10473), .Z(
        P2_U3540) );
  AOI21_X1 U10729 ( .B1(n10444), .B2(n9326), .A(n9325), .ZN(n9327) );
  OAI21_X1 U10730 ( .B1(n9926), .B2(n9328), .A(n9327), .ZN(n9362) );
  MUX2_X1 U10731 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9362), .S(n10473), .Z(
        P2_U3539) );
  AOI22_X1 U10732 ( .A1(n9330), .A2(n10447), .B1(n10444), .B2(n9329), .ZN(
        n9331) );
  OAI211_X1 U10733 ( .C1(n9926), .C2(n9333), .A(n9332), .B(n9331), .ZN(n9363)
         );
  MUX2_X1 U10734 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9363), .S(n10473), .Z(
        P2_U3538) );
  AOI21_X1 U10735 ( .B1(n10444), .B2(n9335), .A(n9334), .ZN(n9336) );
  OAI211_X1 U10736 ( .C1(n9926), .C2(n9338), .A(n9337), .B(n9336), .ZN(n9364)
         );
  MUX2_X1 U10737 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9364), .S(n10473), .Z(
        P2_U3537) );
  INV_X1 U10738 ( .A(n9339), .ZN(n9344) );
  AOI22_X1 U10739 ( .A1(n9341), .A2(n10447), .B1(n10444), .B2(n9340), .ZN(
        n9342) );
  OAI211_X1 U10740 ( .C1(n10428), .C2(n9344), .A(n9343), .B(n9342), .ZN(n9365)
         );
  MUX2_X1 U10741 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9365), .S(n10473), .Z(
        P2_U3536) );
  AOI21_X1 U10742 ( .B1(n10444), .B2(n9346), .A(n9345), .ZN(n9347) );
  OAI211_X1 U10743 ( .C1(n9926), .C2(n9349), .A(n9348), .B(n9347), .ZN(n9366)
         );
  MUX2_X1 U10744 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n9366), .S(n10473), .Z(
        P2_U3535) );
  MUX2_X1 U10745 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9350), .S(n10462), .Z(
        P2_U3519) );
  MUX2_X1 U10746 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9351), .S(n10462), .Z(
        P2_U3518) );
  MUX2_X1 U10747 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9352), .S(n10462), .Z(
        P2_U3517) );
  MUX2_X1 U10748 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9353), .S(n10462), .Z(
        P2_U3516) );
  MUX2_X1 U10749 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9354), .S(n10462), .Z(
        P2_U3515) );
  MUX2_X1 U10750 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9355), .S(n10462), .Z(
        P2_U3514) );
  MUX2_X1 U10751 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9356), .S(n10462), .Z(
        P2_U3513) );
  MUX2_X1 U10752 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9357), .S(n10462), .Z(
        P2_U3512) );
  MUX2_X1 U10753 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9358), .S(n10462), .Z(
        P2_U3511) );
  MUX2_X1 U10754 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9359), .S(n10462), .Z(
        P2_U3510) );
  MUX2_X1 U10755 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9360), .S(n10462), .Z(
        P2_U3509) );
  MUX2_X1 U10756 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9361), .S(n10462), .Z(
        P2_U3508) );
  MUX2_X1 U10757 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9362), .S(n10462), .Z(
        P2_U3507) );
  MUX2_X1 U10758 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9363), .S(n10462), .Z(
        P2_U3505) );
  MUX2_X1 U10759 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9364), .S(n10462), .Z(
        P2_U3502) );
  MUX2_X1 U10760 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9365), .S(n10462), .Z(
        P2_U3499) );
  MUX2_X1 U10761 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n9366), .S(n10462), .Z(
        P2_U3496) );
  INV_X1 U10762 ( .A(n9367), .ZN(n9887) );
  INV_X1 U10763 ( .A(n9368), .ZN(n9370) );
  NOR4_X1 U10764 ( .A1(n9370), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3152), .A4(
        n9369), .ZN(n9371) );
  AOI21_X1 U10765 ( .B1(n9372), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9371), .ZN(
        n9373) );
  OAI21_X1 U10766 ( .B1(n9887), .B2(n9376), .A(n9373), .ZN(P2_U3327) );
  OAI222_X1 U10767 ( .A1(P2_U3152), .A2(n9377), .B1(n9376), .B2(n9375), .C1(
        n9374), .C2(n9382), .ZN(P2_U3329) );
  NAND2_X1 U10768 ( .A1(n9888), .A2(n9378), .ZN(n9380) );
  OAI211_X1 U10769 ( .C1(n9382), .C2(n9381), .A(n9380), .B(n9379), .ZN(
        P2_U3330) );
  INV_X1 U10770 ( .A(n9893), .ZN(n9384) );
  OAI222_X1 U10771 ( .A1(P2_U3152), .A2(n9385), .B1(n9376), .B2(n9384), .C1(
        n9383), .C2(n9382), .ZN(P2_U3331) );
  MUX2_X1 U10772 ( .A(n9386), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  XNOR2_X1 U10773 ( .A(n9388), .B(n9387), .ZN(n9389) );
  XNOR2_X1 U10774 ( .A(n9390), .B(n9389), .ZN(n9395) );
  AOI22_X1 U10775 ( .A1(n9495), .A2(n9627), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n9392) );
  NAND2_X1 U10776 ( .A1(n9507), .A2(n9517), .ZN(n9391) );
  OAI211_X1 U10777 ( .C1(n9510), .C2(n9591), .A(n9392), .B(n9391), .ZN(n9393)
         );
  AOI21_X1 U10778 ( .B1(n9789), .B2(n9512), .A(n9393), .ZN(n9394) );
  OAI21_X1 U10779 ( .B1(n9395), .B2(n9514), .A(n9394), .ZN(P1_U3212) );
  INV_X1 U10780 ( .A(n9396), .ZN(n9400) );
  OR2_X1 U10781 ( .A1(n9397), .A2(n9396), .ZN(n9398) );
  AOI22_X1 U10782 ( .A1(n9401), .A2(n9400), .B1(n9399), .B2(n9398), .ZN(n9406)
         );
  NAND2_X1 U10783 ( .A1(n9662), .A2(n9495), .ZN(n9403) );
  AOI22_X1 U10784 ( .A1(n9507), .A2(n9663), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9402) );
  OAI211_X1 U10785 ( .C1(n9656), .C2(n9510), .A(n9403), .B(n9402), .ZN(n9404)
         );
  AOI21_X1 U10786 ( .B1(n9811), .B2(n9512), .A(n9404), .ZN(n9405) );
  OAI21_X1 U10787 ( .B1(n9406), .B2(n9514), .A(n9405), .ZN(P1_U3214) );
  OAI21_X1 U10788 ( .B1(n9409), .B2(n9408), .A(n9407), .ZN(n9410) );
  NAND2_X1 U10789 ( .A1(n9410), .A2(n9483), .ZN(n9414) );
  NOR2_X1 U10790 ( .A1(n9510), .A2(n9720), .ZN(n9412) );
  NAND2_X1 U10791 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9562) );
  OAI21_X1 U10792 ( .B1(n9718), .B2(n9486), .A(n9562), .ZN(n9411) );
  AOI211_X1 U10793 ( .C1(n9495), .C2(n9752), .A(n9412), .B(n9411), .ZN(n9413)
         );
  OAI211_X1 U10794 ( .C1(n4853), .C2(n9492), .A(n9414), .B(n9413), .ZN(
        P1_U3217) );
  XOR2_X1 U10795 ( .A(n9416), .B(n9415), .Z(n9421) );
  NAND2_X1 U10796 ( .A1(n9662), .A2(n9507), .ZN(n9418) );
  AOI22_X1 U10797 ( .A1(n9519), .A2(n9495), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9417) );
  OAI211_X1 U10798 ( .C1(n9510), .C2(n9692), .A(n9418), .B(n9417), .ZN(n9419)
         );
  AOI21_X1 U10799 ( .B1(n9823), .B2(n9512), .A(n9419), .ZN(n9420) );
  OAI21_X1 U10800 ( .B1(n9421), .B2(n9514), .A(n9420), .ZN(P1_U3221) );
  XOR2_X1 U10801 ( .A(n9423), .B(n9422), .Z(n9428) );
  AOI22_X1 U10802 ( .A1(n9507), .A2(n9627), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9425) );
  NAND2_X1 U10803 ( .A1(n9495), .A2(n9663), .ZN(n9424) );
  OAI211_X1 U10804 ( .C1(n9510), .C2(n9620), .A(n9425), .B(n9424), .ZN(n9426)
         );
  AOI21_X1 U10805 ( .B1(n9799), .B2(n9512), .A(n9426), .ZN(n9427) );
  OAI21_X1 U10806 ( .B1(n9428), .B2(n9514), .A(n9427), .ZN(P1_U3223) );
  INV_X1 U10807 ( .A(n9429), .ZN(n9434) );
  AOI21_X1 U10808 ( .B1(n9432), .B2(n9430), .A(n9431), .ZN(n9433) );
  OAI21_X1 U10809 ( .B1(n9434), .B2(n9433), .A(n9483), .ZN(n9441) );
  INV_X1 U10810 ( .A(n9435), .ZN(n9764) );
  NOR2_X1 U10811 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9436), .ZN(n10119) );
  AOI21_X1 U10812 ( .B1(n9507), .B2(n9771), .A(n10119), .ZN(n9437) );
  OAI21_X1 U10813 ( .B1(n9505), .B2(n9438), .A(n9437), .ZN(n9439) );
  AOI21_X1 U10814 ( .B1(n9466), .B2(n9764), .A(n9439), .ZN(n9440) );
  OAI211_X1 U10815 ( .C1(n9766), .C2(n9492), .A(n9441), .B(n9440), .ZN(
        P1_U3224) );
  OAI21_X1 U10816 ( .B1(n9444), .B2(n9443), .A(n9442), .ZN(n9445) );
  NAND2_X1 U10817 ( .A1(n9445), .A2(n9483), .ZN(n9449) );
  NAND2_X1 U10818 ( .A1(P1_U3084), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10127)
         );
  OAI21_X1 U10819 ( .B1(n9486), .B2(n9717), .A(n10127), .ZN(n9447) );
  NOR2_X1 U10820 ( .A1(n9510), .A2(n9744), .ZN(n9446) );
  AOI211_X1 U10821 ( .C1(n9495), .C2(n9751), .A(n9447), .B(n9446), .ZN(n9448)
         );
  OAI211_X1 U10822 ( .C1(n4834), .C2(n9492), .A(n9449), .B(n9448), .ZN(
        P1_U3226) );
  AOI21_X1 U10823 ( .B1(n4527), .B2(n9451), .A(n9450), .ZN(n9457) );
  AND2_X1 U10824 ( .A1(n9633), .A2(n9849), .ZN(n9806) );
  AOI22_X1 U10825 ( .A1(n9507), .A2(n9518), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9453) );
  NAND2_X1 U10826 ( .A1(n9495), .A2(n9677), .ZN(n9452) );
  OAI211_X1 U10827 ( .C1(n9510), .C2(n9642), .A(n9453), .B(n9452), .ZN(n9454)
         );
  AOI21_X1 U10828 ( .B1(n9806), .B2(n9455), .A(n9454), .ZN(n9456) );
  OAI21_X1 U10829 ( .B1(n9457), .B2(n9514), .A(n9456), .ZN(P1_U3227) );
  NOR2_X1 U10830 ( .A1(n9458), .A2(n4991), .ZN(n9463) );
  AOI21_X1 U10831 ( .B1(n9461), .B2(n9460), .A(n9459), .ZN(n9462) );
  OAI21_X1 U10832 ( .B1(n9463), .B2(n9462), .A(n9483), .ZN(n9468) );
  AOI22_X1 U10833 ( .A1(n9707), .A2(n9507), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9464) );
  OAI21_X1 U10834 ( .B1(n9487), .B2(n9505), .A(n9464), .ZN(n9465) );
  AOI21_X1 U10835 ( .B1(n9701), .B2(n9466), .A(n9465), .ZN(n9467) );
  OAI211_X1 U10836 ( .C1(n9703), .C2(n9492), .A(n9468), .B(n9467), .ZN(
        P1_U3231) );
  NAND2_X1 U10837 ( .A1(n9470), .A2(n9469), .ZN(n9471) );
  XOR2_X1 U10838 ( .A(n9472), .B(n9471), .Z(n9477) );
  NAND2_X1 U10839 ( .A1(n9707), .A2(n9495), .ZN(n9474) );
  AOI22_X1 U10840 ( .A1(n9507), .A2(n9677), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9473) );
  OAI211_X1 U10841 ( .C1(n9510), .C2(n9670), .A(n9474), .B(n9473), .ZN(n9475)
         );
  AOI21_X1 U10842 ( .B1(n9816), .B2(n9512), .A(n9475), .ZN(n9476) );
  OAI21_X1 U10843 ( .B1(n9477), .B2(n9514), .A(n9476), .ZN(P1_U3233) );
  INV_X1 U10844 ( .A(n9838), .ZN(n9733) );
  INV_X1 U10845 ( .A(n9481), .ZN(n9478) );
  NOR2_X1 U10846 ( .A1(n9479), .A2(n9478), .ZN(n9485) );
  AOI21_X1 U10847 ( .B1(n9482), .B2(n9481), .A(n9480), .ZN(n9484) );
  OAI21_X1 U10848 ( .B1(n9485), .B2(n9484), .A(n9483), .ZN(n9491) );
  NAND2_X1 U10849 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10141)
         );
  OAI21_X1 U10850 ( .B1(n9487), .B2(n9486), .A(n10141), .ZN(n9489) );
  NOR2_X1 U10851 ( .A1(n9510), .A2(n9734), .ZN(n9488) );
  AOI211_X1 U10852 ( .C1(n9495), .C2(n9771), .A(n9489), .B(n9488), .ZN(n9490)
         );
  OAI211_X1 U10853 ( .C1(n9733), .C2(n9492), .A(n9491), .B(n9490), .ZN(
        P1_U3236) );
  XOR2_X1 U10854 ( .A(n9494), .B(n9493), .Z(n9500) );
  AOI22_X1 U10855 ( .A1(n9495), .A2(n9518), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9497) );
  NAND2_X1 U10856 ( .A1(n9507), .A2(n9576), .ZN(n9496) );
  OAI211_X1 U10857 ( .C1(n9510), .C2(n9610), .A(n9497), .B(n9496), .ZN(n9498)
         );
  AOI21_X1 U10858 ( .B1(n9796), .B2(n9512), .A(n9498), .ZN(n9499) );
  OAI21_X1 U10859 ( .B1(n9500), .B2(n9514), .A(n9499), .ZN(P1_U3238) );
  NAND2_X1 U10860 ( .A1(n9430), .A2(n9501), .ZN(n9502) );
  XOR2_X1 U10861 ( .A(n9503), .B(n9502), .Z(n9515) );
  AND2_X1 U10862 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10108) );
  NOR2_X1 U10863 ( .A1(n9505), .A2(n9504), .ZN(n9506) );
  AOI211_X1 U10864 ( .C1(n9507), .C2(n9751), .A(n10108), .B(n9506), .ZN(n9508)
         );
  OAI21_X1 U10865 ( .B1(n9510), .B2(n9509), .A(n9508), .ZN(n9511) );
  AOI21_X1 U10866 ( .B1(n9856), .B2(n9512), .A(n9511), .ZN(n9513) );
  OAI21_X1 U10867 ( .B1(n9515), .B2(n9514), .A(n9513), .ZN(P1_U3239) );
  MUX2_X1 U10868 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9516), .S(n9527), .Z(
        P1_U3585) );
  MUX2_X1 U10869 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9577), .S(n9527), .Z(
        P1_U3584) );
  MUX2_X1 U10870 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9517), .S(n9527), .Z(
        P1_U3583) );
  MUX2_X1 U10871 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9576), .S(n9527), .Z(
        P1_U3582) );
  MUX2_X1 U10872 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9627), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10873 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9518), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10874 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9663), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10875 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9662), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10876 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9707), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10877 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9519), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10878 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9727), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10879 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9752), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10880 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9771), .S(n9527), .Z(
        P1_U3572) );
  MUX2_X1 U10881 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9751), .S(n9527), .Z(
        P1_U3571) );
  MUX2_X1 U10882 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9770), .S(n9527), .Z(
        P1_U3570) );
  MUX2_X1 U10883 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9946), .S(n9527), .Z(
        P1_U3569) );
  MUX2_X1 U10884 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9520), .S(n9527), .Z(
        P1_U3568) );
  MUX2_X1 U10885 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9944), .S(n9527), .Z(
        P1_U3567) );
  MUX2_X1 U10886 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n9521), .S(n9527), .Z(
        P1_U3566) );
  MUX2_X1 U10887 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9522), .S(n9527), .Z(
        P1_U3565) );
  MUX2_X1 U10888 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9523), .S(n9527), .Z(
        P1_U3564) );
  MUX2_X1 U10889 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9524), .S(n9527), .Z(
        P1_U3563) );
  MUX2_X1 U10890 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9525), .S(n9527), .Z(
        P1_U3562) );
  MUX2_X1 U10891 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9526), .S(n9527), .Z(
        P1_U3561) );
  MUX2_X1 U10892 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9528), .S(n9527), .Z(
        P1_U3560) );
  MUX2_X1 U10893 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9529), .S(P1_U4006), .Z(
        P1_U3559) );
  MUX2_X1 U10894 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9530), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10895 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n6925), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10896 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n9531), .S(P1_U4006), .Z(
        P1_U3556) );
  NAND2_X1 U10897 ( .A1(n9532), .A2(n9541), .ZN(n9534) );
  INV_X1 U10898 ( .A(n9535), .ZN(n9536) );
  XNOR2_X1 U10899 ( .A(n9535), .B(n9544), .ZN(n10106) );
  NAND2_X1 U10900 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n10120), .ZN(n9537) );
  OAI21_X1 U10901 ( .B1(n10120), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9537), .ZN(
        n10116) );
  NAND2_X1 U10902 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n10133), .ZN(n9538) );
  OAI21_X1 U10903 ( .B1(n10133), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9538), .ZN(
        n10129) );
  NOR2_X1 U10904 ( .A1(n10130), .A2(n10129), .ZN(n10128) );
  NOR2_X1 U10905 ( .A1(n10149), .A2(n9735), .ZN(n9539) );
  AOI21_X1 U10906 ( .B1(n10149), .B2(n9735), .A(n9539), .ZN(n10144) );
  XNOR2_X1 U10907 ( .A(n10149), .B(P1_REG1_REG_18__SCAN_IN), .ZN(n10152) );
  INV_X1 U10908 ( .A(n10133), .ZN(n9549) );
  XOR2_X1 U10909 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10133), .Z(n10137) );
  INV_X1 U10910 ( .A(n10120), .ZN(n9547) );
  XOR2_X1 U10911 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10120), .Z(n10122) );
  AOI21_X1 U10912 ( .B1(n6200), .B2(n9541), .A(n9540), .ZN(n9542) );
  XNOR2_X1 U10913 ( .A(n9542), .B(n10109), .ZN(n10110) );
  INV_X1 U10914 ( .A(n9542), .ZN(n9543) );
  OAI22_X1 U10915 ( .A1(n10110), .A2(n9545), .B1(n9544), .B2(n9543), .ZN(
        n10123) );
  NAND2_X1 U10916 ( .A1(n10122), .A2(n10123), .ZN(n10121) );
  OAI21_X1 U10917 ( .B1(n9547), .B2(n9546), .A(n10121), .ZN(n10136) );
  NAND2_X1 U10918 ( .A1(n10137), .A2(n10136), .ZN(n10134) );
  OAI21_X1 U10919 ( .B1(n9549), .B2(n9548), .A(n10134), .ZN(n10151) );
  NOR2_X1 U10920 ( .A1(n10152), .A2(n10151), .ZN(n10150) );
  AOI21_X1 U10921 ( .B1(n9551), .B2(n9550), .A(n10150), .ZN(n9553) );
  XOR2_X1 U10922 ( .A(n9553), .B(n9552), .Z(n9557) );
  OAI22_X1 U10923 ( .A1(n9556), .A2(n10142), .B1(n9557), .B2(n10154), .ZN(
        n9561) );
  NAND3_X1 U10924 ( .A1(n9556), .A2(n9555), .A3(n9554), .ZN(n9559) );
  AOI21_X1 U10925 ( .B1(n9557), .B2(n10135), .A(n10148), .ZN(n9558) );
  NAND2_X1 U10926 ( .A1(n9559), .A2(n9558), .ZN(n9560) );
  MUX2_X1 U10927 ( .A(n9561), .B(n9560), .S(n4695), .Z(n9564) );
  OAI21_X1 U10928 ( .B1(n10157), .B2(n4979), .A(n9562), .ZN(n9563) );
  XNOR2_X1 U10929 ( .A(n9566), .B(n9565), .ZN(n9983) );
  NAND2_X1 U10930 ( .A1(n9983), .A2(n10163), .ZN(n9569) );
  AOI21_X1 U10931 ( .B1(n9953), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9567), .ZN(
        n9568) );
  OAI211_X1 U10932 ( .C1(n9981), .C2(n10177), .A(n9569), .B(n9568), .ZN(
        P1_U3262) );
  AND2_X1 U10933 ( .A1(n9571), .A2(n9570), .ZN(n9572) );
  XNOR2_X1 U10934 ( .A(n9574), .B(n9573), .ZN(n9575) );
  NAND2_X1 U10935 ( .A1(n9575), .A2(n10172), .ZN(n9579) );
  AOI22_X1 U10936 ( .A1(n9947), .A2(n9577), .B1(n9945), .B2(n9576), .ZN(n9578)
         );
  NAND2_X1 U10937 ( .A1(n9579), .A2(n9578), .ZN(n9786) );
  NAND2_X1 U10938 ( .A1(n9783), .A2(n9590), .ZN(n9580) );
  NAND3_X1 U10939 ( .A1(n9581), .A2(n9984), .A3(n9580), .ZN(n9784) );
  OAI22_X1 U10940 ( .A1(n10181), .A2(n9583), .B1(n9582), .B2(n10178), .ZN(
        n9584) );
  AOI21_X1 U10941 ( .B1(n9783), .B2(n9957), .A(n9584), .ZN(n9585) );
  OAI21_X1 U10942 ( .B1(n9784), .B2(n9586), .A(n9585), .ZN(n9587) );
  AOI21_X1 U10943 ( .B1(n9786), .B2(n10181), .A(n9587), .ZN(n9588) );
  OAI21_X1 U10944 ( .B1(n9788), .B2(n9777), .A(n9588), .ZN(P1_U3263) );
  XNOR2_X1 U10945 ( .A(n9589), .B(n9595), .ZN(n9793) );
  AOI21_X1 U10946 ( .B1(n9789), .B2(n9607), .A(n4845), .ZN(n9790) );
  INV_X1 U10947 ( .A(n9789), .ZN(n9594) );
  INV_X1 U10948 ( .A(n9591), .ZN(n9592) );
  AOI22_X1 U10949 ( .A1(n9953), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n9592), .B2(
        n9763), .ZN(n9593) );
  OAI21_X1 U10950 ( .B1(n9594), .B2(n10177), .A(n9593), .ZN(n9603) );
  AOI21_X1 U10951 ( .B1(n9596), .B2(n9595), .A(n9949), .ZN(n9601) );
  OAI22_X1 U10952 ( .A1(n10170), .A2(n9598), .B1(n9597), .B2(n10167), .ZN(
        n9599) );
  AOI21_X1 U10953 ( .B1(n9601), .B2(n9600), .A(n9599), .ZN(n9792) );
  NOR2_X1 U10954 ( .A1(n9792), .A2(n9953), .ZN(n9602) );
  AOI211_X1 U10955 ( .C1(n9790), .C2(n10163), .A(n9603), .B(n9602), .ZN(n9604)
         );
  OAI21_X1 U10956 ( .B1(n9793), .B2(n9777), .A(n9604), .ZN(P1_U3264) );
  XNOR2_X1 U10957 ( .A(n9606), .B(n9605), .ZN(n9798) );
  AOI22_X1 U10958 ( .A1(n9796), .A2(n9957), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n9953), .ZN(n9617) );
  INV_X1 U10959 ( .A(n9619), .ZN(n9609) );
  INV_X1 U10960 ( .A(n9607), .ZN(n9608) );
  AOI211_X1 U10961 ( .C1(n9796), .C2(n9609), .A(n10228), .B(n9608), .ZN(n9795)
         );
  INV_X1 U10962 ( .A(n9795), .ZN(n9611) );
  OAI22_X1 U10963 ( .A1(n9611), .A2(n4695), .B1(n10178), .B2(n9610), .ZN(n9615) );
  XNOR2_X1 U10964 ( .A(n9612), .B(n4752), .ZN(n9613) );
  OAI222_X1 U10965 ( .A1(n10167), .A2(n9614), .B1(n10170), .B2(n9643), .C1(
        n9949), .C2(n9613), .ZN(n9794) );
  OAI21_X1 U10966 ( .B1(n9615), .B2(n9794), .A(n10181), .ZN(n9616) );
  OAI211_X1 U10967 ( .C1(n9798), .C2(n9777), .A(n9617), .B(n9616), .ZN(
        P1_U3265) );
  XNOR2_X1 U10968 ( .A(n9618), .B(n9626), .ZN(n9803) );
  AOI21_X1 U10969 ( .B1(n9799), .B2(n9634), .A(n9619), .ZN(n9800) );
  INV_X1 U10970 ( .A(n9799), .ZN(n9623) );
  INV_X1 U10971 ( .A(n9620), .ZN(n9621) );
  AOI22_X1 U10972 ( .A1(n9953), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9621), .B2(
        n9763), .ZN(n9622) );
  OAI21_X1 U10973 ( .B1(n9623), .B2(n10177), .A(n9622), .ZN(n9630) );
  OAI21_X1 U10974 ( .B1(n9626), .B2(n9625), .A(n9624), .ZN(n9628) );
  AOI222_X1 U10975 ( .A1(n10172), .A2(n9628), .B1(n9627), .B2(n9947), .C1(
        n9663), .C2(n9945), .ZN(n9802) );
  NOR2_X1 U10976 ( .A1(n9802), .A2(n9953), .ZN(n9629) );
  AOI211_X1 U10977 ( .C1(n9800), .C2(n10163), .A(n9630), .B(n9629), .ZN(n9631)
         );
  OAI21_X1 U10978 ( .B1(n9803), .B2(n9777), .A(n9631), .ZN(P1_U3266) );
  XNOR2_X1 U10979 ( .A(n9632), .B(n9638), .ZN(n9804) );
  INV_X1 U10980 ( .A(n9804), .ZN(n9651) );
  AOI22_X1 U10981 ( .A1(n9633), .A2(n9957), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n9953), .ZN(n9650) );
  AOI21_X1 U10982 ( .B1(n9633), .B2(n9653), .A(n10228), .ZN(n9635) );
  NAND2_X1 U10983 ( .A1(n9635), .A2(n9634), .ZN(n9807) );
  NAND2_X1 U10984 ( .A1(n9637), .A2(n9636), .ZN(n9640) );
  INV_X1 U10985 ( .A(n9638), .ZN(n9639) );
  XNOR2_X1 U10986 ( .A(n9640), .B(n9639), .ZN(n9641) );
  NAND2_X1 U10987 ( .A1(n9641), .A2(n10172), .ZN(n9808) );
  INV_X1 U10988 ( .A(n9642), .ZN(n9646) );
  NAND2_X1 U10989 ( .A1(n9945), .A2(n9677), .ZN(n9645) );
  OR2_X1 U10990 ( .A1(n9643), .A2(n10167), .ZN(n9644) );
  NAND2_X1 U10991 ( .A1(n9645), .A2(n9644), .ZN(n9805) );
  AOI21_X1 U10992 ( .B1(n9646), .B2(n9763), .A(n9805), .ZN(n9647) );
  OAI211_X1 U10993 ( .C1(n4695), .C2(n9807), .A(n9808), .B(n9647), .ZN(n9648)
         );
  NAND2_X1 U10994 ( .A1(n9648), .A2(n10181), .ZN(n9649) );
  OAI211_X1 U10995 ( .C1(n9651), .C2(n9777), .A(n9650), .B(n9649), .ZN(
        P1_U3267) );
  XOR2_X1 U10996 ( .A(n9652), .B(n9660), .Z(n9815) );
  INV_X1 U10997 ( .A(n9669), .ZN(n9655) );
  INV_X1 U10998 ( .A(n9653), .ZN(n9654) );
  AOI21_X1 U10999 ( .B1(n9811), .B2(n9655), .A(n9654), .ZN(n9812) );
  INV_X1 U11000 ( .A(n9656), .ZN(n9657) );
  AOI22_X1 U11001 ( .A1(n9953), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9763), .B2(
        n9657), .ZN(n9658) );
  OAI21_X1 U11002 ( .B1(n9659), .B2(n10177), .A(n9658), .ZN(n9666) );
  XNOR2_X1 U11003 ( .A(n9661), .B(n9660), .ZN(n9664) );
  AOI222_X1 U11004 ( .A1(n10172), .A2(n9664), .B1(n9663), .B2(n9947), .C1(
        n9662), .C2(n9945), .ZN(n9814) );
  NOR2_X1 U11005 ( .A1(n9814), .A2(n9953), .ZN(n9665) );
  AOI211_X1 U11006 ( .C1(n9812), .C2(n10163), .A(n9666), .B(n9665), .ZN(n9667)
         );
  OAI21_X1 U11007 ( .B1(n9815), .B2(n9777), .A(n9667), .ZN(P1_U3268) );
  XNOR2_X1 U11008 ( .A(n9668), .B(n9676), .ZN(n9820) );
  AOI21_X1 U11009 ( .B1(n9816), .B2(n9690), .A(n9669), .ZN(n9817) );
  INV_X1 U11010 ( .A(n9816), .ZN(n9673) );
  INV_X1 U11011 ( .A(n9670), .ZN(n9671) );
  AOI22_X1 U11012 ( .A1(n9671), .A2(n9763), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n9953), .ZN(n9672) );
  OAI21_X1 U11013 ( .B1(n9673), .B2(n10177), .A(n9672), .ZN(n9680) );
  NAND2_X1 U11014 ( .A1(n9684), .A2(n9674), .ZN(n9675) );
  XOR2_X1 U11015 ( .A(n9676), .B(n9675), .Z(n9678) );
  AOI222_X1 U11016 ( .A1(n10172), .A2(n9678), .B1(n9707), .B2(n9945), .C1(
        n9677), .C2(n9947), .ZN(n9819) );
  NOR2_X1 U11017 ( .A1(n9819), .A2(n9953), .ZN(n9679) );
  AOI211_X1 U11018 ( .C1(n9817), .C2(n10163), .A(n9680), .B(n9679), .ZN(n9681)
         );
  OAI21_X1 U11019 ( .B1(n9777), .B2(n9820), .A(n9681), .ZN(P1_U3269) );
  XNOR2_X1 U11020 ( .A(n9682), .B(n9687), .ZN(n9825) );
  AOI22_X1 U11021 ( .A1(n9823), .A2(n9957), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n9953), .ZN(n9696) );
  NAND2_X1 U11022 ( .A1(n9704), .A2(n9683), .ZN(n9686) );
  INV_X1 U11023 ( .A(n9684), .ZN(n9685) );
  AOI21_X1 U11024 ( .B1(n9687), .B2(n9686), .A(n9685), .ZN(n9688) );
  OAI222_X1 U11025 ( .A1(n10167), .A2(n9689), .B1(n10170), .B2(n9718), .C1(
        n9949), .C2(n9688), .ZN(n9821) );
  INV_X1 U11026 ( .A(n9690), .ZN(n9691) );
  AOI211_X1 U11027 ( .C1(n9823), .C2(n9699), .A(n10228), .B(n9691), .ZN(n9822)
         );
  INV_X1 U11028 ( .A(n9822), .ZN(n9693) );
  OAI22_X1 U11029 ( .A1(n9693), .A2(n4695), .B1(n10178), .B2(n9692), .ZN(n9694) );
  OAI21_X1 U11030 ( .B1(n9821), .B2(n9694), .A(n10181), .ZN(n9695) );
  OAI211_X1 U11031 ( .C1(n9825), .C2(n9777), .A(n9696), .B(n9695), .ZN(
        P1_U3270) );
  XNOR2_X1 U11032 ( .A(n9698), .B(n9697), .ZN(n9830) );
  INV_X1 U11033 ( .A(n9699), .ZN(n9700) );
  AOI21_X1 U11034 ( .B1(n9826), .B2(n4855), .A(n9700), .ZN(n9827) );
  AOI22_X1 U11035 ( .A1(n9953), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n9701), .B2(
        n9763), .ZN(n9702) );
  OAI21_X1 U11036 ( .B1(n9703), .B2(n10177), .A(n9702), .ZN(n9711) );
  OAI211_X1 U11037 ( .C1(n9706), .C2(n9705), .A(n9704), .B(n10172), .ZN(n9709)
         );
  AOI22_X1 U11038 ( .A1(n9707), .A2(n9947), .B1(n9945), .B2(n9727), .ZN(n9708)
         );
  AND2_X1 U11039 ( .A1(n9709), .A2(n9708), .ZN(n9829) );
  NOR2_X1 U11040 ( .A1(n9829), .A2(n9953), .ZN(n9710) );
  AOI211_X1 U11041 ( .C1(n9827), .C2(n10163), .A(n9711), .B(n9710), .ZN(n9712)
         );
  OAI21_X1 U11042 ( .B1(n9830), .B2(n9777), .A(n9712), .ZN(P1_U3271) );
  XNOR2_X1 U11043 ( .A(n9713), .B(n9714), .ZN(n9835) );
  XNOR2_X1 U11044 ( .A(n9715), .B(n9714), .ZN(n9716) );
  OAI222_X1 U11045 ( .A1(n10167), .A2(n9718), .B1(n10170), .B2(n9717), .C1(
        n9716), .C2(n9949), .ZN(n9831) );
  AOI211_X1 U11046 ( .C1(n9833), .C2(n9731), .A(n10228), .B(n9719), .ZN(n9832)
         );
  NAND2_X1 U11047 ( .A1(n9832), .A2(n9747), .ZN(n9723) );
  INV_X1 U11048 ( .A(n9720), .ZN(n9721) );
  AOI22_X1 U11049 ( .A1(n9953), .A2(P1_REG2_REG_19__SCAN_IN), .B1(n9721), .B2(
        n9763), .ZN(n9722) );
  OAI211_X1 U11050 ( .C1(n4853), .C2(n10177), .A(n9723), .B(n9722), .ZN(n9724)
         );
  AOI21_X1 U11051 ( .B1(n9831), .B2(n10181), .A(n9724), .ZN(n9725) );
  OAI21_X1 U11052 ( .B1(n9835), .B2(n9777), .A(n9725), .ZN(P1_U3272) );
  OAI21_X1 U11053 ( .B1(n4566), .B2(n4758), .A(n9726), .ZN(n9728) );
  AOI222_X1 U11054 ( .A1(n10172), .A2(n9728), .B1(n9727), .B2(n9947), .C1(
        n9771), .C2(n9945), .ZN(n9841) );
  NAND2_X1 U11055 ( .A1(n9729), .A2(n4758), .ZN(n9836) );
  NAND3_X1 U11056 ( .A1(n9837), .A2(n9836), .A3(n9730), .ZN(n9739) );
  INV_X1 U11057 ( .A(n9731), .ZN(n9732) );
  AOI21_X1 U11058 ( .B1(n9838), .B2(n9741), .A(n9732), .ZN(n9839) );
  NOR2_X1 U11059 ( .A1(n9733), .A2(n10177), .ZN(n9737) );
  OAI22_X1 U11060 ( .A1(n10181), .A2(n9735), .B1(n9734), .B2(n10178), .ZN(
        n9736) );
  AOI211_X1 U11061 ( .C1(n9839), .C2(n10163), .A(n9737), .B(n9736), .ZN(n9738)
         );
  OAI211_X1 U11062 ( .C1(n9953), .C2(n9841), .A(n9739), .B(n9738), .ZN(
        P1_U3273) );
  XOR2_X1 U11063 ( .A(n9740), .B(n9749), .Z(n9847) );
  INV_X1 U11064 ( .A(n9761), .ZN(n9743) );
  INV_X1 U11065 ( .A(n9741), .ZN(n9742) );
  AOI211_X1 U11066 ( .C1(n9845), .C2(n9743), .A(n10228), .B(n9742), .ZN(n9844)
         );
  NOR2_X1 U11067 ( .A1(n4834), .A2(n10177), .ZN(n9746) );
  OAI22_X1 U11068 ( .A1(n10181), .A2(n4600), .B1(n9744), .B2(n10178), .ZN(
        n9745) );
  AOI211_X1 U11069 ( .C1(n9844), .C2(n9747), .A(n9746), .B(n9745), .ZN(n9757)
         );
  NAND2_X1 U11070 ( .A1(n9748), .A2(n10172), .ZN(n9755) );
  AOI21_X1 U11071 ( .B1(n9767), .B2(n9750), .A(n9749), .ZN(n9754) );
  AOI22_X1 U11072 ( .A1(n9752), .A2(n9947), .B1(n9945), .B2(n9751), .ZN(n9753)
         );
  OAI21_X1 U11073 ( .B1(n9755), .B2(n9754), .A(n9753), .ZN(n9843) );
  NAND2_X1 U11074 ( .A1(n9843), .A2(n10181), .ZN(n9756) );
  OAI211_X1 U11075 ( .C1(n9847), .C2(n9777), .A(n9757), .B(n9756), .ZN(
        P1_U3274) );
  XNOR2_X1 U11076 ( .A(n9759), .B(n9758), .ZN(n9854) );
  INV_X1 U11077 ( .A(n9760), .ZN(n9762) );
  AOI211_X1 U11078 ( .C1(n9850), .C2(n9762), .A(n10228), .B(n9761), .ZN(n9848)
         );
  AOI22_X1 U11079 ( .A1(n9953), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9764), .B2(
        n9763), .ZN(n9765) );
  OAI21_X1 U11080 ( .B1(n9766), .B2(n10177), .A(n9765), .ZN(n9774) );
  OAI21_X1 U11081 ( .B1(n9769), .B2(n9768), .A(n9767), .ZN(n9772) );
  AOI222_X1 U11082 ( .A1(n10172), .A2(n9772), .B1(n9771), .B2(n9947), .C1(
        n9770), .C2(n9945), .ZN(n9852) );
  NOR2_X1 U11083 ( .A1(n9852), .A2(n9953), .ZN(n9773) );
  AOI211_X1 U11084 ( .C1(n9848), .C2(n9775), .A(n9774), .B(n9773), .ZN(n9776)
         );
  OAI21_X1 U11085 ( .B1(n9777), .B2(n9854), .A(n9776), .ZN(P1_U3275) );
  AOI22_X1 U11086 ( .A1(n9779), .A2(n9984), .B1(n9778), .B2(n9849), .ZN(n9781)
         );
  MUX2_X1 U11087 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9864), .S(n10245), .Z(
        P1_U3552) );
  OAI21_X1 U11088 ( .B1(n4844), .B2(n10226), .A(n9784), .ZN(n9785) );
  NOR2_X1 U11089 ( .A1(n9786), .A2(n9785), .ZN(n9787) );
  OAI21_X1 U11090 ( .B1(n9788), .B2(n9853), .A(n9787), .ZN(n9865) );
  MUX2_X1 U11091 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9865), .S(n10245), .Z(
        P1_U3551) );
  AOI22_X1 U11092 ( .A1(n9790), .A2(n9984), .B1(n9789), .B2(n9849), .ZN(n9791)
         );
  OAI211_X1 U11093 ( .C1(n9793), .C2(n9853), .A(n9792), .B(n9791), .ZN(n9866)
         );
  MUX2_X1 U11094 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9866), .S(n10245), .Z(
        P1_U3550) );
  AOI211_X1 U11095 ( .C1(n9796), .C2(n9849), .A(n9795), .B(n9794), .ZN(n9797)
         );
  OAI21_X1 U11096 ( .B1(n9798), .B2(n9853), .A(n9797), .ZN(n9867) );
  MUX2_X1 U11097 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9867), .S(n10245), .Z(
        P1_U3549) );
  AOI22_X1 U11098 ( .A1(n9800), .A2(n9984), .B1(n9799), .B2(n9849), .ZN(n9801)
         );
  OAI211_X1 U11099 ( .C1(n9803), .C2(n9853), .A(n9802), .B(n9801), .ZN(n9868)
         );
  MUX2_X1 U11100 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9868), .S(n10245), .Z(
        P1_U3548) );
  NAND2_X1 U11101 ( .A1(n9804), .A2(n4761), .ZN(n9810) );
  NOR2_X1 U11102 ( .A1(n9806), .A2(n9805), .ZN(n9809) );
  NAND4_X1 U11103 ( .A1(n9810), .A2(n9809), .A3(n9808), .A4(n9807), .ZN(n9869)
         );
  MUX2_X1 U11104 ( .A(n9869), .B(P1_REG1_REG_24__SCAN_IN), .S(n10243), .Z(
        P1_U3547) );
  AOI22_X1 U11105 ( .A1(n9812), .A2(n9984), .B1(n9811), .B2(n9849), .ZN(n9813)
         );
  OAI211_X1 U11106 ( .C1(n9815), .C2(n9853), .A(n9814), .B(n9813), .ZN(n9870)
         );
  MUX2_X1 U11107 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9870), .S(n10245), .Z(
        P1_U3546) );
  AOI22_X1 U11108 ( .A1(n9817), .A2(n9984), .B1(n9816), .B2(n9849), .ZN(n9818)
         );
  OAI211_X1 U11109 ( .C1(n9820), .C2(n9853), .A(n9819), .B(n9818), .ZN(n9871)
         );
  MUX2_X1 U11110 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9871), .S(n10245), .Z(
        P1_U3545) );
  AOI211_X1 U11111 ( .C1(n9823), .C2(n9849), .A(n9822), .B(n9821), .ZN(n9824)
         );
  OAI21_X1 U11112 ( .B1(n9853), .B2(n9825), .A(n9824), .ZN(n9872) );
  MUX2_X1 U11113 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9872), .S(n10245), .Z(
        P1_U3544) );
  AOI22_X1 U11114 ( .A1(n9827), .A2(n9984), .B1(n9826), .B2(n9849), .ZN(n9828)
         );
  OAI211_X1 U11115 ( .C1(n9830), .C2(n9853), .A(n9829), .B(n9828), .ZN(n9873)
         );
  MUX2_X1 U11116 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9873), .S(n10245), .Z(
        P1_U3543) );
  AOI211_X1 U11117 ( .C1(n9833), .C2(n9849), .A(n9832), .B(n9831), .ZN(n9834)
         );
  OAI21_X1 U11118 ( .B1(n9835), .B2(n9853), .A(n9834), .ZN(n9874) );
  MUX2_X1 U11119 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9874), .S(n10245), .Z(
        P1_U3542) );
  NAND3_X1 U11120 ( .A1(n9837), .A2(n4761), .A3(n9836), .ZN(n9842) );
  AOI22_X1 U11121 ( .A1(n9839), .A2(n9984), .B1(n9838), .B2(n9849), .ZN(n9840)
         );
  NAND3_X1 U11122 ( .A1(n9842), .A2(n9841), .A3(n9840), .ZN(n9875) );
  MUX2_X1 U11123 ( .A(n9875), .B(P1_REG1_REG_18__SCAN_IN), .S(n10243), .Z(
        P1_U3541) );
  AOI211_X1 U11124 ( .C1(n9845), .C2(n9849), .A(n9844), .B(n9843), .ZN(n9846)
         );
  OAI21_X1 U11125 ( .B1(n9847), .B2(n9853), .A(n9846), .ZN(n9876) );
  MUX2_X1 U11126 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9876), .S(n10245), .Z(
        P1_U3540) );
  AOI21_X1 U11127 ( .B1(n9850), .B2(n9849), .A(n9848), .ZN(n9851) );
  OAI211_X1 U11128 ( .C1(n9854), .C2(n9853), .A(n9852), .B(n9851), .ZN(n9877)
         );
  MUX2_X1 U11129 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9877), .S(n10245), .Z(
        P1_U3539) );
  INV_X1 U11130 ( .A(n9855), .ZN(n9863) );
  INV_X1 U11131 ( .A(n9856), .ZN(n9857) );
  OAI22_X1 U11132 ( .A1(n9858), .A2(n10228), .B1(n9857), .B2(n10226), .ZN(
        n9859) );
  INV_X1 U11133 ( .A(n9859), .ZN(n9860) );
  OAI211_X1 U11134 ( .C1(n9863), .C2(n9862), .A(n9861), .B(n9860), .ZN(n9878)
         );
  MUX2_X1 U11135 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9878), .S(n10245), .Z(
        P1_U3538) );
  MUX2_X1 U11136 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9864), .S(n10236), .Z(
        P1_U3520) );
  MUX2_X1 U11137 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9865), .S(n10236), .Z(
        P1_U3519) );
  MUX2_X1 U11138 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n9866), .S(n10236), .Z(
        P1_U3518) );
  MUX2_X1 U11139 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9867), .S(n10236), .Z(
        P1_U3517) );
  MUX2_X1 U11140 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9868), .S(n10236), .Z(
        P1_U3516) );
  MUX2_X1 U11141 ( .A(n9869), .B(P1_REG0_REG_24__SCAN_IN), .S(n10234), .Z(
        P1_U3515) );
  MUX2_X1 U11142 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9870), .S(n10236), .Z(
        P1_U3514) );
  MUX2_X1 U11143 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9871), .S(n10236), .Z(
        P1_U3513) );
  MUX2_X1 U11144 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9872), .S(n10236), .Z(
        P1_U3512) );
  MUX2_X1 U11145 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9873), .S(n10236), .Z(
        P1_U3511) );
  MUX2_X1 U11146 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9874), .S(n10236), .Z(
        P1_U3510) );
  MUX2_X1 U11147 ( .A(n9875), .B(P1_REG0_REG_18__SCAN_IN), .S(n10234), .Z(
        P1_U3508) );
  MUX2_X1 U11148 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9876), .S(n10236), .Z(
        P1_U3505) );
  MUX2_X1 U11149 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9877), .S(n10236), .Z(
        P1_U3502) );
  MUX2_X1 U11150 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9878), .S(n10236), .Z(
        P1_U3499) );
  MUX2_X1 U11151 ( .A(n9880), .B(P1_D_REG_0__SCAN_IN), .S(n9879), .Z(P1_U3440)
         );
  INV_X1 U11152 ( .A(n9881), .ZN(n9884) );
  NOR4_X1 U11153 ( .A1(P1_U3084), .A2(n5900), .A3(P1_IR_REG_29__SCAN_IN), .A4(
        P1_IR_REG_30__SCAN_IN), .ZN(n9883) );
  AOI22_X1 U11154 ( .A1(n9884), .A2(n9883), .B1(P2_DATAO_REG_31__SCAN_IN), 
        .B2(n9882), .ZN(n9885) );
  OAI21_X1 U11155 ( .B1(n9887), .B2(n9886), .A(n9885), .ZN(P1_U3322) );
  NAND2_X1 U11156 ( .A1(n9888), .A2(n9892), .ZN(n9889) );
  OAI211_X1 U11157 ( .C1(n9891), .C2(n9890), .A(n9889), .B(n10011), .ZN(
        P1_U3325) );
  NAND2_X1 U11158 ( .A1(n9893), .A2(n9892), .ZN(n9894) );
  OAI211_X1 U11159 ( .C1(n9891), .C2(n9895), .A(n9894), .B(n10010), .ZN(
        P1_U3326) );
  INV_X1 U11160 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n9898) );
  AND2_X1 U11161 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10278) );
  INV_X1 U11162 ( .A(n10278), .ZN(n9897) );
  OAI21_X1 U11163 ( .B1(n10304), .B2(n9898), .A(n9897), .ZN(n9899) );
  AOI21_X1 U11164 ( .B1(n10330), .B2(n9900), .A(n9899), .ZN(n9909) );
  OAI211_X1 U11165 ( .C1(n9903), .C2(n9902), .A(n9901), .B(n10336), .ZN(n9908)
         );
  OAI211_X1 U11166 ( .C1(n9906), .C2(n9905), .A(n10332), .B(n9904), .ZN(n9907)
         );
  NAND3_X1 U11167 ( .A1(n9909), .A2(n9908), .A3(n9907), .ZN(P2_U3250) );
  AOI22_X1 U11168 ( .A1(n10328), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n9920) );
  NAND2_X1 U11169 ( .A1(n10330), .A2(n9910), .ZN(n9919) );
  OAI211_X1 U11170 ( .C1(n9913), .C2(n9912), .A(n10336), .B(n9911), .ZN(n9918)
         );
  OAI211_X1 U11171 ( .C1(n9916), .C2(n9915), .A(n10332), .B(n9914), .ZN(n9917)
         );
  NAND4_X1 U11172 ( .A1(n9920), .A2(n9919), .A3(n9918), .A4(n9917), .ZN(
        P2_U3247) );
  OAI21_X1 U11173 ( .B1(n9921), .B2(n10226), .A(n9980), .ZN(n9922) );
  AOI21_X1 U11174 ( .B1(n9923), .B2(n9984), .A(n9922), .ZN(n9925) );
  AOI22_X1 U11175 ( .A1(n10245), .A2(n9925), .B1(n6675), .B2(n10243), .ZN(
        P1_U3554) );
  AOI22_X1 U11176 ( .A1(n10236), .A2(n9925), .B1(n9924), .B2(n10234), .ZN(
        P1_U3522) );
  OAI21_X1 U11177 ( .B1(n9928), .B2(n10453), .A(n9927), .ZN(n9930) );
  AOI211_X1 U11178 ( .C1(n10459), .C2(n9931), .A(n9930), .B(n9929), .ZN(n9933)
         );
  AOI22_X1 U11179 ( .A1(n10473), .A2(n9933), .B1(n5356), .B2(n10471), .ZN(
        P2_U3534) );
  AOI22_X1 U11180 ( .A1(n10462), .A2(n9933), .B1(n9932), .B2(n10461), .ZN(
        P2_U3493) );
  XNOR2_X1 U11181 ( .A(n9935), .B(n9934), .ZN(n9988) );
  OR2_X1 U11182 ( .A1(n9936), .A2(n9985), .ZN(n9937) );
  NAND2_X1 U11183 ( .A1(n9938), .A2(n9937), .ZN(n9986) );
  INV_X1 U11184 ( .A(n9986), .ZN(n9939) );
  AOI22_X1 U11185 ( .A1(n9988), .A2(n10164), .B1(n10163), .B2(n9939), .ZN(
        n9959) );
  OAI22_X1 U11186 ( .A1(n10181), .A2(n9941), .B1(n9940), .B2(n10178), .ZN(
        n9955) );
  XNOR2_X1 U11187 ( .A(n9943), .B(n9942), .ZN(n9950) );
  AOI22_X1 U11188 ( .A1(n9947), .A2(n9946), .B1(n9945), .B2(n9944), .ZN(n9948)
         );
  OAI21_X1 U11189 ( .B1(n9950), .B2(n9949), .A(n9948), .ZN(n9951) );
  AOI21_X1 U11190 ( .B1(n9988), .B2(n9952), .A(n9951), .ZN(n9990) );
  NOR2_X1 U11191 ( .A1(n9990), .A2(n9953), .ZN(n9954) );
  AOI211_X1 U11192 ( .C1(n9957), .C2(n9956), .A(n9955), .B(n9954), .ZN(n9958)
         );
  NAND2_X1 U11193 ( .A1(n9959), .A2(n9958), .ZN(P1_U3278) );
  XNOR2_X1 U11194 ( .A(n9961), .B(n9960), .ZN(n9972) );
  INV_X1 U11195 ( .A(n9972), .ZN(n10001) );
  AND2_X1 U11196 ( .A1(n9962), .A2(n9973), .ZN(n9964) );
  OR2_X1 U11197 ( .A1(n9964), .A2(n9963), .ZN(n9998) );
  INV_X1 U11198 ( .A(n9998), .ZN(n9965) );
  AOI22_X1 U11199 ( .A1(n10001), .A2(n10164), .B1(n10163), .B2(n9965), .ZN(
        n9979) );
  XNOR2_X1 U11200 ( .A(n9967), .B(n9966), .ZN(n9970) );
  OAI22_X1 U11201 ( .A1(n10170), .A2(n10168), .B1(n9968), .B2(n10167), .ZN(
        n9969) );
  AOI21_X1 U11202 ( .B1(n9970), .B2(n10172), .A(n9969), .ZN(n9971) );
  OAI21_X1 U11203 ( .B1(n9972), .B2(n10175), .A(n9971), .ZN(n9999) );
  INV_X1 U11204 ( .A(n9973), .ZN(n9997) );
  NOR2_X1 U11205 ( .A1(n9997), .A2(n10177), .ZN(n9977) );
  OAI22_X1 U11206 ( .A1(n10181), .A2(n9975), .B1(n9974), .B2(n10178), .ZN(
        n9976) );
  AOI211_X1 U11207 ( .C1(n9999), .C2(n10181), .A(n9977), .B(n9976), .ZN(n9978)
         );
  NAND2_X1 U11208 ( .A1(n9979), .A2(n9978), .ZN(P1_U3280) );
  OAI21_X1 U11209 ( .B1(n9981), .B2(n10226), .A(n9980), .ZN(n9982) );
  AOI21_X1 U11210 ( .B1(n9984), .B2(n9983), .A(n9982), .ZN(n10004) );
  AOI22_X1 U11211 ( .A1(n10245), .A2(n10004), .B1(n8016), .B2(n10243), .ZN(
        P1_U3553) );
  OAI22_X1 U11212 ( .A1(n9986), .A2(n10228), .B1(n9985), .B2(n10226), .ZN(
        n9987) );
  AOI21_X1 U11213 ( .B1(n9988), .B2(n10233), .A(n9987), .ZN(n9989) );
  AOI22_X1 U11214 ( .A1(n10245), .A2(n10006), .B1(n7104), .B2(n10243), .ZN(
        P1_U3536) );
  INV_X1 U11215 ( .A(n9991), .ZN(n9996) );
  OAI21_X1 U11216 ( .B1(n9993), .B2(n10226), .A(n9992), .ZN(n9995) );
  AOI211_X1 U11217 ( .C1(n10233), .C2(n9996), .A(n9995), .B(n9994), .ZN(n10008) );
  AOI22_X1 U11218 ( .A1(n10245), .A2(n10008), .B1(n7102), .B2(n10243), .ZN(
        P1_U3535) );
  OAI22_X1 U11219 ( .A1(n9998), .A2(n10228), .B1(n9997), .B2(n10226), .ZN(
        n10000) );
  AOI211_X1 U11220 ( .C1(n10233), .C2(n10001), .A(n10000), .B(n9999), .ZN(
        n10009) );
  AOI22_X1 U11221 ( .A1(n10245), .A2(n10009), .B1(n10002), .B2(n10243), .ZN(
        P1_U3534) );
  INV_X1 U11222 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n10003) );
  AOI22_X1 U11223 ( .A1(n10236), .A2(n10004), .B1(n10003), .B2(n10234), .ZN(
        P1_U3521) );
  INV_X1 U11224 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n10005) );
  AOI22_X1 U11225 ( .A1(n10236), .A2(n10006), .B1(n10005), .B2(n10234), .ZN(
        P1_U3493) );
  INV_X1 U11226 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n10007) );
  AOI22_X1 U11227 ( .A1(n10236), .A2(n10008), .B1(n10007), .B2(n10234), .ZN(
        P1_U3490) );
  AOI22_X1 U11228 ( .A1(n10236), .A2(n10009), .B1(n6139), .B2(n10234), .ZN(
        P1_U3487) );
  XNOR2_X1 U11229 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  XNOR2_X1 U11230 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  INV_X1 U11231 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n10017) );
  OAI21_X1 U11232 ( .B1(n10011), .B2(n10019), .A(n10010), .ZN(n10013) );
  OAI211_X1 U11233 ( .C1(n10014), .C2(n4694), .A(n10013), .B(n10012), .ZN(
        n10015) );
  OAI22_X1 U11234 ( .A1(n10157), .A2(n10017), .B1(n10016), .B2(n10015), .ZN(
        n10018) );
  INV_X1 U11235 ( .A(n10018), .ZN(n10021) );
  OAI211_X1 U11236 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n5941), .A(n10021), .B(
        n10020), .ZN(P1_U3241) );
  INV_X1 U11237 ( .A(n10022), .ZN(n10026) );
  INV_X1 U11238 ( .A(n10023), .ZN(n10025) );
  OAI21_X1 U11239 ( .B1(n10026), .B2(n10025), .A(n10024), .ZN(n10029) );
  INV_X1 U11240 ( .A(n10027), .ZN(n10028) );
  AOI22_X1 U11241 ( .A1(n10058), .A2(n10029), .B1(n10028), .B2(n10148), .ZN(
        n10038) );
  AOI21_X1 U11242 ( .B1(n10032), .B2(n10031), .A(n10030), .ZN(n10033) );
  NOR2_X1 U11243 ( .A1(n10154), .A2(n10033), .ZN(n10034) );
  AOI211_X1 U11244 ( .C1(n10052), .C2(P1_ADDR_REG_4__SCAN_IN), .A(n10035), .B(
        n10034), .ZN(n10037) );
  NAND3_X1 U11245 ( .A1(n10038), .A2(n10037), .A3(n10036), .ZN(P1_U3245) );
  AOI22_X1 U11246 ( .A1(n10052), .A2(P1_ADDR_REG_5__SCAN_IN), .B1(n10039), 
        .B2(n10148), .ZN(n10050) );
  OAI21_X1 U11247 ( .B1(n10042), .B2(n10041), .A(n10040), .ZN(n10043) );
  NAND2_X1 U11248 ( .A1(n10058), .A2(n10043), .ZN(n10048) );
  OAI211_X1 U11249 ( .C1(n10046), .C2(n10045), .A(n10135), .B(n10044), .ZN(
        n10047) );
  NAND4_X1 U11250 ( .A1(n10050), .A2(n10049), .A3(n10048), .A4(n10047), .ZN(
        P1_U3246) );
  AOI22_X1 U11251 ( .A1(n10052), .A2(P1_ADDR_REG_8__SCAN_IN), .B1(n10051), 
        .B2(n10148), .ZN(n10065) );
  INV_X1 U11252 ( .A(n10053), .ZN(n10064) );
  OAI21_X1 U11253 ( .B1(n10056), .B2(n10055), .A(n10054), .ZN(n10057) );
  NAND2_X1 U11254 ( .A1(n10058), .A2(n10057), .ZN(n10063) );
  OAI211_X1 U11255 ( .C1(n10061), .C2(n10060), .A(n10135), .B(n10059), .ZN(
        n10062) );
  NAND4_X1 U11256 ( .A1(n10065), .A2(n10064), .A3(n10063), .A4(n10062), .ZN(
        P1_U3249) );
  AOI21_X1 U11257 ( .B1(n10068), .B2(n10067), .A(n10066), .ZN(n10069) );
  NOR2_X1 U11258 ( .A1(n10069), .A2(n10154), .ZN(n10077) );
  AOI211_X1 U11259 ( .C1(n10072), .C2(n10071), .A(n10070), .B(n10142), .ZN(
        n10076) );
  OAI22_X1 U11260 ( .A1(n10074), .A2(n10073), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7513), .ZN(n10075) );
  NOR3_X1 U11261 ( .A1(n10077), .A2(n10076), .A3(n10075), .ZN(n10078) );
  OAI21_X1 U11262 ( .B1(n10514), .B2(n10157), .A(n10078), .ZN(P1_U3250) );
  INV_X1 U11263 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n10091) );
  AOI211_X1 U11264 ( .C1(n10081), .C2(n10080), .A(n10079), .B(n10142), .ZN(
        n10082) );
  AOI211_X1 U11265 ( .C1(n10148), .C2(n10084), .A(n10083), .B(n10082), .ZN(
        n10090) );
  AOI21_X1 U11266 ( .B1(n10087), .B2(n10086), .A(n10085), .ZN(n10088) );
  OR2_X1 U11267 ( .A1(n10088), .A2(n10154), .ZN(n10089) );
  OAI211_X1 U11268 ( .C1(n10091), .C2(n10157), .A(n10090), .B(n10089), .ZN(
        P1_U3253) );
  INV_X1 U11269 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n10104) );
  AOI211_X1 U11270 ( .C1(n10094), .C2(n10093), .A(n10092), .B(n10142), .ZN(
        n10095) );
  AOI211_X1 U11271 ( .C1(n10148), .C2(n10097), .A(n10096), .B(n10095), .ZN(
        n10103) );
  AOI21_X1 U11272 ( .B1(n10100), .B2(n10099), .A(n10098), .ZN(n10101) );
  OR2_X1 U11273 ( .A1(n10154), .A2(n10101), .ZN(n10102) );
  OAI211_X1 U11274 ( .C1(n10104), .C2(n10157), .A(n10103), .B(n10102), .ZN(
        P1_U3254) );
  INV_X1 U11275 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10114) );
  AOI211_X1 U11276 ( .C1(n7901), .C2(n10106), .A(n10142), .B(n10105), .ZN(
        n10107) );
  AOI211_X1 U11277 ( .C1(n10109), .C2(n10148), .A(n10108), .B(n10107), .ZN(
        n10113) );
  XNOR2_X1 U11278 ( .A(n10110), .B(P1_REG1_REG_15__SCAN_IN), .ZN(n10111) );
  NAND2_X1 U11279 ( .A1(n10111), .A2(n10135), .ZN(n10112) );
  OAI211_X1 U11280 ( .C1(n10114), .C2(n10157), .A(n10113), .B(n10112), .ZN(
        P1_U3256) );
  INV_X1 U11281 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n10126) );
  AOI211_X1 U11282 ( .C1(n10117), .C2(n10116), .A(n10115), .B(n10142), .ZN(
        n10118) );
  AOI211_X1 U11283 ( .C1(n10120), .C2(n10148), .A(n10119), .B(n10118), .ZN(
        n10125) );
  OAI211_X1 U11284 ( .C1(n10123), .C2(n10122), .A(n10135), .B(n10121), .ZN(
        n10124) );
  OAI211_X1 U11285 ( .C1(n10126), .C2(n10157), .A(n10125), .B(n10124), .ZN(
        P1_U3257) );
  INV_X1 U11286 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n10140) );
  INV_X1 U11287 ( .A(n10127), .ZN(n10132) );
  AOI211_X1 U11288 ( .C1(n10130), .C2(n10129), .A(n10128), .B(n10142), .ZN(
        n10131) );
  AOI211_X1 U11289 ( .C1(n10133), .C2(n10148), .A(n10132), .B(n10131), .ZN(
        n10139) );
  OAI211_X1 U11290 ( .C1(n10137), .C2(n10136), .A(n10135), .B(n10134), .ZN(
        n10138) );
  OAI211_X1 U11291 ( .C1(n10140), .C2(n10157), .A(n10139), .B(n10138), .ZN(
        P1_U3258) );
  INV_X1 U11292 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10158) );
  INV_X1 U11293 ( .A(n10141), .ZN(n10147) );
  AOI211_X1 U11294 ( .C1(n10145), .C2(n10144), .A(n10143), .B(n10142), .ZN(
        n10146) );
  AOI211_X1 U11295 ( .C1(n10149), .C2(n10148), .A(n10147), .B(n10146), .ZN(
        n10156) );
  AOI21_X1 U11296 ( .B1(n10152), .B2(n10151), .A(n10150), .ZN(n10153) );
  OR2_X1 U11297 ( .A1(n10154), .A2(n10153), .ZN(n10155) );
  OAI211_X1 U11298 ( .C1(n10158), .C2(n10157), .A(n10156), .B(n10155), .ZN(
        P1_U3259) );
  XOR2_X1 U11299 ( .A(n10159), .B(n10166), .Z(n10176) );
  INV_X1 U11300 ( .A(n10176), .ZN(n10232) );
  OAI21_X1 U11301 ( .B1(n10161), .B2(n10227), .A(n10160), .ZN(n10229) );
  INV_X1 U11302 ( .A(n10229), .ZN(n10162) );
  AOI22_X1 U11303 ( .A1(n10232), .A2(n10164), .B1(n10163), .B2(n10162), .ZN(
        n10185) );
  XOR2_X1 U11304 ( .A(n10166), .B(n10165), .Z(n10173) );
  OAI22_X1 U11305 ( .A1(n10170), .A2(n10169), .B1(n10168), .B2(n10167), .ZN(
        n10171) );
  AOI21_X1 U11306 ( .B1(n10173), .B2(n10172), .A(n10171), .ZN(n10174) );
  OAI21_X1 U11307 ( .B1(n10176), .B2(n10175), .A(n10174), .ZN(n10230) );
  NOR2_X1 U11308 ( .A1(n10227), .A2(n10177), .ZN(n10183) );
  OAI22_X1 U11309 ( .A1(n10181), .A2(n10180), .B1(n10179), .B2(n10178), .ZN(
        n10182) );
  AOI211_X1 U11310 ( .C1(n10230), .C2(n10181), .A(n10183), .B(n10182), .ZN(
        n10184) );
  NAND2_X1 U11311 ( .A1(n10185), .A2(n10184), .ZN(P1_U3282) );
  AND2_X1 U11312 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10193), .ZN(P1_U3292) );
  AND2_X1 U11313 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10193), .ZN(P1_U3293) );
  NOR2_X1 U11314 ( .A1(n10192), .A2(n10186), .ZN(P1_U3294) );
  AND2_X1 U11315 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10193), .ZN(P1_U3295) );
  AND2_X1 U11316 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10193), .ZN(P1_U3296) );
  AND2_X1 U11317 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10193), .ZN(P1_U3297) );
  AND2_X1 U11318 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10193), .ZN(P1_U3298) );
  AND2_X1 U11319 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10193), .ZN(P1_U3299) );
  NOR2_X1 U11320 ( .A1(n10192), .A2(n10187), .ZN(P1_U3300) );
  AND2_X1 U11321 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10193), .ZN(P1_U3301) );
  AND2_X1 U11322 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10193), .ZN(P1_U3302) );
  AND2_X1 U11323 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10193), .ZN(P1_U3303) );
  AND2_X1 U11324 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10193), .ZN(P1_U3304) );
  AND2_X1 U11325 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10193), .ZN(P1_U3305) );
  NOR2_X1 U11326 ( .A1(n10192), .A2(n10188), .ZN(P1_U3306) );
  AND2_X1 U11327 ( .A1(n10193), .A2(P1_D_REG_16__SCAN_IN), .ZN(P1_U3307) );
  AND2_X1 U11328 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10193), .ZN(P1_U3308) );
  AND2_X1 U11329 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10193), .ZN(P1_U3309) );
  AND2_X1 U11330 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10193), .ZN(P1_U3310) );
  NOR2_X1 U11331 ( .A1(n10192), .A2(n10189), .ZN(P1_U3311) );
  AND2_X1 U11332 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10193), .ZN(P1_U3312) );
  AND2_X1 U11333 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10193), .ZN(P1_U3313) );
  AND2_X1 U11334 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10193), .ZN(P1_U3314) );
  AND2_X1 U11335 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10193), .ZN(P1_U3315) );
  AND2_X1 U11336 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10193), .ZN(P1_U3316) );
  AND2_X1 U11337 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10193), .ZN(P1_U3317) );
  AND2_X1 U11338 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10193), .ZN(P1_U3318) );
  NOR2_X1 U11339 ( .A1(n10192), .A2(n10190), .ZN(P1_U3319) );
  NOR2_X1 U11340 ( .A1(n10192), .A2(n10191), .ZN(P1_U3320) );
  AND2_X1 U11341 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10193), .ZN(P1_U3321) );
  INV_X1 U11342 ( .A(n10194), .ZN(n10199) );
  OAI21_X1 U11343 ( .B1(n10226), .B2(n10196), .A(n10195), .ZN(n10198) );
  AOI211_X1 U11344 ( .C1(n10233), .C2(n10199), .A(n10198), .B(n10197), .ZN(
        n10237) );
  INV_X1 U11345 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10200) );
  AOI22_X1 U11346 ( .A1(n10236), .A2(n10237), .B1(n10200), .B2(n10234), .ZN(
        P1_U3457) );
  OAI22_X1 U11347 ( .A1(n10202), .A2(n10228), .B1(n10201), .B2(n10226), .ZN(
        n10204) );
  AOI211_X1 U11348 ( .C1(n10233), .C2(n10205), .A(n10204), .B(n10203), .ZN(
        n10238) );
  AOI22_X1 U11349 ( .A1(n10236), .A2(n10238), .B1(n5919), .B2(n10234), .ZN(
        P1_U3463) );
  OAI21_X1 U11350 ( .B1(n10207), .B2(n10226), .A(n10206), .ZN(n10208) );
  AOI21_X1 U11351 ( .B1(n10209), .B2(n4761), .A(n10208), .ZN(n10211) );
  AND2_X1 U11352 ( .A1(n10211), .A2(n10210), .ZN(n10239) );
  INV_X1 U11353 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U11354 ( .A1(n10236), .A2(n10239), .B1(n10212), .B2(n10234), .ZN(
        P1_U3469) );
  OAI21_X1 U11355 ( .B1(n10214), .B2(n10226), .A(n10213), .ZN(n10216) );
  AOI211_X1 U11356 ( .C1(n4761), .C2(n10217), .A(n10216), .B(n10215), .ZN(
        n10240) );
  INV_X1 U11357 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n10218) );
  AOI22_X1 U11358 ( .A1(n10236), .A2(n10240), .B1(n10218), .B2(n10234), .ZN(
        P1_U3475) );
  INV_X1 U11359 ( .A(n10219), .ZN(n10224) );
  OAI22_X1 U11360 ( .A1(n10221), .A2(n10228), .B1(n10220), .B2(n10226), .ZN(
        n10223) );
  AOI211_X1 U11361 ( .C1(n10233), .C2(n10224), .A(n10223), .B(n10222), .ZN(
        n10242) );
  INV_X1 U11362 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n10225) );
  AOI22_X1 U11363 ( .A1(n10236), .A2(n10242), .B1(n10225), .B2(n10234), .ZN(
        P1_U3478) );
  OAI22_X1 U11364 ( .A1(n10229), .A2(n10228), .B1(n10227), .B2(n10226), .ZN(
        n10231) );
  AOI211_X1 U11365 ( .C1(n10233), .C2(n10232), .A(n10231), .B(n10230), .ZN(
        n10244) );
  INV_X1 U11366 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10235) );
  AOI22_X1 U11367 ( .A1(n10236), .A2(n10244), .B1(n10235), .B2(n10234), .ZN(
        P1_U3481) );
  AOI22_X1 U11368 ( .A1(n10245), .A2(n10237), .B1(n6689), .B2(n10243), .ZN(
        P1_U3524) );
  AOI22_X1 U11369 ( .A1(n10245), .A2(n10238), .B1(n6694), .B2(n10243), .ZN(
        P1_U3526) );
  AOI22_X1 U11370 ( .A1(n10245), .A2(n10239), .B1(n6688), .B2(n10243), .ZN(
        P1_U3528) );
  AOI22_X1 U11371 ( .A1(n10245), .A2(n10240), .B1(n6051), .B2(n10243), .ZN(
        P1_U3530) );
  AOI22_X1 U11372 ( .A1(n10245), .A2(n10242), .B1(n10241), .B2(n10243), .ZN(
        P1_U3531) );
  AOI22_X1 U11373 ( .A1(n10245), .A2(n10244), .B1(n6094), .B2(n10243), .ZN(
        P1_U3532) );
  AOI211_X1 U11374 ( .C1(n10248), .C2(n10247), .A(n10246), .B(n4513), .ZN(
        n10255) );
  INV_X1 U11375 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n10249) );
  NOR2_X1 U11376 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10249), .ZN(n10301) );
  NOR2_X1 U11377 ( .A1(n4871), .A2(n10250), .ZN(n10254) );
  OAI22_X1 U11378 ( .A1(n10252), .A2(n10251), .B1(n4786), .B2(n10260), .ZN(
        n10253) );
  NOR4_X1 U11379 ( .A1(n10255), .A2(n10301), .A3(n10254), .A4(n10253), .ZN(
        n10256) );
  OAI21_X1 U11380 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n10292), .A(n10256), .ZN(
        P2_U3220) );
  NAND2_X1 U11381 ( .A1(n10257), .A2(n10262), .ZN(n10259) );
  OAI211_X1 U11382 ( .C1(n10261), .C2(n10260), .A(n10259), .B(n10258), .ZN(
        n10273) );
  NAND3_X1 U11383 ( .A1(n10264), .A2(n10263), .A3(n10262), .ZN(n10271) );
  INV_X1 U11384 ( .A(n10265), .ZN(n10267) );
  OAI21_X1 U11385 ( .B1(n10267), .B2(n10266), .A(n10287), .ZN(n10270) );
  INV_X1 U11386 ( .A(n10268), .ZN(n10269) );
  AOI21_X1 U11387 ( .B1(n10271), .B2(n10270), .A(n10269), .ZN(n10272) );
  AOI211_X1 U11388 ( .C1(n10286), .C2(n10274), .A(n10273), .B(n10272), .ZN(
        n10275) );
  OAI21_X1 U11389 ( .B1(n10292), .B2(n10276), .A(n10275), .ZN(P2_U3226) );
  INV_X1 U11390 ( .A(n10277), .ZN(n10280) );
  AOI21_X1 U11391 ( .B1(n10280), .B2(n10279), .A(n10278), .ZN(n10290) );
  NAND2_X1 U11392 ( .A1(n10282), .A2(n10281), .ZN(n10284) );
  XOR2_X1 U11393 ( .A(n10284), .B(n10283), .Z(n10288) );
  AOI22_X1 U11394 ( .A1(n10288), .A2(n10287), .B1(n10286), .B2(n10285), .ZN(
        n10289) );
  OAI211_X1 U11395 ( .C1(n10292), .C2(n10291), .A(n10290), .B(n10289), .ZN(
        P2_U3229) );
  AOI22_X1 U11396 ( .A1(n10332), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10336), .ZN(n10300) );
  AOI22_X1 U11397 ( .A1(n10328), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10299) );
  OAI21_X1 U11398 ( .B1(P2_REG1_REG_0__SCAN_IN), .B2(n10294), .A(n10293), .ZN(
        n10297) );
  NOR2_X1 U11399 ( .A1(n10295), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10296) );
  OAI21_X1 U11400 ( .B1(n10297), .B2(n10296), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n10298) );
  OAI211_X1 U11401 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10300), .A(n10299), .B(
        n10298), .ZN(P2_U3245) );
  INV_X1 U11402 ( .A(n10301), .ZN(n10302) );
  OAI21_X1 U11403 ( .B1(n10304), .B2(n10303), .A(n10302), .ZN(n10305) );
  AOI21_X1 U11404 ( .B1(n10330), .B2(n10306), .A(n10305), .ZN(n10315) );
  OAI211_X1 U11405 ( .C1(n10309), .C2(n10308), .A(n10336), .B(n10307), .ZN(
        n10314) );
  OAI211_X1 U11406 ( .C1(n10312), .C2(n10311), .A(n10332), .B(n10310), .ZN(
        n10313) );
  NAND3_X1 U11407 ( .A1(n10315), .A2(n10314), .A3(n10313), .ZN(P2_U3248) );
  AOI22_X1 U11408 ( .A1(n10328), .A2(P2_ADDR_REG_7__SCAN_IN), .B1(
        P2_REG3_REG_7__SCAN_IN), .B2(P2_U3152), .ZN(n10326) );
  NAND2_X1 U11409 ( .A1(n10330), .A2(n10316), .ZN(n10325) );
  OAI211_X1 U11410 ( .C1(n10319), .C2(n10318), .A(n10317), .B(n10336), .ZN(
        n10324) );
  OAI211_X1 U11411 ( .C1(n10322), .C2(n10321), .A(n10332), .B(n10320), .ZN(
        n10323) );
  NAND4_X1 U11412 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        P2_U3252) );
  AOI21_X1 U11413 ( .B1(n10328), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n10327), 
        .ZN(n10342) );
  NAND2_X1 U11414 ( .A1(n10330), .A2(n10329), .ZN(n10341) );
  OAI211_X1 U11415 ( .C1(n10334), .C2(n10333), .A(n10332), .B(n10331), .ZN(
        n10340) );
  OAI211_X1 U11416 ( .C1(n10338), .C2(n10337), .A(n10336), .B(n10335), .ZN(
        n10339) );
  NAND4_X1 U11417 ( .A1(n10342), .A2(n10341), .A3(n10340), .A4(n10339), .ZN(
        P2_U3255) );
  XNOR2_X1 U11418 ( .A(n10344), .B(n10343), .ZN(n10352) );
  NAND2_X1 U11419 ( .A1(n10346), .A2(n10347), .ZN(n10348) );
  NAND2_X1 U11420 ( .A1(n10345), .A2(n10348), .ZN(n10429) );
  NOR2_X1 U11421 ( .A1(n10429), .A2(n10349), .ZN(n10350) );
  AOI211_X1 U11422 ( .C1(n10352), .C2(n10371), .A(n10351), .B(n10350), .ZN(
        n10432) );
  INV_X1 U11423 ( .A(n10353), .ZN(n10354) );
  AOI222_X1 U11424 ( .A1(n10356), .A2(n10355), .B1(P2_REG2_REG_8__SCAN_IN), 
        .B2(n10372), .C1(n10373), .C2(n10354), .ZN(n10363) );
  OAI211_X1 U11425 ( .C1(n10358), .C2(n10431), .A(n10447), .B(n10357), .ZN(
        n10430) );
  OAI22_X1 U11426 ( .A1(n10429), .A2(n10360), .B1(n10359), .B2(n10430), .ZN(
        n10361) );
  INV_X1 U11427 ( .A(n10361), .ZN(n10362) );
  OAI211_X1 U11428 ( .C1(n10372), .C2(n10432), .A(n10363), .B(n10362), .ZN(
        P2_U3288) );
  OAI21_X1 U11429 ( .B1(n10375), .B2(n10365), .A(n10364), .ZN(n10370) );
  AOI222_X1 U11430 ( .A1(n10371), .A2(n10370), .B1(n10369), .B2(n10368), .C1(
        n10367), .C2(n10366), .ZN(n10419) );
  AOI22_X1 U11431 ( .A1(n10374), .A2(n10373), .B1(P2_REG2_REG_6__SCAN_IN), 
        .B2(n10372), .ZN(n10383) );
  XNOR2_X1 U11432 ( .A(n10376), .B(n10375), .ZN(n10422) );
  OAI211_X1 U11433 ( .C1(n4571), .C2(n10379), .A(n10447), .B(n10377), .ZN(
        n10378) );
  OAI21_X1 U11434 ( .B1(n10379), .B2(n10453), .A(n10378), .ZN(n10421) );
  AOI22_X1 U11435 ( .A1(n10422), .A2(n10381), .B1(n10380), .B2(n10421), .ZN(
        n10382) );
  OAI211_X1 U11436 ( .C1(n10372), .C2(n10419), .A(n10383), .B(n10382), .ZN(
        P2_U3290) );
  NOR2_X1 U11437 ( .A1(n10395), .A2(n10386), .ZN(P2_U3297) );
  NOR2_X1 U11438 ( .A1(n10395), .A2(n10387), .ZN(P2_U3298) );
  AND2_X1 U11439 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10398), .ZN(P2_U3299) );
  AND2_X1 U11440 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10398), .ZN(P2_U3300) );
  NOR2_X1 U11441 ( .A1(n10395), .A2(n10388), .ZN(P2_U3301) );
  AND2_X1 U11442 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10398), .ZN(P2_U3302) );
  AND2_X1 U11443 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10398), .ZN(P2_U3303) );
  AND2_X1 U11444 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10398), .ZN(P2_U3304) );
  NOR2_X1 U11445 ( .A1(n10395), .A2(n10389), .ZN(P2_U3305) );
  AND2_X1 U11446 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10398), .ZN(P2_U3306) );
  AND2_X1 U11447 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10398), .ZN(P2_U3307) );
  AND2_X1 U11448 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10398), .ZN(P2_U3308) );
  AND2_X1 U11449 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10398), .ZN(P2_U3309) );
  AND2_X1 U11450 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10398), .ZN(P2_U3310) );
  NOR2_X1 U11451 ( .A1(n10395), .A2(n10390), .ZN(P2_U3311) );
  AND2_X1 U11452 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10398), .ZN(P2_U3312) );
  NOR2_X1 U11453 ( .A1(n10395), .A2(n10391), .ZN(P2_U3313) );
  AND2_X1 U11454 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10398), .ZN(P2_U3314) );
  NOR2_X1 U11455 ( .A1(n10395), .A2(n10392), .ZN(P2_U3315) );
  AND2_X1 U11456 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10398), .ZN(P2_U3316) );
  AND2_X1 U11457 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10398), .ZN(P2_U3317) );
  NOR2_X1 U11458 ( .A1(n10395), .A2(n10393), .ZN(P2_U3318) );
  AND2_X1 U11459 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10398), .ZN(P2_U3319) );
  NOR2_X1 U11460 ( .A1(n10395), .A2(n10394), .ZN(P2_U3320) );
  AND2_X1 U11461 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10398), .ZN(P2_U3321) );
  AND2_X1 U11462 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10398), .ZN(P2_U3322) );
  AND2_X1 U11463 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10398), .ZN(P2_U3323) );
  AND2_X1 U11464 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10398), .ZN(P2_U3324) );
  AND2_X1 U11465 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10398), .ZN(P2_U3325) );
  AND2_X1 U11466 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10398), .ZN(P2_U3326) );
  AOI22_X1 U11467 ( .A1(n10397), .A2(n10400), .B1(n10396), .B2(n10398), .ZN(
        P2_U3437) );
  AOI22_X1 U11468 ( .A1(n10401), .A2(n10400), .B1(n10399), .B2(n10398), .ZN(
        P2_U3438) );
  OAI21_X1 U11469 ( .B1(n10404), .B2(n10403), .A(n10402), .ZN(n10405) );
  AOI21_X1 U11470 ( .B1(n10406), .B2(n10459), .A(n10405), .ZN(n10463) );
  AOI22_X1 U11471 ( .A1(n10462), .A2(n10463), .B1(n5127), .B2(n10461), .ZN(
        P2_U3451) );
  OAI21_X1 U11472 ( .B1(n10408), .B2(n10453), .A(n10407), .ZN(n10410) );
  AOI211_X1 U11473 ( .C1(n10459), .C2(n10411), .A(n10410), .B(n10409), .ZN(
        n10464) );
  INV_X1 U11474 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10412) );
  AOI22_X1 U11475 ( .A1(n10462), .A2(n10464), .B1(n10412), .B2(n10461), .ZN(
        P2_U3457) );
  OAI21_X1 U11476 ( .B1(n10414), .B2(n10453), .A(n10413), .ZN(n10416) );
  AOI211_X1 U11477 ( .C1(n10459), .C2(n10417), .A(n10416), .B(n10415), .ZN(
        n10465) );
  INV_X1 U11478 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10418) );
  AOI22_X1 U11479 ( .A1(n10462), .A2(n10465), .B1(n10418), .B2(n10461), .ZN(
        P2_U3463) );
  INV_X1 U11480 ( .A(n10419), .ZN(n10420) );
  AOI211_X1 U11481 ( .C1(n10422), .C2(n10459), .A(n10421), .B(n10420), .ZN(
        n10466) );
  INV_X1 U11482 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10423) );
  AOI22_X1 U11483 ( .A1(n10462), .A2(n10466), .B1(n10423), .B2(n10461), .ZN(
        P2_U3469) );
  AOI211_X1 U11484 ( .C1(n10459), .C2(n10426), .A(n10425), .B(n10424), .ZN(
        n10467) );
  INV_X1 U11485 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10427) );
  AOI22_X1 U11486 ( .A1(n10462), .A2(n10467), .B1(n10427), .B2(n10461), .ZN(
        P2_U3472) );
  INV_X1 U11487 ( .A(n10428), .ZN(n10440) );
  INV_X1 U11488 ( .A(n10429), .ZN(n10435) );
  OAI21_X1 U11489 ( .B1(n10431), .B2(n10453), .A(n10430), .ZN(n10434) );
  INV_X1 U11490 ( .A(n10432), .ZN(n10433) );
  AOI211_X1 U11491 ( .C1(n10440), .C2(n10435), .A(n10434), .B(n10433), .ZN(
        n10468) );
  AOI22_X1 U11492 ( .A1(n10462), .A2(n10468), .B1(n5243), .B2(n10461), .ZN(
        P2_U3475) );
  INV_X1 U11493 ( .A(n10436), .ZN(n10437) );
  OAI22_X1 U11494 ( .A1(n10438), .A2(n10455), .B1(n10437), .B2(n10453), .ZN(
        n10439) );
  AOI21_X1 U11495 ( .B1(n10441), .B2(n10440), .A(n10439), .ZN(n10442) );
  AND2_X1 U11496 ( .A1(n10443), .A2(n10442), .ZN(n10469) );
  AOI22_X1 U11497 ( .A1(n10462), .A2(n10469), .B1(n5260), .B2(n10461), .ZN(
        P2_U3478) );
  NAND2_X1 U11498 ( .A1(n10445), .A2(n10444), .ZN(n10451) );
  NAND3_X1 U11499 ( .A1(n7738), .A2(n10446), .A3(n10459), .ZN(n10450) );
  NAND2_X1 U11500 ( .A1(n10448), .A2(n10447), .ZN(n10449) );
  AOI22_X1 U11501 ( .A1(n10462), .A2(n10470), .B1(n5277), .B2(n10461), .ZN(
        P2_U3481) );
  OAI22_X1 U11502 ( .A1(n10456), .A2(n10455), .B1(n10454), .B2(n10453), .ZN(
        n10458) );
  AOI211_X1 U11503 ( .C1(n10460), .C2(n10459), .A(n10458), .B(n10457), .ZN(
        n10472) );
  AOI22_X1 U11504 ( .A1(n10462), .A2(n10472), .B1(n5317), .B2(n10461), .ZN(
        P2_U3487) );
  AOI22_X1 U11505 ( .A1(n10473), .A2(n10463), .B1(n6771), .B2(n10471), .ZN(
        P2_U3520) );
  AOI22_X1 U11506 ( .A1(n10473), .A2(n10464), .B1(n6773), .B2(n10471), .ZN(
        P2_U3522) );
  AOI22_X1 U11507 ( .A1(n10473), .A2(n10465), .B1(n6777), .B2(n10471), .ZN(
        P2_U3524) );
  AOI22_X1 U11508 ( .A1(n10473), .A2(n10466), .B1(n6779), .B2(n10471), .ZN(
        P2_U3526) );
  AOI22_X1 U11509 ( .A1(n10473), .A2(n10467), .B1(n6805), .B2(n10471), .ZN(
        P2_U3527) );
  AOI22_X1 U11510 ( .A1(n10473), .A2(n10468), .B1(n6804), .B2(n10471), .ZN(
        P2_U3528) );
  AOI22_X1 U11511 ( .A1(n10473), .A2(n10469), .B1(n6808), .B2(n10471), .ZN(
        P2_U3529) );
  AOI22_X1 U11512 ( .A1(n10473), .A2(n10470), .B1(n6997), .B2(n10471), .ZN(
        P2_U3530) );
  AOI22_X1 U11513 ( .A1(n10473), .A2(n10472), .B1(n7069), .B2(n10471), .ZN(
        P2_U3532) );
  INV_X1 U11514 ( .A(n10474), .ZN(n10475) );
  NAND2_X1 U11515 ( .A1(n10476), .A2(n10475), .ZN(n10477) );
  XNOR2_X1 U11516 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10477), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11517 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11518 ( .B1(n10480), .B2(n10479), .A(n10478), .ZN(ADD_1071_U56) );
  OAI21_X1 U11519 ( .B1(n10483), .B2(n10482), .A(n10481), .ZN(ADD_1071_U57) );
  OAI21_X1 U11520 ( .B1(n10486), .B2(n10485), .A(n10484), .ZN(ADD_1071_U58) );
  OAI21_X1 U11521 ( .B1(n10489), .B2(n10488), .A(n10487), .ZN(ADD_1071_U59) );
  OAI21_X1 U11522 ( .B1(n10492), .B2(n10491), .A(n10490), .ZN(ADD_1071_U60) );
  OAI21_X1 U11523 ( .B1(n10495), .B2(n10494), .A(n10493), .ZN(ADD_1071_U61) );
  AOI21_X1 U11524 ( .B1(n10498), .B2(n10497), .A(n10496), .ZN(ADD_1071_U62) );
  AOI21_X1 U11525 ( .B1(n10501), .B2(n10500), .A(n10499), .ZN(ADD_1071_U63) );
  XOR2_X1 U11526 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10502), .Z(ADD_1071_U50) );
  XOR2_X1 U11527 ( .A(n10504), .B(n10503), .Z(ADD_1071_U54) );
  NOR2_X1 U11528 ( .A1(n10506), .A2(n10505), .ZN(n10507) );
  XOR2_X1 U11529 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10507), .Z(ADD_1071_U51) );
  OAI21_X1 U11530 ( .B1(n10510), .B2(n10509), .A(n10508), .ZN(n10511) );
  XNOR2_X1 U11531 ( .A(n10511), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11532 ( .B1(n10514), .B2(n10513), .A(n10512), .ZN(ADD_1071_U47) );
  XOR2_X1 U11533 ( .A(n10515), .B(P2_ADDR_REG_7__SCAN_IN), .Z(ADD_1071_U49) );
  XOR2_X1 U11534 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10516), .Z(ADD_1071_U48) );
  XOR2_X1 U11535 ( .A(n10518), .B(n10517), .Z(ADD_1071_U53) );
  XNOR2_X1 U11536 ( .A(n10520), .B(n10519), .ZN(ADD_1071_U52) );
  INV_X1 U4997 ( .A(n8011), .ZN(n6123) );
  CLKBUF_X1 U5004 ( .A(n6566), .Z(n8343) );
  CLKBUF_X1 U5166 ( .A(n6524), .Z(n4498) );
endmodule

