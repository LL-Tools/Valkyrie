

module b15_C_SARLock_k_128_10 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006;

  BUF_X2 U3569 ( .A(n3349), .Z(n3439) );
  CLKBUF_X2 U3570 ( .A(n3246), .Z(n4134) );
  BUF_X1 U3571 ( .A(n3354), .Z(n4055) );
  CLKBUF_X2 U3572 ( .A(n3433), .Z(n3120) );
  CLKBUF_X2 U3573 ( .A(n3347), .Z(n5301) );
  CLKBUF_X2 U3574 ( .A(n4137), .Z(n4113) );
  CLKBUF_X2 U3575 ( .A(n3298), .Z(n4081) );
  CLKBUF_X2 U3576 ( .A(n3438), .Z(n4135) );
  CLKBUF_X2 U3577 ( .A(n3392), .Z(n4138) );
  CLKBUF_X2 U3578 ( .A(n3297), .Z(n4106) );
  CLKBUF_X2 U3579 ( .A(n4136), .Z(n4086) );
  AND4_X1 U3580 ( .A1(n3241), .A2(n3240), .A3(n3239), .A4(n3238), .ZN(n3253)
         );
  AND4_X1 U3581 ( .A1(n3245), .A2(n3244), .A3(n3243), .A4(n3242), .ZN(n3252)
         );
  AND4_X1 U3582 ( .A1(n3229), .A2(n3228), .A3(n3227), .A4(n3226), .ZN(n3230)
         );
  AND4_X1 U3583 ( .A1(n3180), .A2(n3179), .A3(n3178), .A4(n3177), .ZN(n3141)
         );
  AND4_X1 U3584 ( .A1(n3172), .A2(n3171), .A3(n3170), .A4(n3169), .ZN(n3143)
         );
  AND4_X1 U3585 ( .A1(n3156), .A2(n3155), .A3(n3154), .A4(n3153), .ZN(n3164)
         );
  AND2_X2 U3586 ( .A1(n5300), .A2(n5309), .ZN(n4136) );
  AOI22_X1 U3587 ( .A1(n6977), .A2(keyinput45), .B1(n5802), .B2(keyinput77), 
        .ZN(n6976) );
  CLKBUF_X2 U3588 ( .A(n3356), .Z(n3121) );
  NOR2_X2 U3589 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3157) );
  OAI221_X1 U3590 ( .B1(n6977), .B2(keyinput45), .C1(n5802), .C2(keyinput77), 
        .A(n6976), .ZN(n6986) );
  OAI22_X1 U3591 ( .A1(n6915), .A2(keyinput1), .B1(n6914), .B2(keyinput96), 
        .ZN(n6913) );
  AOI221_X1 U3592 ( .B1(n6915), .B2(keyinput1), .C1(keyinput96), .C2(n6914), 
        .A(n6913), .ZN(n6928) );
  INV_X1 U3593 ( .A(n4282), .ZN(n4291) );
  MUX2_X1 U3595 ( .A(n4291), .B(n4290), .S(EBX_REG_2__SCAN_IN), .Z(n4212) );
  INV_X1 U3596 ( .A(n4200), .ZN(n5444) );
  INV_X2 U3597 ( .A(n5207), .ZN(n5330) );
  INV_X1 U3598 ( .A(n3552), .ZN(n3556) );
  AND4_X1 U3600 ( .A1(n3250), .A2(n3249), .A3(n3248), .A4(n3247), .ZN(n3251)
         );
  INV_X1 U3601 ( .A(n6193), .ZN(n6203) );
  AND2_X1 U3602 ( .A1(n6073), .A2(n4157), .ZN(n6341) );
  INV_X1 U3603 ( .A(n6258), .ZN(n6254) );
  INV_X2 U3604 ( .A(n4585), .ZN(n3271) );
  NAND2_X2 U3605 ( .A1(n3426), .A2(n3425), .ZN(n4544) );
  INV_X2 U3606 ( .A(n5373), .ZN(n5607) );
  OAI21_X2 U3607 ( .B1(n3663), .B2(n3622), .A(n3454), .ZN(n3456) );
  OAI21_X2 U3608 ( .B1(n5558), .B2(n3561), .A(n3560), .ZN(n5571) );
  CLKBUF_X1 U3609 ( .A(n4485), .Z(n4495) );
  INV_X4 U3610 ( .A(n3556), .ZN(n3119) );
  NAND2_X1 U3611 ( .A1(n6663), .A2(n6480), .ZN(n6477) );
  AOI21_X1 U3612 ( .B1(n4165), .B2(n6329), .A(n4164), .ZN(n4166) );
  NAND4_X1 U3613 ( .A1(n5514), .A2(n5623), .A3(n3556), .A4(n5512), .ZN(n5489)
         );
  NAND2_X1 U3614 ( .A1(n5545), .A2(n5546), .ZN(n5544) );
  NAND2_X1 U3615 ( .A1(n4154), .A2(n4155), .ZN(n4346) );
  CLKBUF_X1 U3616 ( .A(n5689), .Z(n3127) );
  NAND2_X1 U3617 ( .A1(n5409), .A2(n5400), .ZN(n5402) );
  OR2_X1 U3618 ( .A1(n5085), .A2(n3549), .ZN(n3551) );
  NAND2_X1 U3619 ( .A1(n3548), .A2(n3547), .ZN(n5085) );
  INV_X1 U3620 ( .A(n5101), .ZN(n3847) );
  OR2_X2 U3621 ( .A1(n5414), .A2(n5403), .ZN(n5405) );
  AND2_X1 U3622 ( .A1(n5222), .A2(n3555), .ZN(n3125) );
  NOR2_X1 U3623 ( .A1(n4754), .A2(n5735), .ZN(n4778) );
  AOI21_X1 U3624 ( .B1(n3780), .B2(n4905), .A(n3788), .ZN(n4486) );
  NOR2_X2 U3625 ( .A1(n5244), .A2(n5243), .ZN(n6030) );
  NAND2_X1 U3626 ( .A1(n3662), .A2(n3661), .ZN(n4391) );
  OR2_X1 U3627 ( .A1(n3659), .A2(n3660), .ZN(n4399) );
  NOR2_X2 U3628 ( .A1(n5712), .A2(n4249), .ZN(n5716) );
  CLKBUF_X1 U3629 ( .A(n4555), .Z(n4601) );
  NAND2_X1 U3630 ( .A1(n3447), .A2(n3446), .ZN(n4599) );
  NAND2_X1 U3631 ( .A1(n4223), .A2(n4222), .ZN(n4489) );
  NAND2_X1 U3632 ( .A1(n3261), .A2(n3260), .ZN(n4302) );
  BUF_X1 U3633 ( .A(n4209), .Z(n4290) );
  CLKBUF_X1 U3634 ( .A(n3266), .Z(n3638) );
  CLKBUF_X1 U3635 ( .A(n3601), .Z(n3129) );
  OR2_X1 U3636 ( .A1(n3362), .A2(n3361), .ZN(n3372) );
  CLKBUF_X1 U3637 ( .A(n3337), .Z(n4611) );
  INV_X1 U3638 ( .A(n3255), .ZN(n3336) );
  INV_X1 U3639 ( .A(n5203), .ZN(n4296) );
  NAND2_X2 U3640 ( .A1(n3142), .A2(n3230), .ZN(n4642) );
  AND4_X1 U3641 ( .A1(n3237), .A2(n3236), .A3(n3235), .A4(n3234), .ZN(n3254)
         );
  NAND2_X2 U3642 ( .A1(n4160), .A2(n6480), .ZN(n6187) );
  INV_X2 U3643 ( .A(n6344), .ZN(n6329) );
  INV_X2 U3644 ( .A(n6613), .ZN(n6682) );
  AND2_X2 U3645 ( .A1(n3149), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5287)
         );
  AND2_X2 U3646 ( .A1(n3151), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n5285)
         );
  NAND2_X1 U3647 ( .A1(n5377), .A2(n5378), .ZN(n5360) );
  NOR2_X4 U3648 ( .A1(n3517), .A2(n3516), .ZN(n3529) );
  NAND2_X2 U3649 ( .A1(n3491), .A2(n3490), .ZN(n3517) );
  OAI21_X2 U3650 ( .B1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n3341), .A(n3340), 
        .ZN(n3345) );
  NAND2_X1 U3651 ( .A1(n3553), .A2(n3125), .ZN(n3122) );
  AND2_X2 U3652 ( .A1(n3122), .A2(n3123), .ZN(n5558) );
  OR2_X1 U3653 ( .A1(n3124), .A2(n3554), .ZN(n3123) );
  INV_X1 U3654 ( .A(n3555), .ZN(n3124) );
  NAND2_X1 U3655 ( .A1(n5505), .A2(n5622), .ZN(n3126) );
  NAND2_X1 U3656 ( .A1(n3345), .A2(n3380), .ZN(n3128) );
  NAND2_X1 U3657 ( .A1(n5505), .A2(n5622), .ZN(n5490) );
  NAND2_X1 U3658 ( .A1(n3345), .A2(n3380), .ZN(n3382) );
  INV_X1 U3659 ( .A(n3130), .ZN(n4170) );
  AND4_X2 U3660 ( .A1(n3189), .A2(n3188), .A3(n3187), .A4(n3186), .ZN(n3190)
         );
  NOR2_X1 U3661 ( .A1(n5203), .A2(n4585), .ZN(n3601) );
  NOR2_X1 U3662 ( .A1(n4642), .A2(n3220), .ZN(n4382) );
  AND4_X2 U3663 ( .A1(n3199), .A2(n3198), .A3(n3197), .A4(n3196), .ZN(n3146)
         );
  AND2_X2 U3664 ( .A1(n3335), .A2(n3334), .ZN(n3130) );
  INV_X1 U3665 ( .A(n3337), .ZN(n3131) );
  INV_X1 U3666 ( .A(n3337), .ZN(n3221) );
  AND2_X2 U3667 ( .A1(n5285), .A2(n3157), .ZN(n3298) );
  AND2_X2 U3668 ( .A1(n5285), .A2(n3158), .ZN(n3392) );
  AND2_X2 U3669 ( .A1(n5285), .A2(n4538), .ZN(n3246) );
  INV_X1 U3670 ( .A(n6546), .ZN(n3132) );
  NAND2_X1 U3671 ( .A1(n3268), .A2(n3135), .ZN(n3133) );
  AND2_X2 U3672 ( .A1(n3133), .A2(n3134), .ZN(n3329) );
  OR2_X1 U3673 ( .A1(n3269), .A2(n3132), .ZN(n3134) );
  AND2_X1 U3674 ( .A1(n3267), .A2(n3270), .ZN(n3135) );
  OR2_X1 U3675 ( .A1(n5603), .A2(n6073), .ZN(n4353) );
  AND2_X2 U3676 ( .A1(n6030), .A2(n6029), .ZN(n6032) );
  OR2_X4 U3677 ( .A1(n5144), .A2(n5143), .ZN(n5712) );
  NOR2_X2 U3678 ( .A1(n5514), .A2(n3573), .ZN(n5505) );
  NAND2_X2 U3679 ( .A1(n5498), .A2(n5989), .ZN(n4338) );
  NOR2_X2 U3680 ( .A1(n5132), .A2(n5249), .ZN(n5246) );
  AOI211_X2 U3681 ( .C1(INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n5610), .A(n5609), .B(n5608), .ZN(n5611) );
  OAI21_X2 U3682 ( .B1(n5520), .B2(n3571), .A(n3570), .ZN(n5498) );
  NAND2_X2 U3683 ( .A1(n5689), .A2(n6854), .ZN(n5520) );
  NOR2_X2 U3684 ( .A1(n5426), .A2(n5429), .ZN(n5416) );
  OAI21_X2 U3685 ( .B1(n5120), .B2(n5116), .A(n5117), .ZN(n5220) );
  AND2_X2 U3686 ( .A1(n5300), .A2(n5285), .ZN(n3438) );
  AND2_X1 U3687 ( .A1(n3332), .A2(n3331), .ZN(n4183) );
  INV_X1 U3688 ( .A(n5735), .ZN(n4997) );
  CLKBUF_X1 U3689 ( .A(n3304), .Z(n3354) );
  CLKBUF_X1 U3690 ( .A(n3246), .Z(n3307) );
  CLKBUF_X1 U3691 ( .A(n3391), .Z(n3306) );
  NAND2_X1 U3692 ( .A1(n3432), .A2(n3431), .ZN(n3632) );
  INV_X1 U3693 ( .A(n5193), .ZN(n4127) );
  NAND2_X1 U3694 ( .A1(n4642), .A2(n4585), .ZN(n4200) );
  NAND2_X1 U3695 ( .A1(n3414), .A2(n3413), .ZN(n3448) );
  OAI21_X1 U3696 ( .B1(n3412), .B2(n3411), .A(n3410), .ZN(n3414) );
  NAND3_X1 U3697 ( .A1(n3449), .A2(n4599), .A3(n3448), .ZN(n3477) );
  AOI22_X1 U3698 ( .A1(n3297), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3246), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3180) );
  OR2_X1 U3699 ( .A1(n4103), .A2(n4102), .ZN(n4104) );
  NOR2_X1 U3700 ( .A1(n3909), .A2(n5563), .ZN(n3910) );
  NAND2_X1 U3701 ( .A1(n3810), .A2(n3809), .ZN(n5103) );
  OR2_X1 U3702 ( .A1(n3807), .A2(n3808), .ZN(n3809) );
  NAND2_X1 U3703 ( .A1(n5103), .A2(n5102), .ZN(n5101) );
  NAND2_X1 U3704 ( .A1(n3792), .A2(n3791), .ZN(n3807) );
  AND2_X1 U3705 ( .A1(n3790), .A2(n3789), .ZN(n3791) );
  INV_X1 U3706 ( .A(n4485), .ZN(n3792) );
  NOR2_X1 U3707 ( .A1(n4849), .A2(n4486), .ZN(n3789) );
  AND2_X1 U3708 ( .A1(n3781), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3774)
         );
  NAND2_X1 U3709 ( .A1(n5489), .A2(n3575), .ZN(n3577) );
  NAND2_X1 U3710 ( .A1(n3119), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3573) );
  INV_X1 U3711 ( .A(n5544), .ZN(n5524) );
  AND2_X1 U3712 ( .A1(n5559), .A2(n3559), .ZN(n3560) );
  OR2_X1 U3713 ( .A1(n5598), .A2(n3557), .ZN(n3561) );
  INV_X1 U3714 ( .A(n4402), .ZN(n4214) );
  NAND2_X2 U3715 ( .A1(n3140), .A2(n3143), .ZN(n4574) );
  AND2_X1 U3716 ( .A1(n4601), .A2(n4600), .ZN(n5833) );
  CLKBUF_X1 U3717 ( .A(n3325), .Z(n6571) );
  CLKBUF_X1 U3718 ( .A(n4183), .Z(n6572) );
  AND2_X1 U3719 ( .A1(n6271), .A2(n5214), .ZN(n6258) );
  NAND2_X1 U3720 ( .A1(n6271), .A2(n5197), .ZN(n6193) );
  NAND2_X1 U3721 ( .A1(n3323), .A2(n3322), .ZN(n3324) );
  INV_X1 U3722 ( .A(n3321), .ZN(n3322) );
  NAND2_X1 U3723 ( .A1(n3131), .A2(n3255), .ZN(n3266) );
  AND2_X1 U3724 ( .A1(n3746), .A2(n5033), .ZN(n3764) );
  OR2_X1 U3725 ( .A1(n3468), .A2(n3467), .ZN(n3495) );
  OR2_X1 U3726 ( .A1(n3403), .A2(n3402), .ZN(n3405) );
  OR2_X1 U3727 ( .A1(n3445), .A2(n3444), .ZN(n3453) );
  OAI22_X1 U3728 ( .A1(n3627), .A2(n3626), .B1(n3625), .B2(n4174), .ZN(n3628)
         );
  NOR2_X2 U3729 ( .A1(n5360), .A2(n5362), .ZN(n4154) );
  NAND2_X1 U3730 ( .A1(n5431), .A2(n5432), .ZN(n5426) );
  NAND2_X1 U3731 ( .A1(n3847), .A2(n3145), .ZN(n5132) );
  NAND2_X1 U3732 ( .A1(n3679), .A2(n3678), .ZN(n4485) );
  INV_X1 U3733 ( .A(n4492), .ZN(n3678) );
  INV_X1 U3734 ( .A(n4390), .ZN(n3679) );
  INV_X1 U3735 ( .A(n4905), .ZN(n3843) );
  NAND2_X1 U3736 ( .A1(n4391), .A2(n4392), .ZN(n4390) );
  INV_X1 U3737 ( .A(n3405), .ZN(n3417) );
  INV_X1 U3738 ( .A(n4097), .ZN(n4344) );
  INV_X1 U3739 ( .A(n3622), .ZN(n3596) );
  INV_X1 U3740 ( .A(n5569), .ZN(n3562) );
  AND2_X1 U3741 ( .A1(n5586), .A2(n3558), .ZN(n5559) );
  AND2_X1 U3742 ( .A1(n5579), .A2(n5576), .ZN(n5560) );
  AND2_X1 U3743 ( .A1(n4237), .A2(n4236), .ZN(n4991) );
  AND2_X1 U3744 ( .A1(n4290), .A2(n5323), .ZN(n4301) );
  INV_X1 U3745 ( .A(n3542), .ZN(n3539) );
  NAND2_X1 U3746 ( .A1(n4381), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3432) );
  OR2_X1 U3748 ( .A1(n3313), .A2(n3312), .ZN(n3373) );
  NAND2_X1 U3749 ( .A1(n3130), .A2(n3271), .ZN(n4190) );
  NAND2_X1 U3750 ( .A1(n3430), .A2(n3429), .ZN(n4564) );
  AOI21_X1 U3751 ( .B1(n6578), .B2(n4637), .A(n5308), .ZN(n4573) );
  INV_X1 U3752 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6557) );
  OR2_X1 U3753 ( .A1(n5291), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4156) );
  NAND2_X1 U3754 ( .A1(n6671), .A2(n5202), .ZN(n6239) );
  AND2_X1 U3755 ( .A1(n4636), .A2(n4635), .ZN(n6300) );
  OR2_X1 U3757 ( .A1(n3992), .A2(n3991), .ZN(n5417) );
  AND2_X1 U3758 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n3945), .ZN(n3946)
         );
  NAND2_X1 U3759 ( .A1(n3946), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3988)
         );
  CLKBUF_X1 U3760 ( .A(n5426), .Z(n5434) );
  OR2_X1 U3761 ( .A1(n3912), .A2(n3911), .ZN(n5449) );
  INV_X1 U3762 ( .A(n5255), .ZN(n5450) );
  CLKBUF_X1 U3763 ( .A(n5254), .Z(n5255) );
  AND2_X1 U3764 ( .A1(n3875), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3876)
         );
  NAND2_X1 U3765 ( .A1(n3876), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3909)
         );
  CLKBUF_X1 U3766 ( .A(n5246), .Z(n5247) );
  NAND2_X1 U3767 ( .A1(n3828), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3829)
         );
  NOR2_X1 U3768 ( .A1(n6977), .A2(n3829), .ZN(n3875) );
  CLKBUF_X1 U3769 ( .A(n5132), .Z(n5248) );
  AND2_X1 U3770 ( .A1(n3822), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3828)
         );
  XNOR2_X1 U3771 ( .A(n3807), .B(n3808), .ZN(n5599) );
  NOR2_X1 U3772 ( .A1(n6914), .A2(n3696), .ZN(n3822) );
  NAND2_X1 U3773 ( .A1(PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n3712), .ZN(n3696)
         );
  NAND2_X1 U3774 ( .A1(n3747), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3713)
         );
  NOR2_X1 U3775 ( .A1(n6838), .A2(n3767), .ZN(n3747) );
  AND2_X1 U3776 ( .A1(n4985), .A2(n4984), .ZN(n5034) );
  NAND2_X1 U3777 ( .A1(n3774), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3767)
         );
  AND2_X1 U3778 ( .A1(n4910), .A2(n4909), .ZN(n4985) );
  AOI21_X1 U3779 ( .B1(n3779), .B2(n4905), .A(n3778), .ZN(n4849) );
  INV_X1 U3780 ( .A(n3664), .ZN(n3665) );
  AND2_X1 U3781 ( .A1(n4507), .A2(n6583), .ZN(n4632) );
  NOR4_X2 U3782 ( .A1(n5499), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A4(n3552), .ZN(n5506) );
  AND2_X1 U3783 ( .A1(n5437), .A2(n5424), .ZN(n5418) );
  OR2_X1 U3784 ( .A1(n5443), .A2(n4268), .ZN(n5436) );
  NOR2_X2 U3785 ( .A1(n5436), .A2(n5435), .ZN(n5437) );
  AOI21_X1 U3786 ( .B1(n5552), .B2(n5551), .A(n5523), .ZN(n5545) );
  CLKBUF_X1 U3787 ( .A(n5557), .Z(n6002) );
  INV_X1 U3788 ( .A(n4200), .ZN(n3256) );
  AND3_X1 U3789 ( .A1(n4239), .A2(n4279), .A3(n4238), .ZN(n5113) );
  NAND2_X1 U3790 ( .A1(n3551), .A2(n3550), .ZN(n5120) );
  AND2_X1 U3791 ( .A1(n4928), .A2(n4927), .ZN(n4992) );
  INV_X1 U3792 ( .A(n4490), .ZN(n4222) );
  INV_X1 U3793 ( .A(n4488), .ZN(n4223) );
  INV_X1 U3794 ( .A(n4156), .ZN(n4160) );
  NAND2_X1 U3795 ( .A1(n3316), .A2(n3323), .ZN(n3320) );
  INV_X1 U3796 ( .A(n4556), .ZN(n4597) );
  OR2_X1 U3797 ( .A1(n4717), .A2(n4601), .ZN(n6473) );
  NAND2_X1 U3798 ( .A1(n3477), .A2(n3451), .ZN(n3663) );
  AND2_X2 U3799 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5309) );
  CLKBUF_X1 U3800 ( .A(n4526), .Z(n4527) );
  AND2_X2 U3801 ( .A1(n3158), .A2(n5309), .ZN(n3347) );
  INV_X1 U3802 ( .A(n4507), .ZN(n4550) );
  CLKBUF_X1 U3803 ( .A(n4190), .Z(n4514) );
  INV_X1 U3804 ( .A(n6473), .ZN(n5734) );
  AND2_X1 U3805 ( .A1(n5722), .A2(n4997), .ZN(n5733) );
  NOR2_X1 U3806 ( .A1(n6661), .A2(n4573), .ZN(n4654) );
  INV_X1 U3807 ( .A(n4720), .ZN(n4784) );
  INV_X1 U3808 ( .A(n4873), .ZN(n6476) );
  NAND2_X1 U3809 ( .A1(n4375), .A2(n4370), .ZN(n6671) );
  AND2_X1 U3810 ( .A1(n6271), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6245) );
  INV_X1 U3811 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6219) );
  INV_X1 U3812 ( .A(n6220), .ZN(n6261) );
  INV_X1 U3813 ( .A(n6245), .ZN(n6256) );
  CLKBUF_X1 U3814 ( .A(n3649), .Z(n6474) );
  XNOR2_X1 U3815 ( .A(n4295), .B(n5329), .ZN(n5375) );
  INV_X1 U3816 ( .A(n6274), .ZN(n6279) );
  NAND2_X1 U3817 ( .A1(n6284), .A2(n5320), .ZN(n6274) );
  AND2_X1 U3818 ( .A1(n6299), .A2(n4483), .ZN(n6292) );
  AND2_X1 U3819 ( .A1(n6299), .A2(n4482), .ZN(n6289) );
  INV_X1 U3820 ( .A(n6299), .ZN(n6291) );
  OR2_X1 U3821 ( .A1(n6289), .A2(n6292), .ZN(n6295) );
  INV_X1 U3822 ( .A(n6295), .ZN(n5107) );
  BUF_X1 U3824 ( .A(n6316), .Z(n6323) );
  CLKBUF_X2 U3825 ( .A(n4634), .Z(n4457) );
  NOR2_X1 U3826 ( .A1(n4348), .A2(n5352), .ZN(n4349) );
  CLKBUF_X1 U3827 ( .A(n5101), .Z(n5131) );
  INV_X1 U3828 ( .A(n6341), .ZN(n5591) );
  INV_X1 U3829 ( .A(n6335), .ZN(n5593) );
  NAND2_X1 U3830 ( .A1(n3585), .A2(n3138), .ZN(n4196) );
  NOR2_X1 U3831 ( .A1(n5692), .A2(n4313), .ZN(n6014) );
  NAND2_X1 U3832 ( .A1(n6047), .A2(n5234), .ZN(n6348) );
  NAND2_X1 U3833 ( .A1(n4318), .A2(n4364), .ZN(n5235) );
  INV_X1 U3834 ( .A(n5235), .ZN(n6377) );
  INV_X1 U3835 ( .A(n6394), .ZN(n6375) );
  OR2_X1 U3836 ( .A1(n6377), .A2(n6051), .ZN(n6392) );
  CLKBUF_X1 U3837 ( .A(n4562), .Z(n4563) );
  INV_X1 U3838 ( .A(n4597), .ZN(n5722) );
  INV_X1 U3839 ( .A(n4601), .ZN(n5725) );
  CLKBUF_X1 U3840 ( .A(n4511), .Z(n6246) );
  INV_X1 U3841 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6563) );
  INV_X1 U3842 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n5295) );
  INV_X1 U3843 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5317) );
  INV_X1 U3844 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3152) );
  INV_X1 U3845 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5304) );
  NOR2_X1 U3846 ( .A1(n6663), .A2(n4550), .ZN(n5308) );
  INV_X1 U3847 ( .A(n4722), .ZN(n4976) );
  OR2_X1 U3848 ( .A1(n4871), .A2(n4997), .ZN(n4898) );
  AND2_X1 U3849 ( .A1(n4828), .A2(n5735), .ZN(n4845) );
  AND2_X1 U3850 ( .A1(n4828), .A2(n4997), .ZN(n5152) );
  INV_X1 U3851 ( .A(n5840), .ZN(n6470) );
  INV_X1 U3852 ( .A(n6484), .ZN(n5747) );
  INV_X1 U3853 ( .A(n5846), .ZN(n6489) );
  INV_X1 U3854 ( .A(n6490), .ZN(n5751) );
  INV_X1 U3855 ( .A(n6496), .ZN(n5755) );
  INV_X1 U3856 ( .A(n5856), .ZN(n6501) );
  INV_X1 U3857 ( .A(n6502), .ZN(n5759) );
  INV_X1 U3858 ( .A(n5862), .ZN(n6507) );
  INV_X1 U3859 ( .A(n5869), .ZN(n6513) );
  INV_X1 U3860 ( .A(n6514), .ZN(n5768) );
  INV_X1 U3861 ( .A(n6531), .ZN(n5182) );
  NOR2_X1 U3862 ( .A1(n4590), .A2(n4784), .ZN(n6484) );
  NOR2_X1 U3863 ( .A1(n4920), .A2(n4784), .ZN(n6496) );
  NOR2_X1 U3864 ( .A1(n6750), .A2(n4784), .ZN(n6502) );
  NOR2_X1 U3865 ( .A1(n4917), .A2(n4784), .ZN(n6508) );
  NOR2_X1 U3866 ( .A1(n4998), .A2(n4997), .ZN(n5866) );
  INV_X1 U3867 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6585) );
  AND2_X1 U3868 ( .A1(n6574), .A2(n6573), .ZN(n6590) );
  INV_X1 U3869 ( .A(n6590), .ZN(n6662) );
  AND2_X2 U3870 ( .A1(n5287), .A2(n3158), .ZN(n3297) );
  XOR2_X1 U3871 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .B(n5500), .Z(n3136) );
  AND4_X1 U3872 ( .A1(n3195), .A2(n3194), .A3(n3193), .A4(n3192), .ZN(n3137)
         );
  AND2_X1 U3873 ( .A1(n4462), .A2(n4461), .ZN(n3659) );
  INV_X1 U3874 ( .A(n3272), .ZN(n3257) );
  NAND2_X2 U3875 ( .A1(n3541), .A2(n3540), .ZN(n3552) );
  AND2_X1 U3876 ( .A1(n3584), .A2(n3583), .ZN(n3138) );
  AND2_X2 U3877 ( .A1(n5300), .A2(n5287), .ZN(n3433) );
  BUF_X1 U3878 ( .A(n3642), .Z(n4556) );
  NAND2_X1 U3879 ( .A1(n4632), .A2(n6537), .ZN(n6073) );
  INV_X1 U3880 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3575) );
  NOR2_X1 U3881 ( .A1(n6405), .A2(n4596), .ZN(n3139) );
  AND4_X1 U3882 ( .A1(n3168), .A2(n3167), .A3(n3166), .A4(n3165), .ZN(n3140)
         );
  AND4_X1 U3883 ( .A1(n3225), .A2(n3224), .A3(n3223), .A4(n3222), .ZN(n3142)
         );
  NAND2_X1 U3884 ( .A1(n3119), .A2(n3564), .ZN(n3144) );
  INV_X1 U3885 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3576) );
  NAND2_X1 U3886 ( .A1(n3846), .A2(n3845), .ZN(n3145) );
  INV_X1 U3887 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6838) );
  AND2_X1 U3888 ( .A1(n4905), .A2(n3805), .ZN(n3147) );
  NOR2_X1 U3889 ( .A1(n6032), .A2(n6031), .ZN(n3148) );
  NAND2_X1 U3890 ( .A1(n4318), .A2(n4194), .ZN(n6399) );
  OAI21_X1 U3891 ( .B1(n3606), .B2(n3271), .A(n4653), .ZN(n3612) );
  INV_X1 U3892 ( .A(n3372), .ZN(n3366) );
  AND2_X1 U3893 ( .A1(n3258), .A2(n4515), .ZN(n3278) );
  AND2_X1 U3894 ( .A1(n3764), .A2(n4984), .ZN(n3766) );
  NOR2_X1 U3895 ( .A1(n3601), .A2(n3602), .ZN(n3624) );
  NAND2_X1 U3897 ( .A1(n3638), .A2(n3625), .ZN(n3267) );
  AND2_X1 U3898 ( .A1(n4905), .A2(n3766), .ZN(n3765) );
  NAND2_X1 U3899 ( .A1(n3369), .A2(n3368), .ZN(n3410) );
  INV_X1 U3900 ( .A(n3632), .ZN(n3606) );
  INV_X1 U3901 ( .A(n3493), .ZN(n3490) );
  INV_X1 U3902 ( .A(n3407), .ZN(n3408) );
  INV_X2 U3903 ( .A(n3597), .ZN(n3625) );
  OR2_X1 U3904 ( .A1(n3770), .A2(n4907), .ZN(n3771) );
  BUF_X1 U3905 ( .A(n3348), .Z(n4107) );
  INV_X1 U3906 ( .A(n3527), .ZN(n3528) );
  NAND2_X1 U3907 ( .A1(n4296), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3431) );
  OR2_X1 U3908 ( .A1(n3296), .A2(n3295), .ZN(n3542) );
  NAND3_X1 U3909 ( .A1(n4579), .A2(STATE2_REG_0__SCAN_IN), .A3(n5203), .ZN(
        n3597) );
  NAND2_X1 U3910 ( .A1(n4186), .A2(n4642), .ZN(n4304) );
  NOR2_X1 U3911 ( .A1(n6561), .A2(n3594), .ZN(n4177) );
  INV_X1 U3912 ( .A(n5449), .ZN(n3913) );
  INV_X1 U3913 ( .A(n5417), .ZN(n3993) );
  INV_X1 U3914 ( .A(n3944), .ZN(n3945) );
  NAND2_X1 U3915 ( .A1(n3259), .A2(n3286), .ZN(n3260) );
  NAND2_X1 U3916 ( .A1(n3221), .A2(n4574), .ZN(n3647) );
  NOR2_X1 U3917 ( .A1(n4396), .A2(n4394), .ZN(n4497) );
  NAND2_X1 U3918 ( .A1(n3390), .A2(n3389), .ZN(n3425) );
  XNOR2_X1 U3919 ( .A(n4544), .B(n4564), .ZN(n4526) );
  XNOR2_X1 U3920 ( .A(n3415), .B(n3448), .ZN(n4555) );
  AND2_X1 U3921 ( .A1(n4073), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4074)
         );
  NOR2_X1 U3922 ( .A1(n3672), .A2(n6219), .ZN(n3680) );
  INV_X1 U3923 ( .A(n5385), .ZN(n4078) );
  OR2_X1 U3924 ( .A1(n4104), .A2(n5363), .ZN(n4348) );
  AND2_X1 U3925 ( .A1(n3729), .A2(n3728), .ZN(n5109) );
  NAND2_X1 U3926 ( .A1(n3257), .A2(n3256), .ZN(n4515) );
  OAI211_X1 U3927 ( .C1(n3499), .C2(n3498), .A(n3530), .B(n6571), .ZN(n3500)
         );
  INV_X1 U3928 ( .A(n4403), .ZN(n4213) );
  NAND2_X1 U3929 ( .A1(n5094), .A2(n3379), .ZN(n6327) );
  OR2_X1 U3930 ( .A1(n4616), .A2(n5722), .ZN(n4871) );
  INV_X1 U3931 ( .A(n4599), .ZN(n4557) );
  INV_X1 U3932 ( .A(n5812), .ZN(n5822) );
  INV_X1 U3933 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6948) );
  AND2_X1 U3934 ( .A1(n3271), .A2(n5203), .ZN(n3325) );
  NAND2_X1 U3935 ( .A1(n4183), .A2(n5203), .ZN(n4357) );
  NAND2_X1 U3936 ( .A1(n4074), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4103)
         );
  NOR2_X1 U3937 ( .A1(n3988), .A2(n5541), .ZN(n3989) );
  NOR2_X1 U3938 ( .A1(n6825), .A2(n3713), .ZN(n3712) );
  AND2_X1 U3939 ( .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n3680), .ZN(n3781)
         );
  NAND2_X1 U3941 ( .A1(n6032), .A2(n5452), .ZN(n5443) );
  NAND2_X1 U3942 ( .A1(n4992), .A2(n4991), .ZN(n4990) );
  NAND2_X1 U3943 ( .A1(n3646), .A2(n3645), .ZN(n4462) );
  BUF_X1 U3944 ( .A(n4154), .Z(n5361) );
  OR2_X1 U3945 ( .A1(n4031), .A2(n4030), .ZN(n4033) );
  OR2_X1 U3946 ( .A1(n4574), .A2(n4606), .ZN(n4097) );
  OR2_X1 U3947 ( .A1(n5110), .A2(n5109), .ZN(n5139) );
  OR2_X1 U3948 ( .A1(n3635), .A2(n3634), .ZN(n4507) );
  OAI21_X1 U3949 ( .B1(n5490), .B2(n5605), .A(n4341), .ZN(n4342) );
  NAND2_X1 U3950 ( .A1(n5418), .A2(n5419), .ZN(n5421) );
  AND2_X1 U3951 ( .A1(n3119), .A2(n5703), .ZN(n5569) );
  OR2_X1 U3952 ( .A1(n5558), .A2(n5598), .ZN(n5596) );
  CLKBUF_X1 U3953 ( .A(n4488), .Z(n4499) );
  NAND2_X1 U3954 ( .A1(n4214), .A2(n4213), .ZN(n4396) );
  NAND2_X1 U3955 ( .A1(n4465), .A2(n4208), .ZN(n4402) );
  INV_X1 U3956 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3149) );
  OR2_X1 U3957 ( .A1(n4598), .A2(n4601), .ZN(n4754) );
  OR2_X1 U3958 ( .A1(n4871), .A2(n5735), .ZN(n6413) );
  INV_X1 U3959 ( .A(n4845), .ZN(n4813) );
  AND4_X1 U3960 ( .A1(n3203), .A2(n3202), .A3(n3201), .A4(n3200), .ZN(n3219)
         );
  INV_X1 U3961 ( .A(n5152), .ZN(n5188) );
  NOR2_X1 U3962 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4573), .ZN(n4720) );
  AOI21_X1 U3963 ( .B1(n6411), .B2(STATE2_REG_3__SCAN_IN), .A(n4784), .ZN(
        n4873) );
  INV_X1 U3964 ( .A(n4357), .ZN(n4361) );
  AND2_X1 U3965 ( .A1(n5340), .A2(n5919), .ZN(n5906) );
  NAND2_X1 U3966 ( .A1(n3989), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4031)
         );
  AND2_X1 U3967 ( .A1(n5213), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5197) );
  INV_X1 U3968 ( .A(n6671), .ZN(n5212) );
  INV_X1 U3969 ( .A(n6239), .ZN(n6244) );
  NAND2_X1 U3970 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3665), .ZN(n3672)
         );
  INV_X1 U3971 ( .A(n4301), .ZN(n5331) );
  NOR2_X1 U3972 ( .A1(n6674), .A2(n6300), .ZN(n6316) );
  INV_X1 U3973 ( .A(n4476), .ZN(n4448) );
  NOR2_X1 U3974 ( .A1(n4033), .A2(n4032), .ZN(n4073) );
  NAND2_X1 U3975 ( .A1(n3910), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3944)
         );
  AND2_X1 U3976 ( .A1(n5139), .A2(n5111), .ZN(n6155) );
  NAND2_X1 U3977 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3664) );
  INV_X1 U3978 ( .A(n6399), .ZN(n4195) );
  INV_X1 U3979 ( .A(n6021), .ZN(n5642) );
  OAI22_X1 U3980 ( .A1(n5532), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n5539), .B2(n5525), .ZN(n5526) );
  AND2_X1 U3981 ( .A1(n5520), .A2(n5522), .ZN(n5552) );
  AND2_X1 U3982 ( .A1(n4318), .A2(n4309), .ZN(n6051) );
  NAND2_X1 U3983 ( .A1(n4188), .A2(n4187), .ZN(n4318) );
  AND2_X1 U3984 ( .A1(n5833), .A2(n4997), .ZN(n5878) );
  NOR2_X1 U3985 ( .A1(n4754), .A2(n4997), .ZN(n4777) );
  INV_X1 U3986 ( .A(n6413), .ZN(n6443) );
  OR2_X1 U3987 ( .A1(n4786), .A2(n4785), .ZN(n4816) );
  INV_X1 U3988 ( .A(n6535), .ZN(n6518) );
  INV_X1 U3989 ( .A(n5851), .ZN(n6495) );
  NOR2_X1 U3990 ( .A1(n4919), .A2(n4784), .ZN(n6490) );
  NOR2_X1 U3991 ( .A1(n4652), .A2(n4784), .ZN(n6514) );
  NAND2_X1 U3992 ( .A1(n4361), .A2(n4632), .ZN(n4375) );
  INV_X1 U3993 ( .A(n6262), .ZN(n6176) );
  OR2_X1 U3994 ( .A1(n5212), .A2(n5205), .ZN(n6220) );
  OR2_X1 U3995 ( .A1(n6671), .A2(n5196), .ZN(n6271) );
  NAND2_X1 U3996 ( .A1(n4477), .A2(n4476), .ZN(n6299) );
  INV_X1 U3997 ( .A(n6300), .ZN(n6325) );
  AOI21_X1 U3998 ( .B1(n5593), .B2(n5213), .A(n4350), .ZN(n4351) );
  OR2_X1 U3999 ( .A1(n5141), .A2(n5140), .ZN(n6145) );
  NAND2_X1 U4000 ( .A1(n5591), .A2(n6340), .ZN(n6335) );
  AND2_X1 U4001 ( .A1(n5658), .A2(n4330), .ZN(n6021) );
  INV_X1 U4002 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6411) );
  INV_X1 U4003 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6546) );
  NAND2_X1 U4004 ( .A1(n4572), .A2(n5153), .ZN(n6466) );
  INV_X1 U4005 ( .A(n6521), .ZN(n5178) );
  NAND2_X1 U4006 ( .A1(n5734), .A2(n5733), .ZN(n6524) );
  INV_X1 U4007 ( .A(n6508), .ZN(n5763) );
  INV_X1 U4008 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6663) );
  NOR2_X4 U4009 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4548) );
  AND2_X2 U4010 ( .A1(n3157), .A2(n4548), .ZN(n3355) );
  AND2_X2 U4011 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4538) );
  AND2_X2 U4012 ( .A1(n4548), .A2(n4538), .ZN(n3356) );
  AOI22_X1 U4013 ( .A1(n3355), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3156) );
  INV_X1 U4014 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3150) );
  AND2_X2 U4015 ( .A1(n3150), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3158)
         );
  INV_X1 U4016 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3151) );
  AOI22_X1 U4017 ( .A1(n3297), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3246), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3155) );
  AND2_X4 U4018 ( .A1(n3152), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n5300)
         );
  AND2_X2 U4019 ( .A1(n3157), .A2(n5309), .ZN(n3349) );
  AOI22_X1 U4020 ( .A1(n3438), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3154) );
  AOI22_X1 U4021 ( .A1(n3298), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3347), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3153) );
  AND2_X2 U4022 ( .A1(n5287), .A2(n3157), .ZN(n3299) );
  AND2_X2 U4023 ( .A1(n5287), .A2(n4538), .ZN(n3304) );
  AOI22_X1 U4024 ( .A1(n3299), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3162) );
  AOI22_X1 U4025 ( .A1(n3433), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4136), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3161) );
  AND2_X2 U4026 ( .A1(n3158), .A2(n4548), .ZN(n3305) );
  AND2_X4 U4027 ( .A1(n5300), .A2(n4548), .ZN(n3391) );
  AOI22_X1 U4028 ( .A1(n3305), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3160) );
  AND2_X2 U4029 ( .A1(n5309), .A2(n4538), .ZN(n4137) );
  AOI22_X1 U4030 ( .A1(n3392), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4137), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3159) );
  AND4_X2 U4031 ( .A1(n3162), .A2(n3161), .A3(n3160), .A4(n3159), .ZN(n3163)
         );
  NAND2_X2 U4032 ( .A1(n3164), .A2(n3163), .ZN(n3337) );
  AOI22_X1 U4033 ( .A1(n3299), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3168) );
  AOI22_X1 U4034 ( .A1(n3433), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4136), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3167) );
  AOI22_X1 U4035 ( .A1(n3305), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U4036 ( .A1(n3392), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4137), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3165) );
  AOI22_X1 U4037 ( .A1(n3355), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3172) );
  AOI22_X1 U4038 ( .A1(n3438), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3171) );
  AOI22_X1 U4039 ( .A1(n3298), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3347), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3170) );
  AOI22_X1 U4040 ( .A1(n3297), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3246), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3169) );
  AOI22_X1 U4041 ( .A1(n3299), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3176) );
  AOI22_X1 U4042 ( .A1(n3433), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4136), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3175) );
  AOI22_X1 U4043 ( .A1(n3392), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4137), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3174) );
  AOI22_X1 U4044 ( .A1(n3305), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4046 ( .A1(n3438), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3179) );
  AOI22_X1 U4047 ( .A1(n3298), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3347), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3178) );
  AOI22_X1 U4048 ( .A1(n3355), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3177) );
  NAND2_X2 U4049 ( .A1(n3181), .A2(n3141), .ZN(n4579) );
  INV_X2 U4050 ( .A(n4579), .ZN(n3286) );
  AOI22_X1 U4051 ( .A1(n3355), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3185) );
  AOI22_X1 U4052 ( .A1(n3392), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3184) );
  AOI22_X1 U4053 ( .A1(n3438), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3297), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3183) );
  AOI22_X1 U4054 ( .A1(n3299), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4136), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3182) );
  AND4_X2 U4055 ( .A1(n3185), .A2(n3184), .A3(n3183), .A4(n3182), .ZN(n3191)
         );
  AOI22_X1 U4056 ( .A1(n3305), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3189) );
  AOI22_X1 U4057 ( .A1(n3433), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4137), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3188) );
  AOI22_X1 U4058 ( .A1(n3298), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3347), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3187) );
  AOI22_X1 U4059 ( .A1(n3246), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3186) );
  NAND2_X2 U4060 ( .A1(n3191), .A2(n3190), .ZN(n3255) );
  NAND2_X2 U4061 ( .A1(n3336), .A2(n3337), .ZN(n4383) );
  NAND3_X1 U4062 ( .A1(n3647), .A2(n3286), .A3(n4383), .ZN(n3333) );
  AOI22_X1 U4063 ( .A1(n3438), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3246), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3195) );
  AOI22_X1 U4064 ( .A1(n3392), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3194) );
  AOI22_X1 U4065 ( .A1(n3299), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3305), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3193) );
  AOI22_X1 U4066 ( .A1(n3356), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4137), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3192) );
  AOI22_X1 U4067 ( .A1(n3298), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4136), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3199) );
  AOI22_X1 U4068 ( .A1(n3433), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3198) );
  AOI22_X1 U4069 ( .A1(n3297), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3197) );
  AOI22_X1 U4070 ( .A1(n3347), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3355), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3196) );
  NAND2_X2 U4071 ( .A1(n3137), .A2(n3146), .ZN(n3220) );
  NAND2_X1 U4072 ( .A1(n3438), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3203) );
  NAND2_X1 U4073 ( .A1(n3297), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3202) );
  NAND2_X1 U4074 ( .A1(n3246), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3201)
         );
  NAND2_X1 U4075 ( .A1(n3349), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3200) );
  NAND2_X1 U4076 ( .A1(n3433), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3207)
         );
  NAND2_X1 U4077 ( .A1(n4136), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3206)
         );
  NAND2_X1 U4078 ( .A1(n3305), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3205) );
  NAND2_X1 U4079 ( .A1(n3391), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3204) );
  AND4_X2 U4080 ( .A1(n3207), .A2(n3206), .A3(n3205), .A4(n3204), .ZN(n3218)
         );
  NAND2_X1 U4081 ( .A1(n3392), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3211) );
  NAND2_X1 U4082 ( .A1(n3299), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3210) );
  NAND2_X1 U4083 ( .A1(n3304), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3209)
         );
  NAND2_X1 U4084 ( .A1(n4137), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3208)
         );
  AND4_X2 U4085 ( .A1(n3211), .A2(n3210), .A3(n3209), .A4(n3208), .ZN(n3217)
         );
  NAND2_X1 U4086 ( .A1(n3298), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3215) );
  NAND2_X1 U4087 ( .A1(n3347), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3214) );
  NAND2_X1 U4088 ( .A1(n3355), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3213) );
  NAND2_X1 U4089 ( .A1(n3356), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3212)
         );
  AND4_X2 U4090 ( .A1(n3215), .A2(n3214), .A3(n3213), .A4(n3212), .ZN(n3216)
         );
  NAND4_X4 U4091 ( .A1(n3219), .A2(n3218), .A3(n3217), .A4(n3216), .ZN(n4585)
         );
  AOI21_X1 U4092 ( .B1(n3333), .B2(n3220), .A(n4585), .ZN(n3233) );
  NAND2_X1 U4093 ( .A1(n3221), .A2(n4579), .ZN(n3275) );
  INV_X2 U4094 ( .A(n3220), .ZN(n4186) );
  NAND3_X1 U4095 ( .A1(n4383), .A2(n3275), .A3(n4186), .ZN(n3232) );
  AOI22_X1 U4096 ( .A1(n3299), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3304), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3225) );
  AOI22_X1 U4097 ( .A1(n3433), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4136), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3224) );
  AOI22_X1 U4098 ( .A1(n3305), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3223) );
  AOI22_X1 U4099 ( .A1(n3392), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4137), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3222) );
  AOI22_X1 U4100 ( .A1(n3297), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3246), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3229) );
  AOI22_X1 U4101 ( .A1(n3298), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3347), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3228) );
  AOI22_X1 U4102 ( .A1(n3438), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3227) );
  AOI22_X1 U4103 ( .A1(n3355), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3356), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3226) );
  NAND2_X1 U4104 ( .A1(n3266), .A2(n4642), .ZN(n3231) );
  AND3_X2 U4105 ( .A1(n3232), .A2(n3231), .A3(n4574), .ZN(n3334) );
  NAND2_X1 U4106 ( .A1(n3233), .A2(n3334), .ZN(n3273) );
  NAND2_X1 U4107 ( .A1(n4136), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3237)
         );
  NAND2_X1 U4108 ( .A1(n3304), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3236)
         );
  NAND2_X1 U4109 ( .A1(n3305), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3235) );
  NAND2_X1 U4110 ( .A1(n3391), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3234) );
  NAND2_X1 U4111 ( .A1(n3392), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3241) );
  NAND2_X1 U4112 ( .A1(n3298), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U4113 ( .A1(n3433), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3239)
         );
  NAND2_X1 U4114 ( .A1(n3299), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3238) );
  NAND2_X1 U4115 ( .A1(n3297), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3245) );
  NAND2_X1 U4116 ( .A1(n3438), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3244) );
  NAND2_X1 U4117 ( .A1(n3347), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3243) );
  NAND2_X1 U4118 ( .A1(n3355), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3242) );
  NAND2_X1 U4119 ( .A1(n3349), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3250) );
  NAND2_X1 U4120 ( .A1(n3246), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3249)
         );
  NAND2_X1 U4121 ( .A1(n3356), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3248)
         );
  NAND2_X1 U4122 ( .A1(n4137), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3247)
         );
  NAND4_X4 U4123 ( .A1(n3254), .A2(n3253), .A3(n3252), .A4(n3251), .ZN(n5203)
         );
  NAND2_X1 U4124 ( .A1(n3273), .A2(n4296), .ZN(n3264) );
  NAND3_X1 U4125 ( .A1(n4383), .A2(n3286), .A3(n4574), .ZN(n4168) );
  NAND2_X1 U4126 ( .A1(n4168), .A2(n3325), .ZN(n3258) );
  BUF_X4 U4127 ( .A(n3255), .Z(n4653) );
  NAND2_X1 U4128 ( .A1(n3286), .A2(n4653), .ZN(n3272) );
  INV_X1 U4129 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6612) );
  XNOR2_X1 U4130 ( .A(n6612), .B(STATE_REG_1__SCAN_IN), .ZN(n4172) );
  NOR2_X1 U4131 ( .A1(n4585), .A2(n4172), .ZN(n3338) );
  INV_X1 U4132 ( .A(n4304), .ZN(n3639) );
  OAI21_X1 U4133 ( .B1(n3338), .B2(n4653), .A(n3639), .ZN(n3262) );
  AND2_X1 U4134 ( .A1(n4383), .A2(n4574), .ZN(n3261) );
  INV_X1 U4135 ( .A(n3266), .ZN(n3259) );
  NOR2_X1 U4136 ( .A1(n3262), .A2(n4302), .ZN(n3263) );
  NAND3_X1 U4137 ( .A1(n3264), .A2(n3278), .A3(n3263), .ZN(n3265) );
  NAND2_X1 U4138 ( .A1(n3265), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3268) );
  NAND2_X1 U4139 ( .A1(n3268), .A2(n3267), .ZN(n3383) );
  AND2_X1 U4140 ( .A1(n5295), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3636) );
  INV_X1 U4141 ( .A(n3636), .ZN(n3388) );
  NAND2_X1 U4142 ( .A1(n6663), .A2(n5295), .ZN(n5291) );
  MUX2_X1 U4143 ( .A(n3388), .B(n4160), .S(n6411), .Z(n3269) );
  INV_X1 U4144 ( .A(n3269), .ZN(n3270) );
  OAI21_X1 U4145 ( .B1(n3271), .B2(n3272), .A(n3273), .ZN(n3274) );
  MUX2_X1 U4146 ( .A(n4186), .B(n3274), .S(n4296), .Z(n4307) );
  NOR2_X1 U4147 ( .A1(n5291), .A2(n6585), .ZN(n6584) );
  INV_X1 U4148 ( .A(n3275), .ZN(n3276) );
  AOI22_X1 U4149 ( .A1(n3259), .A2(n3325), .B1(n3276), .B2(n4382), .ZN(n3277)
         );
  INV_X1 U4150 ( .A(n4642), .ZN(n3279) );
  NAND2_X1 U4151 ( .A1(n3279), .A2(n5203), .ZN(n4209) );
  NAND4_X1 U4152 ( .A1(n3278), .A2(n6584), .A3(n3277), .A4(n4209), .ZN(n3283)
         );
  INV_X1 U4153 ( .A(n4302), .ZN(n3281) );
  AOI21_X1 U4154 ( .B1(n3638), .B2(n4579), .A(n3279), .ZN(n3280) );
  AOI21_X1 U4155 ( .B1(n3281), .B2(n3280), .A(n3271), .ZN(n3282) );
  NOR2_X1 U4156 ( .A1(n3283), .A2(n3282), .ZN(n3284) );
  NAND2_X1 U4157 ( .A1(n4307), .A2(n3284), .ZN(n3328) );
  INV_X1 U4158 ( .A(n3328), .ZN(n3285) );
  XNOR2_X1 U4159 ( .A(n3329), .B(n3285), .ZN(n3649) );
  NAND2_X1 U4160 ( .A1(n3649), .A2(n6585), .ZN(n3316) );
  INV_X1 U4161 ( .A(n3432), .ZN(n3315) );
  AOI22_X1 U4162 ( .A1(n3120), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3290) );
  BUF_X1 U4163 ( .A(n3305), .Z(n3348) );
  AOI22_X1 U4164 ( .A1(n3348), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3289) );
  AOI22_X1 U4165 ( .A1(n4106), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3288) );
  AOI22_X1 U4167 ( .A1(n5301), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3287) );
  NAND4_X1 U4168 ( .A1(n3290), .A2(n3289), .A3(n3288), .A4(n3287), .ZN(n3296)
         );
  AOI22_X1 U4169 ( .A1(n3307), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3294) );
  AOI22_X1 U4170 ( .A1(n4087), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3293) );
  AOI22_X1 U4171 ( .A1(n4135), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3292) );
  AOI22_X1 U4172 ( .A1(n4138), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3291) );
  NAND4_X1 U4173 ( .A1(n3294), .A2(n3293), .A3(n3292), .A4(n3291), .ZN(n3295)
         );
  AOI22_X1 U4174 ( .A1(n4135), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4175 ( .A1(n4081), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n5301), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3302) );
  BUF_X1 U4176 ( .A(n3299), .Z(n4128) );
  AOI22_X1 U4177 ( .A1(n3120), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3301) );
  AOI22_X1 U4178 ( .A1(n4138), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3300) );
  NAND4_X1 U4179 ( .A1(n3303), .A2(n3302), .A3(n3301), .A4(n3300), .ZN(n3313)
         );
  AOI22_X1 U4180 ( .A1(n3354), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4181 ( .A1(n3348), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3310) );
  AOI22_X1 U4182 ( .A1(n3307), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3309) );
  AOI22_X1 U4183 ( .A1(n3397), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3308) );
  NAND4_X1 U4184 ( .A1(n3311), .A2(n3310), .A3(n3309), .A4(n3308), .ZN(n3312)
         );
  XNOR2_X1 U4185 ( .A(n3539), .B(n3373), .ZN(n3314) );
  NAND2_X1 U4186 ( .A1(n3315), .A2(n3314), .ZN(n3323) );
  INV_X1 U4187 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3319) );
  AOI21_X1 U4188 ( .B1(n4381), .B2(n3542), .A(n6585), .ZN(n3318) );
  NAND2_X1 U4189 ( .A1(n4296), .A2(n3373), .ZN(n3317) );
  OAI211_X1 U4190 ( .C1(n3597), .C2(n3319), .A(n3318), .B(n3317), .ZN(n3321)
         );
  NAND2_X1 U4191 ( .A1(n3320), .A2(n3321), .ZN(n3369) );
  NAND2_X2 U4192 ( .A1(n3369), .A2(n3324), .ZN(n5735) );
  NAND2_X1 U4193 ( .A1(n4653), .A2(n4585), .ZN(n3622) );
  INV_X1 U4194 ( .A(n3373), .ZN(n3326) );
  AND2_X1 U4195 ( .A1(n4296), .A2(n4642), .ZN(n3418) );
  AOI21_X1 U4196 ( .B1(n3326), .B2(n6571), .A(n3418), .ZN(n3327) );
  OAI21_X2 U4197 ( .B1(n5735), .B2(n3622), .A(n3327), .ZN(n4405) );
  NAND2_X1 U4198 ( .A1(n4405), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3378)
         );
  XNOR2_X1 U4199 ( .A(n3378), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5092)
         );
  AND2_X2 U4200 ( .A1(n3329), .A2(n3328), .ZN(n3381) );
  INV_X1 U4201 ( .A(n3381), .ZN(n3346) );
  XNOR2_X1 U4202 ( .A(n6411), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6405)
         );
  AND2_X1 U4203 ( .A1(n3388), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3330)
         );
  AOI21_X1 U4204 ( .B1(n4160), .B2(n6405), .A(n3330), .ZN(n3343) );
  INV_X1 U4205 ( .A(n3343), .ZN(n3341) );
  INV_X1 U4206 ( .A(n4168), .ZN(n3332) );
  NOR2_X1 U4207 ( .A1(n4304), .A2(n4653), .ZN(n3331) );
  NOR2_X1 U4208 ( .A1(n3333), .A2(n5203), .ZN(n3335) );
  NAND3_X1 U4209 ( .A1(n3601), .A2(n4382), .A3(n4478), .ZN(n4512) );
  NAND2_X1 U4210 ( .A1(n4611), .A2(n4574), .ZN(n4479) );
  OR2_X2 U4211 ( .A1(n4512), .A2(n4479), .ZN(n4198) );
  OAI211_X1 U4212 ( .C1(n3338), .C2(n4357), .A(n4190), .B(n4198), .ZN(n3339)
         );
  NAND2_X1 U4213 ( .A1(n3339), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3342) );
  INV_X1 U4214 ( .A(n3342), .ZN(n3340) );
  NAND2_X1 U4215 ( .A1(n3383), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3344) );
  NAND3_X2 U4216 ( .A1(n3344), .A2(n3343), .A3(n3342), .ZN(n3380) );
  XNOR2_X2 U4217 ( .A(n3346), .B(n3128), .ZN(n4562) );
  AOI22_X1 U4218 ( .A1(n4081), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n5301), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4219 ( .A1(n3120), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4220 ( .A1(n4107), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U4221 ( .A1(n4135), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3350) );
  NAND4_X1 U4222 ( .A1(n3353), .A2(n3352), .A3(n3351), .A4(n3350), .ZN(n3362)
         );
  AOI22_X1 U4223 ( .A1(n4106), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4134), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3360) );
  AOI22_X1 U4224 ( .A1(n4055), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3359) );
  AOI22_X1 U4225 ( .A1(n3397), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4226 ( .A1(n4138), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3357) );
  NAND4_X1 U4227 ( .A1(n3360), .A2(n3359), .A3(n3358), .A4(n3357), .ZN(n3361)
         );
  OR2_X1 U4228 ( .A1(n3432), .A2(n3366), .ZN(n3363) );
  OAI21_X4 U4229 ( .B1(n4562), .B2(STATE2_REG_0__SCAN_IN), .A(n3363), .ZN(
        n3412) );
  OR2_X1 U4230 ( .A1(n3432), .A2(n3542), .ZN(n3365) );
  NAND2_X1 U4231 ( .A1(n3625), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3364) );
  OAI211_X1 U4232 ( .C1(n3431), .C2(n3366), .A(n3365), .B(n3364), .ZN(n3411)
         );
  INV_X1 U4233 ( .A(n3411), .ZN(n3367) );
  XNOR2_X1 U4234 ( .A(n3412), .B(n3367), .ZN(n3371) );
  OR2_X1 U4235 ( .A1(n3432), .A2(n3539), .ZN(n3368) );
  INV_X1 U4236 ( .A(n3410), .ZN(n3370) );
  XNOR2_X1 U4237 ( .A(n3371), .B(n3370), .ZN(n3642) );
  NAND2_X1 U4238 ( .A1(n3642), .A2(n3596), .ZN(n3377) );
  NAND2_X1 U4239 ( .A1(n3373), .A2(n3372), .ZN(n3416) );
  OAI211_X1 U4240 ( .C1(n3373), .C2(n3372), .A(n6571), .B(n3416), .ZN(n3375)
         );
  NOR2_X1 U4241 ( .A1(n4304), .A2(n4478), .ZN(n3374) );
  AND2_X1 U4242 ( .A1(n3375), .A2(n3374), .ZN(n3376) );
  NAND2_X1 U4243 ( .A1(n3377), .A2(n3376), .ZN(n5091) );
  NAND2_X1 U4244 ( .A1(n5092), .A2(n5091), .ZN(n5094) );
  INV_X1 U4245 ( .A(n3378), .ZN(n4406) );
  NAND2_X1 U4246 ( .A1(n4406), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3379)
         );
  OAI21_X2 U4247 ( .B1(n3382), .B2(n3381), .A(n3380), .ZN(n3424) );
  NAND2_X1 U4249 ( .A1(n3384), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3390) );
  AND2_X1 U4250 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3385) );
  NAND2_X1 U4251 ( .A1(n3385), .A2(n6557), .ZN(n6468) );
  INV_X1 U4252 ( .A(n3385), .ZN(n3386) );
  NAND2_X1 U4253 ( .A1(n3386), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3387) );
  NAND2_X1 U4254 ( .A1(n6468), .A2(n3387), .ZN(n4607) );
  AOI22_X1 U4255 ( .A1(n4160), .A2(n4607), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3388), .ZN(n3389) );
  XNOR2_X1 U4256 ( .A(n3424), .B(n3425), .ZN(n4511) );
  AOI22_X1 U4257 ( .A1(n4087), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3396) );
  AOI22_X1 U4258 ( .A1(n3120), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3395) );
  INV_X1 U4259 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6930) );
  AOI22_X1 U4260 ( .A1(n4107), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3394) );
  AOI22_X1 U4261 ( .A1(n4138), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3393) );
  NAND4_X1 U4262 ( .A1(n3396), .A2(n3395), .A3(n3394), .A4(n3393), .ZN(n3403)
         );
  AOI22_X1 U4263 ( .A1(n4106), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4134), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4264 ( .A1(n4081), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n5301), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3400) );
  AOI22_X1 U4265 ( .A1(n4135), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3399) );
  BUF_X1 U4266 ( .A(n3397), .Z(n4108) );
  AOI22_X1 U4267 ( .A1(n4108), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3398) );
  NAND4_X1 U4268 ( .A1(n3401), .A2(n3400), .A3(n3399), .A4(n3398), .ZN(n3402)
         );
  NOR2_X1 U4269 ( .A1(n3432), .A2(n3417), .ZN(n3404) );
  AOI21_X2 U4270 ( .B1(n4511), .B2(n6585), .A(n3404), .ZN(n3409) );
  INV_X1 U4271 ( .A(n3431), .ZN(n3406) );
  AOI22_X1 U4272 ( .A1(n3406), .A2(n3405), .B1(n3625), .B2(
        INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3407) );
  XNOR2_X2 U4273 ( .A(n3409), .B(n3408), .ZN(n3449) );
  INV_X1 U4274 ( .A(n3449), .ZN(n3415) );
  NAND2_X1 U4275 ( .A1(n3412), .A2(n3411), .ZN(n3413) );
  NAND2_X1 U4276 ( .A1(n4555), .A2(n3596), .ZN(n3421) );
  NAND2_X1 U4277 ( .A1(n3416), .A2(n3417), .ZN(n3452) );
  OAI21_X1 U4278 ( .B1(n3417), .B2(n3416), .A(n3452), .ZN(n3419) );
  AOI21_X1 U4279 ( .B1(n3419), .B2(n6571), .A(n3418), .ZN(n3420) );
  NAND2_X1 U4280 ( .A1(n3421), .A2(n3420), .ZN(n6326) );
  OAI21_X1 U4281 ( .B1(n6327), .B2(INSTADDRPOINTER_REG_2__SCAN_IN), .A(n6326), 
        .ZN(n3423) );
  NAND2_X1 U4282 ( .A1(n6327), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3422)
         );
  NAND2_X1 U4283 ( .A1(n3423), .A2(n3422), .ZN(n4675) );
  INV_X1 U4284 ( .A(n3424), .ZN(n3426) );
  NAND2_X1 U4285 ( .A1(n3384), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3430) );
  NOR3_X1 U4286 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6557), .A3(n6948), 
        .ZN(n6410) );
  NAND2_X1 U4287 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6410), .ZN(n6449) );
  NAND2_X1 U4288 ( .A1(n6563), .A2(n6449), .ZN(n3427) );
  NOR3_X1 U4289 ( .A1(n6563), .A2(n6557), .A3(n6948), .ZN(n5834) );
  NAND2_X1 U4290 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5834), .ZN(n5868) );
  NAND2_X1 U4291 ( .A1(n3427), .A2(n5868), .ZN(n4783) );
  OAI22_X1 U4292 ( .A1(n4156), .A2(n4783), .B1(n3636), .B2(n6563), .ZN(n3428)
         );
  INV_X1 U4293 ( .A(n3428), .ZN(n3429) );
  NAND2_X1 U4294 ( .A1(n4526), .A2(n6585), .ZN(n3447) );
  AOI22_X1 U4295 ( .A1(n4087), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3437) );
  AOI22_X1 U4296 ( .A1(n3120), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3436) );
  AOI22_X1 U4297 ( .A1(n4107), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3435) );
  AOI22_X1 U4298 ( .A1(n4138), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3434) );
  NAND4_X1 U4299 ( .A1(n3437), .A2(n3436), .A3(n3435), .A4(n3434), .ZN(n3445)
         );
  INV_X1 U4300 ( .A(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n6891) );
  AOI22_X1 U4301 ( .A1(n4106), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4134), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4302 ( .A1(n4081), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n5301), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4303 ( .A1(n4135), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3441) );
  AOI22_X1 U4304 ( .A1(n4108), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3440) );
  NAND4_X1 U4305 ( .A1(n3443), .A2(n3442), .A3(n3441), .A4(n3440), .ZN(n3444)
         );
  AOI22_X1 U4306 ( .A1(n3632), .A2(n3453), .B1(INSTQUEUE_REG_0__3__SCAN_IN), 
        .B2(n3625), .ZN(n3446) );
  NAND2_X1 U4307 ( .A1(n3449), .A2(n3448), .ZN(n3450) );
  NAND2_X1 U4308 ( .A1(n3450), .A2(n4557), .ZN(n3451) );
  NAND2_X1 U4309 ( .A1(n3452), .A2(n3453), .ZN(n3497) );
  OAI211_X1 U4310 ( .C1(n3453), .C2(n3452), .A(n3497), .B(n6571), .ZN(n3454)
         );
  INV_X1 U4311 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3455) );
  XNOR2_X1 U4312 ( .A(n3456), .B(n3455), .ZN(n4674) );
  NAND2_X1 U4313 ( .A1(n4675), .A2(n4674), .ZN(n3458) );
  NAND2_X1 U4314 ( .A1(n3456), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3457)
         );
  NAND2_X1 U4315 ( .A1(n3458), .A2(n3457), .ZN(n4856) );
  AOI22_X1 U4316 ( .A1(n4135), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4134), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3462) );
  AOI22_X1 U4317 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4138), .B1(n4086), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3461) );
  AOI22_X1 U4318 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n3306), .B1(n4107), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3460) );
  AOI22_X1 U4319 ( .A1(n4106), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3459) );
  NAND4_X1 U4320 ( .A1(n3462), .A2(n3461), .A3(n3460), .A4(n3459), .ZN(n3468)
         );
  AOI22_X1 U4321 ( .A1(n4081), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n5301), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3466) );
  AOI22_X1 U4322 ( .A1(n3120), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U4323 ( .A1(n3439), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4324 ( .A1(n4055), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3463) );
  NAND4_X1 U4325 ( .A1(n3466), .A2(n3465), .A3(n3464), .A4(n3463), .ZN(n3467)
         );
  NAND2_X1 U4326 ( .A1(n3632), .A2(n3495), .ZN(n3470) );
  NAND2_X1 U4327 ( .A1(n3625), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3469) );
  NAND2_X1 U4328 ( .A1(n3470), .A2(n3469), .ZN(n3478) );
  XNOR2_X1 U4329 ( .A(n3477), .B(n3478), .ZN(n3677) );
  NAND2_X1 U4330 ( .A1(n3677), .A2(n3596), .ZN(n3473) );
  XNOR2_X1 U4331 ( .A(n3497), .B(n3495), .ZN(n3471) );
  NAND2_X1 U4332 ( .A1(n3471), .A2(n6571), .ZN(n3472) );
  NAND2_X1 U4333 ( .A1(n3473), .A2(n3472), .ZN(n3474) );
  INV_X1 U4334 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6761) );
  XNOR2_X1 U4335 ( .A(n3474), .B(n6761), .ZN(n4857) );
  NAND2_X1 U4336 ( .A1(n4856), .A2(n4857), .ZN(n3476) );
  NAND2_X1 U4337 ( .A1(n3474), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3475)
         );
  NAND2_X1 U4338 ( .A1(n3476), .A2(n3475), .ZN(n4705) );
  INV_X1 U4339 ( .A(n3477), .ZN(n3479) );
  NAND2_X1 U4340 ( .A1(n3479), .A2(n3478), .ZN(n3492) );
  INV_X1 U4341 ( .A(n3492), .ZN(n3491) );
  AOI22_X1 U4342 ( .A1(n4087), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4343 ( .A1(n3120), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4344 ( .A1(n4107), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3481) );
  AOI22_X1 U4345 ( .A1(n4138), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3480) );
  NAND4_X1 U4346 ( .A1(n3483), .A2(n3482), .A3(n3481), .A4(n3480), .ZN(n3489)
         );
  AOI22_X1 U4347 ( .A1(n4106), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4134), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3487) );
  AOI22_X1 U4348 ( .A1(n4081), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n5301), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3486) );
  AOI22_X1 U4349 ( .A1(n4135), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3485) );
  AOI22_X1 U4350 ( .A1(n4108), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3484) );
  NAND4_X1 U4351 ( .A1(n3487), .A2(n3486), .A3(n3485), .A4(n3484), .ZN(n3488)
         );
  OR2_X1 U4352 ( .A1(n3489), .A2(n3488), .ZN(n3498) );
  AOI22_X1 U4353 ( .A1(n3632), .A2(n3498), .B1(INSTQUEUE_REG_0__5__SCAN_IN), 
        .B2(n3625), .ZN(n3493) );
  NAND2_X1 U4354 ( .A1(n3492), .A2(n3493), .ZN(n3494) );
  AND2_X2 U4355 ( .A1(n3517), .A2(n3494), .ZN(n3780) );
  NAND2_X1 U4356 ( .A1(n3780), .A2(n3596), .ZN(n3501) );
  INV_X1 U4357 ( .A(n3495), .ZN(n3496) );
  NOR2_X1 U4358 ( .A1(n3497), .A2(n3496), .ZN(n3499) );
  NAND2_X1 U4359 ( .A1(n3499), .A2(n3498), .ZN(n3530) );
  NAND2_X1 U4360 ( .A1(n3501), .A2(n3500), .ZN(n3503) );
  INV_X1 U4361 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3502) );
  XNOR2_X1 U4362 ( .A(n3503), .B(n3502), .ZN(n4706) );
  NAND2_X1 U4363 ( .A1(n4705), .A2(n4706), .ZN(n3505) );
  NAND2_X1 U4364 ( .A1(n3503), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3504)
         );
  NAND2_X1 U4365 ( .A1(n3505), .A2(n3504), .ZN(n4664) );
  AOI22_X1 U4366 ( .A1(n4135), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4134), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3509) );
  AOI22_X1 U4367 ( .A1(n4128), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3508) );
  AOI22_X1 U4368 ( .A1(n3120), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3507) );
  AOI22_X1 U4369 ( .A1(n4055), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3506) );
  NAND4_X1 U4370 ( .A1(n3509), .A2(n3508), .A3(n3507), .A4(n3506), .ZN(n3515)
         );
  AOI22_X1 U4371 ( .A1(n4081), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n5301), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4372 ( .A1(n4138), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4373 ( .A1(n4106), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4374 ( .A1(n4108), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3510) );
  NAND4_X1 U4375 ( .A1(n3513), .A2(n3512), .A3(n3511), .A4(n3510), .ZN(n3514)
         );
  OR2_X1 U4376 ( .A1(n3515), .A2(n3514), .ZN(n3531) );
  AOI22_X1 U4377 ( .A1(n3632), .A2(n3531), .B1(n3625), .B2(
        INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3516) );
  INV_X1 U4378 ( .A(n3529), .ZN(n3541) );
  NAND2_X1 U4379 ( .A1(n3517), .A2(n3516), .ZN(n3779) );
  NAND3_X1 U4380 ( .A1(n3541), .A2(n3596), .A3(n3779), .ZN(n3520) );
  XNOR2_X1 U4381 ( .A(n3530), .B(n3531), .ZN(n3518) );
  NAND2_X1 U4382 ( .A1(n3518), .A2(n6571), .ZN(n3519) );
  NAND2_X1 U4383 ( .A1(n3520), .A2(n3519), .ZN(n3522) );
  INV_X1 U4384 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3521) );
  XNOR2_X1 U4385 ( .A(n3522), .B(n3521), .ZN(n4665) );
  NAND2_X1 U4386 ( .A1(n4664), .A2(n4665), .ZN(n3524) );
  NAND2_X1 U4387 ( .A1(n3522), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3523)
         );
  NAND2_X1 U4388 ( .A1(n3524), .A2(n3523), .ZN(n5057) );
  INV_X1 U4389 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3526) );
  NAND2_X1 U4390 ( .A1(n3632), .A2(n3542), .ZN(n3525) );
  OAI21_X1 U4391 ( .B1(n3526), .B2(n3597), .A(n3525), .ZN(n3527) );
  XNOR2_X2 U4392 ( .A(n3529), .B(n3528), .ZN(n4906) );
  NAND2_X1 U4393 ( .A1(n4906), .A2(n3596), .ZN(n3535) );
  INV_X1 U4394 ( .A(n3530), .ZN(n3532) );
  NAND2_X1 U4395 ( .A1(n3532), .A2(n3531), .ZN(n3544) );
  XNOR2_X1 U4396 ( .A(n3544), .B(n3542), .ZN(n3533) );
  NAND2_X1 U4397 ( .A1(n3533), .A2(n6571), .ZN(n3534) );
  NAND2_X1 U4398 ( .A1(n3535), .A2(n3534), .ZN(n3536) );
  INV_X1 U4399 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6361) );
  XNOR2_X1 U4400 ( .A(n3536), .B(n6361), .ZN(n5058) );
  NAND2_X1 U4401 ( .A1(n5057), .A2(n5058), .ZN(n3538) );
  NAND2_X1 U4402 ( .A1(n3536), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3537)
         );
  NAND2_X1 U4403 ( .A1(n3538), .A2(n3537), .ZN(n4924) );
  NOR2_X1 U4404 ( .A1(n3622), .A2(n3539), .ZN(n3540) );
  NAND2_X1 U4405 ( .A1(n6571), .A2(n3542), .ZN(n3543) );
  OR2_X1 U4406 ( .A1(n3544), .A2(n3543), .ZN(n3545) );
  NAND2_X1 U4407 ( .A1(n3552), .A2(n3545), .ZN(n3546) );
  INV_X1 U4408 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4230) );
  XNOR2_X1 U4409 ( .A(n3546), .B(n4230), .ZN(n4925) );
  NAND2_X1 U4410 ( .A1(n4924), .A2(n4925), .ZN(n3548) );
  NAND2_X1 U4411 ( .A1(n3546), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3547)
         );
  INV_X1 U4412 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6749) );
  NOR2_X1 U4413 ( .A1(n3119), .A2(n6749), .ZN(n3549) );
  NAND2_X1 U4414 ( .A1(n3119), .A2(n6749), .ZN(n3550) );
  INV_X1 U4415 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5126) );
  AND2_X1 U4416 ( .A1(n3119), .A2(n5126), .ZN(n5116) );
  NAND2_X1 U4417 ( .A1(n3556), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5117) );
  INV_X1 U4418 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6882) );
  NAND2_X1 U4419 ( .A1(n3119), .A2(n6882), .ZN(n5221) );
  NAND2_X1 U4420 ( .A1(n5220), .A2(n5221), .ZN(n3553) );
  NAND2_X1 U4421 ( .A1(n3556), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5222) );
  NAND2_X1 U4422 ( .A1(n3553), .A2(n5222), .ZN(n5227) );
  INV_X1 U4423 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6851) );
  NAND2_X1 U4424 ( .A1(n3119), .A2(n6851), .ZN(n3554) );
  NAND2_X1 U4425 ( .A1(n3556), .A2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3555) );
  INV_X1 U4426 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4311) );
  XNOR2_X1 U4427 ( .A(n3552), .B(n4311), .ZN(n5598) );
  XNOR2_X1 U4428 ( .A(n3119), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5579)
         );
  NAND2_X1 U4429 ( .A1(n3556), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5576) );
  INV_X1 U4430 ( .A(n5560), .ZN(n3557) );
  NAND2_X1 U4431 ( .A1(n3119), .A2(n4311), .ZN(n5586) );
  INV_X1 U4432 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U4433 ( .A1(n3119), .A2(n6056), .ZN(n3558) );
  INV_X1 U4434 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6921) );
  NAND2_X1 U4435 ( .A1(n3119), .A2(n6921), .ZN(n3559) );
  INV_X1 U4436 ( .A(n5571), .ZN(n3563) );
  INV_X1 U4437 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5703) );
  NAND2_X1 U4438 ( .A1(n3563), .A2(n3562), .ZN(n5557) );
  INV_X1 U4439 ( .A(n5557), .ZN(n3565) );
  NAND2_X1 U4440 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3564) );
  NAND2_X1 U4441 ( .A1(n3565), .A2(n3144), .ZN(n5521) );
  NAND2_X1 U4442 ( .A1(n3556), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6001) );
  OAI21_X1 U4443 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n3556), .ZN(n3566) );
  AND2_X1 U4444 ( .A1(n6001), .A2(n3566), .ZN(n3567) );
  NAND2_X1 U4445 ( .A1(n5521), .A2(n3567), .ZN(n3568) );
  INV_X1 U4446 ( .A(n3568), .ZN(n5689) );
  INV_X1 U4447 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6854) );
  NOR2_X1 U4448 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5663) );
  NOR2_X1 U4449 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5648) );
  INV_X1 U4450 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n6799) );
  NAND3_X1 U4451 ( .A1(n5663), .A2(n5648), .A3(n6799), .ZN(n3571) );
  AND2_X1 U4452 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5647) );
  AND2_X1 U4453 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5681) );
  AND2_X1 U4454 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4328) );
  AND3_X1 U4455 ( .A1(n5647), .A2(n5681), .A3(n4328), .ZN(n4312) );
  NAND2_X1 U4456 ( .A1(n3568), .A2(n4312), .ZN(n3569) );
  NAND2_X1 U4457 ( .A1(n3569), .A2(n3119), .ZN(n3570) );
  XNOR2_X1 U4458 ( .A(n3119), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5989)
         );
  INV_X1 U4459 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n6020) );
  NAND2_X1 U4460 ( .A1(n3119), .A2(n6020), .ZN(n3572) );
  NAND2_X2 U4461 ( .A1(n4338), .A2(n3572), .ZN(n5514) );
  INV_X1 U4462 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5512) );
  AND2_X1 U4463 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5622) );
  INV_X1 U4464 ( .A(n3126), .ZN(n3574) );
  NOR2_X1 U4465 ( .A1(n3575), .A2(n3574), .ZN(n3579) );
  NOR2_X1 U4466 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5623) );
  NAND2_X1 U4467 ( .A1(n3577), .A2(n3576), .ZN(n3578) );
  NOR2_X1 U4468 ( .A1(n3579), .A2(n3578), .ZN(n3580) );
  INV_X1 U4469 ( .A(n3580), .ZN(n3585) );
  INV_X1 U4470 ( .A(n5489), .ZN(n3581) );
  NOR3_X1 U4471 ( .A1(n3581), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n3576), 
        .ZN(n3582) );
  INV_X1 U4472 ( .A(n3582), .ZN(n3584) );
  NAND2_X1 U4473 ( .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5605) );
  INV_X1 U4474 ( .A(n5605), .ZN(n5604) );
  NAND2_X1 U4475 ( .A1(n3126), .A2(n5604), .ZN(n3583) );
  INV_X1 U4476 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6063) );
  NAND2_X1 U4477 ( .A1(n6411), .A2(n3132), .ZN(n3603) );
  INV_X1 U4478 ( .A(n3603), .ZN(n3600) );
  XNOR2_X1 U4479 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3598) );
  NAND2_X1 U4480 ( .A1(n3600), .A2(n3598), .ZN(n3587) );
  NAND2_X1 U4481 ( .A1(n6948), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3586) );
  NAND2_X1 U4482 ( .A1(n3587), .A2(n3586), .ZN(n3614) );
  XNOR2_X1 U4483 ( .A(n5317), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3613)
         );
  INV_X1 U4484 ( .A(n3613), .ZN(n3588) );
  NAND2_X1 U4485 ( .A1(n3614), .A2(n3588), .ZN(n3590) );
  NAND2_X1 U4486 ( .A1(n6557), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3589) );
  NAND2_X1 U4487 ( .A1(n3590), .A2(n3589), .ZN(n3621) );
  INV_X1 U4488 ( .A(n3621), .ZN(n3591) );
  XNOR2_X1 U4489 ( .A(n5304), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3620)
         );
  NOR2_X1 U4490 ( .A1(n3591), .A2(n3620), .ZN(n3592) );
  AOI21_X1 U4491 ( .B1(n6563), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3592), 
        .ZN(n3593) );
  OAI222_X1 U4492 ( .A1(n6063), .A2(n3593), .B1(n6063), .B2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C1(n3593), .C2(
        INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n4173) );
  INV_X1 U4493 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6561) );
  NAND2_X1 U4494 ( .A1(n3593), .A2(n6063), .ZN(n3594) );
  AOI22_X1 U4495 ( .A1(n4177), .A2(n3625), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6585), .ZN(n3630) );
  INV_X1 U4496 ( .A(n4177), .ZN(n3595) );
  AOI21_X1 U4497 ( .B1(n3606), .B2(n3596), .A(n3595), .ZN(n3629) );
  NOR2_X1 U4498 ( .A1(n3597), .A2(n3622), .ZN(n3633) );
  INV_X1 U4499 ( .A(n3633), .ZN(n3608) );
  INV_X1 U4500 ( .A(n3598), .ZN(n3599) );
  XNOR2_X1 U4501 ( .A(n3600), .B(n3599), .ZN(n4176) );
  AND2_X1 U4502 ( .A1(n3271), .A2(n4653), .ZN(n3602) );
  OAI21_X1 U4503 ( .B1(n3132), .B2(n6411), .A(n3603), .ZN(n3605) );
  OAI21_X1 U4504 ( .B1(n3257), .B2(n3605), .A(n5203), .ZN(n3604) );
  OAI211_X1 U4505 ( .C1(n3608), .C2(n4176), .A(n3624), .B(n3604), .ZN(n3611)
         );
  NOR2_X1 U4506 ( .A1(n3606), .A2(n3605), .ZN(n3607) );
  OAI21_X1 U4507 ( .B1(n3612), .B2(n4176), .A(n3607), .ZN(n3609) );
  NAND2_X1 U4508 ( .A1(n3609), .A2(n3608), .ZN(n3610) );
  NAND2_X1 U4509 ( .A1(n3611), .A2(n3610), .ZN(n3619) );
  NAND3_X1 U4510 ( .A1(n3612), .A2(STATE2_REG_0__SCAN_IN), .A3(n4176), .ZN(
        n3618) );
  XNOR2_X1 U4511 ( .A(n3614), .B(n3613), .ZN(n4175) );
  INV_X1 U4512 ( .A(n4175), .ZN(n3616) );
  INV_X1 U4513 ( .A(n3624), .ZN(n3615) );
  AOI21_X1 U4514 ( .B1(n3625), .B2(n3616), .A(n3615), .ZN(n3617) );
  NAND2_X1 U4515 ( .A1(n3632), .A2(n4175), .ZN(n3623) );
  AOI22_X1 U4516 ( .A1(n3619), .A2(n3618), .B1(n3617), .B2(n3623), .ZN(n3627)
         );
  XNOR2_X1 U4517 ( .A(n3621), .B(n3620), .ZN(n4174) );
  OAI22_X1 U4518 ( .A1(n3624), .A2(n3623), .B1(n4174), .B2(n3622), .ZN(n3626)
         );
  AOI222_X1 U4519 ( .A1(n3630), .A2(n3629), .B1(n3630), .B2(n3628), .C1(n3629), 
        .C2(n3628), .ZN(n3631) );
  AOI21_X1 U4520 ( .B1(n3632), .B2(n4173), .A(n3631), .ZN(n3635) );
  AND2_X1 U4521 ( .A1(n4173), .A2(n3633), .ZN(n3634) );
  AND2_X1 U4522 ( .A1(n3636), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6583) );
  NAND2_X1 U4523 ( .A1(n4579), .A2(n4574), .ZN(n3637) );
  OR2_X1 U4524 ( .A1(n3638), .A2(n3637), .ZN(n5281) );
  NAND2_X1 U4525 ( .A1(n5281), .A2(n4296), .ZN(n3640) );
  NAND2_X1 U4526 ( .A1(n3640), .A2(n3639), .ZN(n3641) );
  NOR2_X1 U4527 ( .A1(n3641), .A2(n4302), .ZN(n4189) );
  AND2_X1 U4528 ( .A1(n4189), .A2(n3257), .ZN(n6537) );
  NAND2_X1 U4529 ( .A1(n4196), .A2(n6339), .ZN(n4167) );
  INV_X1 U4530 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n4606) );
  NOR2_X2 U4531 ( .A1(n4611), .A2(n4606), .ZN(n4905) );
  NAND2_X1 U4532 ( .A1(n4556), .A2(n4905), .ZN(n3646) );
  INV_X1 U4533 ( .A(n4479), .ZN(n4482) );
  AND2_X1 U4534 ( .A1(n4482), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3670) );
  INV_X1 U4535 ( .A(EAX_REG_1__SCAN_IN), .ZN(n3643) );
  OAI22_X1 U4536 ( .A1(n4097), .A2(n3643), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5099), .ZN(n3644) );
  AOI21_X1 U4537 ( .B1(n3670), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3644), 
        .ZN(n3645) );
  INV_X1 U4538 ( .A(n3647), .ZN(n3648) );
  AOI21_X1 U4539 ( .B1(n5735), .B2(n3648), .A(n6480), .ZN(n4387) );
  NAND2_X1 U4540 ( .A1(n6474), .A2(n4905), .ZN(n3653) );
  INV_X1 U4541 ( .A(EAX_REG_0__SCAN_IN), .ZN(n3650) );
  INV_X1 U4542 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n5215) );
  OAI22_X1 U4543 ( .A1(n4097), .A2(n3650), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5215), .ZN(n3651) );
  AOI21_X1 U4544 ( .B1(n3670), .B2(n3132), .A(n3651), .ZN(n3652) );
  NAND2_X1 U4545 ( .A1(n3653), .A2(n3652), .ZN(n4386) );
  NAND2_X1 U4546 ( .A1(n4387), .A2(n4386), .ZN(n4389) );
  NOR2_X2 U4547 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n5193) );
  OR2_X1 U4548 ( .A1(n4386), .A2(n4127), .ZN(n3654) );
  NAND2_X1 U4549 ( .A1(n4389), .A2(n3654), .ZN(n4461) );
  NAND2_X1 U4550 ( .A1(n4555), .A2(n4905), .ZN(n3655) );
  NAND2_X1 U4551 ( .A1(n6480), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3824) );
  NAND2_X1 U4552 ( .A1(n3655), .A2(n3824), .ZN(n3660) );
  INV_X1 U4553 ( .A(n3670), .ZN(n3658) );
  OAI21_X1 U4554 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3664), .ZN(n6334) );
  INV_X1 U4555 ( .A(n3824), .ZN(n4343) );
  AOI22_X1 U4556 ( .A1(n5193), .A2(n6334), .B1(n4343), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3657) );
  NAND2_X1 U4557 ( .A1(n4344), .A2(EAX_REG_2__SCAN_IN), .ZN(n3656) );
  OAI211_X1 U4558 ( .C1(n3658), .C2(n5317), .A(n3657), .B(n3656), .ZN(n4398)
         );
  NAND2_X1 U4559 ( .A1(n4399), .A2(n4398), .ZN(n3662) );
  NAND2_X1 U4560 ( .A1(n3660), .A2(n3659), .ZN(n3661) );
  INV_X1 U4561 ( .A(EAX_REG_3__SCAN_IN), .ZN(n3667) );
  OAI21_X1 U4562 ( .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n3665), .A(n3672), 
        .ZN(n6243) );
  AOI22_X1 U4563 ( .A1(n5193), .A2(n6243), .B1(n4343), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3666) );
  OAI21_X1 U4564 ( .B1(n4097), .B2(n3667), .A(n3666), .ZN(n3668) );
  AOI21_X1 U4565 ( .B1(n3670), .B2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n3668), 
        .ZN(n3669) );
  OAI21_X1 U4566 ( .B1(n4717), .B2(n3843), .A(n3669), .ZN(n4392) );
  NAND2_X1 U4567 ( .A1(n3670), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3675) );
  AOI21_X1 U4568 ( .B1(n6219), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3671) );
  AOI21_X1 U4569 ( .B1(n4344), .B2(EAX_REG_4__SCAN_IN), .A(n3671), .ZN(n3674)
         );
  NAND2_X1 U4570 ( .A1(n6219), .A2(n3672), .ZN(n3673) );
  INV_X1 U4571 ( .A(n3680), .ZN(n3782) );
  AND2_X1 U4572 ( .A1(n3673), .A2(n3782), .ZN(n5052) );
  AOI22_X1 U4573 ( .A1(n3675), .A2(n3674), .B1(n5193), .B2(n5052), .ZN(n3676)
         );
  AOI21_X1 U4574 ( .B1(n3677), .B2(n4905), .A(n3676), .ZN(n4492) );
  INV_X1 U4575 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n6914) );
  INV_X1 U4576 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6825) );
  AOI21_X1 U4577 ( .B1(n6914), .B2(n3696), .A(n3822), .ZN(n6134) );
  NAND2_X1 U4578 ( .A1(n6134), .A2(n5193), .ZN(n3683) );
  INV_X1 U4579 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5038) );
  INV_X1 U4580 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6072) );
  OAI21_X1 U4581 ( .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n6072), .A(n6480), 
        .ZN(n3681) );
  OAI21_X1 U4582 ( .B1(n4097), .B2(n5038), .A(n3681), .ZN(n3682) );
  NAND2_X1 U4583 ( .A1(n3683), .A2(n3682), .ZN(n3695) );
  AOI22_X1 U4584 ( .A1(n4135), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3687) );
  AOI22_X1 U4585 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3120), .B1(n4086), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3686) );
  AOI22_X1 U4586 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n5301), .B1(n4108), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3685) );
  AOI22_X1 U4587 ( .A1(n4138), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3684) );
  NAND4_X1 U4588 ( .A1(n3687), .A2(n3686), .A3(n3685), .A4(n3684), .ZN(n3693)
         );
  AOI22_X1 U4589 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n4055), .B1(n4128), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3691) );
  AOI22_X1 U4590 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n4107), .B1(n3306), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3690) );
  AOI22_X1 U4591 ( .A1(n4134), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3689) );
  AOI22_X1 U4592 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n4081), .B1(n3121), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3688) );
  NAND4_X1 U4593 ( .A1(n3691), .A2(n3690), .A3(n3689), .A4(n3688), .ZN(n3692)
         );
  OAI21_X1 U4594 ( .B1(n3693), .B2(n3692), .A(n4905), .ZN(n3694) );
  NAND2_X1 U4595 ( .A1(n3695), .A2(n3694), .ZN(n5037) );
  OR2_X1 U4596 ( .A1(n3712), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3697)
         );
  NAND2_X1 U4597 ( .A1(n3697), .A2(n3696), .ZN(n6141) );
  AOI22_X1 U4598 ( .A1(n4138), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4134), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4599 ( .A1(n4055), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3700) );
  AOI22_X1 U4600 ( .A1(n3120), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4601 ( .A1(n4135), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3698) );
  NAND4_X1 U4602 ( .A1(n3701), .A2(n3700), .A3(n3699), .A4(n3698), .ZN(n3707)
         );
  AOI22_X1 U4603 ( .A1(n4128), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3705) );
  AOI22_X1 U4604 ( .A1(n4106), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3704) );
  AOI22_X1 U4605 ( .A1(n5301), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4606 ( .A1(n4081), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3702) );
  NAND4_X1 U4607 ( .A1(n3705), .A2(n3704), .A3(n3703), .A4(n3702), .ZN(n3706)
         );
  NOR2_X1 U4608 ( .A1(n3707), .A2(n3706), .ZN(n3710) );
  NAND2_X1 U4609 ( .A1(n4344), .A2(EAX_REG_11__SCAN_IN), .ZN(n3709) );
  NAND2_X1 U4610 ( .A1(n4343), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3708)
         );
  OAI211_X1 U4611 ( .C1(n3843), .C2(n3710), .A(n3709), .B(n3708), .ZN(n3711)
         );
  AOI21_X1 U4612 ( .B1(n6141), .B2(n5193), .A(n3711), .ZN(n5138) );
  AOI21_X1 U4613 ( .B1(n6825), .B2(n3713), .A(n3712), .ZN(n6154) );
  OR2_X1 U4614 ( .A1(n6154), .A2(n4127), .ZN(n3729) );
  AOI22_X1 U4615 ( .A1(n4135), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4616 ( .A1(n4087), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3716) );
  AOI22_X1 U4617 ( .A1(n3120), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4618 ( .A1(n4055), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3714) );
  NAND4_X1 U4619 ( .A1(n3717), .A2(n3716), .A3(n3715), .A4(n3714), .ZN(n3723)
         );
  AOI22_X1 U4620 ( .A1(n4138), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4621 ( .A1(n4134), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3720) );
  AOI22_X1 U4622 ( .A1(n5301), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4623 ( .A1(n4106), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3718) );
  NAND4_X1 U4624 ( .A1(n3721), .A2(n3720), .A3(n3719), .A4(n3718), .ZN(n3722)
         );
  NOR2_X1 U4625 ( .A1(n3723), .A2(n3722), .ZN(n3726) );
  NAND2_X1 U4626 ( .A1(n4344), .A2(EAX_REG_10__SCAN_IN), .ZN(n3725) );
  NAND2_X1 U4627 ( .A1(n4343), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3724)
         );
  OAI211_X1 U4628 ( .C1(n3843), .C2(n3726), .A(n3725), .B(n3724), .ZN(n3727)
         );
  INV_X1 U4629 ( .A(n3727), .ZN(n3728) );
  NOR2_X1 U4630 ( .A1(n5138), .A2(n5109), .ZN(n5035) );
  AND2_X1 U4631 ( .A1(n5037), .A2(n5035), .ZN(n3746) );
  INV_X1 U4632 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5087) );
  XNOR2_X1 U4633 ( .A(n3747), .B(n5087), .ZN(n6171) );
  OR2_X1 U4634 ( .A1(n6171), .A2(n4127), .ZN(n3745) );
  AOI22_X1 U4635 ( .A1(n4135), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4636 ( .A1(n3120), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3732) );
  AOI22_X1 U4637 ( .A1(n4107), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3731) );
  AOI22_X1 U4638 ( .A1(n5301), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3730) );
  NAND4_X1 U4639 ( .A1(n3733), .A2(n3732), .A3(n3731), .A4(n3730), .ZN(n3739)
         );
  AOI22_X1 U4640 ( .A1(n4138), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4641 ( .A1(n4087), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3736) );
  AOI22_X1 U4642 ( .A1(n4134), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4643 ( .A1(n4108), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3734) );
  NAND4_X1 U4644 ( .A1(n3737), .A2(n3736), .A3(n3735), .A4(n3734), .ZN(n3738)
         );
  NOR2_X1 U4645 ( .A1(n3739), .A2(n3738), .ZN(n3742) );
  NAND2_X1 U4646 ( .A1(n4344), .A2(EAX_REG_9__SCAN_IN), .ZN(n3741) );
  NAND2_X1 U4647 ( .A1(n4343), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3740)
         );
  OAI211_X1 U4648 ( .C1(n3843), .C2(n3742), .A(n3741), .B(n3740), .ZN(n3743)
         );
  INV_X1 U4649 ( .A(n3743), .ZN(n3744) );
  NAND2_X1 U4650 ( .A1(n3745), .A2(n3744), .ZN(n5033) );
  AOI21_X1 U4651 ( .B1(n6838), .B2(n3767), .A(n3747), .ZN(n6179) );
  OR2_X1 U4652 ( .A1(n6179), .A2(n4127), .ZN(n3763) );
  AOI22_X1 U4653 ( .A1(n4138), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4654 ( .A1(n4086), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4655 ( .A1(n4106), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3749) );
  AOI22_X1 U4656 ( .A1(n4081), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3748) );
  NAND4_X1 U4657 ( .A1(n3751), .A2(n3750), .A3(n3749), .A4(n3748), .ZN(n3757)
         );
  AOI22_X1 U4658 ( .A1(n4135), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4134), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4659 ( .A1(n3120), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4660 ( .A1(n5301), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3753) );
  AOI22_X1 U4661 ( .A1(n4055), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3752) );
  NAND4_X1 U4662 ( .A1(n3755), .A2(n3754), .A3(n3753), .A4(n3752), .ZN(n3756)
         );
  NOR2_X1 U4663 ( .A1(n3757), .A2(n3756), .ZN(n3760) );
  NAND2_X1 U4664 ( .A1(n4344), .A2(EAX_REG_8__SCAN_IN), .ZN(n3759) );
  NAND2_X1 U4665 ( .A1(n4343), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3758)
         );
  OAI211_X1 U4666 ( .C1(n3843), .C2(n3760), .A(n3759), .B(n3758), .ZN(n3761)
         );
  INV_X1 U4667 ( .A(n3761), .ZN(n3762) );
  NAND2_X1 U4668 ( .A1(n3763), .A2(n3762), .ZN(n4984) );
  NAND2_X1 U4669 ( .A1(n4906), .A2(n3765), .ZN(n3772) );
  INV_X1 U4670 ( .A(n3766), .ZN(n3770) );
  INV_X1 U4671 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4922) );
  OAI21_X1 U4672 ( .B1(n3774), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3767), 
        .ZN(n6199) );
  AOI22_X1 U4673 ( .A1(n6199), .A2(n5193), .B1(n4343), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3768) );
  OAI21_X1 U4674 ( .B1(n4097), .B2(n4922), .A(n3768), .ZN(n3769) );
  INV_X1 U4675 ( .A(n3769), .ZN(n4907) );
  NAND2_X1 U4676 ( .A1(n3772), .A2(n3771), .ZN(n3790) );
  NOR2_X1 U4677 ( .A1(n3781), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3773)
         );
  NOR2_X1 U4678 ( .A1(n3774), .A2(n3773), .ZN(n6202) );
  INV_X1 U4679 ( .A(EAX_REG_6__SCAN_IN), .ZN(n4853) );
  INV_X1 U4680 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3775) );
  OAI22_X1 U4681 ( .A1(n4097), .A2(n4853), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3775), .ZN(n3776) );
  NAND2_X1 U4682 ( .A1(n3776), .A2(n4127), .ZN(n3777) );
  OAI21_X1 U4683 ( .B1(n6202), .B2(n4127), .A(n3777), .ZN(n3778) );
  INV_X1 U4684 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3787) );
  INV_X1 U4685 ( .A(n3781), .ZN(n3785) );
  INV_X1 U4686 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3783) );
  NAND2_X1 U4687 ( .A1(n3783), .A2(n3782), .ZN(n3784) );
  NAND2_X1 U4688 ( .A1(n3785), .A2(n3784), .ZN(n6218) );
  AOI22_X1 U4689 ( .A1(n6218), .A2(n5193), .B1(n4343), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3786) );
  OAI21_X1 U4690 ( .B1(n4097), .B2(n3787), .A(n3786), .ZN(n3788) );
  XNOR2_X1 U4691 ( .A(n3822), .B(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6124)
         );
  INV_X1 U4692 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6305) );
  INV_X1 U4693 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3793) );
  OAI22_X1 U4694 ( .A1(n4097), .A2(n6305), .B1(n3824), .B2(n3793), .ZN(n3794)
         );
  AOI21_X1 U4695 ( .B1(n6124), .B2(n5193), .A(n3794), .ZN(n3808) );
  INV_X1 U4696 ( .A(n5599), .ZN(n3806) );
  AOI22_X1 U4697 ( .A1(n4128), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4698 ( .A1(n3120), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4699 ( .A1(n4107), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4700 ( .A1(n4138), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3795) );
  NAND4_X1 U4701 ( .A1(n3798), .A2(n3797), .A3(n3796), .A4(n3795), .ZN(n3804)
         );
  AOI22_X1 U4702 ( .A1(n4106), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4134), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4703 ( .A1(n4081), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n5301), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4704 ( .A1(n4135), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3800) );
  AOI22_X1 U4705 ( .A1(n4108), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3799) );
  NAND4_X1 U4706 ( .A1(n3802), .A2(n3801), .A3(n3800), .A4(n3799), .ZN(n3803)
         );
  OR2_X1 U4707 ( .A1(n3804), .A2(n3803), .ZN(n3805) );
  NAND2_X1 U4708 ( .A1(n3806), .A2(n3147), .ZN(n3810) );
  INV_X1 U4709 ( .A(EAX_REG_14__SCAN_IN), .ZN(n5106) );
  AOI22_X1 U4710 ( .A1(n4055), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3814) );
  AOI22_X1 U4711 ( .A1(n4107), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3813) );
  AOI22_X1 U4712 ( .A1(n4135), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3812) );
  AOI22_X1 U4713 ( .A1(n4138), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3811) );
  NAND4_X1 U4714 ( .A1(n3814), .A2(n3813), .A3(n3812), .A4(n3811), .ZN(n3820)
         );
  AOI22_X1 U4715 ( .A1(n4081), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n5301), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3818) );
  AOI22_X1 U4716 ( .A1(n3120), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3817) );
  AOI22_X1 U4717 ( .A1(n4134), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3816) );
  AOI22_X1 U4718 ( .A1(n4106), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3815) );
  NAND4_X1 U4719 ( .A1(n3818), .A2(n3817), .A3(n3816), .A4(n3815), .ZN(n3819)
         );
  OR2_X1 U4720 ( .A1(n3820), .A2(n3819), .ZN(n3821) );
  NAND2_X1 U4721 ( .A1(n4905), .A2(n3821), .ZN(n3827) );
  INV_X1 U4722 ( .A(n3828), .ZN(n3823) );
  XNOR2_X1 U4723 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n3823), .ZN(n6115)
         );
  INV_X1 U4724 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5590) );
  OAI22_X1 U4725 ( .A1(n6115), .A2(n4127), .B1(n3824), .B2(n5590), .ZN(n3825)
         );
  INV_X1 U4726 ( .A(n3825), .ZN(n3826) );
  OAI211_X1 U4727 ( .C1(n5106), .C2(n4097), .A(n3827), .B(n3826), .ZN(n5102)
         );
  INV_X1 U4728 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6977) );
  AOI21_X1 U4729 ( .B1(n6977), .B2(n3829), .A(n3875), .ZN(n5582) );
  OR2_X1 U4730 ( .A1(n5582), .A2(n4127), .ZN(n3846) );
  AOI22_X1 U4731 ( .A1(n4135), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4134), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3833) );
  AOI22_X1 U4732 ( .A1(n4106), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3832) );
  AOI22_X1 U4733 ( .A1(n4107), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4734 ( .A1(n4055), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3830) );
  NAND4_X1 U4735 ( .A1(n3833), .A2(n3832), .A3(n3831), .A4(n3830), .ZN(n3839)
         );
  AOI22_X1 U4736 ( .A1(n4138), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4087), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3837) );
  AOI22_X1 U4737 ( .A1(n3120), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3836) );
  AOI22_X1 U4738 ( .A1(n3439), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3835) );
  AOI22_X1 U4739 ( .A1(n5301), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3834) );
  NAND4_X1 U4740 ( .A1(n3837), .A2(n3836), .A3(n3835), .A4(n3834), .ZN(n3838)
         );
  NOR2_X1 U4741 ( .A1(n3839), .A2(n3838), .ZN(n3842) );
  NAND2_X1 U4742 ( .A1(n4344), .A2(EAX_REG_15__SCAN_IN), .ZN(n3841) );
  NAND2_X1 U4743 ( .A1(n4343), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3840)
         );
  OAI211_X1 U4744 ( .C1(n3843), .C2(n3842), .A(n3841), .B(n3840), .ZN(n3844)
         );
  INV_X1 U4745 ( .A(n3844), .ZN(n3845) );
  XNOR2_X1 U4746 ( .A(n3875), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6106)
         );
  AOI22_X1 U4747 ( .A1(n4055), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4748 ( .A1(n4135), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4749 ( .A1(n4106), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3849) );
  AOI22_X1 U4750 ( .A1(n4138), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3848) );
  NAND4_X1 U4751 ( .A1(n3851), .A2(n3850), .A3(n3849), .A4(n3848), .ZN(n3857)
         );
  AOI22_X1 U4752 ( .A1(n4081), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n5301), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4753 ( .A1(n3120), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3854) );
  AOI22_X1 U4754 ( .A1(n4107), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3853) );
  AOI22_X1 U4755 ( .A1(n4134), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3852) );
  NAND4_X1 U4756 ( .A1(n3855), .A2(n3854), .A3(n3853), .A4(n3852), .ZN(n3856)
         );
  NOR2_X2 U4757 ( .A1(n5281), .A2(n6585), .ZN(n4147) );
  OAI21_X1 U4758 ( .B1(n3857), .B2(n3856), .A(n4147), .ZN(n3859) );
  AOI22_X1 U4759 ( .A1(n4344), .A2(EAX_REG_16__SCAN_IN), .B1(n4343), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3858) );
  NAND2_X1 U4760 ( .A1(n3859), .A2(n3858), .ZN(n3860) );
  AOI21_X1 U4761 ( .B1(n6106), .B2(n5193), .A(n3860), .ZN(n5249) );
  AOI22_X1 U4762 ( .A1(n4135), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4134), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4763 ( .A1(n5301), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4764 ( .A1(n3120), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4128), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3862) );
  AOI22_X1 U4765 ( .A1(n4107), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3861) );
  NAND4_X1 U4766 ( .A1(n3864), .A2(n3863), .A3(n3862), .A4(n3861), .ZN(n3870)
         );
  AOI22_X1 U4767 ( .A1(n4138), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4768 ( .A1(n4106), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4769 ( .A1(n4108), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3866) );
  AOI22_X1 U4770 ( .A1(n4081), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3865) );
  NAND4_X1 U4771 ( .A1(n3868), .A2(n3867), .A3(n3866), .A4(n3865), .ZN(n3869)
         );
  OR2_X1 U4772 ( .A1(n3870), .A2(n3869), .ZN(n3871) );
  NAND2_X1 U4773 ( .A1(n4147), .A2(n3871), .ZN(n3879) );
  INV_X1 U4774 ( .A(EAX_REG_17__SCAN_IN), .ZN(n3873) );
  NAND2_X1 U4775 ( .A1(n6480), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3872)
         );
  OAI211_X1 U4776 ( .C1(n4097), .C2(n3873), .A(n4127), .B(n3872), .ZN(n3874)
         );
  INV_X1 U4777 ( .A(n3874), .ZN(n3878) );
  OAI21_X1 U4778 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3876), .A(n3909), 
        .ZN(n6100) );
  NOR2_X1 U4779 ( .A1(n6100), .A2(n4127), .ZN(n3877) );
  AOI21_X1 U4780 ( .B1(n3879), .B2(n3878), .A(n3877), .ZN(n6008) );
  NAND2_X1 U4781 ( .A1(n5246), .A2(n6008), .ZN(n5252) );
  AOI22_X1 U4782 ( .A1(n4087), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4783 ( .A1(n3120), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3882) );
  AOI22_X1 U4784 ( .A1(n4107), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4785 ( .A1(n4138), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3880) );
  NAND4_X1 U4786 ( .A1(n3883), .A2(n3882), .A3(n3881), .A4(n3880), .ZN(n3889)
         );
  AOI22_X1 U4787 ( .A1(n4106), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n4134), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3887) );
  AOI22_X1 U4788 ( .A1(n4081), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n5301), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4789 ( .A1(n4135), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4790 ( .A1(n4108), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3884) );
  NAND4_X1 U4791 ( .A1(n3887), .A2(n3886), .A3(n3885), .A4(n3884), .ZN(n3888)
         );
  OR2_X1 U4792 ( .A1(n3889), .A2(n3888), .ZN(n3890) );
  NAND2_X1 U4793 ( .A1(n4147), .A2(n3890), .ZN(n3893) );
  INV_X1 U4794 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5563) );
  AOI21_X1 U4795 ( .B1(n5563), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3891) );
  AOI21_X1 U4796 ( .B1(n4344), .B2(EAX_REG_18__SCAN_IN), .A(n3891), .ZN(n3892)
         );
  NAND2_X1 U4797 ( .A1(n3893), .A2(n3892), .ZN(n3895) );
  XNOR2_X1 U4798 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3909), .ZN(n5565)
         );
  NAND2_X1 U4799 ( .A1(n5193), .A2(n5565), .ZN(n3894) );
  NAND2_X1 U4800 ( .A1(n3895), .A2(n3894), .ZN(n5253) );
  NOR2_X2 U4801 ( .A1(n5252), .A2(n5253), .ZN(n5254) );
  AOI22_X1 U4802 ( .A1(n4134), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4803 ( .A1(n4138), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4804 ( .A1(n3120), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4805 ( .A1(n4107), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3896) );
  NAND4_X1 U4806 ( .A1(n3899), .A2(n3898), .A3(n3897), .A4(n3896), .ZN(n3905)
         );
  AOI22_X1 U4807 ( .A1(n4135), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3903) );
  AOI22_X1 U4808 ( .A1(n5301), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3902) );
  AOI22_X1 U4809 ( .A1(n4106), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3901) );
  AOI22_X1 U4810 ( .A1(n4128), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3900) );
  NAND4_X1 U4811 ( .A1(n3903), .A2(n3902), .A3(n3901), .A4(n3900), .ZN(n3904)
         );
  OR2_X1 U4812 ( .A1(n3905), .A2(n3904), .ZN(n3908) );
  INV_X1 U4813 ( .A(EAX_REG_19__SCAN_IN), .ZN(n5071) );
  OAI21_X1 U4814 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n6072), .A(n6480), 
        .ZN(n3906) );
  OAI21_X1 U4815 ( .B1(n4097), .B2(n5071), .A(n3906), .ZN(n3907) );
  AOI21_X1 U4816 ( .B1(n4147), .B2(n3908), .A(n3907), .ZN(n3912) );
  OAI21_X1 U4817 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n3910), .A(n3944), 
        .ZN(n6000) );
  NOR2_X1 U4818 ( .A1(n6000), .A2(n4127), .ZN(n3911) );
  AND2_X2 U4819 ( .A1(n5254), .A2(n3913), .ZN(n5440) );
  AOI22_X1 U4820 ( .A1(n4138), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4821 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n3348), .B1(n3306), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4822 ( .A1(n4135), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4823 ( .A1(n4081), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3914) );
  NAND4_X1 U4824 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n3914), .ZN(n3923)
         );
  AOI22_X1 U4825 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4106), .B1(n4134), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3921) );
  AOI22_X1 U4826 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n3120), .B1(n4086), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3920) );
  AOI22_X1 U4827 ( .A1(n5301), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3919) );
  AOI22_X1 U4828 ( .A1(n4087), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3918) );
  NAND4_X1 U4829 ( .A1(n3921), .A2(n3920), .A3(n3919), .A4(n3918), .ZN(n3922)
         );
  OR2_X1 U4830 ( .A1(n3923), .A2(n3922), .ZN(n3924) );
  NAND2_X1 U4831 ( .A1(n4147), .A2(n3924), .ZN(n3930) );
  INV_X1 U4832 ( .A(EAX_REG_20__SCAN_IN), .ZN(n3926) );
  NAND2_X1 U4833 ( .A1(n6480), .A2(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n3925)
         );
  OAI211_X1 U4834 ( .C1(n4097), .C2(n3926), .A(n4127), .B(n3925), .ZN(n3927)
         );
  INV_X1 U4835 ( .A(n3927), .ZN(n3929) );
  XNOR2_X1 U4836 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n3944), .ZN(n5972)
         );
  AND2_X1 U4837 ( .A1(n5972), .A2(n5193), .ZN(n3928) );
  AOI21_X1 U4838 ( .B1(n3930), .B2(n3929), .A(n3928), .ZN(n5441) );
  AND2_X2 U4839 ( .A1(n5440), .A2(n5441), .ZN(n5431) );
  AOI22_X1 U4840 ( .A1(n4081), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n5301), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3934) );
  AOI22_X1 U4841 ( .A1(n4087), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4842 ( .A1(n4134), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4843 ( .A1(n4106), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3931) );
  NAND4_X1 U4844 ( .A1(n3934), .A2(n3933), .A3(n3932), .A4(n3931), .ZN(n3940)
         );
  AOI22_X1 U4845 ( .A1(n3120), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4846 ( .A1(n3348), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4847 ( .A1(n4135), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3936) );
  AOI22_X1 U4848 ( .A1(n4138), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3935) );
  NAND4_X1 U4849 ( .A1(n3938), .A2(n3937), .A3(n3936), .A4(n3935), .ZN(n3939)
         );
  OR2_X1 U4850 ( .A1(n3940), .A2(n3939), .ZN(n3941) );
  NAND2_X1 U4851 ( .A1(n4147), .A2(n3941), .ZN(n3949) );
  INV_X1 U4852 ( .A(EAX_REG_21__SCAN_IN), .ZN(n6946) );
  OAI21_X1 U4853 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6072), .A(n6480), 
        .ZN(n3942) );
  OAI21_X1 U4854 ( .B1(n4097), .B2(n6946), .A(n3942), .ZN(n3943) );
  INV_X1 U4855 ( .A(n3943), .ZN(n3948) );
  OAI21_X1 U4856 ( .B1(n3946), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n3988), 
        .ZN(n5958) );
  NOR2_X1 U4857 ( .A1(n5958), .A2(n4127), .ZN(n3947) );
  AOI21_X1 U4858 ( .B1(n3949), .B2(n3948), .A(n3947), .ZN(n5432) );
  AOI22_X1 U4859 ( .A1(n4081), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n5301), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3953) );
  AOI22_X1 U4860 ( .A1(n4087), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4861 ( .A1(n4135), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4862 ( .A1(n4106), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3950) );
  NAND4_X1 U4863 ( .A1(n3953), .A2(n3952), .A3(n3951), .A4(n3950), .ZN(n3959)
         );
  AOI22_X1 U4864 ( .A1(n3354), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4865 ( .A1(n3120), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3348), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4866 ( .A1(n4134), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4867 ( .A1(n4138), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3954) );
  NAND4_X1 U4868 ( .A1(n3957), .A2(n3956), .A3(n3955), .A4(n3954), .ZN(n3958)
         );
  OAI21_X1 U4869 ( .B1(n3959), .B2(n3958), .A(n4147), .ZN(n3962) );
  INV_X1 U4870 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5541) );
  OAI21_X1 U4871 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5541), .A(n4127), .ZN(
        n3960) );
  AOI21_X1 U4872 ( .B1(n4344), .B2(EAX_REG_22__SCAN_IN), .A(n3960), .ZN(n3961)
         );
  NAND2_X1 U4873 ( .A1(n3962), .A2(n3961), .ZN(n3964) );
  XNOR2_X1 U4874 ( .A(n3988), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5946)
         );
  NAND2_X1 U4875 ( .A1(n5946), .A2(n5193), .ZN(n3963) );
  NAND2_X1 U4876 ( .A1(n3964), .A2(n3963), .ZN(n5429) );
  AOI22_X1 U4877 ( .A1(n4135), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4134), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4878 ( .A1(n4081), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4879 ( .A1(n4087), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U4880 ( .A1(n5301), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3965) );
  NAND4_X1 U4881 ( .A1(n3968), .A2(n3967), .A3(n3966), .A4(n3965), .ZN(n3974)
         );
  AOI22_X1 U4882 ( .A1(n4138), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4883 ( .A1(n3348), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4884 ( .A1(n4106), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3970) );
  AOI22_X1 U4885 ( .A1(n4108), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3969) );
  NAND4_X1 U4886 ( .A1(n3972), .A2(n3971), .A3(n3970), .A4(n3969), .ZN(n3973)
         );
  NOR2_X1 U4887 ( .A1(n3974), .A2(n3973), .ZN(n3995) );
  AOI22_X1 U4888 ( .A1(n4138), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n5301), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4889 ( .A1(n4128), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4890 ( .A1(n3120), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4891 ( .A1(n4134), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3975) );
  NAND4_X1 U4892 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(n3984)
         );
  AOI22_X1 U4893 ( .A1(n4135), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4894 ( .A1(n4107), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4895 ( .A1(n3397), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4896 ( .A1(n4081), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3979) );
  NAND4_X1 U4897 ( .A1(n3982), .A2(n3981), .A3(n3980), .A4(n3979), .ZN(n3983)
         );
  NOR2_X1 U4898 ( .A1(n3984), .A2(n3983), .ZN(n3994) );
  XOR2_X1 U4899 ( .A(n3995), .B(n3994), .Z(n3987) );
  INV_X1 U4900 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6791) );
  OAI21_X1 U4901 ( .B1(n6072), .B2(PHYADDRPOINTER_REG_23__SCAN_IN), .A(n6480), 
        .ZN(n3985) );
  OAI21_X1 U4902 ( .B1(n4097), .B2(n6791), .A(n3985), .ZN(n3986) );
  AOI21_X1 U4903 ( .B1(n4147), .B2(n3987), .A(n3986), .ZN(n3992) );
  OR2_X1 U4904 ( .A1(n3989), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n3990)
         );
  NAND2_X1 U4905 ( .A1(n4031), .A2(n3990), .ZN(n5945) );
  NOR2_X1 U4906 ( .A1(n5945), .A2(n4127), .ZN(n3991) );
  AND2_X2 U4907 ( .A1(n5416), .A2(n3993), .ZN(n5408) );
  NOR2_X1 U4908 ( .A1(n3995), .A2(n3994), .ZN(n4025) );
  AOI22_X1 U4909 ( .A1(n4128), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4055), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3999) );
  AOI22_X1 U4910 ( .A1(n3120), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4911 ( .A1(n3348), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4912 ( .A1(n4138), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3996) );
  NAND4_X1 U4913 ( .A1(n3999), .A2(n3998), .A3(n3997), .A4(n3996), .ZN(n4005)
         );
  AOI22_X1 U4914 ( .A1(n4106), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4134), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4003) );
  AOI22_X1 U4915 ( .A1(n4081), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n5301), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n4002) );
  AOI22_X1 U4916 ( .A1(n4135), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4001) );
  AOI22_X1 U4917 ( .A1(n4108), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4000) );
  NAND4_X1 U4918 ( .A1(n4003), .A2(n4002), .A3(n4001), .A4(n4000), .ZN(n4004)
         );
  OR2_X1 U4919 ( .A1(n4005), .A2(n4004), .ZN(n4024) );
  INV_X1 U4920 ( .A(n4024), .ZN(n4006) );
  XNOR2_X1 U4921 ( .A(n4025), .B(n4006), .ZN(n4007) );
  NAND2_X1 U4922 ( .A1(n4007), .A2(n4147), .ZN(n4013) );
  INV_X1 U4923 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4010) );
  INV_X1 U4924 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4030) );
  XNOR2_X1 U4925 ( .A(n4031), .B(n4030), .ZN(n5928) );
  NAND2_X1 U4926 ( .A1(n5928), .A2(n5193), .ZN(n4009) );
  NAND2_X1 U4927 ( .A1(n4343), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4008)
         );
  OAI211_X1 U4928 ( .C1(n4097), .C2(n4010), .A(n4009), .B(n4008), .ZN(n4011)
         );
  INV_X1 U4929 ( .A(n4011), .ZN(n4012) );
  NAND2_X1 U4930 ( .A1(n4013), .A2(n4012), .ZN(n5407) );
  AND2_X2 U4931 ( .A1(n5408), .A2(n5407), .ZN(n5409) );
  AOI22_X1 U4932 ( .A1(n4135), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4017) );
  AOI22_X1 U4933 ( .A1(n4128), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4016) );
  AOI22_X1 U4934 ( .A1(n3120), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4935 ( .A1(n3354), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4014) );
  NAND4_X1 U4936 ( .A1(n4017), .A2(n4016), .A3(n4015), .A4(n4014), .ZN(n4023)
         );
  AOI22_X1 U4937 ( .A1(n4138), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4938 ( .A1(n4134), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4020) );
  AOI22_X1 U4939 ( .A1(n5301), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4019) );
  AOI22_X1 U4940 ( .A1(n4081), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4018) );
  NAND4_X1 U4941 ( .A1(n4021), .A2(n4020), .A3(n4019), .A4(n4018), .ZN(n4022)
         );
  NOR2_X1 U4942 ( .A1(n4023), .A2(n4022), .ZN(n4038) );
  NAND2_X1 U4943 ( .A1(n4025), .A2(n4024), .ZN(n4037) );
  XNOR2_X1 U4944 ( .A(n4038), .B(n4037), .ZN(n4029) );
  INV_X1 U4945 ( .A(n4147), .ZN(n4124) );
  INV_X1 U4946 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6829) );
  OAI21_X1 U4947 ( .B1(n6072), .B2(PHYADDRPOINTER_REG_25__SCAN_IN), .A(n6480), 
        .ZN(n4026) );
  OAI21_X1 U4948 ( .B1(n4097), .B2(n6829), .A(n4026), .ZN(n4027) );
  INV_X1 U4949 ( .A(n4027), .ZN(n4028) );
  OAI21_X1 U4950 ( .B1(n4029), .B2(n4124), .A(n4028), .ZN(n4036) );
  INV_X1 U4951 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4032) );
  AND2_X1 U4952 ( .A1(n4033), .A2(n4032), .ZN(n4034) );
  OR2_X1 U4953 ( .A1(n4034), .A2(n4073), .ZN(n5995) );
  INV_X1 U4954 ( .A(n5995), .ZN(n5916) );
  NAND2_X1 U4955 ( .A1(n5916), .A2(n5193), .ZN(n4035) );
  AND2_X1 U4956 ( .A1(n4036), .A2(n4035), .ZN(n5400) );
  OR2_X1 U4957 ( .A1(n4038), .A2(n4037), .ZN(n4066) );
  AOI22_X1 U4958 ( .A1(n4128), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4042) );
  AOI22_X1 U4959 ( .A1(n3120), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U4960 ( .A1(n4135), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U4961 ( .A1(n4108), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4039) );
  NAND4_X1 U4962 ( .A1(n4042), .A2(n4041), .A3(n4040), .A4(n4039), .ZN(n4048)
         );
  AOI22_X1 U4963 ( .A1(n4106), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4134), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U4964 ( .A1(n4138), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U4965 ( .A1(n4086), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U4966 ( .A1(n5301), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4043) );
  NAND4_X1 U4967 ( .A1(n4046), .A2(n4045), .A3(n4044), .A4(n4043), .ZN(n4047)
         );
  NOR2_X1 U4968 ( .A1(n4048), .A2(n4047), .ZN(n4067) );
  XOR2_X1 U4969 ( .A(n4066), .B(n4067), .Z(n4049) );
  NAND2_X1 U4970 ( .A1(n4049), .A2(n4147), .ZN(n4052) );
  INV_X1 U4971 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5904) );
  OAI21_X1 U4972 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5904), .A(n4127), .ZN(
        n4050) );
  AOI21_X1 U4973 ( .B1(n4344), .B2(EAX_REG_26__SCAN_IN), .A(n4050), .ZN(n4051)
         );
  NAND2_X1 U4974 ( .A1(n4052), .A2(n4051), .ZN(n4054) );
  XNOR2_X1 U4975 ( .A(n4073), .B(n5904), .ZN(n5912) );
  NAND2_X1 U4976 ( .A1(n5912), .A2(n5193), .ZN(n4053) );
  NAND2_X1 U4977 ( .A1(n4054), .A2(n4053), .ZN(n5391) );
  NOR2_X2 U4978 ( .A1(n5402), .A2(n5391), .ZN(n5384) );
  AOI22_X1 U4979 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n4086), .B1(n4055), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4059) );
  AOI22_X1 U4980 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n3306), .B1(n4107), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U4981 ( .A1(n4135), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U4982 ( .A1(n4134), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4056) );
  NAND4_X1 U4983 ( .A1(n4059), .A2(n4058), .A3(n4057), .A4(n4056), .ZN(n4065)
         );
  AOI22_X1 U4984 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4138), .B1(n4081), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U4985 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n3120), .B1(n4128), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U4986 ( .A1(n4106), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U4987 ( .A1(n5301), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4060) );
  NAND4_X1 U4988 ( .A1(n4063), .A2(n4062), .A3(n4061), .A4(n4060), .ZN(n4064)
         );
  NOR2_X1 U4989 ( .A1(n4065), .A2(n4064), .ZN(n4080) );
  OR2_X1 U4990 ( .A1(n4067), .A2(n4066), .ZN(n4079) );
  XNOR2_X1 U4991 ( .A(n4080), .B(n4079), .ZN(n4072) );
  INV_X1 U4992 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4069) );
  NAND2_X1 U4993 ( .A1(n6480), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4068)
         );
  OAI211_X1 U4994 ( .C1(n4097), .C2(n4069), .A(n4127), .B(n4068), .ZN(n4070)
         );
  INV_X1 U4995 ( .A(n4070), .ZN(n4071) );
  OAI21_X1 U4996 ( .B1(n4072), .B2(n4124), .A(n4071), .ZN(n4077) );
  OR2_X1 U4997 ( .A1(n4074), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4075)
         );
  NAND2_X1 U4998 ( .A1(n4103), .A2(n4075), .ZN(n5896) );
  OR2_X1 U4999 ( .A1(n5896), .A2(n4127), .ZN(n4076) );
  NAND2_X1 U5000 ( .A1(n4077), .A2(n4076), .ZN(n5385) );
  AND2_X2 U5001 ( .A1(n5384), .A2(n4078), .ZN(n5377) );
  OR2_X1 U5002 ( .A1(n4080), .A2(n4079), .ZN(n4120) );
  AOI22_X1 U5003 ( .A1(n4134), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4081), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4085) );
  AOI22_X1 U5004 ( .A1(n3120), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5005 ( .A1(n4135), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U5006 ( .A1(n4138), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4082) );
  NAND4_X1 U5007 ( .A1(n4085), .A2(n4084), .A3(n4083), .A4(n4082), .ZN(n4093)
         );
  AOI22_X1 U5008 ( .A1(n4087), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4086), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4091) );
  AOI22_X1 U5009 ( .A1(n3348), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4090) );
  AOI22_X1 U5010 ( .A1(n4106), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U5011 ( .A1(n5301), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4108), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4088) );
  NAND4_X1 U5012 ( .A1(n4091), .A2(n4090), .A3(n4089), .A4(n4088), .ZN(n4092)
         );
  NOR2_X1 U5013 ( .A1(n4093), .A2(n4092), .ZN(n4121) );
  XOR2_X1 U5014 ( .A(n4120), .B(n4121), .Z(n4094) );
  NAND2_X1 U5015 ( .A1(n4094), .A2(n4147), .ZN(n4101) );
  INV_X1 U5016 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4096) );
  NAND2_X1 U5017 ( .A1(n4606), .A2(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4095)
         );
  OAI211_X1 U5018 ( .C1(n4097), .C2(n4096), .A(n4127), .B(n4095), .ZN(n4098)
         );
  INV_X1 U5019 ( .A(n4098), .ZN(n4100) );
  XNOR2_X1 U5020 ( .A(n4103), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5887)
         );
  AND2_X1 U5021 ( .A1(n5887), .A2(n5193), .ZN(n4099) );
  AOI21_X1 U5022 ( .B1(n4101), .B2(n4100), .A(n4099), .ZN(n5378) );
  INV_X1 U5023 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n4102) );
  INV_X1 U5024 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U5025 ( .A1(n4104), .A2(n5363), .ZN(n4105) );
  NAND2_X1 U5026 ( .A1(n4348), .A2(n4105), .ZN(n5494) );
  AOI22_X1 U5027 ( .A1(n4135), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4106), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4112) );
  AOI22_X1 U5028 ( .A1(n4128), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4136), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U5029 ( .A1(n3120), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4107), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U5030 ( .A1(n4108), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4109) );
  NAND4_X1 U5031 ( .A1(n4112), .A2(n4111), .A3(n4110), .A4(n4109), .ZN(n4119)
         );
  AOI22_X1 U5032 ( .A1(n4081), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n5301), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U5033 ( .A1(n3354), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3306), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4116) );
  AOI22_X1 U5034 ( .A1(n4134), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4115) );
  AOI22_X1 U5035 ( .A1(n4138), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4114) );
  NAND4_X1 U5036 ( .A1(n4117), .A2(n4116), .A3(n4115), .A4(n4114), .ZN(n4118)
         );
  OR2_X1 U5037 ( .A1(n4119), .A2(n4118), .ZN(n4145) );
  NOR2_X1 U5038 ( .A1(n4121), .A2(n4120), .ZN(n4146) );
  XNOR2_X1 U5039 ( .A(n4145), .B(n4146), .ZN(n4125) );
  AOI21_X1 U5040 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6480), .A(n5193), 
        .ZN(n4123) );
  NAND2_X1 U5041 ( .A1(n4344), .A2(EAX_REG_29__SCAN_IN), .ZN(n4122) );
  OAI211_X1 U5042 ( .C1(n4125), .C2(n4124), .A(n4123), .B(n4122), .ZN(n4126)
         );
  OAI21_X1 U5043 ( .B1(n4127), .B2(n5494), .A(n4126), .ZN(n5362) );
  XNOR2_X1 U5044 ( .A(n4348), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5355)
         );
  INV_X1 U5045 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5352) );
  AOI21_X1 U5046 ( .B1(n5352), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4152) );
  AOI22_X1 U5047 ( .A1(n4128), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U5048 ( .A1(n3348), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3391), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U5049 ( .A1(n4106), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3439), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5050 ( .A1(n4081), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4130) );
  NAND4_X1 U5051 ( .A1(n4133), .A2(n4132), .A3(n4131), .A4(n4130), .ZN(n4144)
         );
  AOI22_X1 U5052 ( .A1(n4135), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4134), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4142) );
  AOI22_X1 U5053 ( .A1(n3120), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n4136), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4141) );
  AOI22_X1 U5054 ( .A1(n5301), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3397), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4140) );
  AOI22_X1 U5055 ( .A1(n4138), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4113), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4139) );
  NAND4_X1 U5056 ( .A1(n4142), .A2(n4141), .A3(n4140), .A4(n4139), .ZN(n4143)
         );
  NOR2_X1 U5057 ( .A1(n4144), .A2(n4143), .ZN(n4150) );
  NAND2_X1 U5058 ( .A1(n4146), .A2(n4145), .ZN(n4149) );
  OAI21_X1 U5059 ( .B1(n4150), .B2(n4149), .A(n4147), .ZN(n4148) );
  AOI21_X1 U5060 ( .B1(n4150), .B2(n4149), .A(n4148), .ZN(n4151) );
  AOI211_X1 U5061 ( .C1(n4344), .C2(EAX_REG_30__SCAN_IN), .A(n4152), .B(n4151), 
        .ZN(n4153) );
  AOI21_X1 U5062 ( .B1(n5355), .B2(n5193), .A(n4153), .ZN(n4155) );
  OAI21_X2 U5063 ( .B1(n5361), .B2(n4155), .A(n4346), .ZN(n5350) );
  INV_X1 U5064 ( .A(n5350), .ZN(n4165) );
  AND2_X1 U5065 ( .A1(n6585), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5194) );
  NAND2_X1 U5066 ( .A1(n5194), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6593) );
  INV_X1 U5067 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6480) );
  OR2_X1 U5068 ( .A1(n6593), .A2(n6477), .ZN(n6344) );
  NAND2_X1 U5069 ( .A1(n4156), .A2(n6477), .ZN(n6672) );
  NAND2_X1 U5070 ( .A1(n6672), .A2(n6585), .ZN(n4157) );
  NAND2_X1 U5071 ( .A1(n6585), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4159) );
  NAND2_X1 U5072 ( .A1(n6072), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4158) );
  NAND2_X1 U5073 ( .A1(n4159), .A2(n4158), .ZN(n6340) );
  INV_X1 U5074 ( .A(n5355), .ZN(n4163) );
  INV_X1 U5075 ( .A(REIP_REG_30__SCAN_IN), .ZN(n4161) );
  NOR2_X1 U5076 ( .A1(n6187), .A2(n4161), .ZN(n4316) );
  AOI21_X1 U5077 ( .B1(n6341), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n4316), 
        .ZN(n4162) );
  OAI21_X1 U5078 ( .B1(n6335), .B2(n4163), .A(n4162), .ZN(n4164) );
  NAND2_X1 U5079 ( .A1(n4167), .A2(n4166), .ZN(U2956) );
  NOR2_X1 U5080 ( .A1(n5281), .A2(n3271), .ZN(n4298) );
  NAND2_X1 U5081 ( .A1(n4550), .A2(n4298), .ZN(n4508) );
  NAND2_X1 U5082 ( .A1(n4168), .A2(n5203), .ZN(n4169) );
  INV_X1 U5083 ( .A(n6571), .ZN(n6676) );
  MUX2_X1 U5084 ( .A(n4169), .B(n6676), .S(n3259), .Z(n4306) );
  NAND2_X1 U5085 ( .A1(n4306), .A2(n4189), .ZN(n4171) );
  NAND2_X1 U5086 ( .A1(n4171), .A2(n4170), .ZN(n4297) );
  INV_X1 U5087 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6606) );
  NAND2_X1 U5088 ( .A1(n4172), .A2(n6606), .ZN(n6601) );
  NAND2_X1 U5089 ( .A1(n4585), .A2(n6601), .ZN(n4180) );
  INV_X1 U5090 ( .A(n4173), .ZN(n4179) );
  NAND3_X1 U5091 ( .A1(n4176), .A2(n4175), .A3(n4174), .ZN(n4178) );
  AOI21_X1 U5092 ( .B1(n4179), .B2(n4178), .A(n4177), .ZN(n4363) );
  NOR2_X1 U5093 ( .A1(n4363), .A2(READY_N), .ZN(n4471) );
  NAND3_X1 U5094 ( .A1(n4180), .A2(n4471), .A3(n3220), .ZN(n4181) );
  NAND3_X1 U5095 ( .A1(n4508), .A2(n4297), .A3(n4181), .ZN(n4182) );
  NAND2_X1 U5096 ( .A1(n4182), .A2(n6583), .ZN(n4188) );
  INV_X1 U5097 ( .A(READY_N), .ZN(n6673) );
  INV_X1 U5098 ( .A(n6601), .ZN(n4635) );
  OR2_X1 U5099 ( .A1(n4585), .A2(n4635), .ZN(n5201) );
  NAND3_X1 U5100 ( .A1(n6572), .A2(n6673), .A3(n5201), .ZN(n4184) );
  NAND3_X1 U5101 ( .A1(n4184), .A2(n5203), .A3(n4479), .ZN(n4185) );
  NAND3_X1 U5102 ( .A1(n4632), .A2(n4186), .A3(n4185), .ZN(n4187) );
  INV_X1 U5103 ( .A(n6537), .ZN(n4193) );
  AND2_X1 U5104 ( .A1(n4189), .A2(n3129), .ZN(n4470) );
  INV_X1 U5105 ( .A(n4470), .ZN(n4518) );
  AND2_X4 U5106 ( .A1(n5203), .A2(n4585), .ZN(n5207) );
  NAND2_X1 U5107 ( .A1(n6572), .A2(n5207), .ZN(n4502) );
  OAI211_X1 U5108 ( .C1(n4381), .C2(n4198), .A(n4514), .B(n4502), .ZN(n4191)
         );
  INV_X1 U5109 ( .A(n4191), .ZN(n4192) );
  NAND3_X1 U5110 ( .A1(n4193), .A2(n4518), .A3(n4192), .ZN(n4194) );
  NAND2_X1 U5111 ( .A1(n4196), .A2(n4195), .ZN(n4337) );
  NAND2_X1 U5112 ( .A1(n6572), .A2(n6571), .ZN(n4197) );
  OAI21_X1 U5113 ( .B1(n4198), .B2(n4579), .A(n4197), .ZN(n4199) );
  NAND2_X1 U5114 ( .A1(n4318), .A2(n4199), .ZN(n6394) );
  OAI22_X1 U5115 ( .A1(n5331), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        EBX_REG_29__SCAN_IN), .B2(n5330), .ZN(n5324) );
  AND2_X2 U5116 ( .A1(n5444), .A2(n5207), .ZN(n4282) );
  INV_X1 U5117 ( .A(EBX_REG_1__SCAN_IN), .ZN(n4467) );
  NAND2_X1 U5118 ( .A1(n4282), .A2(n4467), .ZN(n4205) );
  INV_X1 U5119 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4201) );
  NAND2_X1 U5120 ( .A1(n4209), .A2(n4201), .ZN(n4203) );
  NAND2_X1 U5121 ( .A1(n5207), .A2(n4467), .ZN(n4202) );
  NAND3_X1 U5122 ( .A1(n4203), .A2(n4200), .A3(n4202), .ZN(n4204) );
  NAND2_X1 U5123 ( .A1(n4205), .A2(n4204), .ZN(n4208) );
  NAND2_X1 U5124 ( .A1(n4209), .A2(EBX_REG_0__SCAN_IN), .ZN(n4207) );
  INV_X1 U5125 ( .A(EBX_REG_0__SCAN_IN), .ZN(n6903) );
  NAND2_X1 U5126 ( .A1(n4200), .A2(n6903), .ZN(n4206) );
  NAND2_X1 U5127 ( .A1(n4207), .A2(n4206), .ZN(n4380) );
  XNOR2_X1 U5128 ( .A(n4208), .B(n4380), .ZN(n4464) );
  NAND2_X1 U5129 ( .A1(n4464), .A2(n5207), .ZN(n4465) );
  INV_X1 U5130 ( .A(n4209), .ZN(n4210) );
  NAND2_X1 U5131 ( .A1(n4210), .A2(n5330), .ZN(n4279) );
  NAND2_X1 U5132 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n5330), .ZN(n4211)
         );
  AND3_X2 U5133 ( .A1(n4212), .A2(n4279), .A3(n4211), .ZN(n4403) );
  NAND2_X1 U5134 ( .A1(n5207), .A2(n5323), .ZN(n4287) );
  NAND2_X1 U5135 ( .A1(n5323), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4215)
         );
  OAI211_X1 U5136 ( .C1(n5330), .C2(EBX_REG_3__SCAN_IN), .A(n4290), .B(n4215), 
        .ZN(n4216) );
  OAI21_X1 U5137 ( .B1(n4287), .B2(EBX_REG_3__SCAN_IN), .A(n4216), .ZN(n4394)
         );
  NAND2_X1 U5138 ( .A1(n4290), .A2(n6761), .ZN(n4218) );
  INV_X1 U5139 ( .A(EBX_REG_4__SCAN_IN), .ZN(n6982) );
  NAND2_X1 U5140 ( .A1(n5207), .A2(n6982), .ZN(n4217) );
  NAND3_X1 U5141 ( .A1(n4218), .A2(n5323), .A3(n4217), .ZN(n4219) );
  OAI21_X1 U5142 ( .B1(n4291), .B2(EBX_REG_4__SCAN_IN), .A(n4219), .ZN(n4496)
         );
  NAND2_X1 U5143 ( .A1(n4497), .A2(n4496), .ZN(n4488) );
  NAND2_X1 U5144 ( .A1(n5323), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4220)
         );
  OAI211_X1 U5145 ( .C1(EBX_REG_5__SCAN_IN), .C2(n5330), .A(n4290), .B(n4220), 
        .ZN(n4221) );
  OAI21_X1 U5146 ( .B1(n4287), .B2(EBX_REG_5__SCAN_IN), .A(n4221), .ZN(n4490)
         );
  MUX2_X1 U5147 ( .A(n4287), .B(n5323), .S(EBX_REG_7__SCAN_IN), .Z(n4225) );
  NAND2_X1 U5148 ( .A1(n6361), .A2(n4301), .ZN(n4224) );
  AND2_X1 U5149 ( .A1(n4225), .A2(n4224), .ZN(n4912) );
  MUX2_X1 U5150 ( .A(n4291), .B(n4290), .S(EBX_REG_6__SCAN_IN), .Z(n4228) );
  NAND2_X1 U5151 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n5330), .ZN(n4226)
         );
  AND2_X1 U5152 ( .A1(n4279), .A2(n4226), .ZN(n4227) );
  NAND2_X1 U5153 ( .A1(n4228), .A2(n4227), .ZN(n4913) );
  NAND2_X1 U5154 ( .A1(n4912), .A2(n4913), .ZN(n4229) );
  NOR2_X2 U5155 ( .A1(n4489), .A2(n4229), .ZN(n4928) );
  NAND2_X1 U5156 ( .A1(n4290), .A2(n4230), .ZN(n4233) );
  INV_X1 U5157 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4231) );
  NAND2_X1 U5158 ( .A1(n5207), .A2(n4231), .ZN(n4232) );
  NAND3_X1 U5159 ( .A1(n4233), .A2(n5323), .A3(n4232), .ZN(n4234) );
  OAI21_X1 U5160 ( .B1(n4291), .B2(EBX_REG_8__SCAN_IN), .A(n4234), .ZN(n4927)
         );
  INV_X1 U5161 ( .A(n4287), .ZN(n4274) );
  INV_X1 U5162 ( .A(EBX_REG_9__SCAN_IN), .ZN(n6767) );
  NAND2_X1 U5163 ( .A1(n4274), .A2(n6767), .ZN(n4237) );
  NAND2_X1 U5164 ( .A1(n5323), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4235)
         );
  OAI211_X1 U5165 ( .C1(n5330), .C2(EBX_REG_9__SCAN_IN), .A(n4290), .B(n4235), 
        .ZN(n4236) );
  MUX2_X1 U5166 ( .A(n4291), .B(n4290), .S(EBX_REG_10__SCAN_IN), .Z(n4239) );
  NAND2_X1 U5167 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n5330), .ZN(n4238) );
  OR2_X2 U5168 ( .A1(n4990), .A2(n5113), .ZN(n5144) );
  NAND2_X1 U5169 ( .A1(n5323), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n4240) );
  OAI211_X1 U5170 ( .C1(n5330), .C2(EBX_REG_11__SCAN_IN), .A(n4290), .B(n4240), 
        .ZN(n4241) );
  OAI21_X1 U5171 ( .B1(n4287), .B2(EBX_REG_11__SCAN_IN), .A(n4241), .ZN(n5143)
         );
  INV_X1 U5172 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6277) );
  NAND2_X1 U5173 ( .A1(n4274), .A2(n6277), .ZN(n4244) );
  NAND2_X1 U5174 ( .A1(n5323), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n4242) );
  OAI211_X1 U5175 ( .C1(n5330), .C2(EBX_REG_13__SCAN_IN), .A(n4290), .B(n4242), 
        .ZN(n4243) );
  AND2_X1 U5176 ( .A1(n4244), .A2(n4243), .ZN(n5713) );
  INV_X1 U5177 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6283) );
  NAND2_X1 U5178 ( .A1(n4282), .A2(n6283), .ZN(n4248) );
  NAND2_X1 U5179 ( .A1(n4290), .A2(n6851), .ZN(n4246) );
  NAND2_X1 U5180 ( .A1(n5207), .A2(n6283), .ZN(n4245) );
  NAND3_X1 U5181 ( .A1(n4246), .A2(n5323), .A3(n4245), .ZN(n4247) );
  NAND2_X1 U5182 ( .A1(n4248), .A2(n4247), .ZN(n5714) );
  NAND2_X1 U5183 ( .A1(n5713), .A2(n5714), .ZN(n4249) );
  MUX2_X1 U5184 ( .A(n4291), .B(n4290), .S(EBX_REG_14__SCAN_IN), .Z(n4252) );
  NAND2_X1 U5185 ( .A1(n5330), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4250) );
  AND2_X1 U5186 ( .A1(n4279), .A2(n4250), .ZN(n4251) );
  NAND2_X1 U5187 ( .A1(n4252), .A2(n4251), .ZN(n5104) );
  NAND2_X1 U5188 ( .A1(n5716), .A2(n5104), .ZN(n5134) );
  NAND2_X1 U5189 ( .A1(n5323), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n4253) );
  OAI211_X1 U5190 ( .C1(n5330), .C2(EBX_REG_15__SCAN_IN), .A(n4290), .B(n4253), 
        .ZN(n4254) );
  OAI21_X1 U5191 ( .B1(n4287), .B2(EBX_REG_15__SCAN_IN), .A(n4254), .ZN(n5135)
         );
  OR2_X2 U5192 ( .A1(n5134), .A2(n5135), .ZN(n5244) );
  MUX2_X1 U5193 ( .A(n4291), .B(n4209), .S(EBX_REG_16__SCAN_IN), .Z(n4256) );
  NAND2_X1 U5194 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n5330), .ZN(n4255) );
  AND3_X1 U5195 ( .A1(n4256), .A2(n4279), .A3(n4255), .ZN(n5243) );
  INV_X1 U5196 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6923) );
  NAND2_X1 U5197 ( .A1(n4274), .A2(n6923), .ZN(n4259) );
  NAND2_X1 U5198 ( .A1(n5323), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4257) );
  OAI211_X1 U5199 ( .C1(n5330), .C2(EBX_REG_17__SCAN_IN), .A(n4290), .B(n4257), 
        .ZN(n4258) );
  AND2_X1 U5200 ( .A1(n4259), .A2(n4258), .ZN(n6029) );
  MUX2_X1 U5201 ( .A(n4291), .B(n4290), .S(EBX_REG_19__SCAN_IN), .Z(n4262) );
  NAND2_X1 U5202 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n5330), .ZN(n4260) );
  AND2_X1 U5203 ( .A1(n4279), .A2(n4260), .ZN(n4261) );
  NAND2_X1 U5204 ( .A1(n4262), .A2(n4261), .ZN(n5452) );
  OR2_X1 U5205 ( .A1(n5331), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n4264)
         );
  INV_X1 U5206 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5448) );
  NAND2_X1 U5207 ( .A1(n5207), .A2(n5448), .ZN(n4263) );
  AND2_X1 U5208 ( .A1(n4264), .A2(n4263), .ZN(n5446) );
  OR2_X1 U5209 ( .A1(n5331), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4265)
         );
  INV_X1 U5210 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5280) );
  NAND2_X1 U5211 ( .A1(n5207), .A2(n5280), .ZN(n5262) );
  NAND2_X1 U5212 ( .A1(n4265), .A2(n5262), .ZN(n5261) );
  NAND2_X1 U5213 ( .A1(n5444), .A2(EBX_REG_20__SCAN_IN), .ZN(n4267) );
  NAND2_X1 U5214 ( .A1(n5261), .A2(n5323), .ZN(n4266) );
  OAI211_X1 U5215 ( .C1(n5446), .C2(n5261), .A(n4267), .B(n4266), .ZN(n4268)
         );
  MUX2_X1 U5216 ( .A(n4287), .B(n5323), .S(EBX_REG_21__SCAN_IN), .Z(n4269) );
  OAI21_X1 U5217 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5331), .A(n4269), 
        .ZN(n5435) );
  MUX2_X1 U5218 ( .A(n4291), .B(n4290), .S(EBX_REG_22__SCAN_IN), .Z(n4272) );
  NAND2_X1 U5219 ( .A1(n5330), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4270) );
  AND2_X1 U5220 ( .A1(n4279), .A2(n4270), .ZN(n4271) );
  NAND2_X1 U5221 ( .A1(n4272), .A2(n4271), .ZN(n5424) );
  INV_X1 U5222 ( .A(EBX_REG_23__SCAN_IN), .ZN(n4273) );
  NAND2_X1 U5223 ( .A1(n4274), .A2(n4273), .ZN(n4277) );
  NAND2_X1 U5224 ( .A1(n5323), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4275) );
  OAI211_X1 U5225 ( .C1(n5330), .C2(EBX_REG_23__SCAN_IN), .A(n4209), .B(n4275), 
        .ZN(n4276) );
  AND2_X1 U5226 ( .A1(n4277), .A2(n4276), .ZN(n5419) );
  MUX2_X1 U5227 ( .A(n4291), .B(n4290), .S(EBX_REG_24__SCAN_IN), .Z(n4280) );
  NAND2_X1 U5228 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n5330), .ZN(n4278) );
  AND3_X1 U5229 ( .A1(n4280), .A2(n4279), .A3(n4278), .ZN(n5412) );
  OR2_X2 U5230 ( .A1(n5421), .A2(n5412), .ZN(n5414) );
  MUX2_X1 U5231 ( .A(n4287), .B(n5323), .S(EBX_REG_25__SCAN_IN), .Z(n4281) );
  OAI21_X1 U5232 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5331), .A(n4281), 
        .ZN(n5403) );
  INV_X1 U5233 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5905) );
  NAND2_X1 U5234 ( .A1(n4282), .A2(n5905), .ZN(n4286) );
  NAND2_X1 U5235 ( .A1(n4290), .A2(n5512), .ZN(n4284) );
  NAND2_X1 U5236 ( .A1(n5207), .A2(n5905), .ZN(n4283) );
  NAND3_X1 U5237 ( .A1(n4284), .A2(n5323), .A3(n4283), .ZN(n4285) );
  AND2_X1 U5238 ( .A1(n4286), .A2(n4285), .ZN(n5395) );
  NOR2_X2 U5239 ( .A1(n5405), .A2(n5395), .ZN(n5396) );
  MUX2_X1 U5240 ( .A(n4287), .B(n5323), .S(EBX_REG_27__SCAN_IN), .Z(n4289) );
  OR2_X1 U5241 ( .A1(n5331), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4288)
         );
  AND2_X1 U5242 ( .A1(n4289), .A2(n4288), .ZN(n5387) );
  AND2_X2 U5243 ( .A1(n5396), .A2(n5387), .ZN(n5389) );
  MUX2_X1 U5244 ( .A(n4291), .B(n4290), .S(EBX_REG_28__SCAN_IN), .Z(n4293) );
  NAND2_X1 U5245 ( .A1(n5330), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4292) );
  NAND2_X1 U5246 ( .A1(n4293), .A2(n4292), .ZN(n5381) );
  AND2_X4 U5247 ( .A1(n5389), .A2(n5381), .ZN(n5383) );
  MUX2_X1 U5248 ( .A(n5323), .B(n5324), .S(n5383), .Z(n4295) );
  AND2_X1 U5249 ( .A1(n5330), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4294)
         );
  AOI21_X1 U5250 ( .B1(n5331), .B2(EBX_REG_30__SCAN_IN), .A(n4294), .ZN(n5329)
         );
  INV_X1 U5251 ( .A(n5375), .ZN(n4317) );
  NAND2_X1 U5252 ( .A1(n4296), .A2(n4585), .ZN(n5211) );
  OR2_X1 U5253 ( .A1(n5211), .A2(n3220), .ZN(n4300) );
  AND2_X1 U5254 ( .A1(n4297), .A2(n4300), .ZN(n4504) );
  NAND2_X1 U5255 ( .A1(n4504), .A2(n4298), .ZN(n4519) );
  INV_X1 U5256 ( .A(n4519), .ZN(n4364) );
  NOR2_X1 U5257 ( .A1(n6361), .A2(n4230), .ZN(n5125) );
  NAND3_X1 U5258 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .A3(n5125), .ZN(n4299) );
  INV_X1 U5259 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6372) );
  NAND2_X1 U5260 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6373) );
  NAND2_X1 U5261 ( .A1(n6372), .A2(n6373), .ZN(n6371) );
  NAND3_X1 U5262 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A3(n6371), .ZN(n4707) );
  NOR2_X1 U5263 ( .A1(n3502), .A2(n4707), .ZN(n4670) );
  NAND2_X1 U5264 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4670), .ZN(n4931)
         );
  NOR2_X1 U5265 ( .A1(n4299), .A2(n4931), .ZN(n4320) );
  NAND2_X1 U5266 ( .A1(n6377), .A2(n4320), .ZN(n6047) );
  NOR2_X1 U5267 ( .A1(n6372), .A2(n4201), .ZN(n4668) );
  INV_X1 U5268 ( .A(n4668), .ZN(n4666) );
  NAND2_X1 U5269 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4859) );
  NOR2_X1 U5270 ( .A1(n4666), .A2(n4859), .ZN(n4711) );
  NAND3_X1 U5271 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n4711), .ZN(n4934) );
  NOR2_X1 U5272 ( .A1(n4934), .A2(n4299), .ZN(n4321) );
  NAND3_X1 U5273 ( .A1(n4301), .A2(n4482), .A3(n4300), .ZN(n4303) );
  AOI22_X1 U5274 ( .A1(n4304), .A2(n4303), .B1(n4302), .B2(n5444), .ZN(n4305)
         );
  AND2_X1 U5275 ( .A1(n4306), .A2(n4305), .ZN(n4308) );
  AND2_X1 U5276 ( .A1(n4308), .A2(n4307), .ZN(n4517) );
  OAI21_X1 U5277 ( .B1(n5203), .B2(n4515), .A(n4517), .ZN(n4309) );
  NOR2_X1 U5278 ( .A1(n4170), .A2(n3271), .ZN(n5292) );
  NAND2_X1 U5279 ( .A1(n4318), .A2(n5292), .ZN(n5710) );
  INV_X1 U5280 ( .A(n5710), .ZN(n4409) );
  NOR2_X1 U5281 ( .A1(n6051), .A2(n4409), .ZN(n4322) );
  INV_X1 U5282 ( .A(n4322), .ZN(n4935) );
  INV_X1 U5283 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6391) );
  NAND2_X1 U5284 ( .A1(n5710), .A2(n6391), .ZN(n6388) );
  NAND2_X1 U5285 ( .A1(n4935), .A2(n6388), .ZN(n6378) );
  INV_X1 U5286 ( .A(n6378), .ZN(n4310) );
  NAND2_X1 U5287 ( .A1(n4321), .A2(n4310), .ZN(n5234) );
  NAND2_X1 U5288 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5711) );
  NOR2_X1 U5289 ( .A1(n4311), .A2(n5711), .ZN(n6046) );
  NAND2_X1 U5290 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n6046), .ZN(n5699) );
  NAND2_X1 U5291 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5704) );
  NOR2_X1 U5292 ( .A1(n5699), .A2(n5704), .ZN(n4325) );
  NAND2_X1 U5293 ( .A1(n6348), .A2(n4325), .ZN(n6022) );
  INV_X1 U5294 ( .A(n6022), .ZN(n6036) );
  NAND3_X1 U5295 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n6036), .ZN(n5692) );
  INV_X1 U5296 ( .A(n4312), .ZN(n4313) );
  INV_X1 U5297 ( .A(n6014), .ZN(n4314) );
  NAND2_X1 U5298 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4331) );
  NOR2_X1 U5299 ( .A1(n4314), .A2(n4331), .ZN(n5634) );
  NAND2_X1 U5300 ( .A1(n5634), .A2(n5622), .ZN(n5617) );
  NOR3_X1 U5301 ( .A1(n5617), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n3575), 
        .ZN(n4315) );
  AOI211_X1 U5302 ( .C1(n6375), .C2(n4317), .A(n4316), .B(n4315), .ZN(n4335)
         );
  INV_X1 U5303 ( .A(n6392), .ZN(n4412) );
  NAND2_X1 U5304 ( .A1(n4412), .A2(n5710), .ZN(n6389) );
  INV_X2 U5305 ( .A(n6187), .ZN(n6395) );
  NOR2_X1 U5306 ( .A1(n4318), .A2(n6395), .ZN(n6390) );
  AOI21_X1 U5307 ( .B1(n6051), .B2(n6391), .A(n6390), .ZN(n4319) );
  INV_X1 U5308 ( .A(n4319), .ZN(n4930) );
  OAI22_X1 U5309 ( .A1(n4322), .A2(n4321), .B1(n4320), .B2(n5235), .ZN(n4323)
         );
  NOR2_X1 U5310 ( .A1(n4930), .A2(n4323), .ZN(n6352) );
  NOR2_X1 U5311 ( .A1(n6389), .A2(n4930), .ZN(n4324) );
  AOI21_X1 U5312 ( .B1(n6352), .B2(n4325), .A(n4324), .ZN(n6037) );
  NAND4_X1 U5313 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A3(INSTADDRPOINTER_REG_19__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5646) );
  AND2_X1 U5314 ( .A1(n6389), .A2(n5646), .ZN(n4326) );
  OR2_X1 U5315 ( .A1(n6037), .A2(n4326), .ZN(n5676) );
  INV_X1 U5316 ( .A(n5647), .ZN(n5664) );
  AND2_X1 U5317 ( .A1(n6389), .A2(n5664), .ZN(n4327) );
  NOR2_X1 U5318 ( .A1(n5676), .A2(n4327), .ZN(n5658) );
  NAND2_X1 U5319 ( .A1(n6378), .A2(n5235), .ZN(n4667) );
  INV_X1 U5320 ( .A(n4328), .ZN(n4329) );
  NAND2_X1 U5321 ( .A1(n4667), .A2(n4329), .ZN(n4330) );
  INV_X1 U5322 ( .A(n4331), .ZN(n5628) );
  INV_X1 U5323 ( .A(n6389), .ZN(n5680) );
  AOI21_X1 U5324 ( .B1(n5622), .B2(n5628), .A(n5680), .ZN(n4332) );
  NOR2_X1 U5325 ( .A1(n5642), .A2(n4332), .ZN(n5612) );
  NAND2_X1 U5326 ( .A1(n5612), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4333) );
  OAI211_X1 U5327 ( .C1(n6389), .C2(n5642), .A(n4333), .B(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4334) );
  AND2_X1 U5328 ( .A1(n4335), .A2(n4334), .ZN(n4336) );
  NAND2_X1 U5329 ( .A1(n4337), .A2(n4336), .ZN(U2988) );
  NOR3_X1 U5330 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .A3(INSTADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n4339) );
  NAND3_X1 U5331 ( .A1(n3556), .A2(n5623), .A3(n4339), .ZN(n4340) );
  OR2_X1 U5332 ( .A1(n4338), .A2(n4340), .ZN(n4341) );
  XNOR2_X1 U5333 ( .A(n4342), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5603)
         );
  AOI22_X1 U5334 ( .A1(n4344), .A2(EAX_REG_31__SCAN_IN), .B1(n4343), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4345) );
  XNOR2_X2 U5335 ( .A(n4346), .B(n4345), .ZN(n5319) );
  NOR2_X2 U5336 ( .A1(n5319), .A2(n6344), .ZN(n4347) );
  INV_X1 U5337 ( .A(n4347), .ZN(n4352) );
  INV_X1 U5338 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n6818) );
  XNOR2_X1 U5339 ( .A(n4349), .B(n6818), .ZN(n5213) );
  NAND2_X1 U5340 ( .A1(n6395), .A2(REIP_REG_31__SCAN_IN), .ZN(n5606) );
  OAI21_X1 U5341 ( .B1(n5591), .B2(n6818), .A(n5606), .ZN(n4350) );
  NAND3_X1 U5342 ( .A1(n4353), .A2(n4352), .A3(n4351), .ZN(U2955) );
  OR2_X1 U5343 ( .A1(n4363), .A2(n4170), .ZN(n4358) );
  INV_X1 U5344 ( .A(n4358), .ZN(n4354) );
  NAND2_X1 U5345 ( .A1(n4354), .A2(n6583), .ZN(n4370) );
  INV_X1 U5346 ( .A(n4370), .ZN(n4356) );
  INV_X1 U5347 ( .A(MEMORYFETCH_REG_SCAN_IN), .ZN(n4355) );
  OR2_X1 U5348 ( .A1(n6477), .A2(STATE2_REG_1__SCAN_IN), .ZN(n6068) );
  OAI211_X1 U5349 ( .C1(n4356), .C2(n4355), .A(n4375), .B(n6068), .ZN(U2788)
         );
  NAND2_X1 U5350 ( .A1(n4358), .A2(n4357), .ZN(n4359) );
  OAI21_X1 U5351 ( .B1(n4507), .B2(n3129), .A(n4359), .ZN(n6066) );
  INV_X1 U5352 ( .A(n3129), .ZN(n5198) );
  NAND3_X1 U5353 ( .A1(n5198), .A2(n6601), .A3(n5330), .ZN(n4360) );
  AND2_X1 U5354 ( .A1(n4360), .A2(n6673), .ZN(n6675) );
  OR2_X1 U5355 ( .A1(n6066), .A2(n6675), .ZN(n6541) );
  AND2_X1 U5356 ( .A1(n6541), .A2(n6583), .ZN(n6075) );
  INV_X1 U5357 ( .A(MORE_REG_SCAN_IN), .ZN(n4369) );
  OR2_X1 U5358 ( .A1(n6537), .A2(n4361), .ZN(n4362) );
  NOR2_X1 U5359 ( .A1(n4362), .A2(n4470), .ZN(n4367) );
  NAND2_X1 U5360 ( .A1(n4363), .A2(n3130), .ZN(n4366) );
  NAND2_X1 U5361 ( .A1(n4507), .A2(n4364), .ZN(n4365) );
  OAI211_X1 U5362 ( .C1(n4507), .C2(n4367), .A(n4366), .B(n4365), .ZN(n6538)
         );
  NAND2_X1 U5363 ( .A1(n6075), .A2(n6538), .ZN(n4368) );
  OAI21_X1 U5364 ( .B1(n6075), .B2(n4369), .A(n4368), .ZN(U3471) );
  INV_X1 U5365 ( .A(n6068), .ZN(n4371) );
  OAI21_X1 U5366 ( .B1(n4371), .B2(READREQUEST_REG_SCAN_IN), .A(n5212), .ZN(
        n4373) );
  OAI21_X1 U5367 ( .B1(n3129), .B2(n5207), .A(n6671), .ZN(n4372) );
  NAND2_X1 U5368 ( .A1(n4373), .A2(n4372), .ZN(U3474) );
  INV_X1 U5369 ( .A(n4375), .ZN(n4374) );
  NAND2_X1 U5370 ( .A1(n4374), .A2(n3271), .ZN(n4634) );
  AOI21_X1 U5371 ( .B1(n6676), .B2(READY_N), .A(n4375), .ZN(n4458) );
  INV_X2 U5372 ( .A(n4458), .ZN(n4454) );
  NAND2_X1 U5373 ( .A1(n4454), .A2(UWORD_REG_7__SCAN_IN), .ZN(n4377) );
  NOR2_X1 U5374 ( .A1(n4502), .A2(READY_N), .ZN(n4376) );
  NAND2_X1 U5375 ( .A1(n4632), .A2(n4376), .ZN(n4476) );
  NAND2_X1 U5376 ( .A1(n4448), .A2(DATAI_7_), .ZN(n4428) );
  OAI211_X1 U5377 ( .C1(n4634), .C2(n6791), .A(n4377), .B(n4428), .ZN(U2931)
         );
  NAND2_X1 U5378 ( .A1(n4454), .A2(UWORD_REG_3__SCAN_IN), .ZN(n4378) );
  NAND2_X1 U5379 ( .A1(n4448), .A2(DATAI_3_), .ZN(n4420) );
  OAI211_X1 U5380 ( .C1(n4634), .C2(n5071), .A(n4378), .B(n4420), .ZN(U2927)
         );
  NAND2_X1 U5381 ( .A1(n4454), .A2(UWORD_REG_9__SCAN_IN), .ZN(n4379) );
  NAND2_X1 U5382 ( .A1(n4448), .A2(DATAI_9_), .ZN(n4450) );
  OAI211_X1 U5383 ( .C1(n4634), .C2(n6829), .A(n4379), .B(n4450), .ZN(U2933)
         );
  OAI21_X1 U5384 ( .B1(n5331), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4380), 
        .ZN(n5209) );
  INV_X1 U5385 ( .A(n4574), .ZN(n5320) );
  NAND3_X1 U5386 ( .A1(n4382), .A2(n4381), .A3(n5320), .ZN(n4384) );
  OR2_X1 U5387 ( .A1(n4384), .A2(n4383), .ZN(n4474) );
  OAI22_X1 U5388 ( .A1(n4507), .A2(n4519), .B1(n5330), .B2(n4474), .ZN(n4385)
         );
  AND2_X2 U5389 ( .A1(n4385), .A2(n6583), .ZN(n6284) );
  OR2_X1 U5390 ( .A1(n4387), .A2(n4386), .ZN(n4388) );
  NAND2_X1 U5391 ( .A1(n4389), .A2(n4388), .ZN(n6345) );
  NAND2_X2 U5392 ( .A1(n6284), .A2(n4574), .ZN(n5456) );
  OAI222_X1 U5393 ( .A1(n5209), .A2(n6274), .B1(n6903), .B2(n6284), .C1(n6345), 
        .C2(n5456), .ZN(U2859) );
  CLKBUF_X1 U5394 ( .A(n4390), .Z(n4493) );
  CLKBUF_X1 U5395 ( .A(n4391), .Z(n4401) );
  OR2_X1 U5396 ( .A1(n4401), .A2(n4392), .ZN(n4393) );
  AND2_X1 U5397 ( .A1(n4493), .A2(n4393), .ZN(n6233) );
  INV_X1 U5398 ( .A(n6233), .ZN(n4484) );
  INV_X1 U5399 ( .A(n4394), .ZN(n4395) );
  XNOR2_X1 U5400 ( .A(n4396), .B(n4395), .ZN(n6234) );
  INV_X1 U5401 ( .A(n6284), .ZN(n5422) );
  AOI22_X1 U5402 ( .A1(n6279), .A2(n6234), .B1(EBX_REG_3__SCAN_IN), .B2(n5422), 
        .ZN(n4397) );
  OAI21_X1 U5403 ( .B1(n4484), .B2(n5456), .A(n4397), .ZN(U2856) );
  NOR2_X1 U5404 ( .A1(n4399), .A2(n4398), .ZN(n4400) );
  NOR2_X1 U5405 ( .A1(n4401), .A2(n4400), .ZN(n6330) );
  INV_X1 U5406 ( .A(n6330), .ZN(n4921) );
  XOR2_X1 U5407 ( .A(n4403), .B(n4402), .Z(n6374) );
  AOI22_X1 U5408 ( .A1(n6279), .A2(n6374), .B1(EBX_REG_2__SCAN_IN), .B2(n5422), 
        .ZN(n4404) );
  OAI21_X1 U5409 ( .B1(n4921), .B2(n5456), .A(n4404), .ZN(U2857) );
  INV_X1 U5410 ( .A(n4405), .ZN(n4407) );
  AOI21_X1 U5411 ( .B1(n4407), .B2(n6391), .A(n4406), .ZN(n6338) );
  NAND2_X1 U5412 ( .A1(n6395), .A2(REIP_REG_0__SCAN_IN), .ZN(n6336) );
  OAI21_X1 U5413 ( .B1(n6394), .B2(n5209), .A(n6336), .ZN(n4408) );
  AOI21_X1 U5414 ( .B1(n4195), .B2(n6338), .A(n4408), .ZN(n4411) );
  OAI21_X1 U5415 ( .B1(n6390), .B2(n4409), .A(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4410) );
  OAI211_X1 U5416 ( .C1(n4412), .C2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n4411), 
        .B(n4410), .ZN(U3018) );
  NAND2_X1 U5417 ( .A1(n4454), .A2(UWORD_REG_5__SCAN_IN), .ZN(n4413) );
  NAND2_X1 U5418 ( .A1(n4448), .A2(DATAI_5_), .ZN(n4417) );
  OAI211_X1 U5419 ( .C1(n4457), .C2(n6946), .A(n4413), .B(n4417), .ZN(U2929)
         );
  NAND2_X1 U5420 ( .A1(n4454), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4414) );
  NAND2_X1 U5421 ( .A1(n4448), .A2(DATAI_13_), .ZN(n4442) );
  OAI211_X1 U5422 ( .C1(n4457), .C2(n6305), .A(n4414), .B(n4442), .ZN(U2952)
         );
  INV_X1 U5423 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6860) );
  NAND2_X1 U5424 ( .A1(n4454), .A2(LWORD_REG_11__SCAN_IN), .ZN(n4415) );
  NAND2_X1 U5425 ( .A1(n4448), .A2(DATAI_11_), .ZN(n4446) );
  OAI211_X1 U5426 ( .C1(n6860), .C2(n4457), .A(n4415), .B(n4446), .ZN(U2950)
         );
  NAND2_X1 U5427 ( .A1(n4454), .A2(LWORD_REG_12__SCAN_IN), .ZN(n4416) );
  NAND2_X1 U5428 ( .A1(n4448), .A2(DATAI_12_), .ZN(n4444) );
  OAI211_X1 U5429 ( .C1(n5038), .C2(n4457), .A(n4416), .B(n4444), .ZN(U2951)
         );
  NAND2_X1 U5430 ( .A1(n4454), .A2(LWORD_REG_5__SCAN_IN), .ZN(n4418) );
  OAI211_X1 U5431 ( .C1(n3787), .C2(n4457), .A(n4418), .B(n4417), .ZN(U2944)
         );
  INV_X1 U5432 ( .A(EAX_REG_30__SCAN_IN), .ZN(n5080) );
  NAND2_X1 U5433 ( .A1(n4454), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4419) );
  NAND2_X1 U5434 ( .A1(n4448), .A2(DATAI_14_), .ZN(n4424) );
  OAI211_X1 U5435 ( .C1(n5080), .C2(n4457), .A(n4419), .B(n4424), .ZN(U2938)
         );
  NAND2_X1 U5436 ( .A1(n4454), .A2(LWORD_REG_3__SCAN_IN), .ZN(n4421) );
  OAI211_X1 U5437 ( .C1(n3667), .C2(n4457), .A(n4421), .B(n4420), .ZN(U2942)
         );
  INV_X1 U5438 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U5439 ( .A1(n4454), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4422) );
  NAND2_X1 U5440 ( .A1(n4448), .A2(DATAI_8_), .ZN(n4426) );
  OAI211_X1 U5441 ( .C1(n6313), .C2(n4457), .A(n4422), .B(n4426), .ZN(U2947)
         );
  NAND2_X1 U5442 ( .A1(n4454), .A2(LWORD_REG_1__SCAN_IN), .ZN(n4423) );
  NAND2_X1 U5443 ( .A1(n4448), .A2(DATAI_1_), .ZN(n4455) );
  OAI211_X1 U5444 ( .C1(n3643), .C2(n4457), .A(n4423), .B(n4455), .ZN(U2940)
         );
  NAND2_X1 U5445 ( .A1(n4454), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4425) );
  OAI211_X1 U5446 ( .C1(n5106), .C2(n4457), .A(n4425), .B(n4424), .ZN(U2953)
         );
  NAND2_X1 U5447 ( .A1(n4454), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4427) );
  OAI211_X1 U5448 ( .C1(n4010), .C2(n4457), .A(n4427), .B(n4426), .ZN(U2932)
         );
  NAND2_X1 U5449 ( .A1(n4454), .A2(LWORD_REG_7__SCAN_IN), .ZN(n4429) );
  OAI211_X1 U5450 ( .C1(n4922), .C2(n4457), .A(n4429), .B(n4428), .ZN(U2946)
         );
  NAND2_X1 U5451 ( .A1(n4454), .A2(LWORD_REG_6__SCAN_IN), .ZN(n4430) );
  NAND2_X1 U5452 ( .A1(n4448), .A2(DATAI_6_), .ZN(n4431) );
  OAI211_X1 U5453 ( .C1(n4853), .C2(n4457), .A(n4430), .B(n4431), .ZN(U2945)
         );
  INV_X1 U5454 ( .A(EAX_REG_22__SCAN_IN), .ZN(n5077) );
  NAND2_X1 U5455 ( .A1(n4454), .A2(UWORD_REG_6__SCAN_IN), .ZN(n4432) );
  OAI211_X1 U5456 ( .C1(n5077), .C2(n4457), .A(n4432), .B(n4431), .ZN(U2930)
         );
  INV_X1 U5457 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6939) );
  NAND2_X1 U5458 ( .A1(n4454), .A2(LWORD_REG_4__SCAN_IN), .ZN(n4433) );
  NAND2_X1 U5459 ( .A1(n4448), .A2(DATAI_4_), .ZN(n4434) );
  OAI211_X1 U5460 ( .C1(n6939), .C2(n4457), .A(n4433), .B(n4434), .ZN(U2943)
         );
  NAND2_X1 U5461 ( .A1(n4454), .A2(UWORD_REG_4__SCAN_IN), .ZN(n4435) );
  OAI211_X1 U5462 ( .C1(n3926), .C2(n4457), .A(n4435), .B(n4434), .ZN(U2928)
         );
  INV_X1 U5463 ( .A(EAX_REG_2__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U5464 ( .A1(n4454), .A2(LWORD_REG_2__SCAN_IN), .ZN(n4436) );
  NAND2_X1 U5465 ( .A1(n4448), .A2(DATAI_2_), .ZN(n4437) );
  OAI211_X1 U5466 ( .C1(n6321), .C2(n4457), .A(n4436), .B(n4437), .ZN(U2941)
         );
  INV_X1 U5467 ( .A(EAX_REG_18__SCAN_IN), .ZN(n5069) );
  NAND2_X1 U5468 ( .A1(n4454), .A2(UWORD_REG_2__SCAN_IN), .ZN(n4438) );
  OAI211_X1 U5469 ( .C1(n5069), .C2(n4457), .A(n4438), .B(n4437), .ZN(U2926)
         );
  NAND2_X1 U5470 ( .A1(n4454), .A2(LWORD_REG_0__SCAN_IN), .ZN(n4439) );
  NAND2_X1 U5471 ( .A1(n4448), .A2(DATAI_0_), .ZN(n4440) );
  OAI211_X1 U5472 ( .C1(n3650), .C2(n4457), .A(n4439), .B(n4440), .ZN(U2939)
         );
  INV_X1 U5473 ( .A(EAX_REG_16__SCAN_IN), .ZN(n6962) );
  NAND2_X1 U5474 ( .A1(n4454), .A2(UWORD_REG_0__SCAN_IN), .ZN(n4441) );
  OAI211_X1 U5475 ( .C1(n6962), .C2(n4457), .A(n4441), .B(n4440), .ZN(U2924)
         );
  INV_X1 U5476 ( .A(EAX_REG_29__SCAN_IN), .ZN(n6933) );
  NAND2_X1 U5477 ( .A1(n4454), .A2(UWORD_REG_13__SCAN_IN), .ZN(n4443) );
  OAI211_X1 U5478 ( .C1(n6933), .C2(n4457), .A(n4443), .B(n4442), .ZN(U2937)
         );
  NAND2_X1 U5479 ( .A1(n4454), .A2(UWORD_REG_12__SCAN_IN), .ZN(n4445) );
  OAI211_X1 U5480 ( .C1(n4096), .C2(n4457), .A(n4445), .B(n4444), .ZN(U2936)
         );
  NAND2_X1 U5481 ( .A1(n4454), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4447) );
  OAI211_X1 U5482 ( .C1(n4069), .C2(n4457), .A(n4447), .B(n4446), .ZN(U2935)
         );
  INV_X1 U5483 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6809) );
  NAND2_X1 U5484 ( .A1(n4454), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4449) );
  NAND2_X1 U5485 ( .A1(n4448), .A2(DATAI_10_), .ZN(n4452) );
  OAI211_X1 U5486 ( .C1(n6809), .C2(n4457), .A(n4449), .B(n4452), .ZN(U2934)
         );
  INV_X1 U5487 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6311) );
  NAND2_X1 U5488 ( .A1(n4454), .A2(LWORD_REG_9__SCAN_IN), .ZN(n4451) );
  OAI211_X1 U5489 ( .C1(n6311), .C2(n4457), .A(n4451), .B(n4450), .ZN(U2948)
         );
  INV_X1 U5490 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6309) );
  NAND2_X1 U5491 ( .A1(n4454), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4453) );
  OAI211_X1 U5492 ( .C1(n6309), .C2(n4457), .A(n4453), .B(n4452), .ZN(U2949)
         );
  NAND2_X1 U5493 ( .A1(n4454), .A2(UWORD_REG_1__SCAN_IN), .ZN(n4456) );
  OAI211_X1 U5494 ( .C1(n3873), .C2(n4457), .A(n4456), .B(n4455), .ZN(U2925)
         );
  INV_X1 U5495 ( .A(DATAI_15_), .ZN(n4460) );
  INV_X1 U5496 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4459) );
  INV_X1 U5497 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6302) );
  OAI222_X1 U5498 ( .A1(n4460), .A2(n4476), .B1(n4459), .B2(n4458), .C1(n4457), 
        .C2(n6302), .ZN(U2954) );
  INV_X1 U5499 ( .A(n5456), .ZN(n6280) );
  NOR2_X1 U5500 ( .A1(n4462), .A2(n4461), .ZN(n4463) );
  OR2_X1 U5501 ( .A1(n3659), .A2(n4463), .ZN(n5095) );
  INV_X1 U5502 ( .A(n5095), .ZN(n6263) );
  OR2_X1 U5503 ( .A1(n4464), .A2(n5207), .ZN(n4466) );
  AND2_X1 U5504 ( .A1(n4466), .A2(n4465), .ZN(n6393) );
  OAI22_X1 U5505 ( .A1(n6274), .A2(n6393), .B1(n4467), .B2(n6284), .ZN(n4468)
         );
  AOI21_X1 U5506 ( .B1(n6280), .B2(n6263), .A(n4468), .ZN(n4469) );
  INV_X1 U5507 ( .A(n4469), .ZN(U2858) );
  NAND2_X1 U5508 ( .A1(n4507), .A2(n4470), .ZN(n4473) );
  INV_X1 U5509 ( .A(n4514), .ZN(n6060) );
  NAND2_X1 U5510 ( .A1(n6060), .A2(n4471), .ZN(n4472) );
  NAND2_X1 U5511 ( .A1(n4473), .A2(n4472), .ZN(n4501) );
  NOR2_X1 U5512 ( .A1(n4474), .A2(n5198), .ZN(n4475) );
  OAI21_X1 U5513 ( .B1(n4501), .B2(n4475), .A(n6583), .ZN(n4477) );
  AND2_X1 U5514 ( .A1(n4478), .A2(n4574), .ZN(n4483) );
  INV_X1 U5515 ( .A(n4483), .ZN(n4480) );
  AND2_X1 U5516 ( .A1(n4480), .A2(n4479), .ZN(n4481) );
  NAND2_X2 U5517 ( .A1(n6299), .A2(n4481), .ZN(n6285) );
  INV_X1 U5518 ( .A(DATAI_3_), .ZN(n6750) );
  OAI222_X1 U5519 ( .A1(n4484), .A2(n6285), .B1(n5107), .B2(n6750), .C1(n6299), 
        .C2(n3667), .ZN(U2888) );
  INV_X1 U5520 ( .A(DATAI_0_), .ZN(n4590) );
  OAI222_X1 U5521 ( .A1(n6345), .A2(n6285), .B1(n5107), .B2(n4590), .C1(n6299), 
        .C2(n3650), .ZN(U2891) );
  OR2_X1 U5522 ( .A1(n4495), .A2(n4486), .ZN(n4850) );
  NAND2_X1 U5523 ( .A1(n4495), .A2(n4486), .ZN(n4487) );
  NAND2_X1 U5524 ( .A1(n4850), .A2(n4487), .ZN(n5040) );
  INV_X1 U5525 ( .A(DATAI_5_), .ZN(n4652) );
  OAI222_X1 U5526 ( .A1(n5040), .A2(n6285), .B1(n5107), .B2(n4652), .C1(n6299), 
        .C2(n3787), .ZN(U2886) );
  INV_X1 U5527 ( .A(n4489), .ZN(n4914) );
  AOI21_X1 U5528 ( .B1(n4490), .B2(n4499), .A(n4914), .ZN(n6211) );
  AOI22_X1 U5529 ( .A1(n6279), .A2(n6211), .B1(EBX_REG_5__SCAN_IN), .B2(n5422), 
        .ZN(n4491) );
  OAI21_X1 U5530 ( .B1(n5040), .B2(n5456), .A(n4491), .ZN(U2854) );
  NAND2_X1 U5531 ( .A1(n4493), .A2(n4492), .ZN(n4494) );
  AND2_X1 U5532 ( .A1(n4495), .A2(n4494), .ZN(n6223) );
  INV_X1 U5533 ( .A(n6223), .ZN(n4918) );
  OR2_X1 U5534 ( .A1(n4497), .A2(n4496), .ZN(n4498) );
  NAND2_X1 U5535 ( .A1(n4499), .A2(n4498), .ZN(n4858) );
  INV_X1 U5536 ( .A(n4858), .ZN(n6224) );
  AOI22_X1 U5537 ( .A1(n6279), .A2(n6224), .B1(EBX_REG_4__SCAN_IN), .B2(n5422), 
        .ZN(n4500) );
  OAI21_X1 U5538 ( .B1(n4918), .B2(n5456), .A(n4500), .ZN(U2855) );
  INV_X1 U5539 ( .A(n4501), .ZN(n4510) );
  OAI21_X1 U5540 ( .B1(n5292), .B2(n6572), .A(n4635), .ZN(n4503) );
  AOI21_X1 U5541 ( .B1(n4503), .B2(n4502), .A(READY_N), .ZN(n4506) );
  INV_X1 U5542 ( .A(n4504), .ZN(n4505) );
  AOI21_X1 U5543 ( .B1(n4507), .B2(n4506), .A(n4505), .ZN(n4509) );
  NAND3_X1 U5544 ( .A1(n4510), .A2(n4509), .A3(n4508), .ZN(n6548) );
  OR2_X1 U5545 ( .A1(n6548), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4525)
         );
  INV_X1 U5546 ( .A(n6572), .ZN(n4513) );
  AND4_X1 U5547 ( .A1(n4515), .A2(n4514), .A3(n4513), .A4(n4512), .ZN(n4516)
         );
  NAND2_X1 U5548 ( .A1(n4517), .A2(n4516), .ZN(n5294) );
  NAND2_X1 U5549 ( .A1(n6246), .A2(n5294), .ZN(n4523) );
  NAND2_X1 U5550 ( .A1(n4519), .A2(n4518), .ZN(n4533) );
  INV_X1 U5551 ( .A(n5309), .ZN(n5303) );
  NAND2_X1 U5552 ( .A1(n5303), .A2(n5317), .ZN(n4528) );
  OAI21_X1 U5553 ( .B1(n5317), .B2(n5303), .A(n4528), .ZN(n4521) );
  INV_X1 U5554 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n5290) );
  XNOR2_X1 U5555 ( .A(n5290), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4520)
         );
  AOI22_X1 U5556 ( .A1(n4533), .A2(n4521), .B1(n5292), .B2(n4520), .ZN(n4522)
         );
  AND2_X1 U5557 ( .A1(n4523), .A2(n4522), .ZN(n5307) );
  NAND2_X1 U5558 ( .A1(n6548), .A2(n5307), .ZN(n4524) );
  AND2_X1 U5559 ( .A1(n4525), .A2(n4524), .ZN(n6553) );
  OR2_X1 U5560 ( .A1(n6548), .A2(n5304), .ZN(n4537) );
  NAND2_X1 U5561 ( .A1(n4527), .A2(n5294), .ZN(n4535) );
  XNOR2_X1 U5562 ( .A(n4528), .B(n5304), .ZN(n4532) );
  AND2_X1 U5563 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4530) );
  INV_X1 U5564 ( .A(n4530), .ZN(n4529) );
  MUX2_X1 U5565 ( .A(n4530), .B(n4529), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4531) );
  AOI22_X1 U5566 ( .A1(n4533), .A2(n4532), .B1(n5292), .B2(n4531), .ZN(n4534)
         );
  NAND2_X1 U5567 ( .A1(n4535), .A2(n4534), .ZN(n5302) );
  NAND2_X1 U5568 ( .A1(n6548), .A2(n5302), .ZN(n4536) );
  NAND2_X1 U5569 ( .A1(n4537), .A2(n4536), .ZN(n6564) );
  NAND3_X1 U5570 ( .A1(n6553), .A2(n5295), .A3(n6564), .ZN(n4541) );
  INV_X1 U5571 ( .A(FLUSH_REG_SCAN_IN), .ZN(n6074) );
  AND2_X1 U5572 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6074), .ZN(n4539) );
  NAND2_X1 U5573 ( .A1(n4539), .A2(n4538), .ZN(n4540) );
  NAND2_X1 U5574 ( .A1(n4541), .A2(n4540), .ZN(n6543) );
  INV_X1 U5575 ( .A(n6543), .ZN(n4549) );
  MUX2_X1 U5576 ( .A(n6548), .B(FLUSH_REG_SCAN_IN), .S(STATE2_REG_1__SCAN_IN), 
        .Z(n4542) );
  INV_X1 U5577 ( .A(n4542), .ZN(n4543) );
  NAND2_X1 U5578 ( .A1(n4543), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4547) );
  INV_X1 U5579 ( .A(n4564), .ZN(n4618) );
  NOR2_X1 U5580 ( .A1(n4544), .A2(n4618), .ZN(n4545) );
  XNOR2_X1 U5581 ( .A(n4545), .B(n6063), .ZN(n6225) );
  NAND3_X1 U5582 ( .A1(n6225), .A2(n6060), .A3(n5295), .ZN(n4546) );
  AND2_X1 U5583 ( .A1(n4547), .A2(n4546), .ZN(n6566) );
  OAI21_X1 U5584 ( .B1(n4549), .B2(n4548), .A(n6566), .ZN(n4552) );
  NAND2_X1 U5585 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .ZN(n4637) );
  NOR2_X1 U5586 ( .A1(n6585), .A2(n4637), .ZN(n6591) );
  OAI21_X1 U5587 ( .B1(n4552), .B2(FLUSH_REG_SCAN_IN), .A(n6591), .ZN(n4551)
         );
  NOR2_X1 U5588 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6677) );
  INV_X1 U5589 ( .A(n6677), .ZN(n6578) );
  NAND2_X1 U5590 ( .A1(n4551), .A2(n4784), .ZN(n6404) );
  NOR2_X1 U5591 ( .A1(n4552), .A2(n4637), .ZN(n6576) );
  INV_X1 U5592 ( .A(n6474), .ZN(n4943) );
  AND2_X1 U5593 ( .A1(n6663), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5726) );
  OAI22_X1 U5594 ( .A1(n5735), .A2(n6477), .B1(n4943), .B2(n5726), .ZN(n4553)
         );
  OAI21_X1 U5595 ( .B1(n6576), .B2(n4553), .A(n6404), .ZN(n4554) );
  OAI21_X1 U5596 ( .B1(n6404), .B2(n6411), .A(n4554), .ZN(U3465) );
  NOR3_X1 U5597 ( .A1(n5725), .A2(n4557), .A3(n5722), .ZN(n5736) );
  NAND2_X1 U5598 ( .A1(n5736), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5783) );
  AND2_X1 U5599 ( .A1(n5783), .A2(n6473), .ZN(n4941) );
  NAND2_X1 U5600 ( .A1(n4601), .A2(n4557), .ZN(n4616) );
  NAND2_X1 U5601 ( .A1(n5722), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6472) );
  OR2_X1 U5602 ( .A1(n4616), .A2(n6472), .ZN(n4561) );
  AOI21_X1 U5603 ( .B1(n4941), .B2(n4561), .A(n6477), .ZN(n4559) );
  OR2_X1 U5604 ( .A1(n6477), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5832) );
  INV_X1 U5605 ( .A(n4527), .ZN(n5731) );
  OAI22_X1 U5606 ( .A1(n4717), .A2(n5832), .B1(n5731), .B2(n5726), .ZN(n4558)
         );
  OAI21_X1 U5607 ( .B1(n4559), .B2(n4558), .A(n6404), .ZN(n4560) );
  OAI21_X1 U5608 ( .B1(n6404), .B2(n6563), .A(n4560), .ZN(U3462) );
  INV_X1 U5609 ( .A(n6477), .ZN(n6471) );
  NAND2_X1 U5610 ( .A1(n4561), .A2(n6471), .ZN(n4569) );
  INV_X1 U5611 ( .A(n4563), .ZN(n6259) );
  NAND2_X1 U5612 ( .A1(n6246), .A2(n6259), .ZN(n6408) );
  OR2_X1 U5613 ( .A1(n6408), .A2(n4564), .ZN(n6415) );
  OAI21_X1 U5614 ( .B1(n6415), .B2(n4943), .A(n6449), .ZN(n4567) );
  INV_X1 U5615 ( .A(n6410), .ZN(n4565) );
  NAND2_X1 U5616 ( .A1(n6477), .A2(n4565), .ZN(n4566) );
  OAI211_X1 U5617 ( .C1(n4569), .C2(n4567), .A(n4873), .B(n4566), .ZN(n6463)
         );
  INV_X1 U5618 ( .A(n6463), .ZN(n4595) );
  INV_X1 U5619 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4578) );
  AND2_X1 U5620 ( .A1(DATAI_7_), .A2(n4720), .ZN(n6531) );
  INV_X1 U5621 ( .A(n4567), .ZN(n4568) );
  OR2_X1 U5622 ( .A1(n4569), .A2(n4568), .ZN(n4571) );
  NAND2_X1 U5623 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6410), .ZN(n4570) );
  NAND2_X1 U5624 ( .A1(n4571), .A2(n4570), .ZN(n6462) );
  NAND2_X1 U5625 ( .A1(n6329), .A2(DATAI_31_), .ZN(n6536) );
  INV_X1 U5626 ( .A(n4616), .ZN(n4572) );
  AND2_X1 U5627 ( .A1(n5722), .A2(n5735), .ZN(n5153) );
  NAND2_X1 U5628 ( .A1(n4572), .A2(n5733), .ZN(n6450) );
  NAND2_X1 U5629 ( .A1(n6329), .A2(DATAI_23_), .ZN(n6448) );
  OAI22_X1 U5630 ( .A1(n6536), .A2(n6466), .B1(n6450), .B2(n6448), .ZN(n4576)
         );
  NAND2_X1 U5631 ( .A1(n6585), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6661) );
  NAND2_X1 U5632 ( .A1(n4654), .A2(n4574), .ZN(n5780) );
  NOR2_X1 U5633 ( .A1(n5780), .A2(n6449), .ZN(n4575) );
  AOI211_X1 U5634 ( .C1(n6531), .C2(n6462), .A(n4576), .B(n4575), .ZN(n4577)
         );
  OAI21_X1 U5635 ( .B1(n4595), .B2(n4578), .A(n4577), .ZN(U3083) );
  INV_X1 U5636 ( .A(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4584) );
  INV_X1 U5637 ( .A(DATAI_4_), .ZN(n4917) );
  NAND2_X1 U5638 ( .A1(n4654), .A2(n4579), .ZN(n5862) );
  NOR2_X1 U5639 ( .A1(n5862), .A2(n6449), .ZN(n4582) );
  INV_X1 U5640 ( .A(DATAI_28_), .ZN(n4580) );
  NOR2_X1 U5641 ( .A1(n6344), .A2(n4580), .ZN(n6506) );
  INV_X1 U5642 ( .A(n6506), .ZN(n5807) );
  NAND2_X1 U5643 ( .A1(n6329), .A2(DATAI_20_), .ZN(n6511) );
  OAI22_X1 U5644 ( .A1(n5807), .A2(n6466), .B1(n6450), .B2(n6511), .ZN(n4581)
         );
  AOI211_X1 U5645 ( .C1(n6508), .C2(n6462), .A(n4582), .B(n4581), .ZN(n4583)
         );
  OAI21_X1 U5646 ( .B1(n4595), .B2(n4584), .A(n4583), .ZN(U3080) );
  INV_X1 U5647 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4589) );
  INV_X1 U5648 ( .A(DATAI_1_), .ZN(n4919) );
  NAND2_X1 U5649 ( .A1(n4654), .A2(n4585), .ZN(n5846) );
  NOR2_X1 U5650 ( .A1(n5846), .A2(n6449), .ZN(n4587) );
  INV_X1 U5651 ( .A(DATAI_25_), .ZN(n6959) );
  NOR2_X1 U5652 ( .A1(n6344), .A2(n6959), .ZN(n6488) );
  INV_X1 U5653 ( .A(n6488), .ZN(n5794) );
  NAND2_X1 U5654 ( .A1(n6329), .A2(DATAI_17_), .ZN(n6493) );
  OAI22_X1 U5655 ( .A1(n5794), .A2(n6466), .B1(n6450), .B2(n6493), .ZN(n4586)
         );
  AOI211_X1 U5656 ( .C1(n6490), .C2(n6462), .A(n4587), .B(n4586), .ZN(n4588)
         );
  OAI21_X1 U5657 ( .B1(n4595), .B2(n4589), .A(n4588), .ZN(U3077) );
  INV_X1 U5658 ( .A(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4594) );
  NAND2_X1 U5659 ( .A1(n4654), .A2(n5203), .ZN(n5840) );
  NOR2_X1 U5660 ( .A1(n5840), .A2(n6449), .ZN(n4592) );
  NAND2_X1 U5661 ( .A1(n6329), .A2(DATAI_24_), .ZN(n6487) );
  NAND2_X1 U5662 ( .A1(n6329), .A2(DATAI_16_), .ZN(n6424) );
  OAI22_X1 U5663 ( .A1(n6487), .A2(n6466), .B1(n6450), .B2(n6424), .ZN(n4591)
         );
  AOI211_X1 U5664 ( .C1(n6484), .C2(n6462), .A(n4592), .B(n4591), .ZN(n4593)
         );
  OAI21_X1 U5665 ( .B1(n4595), .B2(n4594), .A(n4593), .ZN(U3076) );
  NAND3_X1 U5666 ( .A1(n6563), .A2(n6557), .A3(n6948), .ZN(n4758) );
  NOR2_X1 U5667 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4758), .ZN(n4695)
         );
  INV_X1 U5668 ( .A(n4695), .ZN(n4615) );
  AND2_X1 U5669 ( .A1(n4607), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6406) );
  INV_X1 U5670 ( .A(n4783), .ZN(n4596) );
  OAI21_X1 U5671 ( .B1(n3139), .B2(n4606), .A(n4720), .ZN(n4619) );
  AOI211_X1 U5672 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4615), .A(n6406), .B(
        n4619), .ZN(n4604) );
  NAND2_X1 U5673 ( .A1(n4717), .A2(n4597), .ZN(n4598) );
  AND2_X1 U5674 ( .A1(n4599), .A2(n5722), .ZN(n4600) );
  OAI21_X1 U5675 ( .B1(n4777), .B2(n5878), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4602) );
  NOR2_X1 U5676 ( .A1(n6246), .A2(n6259), .ZN(n4821) );
  NAND2_X1 U5677 ( .A1(n5731), .A2(n4821), .ZN(n4605) );
  NAND3_X1 U5678 ( .A1(n4602), .A2(n6471), .A3(n4605), .ZN(n4603) );
  NAND2_X1 U5679 ( .A1(n4604), .A2(n4603), .ZN(n4691) );
  NAND2_X1 U5680 ( .A1(n4691), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4610) );
  INV_X1 U5681 ( .A(n6536), .ZN(n6444) );
  INV_X1 U5682 ( .A(n4777), .ZN(n4693) );
  INV_X1 U5683 ( .A(n4605), .ZN(n4753) );
  NOR2_X1 U5684 ( .A1(n4607), .A2(n4606), .ZN(n5156) );
  AOI22_X1 U5685 ( .A1(n4753), .A2(n6471), .B1(n5156), .B2(n3139), .ZN(n4698)
         );
  OAI22_X1 U5686 ( .A1(n4693), .A2(n6448), .B1(n4698), .B2(n5182), .ZN(n4608)
         );
  AOI21_X1 U5687 ( .B1(n6444), .B2(n5878), .A(n4608), .ZN(n4609) );
  OAI211_X1 U5688 ( .C1(n4615), .C2(n5780), .A(n4610), .B(n4609), .ZN(U3027)
         );
  NAND2_X1 U5689 ( .A1(n4654), .A2(n4611), .ZN(n5773) );
  NAND2_X1 U5690 ( .A1(n4691), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4614) );
  NAND2_X1 U5691 ( .A1(n6329), .A2(DATAI_30_), .ZN(n6467) );
  INV_X1 U5692 ( .A(n6467), .ZN(n6519) );
  NAND2_X1 U5693 ( .A1(n6329), .A2(DATAI_22_), .ZN(n6525) );
  AND2_X1 U5694 ( .A1(DATAI_6_), .A2(n4720), .ZN(n6521) );
  OAI22_X1 U5695 ( .A1(n4693), .A2(n6525), .B1(n4698), .B2(n5178), .ZN(n4612)
         );
  AOI21_X1 U5696 ( .B1(n6519), .B2(n5878), .A(n4612), .ZN(n4613) );
  OAI211_X1 U5697 ( .C1(n4615), .C2(n5773), .A(n4614), .B(n4613), .ZN(U3026)
         );
  NAND2_X1 U5698 ( .A1(n6948), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5788) );
  OR2_X1 U5699 ( .A1(n5788), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4874)
         );
  NOR2_X1 U5700 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4874), .ZN(n4701)
         );
  INV_X1 U5701 ( .A(n4701), .ZN(n4631) );
  OR2_X1 U5702 ( .A1(n4871), .A2(n6072), .ZN(n4617) );
  NAND2_X1 U5703 ( .A1(n4617), .A2(n6471), .ZN(n4877) );
  NAND3_X1 U5704 ( .A1(n5725), .A2(n5733), .A3(n4717), .ZN(n4975) );
  INV_X1 U5705 ( .A(n5832), .ZN(n6416) );
  AND2_X1 U5706 ( .A1(n6246), .A2(n4563), .ZN(n5782) );
  NAND2_X1 U5707 ( .A1(n5782), .A2(n4618), .ZN(n4866) );
  OAI21_X1 U5708 ( .B1(n4975), .B2(n6416), .A(n4866), .ZN(n4621) );
  AOI211_X1 U5709 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4631), .A(n5156), .B(
        n4619), .ZN(n4620) );
  OAI21_X1 U5710 ( .B1(n4877), .B2(n4621), .A(n4620), .ZN(n4699) );
  NAND2_X1 U5711 ( .A1(n4699), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4626) );
  INV_X1 U5712 ( .A(n6525), .ZN(n6460) );
  INV_X1 U5713 ( .A(n4898), .ZN(n4628) );
  OR2_X1 U5714 ( .A1(n4527), .A2(n6477), .ZN(n6409) );
  INV_X1 U5715 ( .A(n6409), .ZN(n4623) );
  AND2_X1 U5716 ( .A1(n3139), .A2(n6406), .ZN(n4622) );
  AOI21_X1 U5717 ( .B1(n4623), .B2(n5782), .A(n4622), .ZN(n4704) );
  OAI22_X1 U5718 ( .A1(n4975), .A2(n6467), .B1(n4704), .B2(n5178), .ZN(n4624)
         );
  AOI21_X1 U5719 ( .B1(n6460), .B2(n4628), .A(n4624), .ZN(n4625) );
  OAI211_X1 U5720 ( .C1(n4631), .C2(n5773), .A(n4626), .B(n4625), .ZN(U3058)
         );
  NAND2_X1 U5721 ( .A1(n4699), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4630) );
  INV_X1 U5722 ( .A(n6448), .ZN(n6527) );
  OAI22_X1 U5723 ( .A1(n4975), .A2(n6536), .B1(n4704), .B2(n5182), .ZN(n4627)
         );
  AOI21_X1 U5724 ( .B1(n6527), .B2(n4628), .A(n4627), .ZN(n4629) );
  OAI211_X1 U5725 ( .C1(n4631), .C2(n5780), .A(n4630), .B(n4629), .ZN(U3059)
         );
  NAND2_X1 U5726 ( .A1(n4632), .A2(n5292), .ZN(n4633) );
  NAND2_X1 U5727 ( .A1(n4634), .A2(n4633), .ZN(n4636) );
  NAND2_X1 U5728 ( .A1(n6300), .A2(n5203), .ZN(n5084) );
  NOR2_X1 U5729 ( .A1(n4637), .A2(STATE2_REG_0__SCAN_IN), .ZN(n5082) );
  AOI22_X1 U5730 ( .A1(n5082), .A2(UWORD_REG_12__SCAN_IN), .B1(n6316), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4638) );
  OAI21_X1 U5731 ( .B1(n4096), .B2(n5084), .A(n4638), .ZN(U2895) );
  AOI22_X1 U5732 ( .A1(n5082), .A2(UWORD_REG_13__SCAN_IN), .B1(n6316), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4639) );
  OAI21_X1 U5733 ( .B1(n6933), .B2(n5084), .A(n4639), .ZN(U2894) );
  AOI22_X1 U5734 ( .A1(n5082), .A2(UWORD_REG_10__SCAN_IN), .B1(n6316), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4640) );
  OAI21_X1 U5735 ( .B1(n6809), .B2(n5084), .A(n4640), .ZN(U2897) );
  AOI22_X1 U5736 ( .A1(n5082), .A2(UWORD_REG_8__SCAN_IN), .B1(n6316), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4641) );
  OAI21_X1 U5737 ( .B1(n4010), .B2(n5084), .A(n4641), .ZN(U2899) );
  NAND2_X1 U5738 ( .A1(n4699), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4645) );
  NAND2_X1 U5739 ( .A1(n4654), .A2(n4642), .ZN(n5856) );
  NAND2_X1 U5740 ( .A1(n6329), .A2(DATAI_19_), .ZN(n6434) );
  NAND2_X1 U5741 ( .A1(n6329), .A2(DATAI_27_), .ZN(n6505) );
  OAI22_X1 U5742 ( .A1(n4898), .A2(n6434), .B1(n4975), .B2(n6505), .ZN(n4643)
         );
  AOI21_X1 U5743 ( .B1(n6501), .B2(n4701), .A(n4643), .ZN(n4644) );
  OAI211_X1 U5744 ( .C1(n4704), .C2(n5759), .A(n4645), .B(n4644), .ZN(U3055)
         );
  NAND2_X1 U5745 ( .A1(n4691), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4648) );
  INV_X1 U5746 ( .A(n5878), .ZN(n4692) );
  OAI22_X1 U5747 ( .A1(n4693), .A2(n6434), .B1(n4692), .B2(n6505), .ZN(n4646)
         );
  AOI21_X1 U5748 ( .B1(n6501), .B2(n4695), .A(n4646), .ZN(n4647) );
  OAI211_X1 U5749 ( .C1(n4698), .C2(n5759), .A(n4648), .B(n4647), .ZN(U3023)
         );
  INV_X1 U5750 ( .A(DATAI_2_), .ZN(n4920) );
  NAND2_X1 U5751 ( .A1(n4699), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4651) );
  NAND2_X1 U5752 ( .A1(n4654), .A2(n3220), .ZN(n5851) );
  NAND2_X1 U5753 ( .A1(n6329), .A2(DATAI_18_), .ZN(n6430) );
  NAND2_X1 U5754 ( .A1(n6329), .A2(DATAI_26_), .ZN(n6499) );
  OAI22_X1 U5755 ( .A1(n4898), .A2(n6430), .B1(n4975), .B2(n6499), .ZN(n4649)
         );
  AOI21_X1 U5756 ( .B1(n6495), .B2(n4701), .A(n4649), .ZN(n4650) );
  OAI211_X1 U5757 ( .C1(n4704), .C2(n5755), .A(n4651), .B(n4650), .ZN(U3054)
         );
  NAND2_X1 U5758 ( .A1(n4691), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4657) );
  NAND2_X1 U5759 ( .A1(n4654), .A2(n4653), .ZN(n5869) );
  NAND2_X1 U5760 ( .A1(n6329), .A2(DATAI_21_), .ZN(n6517) );
  NAND2_X1 U5761 ( .A1(n6329), .A2(DATAI_29_), .ZN(n6458) );
  OAI22_X1 U5762 ( .A1(n4693), .A2(n6517), .B1(n4692), .B2(n6458), .ZN(n4655)
         );
  AOI21_X1 U5763 ( .B1(n6513), .B2(n4695), .A(n4655), .ZN(n4656) );
  OAI211_X1 U5764 ( .C1(n4698), .C2(n5768), .A(n4657), .B(n4656), .ZN(U3025)
         );
  NAND2_X1 U5765 ( .A1(n4699), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4660) );
  OAI22_X1 U5766 ( .A1(n4898), .A2(n6517), .B1(n4975), .B2(n6458), .ZN(n4658)
         );
  AOI21_X1 U5767 ( .B1(n6513), .B2(n4701), .A(n4658), .ZN(n4659) );
  OAI211_X1 U5768 ( .C1(n4704), .C2(n5768), .A(n4660), .B(n4659), .ZN(U3057)
         );
  NAND2_X1 U5769 ( .A1(n4691), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4663) );
  OAI22_X1 U5770 ( .A1(n4693), .A2(n6430), .B1(n4692), .B2(n6499), .ZN(n4661)
         );
  AOI21_X1 U5771 ( .B1(n6495), .B2(n4695), .A(n4661), .ZN(n4662) );
  OAI211_X1 U5772 ( .C1(n4698), .C2(n5755), .A(n4663), .B(n4662), .ZN(U3022)
         );
  XNOR2_X1 U5773 ( .A(n4664), .B(n4665), .ZN(n5051) );
  AOI21_X1 U5774 ( .B1(n4935), .B2(n4666), .A(n4930), .ZN(n6379) );
  OAI21_X1 U5775 ( .B1(n5680), .B2(n4670), .A(n6379), .ZN(n4709) );
  OAI21_X1 U5776 ( .B1(n6377), .B2(n4668), .A(n4667), .ZN(n4926) );
  NOR2_X1 U5777 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4926), .ZN(n4669)
         );
  AOI22_X1 U5778 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4709), .B1(n4670), 
        .B2(n4669), .ZN(n4673) );
  XNOR2_X1 U5779 ( .A(n4489), .B(n4913), .ZN(n6201) );
  INV_X1 U5780 ( .A(REIP_REG_6__SCAN_IN), .ZN(n4671) );
  NOR2_X1 U5781 ( .A1(n6187), .A2(n4671), .ZN(n5046) );
  AOI21_X1 U5782 ( .B1(n6375), .B2(n6201), .A(n5046), .ZN(n4672) );
  OAI211_X1 U5783 ( .C1(n6399), .C2(n5051), .A(n4673), .B(n4672), .ZN(U3012)
         );
  XNOR2_X1 U5784 ( .A(n4675), .B(n4674), .ZN(n5067) );
  OAI21_X1 U5785 ( .B1(n5235), .B2(n6371), .A(n6379), .ZN(n4864) );
  INV_X1 U5786 ( .A(n6371), .ZN(n4676) );
  NOR2_X1 U5787 ( .A1(n4676), .A2(n4926), .ZN(n4860) );
  AOI22_X1 U5788 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4864), .B1(n4860), 
        .B2(n3455), .ZN(n4678) );
  INV_X1 U5789 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6615) );
  NOR2_X1 U5790 ( .A1(n6187), .A2(n6615), .ZN(n5063) );
  AOI21_X1 U5791 ( .B1(n6375), .B2(n6234), .A(n5063), .ZN(n4677) );
  OAI211_X1 U5792 ( .C1(n6399), .C2(n5067), .A(n4678), .B(n4677), .ZN(U3015)
         );
  NAND2_X1 U5793 ( .A1(n4699), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4681) );
  OAI22_X1 U5794 ( .A1(n4898), .A2(n6511), .B1(n4975), .B2(n5807), .ZN(n4679)
         );
  AOI21_X1 U5795 ( .B1(n6507), .B2(n4701), .A(n4679), .ZN(n4680) );
  OAI211_X1 U5796 ( .C1(n4704), .C2(n5763), .A(n4681), .B(n4680), .ZN(U3056)
         );
  NAND2_X1 U5797 ( .A1(n4691), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4684) );
  OAI22_X1 U5798 ( .A1(n4693), .A2(n6493), .B1(n4692), .B2(n5794), .ZN(n4682)
         );
  AOI21_X1 U5799 ( .B1(n6489), .B2(n4695), .A(n4682), .ZN(n4683) );
  OAI211_X1 U5800 ( .C1(n4698), .C2(n5751), .A(n4684), .B(n4683), .ZN(U3021)
         );
  NAND2_X1 U5801 ( .A1(n4691), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4687) );
  OAI22_X1 U5802 ( .A1(n4693), .A2(n6511), .B1(n4692), .B2(n5807), .ZN(n4685)
         );
  AOI21_X1 U5803 ( .B1(n6507), .B2(n4695), .A(n4685), .ZN(n4686) );
  OAI211_X1 U5804 ( .C1(n4698), .C2(n5763), .A(n4687), .B(n4686), .ZN(U3024)
         );
  NAND2_X1 U5805 ( .A1(n4699), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4690) );
  OAI22_X1 U5806 ( .A1(n4898), .A2(n6493), .B1(n4975), .B2(n5794), .ZN(n4688)
         );
  AOI21_X1 U5807 ( .B1(n6489), .B2(n4701), .A(n4688), .ZN(n4689) );
  OAI211_X1 U5808 ( .C1(n4704), .C2(n5751), .A(n4690), .B(n4689), .ZN(U3053)
         );
  NAND2_X1 U5809 ( .A1(n4691), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4697) );
  OAI22_X1 U5810 ( .A1(n4693), .A2(n6424), .B1(n4692), .B2(n6487), .ZN(n4694)
         );
  AOI21_X1 U5811 ( .B1(n6470), .B2(n4695), .A(n4694), .ZN(n4696) );
  OAI211_X1 U5812 ( .C1(n4698), .C2(n5747), .A(n4697), .B(n4696), .ZN(U3020)
         );
  NAND2_X1 U5813 ( .A1(n4699), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4703) );
  OAI22_X1 U5814 ( .A1(n4898), .A2(n6424), .B1(n4975), .B2(n6487), .ZN(n4700)
         );
  AOI21_X1 U5815 ( .B1(n6470), .B2(n4701), .A(n4700), .ZN(n4702) );
  OAI211_X1 U5816 ( .C1(n4704), .C2(n5747), .A(n4703), .B(n4702), .ZN(U3052)
         );
  XNOR2_X1 U5817 ( .A(n4706), .B(n4705), .ZN(n5045) );
  NOR2_X1 U5818 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n6378), .ZN(n4710)
         );
  OAI21_X1 U5819 ( .B1(n5235), .B2(n4707), .A(n3502), .ZN(n4708) );
  AOI22_X1 U5820 ( .A1(n4711), .A2(n4710), .B1(n4709), .B2(n4708), .ZN(n4713)
         );
  INV_X1 U5821 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6620) );
  NOR2_X1 U5822 ( .A1(n6187), .A2(n6620), .ZN(n5041) );
  AOI21_X1 U5823 ( .B1(n6375), .B2(n6211), .A(n5041), .ZN(n4712) );
  OAI211_X1 U5824 ( .C1(n6399), .C2(n5045), .A(n4713), .B(n4712), .ZN(U3013)
         );
  NOR2_X1 U5825 ( .A1(n6246), .A2(n4563), .ZN(n5155) );
  NAND2_X1 U5826 ( .A1(n5731), .A2(n5155), .ZN(n4944) );
  INV_X1 U5827 ( .A(n4944), .ZN(n4714) );
  NAND2_X1 U5828 ( .A1(n4714), .A2(n6471), .ZN(n4716) );
  NAND3_X1 U5829 ( .A1(n5156), .A2(n6405), .A3(n6563), .ZN(n4715) );
  AND2_X1 U5830 ( .A1(n4716), .A2(n4715), .ZN(n4751) );
  NAND3_X1 U5831 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6563), .A3(n6557), .ZN(n4951) );
  NOR2_X1 U5832 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4951), .ZN(n4748)
         );
  AND2_X1 U5833 ( .A1(n4717), .A2(n5153), .ZN(n4718) );
  AND2_X1 U5834 ( .A1(n4718), .A2(n5725), .ZN(n4722) );
  OAI21_X1 U5835 ( .B1(n4778), .B2(n4722), .A(n5832), .ZN(n4719) );
  AOI21_X1 U5836 ( .B1(n4719), .B2(n4944), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4721) );
  OAI21_X1 U5837 ( .B1(n6405), .B2(n6480), .A(n4720), .ZN(n5003) );
  NOR2_X1 U5838 ( .A1(n6406), .A2(n5003), .ZN(n5162) );
  OAI21_X1 U5839 ( .B1(n4748), .B2(n4721), .A(n5162), .ZN(n4745) );
  NAND2_X1 U5840 ( .A1(n4745), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4725) );
  INV_X1 U5841 ( .A(n4778), .ZN(n4746) );
  OAI22_X1 U5842 ( .A1(n4746), .A2(n5807), .B1(n6511), .B2(n4976), .ZN(n4723)
         );
  AOI21_X1 U5843 ( .B1(n6507), .B2(n4748), .A(n4723), .ZN(n4724) );
  OAI211_X1 U5844 ( .C1(n5763), .C2(n4751), .A(n4725), .B(n4724), .ZN(U3040)
         );
  NAND2_X1 U5845 ( .A1(n4745), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4728) );
  OAI22_X1 U5846 ( .A1(n4746), .A2(n6487), .B1(n6424), .B2(n4976), .ZN(n4726)
         );
  AOI21_X1 U5847 ( .B1(n6470), .B2(n4748), .A(n4726), .ZN(n4727) );
  OAI211_X1 U5848 ( .C1(n5747), .C2(n4751), .A(n4728), .B(n4727), .ZN(U3036)
         );
  NAND2_X1 U5849 ( .A1(n4745), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4731) );
  OAI22_X1 U5850 ( .A1(n4746), .A2(n6458), .B1(n6517), .B2(n4976), .ZN(n4729)
         );
  AOI21_X1 U5851 ( .B1(n6513), .B2(n4748), .A(n4729), .ZN(n4730) );
  OAI211_X1 U5852 ( .C1(n5768), .C2(n4751), .A(n4731), .B(n4730), .ZN(U3041)
         );
  NAND2_X1 U5853 ( .A1(n4745), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4734) );
  OAI22_X1 U5854 ( .A1(n4746), .A2(n6499), .B1(n6430), .B2(n4976), .ZN(n4732)
         );
  AOI21_X1 U5855 ( .B1(n6495), .B2(n4748), .A(n4732), .ZN(n4733) );
  OAI211_X1 U5856 ( .C1(n5755), .C2(n4751), .A(n4734), .B(n4733), .ZN(U3038)
         );
  NAND2_X1 U5857 ( .A1(n4745), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4737) );
  OAI22_X1 U5858 ( .A1(n4746), .A2(n6505), .B1(n6434), .B2(n4976), .ZN(n4735)
         );
  AOI21_X1 U5859 ( .B1(n6501), .B2(n4748), .A(n4735), .ZN(n4736) );
  OAI211_X1 U5860 ( .C1(n5759), .C2(n4751), .A(n4737), .B(n4736), .ZN(U3039)
         );
  INV_X1 U5861 ( .A(n4748), .ZN(n4744) );
  NAND2_X1 U5862 ( .A1(n4745), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4740) );
  OAI22_X1 U5863 ( .A1(n4976), .A2(n6525), .B1(n4751), .B2(n5178), .ZN(n4738)
         );
  AOI21_X1 U5864 ( .B1(n4778), .B2(n6519), .A(n4738), .ZN(n4739) );
  OAI211_X1 U5865 ( .C1(n4744), .C2(n5773), .A(n4740), .B(n4739), .ZN(U3042)
         );
  NAND2_X1 U5866 ( .A1(n4745), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4743) );
  OAI22_X1 U5867 ( .A1(n4976), .A2(n6448), .B1(n4751), .B2(n5182), .ZN(n4741)
         );
  AOI21_X1 U5868 ( .B1(n6444), .B2(n4778), .A(n4741), .ZN(n4742) );
  OAI211_X1 U5869 ( .C1(n4744), .C2(n5780), .A(n4743), .B(n4742), .ZN(U3043)
         );
  NAND2_X1 U5870 ( .A1(n4745), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4750) );
  OAI22_X1 U5871 ( .A1(n4746), .A2(n5794), .B1(n6493), .B2(n4976), .ZN(n4747)
         );
  AOI21_X1 U5872 ( .B1(n6489), .B2(n4748), .A(n4747), .ZN(n4749) );
  OAI211_X1 U5873 ( .C1(n5751), .C2(n4751), .A(n4750), .B(n4749), .ZN(U3037)
         );
  NOR2_X1 U5874 ( .A1(n6411), .A2(n4758), .ZN(n4752) );
  INV_X1 U5875 ( .A(n4752), .ZN(n4781) );
  AOI21_X1 U5876 ( .B1(n4753), .B2(n6474), .A(n4752), .ZN(n4760) );
  INV_X1 U5877 ( .A(n4754), .ZN(n4755) );
  AOI21_X1 U5878 ( .B1(n4755), .B2(STATEBS16_REG_SCAN_IN), .A(n6477), .ZN(
        n4757) );
  AOI22_X1 U5879 ( .A1(n4760), .A2(n4757), .B1(n6477), .B2(n4758), .ZN(n4756)
         );
  NAND2_X1 U5880 ( .A1(n4873), .A2(n4756), .ZN(n4776) );
  INV_X1 U5881 ( .A(n4757), .ZN(n4759) );
  OAI22_X1 U5882 ( .A1(n4760), .A2(n4759), .B1(n6480), .B2(n4758), .ZN(n4775)
         );
  AOI22_X1 U5883 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4776), .B1(n6521), 
        .B2(n4775), .ZN(n4762) );
  AOI22_X1 U5884 ( .A1(n6460), .A2(n4778), .B1(n4777), .B2(n6519), .ZN(n4761)
         );
  OAI211_X1 U5885 ( .C1(n5773), .C2(n4781), .A(n4762), .B(n4761), .ZN(U3034)
         );
  AOI22_X1 U5886 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4776), .B1(n6531), 
        .B2(n4775), .ZN(n4764) );
  AOI22_X1 U5887 ( .A1(n6527), .A2(n4778), .B1(n4777), .B2(n6444), .ZN(n4763)
         );
  OAI211_X1 U5888 ( .C1(n5780), .C2(n4781), .A(n4764), .B(n4763), .ZN(U3035)
         );
  AOI22_X1 U5889 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4776), .B1(n6502), 
        .B2(n4775), .ZN(n4766) );
  INV_X1 U5890 ( .A(n6434), .ZN(n6500) );
  INV_X1 U5891 ( .A(n6505), .ZN(n6431) );
  AOI22_X1 U5892 ( .A1(n6500), .A2(n4778), .B1(n4777), .B2(n6431), .ZN(n4765)
         );
  OAI211_X1 U5893 ( .C1(n5856), .C2(n4781), .A(n4766), .B(n4765), .ZN(U3031)
         );
  AOI22_X1 U5894 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4776), .B1(n6514), 
        .B2(n4775), .ZN(n4768) );
  INV_X1 U5895 ( .A(n6517), .ZN(n6455) );
  INV_X1 U5896 ( .A(n6458), .ZN(n6512) );
  AOI22_X1 U5897 ( .A1(n6455), .A2(n4778), .B1(n4777), .B2(n6512), .ZN(n4767)
         );
  OAI211_X1 U5898 ( .C1(n5869), .C2(n4781), .A(n4768), .B(n4767), .ZN(U3033)
         );
  AOI22_X1 U5899 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4776), .B1(n6496), 
        .B2(n4775), .ZN(n4770) );
  INV_X1 U5900 ( .A(n6430), .ZN(n6494) );
  INV_X1 U5901 ( .A(n6499), .ZN(n6427) );
  AOI22_X1 U5902 ( .A1(n6494), .A2(n4778), .B1(n4777), .B2(n6427), .ZN(n4769)
         );
  OAI211_X1 U5903 ( .C1(n5851), .C2(n4781), .A(n4770), .B(n4769), .ZN(U3030)
         );
  AOI22_X1 U5904 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4776), .B1(n6484), 
        .B2(n4775), .ZN(n4772) );
  INV_X1 U5905 ( .A(n6424), .ZN(n6469) );
  INV_X1 U5906 ( .A(n6487), .ZN(n6421) );
  AOI22_X1 U5907 ( .A1(n6469), .A2(n4778), .B1(n4777), .B2(n6421), .ZN(n4771)
         );
  OAI211_X1 U5908 ( .C1(n5840), .C2(n4781), .A(n4772), .B(n4771), .ZN(U3028)
         );
  AOI22_X1 U5909 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4776), .B1(n6490), 
        .B2(n4775), .ZN(n4774) );
  INV_X1 U5910 ( .A(n6493), .ZN(n5844) );
  AOI22_X1 U5911 ( .A1(n5844), .A2(n4778), .B1(n4777), .B2(n6488), .ZN(n4773)
         );
  OAI211_X1 U5912 ( .C1(n5846), .C2(n4781), .A(n4774), .B(n4773), .ZN(U3029)
         );
  AOI22_X1 U5913 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4776), .B1(n6508), 
        .B2(n4775), .ZN(n4780) );
  INV_X1 U5914 ( .A(n6511), .ZN(n5860) );
  AOI22_X1 U5915 ( .A1(n5860), .A2(n4778), .B1(n4777), .B2(n6506), .ZN(n4779)
         );
  OAI211_X1 U5916 ( .C1(n5862), .C2(n4781), .A(n4780), .B(n4779), .ZN(U3032)
         );
  NAND3_X1 U5917 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6557), .A3(n6948), .ZN(n4825) );
  NOR2_X1 U5918 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4825), .ZN(n4815)
         );
  INV_X1 U5919 ( .A(n4815), .ZN(n4797) );
  NOR2_X1 U5920 ( .A1(n6473), .A2(n5722), .ZN(n4828) );
  NAND3_X1 U5921 ( .A1(n4813), .A2(n6471), .A3(n6450), .ZN(n4782) );
  AND2_X1 U5922 ( .A1(n4821), .A2(n4527), .ZN(n4787) );
  AOI21_X1 U5923 ( .B1(n4782), .B2(n5832), .A(n4787), .ZN(n4786) );
  INV_X1 U5924 ( .A(n6406), .ZN(n4994) );
  OR2_X1 U5925 ( .A1(n6405), .A2(n4783), .ZN(n4788) );
  AOI21_X1 U5926 ( .B1(n4788), .B2(STATE2_REG_2__SCAN_IN), .A(n4784), .ZN(
        n5739) );
  OAI211_X1 U5927 ( .C1(n6663), .C2(n4815), .A(n4994), .B(n5739), .ZN(n4785)
         );
  NAND2_X1 U5928 ( .A1(n4816), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4793) );
  NAND2_X1 U5929 ( .A1(n4787), .A2(n6471), .ZN(n4790) );
  INV_X1 U5930 ( .A(n4788), .ZN(n5732) );
  NAND2_X1 U5931 ( .A1(n5156), .A2(n5732), .ZN(n4789) );
  AND2_X1 U5932 ( .A1(n4790), .A2(n4789), .ZN(n4819) );
  OAI22_X1 U5933 ( .A1(n6450), .A2(n6536), .B1(n4819), .B2(n5182), .ZN(n4791)
         );
  AOI21_X1 U5934 ( .B1(n4845), .B2(n6527), .A(n4791), .ZN(n4792) );
  OAI211_X1 U5935 ( .C1(n4797), .C2(n5780), .A(n4793), .B(n4792), .ZN(U3091)
         );
  NAND2_X1 U5936 ( .A1(n4816), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4796) );
  OAI22_X1 U5937 ( .A1(n6450), .A2(n6467), .B1(n4819), .B2(n5178), .ZN(n4794)
         );
  AOI21_X1 U5938 ( .B1(n4845), .B2(n6460), .A(n4794), .ZN(n4795) );
  OAI211_X1 U5939 ( .C1(n4797), .C2(n5773), .A(n4796), .B(n4795), .ZN(U3090)
         );
  OAI22_X1 U5940 ( .A1(n4813), .A2(n6493), .B1(n5794), .B2(n6450), .ZN(n4798)
         );
  AOI21_X1 U5941 ( .B1(n6489), .B2(n4815), .A(n4798), .ZN(n4800) );
  NAND2_X1 U5942 ( .A1(n4816), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4799) );
  OAI211_X1 U5943 ( .C1(n5751), .C2(n4819), .A(n4800), .B(n4799), .ZN(U3085)
         );
  OAI22_X1 U5944 ( .A1(n4813), .A2(n6434), .B1(n6505), .B2(n6450), .ZN(n4801)
         );
  AOI21_X1 U5945 ( .B1(n6501), .B2(n4815), .A(n4801), .ZN(n4803) );
  NAND2_X1 U5946 ( .A1(n4816), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4802) );
  OAI211_X1 U5947 ( .C1(n5759), .C2(n4819), .A(n4803), .B(n4802), .ZN(U3087)
         );
  OAI22_X1 U5948 ( .A1(n4813), .A2(n6424), .B1(n6487), .B2(n6450), .ZN(n4804)
         );
  AOI21_X1 U5949 ( .B1(n6470), .B2(n4815), .A(n4804), .ZN(n4806) );
  NAND2_X1 U5950 ( .A1(n4816), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4805) );
  OAI211_X1 U5951 ( .C1(n5747), .C2(n4819), .A(n4806), .B(n4805), .ZN(U3084)
         );
  OAI22_X1 U5952 ( .A1(n4813), .A2(n6430), .B1(n6499), .B2(n6450), .ZN(n4807)
         );
  AOI21_X1 U5953 ( .B1(n6495), .B2(n4815), .A(n4807), .ZN(n4809) );
  NAND2_X1 U5954 ( .A1(n4816), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4808) );
  OAI211_X1 U5955 ( .C1(n5755), .C2(n4819), .A(n4809), .B(n4808), .ZN(U3086)
         );
  OAI22_X1 U5956 ( .A1(n4813), .A2(n6511), .B1(n5807), .B2(n6450), .ZN(n4810)
         );
  AOI21_X1 U5957 ( .B1(n6507), .B2(n4815), .A(n4810), .ZN(n4812) );
  NAND2_X1 U5958 ( .A1(n4816), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4811) );
  OAI211_X1 U5959 ( .C1(n5763), .C2(n4819), .A(n4812), .B(n4811), .ZN(U3088)
         );
  OAI22_X1 U5960 ( .A1(n4813), .A2(n6517), .B1(n6458), .B2(n6450), .ZN(n4814)
         );
  AOI21_X1 U5961 ( .B1(n6513), .B2(n4815), .A(n4814), .ZN(n4818) );
  NAND2_X1 U5962 ( .A1(n4816), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4817) );
  OAI211_X1 U5963 ( .C1(n5768), .C2(n4819), .A(n4818), .B(n4817), .ZN(U3089)
         );
  NOR2_X1 U5964 ( .A1(n6411), .A2(n4825), .ZN(n4820) );
  INV_X1 U5965 ( .A(n4820), .ZN(n4848) );
  AND2_X1 U5966 ( .A1(n4527), .A2(n6474), .ZN(n5831) );
  AOI21_X1 U5967 ( .B1(n5831), .B2(n4821), .A(n4820), .ZN(n4827) );
  NOR2_X1 U5968 ( .A1(n5722), .A2(n6072), .ZN(n4822) );
  AOI21_X1 U5969 ( .B1(n5734), .B2(n4822), .A(n6477), .ZN(n4824) );
  AOI22_X1 U5970 ( .A1(n4827), .A2(n4824), .B1(n6477), .B2(n4825), .ZN(n4823)
         );
  NAND2_X1 U5971 ( .A1(n4873), .A2(n4823), .ZN(n4844) );
  INV_X1 U5972 ( .A(n4824), .ZN(n4826) );
  OAI22_X1 U5973 ( .A1(n4827), .A2(n4826), .B1(n4606), .B2(n4825), .ZN(n4843)
         );
  AOI22_X1 U5974 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4844), .B1(n6531), 
        .B2(n4843), .ZN(n4830) );
  AOI22_X1 U5975 ( .A1(n5152), .A2(n6527), .B1(n4845), .B2(n6444), .ZN(n4829)
         );
  OAI211_X1 U5976 ( .C1(n4848), .C2(n5780), .A(n4830), .B(n4829), .ZN(U3099)
         );
  AOI22_X1 U5977 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4844), .B1(n6521), 
        .B2(n4843), .ZN(n4832) );
  AOI22_X1 U5978 ( .A1(n5152), .A2(n6460), .B1(n4845), .B2(n6519), .ZN(n4831)
         );
  OAI211_X1 U5979 ( .C1(n4848), .C2(n5773), .A(n4832), .B(n4831), .ZN(U3098)
         );
  AOI22_X1 U5980 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4844), .B1(n6502), 
        .B2(n4843), .ZN(n4834) );
  AOI22_X1 U5981 ( .A1(n5152), .A2(n6500), .B1(n4845), .B2(n6431), .ZN(n4833)
         );
  OAI211_X1 U5982 ( .C1(n4848), .C2(n5856), .A(n4834), .B(n4833), .ZN(U3095)
         );
  AOI22_X1 U5983 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4844), .B1(n6514), 
        .B2(n4843), .ZN(n4836) );
  AOI22_X1 U5984 ( .A1(n5152), .A2(n6455), .B1(n4845), .B2(n6512), .ZN(n4835)
         );
  OAI211_X1 U5985 ( .C1(n4848), .C2(n5869), .A(n4836), .B(n4835), .ZN(U3097)
         );
  AOI22_X1 U5986 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4844), .B1(n6496), 
        .B2(n4843), .ZN(n4838) );
  AOI22_X1 U5987 ( .A1(n5152), .A2(n6494), .B1(n4845), .B2(n6427), .ZN(n4837)
         );
  OAI211_X1 U5988 ( .C1(n4848), .C2(n5851), .A(n4838), .B(n4837), .ZN(U3094)
         );
  AOI22_X1 U5989 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4844), .B1(n6508), 
        .B2(n4843), .ZN(n4840) );
  AOI22_X1 U5990 ( .A1(n5152), .A2(n5860), .B1(n4845), .B2(n6506), .ZN(n4839)
         );
  OAI211_X1 U5991 ( .C1(n4848), .C2(n5862), .A(n4840), .B(n4839), .ZN(U3096)
         );
  AOI22_X1 U5992 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4844), .B1(n6490), 
        .B2(n4843), .ZN(n4842) );
  AOI22_X1 U5993 ( .A1(n5152), .A2(n5844), .B1(n4845), .B2(n6488), .ZN(n4841)
         );
  OAI211_X1 U5994 ( .C1(n4848), .C2(n5846), .A(n4842), .B(n4841), .ZN(U3093)
         );
  AOI22_X1 U5995 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4844), .B1(n6484), 
        .B2(n4843), .ZN(n4847) );
  AOI22_X1 U5996 ( .A1(n6469), .A2(n5152), .B1(n4845), .B2(n6421), .ZN(n4846)
         );
  OAI211_X1 U5997 ( .C1(n4848), .C2(n5840), .A(n4847), .B(n4846), .ZN(U3092)
         );
  NOR2_X1 U5998 ( .A1(n4850), .A2(n4849), .ZN(n4910) );
  AND2_X1 U5999 ( .A1(n4850), .A2(n4849), .ZN(n4851) );
  NOR2_X1 U6000 ( .A1(n4910), .A2(n4851), .ZN(n6204) );
  INV_X1 U6001 ( .A(n6204), .ZN(n4855) );
  AOI22_X1 U6002 ( .A1(n6279), .A2(n6201), .B1(EBX_REG_6__SCAN_IN), .B2(n5422), 
        .ZN(n4852) );
  OAI21_X1 U6003 ( .B1(n4855), .B2(n5456), .A(n4852), .ZN(U2853) );
  INV_X1 U6004 ( .A(DATAI_6_), .ZN(n4854) );
  OAI222_X1 U6005 ( .A1(n4855), .A2(n6285), .B1(n4854), .B2(n5107), .C1(n4853), 
        .C2(n6299), .ZN(U2885) );
  XNOR2_X1 U6006 ( .A(n4857), .B(n4856), .ZN(n5056) );
  INV_X1 U6007 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6617) );
  OAI22_X1 U6008 ( .A1(n6394), .A2(n4858), .B1(n6617), .B2(n6187), .ZN(n4863)
         );
  OAI211_X1 U6009 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n4860), .B(n4859), .ZN(n4861) );
  INV_X1 U6010 ( .A(n4861), .ZN(n4862) );
  AOI211_X1 U6011 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n4864), .A(n4863), 
        .B(n4862), .ZN(n4865) );
  OAI21_X1 U6012 ( .B1(n6399), .B2(n5056), .A(n4865), .ZN(U3014) );
  INV_X1 U6013 ( .A(n4877), .ZN(n4870) );
  OR2_X1 U6014 ( .A1(n4866), .A2(n4943), .ZN(n4868) );
  NOR2_X1 U6015 ( .A1(n6411), .A2(n4874), .ZN(n4900) );
  INV_X1 U6016 ( .A(n4900), .ZN(n4867) );
  NAND2_X1 U6017 ( .A1(n4868), .A2(n4867), .ZN(n4876) );
  INV_X1 U6018 ( .A(n4874), .ZN(n4869) );
  AOI22_X1 U6019 ( .A1(n4870), .A2(n4876), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4869), .ZN(n4904) );
  INV_X1 U6020 ( .A(n5780), .ZN(n6529) );
  OAI22_X1 U6021 ( .A1(n6448), .A2(n6413), .B1(n4898), .B2(n6536), .ZN(n4872)
         );
  AOI21_X1 U6022 ( .B1(n6529), .B2(n4900), .A(n4872), .ZN(n4879) );
  AOI21_X1 U6023 ( .B1(n6477), .B2(n4874), .A(n6476), .ZN(n4875) );
  OAI21_X1 U6024 ( .B1(n4877), .B2(n4876), .A(n4875), .ZN(n4901) );
  NAND2_X1 U6025 ( .A1(n4901), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4878) );
  OAI211_X1 U6026 ( .C1(n4904), .C2(n5182), .A(n4879), .B(n4878), .ZN(U3067)
         );
  OAI22_X1 U6027 ( .A1(n6493), .A2(n6413), .B1(n4898), .B2(n5794), .ZN(n4880)
         );
  AOI21_X1 U6028 ( .B1(n6489), .B2(n4900), .A(n4880), .ZN(n4882) );
  NAND2_X1 U6029 ( .A1(n4901), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4881) );
  OAI211_X1 U6030 ( .C1(n5751), .C2(n4904), .A(n4882), .B(n4881), .ZN(U3061)
         );
  INV_X1 U6031 ( .A(n5773), .ZN(n6520) );
  OAI22_X1 U6032 ( .A1(n6525), .A2(n6413), .B1(n4898), .B2(n6467), .ZN(n4883)
         );
  AOI21_X1 U6033 ( .B1(n6520), .B2(n4900), .A(n4883), .ZN(n4885) );
  NAND2_X1 U6034 ( .A1(n4901), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4884) );
  OAI211_X1 U6035 ( .C1(n4904), .C2(n5178), .A(n4885), .B(n4884), .ZN(U3066)
         );
  OAI22_X1 U6036 ( .A1(n6511), .A2(n6413), .B1(n4898), .B2(n5807), .ZN(n4886)
         );
  AOI21_X1 U6037 ( .B1(n6507), .B2(n4900), .A(n4886), .ZN(n4888) );
  NAND2_X1 U6038 ( .A1(n4901), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4887) );
  OAI211_X1 U6039 ( .C1(n5763), .C2(n4904), .A(n4888), .B(n4887), .ZN(U3064)
         );
  OAI22_X1 U6040 ( .A1(n6517), .A2(n6413), .B1(n4898), .B2(n6458), .ZN(n4889)
         );
  AOI21_X1 U6041 ( .B1(n6513), .B2(n4900), .A(n4889), .ZN(n4891) );
  NAND2_X1 U6042 ( .A1(n4901), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4890) );
  OAI211_X1 U6043 ( .C1(n5768), .C2(n4904), .A(n4891), .B(n4890), .ZN(U3065)
         );
  OAI22_X1 U6044 ( .A1(n6434), .A2(n6413), .B1(n4898), .B2(n6505), .ZN(n4892)
         );
  AOI21_X1 U6045 ( .B1(n6501), .B2(n4900), .A(n4892), .ZN(n4894) );
  NAND2_X1 U6046 ( .A1(n4901), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4893) );
  OAI211_X1 U6047 ( .C1(n5759), .C2(n4904), .A(n4894), .B(n4893), .ZN(U3063)
         );
  OAI22_X1 U6048 ( .A1(n6430), .A2(n6413), .B1(n4898), .B2(n6499), .ZN(n4895)
         );
  AOI21_X1 U6049 ( .B1(n6495), .B2(n4900), .A(n4895), .ZN(n4897) );
  NAND2_X1 U6050 ( .A1(n4901), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4896) );
  OAI211_X1 U6051 ( .C1(n5755), .C2(n4904), .A(n4897), .B(n4896), .ZN(U3062)
         );
  OAI22_X1 U6052 ( .A1(n6424), .A2(n6413), .B1(n4898), .B2(n6487), .ZN(n4899)
         );
  AOI21_X1 U6053 ( .B1(n6470), .B2(n4900), .A(n4899), .ZN(n4903) );
  NAND2_X1 U6054 ( .A1(n4901), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4902) );
  OAI211_X1 U6055 ( .C1(n5747), .C2(n4904), .A(n4903), .B(n4902), .ZN(U3060)
         );
  NAND2_X1 U6056 ( .A1(n4906), .A2(n4905), .ZN(n4908) );
  NAND2_X1 U6057 ( .A1(n4908), .A2(n4907), .ZN(n4909) );
  NOR2_X1 U6058 ( .A1(n4910), .A2(n4909), .ZN(n4911) );
  OR2_X1 U6059 ( .A1(n4985), .A2(n4911), .ZN(n6194) );
  INV_X1 U6060 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4916) );
  AOI21_X1 U6061 ( .B1(n4914), .B2(n4913), .A(n4912), .ZN(n4915) );
  OR2_X1 U6062 ( .A1(n4915), .A2(n4928), .ZN(n6186) );
  OAI222_X1 U6063 ( .A1(n6194), .A2(n5456), .B1(n4916), .B2(n6284), .C1(n6274), 
        .C2(n6186), .ZN(U2852) );
  OAI222_X1 U6064 ( .A1(n4918), .A2(n6285), .B1(n5107), .B2(n4917), .C1(n6299), 
        .C2(n6939), .ZN(U2887) );
  OAI222_X1 U6065 ( .A1(n5095), .A2(n6285), .B1(n5107), .B2(n4919), .C1(n6299), 
        .C2(n3643), .ZN(U2890) );
  OAI222_X1 U6066 ( .A1(n4921), .A2(n6285), .B1(n5107), .B2(n4920), .C1(n6299), 
        .C2(n6321), .ZN(U2889) );
  INV_X1 U6067 ( .A(DATAI_7_), .ZN(n4923) );
  OAI222_X1 U6068 ( .A1(n6194), .A2(n6285), .B1(n4923), .B2(n5107), .C1(n4922), 
        .C2(n6299), .ZN(U2884) );
  XNOR2_X1 U6069 ( .A(n4924), .B(n4925), .ZN(n5151) );
  AOI21_X1 U6070 ( .B1(n6361), .B2(n4230), .A(n5125), .ZN(n4938) );
  NOR2_X1 U6071 ( .A1(n4931), .A2(n4926), .ZN(n6362) );
  NOR2_X1 U6072 ( .A1(n4928), .A2(n4927), .ZN(n4929) );
  OR2_X1 U6073 ( .A1(n4992), .A2(n4929), .ZN(n6175) );
  NAND2_X1 U6074 ( .A1(n6395), .A2(REIP_REG_8__SCAN_IN), .ZN(n5147) );
  OAI21_X1 U6075 ( .B1(n6394), .B2(n6175), .A(n5147), .ZN(n4937) );
  AOI21_X1 U6076 ( .B1(n4931), .B2(n6377), .A(n4930), .ZN(n4932) );
  INV_X1 U6077 ( .A(n4932), .ZN(n4933) );
  AOI21_X1 U6078 ( .B1(n4935), .B2(n4934), .A(n4933), .ZN(n6370) );
  NOR2_X1 U6079 ( .A1(n6370), .A2(n4230), .ZN(n4936) );
  AOI211_X1 U6080 ( .C1(n4938), .C2(n6362), .A(n4937), .B(n4936), .ZN(n4939)
         );
  OAI21_X1 U6081 ( .B1(n6399), .B2(n5151), .A(n4939), .ZN(U3010) );
  INV_X1 U6082 ( .A(n6472), .ZN(n4940) );
  NAND3_X1 U6083 ( .A1(n4941), .A2(n5725), .A3(n4940), .ZN(n4942) );
  NAND2_X1 U6084 ( .A1(n4942), .A2(n6471), .ZN(n4954) );
  INV_X1 U6085 ( .A(n4954), .ZN(n4948) );
  OR2_X1 U6086 ( .A1(n4944), .A2(n4943), .ZN(n4946) );
  INV_X1 U6087 ( .A(n6468), .ZN(n4945) );
  NAND2_X1 U6088 ( .A1(n4945), .A2(n6563), .ZN(n4949) );
  NAND2_X1 U6089 ( .A1(n4946), .A2(n4949), .ZN(n4953) );
  INV_X1 U6090 ( .A(n4951), .ZN(n4947) );
  AOI22_X1 U6091 ( .A1(n4948), .A2(n4953), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4947), .ZN(n4982) );
  INV_X1 U6092 ( .A(n4949), .ZN(n4978) );
  OAI22_X1 U6093 ( .A1(n4976), .A2(n6487), .B1(n6424), .B2(n4975), .ZN(n4950)
         );
  AOI21_X1 U6094 ( .B1(n6470), .B2(n4978), .A(n4950), .ZN(n4956) );
  AOI21_X1 U6095 ( .B1(n6477), .B2(n4951), .A(n6476), .ZN(n4952) );
  OAI21_X1 U6096 ( .B1(n4954), .B2(n4953), .A(n4952), .ZN(n4979) );
  NAND2_X1 U6097 ( .A1(n4979), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4955) );
  OAI211_X1 U6098 ( .C1(n5747), .C2(n4982), .A(n4956), .B(n4955), .ZN(U3044)
         );
  OAI22_X1 U6099 ( .A1(n4976), .A2(n5794), .B1(n6493), .B2(n4975), .ZN(n4957)
         );
  AOI21_X1 U6100 ( .B1(n6489), .B2(n4978), .A(n4957), .ZN(n4959) );
  NAND2_X1 U6101 ( .A1(n4979), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4958) );
  OAI211_X1 U6102 ( .C1(n5751), .C2(n4982), .A(n4959), .B(n4958), .ZN(U3045)
         );
  OAI22_X1 U6103 ( .A1(n4976), .A2(n6536), .B1(n6448), .B2(n4975), .ZN(n4960)
         );
  AOI21_X1 U6104 ( .B1(n6529), .B2(n4978), .A(n4960), .ZN(n4962) );
  NAND2_X1 U6105 ( .A1(n4979), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4961) );
  OAI211_X1 U6106 ( .C1(n4982), .C2(n5182), .A(n4962), .B(n4961), .ZN(U3051)
         );
  OAI22_X1 U6107 ( .A1(n4976), .A2(n6458), .B1(n6517), .B2(n4975), .ZN(n4963)
         );
  AOI21_X1 U6108 ( .B1(n6513), .B2(n4978), .A(n4963), .ZN(n4965) );
  NAND2_X1 U6109 ( .A1(n4979), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4964) );
  OAI211_X1 U6110 ( .C1(n5768), .C2(n4982), .A(n4965), .B(n4964), .ZN(U3049)
         );
  OAI22_X1 U6111 ( .A1(n4976), .A2(n5807), .B1(n6511), .B2(n4975), .ZN(n4966)
         );
  AOI21_X1 U6112 ( .B1(n6507), .B2(n4978), .A(n4966), .ZN(n4968) );
  NAND2_X1 U6113 ( .A1(n4979), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4967) );
  OAI211_X1 U6114 ( .C1(n5763), .C2(n4982), .A(n4968), .B(n4967), .ZN(U3048)
         );
  OAI22_X1 U6115 ( .A1(n4976), .A2(n6505), .B1(n6434), .B2(n4975), .ZN(n4969)
         );
  AOI21_X1 U6116 ( .B1(n6501), .B2(n4978), .A(n4969), .ZN(n4971) );
  NAND2_X1 U6117 ( .A1(n4979), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4970) );
  OAI211_X1 U6118 ( .C1(n5759), .C2(n4982), .A(n4971), .B(n4970), .ZN(U3047)
         );
  OAI22_X1 U6119 ( .A1(n4976), .A2(n6499), .B1(n6430), .B2(n4975), .ZN(n4972)
         );
  AOI21_X1 U6120 ( .B1(n6495), .B2(n4978), .A(n4972), .ZN(n4974) );
  NAND2_X1 U6121 ( .A1(n4979), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4973) );
  OAI211_X1 U6122 ( .C1(n5755), .C2(n4982), .A(n4974), .B(n4973), .ZN(U3046)
         );
  OAI22_X1 U6123 ( .A1(n4976), .A2(n6467), .B1(n6525), .B2(n4975), .ZN(n4977)
         );
  AOI21_X1 U6124 ( .B1(n6520), .B2(n4978), .A(n4977), .ZN(n4981) );
  NAND2_X1 U6125 ( .A1(n4979), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4980) );
  OAI211_X1 U6126 ( .C1(n4982), .C2(n5178), .A(n4981), .B(n4980), .ZN(U3050)
         );
  INV_X1 U6127 ( .A(n5034), .ZN(n4983) );
  OAI21_X1 U6128 ( .B1(n4985), .B2(n4984), .A(n4983), .ZN(n6178) );
  AOI22_X1 U6129 ( .A1(n6295), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n6291), .ZN(n4986) );
  OAI21_X1 U6130 ( .B1(n6178), .B2(n6285), .A(n4986), .ZN(U2883) );
  INV_X1 U6131 ( .A(n6175), .ZN(n4987) );
  AOI22_X1 U6132 ( .A1(n6279), .A2(n4987), .B1(EBX_REG_8__SCAN_IN), .B2(n5422), 
        .ZN(n4988) );
  OAI21_X1 U6133 ( .B1(n6178), .B2(n5456), .A(n4988), .ZN(U2851) );
  NAND2_X1 U6134 ( .A1(n5034), .A2(n5033), .ZN(n5110) );
  OAI21_X1 U6135 ( .B1(n5034), .B2(n5033), .A(n5110), .ZN(n6169) );
  AOI22_X1 U6136 ( .A1(n6295), .A2(DATAI_9_), .B1(EAX_REG_9__SCAN_IN), .B2(
        n6291), .ZN(n4989) );
  OAI21_X1 U6137 ( .B1(n6169), .B2(n6285), .A(n4989), .ZN(U2882) );
  OAI21_X1 U6138 ( .B1(n4992), .B2(n4991), .A(n4990), .ZN(n6166) );
  INV_X1 U6139 ( .A(n6166), .ZN(n6355) );
  AOI22_X1 U6140 ( .A1(n6279), .A2(n6355), .B1(EBX_REG_9__SCAN_IN), .B2(n5422), 
        .ZN(n4993) );
  OAI21_X1 U6141 ( .B1(n6169), .B2(n5456), .A(n4993), .ZN(U2850) );
  INV_X1 U6142 ( .A(n6408), .ZN(n5830) );
  NAND2_X1 U6143 ( .A1(n5830), .A2(n4527), .ZN(n5001) );
  INV_X1 U6144 ( .A(n5001), .ZN(n4996) );
  NOR2_X1 U6145 ( .A1(n4994), .A2(n6563), .ZN(n4995) );
  AOI22_X1 U6146 ( .A1(n4996), .A2(n6471), .B1(n6405), .B2(n4995), .ZN(n5028)
         );
  INV_X1 U6147 ( .A(n5834), .ZN(n5837) );
  NOR2_X1 U6148 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5837), .ZN(n5021)
         );
  NAND2_X1 U6149 ( .A1(n5736), .A2(n4997), .ZN(n5824) );
  INV_X1 U6150 ( .A(n5833), .ZN(n4998) );
  INV_X1 U6151 ( .A(n5866), .ZN(n5880) );
  OAI22_X1 U6152 ( .A1(n5824), .A2(n6487), .B1(n6424), .B2(n5880), .ZN(n4999)
         );
  AOI21_X1 U6153 ( .B1(n6470), .B2(n5021), .A(n4999), .ZN(n5007) );
  INV_X1 U6154 ( .A(n5824), .ZN(n5000) );
  NOR3_X1 U6155 ( .A1(n5000), .A2(n5866), .A3(n6477), .ZN(n5002) );
  OAI21_X1 U6156 ( .B1(n5002), .B2(n6416), .A(n5001), .ZN(n5005) );
  NOR2_X1 U6157 ( .A1(n5156), .A2(n5003), .ZN(n6420) );
  INV_X1 U6158 ( .A(n5021), .ZN(n5032) );
  AOI21_X1 U6159 ( .B1(n5032), .B2(STATE2_REG_3__SCAN_IN), .A(n6563), .ZN(
        n5004) );
  NAND3_X1 U6160 ( .A1(n5005), .A2(n6420), .A3(n5004), .ZN(n5027) );
  NAND2_X1 U6161 ( .A1(n5027), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n5006)
         );
  OAI211_X1 U6162 ( .C1(n5747), .C2(n5028), .A(n5007), .B(n5006), .ZN(U3132)
         );
  OAI22_X1 U6163 ( .A1(n5824), .A2(n5807), .B1(n6511), .B2(n5880), .ZN(n5008)
         );
  AOI21_X1 U6164 ( .B1(n6507), .B2(n5021), .A(n5008), .ZN(n5010) );
  NAND2_X1 U6165 ( .A1(n5027), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n5009)
         );
  OAI211_X1 U6166 ( .C1(n5763), .C2(n5028), .A(n5010), .B(n5009), .ZN(U3136)
         );
  OAI22_X1 U6167 ( .A1(n5824), .A2(n6458), .B1(n6517), .B2(n5880), .ZN(n5011)
         );
  AOI21_X1 U6168 ( .B1(n6513), .B2(n5021), .A(n5011), .ZN(n5013) );
  NAND2_X1 U6169 ( .A1(n5027), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n5012)
         );
  OAI211_X1 U6170 ( .C1(n5768), .C2(n5028), .A(n5013), .B(n5012), .ZN(U3137)
         );
  OAI22_X1 U6171 ( .A1(n5824), .A2(n6499), .B1(n6430), .B2(n5880), .ZN(n5014)
         );
  AOI21_X1 U6172 ( .B1(n6495), .B2(n5021), .A(n5014), .ZN(n5016) );
  NAND2_X1 U6173 ( .A1(n5027), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n5015)
         );
  OAI211_X1 U6174 ( .C1(n5755), .C2(n5028), .A(n5016), .B(n5015), .ZN(U3134)
         );
  OAI22_X1 U6175 ( .A1(n5824), .A2(n6505), .B1(n6434), .B2(n5880), .ZN(n5017)
         );
  AOI21_X1 U6176 ( .B1(n6501), .B2(n5021), .A(n5017), .ZN(n5019) );
  NAND2_X1 U6177 ( .A1(n5027), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n5018)
         );
  OAI211_X1 U6178 ( .C1(n5759), .C2(n5028), .A(n5019), .B(n5018), .ZN(U3135)
         );
  OAI22_X1 U6179 ( .A1(n5824), .A2(n5794), .B1(n6493), .B2(n5880), .ZN(n5020)
         );
  AOI21_X1 U6180 ( .B1(n6489), .B2(n5021), .A(n5020), .ZN(n5023) );
  NAND2_X1 U6181 ( .A1(n5027), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n5022)
         );
  OAI211_X1 U6182 ( .C1(n5751), .C2(n5028), .A(n5023), .B(n5022), .ZN(U3133)
         );
  NAND2_X1 U6183 ( .A1(n5027), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n5026)
         );
  OAI22_X1 U6184 ( .A1(n5824), .A2(n6467), .B1(n5028), .B2(n5178), .ZN(n5024)
         );
  AOI21_X1 U6185 ( .B1(n6460), .B2(n5866), .A(n5024), .ZN(n5025) );
  OAI211_X1 U6186 ( .C1(n5032), .C2(n5773), .A(n5026), .B(n5025), .ZN(U3138)
         );
  NAND2_X1 U6187 ( .A1(n5027), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n5031)
         );
  OAI22_X1 U6188 ( .A1(n5824), .A2(n6536), .B1(n5028), .B2(n5182), .ZN(n5029)
         );
  AOI21_X1 U6189 ( .B1(n6527), .B2(n5866), .A(n5029), .ZN(n5030) );
  OAI211_X1 U6190 ( .C1(n5032), .C2(n5780), .A(n5031), .B(n5030), .ZN(U3139)
         );
  AND2_X1 U6191 ( .A1(n5034), .A2(n5033), .ZN(n5036) );
  AND2_X1 U6192 ( .A1(n5036), .A2(n5035), .ZN(n5140) );
  OAI21_X1 U6193 ( .B1(n5140), .B2(n5037), .A(n3807), .ZN(n6133) );
  INV_X1 U6194 ( .A(DATAI_12_), .ZN(n5039) );
  OAI222_X1 U6195 ( .A1(n6133), .A2(n6285), .B1(n5039), .B2(n5107), .C1(n5038), 
        .C2(n6299), .ZN(U2879) );
  INV_X1 U6196 ( .A(n5040), .ZN(n6213) );
  AOI21_X1 U6197 ( .B1(n6341), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n5041), 
        .ZN(n5042) );
  OAI21_X1 U6198 ( .B1(n6335), .B2(n6218), .A(n5042), .ZN(n5043) );
  AOI21_X1 U6199 ( .B1(n6213), .B2(n6329), .A(n5043), .ZN(n5044) );
  OAI21_X1 U6200 ( .B1(n6073), .B2(n5045), .A(n5044), .ZN(U2981) );
  INV_X1 U6201 ( .A(n6202), .ZN(n5048) );
  AOI21_X1 U6202 ( .B1(n6341), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n5046), 
        .ZN(n5047) );
  OAI21_X1 U6203 ( .B1(n6335), .B2(n5048), .A(n5047), .ZN(n5049) );
  AOI21_X1 U6204 ( .B1(n6204), .B2(n6329), .A(n5049), .ZN(n5050) );
  OAI21_X1 U6205 ( .B1(n6073), .B2(n5051), .A(n5050), .ZN(U2980) );
  INV_X1 U6206 ( .A(n5052), .ZN(n6232) );
  AOI22_X1 U6207 ( .A1(n6341), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6395), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n5053) );
  OAI21_X1 U6208 ( .B1(n6335), .B2(n6232), .A(n5053), .ZN(n5054) );
  AOI21_X1 U6209 ( .B1(n6223), .B2(n6329), .A(n5054), .ZN(n5055) );
  OAI21_X1 U6210 ( .B1(n6073), .B2(n5056), .A(n5055), .ZN(U2982) );
  XNOR2_X1 U6211 ( .A(n5057), .B(n5058), .ZN(n6367) );
  INV_X1 U6212 ( .A(n6194), .ZN(n5061) );
  INV_X1 U6213 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6623) );
  NOR2_X1 U6214 ( .A1(n6187), .A2(n6623), .ZN(n6363) );
  AOI21_X1 U6215 ( .B1(n6341), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n6363), 
        .ZN(n5059) );
  OAI21_X1 U6216 ( .B1(n6335), .B2(n6199), .A(n5059), .ZN(n5060) );
  AOI21_X1 U6217 ( .B1(n5061), .B2(n6329), .A(n5060), .ZN(n5062) );
  OAI21_X1 U6218 ( .B1(n6073), .B2(n6367), .A(n5062), .ZN(U2979) );
  AOI21_X1 U6219 ( .B1(n6341), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n5063), 
        .ZN(n5064) );
  OAI21_X1 U6220 ( .B1(n6335), .B2(n6243), .A(n5064), .ZN(n5065) );
  AOI21_X1 U6221 ( .B1(n6329), .B2(n6233), .A(n5065), .ZN(n5066) );
  OAI21_X1 U6222 ( .B1(n6073), .B2(n5067), .A(n5066), .ZN(U2983) );
  AOI22_X1 U6223 ( .A1(n6674), .A2(UWORD_REG_2__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n5068) );
  OAI21_X1 U6224 ( .B1(n5069), .B2(n5084), .A(n5068), .ZN(U2905) );
  AOI22_X1 U6225 ( .A1(n6674), .A2(UWORD_REG_3__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n5070) );
  OAI21_X1 U6226 ( .B1(n5071), .B2(n5084), .A(n5070), .ZN(U2904) );
  AOI22_X1 U6227 ( .A1(n6674), .A2(UWORD_REG_0__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n5072) );
  OAI21_X1 U6228 ( .B1(n6962), .B2(n5084), .A(n5072), .ZN(U2907) );
  AOI22_X1 U6229 ( .A1(n6674), .A2(UWORD_REG_4__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n5073) );
  OAI21_X1 U6230 ( .B1(n3926), .B2(n5084), .A(n5073), .ZN(U2903) );
  AOI22_X1 U6231 ( .A1(n6674), .A2(UWORD_REG_1__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n5074) );
  OAI21_X1 U6232 ( .B1(n3873), .B2(n5084), .A(n5074), .ZN(U2906) );
  AOI22_X1 U6233 ( .A1(n5082), .A2(UWORD_REG_9__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n5075) );
  OAI21_X1 U6234 ( .B1(n6829), .B2(n5084), .A(n5075), .ZN(U2898) );
  AOI22_X1 U6235 ( .A1(n5082), .A2(UWORD_REG_6__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n5076) );
  OAI21_X1 U6236 ( .B1(n5077), .B2(n5084), .A(n5076), .ZN(U2901) );
  AOI22_X1 U6237 ( .A1(n5082), .A2(UWORD_REG_11__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n5078) );
  OAI21_X1 U6238 ( .B1(n4069), .B2(n5084), .A(n5078), .ZN(U2896) );
  AOI22_X1 U6239 ( .A1(n5082), .A2(UWORD_REG_14__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n5079) );
  OAI21_X1 U6240 ( .B1(n5080), .B2(n5084), .A(n5079), .ZN(U2893) );
  AOI22_X1 U6241 ( .A1(n5082), .A2(UWORD_REG_5__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n5081) );
  OAI21_X1 U6242 ( .B1(n6946), .B2(n5084), .A(n5081), .ZN(U2902) );
  AOI22_X1 U6243 ( .A1(n5082), .A2(UWORD_REG_7__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n5083) );
  OAI21_X1 U6244 ( .B1(n6791), .B2(n5084), .A(n5083), .ZN(U2900) );
  XNOR2_X1 U6245 ( .A(n3552), .B(n6749), .ZN(n5086) );
  XNOR2_X1 U6246 ( .A(n5085), .B(n5086), .ZN(n6356) );
  INV_X1 U6247 ( .A(n6073), .ZN(n6339) );
  NAND2_X1 U6248 ( .A1(n6356), .A2(n6339), .ZN(n5090) );
  NAND2_X1 U6249 ( .A1(n6395), .A2(REIP_REG_9__SCAN_IN), .ZN(n6353) );
  OAI21_X1 U6250 ( .B1(n5591), .B2(n5087), .A(n6353), .ZN(n5088) );
  AOI21_X1 U6251 ( .B1(n5593), .B2(n6171), .A(n5088), .ZN(n5089) );
  OAI211_X1 U6252 ( .C1(n6344), .C2(n6169), .A(n5090), .B(n5089), .ZN(U2977)
         );
  OR2_X1 U6253 ( .A1(n5092), .A2(n5091), .ZN(n5093) );
  NAND2_X1 U6254 ( .A1(n5094), .A2(n5093), .ZN(n6398) );
  INV_X1 U6255 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5099) );
  NOR2_X1 U6256 ( .A1(n5095), .A2(n6344), .ZN(n5098) );
  INV_X1 U6257 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5096) );
  OAI22_X1 U6258 ( .A1(n5591), .A2(n5099), .B1(n6187), .B2(n5096), .ZN(n5097)
         );
  AOI211_X1 U6259 ( .C1(n5593), .C2(n5099), .A(n5098), .B(n5097), .ZN(n5100)
         );
  OAI21_X1 U6260 ( .B1(n6073), .B2(n6398), .A(n5100), .ZN(U2985) );
  OAI21_X1 U6261 ( .B1(n5103), .B2(n5102), .A(n5131), .ZN(n6113) );
  INV_X1 U6262 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5105) );
  OAI21_X1 U6263 ( .B1(n5716), .B2(n5104), .A(n5134), .ZN(n6112) );
  OAI222_X1 U6264 ( .A1(n6113), .A2(n5456), .B1(n6284), .B2(n5105), .C1(n6112), 
        .C2(n6274), .ZN(U2845) );
  INV_X1 U6265 ( .A(DATAI_14_), .ZN(n5108) );
  OAI222_X1 U6266 ( .A1(n6113), .A2(n6285), .B1(n5108), .B2(n5107), .C1(n5106), 
        .C2(n6299), .ZN(U2877) );
  NAND2_X1 U6267 ( .A1(n5110), .A2(n5109), .ZN(n5111) );
  INV_X1 U6268 ( .A(n6155), .ZN(n5115) );
  AOI22_X1 U6269 ( .A1(n6295), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n6291), .ZN(n5112) );
  OAI21_X1 U6270 ( .B1(n5115), .B2(n6285), .A(n5112), .ZN(U2881) );
  INV_X1 U6271 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U6272 ( .A1(n4990), .A2(n5113), .ZN(n5114) );
  NAND2_X1 U6273 ( .A1(n5144), .A2(n5114), .ZN(n6151) );
  OAI222_X1 U6274 ( .A1(n5115), .A2(n5456), .B1(n6284), .B2(n6152), .C1(n6151), 
        .C2(n6274), .ZN(U2849) );
  INV_X1 U6275 ( .A(n5116), .ZN(n5118) );
  NAND2_X1 U6276 ( .A1(n5118), .A2(n5117), .ZN(n5119) );
  XNOR2_X1 U6277 ( .A(n5120), .B(n5119), .ZN(n5130) );
  INV_X1 U6278 ( .A(n6154), .ZN(n5122) );
  AOI22_X1 U6279 ( .A1(n6341), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .B1(n6395), 
        .B2(REIP_REG_10__SCAN_IN), .ZN(n5121) );
  OAI21_X1 U6280 ( .B1(n6335), .B2(n5122), .A(n5121), .ZN(n5123) );
  AOI21_X1 U6281 ( .B1(n6155), .B2(n6329), .A(n5123), .ZN(n5124) );
  OAI21_X1 U6282 ( .B1(n5130), .B2(n6073), .A(n5124), .ZN(U2976) );
  OAI21_X1 U6283 ( .B1(n5680), .B2(n5125), .A(n6370), .ZN(n6357) );
  INV_X1 U6284 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6159) );
  OAI22_X1 U6285 ( .A1(n6394), .A2(n6151), .B1(n6159), .B2(n6187), .ZN(n5128)
         );
  NAND2_X1 U6286 ( .A1(n5125), .A2(n6362), .ZN(n6360) );
  AOI221_X1 U6287 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .C1(n6749), .C2(n5126), .A(n6360), 
        .ZN(n5127) );
  AOI211_X1 U6288 ( .C1(INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n6357), .A(n5128), .B(n5127), .ZN(n5129) );
  OAI21_X1 U6289 ( .B1(n6399), .B2(n5130), .A(n5129), .ZN(U3008) );
  OAI21_X1 U6290 ( .B1(n3847), .B2(n3145), .A(n5248), .ZN(n5585) );
  INV_X1 U6291 ( .A(n5244), .ZN(n5133) );
  AOI21_X1 U6292 ( .B1(n5135), .B2(n5134), .A(n5133), .ZN(n6041) );
  AOI22_X1 U6293 ( .A1(n6041), .A2(n6279), .B1(EBX_REG_15__SCAN_IN), .B2(n5422), .ZN(n5136) );
  OAI21_X1 U6294 ( .B1(n5585), .B2(n5456), .A(n5136), .ZN(U2844) );
  AOI22_X1 U6295 ( .A1(n6295), .A2(DATAI_15_), .B1(EAX_REG_15__SCAN_IN), .B2(
        n6291), .ZN(n5137) );
  OAI21_X1 U6296 ( .B1(n5585), .B2(n6285), .A(n5137), .ZN(U2876) );
  AND2_X1 U6297 ( .A1(n5139), .A2(n5138), .ZN(n5141) );
  AOI22_X1 U6298 ( .A1(n6295), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6291), .ZN(n5142) );
  OAI21_X1 U6299 ( .B1(n6145), .B2(n6285), .A(n5142), .ZN(U2880) );
  NAND2_X1 U6300 ( .A1(n5144), .A2(n5143), .ZN(n5145) );
  NAND2_X1 U6301 ( .A1(n5712), .A2(n5145), .ZN(n6142) );
  INV_X1 U6302 ( .A(n6142), .ZN(n6347) );
  AOI22_X1 U6303 ( .A1(n6279), .A2(n6347), .B1(EBX_REG_11__SCAN_IN), .B2(n5422), .ZN(n5146) );
  OAI21_X1 U6304 ( .B1(n6145), .B2(n5456), .A(n5146), .ZN(U2848) );
  OAI21_X1 U6305 ( .B1(n5591), .B2(n6838), .A(n5147), .ZN(n5149) );
  NOR2_X1 U6306 ( .A1(n6178), .A2(n6344), .ZN(n5148) );
  AOI211_X1 U6307 ( .C1(n5593), .C2(n6179), .A(n5149), .B(n5148), .ZN(n5150)
         );
  OAI21_X1 U6308 ( .B1(n6073), .B2(n5151), .A(n5150), .ZN(U2978) );
  NAND2_X1 U6309 ( .A1(n5734), .A2(n5153), .ZN(n6535) );
  AOI21_X1 U6310 ( .B1(n5188), .B2(n6535), .A(n6072), .ZN(n5154) );
  NOR2_X1 U6311 ( .A1(n5154), .A2(n6477), .ZN(n5159) );
  AND2_X1 U6312 ( .A1(n5155), .A2(n4527), .ZN(n6475) );
  INV_X1 U6313 ( .A(n5156), .ZN(n5742) );
  NOR2_X1 U6314 ( .A1(n5742), .A2(n6563), .ZN(n5157) );
  AOI22_X1 U6315 ( .A1(n5159), .A2(n6475), .B1(n6405), .B2(n5157), .ZN(n5192)
         );
  NAND3_X1 U6316 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n6557), .ZN(n6481) );
  NOR2_X1 U6317 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6481), .ZN(n5190)
         );
  INV_X1 U6318 ( .A(n5190), .ZN(n5160) );
  INV_X1 U6319 ( .A(n6475), .ZN(n5158) );
  AOI22_X1 U6320 ( .A1(STATE2_REG_3__SCAN_IN), .A2(n5160), .B1(n5159), .B2(
        n5158), .ZN(n5161) );
  OAI211_X1 U6321 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n4606), .A(n5162), .B(n5161), .ZN(n5186) );
  AOI22_X1 U6322 ( .A1(n6518), .A2(n6455), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5186), .ZN(n5163) );
  OAI21_X1 U6323 ( .B1(n5188), .B2(n6458), .A(n5163), .ZN(n5164) );
  AOI21_X1 U6324 ( .B1(n6513), .B2(n5190), .A(n5164), .ZN(n5165) );
  OAI21_X1 U6325 ( .B1(n5768), .B2(n5192), .A(n5165), .ZN(U3105) );
  AOI22_X1 U6326 ( .A1(n6518), .A2(n6494), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5186), .ZN(n5166) );
  OAI21_X1 U6327 ( .B1(n5188), .B2(n6499), .A(n5166), .ZN(n5167) );
  AOI21_X1 U6328 ( .B1(n6495), .B2(n5190), .A(n5167), .ZN(n5168) );
  OAI21_X1 U6329 ( .B1(n5755), .B2(n5192), .A(n5168), .ZN(U3102) );
  AOI22_X1 U6330 ( .A1(n6518), .A2(n6500), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5186), .ZN(n5169) );
  OAI21_X1 U6331 ( .B1(n5188), .B2(n6505), .A(n5169), .ZN(n5170) );
  AOI21_X1 U6332 ( .B1(n6501), .B2(n5190), .A(n5170), .ZN(n5171) );
  OAI21_X1 U6333 ( .B1(n5759), .B2(n5192), .A(n5171), .ZN(U3103) );
  AOI22_X1 U6334 ( .A1(n6518), .A2(n6469), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5186), .ZN(n5172) );
  OAI21_X1 U6335 ( .B1(n5188), .B2(n6487), .A(n5172), .ZN(n5173) );
  AOI21_X1 U6336 ( .B1(n6470), .B2(n5190), .A(n5173), .ZN(n5174) );
  OAI21_X1 U6337 ( .B1(n5747), .B2(n5192), .A(n5174), .ZN(U3100) );
  AOI22_X1 U6338 ( .A1(n6518), .A2(n6460), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5186), .ZN(n5175) );
  OAI21_X1 U6339 ( .B1(n5188), .B2(n6467), .A(n5175), .ZN(n5176) );
  AOI21_X1 U6340 ( .B1(n6520), .B2(n5190), .A(n5176), .ZN(n5177) );
  OAI21_X1 U6341 ( .B1(n5192), .B2(n5178), .A(n5177), .ZN(U3106) );
  AOI22_X1 U6342 ( .A1(n6518), .A2(n6527), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5186), .ZN(n5179) );
  OAI21_X1 U6343 ( .B1(n5188), .B2(n6536), .A(n5179), .ZN(n5180) );
  AOI21_X1 U6344 ( .B1(n6529), .B2(n5190), .A(n5180), .ZN(n5181) );
  OAI21_X1 U6345 ( .B1(n5192), .B2(n5182), .A(n5181), .ZN(U3107) );
  AOI22_X1 U6346 ( .A1(n6518), .A2(n5844), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5186), .ZN(n5183) );
  OAI21_X1 U6347 ( .B1(n5188), .B2(n5794), .A(n5183), .ZN(n5184) );
  AOI21_X1 U6348 ( .B1(n6489), .B2(n5190), .A(n5184), .ZN(n5185) );
  OAI21_X1 U6349 ( .B1(n5751), .B2(n5192), .A(n5185), .ZN(U3101) );
  AOI22_X1 U6350 ( .A1(n6518), .A2(n5860), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5186), .ZN(n5187) );
  OAI21_X1 U6351 ( .B1(n5188), .B2(n5807), .A(n5187), .ZN(n5189) );
  AOI21_X1 U6352 ( .B1(n6507), .B2(n5190), .A(n5189), .ZN(n5191) );
  OAI21_X1 U6353 ( .B1(n5763), .B2(n5192), .A(n5191), .ZN(U3104) );
  NOR3_X1 U6354 ( .A1(n6585), .A2(n6663), .A3(n6578), .ZN(n6575) );
  NAND2_X1 U6355 ( .A1(n5194), .A2(n5193), .ZN(n6588) );
  NAND2_X1 U6356 ( .A1(n6187), .A2(n6588), .ZN(n5195) );
  OR2_X1 U6357 ( .A1(n6575), .A2(n5195), .ZN(n5196) );
  OAI21_X1 U6358 ( .B1(n5212), .B2(n5198), .A(n6193), .ZN(n6264) );
  INV_X1 U6359 ( .A(n6264), .ZN(n5219) );
  NAND2_X1 U6360 ( .A1(n6673), .A2(n6072), .ZN(n5206) );
  INV_X1 U6361 ( .A(n5206), .ZN(n5199) );
  AND2_X1 U6362 ( .A1(n5203), .A2(n5199), .ZN(n5200) );
  AND2_X1 U6363 ( .A1(n5201), .A2(n5200), .ZN(n5202) );
  NAND2_X1 U6364 ( .A1(n6239), .A2(n6271), .ZN(n5919) );
  NOR2_X1 U6365 ( .A1(n6601), .A2(n5206), .ZN(n6570) );
  NOR2_X1 U6366 ( .A1(n6676), .A2(n6570), .ZN(n5334) );
  INV_X1 U6367 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5374) );
  AND3_X1 U6368 ( .A1(n5203), .A2(n5374), .A3(n5206), .ZN(n5204) );
  NOR2_X1 U6369 ( .A1(n5334), .A2(n5204), .ZN(n5205) );
  NAND3_X1 U6370 ( .A1(n5207), .A2(EBX_REG_31__SCAN_IN), .A3(n5206), .ZN(n5208) );
  NOR2_X2 U6371 ( .A1(n5212), .A2(n5208), .ZN(n6262) );
  OAI22_X1 U6372 ( .A1(n6903), .A2(n6220), .B1(n6176), .B2(n5209), .ZN(n5210)
         );
  AOI21_X1 U6373 ( .B1(REIP_REG_0__SCAN_IN), .B2(n5919), .A(n5210), .ZN(n5218)
         );
  NOR2_X1 U6374 ( .A1(n5212), .A2(n5211), .ZN(n6260) );
  NOR2_X1 U6375 ( .A1(n5213), .A2(n5295), .ZN(n5214) );
  AOI21_X1 U6376 ( .B1(n6256), .B2(n6254), .A(n5215), .ZN(n5216) );
  AOI21_X1 U6377 ( .B1(n6260), .B2(n6474), .A(n5216), .ZN(n5217) );
  OAI211_X1 U6378 ( .C1(n5219), .C2(n6345), .A(n5218), .B(n5217), .ZN(U2827)
         );
  NAND2_X1 U6379 ( .A1(n5222), .A2(n5221), .ZN(n5223) );
  XNOR2_X1 U6380 ( .A(n5220), .B(n5223), .ZN(n6349) );
  NAND2_X1 U6381 ( .A1(n6349), .A2(n6339), .ZN(n5226) );
  AND2_X1 U6382 ( .A1(n6395), .A2(REIP_REG_11__SCAN_IN), .ZN(n6346) );
  NOR2_X1 U6383 ( .A1(n6335), .A2(n6141), .ZN(n5224) );
  AOI211_X1 U6384 ( .C1(n6341), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6346), 
        .B(n5224), .ZN(n5225) );
  OAI211_X1 U6385 ( .C1(n6344), .C2(n6145), .A(n5226), .B(n5225), .ZN(U2975)
         );
  XNOR2_X1 U6386 ( .A(n3552), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n5228)
         );
  XNOR2_X1 U6387 ( .A(n5227), .B(n5228), .ZN(n5242) );
  INV_X1 U6388 ( .A(REIP_REG_12__SCAN_IN), .ZN(n5229) );
  OAI22_X1 U6389 ( .A1(n5591), .A2(n6914), .B1(n6187), .B2(n5229), .ZN(n5231)
         );
  NOR2_X1 U6390 ( .A1(n6133), .A2(n6344), .ZN(n5230) );
  AOI211_X1 U6391 ( .C1(n5593), .C2(n6134), .A(n5231), .B(n5230), .ZN(n5232)
         );
  OAI21_X1 U6392 ( .B1(n5242), .B2(n6073), .A(n5232), .ZN(U2974) );
  XNOR2_X1 U6393 ( .A(n5712), .B(n5714), .ZN(n6278) );
  NOR2_X1 U6394 ( .A1(n6187), .A2(n5229), .ZN(n5240) );
  INV_X1 U6395 ( .A(n6348), .ZN(n5233) );
  NOR2_X1 U6396 ( .A1(n5233), .A2(n6882), .ZN(n5238) );
  NAND2_X1 U6397 ( .A1(n5235), .A2(n5234), .ZN(n5679) );
  INV_X1 U6398 ( .A(n6352), .ZN(n5698) );
  AOI21_X1 U6399 ( .B1(n6882), .B2(n5679), .A(n5698), .ZN(n5236) );
  INV_X1 U6400 ( .A(n5236), .ZN(n5237) );
  MUX2_X1 U6401 ( .A(n5238), .B(n5237), .S(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .Z(n5239) );
  AOI211_X1 U6402 ( .C1(n6375), .C2(n6278), .A(n5240), .B(n5239), .ZN(n5241)
         );
  OAI21_X1 U6403 ( .B1(n5242), .B2(n6399), .A(n5241), .ZN(U3006) );
  AND2_X1 U6404 ( .A1(n5244), .A2(n5243), .ZN(n5245) );
  OR2_X1 U6405 ( .A1(n5245), .A2(n6030), .ZN(n6110) );
  INV_X1 U6406 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5251) );
  AOI21_X1 U6407 ( .B1(n5249), .B2(n5248), .A(n5247), .ZN(n6290) );
  INV_X1 U6408 ( .A(n6290), .ZN(n5250) );
  OAI222_X1 U6409 ( .A1(n6110), .A2(n6274), .B1(n6284), .B2(n5251), .C1(n5250), 
        .C2(n5456), .ZN(U2843) );
  INV_X1 U6410 ( .A(n5252), .ZN(n6009) );
  INV_X1 U6411 ( .A(n5253), .ZN(n5256) );
  OAI21_X1 U6412 ( .B1(n6009), .B2(n5256), .A(n5450), .ZN(n5568) );
  INV_X1 U6413 ( .A(n6271), .ZN(n5258) );
  INV_X1 U6414 ( .A(REIP_REG_13__SCAN_IN), .ZN(n5257) );
  INV_X1 U6415 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6629) );
  INV_X1 U6416 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6626) );
  INV_X1 U6417 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6387) );
  NOR3_X1 U6418 ( .A1(n5096), .A2(n6387), .A3(n6615), .ZN(n6222) );
  NAND2_X1 U6419 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6222), .ZN(n6212) );
  NOR2_X1 U6420 ( .A1(n6620), .A2(n6212), .ZN(n6196) );
  NAND2_X1 U6421 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6196), .ZN(n6185) );
  NOR2_X1 U6422 ( .A1(n6623), .A2(n6185), .ZN(n6174) );
  NAND2_X1 U6423 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6174), .ZN(n6157) );
  NOR2_X1 U6424 ( .A1(n6626), .A2(n6157), .ZN(n6158) );
  NAND2_X1 U6425 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6158), .ZN(n6138) );
  NOR2_X1 U6426 ( .A1(n6629), .A2(n6138), .ZN(n6131) );
  NAND2_X1 U6427 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6131), .ZN(n6121) );
  NOR2_X1 U6428 ( .A1(n5257), .A2(n6121), .ZN(n6116) );
  NAND2_X1 U6429 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6116), .ZN(n5260) );
  NOR2_X1 U6430 ( .A1(n5258), .A2(n5260), .ZN(n5272) );
  NAND4_X1 U6431 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .A4(n5272), .ZN(n5336) );
  AND2_X1 U6432 ( .A1(n5919), .A2(n5336), .ZN(n6097) );
  AOI22_X1 U6433 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6261), .B1(
        REIP_REG_18__SCAN_IN), .B2(n6097), .ZN(n5259) );
  OAI211_X1 U6434 ( .C1(n6256), .C2(n5563), .A(n5259), .B(n6187), .ZN(n5268)
         );
  INV_X1 U6435 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6979) );
  INV_X1 U6436 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6636) );
  NOR2_X1 U6437 ( .A1(n6239), .A2(n5260), .ZN(n6102) );
  NAND3_X1 U6438 ( .A1(n6102), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n6093) );
  NOR2_X1 U6439 ( .A1(n6636), .A2(n6093), .ZN(n5977) );
  AND2_X1 U6440 ( .A1(n6979), .A2(n5977), .ZN(n5985) );
  INV_X1 U6441 ( .A(n5261), .ZN(n5445) );
  INV_X1 U6442 ( .A(n5262), .ZN(n5263) );
  MUX2_X1 U6443 ( .A(n5445), .B(n5263), .S(n5444), .Z(n5264) );
  NAND2_X1 U6444 ( .A1(n6032), .A2(n5264), .ZN(n5454) );
  OR2_X1 U6445 ( .A1(n6032), .A2(n5264), .ZN(n5265) );
  AND2_X1 U6446 ( .A1(n5454), .A2(n5265), .ZN(n6024) );
  INV_X1 U6447 ( .A(n6024), .ZN(n5279) );
  INV_X1 U6448 ( .A(n5565), .ZN(n5266) );
  OAI22_X1 U6449 ( .A1(n5279), .A2(n6176), .B1(n5266), .B2(n6254), .ZN(n5267)
         );
  NOR3_X1 U6450 ( .A1(n5268), .A2(n5985), .A3(n5267), .ZN(n5269) );
  OAI21_X1 U6451 ( .B1(n5568), .B2(n6193), .A(n5269), .ZN(U2809) );
  INV_X1 U6452 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6634) );
  INV_X1 U6453 ( .A(n6041), .ZN(n5271) );
  INV_X1 U6454 ( .A(n5582), .ZN(n5270) );
  OAI22_X1 U6455 ( .A1(n6176), .A2(n5271), .B1(n6254), .B2(n5270), .ZN(n5275)
         );
  INV_X1 U6456 ( .A(n5919), .ZN(n5948) );
  NOR2_X1 U6457 ( .A1(n5948), .A2(n5272), .ZN(n6111) );
  AOI22_X1 U6458 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6261), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6111), .ZN(n5273) );
  OAI211_X1 U6459 ( .C1(n6256), .C2(n6977), .A(n5273), .B(n6187), .ZN(n5274)
         );
  AOI211_X1 U6460 ( .C1(n6102), .C2(n6634), .A(n5275), .B(n5274), .ZN(n5276)
         );
  OAI21_X1 U6461 ( .B1(n5585), .B2(n6193), .A(n5276), .ZN(U2812) );
  AOI22_X1 U6462 ( .A1(n6289), .A2(DATAI_18_), .B1(n6291), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5278) );
  NAND2_X1 U6463 ( .A1(n6292), .A2(DATAI_2_), .ZN(n5277) );
  OAI211_X1 U6464 ( .C1(n5568), .C2(n6285), .A(n5278), .B(n5277), .ZN(U2873)
         );
  OAI222_X1 U6465 ( .A1(n5568), .A2(n5456), .B1(n5280), .B2(n6284), .C1(n6274), 
        .C2(n5279), .ZN(U2841) );
  AOI22_X1 U6466 ( .A1(n6548), .A2(n6583), .B1(FLUSH_REG_SCAN_IN), .B2(n6591), 
        .ZN(n6058) );
  NAND2_X1 U6467 ( .A1(n6661), .A2(n6058), .ZN(n6064) );
  INV_X1 U6468 ( .A(n5292), .ZN(n6545) );
  INV_X1 U6469 ( .A(n5281), .ZN(n5293) );
  OAI21_X1 U6470 ( .B1(n5285), .B2(n5287), .A(n5293), .ZN(n5282) );
  OAI21_X1 U6471 ( .B1(n6545), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n5282), 
        .ZN(n5283) );
  AOI21_X1 U6472 ( .B1(n6259), .B2(n5294), .A(n5283), .ZN(n6547) );
  INV_X1 U6473 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5284) );
  AOI22_X1 U6474 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5284), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4201), .ZN(n5312) );
  NOR2_X1 U6475 ( .A1(n5295), .A2(n6391), .ZN(n5296) );
  AOI22_X1 U6476 ( .A1(n5312), .A2(n5296), .B1(n5285), .B2(n5308), .ZN(n5286)
         );
  OAI21_X1 U6477 ( .B1(n6547), .B2(n5291), .A(n5286), .ZN(n5288) );
  AOI22_X1 U6478 ( .A1(n6064), .A2(n5288), .B1(n5287), .B2(n5308), .ZN(n5289)
         );
  OAI21_X1 U6479 ( .B1(n6064), .B2(n5290), .A(n5289), .ZN(U3460) );
  INV_X1 U6480 ( .A(n5291), .ZN(n6059) );
  INV_X1 U6481 ( .A(n6064), .ZN(n5315) );
  AOI21_X1 U6482 ( .B1(n6059), .B2(n5292), .A(n5315), .ZN(n5299) );
  AOI22_X1 U6483 ( .A1(n6474), .A2(n5294), .B1(n5293), .B2(n6546), .ZN(n6544)
         );
  OAI21_X1 U6484 ( .B1(n6544), .B2(STATE2_REG_3__SCAN_IN), .A(n5295), .ZN(
        n5297) );
  INV_X1 U6485 ( .A(n5296), .ZN(n5311) );
  AOI22_X1 U6486 ( .A1(n5297), .A2(n5311), .B1(n5308), .B2(n6546), .ZN(n5298)
         );
  OAI22_X1 U6487 ( .A1(n5299), .A2(n6546), .B1(n5298), .B2(n5315), .ZN(U3461)
         );
  INV_X1 U6488 ( .A(n5308), .ZN(n6577) );
  INV_X1 U6489 ( .A(n5300), .ZN(n5306) );
  AOI22_X1 U6490 ( .A1(n5302), .A2(n6059), .B1(n5301), .B2(n5308), .ZN(n5305)
         );
  AOI21_X1 U6491 ( .B1(n5308), .B2(n5303), .A(n5315), .ZN(n5318) );
  OAI222_X1 U6492 ( .A1(n6577), .A2(n5306), .B1(n5315), .B2(n5305), .C1(n5304), 
        .C2(n5318), .ZN(U3456) );
  INV_X1 U6493 ( .A(n5307), .ZN(n5314) );
  NAND3_X1 U6494 ( .A1(n5309), .A2(n5308), .A3(n5317), .ZN(n5310) );
  OAI21_X1 U6495 ( .B1(n5312), .B2(n5311), .A(n5310), .ZN(n5313) );
  AOI21_X1 U6496 ( .B1(n5314), .B2(n6059), .A(n5313), .ZN(n5316) );
  OAI22_X1 U6497 ( .A1(n5318), .A2(n5317), .B1(n5316), .B2(n5315), .ZN(U3459)
         );
  BUF_X2 U6498 ( .A(n5319), .Z(n5349) );
  NAND2_X1 U6499 ( .A1(n6299), .A2(n5320), .ZN(n5322) );
  AOI22_X1 U6500 ( .A1(n6289), .A2(DATAI_31_), .B1(n6291), .B2(
        EAX_REG_31__SCAN_IN), .ZN(n5321) );
  OAI21_X1 U6501 ( .B1(n5349), .B2(n5322), .A(n5321), .ZN(U2860) );
  INV_X1 U6502 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5376) );
  NOR2_X1 U6503 ( .A1(n5323), .A2(n5376), .ZN(n5326) );
  AOI21_X1 U6504 ( .B1(n5324), .B2(n5323), .A(n5326), .ZN(n5365) );
  NAND2_X1 U6505 ( .A1(n5383), .A2(n5365), .ZN(n5364) );
  INV_X1 U6506 ( .A(n5383), .ZN(n5325) );
  NAND2_X1 U6507 ( .A1(n5325), .A2(n5444), .ZN(n5328) );
  INV_X1 U6508 ( .A(n5326), .ZN(n5327) );
  OAI211_X1 U6509 ( .C1(n5364), .C2(n5329), .A(n5328), .B(n5327), .ZN(n5333)
         );
  OAI22_X1 U6510 ( .A1(n5331), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n5330), .ZN(n5332) );
  XNOR2_X1 U6511 ( .A(n5333), .B(n5332), .ZN(n5373) );
  NAND3_X1 U6512 ( .A1(n6671), .A2(EBX_REG_31__SCAN_IN), .A3(n5334), .ZN(n5335) );
  OAI21_X1 U6513 ( .B1(n6256), .B2(n6818), .A(n5335), .ZN(n5343) );
  INV_X1 U6514 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6641) );
  NAND2_X1 U6515 ( .A1(REIP_REG_18__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n5337) );
  NOR3_X1 U6516 ( .A1(n6641), .A2(n5337), .A3(n5336), .ZN(n5947) );
  NAND4_X1 U6517 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5947), .ZN(n5918) );
  INV_X1 U6518 ( .A(n5918), .ZN(n5339) );
  NAND3_X1 U6519 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5344) );
  INV_X1 U6520 ( .A(n5344), .ZN(n5338) );
  NAND2_X1 U6521 ( .A1(n5339), .A2(n5338), .ZN(n5340) );
  AND2_X1 U6522 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5345) );
  NOR2_X1 U6523 ( .A1(n6239), .A2(n5345), .ZN(n5341) );
  OR2_X1 U6524 ( .A1(n5906), .A2(n5341), .ZN(n5886) );
  INV_X1 U6525 ( .A(REIP_REG_29__SCAN_IN), .ZN(n5492) );
  NOR2_X1 U6526 ( .A1(n5886), .A2(n5492), .ZN(n5368) );
  INV_X1 U6527 ( .A(REIP_REG_31__SCAN_IN), .ZN(n5346) );
  NOR2_X1 U6528 ( .A1(n5906), .A2(n6244), .ZN(n5351) );
  AOI211_X1 U6529 ( .C1(n5368), .C2(REIP_REG_30__SCAN_IN), .A(n5346), .B(n5351), .ZN(n5342) );
  AOI211_X1 U6530 ( .C1(n6262), .C2(n5373), .A(n5343), .B(n5342), .ZN(n5348)
         );
  NAND3_X1 U6531 ( .A1(n5977), .A2(REIP_REG_18__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .ZN(n5969) );
  NOR2_X1 U6532 ( .A1(n6641), .A2(n5969), .ZN(n5960) );
  NAND4_X1 U6533 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5960), .ZN(n5920) );
  NOR2_X1 U6534 ( .A1(n5920), .A2(n5344), .ZN(n5898) );
  AND2_X1 U6535 ( .A1(n5898), .A2(n5345), .ZN(n5370) );
  NAND4_X1 U6536 ( .A1(n5370), .A2(REIP_REG_29__SCAN_IN), .A3(
        REIP_REG_30__SCAN_IN), .A4(n5346), .ZN(n5347) );
  OAI211_X1 U6537 ( .C1(n5349), .C2(n6193), .A(n5348), .B(n5347), .ZN(U2796)
         );
  NAND3_X1 U6538 ( .A1(n5370), .A2(REIP_REG_29__SCAN_IN), .A3(n4161), .ZN(
        n5357) );
  NOR3_X1 U6539 ( .A1(n5351), .A2(n5368), .A3(n4161), .ZN(n5354) );
  INV_X1 U6540 ( .A(EBX_REG_30__SCAN_IN), .ZN(n6951) );
  OAI22_X1 U6541 ( .A1(n6951), .A2(n6220), .B1(n5352), .B2(n6256), .ZN(n5353)
         );
  AOI211_X1 U6542 ( .C1(n6258), .C2(n5355), .A(n5354), .B(n5353), .ZN(n5356)
         );
  OAI211_X1 U6543 ( .C1(n5375), .C2(n6176), .A(n5357), .B(n5356), .ZN(n5358)
         );
  INV_X1 U6544 ( .A(n5358), .ZN(n5359) );
  OAI21_X1 U6545 ( .B1(n5350), .B2(n6193), .A(n5359), .ZN(U2797) );
  AOI21_X1 U6546 ( .B1(n5362), .B2(n5380), .A(n5361), .ZN(n5496) );
  INV_X1 U6547 ( .A(n5496), .ZN(n5461) );
  OAI22_X1 U6548 ( .A1(n5363), .A2(n6256), .B1(n6254), .B2(n5494), .ZN(n5367)
         );
  OAI21_X1 U6549 ( .B1(n5383), .B2(n5365), .A(n5364), .ZN(n5613) );
  NOR2_X1 U6550 ( .A1(n5613), .A2(n6176), .ZN(n5366) );
  AOI211_X1 U6551 ( .C1(EBX_REG_29__SCAN_IN), .C2(n6261), .A(n5367), .B(n5366), 
        .ZN(n5372) );
  INV_X1 U6552 ( .A(n5368), .ZN(n5369) );
  OAI21_X1 U6553 ( .B1(n5370), .B2(REIP_REG_29__SCAN_IN), .A(n5369), .ZN(n5371) );
  OAI211_X1 U6554 ( .C1(n5461), .C2(n6193), .A(n5372), .B(n5371), .ZN(U2798)
         );
  OAI22_X1 U6555 ( .A1(n5607), .A2(n6274), .B1(n6284), .B2(n5374), .ZN(U2828)
         );
  OAI222_X1 U6556 ( .A1(n5350), .A2(n5456), .B1(n6284), .B2(n6951), .C1(n6274), 
        .C2(n5375), .ZN(U2829) );
  OAI222_X1 U6557 ( .A1(n5456), .A2(n5461), .B1(n5376), .B2(n6284), .C1(n5613), 
        .C2(n6274), .ZN(U2830) );
  OR2_X1 U6558 ( .A1(n5377), .A2(n5378), .ZN(n5379) );
  AND2_X1 U6559 ( .A1(n5380), .A2(n5379), .ZN(n5890) );
  INV_X1 U6560 ( .A(n5890), .ZN(n5464) );
  INV_X1 U6561 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6890) );
  NOR2_X1 U6562 ( .A1(n5389), .A2(n5381), .ZN(n5382) );
  OR2_X1 U6563 ( .A1(n5383), .A2(n5382), .ZN(n5888) );
  OAI222_X1 U6564 ( .A1(n5456), .A2(n5464), .B1(n6284), .B2(n6890), .C1(n5888), 
        .C2(n6274), .ZN(U2831) );
  INV_X1 U6565 ( .A(n5384), .ZN(n5392) );
  AND2_X1 U6566 ( .A1(n5392), .A2(n5385), .ZN(n5386) );
  OR2_X1 U6567 ( .A1(n5377), .A2(n5386), .ZN(n5900) );
  INV_X1 U6568 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5390) );
  NOR2_X1 U6569 ( .A1(n5396), .A2(n5387), .ZN(n5388) );
  OR2_X1 U6570 ( .A1(n5389), .A2(n5388), .ZN(n5899) );
  OAI222_X1 U6571 ( .A1(n5456), .A2(n5900), .B1(n5390), .B2(n6284), .C1(n5899), 
        .C2(n6274), .ZN(U2832) );
  INV_X1 U6572 ( .A(n5402), .ZN(n5394) );
  INV_X1 U6573 ( .A(n5391), .ZN(n5393) );
  OAI21_X1 U6574 ( .B1(n5394), .B2(n5393), .A(n5392), .ZN(n5909) );
  AND2_X1 U6575 ( .A1(n5405), .A2(n5395), .ZN(n5397) );
  OR2_X1 U6576 ( .A1(n5397), .A2(n5396), .ZN(n5914) );
  OAI22_X1 U6577 ( .A1(n5914), .A2(n6274), .B1(n5905), .B2(n6284), .ZN(n5398)
         );
  INV_X1 U6578 ( .A(n5398), .ZN(n5399) );
  OAI21_X1 U6579 ( .B1(n5909), .B2(n5456), .A(n5399), .ZN(U2833) );
  OR2_X1 U6580 ( .A1(n5409), .A2(n5400), .ZN(n5401) );
  AND2_X1 U6581 ( .A1(n5402), .A2(n5401), .ZN(n5992) );
  INV_X1 U6582 ( .A(n5992), .ZN(n5471) );
  INV_X1 U6583 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5406) );
  NAND2_X1 U6584 ( .A1(n5414), .A2(n5403), .ZN(n5404) );
  NAND2_X1 U6585 ( .A1(n5405), .A2(n5404), .ZN(n6015) );
  OAI222_X1 U6586 ( .A1(n5471), .A2(n5456), .B1(n5406), .B2(n6284), .C1(n6274), 
        .C2(n6015), .ZN(U2834) );
  INV_X1 U6587 ( .A(n5407), .ZN(n5411) );
  INV_X1 U6588 ( .A(n5408), .ZN(n5410) );
  AOI21_X1 U6589 ( .B1(n5411), .B2(n5410), .A(n5409), .ZN(n5930) );
  INV_X1 U6590 ( .A(n5930), .ZN(n5474) );
  INV_X1 U6591 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5415) );
  NAND2_X1 U6592 ( .A1(n5421), .A2(n5412), .ZN(n5413) );
  NAND2_X1 U6593 ( .A1(n5414), .A2(n5413), .ZN(n5935) );
  OAI222_X1 U6594 ( .A1(n5456), .A2(n5474), .B1(n6284), .B2(n5415), .C1(n5935), 
        .C2(n6274), .ZN(U2835) );
  INV_X1 U6595 ( .A(n5416), .ZN(n5427) );
  AOI21_X1 U6596 ( .B1(n5417), .B2(n5427), .A(n5408), .ZN(n5942) );
  INV_X1 U6597 ( .A(n5942), .ZN(n5477) );
  OR2_X1 U6598 ( .A1(n5418), .A2(n5419), .ZN(n5420) );
  AND2_X1 U6599 ( .A1(n5421), .A2(n5420), .ZN(n5937) );
  AOI22_X1 U6600 ( .A1(n5937), .A2(n6279), .B1(EBX_REG_23__SCAN_IN), .B2(n5422), .ZN(n5423) );
  OAI21_X1 U6601 ( .B1(n5477), .B2(n5456), .A(n5423), .ZN(U2836) );
  NOR2_X1 U6602 ( .A1(n5437), .A2(n5424), .ZN(n5425) );
  OR2_X1 U6603 ( .A1(n5418), .A2(n5425), .ZN(n5949) );
  INV_X1 U6604 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5430) );
  INV_X1 U6605 ( .A(n5427), .ZN(n5428) );
  AOI21_X1 U6606 ( .B1(n5429), .B2(n5434), .A(n5428), .ZN(n5951) );
  INV_X1 U6607 ( .A(n5951), .ZN(n5480) );
  OAI222_X1 U6608 ( .A1(n6274), .A2(n5949), .B1(n6284), .B2(n5430), .C1(n5480), 
        .C2(n5456), .ZN(U2837) );
  OR2_X1 U6609 ( .A1(n5431), .A2(n5432), .ZN(n5433) );
  AND2_X1 U6610 ( .A1(n5434), .A2(n5433), .ZN(n5963) );
  INV_X1 U6611 ( .A(n5963), .ZN(n5483) );
  INV_X1 U6612 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5439) );
  AND2_X1 U6613 ( .A1(n5436), .A2(n5435), .ZN(n5438) );
  OR2_X1 U6614 ( .A1(n5438), .A2(n5437), .ZN(n5961) );
  OAI222_X1 U6615 ( .A1(n5483), .A2(n5456), .B1(n5439), .B2(n6284), .C1(n6274), 
        .C2(n5961), .ZN(U2838) );
  NOR2_X1 U6616 ( .A1(n5440), .A2(n5441), .ZN(n5442) );
  OR2_X1 U6617 ( .A1(n5431), .A2(n5442), .ZN(n5967) );
  MUX2_X1 U6618 ( .A(n5445), .B(n5444), .S(n5443), .Z(n5447) );
  XNOR2_X1 U6619 ( .A(n5447), .B(n5446), .ZN(n5966) );
  OAI222_X1 U6620 ( .A1(n5967), .A2(n5456), .B1(n5448), .B2(n6284), .C1(n6274), 
        .C2(n5966), .ZN(U2839) );
  AND2_X1 U6621 ( .A1(n5450), .A2(n5449), .ZN(n5451) );
  NOR2_X1 U6622 ( .A1(n5440), .A2(n5451), .ZN(n5996) );
  INV_X1 U6623 ( .A(n5996), .ZN(n5488) );
  INV_X1 U6624 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5455) );
  INV_X1 U6625 ( .A(n5452), .ZN(n5453) );
  XNOR2_X1 U6626 ( .A(n5454), .B(n5453), .ZN(n5988) );
  OAI222_X1 U6627 ( .A1(n5456), .A2(n5488), .B1(n6284), .B2(n5455), .C1(n6274), 
        .C2(n5988), .ZN(U2840) );
  AOI22_X1 U6628 ( .A1(n6289), .A2(DATAI_30_), .B1(n6291), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U6629 ( .A1(n6292), .A2(DATAI_14_), .ZN(n5457) );
  OAI211_X1 U6630 ( .C1(n5350), .C2(n6285), .A(n5458), .B(n5457), .ZN(U2861)
         );
  AOI22_X1 U6631 ( .A1(n6289), .A2(DATAI_29_), .B1(n6291), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5460) );
  NAND2_X1 U6632 ( .A1(n6292), .A2(DATAI_13_), .ZN(n5459) );
  OAI211_X1 U6633 ( .C1(n5461), .C2(n6285), .A(n5460), .B(n5459), .ZN(U2862)
         );
  AOI22_X1 U6634 ( .A1(n6289), .A2(DATAI_28_), .B1(n6291), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5463) );
  NAND2_X1 U6635 ( .A1(n6292), .A2(DATAI_12_), .ZN(n5462) );
  OAI211_X1 U6636 ( .C1(n5464), .C2(n6285), .A(n5463), .B(n5462), .ZN(U2863)
         );
  AOI22_X1 U6637 ( .A1(n6289), .A2(DATAI_27_), .B1(n6291), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5466) );
  NAND2_X1 U6638 ( .A1(n6292), .A2(DATAI_11_), .ZN(n5465) );
  OAI211_X1 U6639 ( .C1(n5900), .C2(n6285), .A(n5466), .B(n5465), .ZN(U2864)
         );
  AOI22_X1 U6640 ( .A1(n6289), .A2(DATAI_26_), .B1(n6291), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5468) );
  NAND2_X1 U6641 ( .A1(n6292), .A2(DATAI_10_), .ZN(n5467) );
  OAI211_X1 U6642 ( .C1(n5909), .C2(n6285), .A(n5468), .B(n5467), .ZN(U2865)
         );
  AOI22_X1 U6643 ( .A1(n6289), .A2(DATAI_25_), .B1(n6291), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U6644 ( .A1(n6292), .A2(DATAI_9_), .ZN(n5469) );
  OAI211_X1 U6645 ( .C1(n5471), .C2(n6285), .A(n5470), .B(n5469), .ZN(U2866)
         );
  AOI22_X1 U6646 ( .A1(n6289), .A2(DATAI_24_), .B1(n6291), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5473) );
  NAND2_X1 U6647 ( .A1(n6292), .A2(DATAI_8_), .ZN(n5472) );
  OAI211_X1 U6648 ( .C1(n5474), .C2(n6285), .A(n5473), .B(n5472), .ZN(U2867)
         );
  AOI22_X1 U6649 ( .A1(n6289), .A2(DATAI_23_), .B1(n6291), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5476) );
  NAND2_X1 U6650 ( .A1(n6292), .A2(DATAI_7_), .ZN(n5475) );
  OAI211_X1 U6651 ( .C1(n5477), .C2(n6285), .A(n5476), .B(n5475), .ZN(U2868)
         );
  AOI22_X1 U6652 ( .A1(n6289), .A2(DATAI_22_), .B1(n6291), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5479) );
  NAND2_X1 U6653 ( .A1(n6292), .A2(DATAI_6_), .ZN(n5478) );
  OAI211_X1 U6654 ( .C1(n5480), .C2(n6285), .A(n5479), .B(n5478), .ZN(U2869)
         );
  AOI22_X1 U6655 ( .A1(n6289), .A2(DATAI_21_), .B1(n6291), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5482) );
  NAND2_X1 U6656 ( .A1(n6292), .A2(DATAI_5_), .ZN(n5481) );
  OAI211_X1 U6657 ( .C1(n5483), .C2(n6285), .A(n5482), .B(n5481), .ZN(U2870)
         );
  AOI22_X1 U6658 ( .A1(n6289), .A2(DATAI_20_), .B1(n6291), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5485) );
  NAND2_X1 U6659 ( .A1(n6292), .A2(DATAI_4_), .ZN(n5484) );
  OAI211_X1 U6660 ( .C1(n5967), .C2(n6285), .A(n5485), .B(n5484), .ZN(U2871)
         );
  AOI22_X1 U6661 ( .A1(n6289), .A2(DATAI_19_), .B1(n6291), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5487) );
  NAND2_X1 U6662 ( .A1(n6292), .A2(DATAI_3_), .ZN(n5486) );
  OAI211_X1 U6663 ( .C1(n5488), .C2(n6285), .A(n5487), .B(n5486), .ZN(U2872)
         );
  NAND2_X1 U6664 ( .A1(n3126), .A2(n5489), .ZN(n5491) );
  XNOR2_X1 U6665 ( .A(n5491), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5621)
         );
  NOR2_X1 U6666 ( .A1(n6187), .A2(n5492), .ZN(n5614) );
  AOI21_X1 U6667 ( .B1(n6341), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5614), 
        .ZN(n5493) );
  OAI21_X1 U6668 ( .B1(n6335), .B2(n5494), .A(n5493), .ZN(n5495) );
  AOI21_X1 U6669 ( .B1(n5496), .B2(n6329), .A(n5495), .ZN(n5497) );
  OAI21_X1 U6670 ( .B1(n5621), .B2(n6073), .A(n5497), .ZN(U2957) );
  INV_X1 U6672 ( .A(n5990), .ZN(n5499) );
  INV_X1 U6673 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5633) );
  AOI22_X1 U6674 ( .A1(n5506), .A2(n5633), .B1(n5505), .B2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5500) );
  INV_X1 U6675 ( .A(n5887), .ZN(n5502) );
  INV_X1 U6676 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6859) );
  NOR2_X1 U6677 ( .A1(n6187), .A2(n6859), .ZN(n5626) );
  AOI21_X1 U6678 ( .B1(n6341), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5626), 
        .ZN(n5501) );
  OAI21_X1 U6679 ( .B1(n6335), .B2(n5502), .A(n5501), .ZN(n5503) );
  AOI21_X1 U6680 ( .B1(n5890), .B2(n6329), .A(n5503), .ZN(n5504) );
  OAI21_X1 U6681 ( .B1(n3136), .B2(n6073), .A(n5504), .ZN(U2958) );
  NOR2_X1 U6682 ( .A1(n5506), .A2(n5505), .ZN(n5507) );
  XNOR2_X1 U6683 ( .A(n5507), .B(n5633), .ZN(n5638) );
  INV_X1 U6684 ( .A(n5900), .ZN(n5510) );
  INV_X1 U6685 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6949) );
  NOR2_X1 U6686 ( .A1(n6187), .A2(n6949), .ZN(n5632) );
  AOI21_X1 U6687 ( .B1(n6341), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5632), 
        .ZN(n5508) );
  OAI21_X1 U6688 ( .B1(n6335), .B2(n5896), .A(n5508), .ZN(n5509) );
  AOI21_X1 U6689 ( .B1(n5510), .B2(n6329), .A(n5509), .ZN(n5511) );
  OAI21_X1 U6690 ( .B1(n5638), .B2(n6073), .A(n5511), .ZN(U2959) );
  XNOR2_X1 U6691 ( .A(n3119), .B(n5512), .ZN(n5513) );
  XNOR2_X1 U6692 ( .A(n5514), .B(n5513), .ZN(n5645) );
  INV_X1 U6693 ( .A(n5909), .ZN(n5518) );
  INV_X1 U6694 ( .A(n5912), .ZN(n5516) );
  INV_X1 U6695 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6869) );
  NOR2_X1 U6696 ( .A1(n6187), .A2(n6869), .ZN(n5640) );
  AOI21_X1 U6697 ( .B1(n6341), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5640), 
        .ZN(n5515) );
  OAI21_X1 U6698 ( .B1(n6335), .B2(n5516), .A(n5515), .ZN(n5517) );
  AOI21_X1 U6699 ( .B1(n5518), .B2(n6329), .A(n5517), .ZN(n5519) );
  OAI21_X1 U6700 ( .B1(n6073), .B2(n5645), .A(n5519), .ZN(U2960) );
  OAI21_X1 U6701 ( .B1(n5521), .B2(n6854), .A(n3119), .ZN(n5522) );
  XNOR2_X1 U6702 ( .A(n3552), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5551)
         );
  NOR2_X1 U6703 ( .A1(n3119), .A2(n6799), .ZN(n5523) );
  XNOR2_X1 U6704 ( .A(n3552), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5546)
         );
  NOR2_X1 U6705 ( .A1(n3119), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5537)
         );
  NAND2_X1 U6706 ( .A1(n5524), .A2(n5537), .ZN(n5532) );
  OAI21_X1 U6707 ( .B1(n3556), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5544), 
        .ZN(n5539) );
  NAND3_X1 U6708 ( .A1(n3119), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5525) );
  XNOR2_X1 U6709 ( .A(n5526), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5654)
         );
  INV_X1 U6710 ( .A(REIP_REG_24__SCAN_IN), .ZN(n5527) );
  NOR2_X1 U6711 ( .A1(n6187), .A2(n5527), .ZN(n5651) );
  AOI21_X1 U6712 ( .B1(n6341), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5651), 
        .ZN(n5528) );
  OAI21_X1 U6713 ( .B1(n6335), .B2(n5928), .A(n5528), .ZN(n5529) );
  AOI21_X1 U6714 ( .B1(n5930), .B2(n6329), .A(n5529), .ZN(n5530) );
  OAI21_X1 U6715 ( .B1(n5654), .B2(n6073), .A(n5530), .ZN(U2962) );
  NAND4_X1 U6716 ( .A1(n5552), .A2(n5647), .A3(INSTADDRPOINTER_REG_20__SCAN_IN), .A4(n3119), .ZN(n5531) );
  NAND2_X1 U6717 ( .A1(n5532), .A2(n5531), .ZN(n5533) );
  XNOR2_X1 U6718 ( .A(n5533), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5662)
         );
  NAND2_X1 U6719 ( .A1(n6395), .A2(REIP_REG_23__SCAN_IN), .ZN(n5655) );
  NAND2_X1 U6720 ( .A1(n6341), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5534)
         );
  OAI211_X1 U6721 ( .C1(n6335), .C2(n5945), .A(n5655), .B(n5534), .ZN(n5535)
         );
  AOI21_X1 U6722 ( .B1(n5942), .B2(n6329), .A(n5535), .ZN(n5536) );
  OAI21_X1 U6723 ( .B1(n5662), .B2(n6073), .A(n5536), .ZN(U2963) );
  AOI21_X1 U6724 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n3119), .A(n5537), 
        .ZN(n5538) );
  XNOR2_X1 U6725 ( .A(n5539), .B(n5538), .ZN(n5670) );
  NAND2_X1 U6726 ( .A1(n5593), .A2(n5946), .ZN(n5540) );
  NAND2_X1 U6727 ( .A1(n6395), .A2(REIP_REG_22__SCAN_IN), .ZN(n5667) );
  OAI211_X1 U6728 ( .C1(n5591), .C2(n5541), .A(n5540), .B(n5667), .ZN(n5542)
         );
  AOI21_X1 U6729 ( .B1(n5951), .B2(n6329), .A(n5542), .ZN(n5543) );
  OAI21_X1 U6730 ( .B1(n5670), .B2(n6073), .A(n5543), .ZN(U2964) );
  OAI21_X1 U6731 ( .B1(n5546), .B2(n5545), .A(n5544), .ZN(n5547) );
  INV_X1 U6732 ( .A(n5547), .ZN(n5678) );
  NAND2_X1 U6733 ( .A1(n6395), .A2(REIP_REG_21__SCAN_IN), .ZN(n5674) );
  NAND2_X1 U6734 ( .A1(n6341), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5548)
         );
  OAI211_X1 U6735 ( .C1(n6335), .C2(n5958), .A(n5674), .B(n5548), .ZN(n5549)
         );
  AOI21_X1 U6736 ( .B1(n5963), .B2(n6329), .A(n5549), .ZN(n5550) );
  OAI21_X1 U6737 ( .B1(n5678), .B2(n6073), .A(n5550), .ZN(U2965) );
  XNOR2_X1 U6738 ( .A(n5552), .B(n5551), .ZN(n5688) );
  INV_X1 U6739 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5553) );
  NAND2_X1 U6740 ( .A1(n6395), .A2(REIP_REG_20__SCAN_IN), .ZN(n5685) );
  OAI21_X1 U6741 ( .B1(n5591), .B2(n5553), .A(n5685), .ZN(n5555) );
  NOR2_X1 U6742 ( .A1(n5967), .A2(n6344), .ZN(n5554) );
  AOI211_X1 U6743 ( .C1(n5593), .C2(n5972), .A(n5555), .B(n5554), .ZN(n5556)
         );
  OAI21_X1 U6744 ( .B1(n6073), .B2(n5688), .A(n5556), .ZN(U2966) );
  NAND2_X1 U6745 ( .A1(n3552), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6006) );
  NAND2_X1 U6746 ( .A1(n5596), .A2(n5559), .ZN(n5577) );
  NAND2_X1 U6747 ( .A1(n5577), .A2(n5560), .ZN(n5578) );
  INV_X1 U6748 ( .A(n5578), .ZN(n5561) );
  INV_X1 U6749 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6035) );
  NAND4_X1 U6750 ( .A1(n5561), .A2(n3556), .A3(n5703), .A4(n6035), .ZN(n6004)
         );
  OAI21_X1 U6751 ( .B1(n6002), .B2(n6006), .A(n6004), .ZN(n5562) );
  XOR2_X1 U6752 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n5562), .Z(n6025) );
  NAND2_X1 U6753 ( .A1(n6025), .A2(n6339), .ZN(n5567) );
  OAI22_X1 U6754 ( .A1(n5591), .A2(n5563), .B1(n6187), .B2(n6979), .ZN(n5564)
         );
  AOI21_X1 U6755 ( .B1(n5593), .B2(n5565), .A(n5564), .ZN(n5566) );
  OAI211_X1 U6756 ( .C1(n6344), .C2(n5568), .A(n5567), .B(n5566), .ZN(U2968)
         );
  INV_X1 U6757 ( .A(n6001), .ZN(n5570) );
  NOR2_X1 U6758 ( .A1(n5570), .A2(n5569), .ZN(n5572) );
  XOR2_X1 U6759 ( .A(n5572), .B(n5571), .Z(n5708) );
  NAND2_X1 U6760 ( .A1(n6395), .A2(REIP_REG_16__SCAN_IN), .ZN(n5701) );
  NAND2_X1 U6761 ( .A1(n6341), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5573)
         );
  OAI211_X1 U6762 ( .C1(n6335), .C2(n6106), .A(n5701), .B(n5573), .ZN(n5574)
         );
  AOI21_X1 U6763 ( .B1(n6290), .B2(n6329), .A(n5574), .ZN(n5575) );
  OAI21_X1 U6764 ( .B1(n5708), .B2(n6073), .A(n5575), .ZN(U2970) );
  AND2_X1 U6765 ( .A1(n5577), .A2(n5576), .ZN(n5580) );
  OAI21_X1 U6766 ( .B1(n5580), .B2(n5579), .A(n5578), .ZN(n6042) );
  NAND2_X1 U6767 ( .A1(n6042), .A2(n6339), .ZN(n5584) );
  OAI22_X1 U6768 ( .A1(n5591), .A2(n6977), .B1(n6187), .B2(n6634), .ZN(n5581)
         );
  AOI21_X1 U6769 ( .B1(n5593), .B2(n5582), .A(n5581), .ZN(n5583) );
  OAI211_X1 U6770 ( .C1(n6344), .C2(n5585), .A(n5584), .B(n5583), .ZN(U2971)
         );
  NAND2_X1 U6771 ( .A1(n5596), .A2(n5586), .ZN(n5588) );
  XNOR2_X1 U6772 ( .A(n3119), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5587)
         );
  XNOR2_X1 U6773 ( .A(n5588), .B(n5587), .ZN(n6053) );
  NAND2_X1 U6774 ( .A1(n6053), .A2(n6339), .ZN(n5595) );
  INV_X1 U6775 ( .A(REIP_REG_14__SCAN_IN), .ZN(n5589) );
  OAI22_X1 U6776 ( .A1(n5591), .A2(n5590), .B1(n6187), .B2(n5589), .ZN(n5592)
         );
  AOI21_X1 U6777 ( .B1(n5593), .B2(n6115), .A(n5592), .ZN(n5594) );
  OAI211_X1 U6778 ( .C1(n6344), .C2(n6113), .A(n5595), .B(n5594), .ZN(U2972)
         );
  INV_X1 U6779 ( .A(n5596), .ZN(n5597) );
  AOI21_X1 U6780 ( .B1(n5598), .B2(n5558), .A(n5597), .ZN(n5721) );
  XNOR2_X1 U6781 ( .A(n5599), .B(n3147), .ZN(n6297) );
  NOR2_X1 U6782 ( .A1(n6187), .A2(n5257), .ZN(n5718) );
  AOI21_X1 U6783 ( .B1(n6341), .B2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n5718), 
        .ZN(n5600) );
  OAI21_X1 U6784 ( .B1(n6335), .B2(n6124), .A(n5600), .ZN(n5601) );
  AOI21_X1 U6785 ( .B1(n6297), .B2(n6329), .A(n5601), .ZN(n5602) );
  OAI21_X1 U6786 ( .B1(n5721), .B2(n6073), .A(n5602), .ZN(U2973) );
  OAI21_X1 U6787 ( .B1(n5604), .B2(n5680), .A(n5612), .ZN(n5610) );
  NOR3_X1 U6788 ( .A1(n5617), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5605), 
        .ZN(n5609) );
  OAI21_X1 U6789 ( .B1(n5607), .B2(n6394), .A(n5606), .ZN(n5608) );
  OAI21_X1 U6790 ( .B1(n5603), .B2(n6399), .A(n5611), .ZN(U2987) );
  INV_X1 U6791 ( .A(n5612), .ZN(n5619) );
  INV_X1 U6792 ( .A(n5613), .ZN(n5615) );
  AOI21_X1 U6793 ( .B1(n5615), .B2(n6375), .A(n5614), .ZN(n5616) );
  OAI21_X1 U6794 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5617), .A(n5616), 
        .ZN(n5618) );
  AOI21_X1 U6795 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5619), .A(n5618), 
        .ZN(n5620) );
  OAI21_X1 U6796 ( .B1(n5621), .B2(n6399), .A(n5620), .ZN(U2989) );
  INV_X1 U6797 ( .A(n5888), .ZN(n5627) );
  INV_X1 U6798 ( .A(n5634), .ZN(n5624) );
  NOR3_X1 U6799 ( .A1(n5624), .A2(n5623), .A3(n5622), .ZN(n5625) );
  AOI211_X1 U6800 ( .C1(n6375), .C2(n5627), .A(n5626), .B(n5625), .ZN(n5630)
         );
  OAI21_X1 U6801 ( .B1(n5680), .B2(n5628), .A(n6021), .ZN(n5635) );
  NAND2_X1 U6802 ( .A1(n5635), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5629) );
  OAI211_X1 U6803 ( .C1(n3136), .C2(n6399), .A(n5630), .B(n5629), .ZN(U2990)
         );
  NOR2_X1 U6804 ( .A1(n5899), .A2(n6394), .ZN(n5631) );
  AOI211_X1 U6805 ( .C1(n5634), .C2(n5633), .A(n5632), .B(n5631), .ZN(n5637)
         );
  NAND2_X1 U6806 ( .A1(n5635), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5636) );
  OAI211_X1 U6807 ( .C1(n5638), .C2(n6399), .A(n5637), .B(n5636), .ZN(U2991)
         );
  XNOR2_X1 U6808 ( .A(n6020), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5641)
         );
  NOR2_X1 U6809 ( .A1(n5914), .A2(n6394), .ZN(n5639) );
  AOI211_X1 U6810 ( .C1(n5641), .C2(n6014), .A(n5640), .B(n5639), .ZN(n5644)
         );
  NAND2_X1 U6811 ( .A1(n5642), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5643) );
  OAI211_X1 U6812 ( .C1(n5645), .C2(n6399), .A(n5644), .B(n5643), .ZN(U2992)
         );
  INV_X1 U6813 ( .A(n5935), .ZN(n5652) );
  INV_X1 U6814 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5649) );
  NOR2_X1 U6815 ( .A1(n5646), .A2(n6022), .ZN(n5671) );
  NAND2_X1 U6816 ( .A1(n5647), .A2(n5671), .ZN(n5656) );
  AOI211_X1 U6817 ( .C1(n5649), .C2(n5656), .A(n5648), .B(n6021), .ZN(n5650)
         );
  AOI211_X1 U6818 ( .C1(n6375), .C2(n5652), .A(n5651), .B(n5650), .ZN(n5653)
         );
  OAI21_X1 U6819 ( .B1(n5654), .B2(n6399), .A(n5653), .ZN(U2994) );
  OAI21_X1 U6820 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5656), .A(n5655), 
        .ZN(n5660) );
  INV_X1 U6821 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5657) );
  NOR2_X1 U6822 ( .A1(n5658), .A2(n5657), .ZN(n5659) );
  AOI211_X1 U6823 ( .C1(n6375), .C2(n5937), .A(n5660), .B(n5659), .ZN(n5661)
         );
  OAI21_X1 U6824 ( .B1(n5662), .B2(n6399), .A(n5661), .ZN(U2995) );
  INV_X1 U6825 ( .A(n5663), .ZN(n5665) );
  NAND3_X1 U6826 ( .A1(n5665), .A2(n5671), .A3(n5664), .ZN(n5666) );
  OAI211_X1 U6827 ( .C1(n5949), .C2(n6394), .A(n5667), .B(n5666), .ZN(n5668)
         );
  AOI21_X1 U6828 ( .B1(n5676), .B2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5668), 
        .ZN(n5669) );
  OAI21_X1 U6829 ( .B1(n5670), .B2(n6399), .A(n5669), .ZN(U2996) );
  INV_X1 U6830 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5672) );
  NAND2_X1 U6831 ( .A1(n5672), .A2(n5671), .ZN(n5673) );
  OAI211_X1 U6832 ( .C1(n5961), .C2(n6394), .A(n5674), .B(n5673), .ZN(n5675)
         );
  AOI21_X1 U6833 ( .B1(n5676), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5675), 
        .ZN(n5677) );
  OAI21_X1 U6834 ( .B1(n5678), .B2(n6399), .A(n5677), .ZN(U2997) );
  AOI21_X1 U6835 ( .B1(n6035), .B2(n5679), .A(n6037), .ZN(n6028) );
  OAI21_X1 U6836 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5680), .A(n6028), 
        .ZN(n5695) );
  INV_X1 U6837 ( .A(n5681), .ZN(n5683) );
  AOI21_X1 U6838 ( .B1(n6854), .B2(n6799), .A(n5692), .ZN(n5682) );
  NAND2_X1 U6839 ( .A1(n5683), .A2(n5682), .ZN(n5684) );
  OAI211_X1 U6840 ( .C1(n5966), .C2(n6394), .A(n5685), .B(n5684), .ZN(n5686)
         );
  AOI21_X1 U6841 ( .B1(n5695), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5686), 
        .ZN(n5687) );
  OAI21_X1 U6842 ( .B1(n5688), .B2(n6399), .A(n5687), .ZN(U2998) );
  OAI21_X1 U6843 ( .B1(n3127), .B2(n6854), .A(n5520), .ZN(n5690) );
  XNOR2_X1 U6844 ( .A(n5690), .B(n3556), .ZN(n5997) );
  INV_X1 U6845 ( .A(n5997), .ZN(n5697) );
  INV_X1 U6846 ( .A(REIP_REG_19__SCAN_IN), .ZN(n5691) );
  OAI22_X1 U6847 ( .A1(n5988), .A2(n6394), .B1(n6187), .B2(n5691), .ZN(n5694)
         );
  NOR2_X1 U6848 ( .A1(n5692), .A2(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5693)
         );
  AOI211_X1 U6849 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5695), .A(n5694), .B(n5693), .ZN(n5696) );
  OAI21_X1 U6850 ( .B1(n5697), .B2(n6399), .A(n5696), .ZN(U2999) );
  AOI21_X1 U6851 ( .B1(n6389), .B2(n5699), .A(n5698), .ZN(n5700) );
  INV_X1 U6852 ( .A(n5700), .ZN(n6040) );
  OAI21_X1 U6853 ( .B1(n6110), .B2(n6394), .A(n5701), .ZN(n5702) );
  AOI21_X1 U6854 ( .B1(n6040), .B2(INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5702), 
        .ZN(n5707) );
  NAND3_X1 U6855 ( .A1(n6046), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n6348), .ZN(n6045) );
  AOI21_X1 U6856 ( .B1(n6921), .B2(n5703), .A(n6045), .ZN(n5705) );
  NAND2_X1 U6857 ( .A1(n5705), .A2(n5704), .ZN(n5706) );
  OAI211_X1 U6858 ( .C1(n5708), .C2(n6399), .A(n5707), .B(n5706), .ZN(U3002)
         );
  NAND2_X1 U6859 ( .A1(n6392), .A2(n5711), .ZN(n5709) );
  OAI211_X1 U6860 ( .C1(n6046), .C2(n5710), .A(n6352), .B(n5709), .ZN(n6048)
         );
  NOR2_X1 U6861 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5711), .ZN(n6050)
         );
  AOI22_X1 U6862 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n6048), .B1(n6050), .B2(n6348), .ZN(n5720) );
  INV_X1 U6863 ( .A(n5712), .ZN(n5715) );
  AOI21_X1 U6864 ( .B1(n5715), .B2(n5714), .A(n5713), .ZN(n5717) );
  OR2_X1 U6865 ( .A1(n5717), .A2(n5716), .ZN(n6273) );
  INV_X1 U6866 ( .A(n6273), .ZN(n6123) );
  AOI21_X1 U6867 ( .B1(n6375), .B2(n6123), .A(n5718), .ZN(n5719) );
  OAI211_X1 U6868 ( .C1(n5721), .C2(n6399), .A(n5720), .B(n5719), .ZN(U3005)
         );
  OAI211_X1 U6869 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5722), .A(n6472), .B(
        n6471), .ZN(n5723) );
  OAI21_X1 U6870 ( .B1(n5726), .B2(n4563), .A(n5723), .ZN(n5724) );
  MUX2_X1 U6871 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5724), .S(n6404), 
        .Z(U3464) );
  XNOR2_X1 U6872 ( .A(n5725), .B(n6472), .ZN(n5728) );
  INV_X1 U6873 ( .A(n6246), .ZN(n5727) );
  OAI22_X1 U6874 ( .A1(n5728), .A2(n6477), .B1(n5727), .B2(n5726), .ZN(n5729)
         );
  MUX2_X1 U6875 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5729), .S(n6404), 
        .Z(U3463) );
  INV_X1 U6876 ( .A(n5782), .ZN(n5730) );
  NOR2_X1 U6877 ( .A1(n5731), .A2(n5730), .ZN(n5738) );
  AOI22_X1 U6878 ( .A1(n5738), .A2(n6471), .B1(n6406), .B2(n5732), .ZN(n5769)
         );
  NOR2_X1 U6879 ( .A1(n6563), .A2(n5788), .ZN(n5781) );
  NAND2_X1 U6880 ( .A1(n6411), .A2(n5781), .ZN(n5779) );
  INV_X1 U6881 ( .A(n5779), .ZN(n5766) );
  NAND2_X1 U6882 ( .A1(n5736), .A2(n5735), .ZN(n5812) );
  AOI21_X1 U6883 ( .B1(n5812), .B2(n6524), .A(n6072), .ZN(n5737) );
  NOR3_X1 U6884 ( .A1(n5738), .A2(n5737), .A3(n6477), .ZN(n5741) );
  INV_X1 U6885 ( .A(n5739), .ZN(n5740) );
  AOI211_X1 U6886 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n5779), .A(n5741), .B(
        n5740), .ZN(n5743) );
  NAND2_X1 U6887 ( .A1(n5743), .A2(n5742), .ZN(n5774) );
  AOI22_X1 U6888 ( .A1(n5822), .A2(n6469), .B1(INSTQUEUE_REG_12__0__SCAN_IN), 
        .B2(n5774), .ZN(n5744) );
  OAI21_X1 U6889 ( .B1(n6487), .B2(n6524), .A(n5744), .ZN(n5745) );
  AOI21_X1 U6890 ( .B1(n6470), .B2(n5766), .A(n5745), .ZN(n5746) );
  OAI21_X1 U6891 ( .B1(n5747), .B2(n5769), .A(n5746), .ZN(U3116) );
  AOI22_X1 U6892 ( .A1(n5822), .A2(n5844), .B1(INSTQUEUE_REG_12__1__SCAN_IN), 
        .B2(n5774), .ZN(n5748) );
  OAI21_X1 U6893 ( .B1(n5794), .B2(n6524), .A(n5748), .ZN(n5749) );
  AOI21_X1 U6894 ( .B1(n6489), .B2(n5766), .A(n5749), .ZN(n5750) );
  OAI21_X1 U6895 ( .B1(n5751), .B2(n5769), .A(n5750), .ZN(U3117) );
  AOI22_X1 U6896 ( .A1(n5822), .A2(n6494), .B1(INSTQUEUE_REG_12__2__SCAN_IN), 
        .B2(n5774), .ZN(n5752) );
  OAI21_X1 U6897 ( .B1(n6499), .B2(n6524), .A(n5752), .ZN(n5753) );
  AOI21_X1 U6898 ( .B1(n6495), .B2(n5766), .A(n5753), .ZN(n5754) );
  OAI21_X1 U6899 ( .B1(n5755), .B2(n5769), .A(n5754), .ZN(U3118) );
  AOI22_X1 U6900 ( .A1(n5822), .A2(n6500), .B1(INSTQUEUE_REG_12__3__SCAN_IN), 
        .B2(n5774), .ZN(n5756) );
  OAI21_X1 U6901 ( .B1(n6505), .B2(n6524), .A(n5756), .ZN(n5757) );
  AOI21_X1 U6902 ( .B1(n6501), .B2(n5766), .A(n5757), .ZN(n5758) );
  OAI21_X1 U6903 ( .B1(n5759), .B2(n5769), .A(n5758), .ZN(U3119) );
  AOI22_X1 U6904 ( .A1(n5822), .A2(n5860), .B1(INSTQUEUE_REG_12__4__SCAN_IN), 
        .B2(n5774), .ZN(n5760) );
  OAI21_X1 U6905 ( .B1(n5807), .B2(n6524), .A(n5760), .ZN(n5761) );
  AOI21_X1 U6906 ( .B1(n6507), .B2(n5766), .A(n5761), .ZN(n5762) );
  OAI21_X1 U6907 ( .B1(n5763), .B2(n5769), .A(n5762), .ZN(U3120) );
  AOI22_X1 U6908 ( .A1(n5822), .A2(n6455), .B1(INSTQUEUE_REG_12__5__SCAN_IN), 
        .B2(n5774), .ZN(n5764) );
  OAI21_X1 U6909 ( .B1(n6458), .B2(n6524), .A(n5764), .ZN(n5765) );
  AOI21_X1 U6910 ( .B1(n6513), .B2(n5766), .A(n5765), .ZN(n5767) );
  OAI21_X1 U6911 ( .B1(n5768), .B2(n5769), .A(n5767), .ZN(U3121) );
  INV_X1 U6912 ( .A(n6524), .ZN(n6526) );
  INV_X1 U6913 ( .A(n5769), .ZN(n5775) );
  AOI22_X1 U6914 ( .A1(n5775), .A2(n6521), .B1(INSTQUEUE_REG_12__6__SCAN_IN), 
        .B2(n5774), .ZN(n5770) );
  OAI21_X1 U6915 ( .B1(n5812), .B2(n6525), .A(n5770), .ZN(n5771) );
  AOI21_X1 U6916 ( .B1(n6519), .B2(n6526), .A(n5771), .ZN(n5772) );
  OAI21_X1 U6917 ( .B1(n5773), .B2(n5779), .A(n5772), .ZN(U3122) );
  AOI22_X1 U6918 ( .A1(n5775), .A2(n6531), .B1(INSTQUEUE_REG_12__7__SCAN_IN), 
        .B2(n5774), .ZN(n5776) );
  OAI21_X1 U6919 ( .B1(n5812), .B2(n6448), .A(n5776), .ZN(n5777) );
  AOI21_X1 U6920 ( .B1(n6444), .B2(n6526), .A(n5777), .ZN(n5778) );
  OAI21_X1 U6921 ( .B1(n5780), .B2(n5779), .A(n5778), .ZN(U3123) );
  INV_X1 U6922 ( .A(n5781), .ZN(n5786) );
  AND2_X1 U6923 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5781), .ZN(n5826)
         );
  AOI21_X1 U6924 ( .B1(n5831), .B2(n5782), .A(n5826), .ZN(n5790) );
  NAND2_X1 U6925 ( .A1(n5790), .A2(n5783), .ZN(n5784) );
  NOR2_X1 U6926 ( .A1(n6477), .A2(n5784), .ZN(n5785) );
  INV_X1 U6927 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n5793) );
  OAI22_X1 U6928 ( .A1(n6424), .A2(n5824), .B1(n5812), .B2(n6487), .ZN(n5787)
         );
  AOI21_X1 U6929 ( .B1(n6470), .B2(n5826), .A(n5787), .ZN(n5792) );
  NAND2_X1 U6930 ( .A1(STATE2_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n5789) );
  OAI22_X1 U6931 ( .A1(n5790), .A2(n6477), .B1(n5789), .B2(n5788), .ZN(n5821)
         );
  NAND2_X1 U6932 ( .A1(n6484), .A2(n5821), .ZN(n5791) );
  OAI211_X1 U6933 ( .C1(n5829), .C2(n5793), .A(n5792), .B(n5791), .ZN(U3124)
         );
  INV_X1 U6934 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n5798) );
  OAI22_X1 U6935 ( .A1(n6493), .A2(n5824), .B1(n5812), .B2(n5794), .ZN(n5795)
         );
  AOI21_X1 U6936 ( .B1(n6489), .B2(n5826), .A(n5795), .ZN(n5797) );
  NAND2_X1 U6937 ( .A1(n6490), .A2(n5821), .ZN(n5796) );
  OAI211_X1 U6938 ( .C1(n5829), .C2(n5798), .A(n5797), .B(n5796), .ZN(U3125)
         );
  INV_X1 U6939 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n5802) );
  OAI22_X1 U6940 ( .A1(n6430), .A2(n5824), .B1(n5812), .B2(n6499), .ZN(n5799)
         );
  AOI21_X1 U6941 ( .B1(n6495), .B2(n5826), .A(n5799), .ZN(n5801) );
  NAND2_X1 U6942 ( .A1(n6496), .A2(n5821), .ZN(n5800) );
  OAI211_X1 U6943 ( .C1(n5829), .C2(n5802), .A(n5801), .B(n5800), .ZN(U3126)
         );
  INV_X1 U6944 ( .A(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n5806) );
  OAI22_X1 U6945 ( .A1(n6434), .A2(n5824), .B1(n5812), .B2(n6505), .ZN(n5803)
         );
  AOI21_X1 U6946 ( .B1(n6501), .B2(n5826), .A(n5803), .ZN(n5805) );
  NAND2_X1 U6947 ( .A1(n6502), .A2(n5821), .ZN(n5804) );
  OAI211_X1 U6948 ( .C1(n5829), .C2(n5806), .A(n5805), .B(n5804), .ZN(U3127)
         );
  INV_X1 U6949 ( .A(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n5811) );
  OAI22_X1 U6950 ( .A1(n6511), .A2(n5824), .B1(n5812), .B2(n5807), .ZN(n5808)
         );
  AOI21_X1 U6951 ( .B1(n6507), .B2(n5826), .A(n5808), .ZN(n5810) );
  NAND2_X1 U6952 ( .A1(n6508), .A2(n5821), .ZN(n5809) );
  OAI211_X1 U6953 ( .C1(n5829), .C2(n5811), .A(n5810), .B(n5809), .ZN(U3128)
         );
  INV_X1 U6954 ( .A(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n5816) );
  OAI22_X1 U6955 ( .A1(n6517), .A2(n5824), .B1(n5812), .B2(n6458), .ZN(n5813)
         );
  AOI21_X1 U6956 ( .B1(n6513), .B2(n5826), .A(n5813), .ZN(n5815) );
  NAND2_X1 U6957 ( .A1(n6514), .A2(n5821), .ZN(n5814) );
  OAI211_X1 U6958 ( .C1(n5829), .C2(n5816), .A(n5815), .B(n5814), .ZN(U3129)
         );
  INV_X1 U6959 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n5820) );
  AOI22_X1 U6960 ( .A1(n5822), .A2(n6519), .B1(n6521), .B2(n5821), .ZN(n5817)
         );
  OAI21_X1 U6961 ( .B1(n6525), .B2(n5824), .A(n5817), .ZN(n5818) );
  AOI21_X1 U6962 ( .B1(n6520), .B2(n5826), .A(n5818), .ZN(n5819) );
  OAI21_X1 U6963 ( .B1(n5829), .B2(n5820), .A(n5819), .ZN(U3130) );
  INV_X1 U6964 ( .A(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n5828) );
  AOI22_X1 U6965 ( .A1(n5822), .A2(n6444), .B1(n6531), .B2(n5821), .ZN(n5823)
         );
  OAI21_X1 U6966 ( .B1(n6448), .B2(n5824), .A(n5823), .ZN(n5825) );
  AOI21_X1 U6967 ( .B1(n6529), .B2(n5826), .A(n5825), .ZN(n5827) );
  OAI21_X1 U6968 ( .B1(n5829), .B2(n5828), .A(n5827), .ZN(U3131) );
  INV_X1 U6969 ( .A(n5868), .ZN(n5882) );
  AOI21_X1 U6970 ( .B1(n5831), .B2(n5830), .A(n5882), .ZN(n5838) );
  OAI21_X1 U6971 ( .B1(n5833), .B2(n6344), .A(n5832), .ZN(n5836) );
  NOR2_X1 U6972 ( .A1(n6471), .A2(n5834), .ZN(n5835) );
  AOI211_X2 U6973 ( .C1(n5838), .C2(n5836), .A(n5835), .B(n6476), .ZN(n5885)
         );
  INV_X1 U6974 ( .A(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n5843) );
  OAI22_X1 U6975 ( .A1(n5838), .A2(n6477), .B1(n6480), .B2(n5837), .ZN(n5877)
         );
  AOI22_X1 U6976 ( .A1(n6421), .A2(n5866), .B1(n5878), .B2(n6469), .ZN(n5839)
         );
  OAI21_X1 U6977 ( .B1(n5840), .B2(n5868), .A(n5839), .ZN(n5841) );
  AOI21_X1 U6978 ( .B1(n6484), .B2(n5877), .A(n5841), .ZN(n5842) );
  OAI21_X1 U6979 ( .B1(n5885), .B2(n5843), .A(n5842), .ZN(U3140) );
  INV_X1 U6980 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n5849) );
  AOI22_X1 U6981 ( .A1(n6488), .A2(n5866), .B1(n5878), .B2(n5844), .ZN(n5845)
         );
  OAI21_X1 U6982 ( .B1(n5846), .B2(n5868), .A(n5845), .ZN(n5847) );
  AOI21_X1 U6983 ( .B1(n6490), .B2(n5877), .A(n5847), .ZN(n5848) );
  OAI21_X1 U6984 ( .B1(n5885), .B2(n5849), .A(n5848), .ZN(U3141) );
  INV_X1 U6985 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n5854) );
  AOI22_X1 U6986 ( .A1(n6427), .A2(n5866), .B1(n5878), .B2(n6494), .ZN(n5850)
         );
  OAI21_X1 U6987 ( .B1(n5851), .B2(n5868), .A(n5850), .ZN(n5852) );
  AOI21_X1 U6988 ( .B1(n6496), .B2(n5877), .A(n5852), .ZN(n5853) );
  OAI21_X1 U6989 ( .B1(n5885), .B2(n5854), .A(n5853), .ZN(U3142) );
  INV_X1 U6990 ( .A(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n5859) );
  AOI22_X1 U6991 ( .A1(n6431), .A2(n5866), .B1(n5878), .B2(n6500), .ZN(n5855)
         );
  OAI21_X1 U6992 ( .B1(n5856), .B2(n5868), .A(n5855), .ZN(n5857) );
  AOI21_X1 U6993 ( .B1(n6502), .B2(n5877), .A(n5857), .ZN(n5858) );
  OAI21_X1 U6994 ( .B1(n5885), .B2(n5859), .A(n5858), .ZN(U3143) );
  INV_X1 U6995 ( .A(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n5865) );
  AOI22_X1 U6996 ( .A1(n6506), .A2(n5866), .B1(n5878), .B2(n5860), .ZN(n5861)
         );
  OAI21_X1 U6997 ( .B1(n5862), .B2(n5868), .A(n5861), .ZN(n5863) );
  AOI21_X1 U6998 ( .B1(n6508), .B2(n5877), .A(n5863), .ZN(n5864) );
  OAI21_X1 U6999 ( .B1(n5885), .B2(n5865), .A(n5864), .ZN(U3144) );
  INV_X1 U7000 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n5872) );
  AOI22_X1 U7001 ( .A1(n6512), .A2(n5866), .B1(n5878), .B2(n6455), .ZN(n5867)
         );
  OAI21_X1 U7002 ( .B1(n5869), .B2(n5868), .A(n5867), .ZN(n5870) );
  AOI21_X1 U7003 ( .B1(n6514), .B2(n5877), .A(n5870), .ZN(n5871) );
  OAI21_X1 U7004 ( .B1(n5885), .B2(n5872), .A(n5871), .ZN(U3145) );
  INV_X1 U7005 ( .A(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n5876) );
  AOI22_X1 U7006 ( .A1(n5878), .A2(n6460), .B1(n6521), .B2(n5877), .ZN(n5873)
         );
  OAI21_X1 U7007 ( .B1(n5880), .B2(n6467), .A(n5873), .ZN(n5874) );
  AOI21_X1 U7008 ( .B1(n6520), .B2(n5882), .A(n5874), .ZN(n5875) );
  OAI21_X1 U7009 ( .B1(n5885), .B2(n5876), .A(n5875), .ZN(U3146) );
  INV_X1 U7010 ( .A(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n5884) );
  AOI22_X1 U7011 ( .A1(n5878), .A2(n6527), .B1(n6531), .B2(n5877), .ZN(n5879)
         );
  OAI21_X1 U7012 ( .B1(n5880), .B2(n6536), .A(n5879), .ZN(n5881) );
  AOI21_X1 U7013 ( .B1(n6529), .B2(n5882), .A(n5881), .ZN(n5883) );
  OAI21_X1 U7014 ( .B1(n5885), .B2(n5884), .A(n5883), .ZN(U3147) );
  AND2_X1 U7015 ( .A1(n6323), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U7016 ( .A1(EBX_REG_28__SCAN_IN), .A2(n6261), .B1(
        PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n6245), .ZN(n5894) );
  AOI22_X1 U7017 ( .A1(n5887), .A2(n6258), .B1(REIP_REG_28__SCAN_IN), .B2(
        n5886), .ZN(n5893) );
  NOR2_X1 U7018 ( .A1(n5888), .A2(n6176), .ZN(n5889) );
  AOI21_X1 U7019 ( .B1(n5890), .B2(n6203), .A(n5889), .ZN(n5892) );
  NAND3_X1 U7020 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5898), .A3(n6859), .ZN(
        n5891) );
  NAND4_X1 U7021 ( .A1(n5894), .A2(n5893), .A3(n5892), .A4(n5891), .ZN(U2799)
         );
  AOI22_X1 U7022 ( .A1(EBX_REG_27__SCAN_IN), .A2(n6261), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6245), .ZN(n5895) );
  OAI21_X1 U7023 ( .B1(n5896), .B2(n6254), .A(n5895), .ZN(n5897) );
  AOI221_X1 U7024 ( .B1(n5906), .B2(REIP_REG_27__SCAN_IN), .C1(n5898), .C2(
        n6949), .A(n5897), .ZN(n5903) );
  OAI22_X1 U7025 ( .A1(n5900), .A2(n6193), .B1(n6176), .B2(n5899), .ZN(n5901)
         );
  INV_X1 U7026 ( .A(n5901), .ZN(n5902) );
  NAND2_X1 U7027 ( .A1(n5903), .A2(n5902), .ZN(U2800) );
  OAI22_X1 U7028 ( .A1(n5905), .A2(n6220), .B1(n5904), .B2(n6256), .ZN(n5911)
         );
  NOR2_X1 U7029 ( .A1(n5527), .A2(n5920), .ZN(n5915) );
  AOI21_X1 U7030 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5915), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5908) );
  INV_X1 U7031 ( .A(n5906), .ZN(n5907) );
  OAI22_X1 U7032 ( .A1(n5909), .A2(n6193), .B1(n5908), .B2(n5907), .ZN(n5910)
         );
  AOI211_X1 U7033 ( .C1(n5912), .C2(n6258), .A(n5911), .B(n5910), .ZN(n5913)
         );
  OAI21_X1 U7034 ( .B1(n5914), .B2(n6176), .A(n5913), .ZN(U2801) );
  AOI22_X1 U7035 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6261), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6245), .ZN(n5924) );
  INV_X1 U7036 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6647) );
  AOI22_X1 U7037 ( .A1(n5916), .A2(n6258), .B1(n5915), .B2(n6647), .ZN(n5923)
         );
  NOR2_X1 U7038 ( .A1(n6015), .A2(n6176), .ZN(n5917) );
  AOI21_X1 U7039 ( .B1(n5992), .B2(n6203), .A(n5917), .ZN(n5922) );
  NAND2_X1 U7040 ( .A1(n5919), .A2(n5918), .ZN(n5939) );
  INV_X1 U7041 ( .A(n5939), .ZN(n5925) );
  NOR2_X1 U7042 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5920), .ZN(n5932) );
  OAI21_X1 U7043 ( .B1(n5925), .B2(n5932), .A(REIP_REG_25__SCAN_IN), .ZN(n5921) );
  NAND4_X1 U7044 ( .A1(n5924), .A2(n5923), .A3(n5922), .A4(n5921), .ZN(U2802)
         );
  NAND2_X1 U7045 ( .A1(n6261), .A2(EBX_REG_24__SCAN_IN), .ZN(n5927) );
  AOI22_X1 U7046 ( .A1(n6245), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        REIP_REG_24__SCAN_IN), .B2(n5925), .ZN(n5926) );
  OAI211_X1 U7047 ( .C1(n6254), .C2(n5928), .A(n5927), .B(n5926), .ZN(n5929)
         );
  AOI21_X1 U7048 ( .B1(n5930), .B2(n6203), .A(n5929), .ZN(n5931) );
  INV_X1 U7049 ( .A(n5931), .ZN(n5933) );
  NOR2_X1 U7050 ( .A1(n5933), .A2(n5932), .ZN(n5934) );
  OAI21_X1 U7051 ( .B1(n5935), .B2(n6176), .A(n5934), .ZN(U2803) );
  AOI22_X1 U7052 ( .A1(EBX_REG_23__SCAN_IN), .A2(n6261), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6245), .ZN(n5944) );
  NAND2_X1 U7053 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .ZN(
        n5952) );
  INV_X1 U7054 ( .A(n5952), .ZN(n5936) );
  AOI21_X1 U7055 ( .B1(n5960), .B2(n5936), .A(REIP_REG_23__SCAN_IN), .ZN(n5940) );
  INV_X1 U7056 ( .A(n5937), .ZN(n5938) );
  OAI22_X1 U7057 ( .A1(n5940), .A2(n5939), .B1(n6176), .B2(n5938), .ZN(n5941)
         );
  AOI21_X1 U7058 ( .B1(n5942), .B2(n6203), .A(n5941), .ZN(n5943) );
  OAI211_X1 U7059 ( .C1(n5945), .C2(n6254), .A(n5944), .B(n5943), .ZN(U2804)
         );
  AOI22_X1 U7060 ( .A1(EBX_REG_22__SCAN_IN), .A2(n6261), .B1(n5946), .B2(n6258), .ZN(n5956) );
  NOR2_X1 U7061 ( .A1(n5948), .A2(n5947), .ZN(n5970) );
  AOI22_X1 U7062 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n6245), .B1(
        REIP_REG_22__SCAN_IN), .B2(n5970), .ZN(n5955) );
  INV_X1 U7063 ( .A(n5949), .ZN(n5950) );
  AOI22_X1 U7064 ( .A1(n5951), .A2(n6203), .B1(n6262), .B2(n5950), .ZN(n5954)
         );
  OAI211_X1 U7065 ( .C1(REIP_REG_22__SCAN_IN), .C2(REIP_REG_21__SCAN_IN), .A(
        n5960), .B(n5952), .ZN(n5953) );
  NAND4_X1 U7066 ( .A1(n5956), .A2(n5955), .A3(n5954), .A4(n5953), .ZN(U2805)
         );
  INV_X1 U7067 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6935) );
  AOI22_X1 U7068 ( .A1(EBX_REG_21__SCAN_IN), .A2(n6261), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6245), .ZN(n5957) );
  OAI21_X1 U7069 ( .B1(n5958), .B2(n6254), .A(n5957), .ZN(n5959) );
  AOI221_X1 U7070 ( .B1(n5970), .B2(REIP_REG_21__SCAN_IN), .C1(n5960), .C2(
        n6935), .A(n5959), .ZN(n5965) );
  NOR2_X1 U7071 ( .A1(n5961), .A2(n6176), .ZN(n5962) );
  AOI21_X1 U7072 ( .B1(n5963), .B2(n6203), .A(n5962), .ZN(n5964) );
  NAND2_X1 U7073 ( .A1(n5965), .A2(n5964), .ZN(U2806) );
  AOI22_X1 U7074 ( .A1(EBX_REG_20__SCAN_IN), .A2(n6261), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6245), .ZN(n5976) );
  OAI22_X1 U7075 ( .A1(n5967), .A2(n6193), .B1(n6176), .B2(n5966), .ZN(n5968)
         );
  INV_X1 U7076 ( .A(n5968), .ZN(n5975) );
  INV_X1 U7077 ( .A(n5969), .ZN(n5971) );
  OAI21_X1 U7078 ( .B1(REIP_REG_20__SCAN_IN), .B2(n5971), .A(n5970), .ZN(n5974) );
  NAND2_X1 U7079 ( .A1(n5972), .A2(n6258), .ZN(n5973) );
  NAND4_X1 U7080 ( .A1(n5976), .A2(n5975), .A3(n5974), .A4(n5973), .ZN(U2807)
         );
  NAND3_X1 U7081 ( .A1(REIP_REG_18__SCAN_IN), .A2(n5977), .A3(n5691), .ZN(
        n5983) );
  NAND2_X1 U7082 ( .A1(n6245), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5980)
         );
  INV_X1 U7083 ( .A(n6000), .ZN(n5978) );
  NAND2_X1 U7084 ( .A1(n6258), .A2(n5978), .ZN(n5979) );
  NAND3_X1 U7085 ( .A1(n5980), .A2(n5979), .A3(n6187), .ZN(n5981) );
  AOI21_X1 U7086 ( .B1(n6261), .B2(EBX_REG_19__SCAN_IN), .A(n5981), .ZN(n5982)
         );
  NAND2_X1 U7087 ( .A1(n5983), .A2(n5982), .ZN(n5984) );
  AOI21_X1 U7088 ( .B1(n5996), .B2(n6203), .A(n5984), .ZN(n5987) );
  OAI21_X1 U7089 ( .B1(n6097), .B2(n5985), .A(REIP_REG_19__SCAN_IN), .ZN(n5986) );
  OAI211_X1 U7090 ( .C1(n5988), .C2(n6176), .A(n5987), .B(n5986), .ZN(U2808)
         );
  AOI22_X1 U7091 ( .A1(n6395), .A2(REIP_REG_25__SCAN_IN), .B1(n6341), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5994) );
  OR2_X1 U7092 ( .A1(n5990), .A2(n5989), .ZN(n5991) );
  NAND2_X1 U7093 ( .A1(n4338), .A2(n5991), .ZN(n6017) );
  AOI22_X1 U7094 ( .A1(n5992), .A2(n6329), .B1(n6339), .B2(n6017), .ZN(n5993)
         );
  OAI211_X1 U7095 ( .C1(n6335), .C2(n5995), .A(n5994), .B(n5993), .ZN(U2961)
         );
  AOI22_X1 U7096 ( .A1(n6395), .A2(REIP_REG_19__SCAN_IN), .B1(n6341), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5999) );
  AOI22_X1 U7097 ( .A1(n5997), .A2(n6339), .B1(n6329), .B2(n5996), .ZN(n5998)
         );
  OAI211_X1 U7098 ( .C1(n6335), .C2(n6000), .A(n5999), .B(n5998), .ZN(U2967)
         );
  AOI22_X1 U7099 ( .A1(n6395), .A2(REIP_REG_17__SCAN_IN), .B1(n6341), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6013) );
  INV_X1 U7100 ( .A(n6002), .ZN(n6007) );
  NAND2_X1 U7101 ( .A1(n6002), .A2(n6001), .ZN(n6003) );
  OAI211_X1 U7102 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n3119), .A(n6003), .B(n6006), .ZN(n6005) );
  OAI211_X1 U7103 ( .C1(n6007), .C2(n6006), .A(n6005), .B(n6004), .ZN(n6033)
         );
  INV_X1 U7104 ( .A(n6008), .ZN(n6011) );
  INV_X1 U7105 ( .A(n5247), .ZN(n6010) );
  AOI21_X1 U7106 ( .B1(n6011), .B2(n6010), .A(n6009), .ZN(n6286) );
  AOI22_X1 U7107 ( .A1(n6033), .A2(n6339), .B1(n6286), .B2(n6329), .ZN(n6012)
         );
  OAI211_X1 U7108 ( .C1(n6335), .C2(n6100), .A(n6013), .B(n6012), .ZN(U2969)
         );
  AOI22_X1 U7109 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6395), .B1(n6014), .B2(
        n6020), .ZN(n6019) );
  INV_X1 U7110 ( .A(n6015), .ZN(n6016) );
  AOI22_X1 U7111 ( .A1(n6017), .A2(n4195), .B1(n6375), .B2(n6016), .ZN(n6018)
         );
  OAI211_X1 U7112 ( .C1(n6021), .C2(n6020), .A(n6019), .B(n6018), .ZN(U2993)
         );
  INV_X1 U7113 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6776) );
  NOR3_X1 U7114 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6035), .A3(n6022), 
        .ZN(n6023) );
  AOI21_X1 U7115 ( .B1(REIP_REG_18__SCAN_IN), .B2(n6395), .A(n6023), .ZN(n6027) );
  AOI22_X1 U7116 ( .A1(n6025), .A2(n4195), .B1(n6375), .B2(n6024), .ZN(n6026)
         );
  OAI211_X1 U7117 ( .C1(n6028), .C2(n6776), .A(n6027), .B(n6026), .ZN(U3000)
         );
  NOR2_X1 U7118 ( .A1(n6030), .A2(n6029), .ZN(n6031) );
  AOI22_X1 U7119 ( .A1(n6033), .A2(n4195), .B1(n6375), .B2(n3148), .ZN(n6039)
         );
  NOR2_X1 U7120 ( .A1(n6187), .A2(n6636), .ZN(n6034) );
  AOI221_X1 U7121 ( .B1(n6037), .B2(INSTADDRPOINTER_REG_17__SCAN_IN), .C1(
        n6036), .C2(n6035), .A(n6034), .ZN(n6038) );
  NAND2_X1 U7122 ( .A1(n6039), .A2(n6038), .ZN(U3001) );
  AOI22_X1 U7123 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n6040), .B1(n6395), .B2(REIP_REG_15__SCAN_IN), .ZN(n6044) );
  AOI22_X1 U7124 ( .A1(n6042), .A2(n4195), .B1(n6375), .B2(n6041), .ZN(n6043)
         );
  OAI211_X1 U7125 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n6045), .A(n6044), .B(n6043), .ZN(U3003) );
  NAND2_X1 U7126 ( .A1(n6046), .A2(n6348), .ZN(n6057) );
  INV_X1 U7127 ( .A(n6047), .ZN(n6049) );
  AOI221_X1 U7128 ( .B1(n6051), .B2(n6050), .C1(n6049), .C2(n6050), .A(n6048), 
        .ZN(n6055) );
  OAI22_X1 U7129 ( .A1(n6394), .A2(n6112), .B1(n5589), .B2(n6187), .ZN(n6052)
         );
  AOI21_X1 U7130 ( .B1(n6053), .B2(n4195), .A(n6052), .ZN(n6054) );
  OAI221_X1 U7131 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n6057), .C1(
        n6056), .C2(n6055), .A(n6054), .ZN(U3004) );
  INV_X1 U7132 ( .A(n6058), .ZN(n6061) );
  NAND4_X1 U7133 ( .A1(n6061), .A2(n6060), .A3(n6059), .A4(n6225), .ZN(n6062)
         );
  OAI21_X1 U7134 ( .B1(n6064), .B2(n6063), .A(n6062), .ZN(U3455) );
  AOI21_X1 U7135 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6612), .A(n6606), .ZN(n6070) );
  INV_X1 U7136 ( .A(ADS_N_REG_SCAN_IN), .ZN(n6065) );
  INV_X1 U7137 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6602) );
  NOR2_X1 U7138 ( .A1(n6602), .A2(STATE_REG_0__SCAN_IN), .ZN(n6613) );
  AOI21_X1 U7139 ( .B1(n6070), .B2(n6065), .A(n6613), .ZN(U2789) );
  INV_X1 U7140 ( .A(n6583), .ZN(n6581) );
  OAI21_X1 U7141 ( .B1(n6066), .B2(n6581), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n6067) );
  OAI21_X1 U7142 ( .B1(n6068), .B2(n6585), .A(n6067), .ZN(U2790) );
  NOR2_X1 U7143 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6071) );
  OAI21_X1 U7144 ( .B1(n6071), .B2(D_C_N_REG_SCAN_IN), .A(n6682), .ZN(n6069)
         );
  OAI21_X1 U7145 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6682), .A(n6069), .ZN(
        U2791) );
  NOR2_X1 U7146 ( .A1(n6613), .A2(n6070), .ZN(n6659) );
  OAI21_X1 U7147 ( .B1(n6071), .B2(BS16_N), .A(n6659), .ZN(n6657) );
  OAI21_X1 U7148 ( .B1(n6659), .B2(n6072), .A(n6657), .ZN(U2792) );
  OAI21_X1 U7149 ( .B1(n6075), .B2(n6074), .A(n6073), .ZN(U2793) );
  NOR4_X1 U7150 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_21__SCAN_IN), .A3(DATAWIDTH_REG_22__SCAN_IN), .A4(
        DATAWIDTH_REG_23__SCAN_IN), .ZN(n6079) );
  NOR4_X1 U7151 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_16__SCAN_IN), .A3(DATAWIDTH_REG_17__SCAN_IN), .A4(
        DATAWIDTH_REG_18__SCAN_IN), .ZN(n6078) );
  NOR4_X1 U7152 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n6077) );
  NOR4_X1 U7153 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n6076) );
  NAND4_X1 U7154 ( .A1(n6079), .A2(n6078), .A3(n6077), .A4(n6076), .ZN(n6085)
         );
  NOR4_X1 U7155 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(DATAWIDTH_REG_8__SCAN_IN), .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6083) );
  AOI211_X1 U7156 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_20__SCAN_IN), .B(
        DATAWIDTH_REG_13__SCAN_IN), .ZN(n6082) );
  NOR4_X1 U7157 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6081)
         );
  NOR4_X1 U7158 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_5__SCAN_IN), 
        .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n6080) );
  NAND4_X1 U7159 ( .A1(n6083), .A2(n6082), .A3(n6081), .A4(n6080), .ZN(n6084)
         );
  NOR2_X1 U7160 ( .A1(n6085), .A2(n6084), .ZN(n6669) );
  INV_X1 U7161 ( .A(n6669), .ZN(n6088) );
  INV_X1 U7162 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6658) );
  NAND2_X1 U7163 ( .A1(n6669), .A2(n6658), .ZN(n6090) );
  NOR3_X1 U7164 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .A3(n6090), .ZN(n6086) );
  AOI21_X1 U7165 ( .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(n6088), .A(n6086), .ZN(
        n6087) );
  OAI21_X1 U7166 ( .B1(n5096), .B2(n6088), .A(n6087), .ZN(U2794) );
  INV_X1 U7167 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n6092) );
  NOR2_X1 U7168 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_0__SCAN_IN), 
        .ZN(n6089) );
  NOR2_X1 U7169 ( .A1(n6089), .A2(n5096), .ZN(n6091) );
  OAI22_X1 U7170 ( .A1(n6669), .A2(n6092), .B1(n6091), .B2(n6090), .ZN(U2795)
         );
  NAND2_X1 U7171 ( .A1(n6636), .A2(n6093), .ZN(n6096) );
  AOI22_X1 U7172 ( .A1(EBX_REG_17__SCAN_IN), .A2(n6261), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6245), .ZN(n6094) );
  INV_X1 U7173 ( .A(n6094), .ZN(n6095) );
  AOI211_X1 U7174 ( .C1(n6097), .C2(n6096), .A(n6395), .B(n6095), .ZN(n6099)
         );
  AOI22_X1 U7175 ( .A1(n6286), .A2(n6203), .B1(n6262), .B2(n3148), .ZN(n6098)
         );
  OAI211_X1 U7176 ( .C1(n6100), .C2(n6254), .A(n6099), .B(n6098), .ZN(U2810)
         );
  INV_X1 U7177 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6104) );
  XOR2_X1 U7178 ( .A(REIP_REG_16__SCAN_IN), .B(REIP_REG_15__SCAN_IN), .Z(n6101) );
  AOI22_X1 U7179 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6111), .B1(n6102), .B2(
        n6101), .ZN(n6103) );
  OAI211_X1 U7180 ( .C1(n6256), .C2(n6104), .A(n6103), .B(n6187), .ZN(n6105)
         );
  AOI21_X1 U7181 ( .B1(EBX_REG_16__SCAN_IN), .B2(n6261), .A(n6105), .ZN(n6109)
         );
  INV_X1 U7182 ( .A(n6106), .ZN(n6107) );
  AOI22_X1 U7183 ( .A1(n6290), .A2(n6203), .B1(n6107), .B2(n6258), .ZN(n6108)
         );
  OAI211_X1 U7184 ( .C1(n6176), .C2(n6110), .A(n6109), .B(n6108), .ZN(U2811)
         );
  AOI21_X1 U7185 ( .B1(n6245), .B2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n6395), 
        .ZN(n6120) );
  AOI22_X1 U7186 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6261), .B1(
        REIP_REG_14__SCAN_IN), .B2(n6111), .ZN(n6119) );
  OAI22_X1 U7187 ( .A1(n6113), .A2(n6193), .B1(n6176), .B2(n6112), .ZN(n6114)
         );
  AOI21_X1 U7188 ( .B1(n6115), .B2(n6258), .A(n6114), .ZN(n6118) );
  NAND3_X1 U7189 ( .A1(n6244), .A2(n5589), .A3(n6116), .ZN(n6117) );
  NAND4_X1 U7190 ( .A1(n6120), .A2(n6119), .A3(n6118), .A4(n6117), .ZN(U2813)
         );
  NOR3_X1 U7191 ( .A1(n6239), .A2(REIP_REG_13__SCAN_IN), .A3(n6121), .ZN(n6122) );
  AOI211_X1 U7192 ( .C1(n6245), .C2(PHYADDRPOINTER_REG_13__SCAN_IN), .A(n6395), 
        .B(n6122), .ZN(n6129) );
  AOI22_X1 U7193 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6261), .B1(n6262), .B2(n6123), .ZN(n6128) );
  INV_X1 U7194 ( .A(n6124), .ZN(n6125) );
  AOI22_X1 U7195 ( .A1(n6297), .A2(n6203), .B1(n6125), .B2(n6258), .ZN(n6127)
         );
  OAI21_X1 U7196 ( .B1(n6239), .B2(n6131), .A(n6271), .ZN(n6139) );
  NOR2_X1 U7197 ( .A1(n6239), .A2(REIP_REG_12__SCAN_IN), .ZN(n6130) );
  OAI21_X1 U7198 ( .B1(n6139), .B2(n6130), .A(REIP_REG_13__SCAN_IN), .ZN(n6126) );
  NAND4_X1 U7199 ( .A1(n6129), .A2(n6128), .A3(n6127), .A4(n6126), .ZN(U2814)
         );
  AOI22_X1 U7200 ( .A1(n6262), .A2(n6278), .B1(n6131), .B2(n6130), .ZN(n6137)
         );
  OAI22_X1 U7201 ( .A1(n6283), .A2(n6220), .B1(n6914), .B2(n6256), .ZN(n6132)
         );
  AOI211_X1 U7202 ( .C1(REIP_REG_12__SCAN_IN), .C2(n6139), .A(n6395), .B(n6132), .ZN(n6136) );
  INV_X1 U7203 ( .A(n6133), .ZN(n6281) );
  AOI22_X1 U7204 ( .A1(n6281), .A2(n6203), .B1(n6134), .B2(n6258), .ZN(n6135)
         );
  NAND3_X1 U7205 ( .A1(n6137), .A2(n6136), .A3(n6135), .ZN(U2815) );
  INV_X1 U7206 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6150) );
  OAI21_X1 U7207 ( .B1(n6239), .B2(n6138), .A(n6629), .ZN(n6140) );
  NAND2_X1 U7208 ( .A1(n6140), .A2(n6139), .ZN(n6149) );
  INV_X1 U7209 ( .A(n6141), .ZN(n6147) );
  NOR2_X1 U7210 ( .A1(n6176), .A2(n6142), .ZN(n6143) );
  AOI211_X1 U7211 ( .C1(n6245), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6395), 
        .B(n6143), .ZN(n6144) );
  OAI21_X1 U7212 ( .B1(n6145), .B2(n6193), .A(n6144), .ZN(n6146) );
  AOI21_X1 U7213 ( .B1(n6147), .B2(n6258), .A(n6146), .ZN(n6148) );
  OAI211_X1 U7214 ( .C1(n6150), .C2(n6220), .A(n6149), .B(n6148), .ZN(U2816)
         );
  OAI22_X1 U7215 ( .A1(n6152), .A2(n6220), .B1(n6176), .B2(n6151), .ZN(n6153)
         );
  AOI211_X1 U7216 ( .C1(n6245), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6395), 
        .B(n6153), .ZN(n6163) );
  AOI22_X1 U7217 ( .A1(n6155), .A2(n6203), .B1(n6258), .B2(n6154), .ZN(n6162)
         );
  NAND2_X1 U7218 ( .A1(n6244), .A2(n6157), .ZN(n6156) );
  AND2_X1 U7219 ( .A1(n6156), .A2(n6271), .ZN(n6183) );
  INV_X1 U7220 ( .A(n6183), .ZN(n6165) );
  NOR3_X1 U7221 ( .A1(n6239), .A2(REIP_REG_9__SCAN_IN), .A3(n6157), .ZN(n6164)
         );
  OAI21_X1 U7222 ( .B1(n6165), .B2(n6164), .A(REIP_REG_10__SCAN_IN), .ZN(n6161) );
  NAND3_X1 U7223 ( .A1(n6244), .A2(n6159), .A3(n6158), .ZN(n6160) );
  NAND4_X1 U7224 ( .A1(n6163), .A2(n6162), .A3(n6161), .A4(n6160), .ZN(U2817)
         );
  AOI21_X1 U7225 ( .B1(n6165), .B2(REIP_REG_9__SCAN_IN), .A(n6164), .ZN(n6173)
         );
  NOR2_X1 U7226 ( .A1(n6176), .A2(n6166), .ZN(n6167) );
  AOI211_X1 U7227 ( .C1(n6245), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n6395), 
        .B(n6167), .ZN(n6168) );
  OAI21_X1 U7228 ( .B1(n6169), .B2(n6193), .A(n6168), .ZN(n6170) );
  AOI21_X1 U7229 ( .B1(n6171), .B2(n6258), .A(n6170), .ZN(n6172) );
  OAI211_X1 U7230 ( .C1(n6767), .C2(n6220), .A(n6173), .B(n6172), .ZN(U2818)
         );
  AOI21_X1 U7231 ( .B1(n6244), .B2(n6174), .A(REIP_REG_8__SCAN_IN), .ZN(n6184)
         );
  OAI22_X1 U7232 ( .A1(n6838), .A2(n6256), .B1(n6176), .B2(n6175), .ZN(n6177)
         );
  AOI211_X1 U7233 ( .C1(n6261), .C2(EBX_REG_8__SCAN_IN), .A(n6395), .B(n6177), 
        .ZN(n6182) );
  INV_X1 U7234 ( .A(n6178), .ZN(n6180) );
  AOI22_X1 U7235 ( .A1(n6180), .A2(n6203), .B1(n6258), .B2(n6179), .ZN(n6181)
         );
  OAI211_X1 U7236 ( .C1(n6184), .C2(n6183), .A(n6182), .B(n6181), .ZN(U2819)
         );
  NOR2_X1 U7237 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6185), .ZN(n6191) );
  NAND2_X1 U7238 ( .A1(n6245), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n6189)
         );
  INV_X1 U7239 ( .A(n6186), .ZN(n6364) );
  AOI22_X1 U7240 ( .A1(EBX_REG_7__SCAN_IN), .A2(n6261), .B1(n6262), .B2(n6364), 
        .ZN(n6188) );
  NAND3_X1 U7241 ( .A1(n6189), .A2(n6188), .A3(n6187), .ZN(n6190) );
  AOI21_X1 U7242 ( .B1(n6244), .B2(n6191), .A(n6190), .ZN(n6192) );
  OAI21_X1 U7243 ( .B1(n6194), .B2(n6193), .A(n6192), .ZN(n6195) );
  INV_X1 U7244 ( .A(n6195), .ZN(n6198) );
  OAI21_X1 U7245 ( .B1(n6239), .B2(n6196), .A(n6271), .ZN(n6215) );
  NOR4_X1 U7246 ( .A1(n6239), .A2(n6620), .A3(REIP_REG_6__SCAN_IN), .A4(n6212), 
        .ZN(n6200) );
  OAI21_X1 U7247 ( .B1(n6215), .B2(n6200), .A(REIP_REG_7__SCAN_IN), .ZN(n6197)
         );
  OAI211_X1 U7248 ( .C1(n6254), .C2(n6199), .A(n6198), .B(n6197), .ZN(U2820)
         );
  AOI21_X1 U7249 ( .B1(n6201), .B2(n6262), .A(n6200), .ZN(n6208) );
  AOI22_X1 U7250 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n6245), .B1(
        REIP_REG_6__SCAN_IN), .B2(n6215), .ZN(n6207) );
  AOI21_X1 U7251 ( .B1(n6261), .B2(EBX_REG_6__SCAN_IN), .A(n6395), .ZN(n6206)
         );
  AOI22_X1 U7252 ( .A1(n6204), .A2(n6203), .B1(n6202), .B2(n6258), .ZN(n6205)
         );
  NAND4_X1 U7253 ( .A1(n6208), .A2(n6207), .A3(n6206), .A4(n6205), .ZN(U2821)
         );
  AOI22_X1 U7254 ( .A1(EBX_REG_5__SCAN_IN), .A2(n6261), .B1(
        PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n6245), .ZN(n6209) );
  INV_X1 U7255 ( .A(n6209), .ZN(n6210) );
  AOI211_X1 U7256 ( .C1(n6262), .C2(n6211), .A(n6395), .B(n6210), .ZN(n6217)
         );
  OAI21_X1 U7257 ( .B1(n6239), .B2(n6212), .A(n6620), .ZN(n6214) );
  AOI22_X1 U7258 ( .A1(n6215), .A2(n6214), .B1(n6213), .B2(n6264), .ZN(n6216)
         );
  OAI211_X1 U7259 ( .C1(n6218), .C2(n6254), .A(n6217), .B(n6216), .ZN(U2822)
         );
  OAI21_X1 U7260 ( .B1(n6239), .B2(n6222), .A(n6271), .ZN(n6240) );
  OAI22_X1 U7261 ( .A1(n6982), .A2(n6220), .B1(n6219), .B2(n6256), .ZN(n6221)
         );
  AOI211_X1 U7262 ( .C1(REIP_REG_4__SCAN_IN), .C2(n6240), .A(n6395), .B(n6221), 
        .ZN(n6231) );
  NAND3_X1 U7263 ( .A1(n6244), .A2(n6617), .A3(n6222), .ZN(n6229) );
  NAND2_X1 U7264 ( .A1(n6223), .A2(n6264), .ZN(n6228) );
  NAND2_X1 U7265 ( .A1(n6262), .A2(n6224), .ZN(n6227) );
  NAND2_X1 U7266 ( .A1(n6260), .A2(n6225), .ZN(n6226) );
  AND4_X1 U7267 ( .A1(n6229), .A2(n6228), .A3(n6227), .A4(n6226), .ZN(n6230)
         );
  OAI211_X1 U7268 ( .C1(n6232), .C2(n6254), .A(n6231), .B(n6230), .ZN(U2823)
         );
  INV_X1 U7269 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6885) );
  AOI22_X1 U7270 ( .A1(n6260), .A2(n4527), .B1(n6245), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U7271 ( .A1(n6264), .A2(n6233), .ZN(n6237) );
  NAND2_X1 U7272 ( .A1(n6262), .A2(n6234), .ZN(n6236) );
  NAND2_X1 U7273 ( .A1(n6261), .A2(EBX_REG_3__SCAN_IN), .ZN(n6235) );
  AND4_X1 U7274 ( .A1(n6238), .A2(n6237), .A3(n6236), .A4(n6235), .ZN(n6242)
         );
  OR2_X1 U7275 ( .A1(n6239), .A2(REIP_REG_1__SCAN_IN), .ZN(n6255) );
  AND3_X1 U7276 ( .A1(n6255), .A2(n6271), .A3(REIP_REG_2__SCAN_IN), .ZN(n6250)
         );
  OAI21_X1 U7277 ( .B1(REIP_REG_3__SCAN_IN), .B2(n6250), .A(n6240), .ZN(n6241)
         );
  OAI211_X1 U7278 ( .C1(n6254), .C2(n6243), .A(n6242), .B(n6241), .ZN(U2824)
         );
  AOI22_X1 U7279 ( .A1(EBX_REG_2__SCAN_IN), .A2(n6261), .B1(n6262), .B2(n6374), 
        .ZN(n6253) );
  AOI21_X1 U7280 ( .B1(n6244), .B2(REIP_REG_1__SCAN_IN), .A(
        REIP_REG_2__SCAN_IN), .ZN(n6249) );
  AOI22_X1 U7281 ( .A1(n6260), .A2(n6246), .B1(n6245), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6248) );
  NAND2_X1 U7282 ( .A1(n6264), .A2(n6330), .ZN(n6247) );
  OAI211_X1 U7283 ( .C1(n6250), .C2(n6249), .A(n6248), .B(n6247), .ZN(n6251)
         );
  INV_X1 U7284 ( .A(n6251), .ZN(n6252) );
  OAI211_X1 U7285 ( .C1(n6334), .C2(n6254), .A(n6253), .B(n6252), .ZN(U2825)
         );
  OAI21_X1 U7286 ( .B1(n6256), .B2(n5099), .A(n6255), .ZN(n6257) );
  INV_X1 U7287 ( .A(n6257), .ZN(n6270) );
  AOI22_X1 U7288 ( .A1(n6260), .A2(n6259), .B1(n6258), .B2(n5099), .ZN(n6268)
         );
  NAND2_X1 U7289 ( .A1(n6261), .A2(EBX_REG_1__SCAN_IN), .ZN(n6267) );
  NAND2_X1 U7290 ( .A1(n6262), .A2(n4464), .ZN(n6266) );
  NAND2_X1 U7291 ( .A1(n6264), .A2(n6263), .ZN(n6265) );
  AND4_X1 U7292 ( .A1(n6268), .A2(n6267), .A3(n6266), .A4(n6265), .ZN(n6269)
         );
  OAI211_X1 U7293 ( .C1(n6271), .C2(n5096), .A(n6270), .B(n6269), .ZN(U2826)
         );
  AOI22_X1 U7294 ( .A1(n6286), .A2(n6280), .B1(n6279), .B2(n3148), .ZN(n6272)
         );
  OAI21_X1 U7295 ( .B1(n6284), .B2(n6923), .A(n6272), .ZN(U2842) );
  NOR2_X1 U7296 ( .A1(n6274), .A2(n6273), .ZN(n6275) );
  AOI21_X1 U7297 ( .B1(n6297), .B2(n6280), .A(n6275), .ZN(n6276) );
  OAI21_X1 U7298 ( .B1(n6284), .B2(n6277), .A(n6276), .ZN(U2846) );
  AOI22_X1 U7299 ( .A1(n6281), .A2(n6280), .B1(n6279), .B2(n6278), .ZN(n6282)
         );
  OAI21_X1 U7300 ( .B1(n6284), .B2(n6283), .A(n6282), .ZN(U2847) );
  INV_X1 U7301 ( .A(n6285), .ZN(n6296) );
  AOI22_X1 U7302 ( .A1(n6286), .A2(n6296), .B1(n6289), .B2(DATAI_17_), .ZN(
        n6288) );
  AOI22_X1 U7303 ( .A1(n6292), .A2(DATAI_1_), .B1(n6291), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U7304 ( .A1(n6288), .A2(n6287), .ZN(U2874) );
  AOI22_X1 U7305 ( .A1(n6290), .A2(n6296), .B1(n6289), .B2(DATAI_16_), .ZN(
        n6294) );
  AOI22_X1 U7306 ( .A1(n6292), .A2(DATAI_0_), .B1(n6291), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6293) );
  NAND2_X1 U7307 ( .A1(n6294), .A2(n6293), .ZN(U2875) );
  AOI22_X1 U7308 ( .A1(n6297), .A2(n6296), .B1(DATAI_13_), .B2(n6295), .ZN(
        n6298) );
  OAI21_X1 U7309 ( .B1(n6305), .B2(n6299), .A(n6298), .ZN(U2878) );
  AOI22_X1 U7310 ( .A1(n6674), .A2(LWORD_REG_15__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6301) );
  OAI21_X1 U7311 ( .B1(n6302), .B2(n6325), .A(n6301), .ZN(U2908) );
  AOI22_X1 U7312 ( .A1(n6674), .A2(LWORD_REG_14__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6303) );
  OAI21_X1 U7313 ( .B1(n5106), .B2(n6325), .A(n6303), .ZN(U2909) );
  AOI22_X1 U7314 ( .A1(n6674), .A2(LWORD_REG_13__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6304) );
  OAI21_X1 U7315 ( .B1(n6305), .B2(n6325), .A(n6304), .ZN(U2910) );
  AOI22_X1 U7316 ( .A1(n6674), .A2(LWORD_REG_12__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6306) );
  OAI21_X1 U7317 ( .B1(n5038), .B2(n6325), .A(n6306), .ZN(U2911) );
  AOI22_X1 U7318 ( .A1(n6674), .A2(LWORD_REG_11__SCAN_IN), .B1(n6316), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6307) );
  OAI21_X1 U7319 ( .B1(n6860), .B2(n6325), .A(n6307), .ZN(U2912) );
  AOI22_X1 U7320 ( .A1(n6674), .A2(LWORD_REG_10__SCAN_IN), .B1(n6316), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6308) );
  OAI21_X1 U7321 ( .B1(n6309), .B2(n6325), .A(n6308), .ZN(U2913) );
  AOI22_X1 U7322 ( .A1(n6674), .A2(LWORD_REG_9__SCAN_IN), .B1(n6316), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6310) );
  OAI21_X1 U7323 ( .B1(n6311), .B2(n6325), .A(n6310), .ZN(U2914) );
  AOI22_X1 U7324 ( .A1(n6674), .A2(LWORD_REG_8__SCAN_IN), .B1(n6316), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6312) );
  OAI21_X1 U7325 ( .B1(n6313), .B2(n6325), .A(n6312), .ZN(U2915) );
  AOI22_X1 U7326 ( .A1(n6674), .A2(LWORD_REG_7__SCAN_IN), .B1(n6316), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6314) );
  OAI21_X1 U7327 ( .B1(n4922), .B2(n6325), .A(n6314), .ZN(U2916) );
  AOI22_X1 U7328 ( .A1(n6674), .A2(LWORD_REG_6__SCAN_IN), .B1(n6316), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6315) );
  OAI21_X1 U7329 ( .B1(n4853), .B2(n6325), .A(n6315), .ZN(U2917) );
  AOI22_X1 U7330 ( .A1(n6674), .A2(LWORD_REG_5__SCAN_IN), .B1(n6316), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6317) );
  OAI21_X1 U7331 ( .B1(n3787), .B2(n6325), .A(n6317), .ZN(U2918) );
  AOI22_X1 U7332 ( .A1(n6674), .A2(LWORD_REG_4__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6318) );
  OAI21_X1 U7333 ( .B1(n6939), .B2(n6325), .A(n6318), .ZN(U2919) );
  AOI22_X1 U7334 ( .A1(n6674), .A2(LWORD_REG_3__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6319) );
  OAI21_X1 U7335 ( .B1(n3667), .B2(n6325), .A(n6319), .ZN(U2920) );
  AOI22_X1 U7336 ( .A1(n6674), .A2(LWORD_REG_2__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6320) );
  OAI21_X1 U7337 ( .B1(n6321), .B2(n6325), .A(n6320), .ZN(U2921) );
  AOI22_X1 U7338 ( .A1(n6674), .A2(LWORD_REG_1__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6322) );
  OAI21_X1 U7339 ( .B1(n3643), .B2(n6325), .A(n6322), .ZN(U2922) );
  AOI22_X1 U7340 ( .A1(n6674), .A2(LWORD_REG_0__SCAN_IN), .B1(n6323), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6324) );
  OAI21_X1 U7341 ( .B1(n3650), .B2(n6325), .A(n6324), .ZN(U2923) );
  AOI22_X1 U7342 ( .A1(n6395), .A2(REIP_REG_2__SCAN_IN), .B1(n6341), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6333) );
  XNOR2_X1 U7343 ( .A(n6326), .B(n6372), .ZN(n6328) );
  XNOR2_X1 U7344 ( .A(n6328), .B(n6327), .ZN(n6382) );
  INV_X1 U7345 ( .A(n6382), .ZN(n6331) );
  AOI22_X1 U7346 ( .A1(n6339), .A2(n6331), .B1(n6330), .B2(n6329), .ZN(n6332)
         );
  OAI211_X1 U7347 ( .C1(n6335), .C2(n6334), .A(n6333), .B(n6332), .ZN(U2984)
         );
  INV_X1 U7348 ( .A(n6336), .ZN(n6337) );
  AOI21_X1 U7349 ( .B1(n6339), .B2(n6338), .A(n6337), .ZN(n6343) );
  OAI21_X1 U7350 ( .B1(n6341), .B2(n6340), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n6342) );
  OAI211_X1 U7351 ( .C1(n6345), .C2(n6344), .A(n6343), .B(n6342), .ZN(U2986)
         );
  AOI21_X1 U7352 ( .B1(n6375), .B2(n6347), .A(n6346), .ZN(n6351) );
  AOI22_X1 U7353 ( .A1(n6349), .A2(n4195), .B1(n6348), .B2(n6882), .ZN(n6350)
         );
  OAI211_X1 U7354 ( .C1(n6352), .C2(n6882), .A(n6351), .B(n6350), .ZN(U3007)
         );
  INV_X1 U7355 ( .A(n6353), .ZN(n6354) );
  AOI21_X1 U7356 ( .B1(n6375), .B2(n6355), .A(n6354), .ZN(n6359) );
  AOI22_X1 U7357 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n6357), .B1(n6356), 
        .B2(n4195), .ZN(n6358) );
  OAI211_X1 U7358 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6360), .A(n6359), 
        .B(n6358), .ZN(U3009) );
  NAND2_X1 U7359 ( .A1(n6362), .A2(n6361), .ZN(n6366) );
  AOI21_X1 U7360 ( .B1(n6375), .B2(n6364), .A(n6363), .ZN(n6365) );
  OAI211_X1 U7361 ( .C1(n6367), .C2(n6399), .A(n6366), .B(n6365), .ZN(n6368)
         );
  INV_X1 U7362 ( .A(n6368), .ZN(n6369) );
  OAI21_X1 U7363 ( .B1(n6370), .B2(n6361), .A(n6369), .ZN(U3011) );
  OAI21_X1 U7364 ( .B1(n6373), .B2(n6372), .A(n6371), .ZN(n6376) );
  AOI22_X1 U7365 ( .A1(n6377), .A2(n6376), .B1(n6375), .B2(n6374), .ZN(n6386)
         );
  NOR2_X1 U7366 ( .A1(n4201), .A2(n6378), .ZN(n6381) );
  INV_X1 U7367 ( .A(n6379), .ZN(n6380) );
  MUX2_X1 U7368 ( .A(n6381), .B(n6380), .S(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .Z(n6384) );
  NOR2_X1 U7369 ( .A1(n6382), .A2(n6399), .ZN(n6383) );
  NOR2_X1 U7370 ( .A1(n6384), .A2(n6383), .ZN(n6385) );
  OAI211_X1 U7371 ( .C1(n6187), .C2(n6387), .A(n6386), .B(n6385), .ZN(U3016)
         );
  NAND2_X1 U7372 ( .A1(n6389), .A2(n6388), .ZN(n6403) );
  AOI21_X1 U7373 ( .B1(n6392), .B2(n6391), .A(n6390), .ZN(n6402) );
  OR2_X1 U7374 ( .A1(n6394), .A2(n6393), .ZN(n6397) );
  NAND2_X1 U7375 ( .A1(n6395), .A2(REIP_REG_1__SCAN_IN), .ZN(n6396) );
  OAI211_X1 U7376 ( .C1(n6399), .C2(n6398), .A(n6397), .B(n6396), .ZN(n6400)
         );
  INV_X1 U7377 ( .A(n6400), .ZN(n6401) );
  OAI221_X1 U7378 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n6403), .C1(n4201), .C2(n6402), .A(n6401), .ZN(U3017) );
  NOR2_X1 U7379 ( .A1(n6561), .A2(n6404), .ZN(U3019) );
  NAND3_X1 U7380 ( .A1(n6406), .A2(n6405), .A3(n6563), .ZN(n6407) );
  OAI21_X1 U7381 ( .B1(n6409), .B2(n6408), .A(n6407), .ZN(n6441) );
  NAND2_X1 U7382 ( .A1(n6411), .A2(n6410), .ZN(n6412) );
  INV_X1 U7383 ( .A(n6412), .ZN(n6442) );
  AOI22_X1 U7384 ( .A1(n6484), .A2(n6441), .B1(n6470), .B2(n6442), .ZN(n6423)
         );
  AOI21_X1 U7385 ( .B1(n6412), .B2(STATE2_REG_3__SCAN_IN), .A(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6419) );
  INV_X1 U7386 ( .A(n6466), .ZN(n6414) );
  NOR3_X1 U7387 ( .A1(n6443), .A2(n6414), .A3(n6477), .ZN(n6417) );
  OAI21_X1 U7388 ( .B1(n6417), .B2(n6416), .A(n6415), .ZN(n6418) );
  NAND3_X1 U7389 ( .A1(n6420), .A2(n6419), .A3(n6418), .ZN(n6445) );
  AOI22_X1 U7390 ( .A1(n6445), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6421), 
        .B2(n6443), .ZN(n6422) );
  OAI211_X1 U7391 ( .C1(n6424), .C2(n6466), .A(n6423), .B(n6422), .ZN(U3068)
         );
  AOI22_X1 U7392 ( .A1(n6490), .A2(n6441), .B1(n6489), .B2(n6442), .ZN(n6426)
         );
  AOI22_X1 U7393 ( .A1(n6445), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6488), 
        .B2(n6443), .ZN(n6425) );
  OAI211_X1 U7394 ( .C1(n6493), .C2(n6466), .A(n6426), .B(n6425), .ZN(U3069)
         );
  AOI22_X1 U7395 ( .A1(n6496), .A2(n6441), .B1(n6495), .B2(n6442), .ZN(n6429)
         );
  AOI22_X1 U7396 ( .A1(n6445), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6427), 
        .B2(n6443), .ZN(n6428) );
  OAI211_X1 U7397 ( .C1(n6430), .C2(n6466), .A(n6429), .B(n6428), .ZN(U3070)
         );
  AOI22_X1 U7398 ( .A1(n6502), .A2(n6441), .B1(n6501), .B2(n6442), .ZN(n6433)
         );
  AOI22_X1 U7399 ( .A1(n6445), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6431), 
        .B2(n6443), .ZN(n6432) );
  OAI211_X1 U7400 ( .C1(n6434), .C2(n6466), .A(n6433), .B(n6432), .ZN(U3071)
         );
  AOI22_X1 U7401 ( .A1(n6508), .A2(n6441), .B1(n6507), .B2(n6442), .ZN(n6436)
         );
  AOI22_X1 U7402 ( .A1(n6445), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6506), 
        .B2(n6443), .ZN(n6435) );
  OAI211_X1 U7403 ( .C1(n6511), .C2(n6466), .A(n6436), .B(n6435), .ZN(U3072)
         );
  AOI22_X1 U7404 ( .A1(n6514), .A2(n6441), .B1(n6513), .B2(n6442), .ZN(n6438)
         );
  AOI22_X1 U7405 ( .A1(n6445), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6512), 
        .B2(n6443), .ZN(n6437) );
  OAI211_X1 U7406 ( .C1(n6517), .C2(n6466), .A(n6438), .B(n6437), .ZN(U3073)
         );
  AOI22_X1 U7407 ( .A1(n6520), .A2(n6442), .B1(n6521), .B2(n6441), .ZN(n6440)
         );
  AOI22_X1 U7408 ( .A1(n6445), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6519), 
        .B2(n6443), .ZN(n6439) );
  OAI211_X1 U7409 ( .C1(n6525), .C2(n6466), .A(n6440), .B(n6439), .ZN(U3074)
         );
  AOI22_X1 U7410 ( .A1(n6529), .A2(n6442), .B1(n6531), .B2(n6441), .ZN(n6447)
         );
  AOI22_X1 U7411 ( .A1(n6445), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6444), 
        .B2(n6443), .ZN(n6446) );
  OAI211_X1 U7412 ( .C1(n6448), .C2(n6466), .A(n6447), .B(n6446), .ZN(U3075)
         );
  INV_X1 U7413 ( .A(n6449), .ZN(n6461) );
  INV_X1 U7414 ( .A(n6450), .ZN(n6459) );
  AOI22_X1 U7415 ( .A1(n6495), .A2(n6461), .B1(n6494), .B2(n6459), .ZN(n6452)
         );
  AOI22_X1 U7416 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6463), .B1(n6496), 
        .B2(n6462), .ZN(n6451) );
  OAI211_X1 U7417 ( .C1(n6499), .C2(n6466), .A(n6452), .B(n6451), .ZN(U3078)
         );
  AOI22_X1 U7418 ( .A1(n6501), .A2(n6461), .B1(n6500), .B2(n6459), .ZN(n6454)
         );
  AOI22_X1 U7419 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6463), .B1(n6502), 
        .B2(n6462), .ZN(n6453) );
  OAI211_X1 U7420 ( .C1(n6505), .C2(n6466), .A(n6454), .B(n6453), .ZN(U3079)
         );
  AOI22_X1 U7421 ( .A1(n6513), .A2(n6461), .B1(n6455), .B2(n6459), .ZN(n6457)
         );
  AOI22_X1 U7422 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6463), .B1(n6514), 
        .B2(n6462), .ZN(n6456) );
  OAI211_X1 U7423 ( .C1(n6458), .C2(n6466), .A(n6457), .B(n6456), .ZN(U3081)
         );
  AOI22_X1 U7424 ( .A1(n6520), .A2(n6461), .B1(n6460), .B2(n6459), .ZN(n6465)
         );
  AOI22_X1 U7425 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6463), .B1(n6521), 
        .B2(n6462), .ZN(n6464) );
  OAI211_X1 U7426 ( .C1(n6467), .C2(n6466), .A(n6465), .B(n6464), .ZN(U3082)
         );
  NOR2_X1 U7427 ( .A1(n6468), .A2(n6563), .ZN(n6528) );
  AOI22_X1 U7428 ( .A1(n6470), .A2(n6528), .B1(n6469), .B2(n6526), .ZN(n6486)
         );
  OAI21_X1 U7429 ( .B1(n6473), .B2(n6472), .A(n6471), .ZN(n6483) );
  AOI21_X1 U7430 ( .B1(n6475), .B2(n6474), .A(n6528), .ZN(n6482) );
  INV_X1 U7431 ( .A(n6482), .ZN(n6479) );
  AOI21_X1 U7432 ( .B1(n6477), .B2(n6481), .A(n6476), .ZN(n6478) );
  OAI21_X1 U7433 ( .B1(n6483), .B2(n6479), .A(n6478), .ZN(n6532) );
  OAI22_X1 U7434 ( .A1(n6483), .A2(n6482), .B1(n6481), .B2(n6480), .ZN(n6530)
         );
  AOI22_X1 U7435 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6532), .B1(n6484), 
        .B2(n6530), .ZN(n6485) );
  OAI211_X1 U7436 ( .C1(n6487), .C2(n6535), .A(n6486), .B(n6485), .ZN(U3108)
         );
  AOI22_X1 U7437 ( .A1(n6489), .A2(n6528), .B1(n6488), .B2(n6518), .ZN(n6492)
         );
  AOI22_X1 U7438 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6532), .B1(n6490), 
        .B2(n6530), .ZN(n6491) );
  OAI211_X1 U7439 ( .C1(n6493), .C2(n6524), .A(n6492), .B(n6491), .ZN(U3109)
         );
  AOI22_X1 U7440 ( .A1(n6495), .A2(n6528), .B1(n6494), .B2(n6526), .ZN(n6498)
         );
  AOI22_X1 U7441 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6532), .B1(n6496), 
        .B2(n6530), .ZN(n6497) );
  OAI211_X1 U7442 ( .C1(n6499), .C2(n6535), .A(n6498), .B(n6497), .ZN(U3110)
         );
  AOI22_X1 U7443 ( .A1(n6501), .A2(n6528), .B1(n6500), .B2(n6526), .ZN(n6504)
         );
  AOI22_X1 U7444 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6532), .B1(n6502), 
        .B2(n6530), .ZN(n6503) );
  OAI211_X1 U7445 ( .C1(n6505), .C2(n6535), .A(n6504), .B(n6503), .ZN(U3111)
         );
  AOI22_X1 U7446 ( .A1(n6507), .A2(n6528), .B1(n6506), .B2(n6518), .ZN(n6510)
         );
  AOI22_X1 U7447 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6532), .B1(n6508), 
        .B2(n6530), .ZN(n6509) );
  OAI211_X1 U7448 ( .C1(n6511), .C2(n6524), .A(n6510), .B(n6509), .ZN(U3112)
         );
  AOI22_X1 U7449 ( .A1(n6513), .A2(n6528), .B1(n6512), .B2(n6518), .ZN(n6516)
         );
  AOI22_X1 U7450 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6532), .B1(n6514), 
        .B2(n6530), .ZN(n6515) );
  OAI211_X1 U7451 ( .C1(n6517), .C2(n6524), .A(n6516), .B(n6515), .ZN(U3113)
         );
  AOI22_X1 U7452 ( .A1(n6520), .A2(n6528), .B1(n6519), .B2(n6518), .ZN(n6523)
         );
  AOI22_X1 U7453 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6532), .B1(n6521), 
        .B2(n6530), .ZN(n6522) );
  OAI211_X1 U7454 ( .C1(n6525), .C2(n6524), .A(n6523), .B(n6522), .ZN(U3114)
         );
  AOI22_X1 U7455 ( .A1(n6529), .A2(n6528), .B1(n6527), .B2(n6526), .ZN(n6534)
         );
  AOI22_X1 U7456 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6532), .B1(n6531), 
        .B2(n6530), .ZN(n6533) );
  OAI211_X1 U7457 ( .C1(n6536), .C2(n6535), .A(n6534), .B(n6533), .ZN(U3115)
         );
  NOR2_X1 U7458 ( .A1(FLUSH_REG_SCAN_IN), .A2(MORE_REG_SCAN_IN), .ZN(n6540) );
  NOR2_X1 U7459 ( .A1(n6538), .A2(n6537), .ZN(n6539) );
  OAI21_X1 U7460 ( .B1(n6541), .B2(n6540), .A(n6539), .ZN(n6542) );
  NOR2_X1 U7461 ( .A1(n6543), .A2(n6542), .ZN(n6567) );
  OAI211_X1 U7462 ( .C1(n6546), .C2(n6545), .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n6544), .ZN(n6550) );
  INV_X1 U7463 ( .A(n6547), .ZN(n6549) );
  OAI211_X1 U7464 ( .C1(n6948), .C2(n6550), .A(n6549), .B(n6548), .ZN(n6552)
         );
  NAND2_X1 U7465 ( .A1(n6948), .A2(n6550), .ZN(n6551) );
  NAND2_X1 U7466 ( .A1(n6552), .A2(n6551), .ZN(n6558) );
  INV_X1 U7467 ( .A(n6553), .ZN(n6555) );
  NAND2_X1 U7468 ( .A1(n6557), .A2(n6558), .ZN(n6554) );
  NAND2_X1 U7469 ( .A1(n6555), .A2(n6554), .ZN(n6556) );
  OAI21_X1 U7470 ( .B1(n6558), .B2(n6557), .A(n6556), .ZN(n6560) );
  NAND2_X1 U7471 ( .A1(n6564), .A2(n6563), .ZN(n6559) );
  NAND2_X1 U7472 ( .A1(n6560), .A2(n6559), .ZN(n6562) );
  OAI211_X1 U7473 ( .C1(n6564), .C2(n6563), .A(n6562), .B(n6561), .ZN(n6565)
         );
  AND3_X1 U7474 ( .A1(n6567), .A2(n6566), .A3(n6565), .ZN(n6582) );
  NAND2_X1 U7475 ( .A1(n6582), .A2(n6583), .ZN(n6569) );
  NAND2_X1 U7476 ( .A1(READY_N), .A2(n6674), .ZN(n6568) );
  NAND2_X1 U7477 ( .A1(n6569), .A2(n6568), .ZN(n6574) );
  NAND3_X1 U7478 ( .A1(n6572), .A2(n6571), .A3(n6570), .ZN(n6573) );
  OAI21_X1 U7479 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6673), .A(n6662), .ZN(
        n6586) );
  AOI221_X1 U7480 ( .B1(n6576), .B2(STATE2_REG_0__SCAN_IN), .C1(n6586), .C2(
        STATE2_REG_0__SCAN_IN), .A(n6575), .ZN(n6580) );
  OAI211_X1 U7481 ( .C1(n6578), .C2(n6577), .A(n6585), .B(n6662), .ZN(n6579)
         );
  OAI211_X1 U7482 ( .C1(n6582), .C2(n6581), .A(n6580), .B(n6579), .ZN(U3148)
         );
  AOI21_X1 U7483 ( .B1(n6584), .B2(n6673), .A(n6583), .ZN(n6589) );
  NAND2_X1 U7484 ( .A1(n6585), .A2(n6480), .ZN(n6592) );
  NAND3_X1 U7485 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6592), .A3(n6586), .ZN(
        n6587) );
  OAI211_X1 U7486 ( .C1(n6590), .C2(n6589), .A(n6588), .B(n6587), .ZN(U3149)
         );
  INV_X1 U7487 ( .A(n6591), .ZN(n6660) );
  OAI211_X1 U7488 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6673), .A(n6660), .B(
        n6592), .ZN(n6594) );
  OAI21_X1 U7489 ( .B1(n6677), .B2(n6594), .A(n6593), .ZN(U3150) );
  INV_X1 U7490 ( .A(n6659), .ZN(n6595) );
  AND2_X1 U7491 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6595), .ZN(U3151) );
  AND2_X1 U7492 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6595), .ZN(U3152) );
  AND2_X1 U7493 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6595), .ZN(U3153) );
  AND2_X1 U7494 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6595), .ZN(U3154) );
  AND2_X1 U7495 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6595), .ZN(U3155) );
  AND2_X1 U7496 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6595), .ZN(U3156) );
  AND2_X1 U7497 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6595), .ZN(U3157) );
  AND2_X1 U7498 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6595), .ZN(U3158) );
  AND2_X1 U7499 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6595), .ZN(U3159) );
  AND2_X1 U7500 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6595), .ZN(U3160) );
  AND2_X1 U7501 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6595), .ZN(U3161) );
  AND2_X1 U7502 ( .A1(n6595), .A2(DATAWIDTH_REG_20__SCAN_IN), .ZN(U3162) );
  AND2_X1 U7503 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6595), .ZN(U3163) );
  AND2_X1 U7504 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6595), .ZN(U3164) );
  AND2_X1 U7505 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6595), .ZN(U3165) );
  AND2_X1 U7506 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6595), .ZN(U3166) );
  AND2_X1 U7507 ( .A1(n6595), .A2(DATAWIDTH_REG_15__SCAN_IN), .ZN(U3167) );
  AND2_X1 U7508 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6595), .ZN(U3168) );
  AND2_X1 U7509 ( .A1(n6595), .A2(DATAWIDTH_REG_13__SCAN_IN), .ZN(U3169) );
  AND2_X1 U7510 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6595), .ZN(U3170) );
  AND2_X1 U7511 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6595), .ZN(U3171) );
  AND2_X1 U7512 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6595), .ZN(U3172) );
  AND2_X1 U7513 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6595), .ZN(U3173) );
  INV_X1 U7514 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6857) );
  NOR2_X1 U7515 ( .A1(n6659), .A2(n6857), .ZN(U3174) );
  AND2_X1 U7516 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6595), .ZN(U3175) );
  AND2_X1 U7517 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6595), .ZN(U3176) );
  AND2_X1 U7518 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6595), .ZN(U3177) );
  AND2_X1 U7519 ( .A1(n6595), .A2(DATAWIDTH_REG_4__SCAN_IN), .ZN(U3178) );
  AND2_X1 U7520 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6595), .ZN(U3179) );
  AND2_X1 U7521 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6595), .ZN(U3180) );
  NOR2_X1 U7522 ( .A1(n6602), .A2(n6612), .ZN(n6603) );
  AOI22_X1 U7523 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6611) );
  AND2_X1 U7524 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6599) );
  INV_X1 U7525 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6597) );
  INV_X1 U7526 ( .A(NA_N), .ZN(n6604) );
  AOI221_X1 U7527 ( .B1(STATE_REG_1__SCAN_IN), .B2(STATE_REG_2__SCAN_IN), .C1(
        n6604), .C2(STATE_REG_2__SCAN_IN), .A(STATE_REG_0__SCAN_IN), .ZN(n6608) );
  AOI221_X1 U7528 ( .B1(n6599), .B2(n6682), .C1(n6597), .C2(n6682), .A(n6608), 
        .ZN(n6596) );
  OAI21_X1 U7529 ( .B1(n6603), .B2(n6611), .A(n6596), .ZN(U3181) );
  NOR2_X1 U7530 ( .A1(n6606), .A2(n6597), .ZN(n6605) );
  NAND2_X1 U7531 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6598) );
  OAI21_X1 U7532 ( .B1(n6605), .B2(n6599), .A(n6598), .ZN(n6600) );
  OAI211_X1 U7533 ( .C1(n6602), .C2(n6673), .A(n6601), .B(n6600), .ZN(U3182)
         );
  AOI21_X1 U7534 ( .B1(n6605), .B2(n6604), .A(n6603), .ZN(n6610) );
  AOI221_X1 U7535 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6673), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6607) );
  AOI221_X1 U7536 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6607), .C2(HOLD), .A(n6606), .ZN(n6609) );
  OAI22_X1 U7537 ( .A1(n6611), .A2(n6610), .B1(n6609), .B2(n6608), .ZN(U3183)
         );
  NAND2_X1 U7538 ( .A1(n6612), .A2(n6613), .ZN(n6653) );
  NAND2_X1 U7539 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6613), .ZN(n6655) );
  INV_X1 U7540 ( .A(n6655), .ZN(n7003) );
  AOI22_X1 U7541 ( .A1(REIP_REG_2__SCAN_IN), .A2(n7003), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6682), .ZN(n6614) );
  OAI21_X1 U7542 ( .B1(n6615), .B2(n6653), .A(n6614), .ZN(U3185) );
  AOI22_X1 U7543 ( .A1(REIP_REG_3__SCAN_IN), .A2(n7003), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6682), .ZN(n6616) );
  OAI21_X1 U7544 ( .B1(n6617), .B2(n6653), .A(n6616), .ZN(U3186) );
  AOI22_X1 U7545 ( .A1(REIP_REG_4__SCAN_IN), .A2(n7003), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6682), .ZN(n6618) );
  OAI21_X1 U7546 ( .B1(n6620), .B2(n6653), .A(n6618), .ZN(U3187) );
  INV_X1 U7547 ( .A(n6653), .ZN(n7004) );
  AOI22_X1 U7548 ( .A1(REIP_REG_6__SCAN_IN), .A2(n7004), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6682), .ZN(n6619) );
  OAI21_X1 U7549 ( .B1(n6620), .B2(n6655), .A(n6619), .ZN(U3188) );
  AOI22_X1 U7550 ( .A1(REIP_REG_6__SCAN_IN), .A2(n7003), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6682), .ZN(n6621) );
  OAI21_X1 U7551 ( .B1(n6623), .B2(n6653), .A(n6621), .ZN(U3189) );
  AOI22_X1 U7552 ( .A1(REIP_REG_8__SCAN_IN), .A2(n7004), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6682), .ZN(n6622) );
  OAI21_X1 U7553 ( .B1(n6623), .B2(n6655), .A(n6622), .ZN(U3190) );
  AOI22_X1 U7554 ( .A1(REIP_REG_8__SCAN_IN), .A2(n7003), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6682), .ZN(n6624) );
  OAI21_X1 U7555 ( .B1(n6626), .B2(n6653), .A(n6624), .ZN(U3191) );
  AOI22_X1 U7556 ( .A1(REIP_REG_10__SCAN_IN), .A2(n7004), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6682), .ZN(n6625) );
  OAI21_X1 U7557 ( .B1(n6626), .B2(n6655), .A(n6625), .ZN(U3192) );
  AOI22_X1 U7558 ( .A1(REIP_REG_10__SCAN_IN), .A2(n7003), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6682), .ZN(n6627) );
  OAI21_X1 U7559 ( .B1(n6629), .B2(n6653), .A(n6627), .ZN(U3193) );
  AOI22_X1 U7560 ( .A1(REIP_REG_12__SCAN_IN), .A2(n7004), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6682), .ZN(n6628) );
  OAI21_X1 U7561 ( .B1(n6629), .B2(n6655), .A(n6628), .ZN(U3194) );
  AOI22_X1 U7562 ( .A1(REIP_REG_13__SCAN_IN), .A2(n7004), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6682), .ZN(n6630) );
  OAI21_X1 U7563 ( .B1(n5229), .B2(n6655), .A(n6630), .ZN(U3195) );
  AOI222_X1 U7564 ( .A1(n7003), .A2(REIP_REG_13__SCAN_IN), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6682), .C1(REIP_REG_14__SCAN_IN), .C2(
        n7004), .ZN(n6631) );
  INV_X1 U7565 ( .A(n6631), .ZN(U3196) );
  AOI22_X1 U7566 ( .A1(REIP_REG_15__SCAN_IN), .A2(n7004), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6682), .ZN(n6632) );
  OAI21_X1 U7567 ( .B1(n5589), .B2(n6655), .A(n6632), .ZN(U3197) );
  AOI22_X1 U7568 ( .A1(REIP_REG_16__SCAN_IN), .A2(n7004), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6682), .ZN(n6633) );
  OAI21_X1 U7569 ( .B1(n6634), .B2(n6655), .A(n6633), .ZN(U3198) );
  AOI22_X1 U7570 ( .A1(REIP_REG_16__SCAN_IN), .A2(n7003), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6682), .ZN(n6635) );
  OAI21_X1 U7571 ( .B1(n6636), .B2(n6653), .A(n6635), .ZN(U3199) );
  AOI222_X1 U7572 ( .A1(n7004), .A2(REIP_REG_18__SCAN_IN), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6682), .C1(REIP_REG_17__SCAN_IN), .C2(
        n7003), .ZN(n6637) );
  INV_X1 U7573 ( .A(n6637), .ZN(U3200) );
  AOI222_X1 U7574 ( .A1(n7004), .A2(REIP_REG_19__SCAN_IN), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6682), .C1(REIP_REG_18__SCAN_IN), .C2(
        n7003), .ZN(n6638) );
  INV_X1 U7575 ( .A(n6638), .ZN(U3201) );
  AOI22_X1 U7576 ( .A1(REIP_REG_19__SCAN_IN), .A2(n7003), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6682), .ZN(n6639) );
  OAI21_X1 U7577 ( .B1(n6641), .B2(n6653), .A(n6639), .ZN(U3202) );
  AOI22_X1 U7578 ( .A1(REIP_REG_21__SCAN_IN), .A2(n7004), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6682), .ZN(n6640) );
  OAI21_X1 U7579 ( .B1(n6641), .B2(n6655), .A(n6640), .ZN(U3203) );
  AOI222_X1 U7580 ( .A1(n7003), .A2(REIP_REG_21__SCAN_IN), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6682), .C1(REIP_REG_22__SCAN_IN), .C2(
        n7004), .ZN(n6642) );
  INV_X1 U7581 ( .A(n6642), .ZN(U3204) );
  INV_X1 U7582 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6644) );
  AOI22_X1 U7583 ( .A1(REIP_REG_23__SCAN_IN), .A2(n7004), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6682), .ZN(n6643) );
  OAI21_X1 U7584 ( .B1(n6644), .B2(n6655), .A(n6643), .ZN(U3205) );
  AOI22_X1 U7585 ( .A1(REIP_REG_23__SCAN_IN), .A2(n7003), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6682), .ZN(n6645) );
  OAI21_X1 U7586 ( .B1(n5527), .B2(n6653), .A(n6645), .ZN(U3206) );
  AOI22_X1 U7587 ( .A1(REIP_REG_24__SCAN_IN), .A2(n7003), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6682), .ZN(n6646) );
  OAI21_X1 U7588 ( .B1(n6647), .B2(n6653), .A(n6646), .ZN(U3207) );
  AOI22_X1 U7589 ( .A1(REIP_REG_25__SCAN_IN), .A2(n7003), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6682), .ZN(n6648) );
  OAI21_X1 U7590 ( .B1(n6869), .B2(n6653), .A(n6648), .ZN(U3208) );
  AOI222_X1 U7591 ( .A1(n7003), .A2(REIP_REG_26__SCAN_IN), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6682), .C1(REIP_REG_27__SCAN_IN), .C2(
        n7004), .ZN(n6649) );
  INV_X1 U7592 ( .A(n6649), .ZN(U3209) );
  AOI22_X1 U7593 ( .A1(REIP_REG_27__SCAN_IN), .A2(n7003), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6682), .ZN(n6650) );
  OAI21_X1 U7594 ( .B1(n6859), .B2(n6653), .A(n6650), .ZN(U3210) );
  AOI22_X1 U7595 ( .A1(REIP_REG_29__SCAN_IN), .A2(n7004), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6682), .ZN(n6651) );
  OAI21_X1 U7596 ( .B1(n6859), .B2(n6655), .A(n6651), .ZN(U3211) );
  AOI22_X1 U7597 ( .A1(REIP_REG_29__SCAN_IN), .A2(n7003), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6682), .ZN(n6652) );
  OAI21_X1 U7598 ( .B1(n4161), .B2(n6653), .A(n6652), .ZN(U3212) );
  AOI22_X1 U7599 ( .A1(REIP_REG_31__SCAN_IN), .A2(n7004), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6682), .ZN(n6654) );
  OAI21_X1 U7600 ( .B1(n4161), .B2(n6655), .A(n6654), .ZN(U3213) );
  MUX2_X1 U7601 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6682), .Z(U3445) );
  MUX2_X1 U7602 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6682), .Z(U3446) );
  MUX2_X1 U7603 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6682), .Z(U3447) );
  MUX2_X1 U7604 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6682), .Z(U3448) );
  OAI21_X1 U7605 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6659), .A(n6657), .ZN(
        n6656) );
  INV_X1 U7606 ( .A(n6656), .ZN(U3451) );
  OAI21_X1 U7607 ( .B1(n6659), .B2(n6658), .A(n6657), .ZN(U3452) );
  OAI211_X1 U7608 ( .C1(n6663), .C2(n6662), .A(n6661), .B(n6660), .ZN(U3453)
         );
  INV_X1 U7609 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6666) );
  AOI21_X1 U7610 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6664) );
  OAI221_X1 U7611 ( .B1(REIP_REG_1__SCAN_IN), .B2(n6664), .C1(n5096), .C2(
        REIP_REG_0__SCAN_IN), .A(n6669), .ZN(n6665) );
  OAI21_X1 U7612 ( .B1(n6669), .B2(n6666), .A(n6665), .ZN(U3468) );
  INV_X1 U7613 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6668) );
  OAI21_X1 U7614 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6669), .ZN(n6667) );
  OAI21_X1 U7615 ( .B1(n6669), .B2(n6668), .A(n6667), .ZN(U3469) );
  NAND2_X1 U7616 ( .A1(n6682), .A2(W_R_N_REG_SCAN_IN), .ZN(n6670) );
  OAI21_X1 U7617 ( .B1(n6682), .B2(READREQUEST_REG_SCAN_IN), .A(n6670), .ZN(
        U3470) );
  AOI211_X1 U7618 ( .C1(n6674), .C2(n6673), .A(n6672), .B(n6671), .ZN(n6681)
         );
  OAI211_X1 U7619 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6676), .A(n6675), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6678) );
  AOI21_X1 U7620 ( .B1(n6678), .B2(STATE2_REG_0__SCAN_IN), .A(n6677), .ZN(
        n6680) );
  NAND2_X1 U7621 ( .A1(n6681), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6679) );
  OAI21_X1 U7622 ( .B1(n6681), .B2(n6680), .A(n6679), .ZN(U3472) );
  MUX2_X1 U7623 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6682), .Z(U3473) );
  INV_X1 U7624 ( .A(keyinput95), .ZN(n6683) );
  NAND4_X1 U7625 ( .A1(keyinput83), .A2(keyinput16), .A3(keyinput68), .A4(
        n6683), .ZN(n6684) );
  NOR4_X1 U7626 ( .A1(keyinput88), .A2(keyinput105), .A3(keyinput38), .A4(
        n6684), .ZN(n6695) );
  NOR4_X1 U7627 ( .A1(keyinput10), .A2(keyinput63), .A3(keyinput26), .A4(
        keyinput56), .ZN(n6694) );
  NAND2_X1 U7628 ( .A1(keyinput125), .A2(keyinput108), .ZN(n6685) );
  NOR3_X1 U7629 ( .A1(keyinput92), .A2(keyinput5), .A3(n6685), .ZN(n6693) );
  NAND4_X1 U7630 ( .A1(keyinput47), .A2(keyinput53), .A3(keyinput127), .A4(
        keyinput33), .ZN(n6691) );
  NAND4_X1 U7631 ( .A1(keyinput112), .A2(keyinput30), .A3(keyinput113), .A4(
        keyinput6), .ZN(n6690) );
  NOR2_X1 U7632 ( .A1(keyinput67), .A2(keyinput49), .ZN(n6686) );
  NAND3_X1 U7633 ( .A1(keyinput100), .A2(keyinput65), .A3(n6686), .ZN(n6689)
         );
  INV_X1 U7634 ( .A(keyinput54), .ZN(n6687) );
  NAND4_X1 U7635 ( .A1(keyinput69), .A2(keyinput103), .A3(keyinput57), .A4(
        n6687), .ZN(n6688) );
  NOR4_X1 U7636 ( .A1(n6691), .A2(n6690), .A3(n6689), .A4(n6688), .ZN(n6692)
         );
  NAND4_X1 U7637 ( .A1(n6695), .A2(n6694), .A3(n6693), .A4(n6692), .ZN(n6744)
         );
  NAND3_X1 U7638 ( .A1(keyinput82), .A2(keyinput22), .A3(keyinput96), .ZN(
        n6696) );
  NOR2_X1 U7639 ( .A1(keyinput76), .A2(n6696), .ZN(n6742) );
  INV_X1 U7640 ( .A(keyinput41), .ZN(n6917) );
  NOR4_X1 U7641 ( .A1(keyinput37), .A2(keyinput122), .A3(keyinput1), .A4(n6917), .ZN(n6741) );
  NAND2_X1 U7642 ( .A1(keyinput11), .A2(keyinput109), .ZN(n6697) );
  NOR3_X1 U7643 ( .A1(keyinput115), .A2(keyinput124), .A3(n6697), .ZN(n6698)
         );
  NAND3_X1 U7644 ( .A1(keyinput73), .A2(keyinput94), .A3(n6698), .ZN(n6706) );
  NAND2_X1 U7645 ( .A1(keyinput50), .A2(keyinput77), .ZN(n6699) );
  NOR3_X1 U7646 ( .A1(keyinput75), .A2(keyinput120), .A3(n6699), .ZN(n6704) );
  NOR4_X1 U7647 ( .A1(keyinput14), .A2(keyinput45), .A3(keyinput36), .A4(
        keyinput106), .ZN(n6703) );
  NAND3_X1 U7648 ( .A1(keyinput60), .A2(keyinput102), .A3(keyinput15), .ZN(
        n6700) );
  NOR2_X1 U7649 ( .A1(keyinput8), .A2(n6700), .ZN(n6702) );
  NOR4_X1 U7650 ( .A1(keyinput17), .A2(keyinput81), .A3(keyinput87), .A4(
        keyinput31), .ZN(n6701) );
  NAND4_X1 U7651 ( .A1(n6704), .A2(n6703), .A3(n6702), .A4(n6701), .ZN(n6705)
         );
  NOR4_X1 U7652 ( .A1(keyinput52), .A2(keyinput29), .A3(n6706), .A4(n6705), 
        .ZN(n6740) );
  NOR2_X1 U7653 ( .A1(keyinput114), .A2(keyinput119), .ZN(n6707) );
  NAND3_X1 U7654 ( .A1(keyinput34), .A2(keyinput39), .A3(n6707), .ZN(n6708) );
  NOR3_X1 U7655 ( .A1(keyinput71), .A2(keyinput101), .A3(n6708), .ZN(n6720) );
  NAND2_X1 U7656 ( .A1(keyinput12), .A2(keyinput104), .ZN(n6709) );
  NOR3_X1 U7657 ( .A1(keyinput78), .A2(keyinput116), .A3(n6709), .ZN(n6710) );
  NAND3_X1 U7658 ( .A1(keyinput4), .A2(keyinput64), .A3(n6710), .ZN(n6718) );
  NOR4_X1 U7659 ( .A1(keyinput13), .A2(keyinput123), .A3(keyinput18), .A4(
        keyinput61), .ZN(n6716) );
  NAND3_X1 U7660 ( .A1(keyinput86), .A2(keyinput118), .A3(keyinput25), .ZN(
        n6711) );
  NOR2_X1 U7661 ( .A1(keyinput24), .A2(n6711), .ZN(n6715) );
  NAND3_X1 U7662 ( .A1(keyinput93), .A2(keyinput58), .A3(keyinput99), .ZN(
        n6712) );
  NOR2_X1 U7663 ( .A1(keyinput74), .A2(n6712), .ZN(n6714) );
  INV_X1 U7664 ( .A(keyinput98), .ZN(n6853) );
  NOR4_X1 U7665 ( .A1(keyinput51), .A2(keyinput126), .A3(keyinput62), .A4(
        n6853), .ZN(n6713) );
  NAND4_X1 U7666 ( .A1(n6716), .A2(n6715), .A3(n6714), .A4(n6713), .ZN(n6717)
         );
  NOR4_X1 U7667 ( .A1(keyinput27), .A2(keyinput9), .A3(n6718), .A4(n6717), 
        .ZN(n6719) );
  NAND4_X1 U7668 ( .A1(keyinput32), .A2(keyinput35), .A3(n6720), .A4(n6719), 
        .ZN(n6738) );
  NOR2_X1 U7669 ( .A1(keyinput48), .A2(keyinput66), .ZN(n6721) );
  NAND3_X1 U7670 ( .A1(keyinput2), .A2(keyinput72), .A3(n6721), .ZN(n6737) );
  INV_X1 U7671 ( .A(keyinput59), .ZN(n6722) );
  NAND4_X1 U7672 ( .A1(keyinput91), .A2(keyinput21), .A3(keyinput23), .A4(
        n6722), .ZN(n6736) );
  INV_X1 U7673 ( .A(keyinput80), .ZN(n6723) );
  NOR4_X1 U7674 ( .A1(keyinput70), .A2(keyinput90), .A3(keyinput55), .A4(n6723), .ZN(n6734) );
  NAND2_X1 U7675 ( .A1(keyinput3), .A2(keyinput46), .ZN(n6724) );
  NOR3_X1 U7676 ( .A1(keyinput7), .A2(keyinput85), .A3(n6724), .ZN(n6733) );
  INV_X1 U7677 ( .A(keyinput110), .ZN(n6725) );
  NAND4_X1 U7678 ( .A1(keyinput19), .A2(keyinput43), .A3(keyinput79), .A4(
        n6725), .ZN(n6731) );
  NOR2_X1 U7679 ( .A1(keyinput40), .A2(keyinput89), .ZN(n6726) );
  NAND3_X1 U7680 ( .A1(keyinput107), .A2(keyinput121), .A3(n6726), .ZN(n6730)
         );
  NAND4_X1 U7681 ( .A1(keyinput117), .A2(keyinput44), .A3(keyinput111), .A4(
        keyinput42), .ZN(n6729) );
  NOR2_X1 U7682 ( .A1(keyinput97), .A2(keyinput28), .ZN(n6727) );
  NAND3_X1 U7683 ( .A1(keyinput84), .A2(keyinput0), .A3(n6727), .ZN(n6728) );
  NOR4_X1 U7684 ( .A1(n6731), .A2(n6730), .A3(n6729), .A4(n6728), .ZN(n6732)
         );
  NAND3_X1 U7685 ( .A1(n6734), .A2(n6733), .A3(n6732), .ZN(n6735) );
  NOR4_X1 U7686 ( .A1(n6738), .A2(n6737), .A3(n6736), .A4(n6735), .ZN(n6739)
         );
  NAND4_X1 U7687 ( .A1(n6742), .A2(n6741), .A3(n6740), .A4(n6739), .ZN(n6743)
         );
  OAI21_X1 U7688 ( .B1(n6744), .B2(n6743), .A(keyinput20), .ZN(n7002) );
  INV_X1 U7689 ( .A(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n6747) );
  INV_X1 U7690 ( .A(keyinput91), .ZN(n6746) );
  AOI22_X1 U7691 ( .A1(n6747), .A2(keyinput59), .B1(DATAO_REG_9__SCAN_IN), 
        .B2(n6746), .ZN(n6745) );
  OAI221_X1 U7692 ( .B1(n6747), .B2(keyinput59), .C1(n6746), .C2(
        DATAO_REG_9__SCAN_IN), .A(n6745), .ZN(n6758) );
  AOI22_X1 U7693 ( .A1(n6750), .A2(keyinput23), .B1(n6749), .B2(keyinput48), 
        .ZN(n6748) );
  OAI221_X1 U7694 ( .B1(n6750), .B2(keyinput23), .C1(n6749), .C2(keyinput48), 
        .A(n6748), .ZN(n6757) );
  INV_X1 U7695 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n6753) );
  INV_X1 U7696 ( .A(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n6752) );
  AOI22_X1 U7697 ( .A1(n6753), .A2(keyinput2), .B1(keyinput66), .B2(n6752), 
        .ZN(n6751) );
  OAI221_X1 U7698 ( .B1(n6753), .B2(keyinput2), .C1(n6752), .C2(keyinput66), 
        .A(n6751), .ZN(n6756) );
  AOI22_X1 U7699 ( .A1(n5872), .A2(keyinput72), .B1(keyinput40), .B2(n4161), 
        .ZN(n6754) );
  OAI221_X1 U7700 ( .B1(n5872), .B2(keyinput72), .C1(n4161), .C2(keyinput40), 
        .A(n6754), .ZN(n6755) );
  NOR4_X1 U7701 ( .A1(n6758), .A2(n6757), .A3(n6756), .A4(n6755), .ZN(n6807)
         );
  INV_X1 U7702 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n6760) );
  AOI22_X1 U7703 ( .A1(n6761), .A2(keyinput110), .B1(keyinput43), .B2(n6760), 
        .ZN(n6759) );
  OAI221_X1 U7704 ( .B1(n6761), .B2(keyinput110), .C1(n6760), .C2(keyinput43), 
        .A(n6759), .ZN(n6774) );
  INV_X1 U7705 ( .A(DATAI_27_), .ZN(n6764) );
  INV_X1 U7706 ( .A(keyinput107), .ZN(n6763) );
  AOI22_X1 U7707 ( .A1(n6764), .A2(keyinput121), .B1(DATAO_REG_18__SCAN_IN), 
        .B2(n6763), .ZN(n6762) );
  OAI221_X1 U7708 ( .B1(n6764), .B2(keyinput121), .C1(n6763), .C2(
        DATAO_REG_18__SCAN_IN), .A(n6762), .ZN(n6773) );
  INV_X1 U7709 ( .A(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n6766) );
  AOI22_X1 U7710 ( .A1(n6767), .A2(keyinput89), .B1(n6766), .B2(keyinput19), 
        .ZN(n6765) );
  OAI221_X1 U7711 ( .B1(n6767), .B2(keyinput89), .C1(n6766), .C2(keyinput19), 
        .A(n6765), .ZN(n6772) );
  INV_X1 U7712 ( .A(DATAI_8_), .ZN(n6768) );
  XOR2_X1 U7713 ( .A(n6768), .B(keyinput84), .Z(n6770) );
  XNOR2_X1 U7714 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput79), .ZN(
        n6769) );
  NAND2_X1 U7715 ( .A1(n6770), .A2(n6769), .ZN(n6771) );
  NOR4_X1 U7716 ( .A1(n6774), .A2(n6773), .A3(n6772), .A4(n6771), .ZN(n6806)
         );
  INV_X1 U7717 ( .A(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n6777) );
  AOI22_X1 U7718 ( .A1(n6777), .A2(keyinput97), .B1(keyinput117), .B2(n6776), 
        .ZN(n6775) );
  OAI221_X1 U7719 ( .B1(n6777), .B2(keyinput97), .C1(n6776), .C2(keyinput117), 
        .A(n6775), .ZN(n6789) );
  INV_X1 U7720 ( .A(keyinput44), .ZN(n6780) );
  INV_X1 U7721 ( .A(keyinput0), .ZN(n6779) );
  AOI22_X1 U7722 ( .A1(n6780), .A2(ADDRESS_REG_20__SCAN_IN), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6779), .ZN(n6778) );
  OAI221_X1 U7723 ( .B1(n6780), .B2(ADDRESS_REG_20__SCAN_IN), .C1(n6779), .C2(
        ADDRESS_REG_16__SCAN_IN), .A(n6778), .ZN(n6788) );
  INV_X1 U7724 ( .A(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n6783) );
  INV_X1 U7725 ( .A(DATAI_26_), .ZN(n6782) );
  AOI22_X1 U7726 ( .A1(n6783), .A2(keyinput28), .B1(keyinput111), .B2(n6782), 
        .ZN(n6781) );
  OAI221_X1 U7727 ( .B1(n6783), .B2(keyinput28), .C1(n6782), .C2(keyinput111), 
        .A(n6781), .ZN(n6787) );
  INV_X1 U7728 ( .A(keyinput42), .ZN(n6785) );
  AOI22_X1 U7729 ( .A1(n4355), .A2(keyinput7), .B1(ADDRESS_REG_1__SCAN_IN), 
        .B2(n6785), .ZN(n6784) );
  OAI221_X1 U7730 ( .B1(n4355), .B2(keyinput7), .C1(n6785), .C2(
        ADDRESS_REG_1__SCAN_IN), .A(n6784), .ZN(n6786) );
  NOR4_X1 U7731 ( .A1(n6789), .A2(n6788), .A3(n6787), .A4(n6786), .ZN(n6805)
         );
  AOI22_X1 U7732 ( .A1(n5406), .A2(keyinput46), .B1(keyinput3), .B2(n6791), 
        .ZN(n6790) );
  OAI221_X1 U7733 ( .B1(n5406), .B2(keyinput46), .C1(n6791), .C2(keyinput3), 
        .A(n6790), .ZN(n6803) );
  INV_X1 U7734 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n6794) );
  INV_X1 U7735 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n6793) );
  AOI22_X1 U7736 ( .A1(n6794), .A2(keyinput85), .B1(keyinput70), .B2(n6793), 
        .ZN(n6792) );
  OAI221_X1 U7737 ( .B1(n6794), .B2(keyinput85), .C1(n6793), .C2(keyinput70), 
        .A(n6792), .ZN(n6802) );
  INV_X1 U7738 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6797) );
  INV_X1 U7739 ( .A(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n6796) );
  AOI22_X1 U7740 ( .A1(n6797), .A2(keyinput80), .B1(n6796), .B2(keyinput90), 
        .ZN(n6795) );
  OAI221_X1 U7741 ( .B1(n6797), .B2(keyinput80), .C1(n6796), .C2(keyinput90), 
        .A(n6795), .ZN(n6801) );
  AOI22_X1 U7742 ( .A1(n5096), .A2(keyinput88), .B1(n6799), .B2(keyinput55), 
        .ZN(n6798) );
  OAI221_X1 U7743 ( .B1(n5096), .B2(keyinput88), .C1(n6799), .C2(keyinput55), 
        .A(n6798), .ZN(n6800) );
  NOR4_X1 U7744 ( .A1(n6803), .A2(n6802), .A3(n6801), .A4(n6800), .ZN(n6804)
         );
  NAND4_X1 U7745 ( .A1(n6807), .A2(n6806), .A3(n6805), .A4(n6804), .ZN(n7001)
         );
  INV_X1 U7746 ( .A(LWORD_REG_8__SCAN_IN), .ZN(n6810) );
  AOI22_X1 U7747 ( .A1(n6810), .A2(keyinput34), .B1(n6809), .B2(keyinput32), 
        .ZN(n6808) );
  OAI221_X1 U7748 ( .B1(n6810), .B2(keyinput34), .C1(n6809), .C2(keyinput32), 
        .A(n6808), .ZN(n6822) );
  INV_X1 U7749 ( .A(DATAI_18_), .ZN(n6813) );
  INV_X1 U7750 ( .A(keyinput71), .ZN(n6812) );
  AOI22_X1 U7751 ( .A1(n6813), .A2(keyinput35), .B1(HOLD), .B2(n6812), .ZN(
        n6811) );
  OAI221_X1 U7752 ( .B1(n6813), .B2(keyinput35), .C1(n6812), .C2(HOLD), .A(
        n6811), .ZN(n6821) );
  INV_X1 U7753 ( .A(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n6815) );
  AOI22_X1 U7754 ( .A1(n5884), .A2(keyinput101), .B1(keyinput119), .B2(n6815), 
        .ZN(n6814) );
  OAI221_X1 U7755 ( .B1(n5884), .B2(keyinput101), .C1(n6815), .C2(keyinput119), 
        .A(n6814), .ZN(n6820) );
  INV_X1 U7756 ( .A(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n6817) );
  AOI22_X1 U7757 ( .A1(n6818), .A2(keyinput39), .B1(n6817), .B2(keyinput118), 
        .ZN(n6816) );
  OAI221_X1 U7758 ( .B1(n6818), .B2(keyinput39), .C1(n6817), .C2(keyinput118), 
        .A(n6816), .ZN(n6819) );
  NOR4_X1 U7759 ( .A1(n6822), .A2(n6821), .A3(n6820), .A4(n6819), .ZN(n6999)
         );
  INV_X1 U7760 ( .A(keyinput25), .ZN(n6824) );
  AOI22_X1 U7761 ( .A1(n6825), .A2(keyinput13), .B1(DATAO_REG_27__SCAN_IN), 
        .B2(n6824), .ZN(n6823) );
  OAI221_X1 U7762 ( .B1(n6825), .B2(keyinput13), .C1(n6824), .C2(
        DATAO_REG_27__SCAN_IN), .A(n6823), .ZN(n6836) );
  AOI22_X1 U7763 ( .A1(n5439), .A2(keyinput123), .B1(keyinput18), .B2(n3787), 
        .ZN(n6826) );
  OAI221_X1 U7764 ( .B1(n5439), .B2(keyinput123), .C1(n3787), .C2(keyinput18), 
        .A(n6826), .ZN(n6835) );
  INV_X1 U7765 ( .A(DATAI_13_), .ZN(n6828) );
  AOI22_X1 U7766 ( .A1(n6829), .A2(keyinput61), .B1(keyinput24), .B2(n6828), 
        .ZN(n6827) );
  OAI221_X1 U7767 ( .B1(n6829), .B2(keyinput61), .C1(n6828), .C2(keyinput24), 
        .A(n6827), .ZN(n6834) );
  INV_X1 U7768 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n6832) );
  INV_X1 U7769 ( .A(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n6831) );
  AOI22_X1 U7770 ( .A1(n6832), .A2(keyinput86), .B1(n6831), .B2(keyinput4), 
        .ZN(n6830) );
  OAI221_X1 U7771 ( .B1(n6832), .B2(keyinput86), .C1(n6831), .C2(keyinput4), 
        .A(n6830), .ZN(n6833) );
  NOR4_X1 U7772 ( .A1(n6836), .A2(n6835), .A3(n6834), .A4(n6833), .ZN(n6998)
         );
  AOI22_X1 U7773 ( .A1(n6838), .A2(keyinput9), .B1(n3576), .B2(keyinput51), 
        .ZN(n6837) );
  OAI221_X1 U7774 ( .B1(n6838), .B2(keyinput9), .C1(n3576), .C2(keyinput51), 
        .A(n6837), .ZN(n6867) );
  INV_X1 U7775 ( .A(keyinput64), .ZN(n6841) );
  INV_X1 U7776 ( .A(keyinput78), .ZN(n6840) );
  OAI22_X1 U7777 ( .A1(n6841), .A2(ADDRESS_REG_12__SCAN_IN), .B1(n6840), .B2(
        DATAWIDTH_REG_15__SCAN_IN), .ZN(n6839) );
  AOI221_X1 U7778 ( .B1(n6841), .B2(ADDRESS_REG_12__SCAN_IN), .C1(
        DATAWIDTH_REG_15__SCAN_IN), .C2(n6840), .A(n6839), .ZN(n6849) );
  INV_X1 U7779 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n6844) );
  INV_X1 U7780 ( .A(UWORD_REG_9__SCAN_IN), .ZN(n6843) );
  OAI22_X1 U7781 ( .A1(n6844), .A2(keyinput104), .B1(n6843), .B2(keyinput116), 
        .ZN(n6842) );
  AOI221_X1 U7782 ( .B1(n6844), .B2(keyinput104), .C1(keyinput116), .C2(n6843), 
        .A(n6842), .ZN(n6848) );
  INV_X1 U7783 ( .A(keyinput12), .ZN(n6846) );
  OAI22_X1 U7784 ( .A1(n5589), .A2(keyinput27), .B1(n6846), .B2(
        ADDRESS_REG_22__SCAN_IN), .ZN(n6845) );
  AOI221_X1 U7785 ( .B1(n5589), .B2(keyinput27), .C1(ADDRESS_REG_22__SCAN_IN), 
        .C2(n6846), .A(n6845), .ZN(n6847) );
  NAND3_X1 U7786 ( .A1(n6849), .A2(n6848), .A3(n6847), .ZN(n6866) );
  AOI22_X1 U7787 ( .A1(n5108), .A2(keyinput62), .B1(n6851), .B2(keyinput58), 
        .ZN(n6850) );
  OAI221_X1 U7788 ( .B1(n5108), .B2(keyinput62), .C1(n6851), .C2(keyinput58), 
        .A(n6850), .ZN(n6865) );
  OAI22_X1 U7789 ( .A1(n6854), .A2(keyinput126), .B1(n6853), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6852) );
  AOI221_X1 U7790 ( .B1(n6854), .B2(keyinput126), .C1(DATAO_REG_10__SCAN_IN), 
        .C2(n6853), .A(n6852), .ZN(n6863) );
  INV_X1 U7791 ( .A(keyinput74), .ZN(n6856) );
  OAI22_X1 U7792 ( .A1(keyinput99), .A2(n6857), .B1(n6856), .B2(
        ADDRESS_REG_21__SCAN_IN), .ZN(n6855) );
  AOI221_X1 U7793 ( .B1(n6857), .B2(keyinput99), .C1(n6856), .C2(
        ADDRESS_REG_21__SCAN_IN), .A(n6855), .ZN(n6862) );
  OAI22_X1 U7794 ( .A1(n6860), .A2(keyinput93), .B1(n6859), .B2(keyinput21), 
        .ZN(n6858) );
  AOI221_X1 U7795 ( .B1(n6860), .B2(keyinput93), .C1(keyinput21), .C2(n6859), 
        .A(n6858), .ZN(n6861) );
  NAND3_X1 U7796 ( .A1(n6863), .A2(n6862), .A3(n6861), .ZN(n6864) );
  NOR4_X1 U7797 ( .A1(n6867), .A2(n6866), .A3(n6865), .A4(n6864), .ZN(n6997)
         );
  INV_X1 U7798 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n6873) );
  XOR2_X1 U7799 ( .A(EBX_REG_20__SCAN_IN), .B(keyinput105), .Z(n6872) );
  INV_X1 U7800 ( .A(DATAI_16_), .ZN(n6870) );
  AOI22_X1 U7801 ( .A1(n6870), .A2(keyinput38), .B1(n6869), .B2(keyinput16), 
        .ZN(n6868) );
  OAI221_X1 U7802 ( .B1(n6870), .B2(keyinput38), .C1(n6869), .C2(keyinput16), 
        .A(n6868), .ZN(n6871) );
  AOI211_X1 U7803 ( .C1(keyinput20), .C2(n6873), .A(n6872), .B(n6871), .ZN(
        n6899) );
  INV_X1 U7804 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6876) );
  INV_X1 U7805 ( .A(DATAI_21_), .ZN(n6875) );
  OAI22_X1 U7806 ( .A1(n6876), .A2(keyinput95), .B1(n6875), .B2(keyinput108), 
        .ZN(n6874) );
  AOI221_X1 U7807 ( .B1(n6876), .B2(keyinput95), .C1(keyinput108), .C2(n6875), 
        .A(n6874), .ZN(n6898) );
  INV_X1 U7808 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6879) );
  INV_X1 U7809 ( .A(keyinput83), .ZN(n6878) );
  OAI22_X1 U7810 ( .A1(n6879), .A2(keyinput68), .B1(n6878), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6877) );
  AOI221_X1 U7811 ( .B1(n6879), .B2(keyinput68), .C1(DATAO_REG_14__SCAN_IN), 
        .C2(n6878), .A(n6877), .ZN(n6897) );
  INV_X1 U7812 ( .A(keyinput63), .ZN(n6881) );
  AOI22_X1 U7813 ( .A1(n6882), .A2(keyinput125), .B1(BYTEENABLE_REG_1__SCAN_IN), .B2(n6881), .ZN(n6880) );
  OAI221_X1 U7814 ( .B1(n6882), .B2(keyinput125), .C1(n6881), .C2(
        BYTEENABLE_REG_1__SCAN_IN), .A(n6880), .ZN(n6895) );
  INV_X1 U7815 ( .A(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n6884) );
  AOI22_X1 U7816 ( .A1(n6885), .A2(keyinput92), .B1(n6884), .B2(keyinput10), 
        .ZN(n6883) );
  OAI221_X1 U7817 ( .B1(n6885), .B2(keyinput92), .C1(n6884), .C2(keyinput10), 
        .A(n6883), .ZN(n6894) );
  INV_X1 U7818 ( .A(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n6888) );
  INV_X1 U7819 ( .A(keyinput56), .ZN(n6887) );
  AOI22_X1 U7820 ( .A1(n6888), .A2(keyinput112), .B1(DATAO_REG_13__SCAN_IN), 
        .B2(n6887), .ZN(n6886) );
  OAI221_X1 U7821 ( .B1(n6888), .B2(keyinput112), .C1(n6887), .C2(
        DATAO_REG_13__SCAN_IN), .A(n6886), .ZN(n6893) );
  AOI22_X1 U7822 ( .A1(n6891), .A2(keyinput5), .B1(keyinput26), .B2(n6890), 
        .ZN(n6889) );
  OAI221_X1 U7823 ( .B1(n6891), .B2(keyinput5), .C1(n6890), .C2(keyinput26), 
        .A(n6889), .ZN(n6892) );
  NOR4_X1 U7824 ( .A1(n6895), .A2(n6894), .A3(n6893), .A4(n6892), .ZN(n6896)
         );
  NAND4_X1 U7825 ( .A1(n6899), .A2(n6898), .A3(n6897), .A4(n6896), .ZN(n6995)
         );
  INV_X1 U7826 ( .A(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n6901) );
  OAI22_X1 U7827 ( .A1(n6901), .A2(keyinput109), .B1(n4096), .B2(keyinput11), 
        .ZN(n6900) );
  AOI221_X1 U7828 ( .B1(n6901), .B2(keyinput109), .C1(keyinput11), .C2(n4096), 
        .A(n6900), .ZN(n6912) );
  OAI22_X1 U7829 ( .A1(n6903), .A2(keyinput52), .B1(n4853), .B2(keyinput29), 
        .ZN(n6902) );
  AOI221_X1 U7830 ( .B1(n6903), .B2(keyinput52), .C1(keyinput29), .C2(n4853), 
        .A(n6902), .ZN(n6911) );
  INV_X1 U7831 ( .A(keyinput124), .ZN(n6905) );
  OAI22_X1 U7832 ( .A1(n5816), .A2(keyinput73), .B1(n6905), .B2(
        DATAWIDTH_REG_20__SCAN_IN), .ZN(n6904) );
  AOI221_X1 U7833 ( .B1(n5816), .B2(keyinput73), .C1(DATAWIDTH_REG_20__SCAN_IN), .C2(n6905), .A(n6904), .ZN(n6910) );
  INV_X1 U7834 ( .A(keyinput94), .ZN(n6906) );
  XNOR2_X1 U7835 ( .A(n6906), .B(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6908) );
  XOR2_X1 U7836 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .B(keyinput14), .Z(n6907)
         );
  NOR2_X1 U7837 ( .A1(n6908), .A2(n6907), .ZN(n6909) );
  NAND4_X1 U7838 ( .A1(n6912), .A2(n6911), .A3(n6910), .A4(n6909), .ZN(n6994)
         );
  INV_X1 U7839 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n6915) );
  INV_X1 U7840 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n6918) );
  OAI22_X1 U7841 ( .A1(n6918), .A2(keyinput122), .B1(n6917), .B2(
        ADDRESS_REG_15__SCAN_IN), .ZN(n6916) );
  AOI221_X1 U7842 ( .B1(n6918), .B2(keyinput122), .C1(ADDRESS_REG_15__SCAN_IN), 
        .C2(n6917), .A(n6916), .ZN(n6927) );
  INV_X1 U7843 ( .A(keyinput22), .ZN(n6920) );
  OAI22_X1 U7844 ( .A1(n6921), .A2(keyinput115), .B1(n6920), .B2(
        ADDRESS_REG_17__SCAN_IN), .ZN(n6919) );
  AOI221_X1 U7845 ( .B1(n6921), .B2(keyinput115), .C1(ADDRESS_REG_17__SCAN_IN), 
        .C2(n6920), .A(n6919), .ZN(n6926) );
  INV_X1 U7846 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6924) );
  OAI22_X1 U7847 ( .A1(n6924), .A2(keyinput76), .B1(n6923), .B2(keyinput82), 
        .ZN(n6922) );
  AOI221_X1 U7848 ( .B1(n6924), .B2(keyinput76), .C1(keyinput82), .C2(n6923), 
        .A(n6922), .ZN(n6925) );
  NAND4_X1 U7849 ( .A1(n6928), .A2(n6927), .A3(n6926), .A4(n6925), .ZN(n6993)
         );
  AOI22_X1 U7850 ( .A1(n6930), .A2(keyinput57), .B1(keyinput67), .B2(n5215), 
        .ZN(n6929) );
  OAI221_X1 U7851 ( .B1(n6930), .B2(keyinput57), .C1(n5215), .C2(keyinput67), 
        .A(n6929), .ZN(n6943) );
  INV_X1 U7852 ( .A(keyinput69), .ZN(n6932) );
  AOI22_X1 U7853 ( .A1(n6933), .A2(keyinput103), .B1(ADDRESS_REG_25__SCAN_IN), 
        .B2(n6932), .ZN(n6931) );
  OAI221_X1 U7854 ( .B1(n6933), .B2(keyinput103), .C1(n6932), .C2(
        ADDRESS_REG_25__SCAN_IN), .A(n6931), .ZN(n6942) );
  INV_X1 U7855 ( .A(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n6936) );
  AOI22_X1 U7856 ( .A1(n6936), .A2(keyinput49), .B1(keyinput37), .B2(n6935), 
        .ZN(n6934) );
  OAI221_X1 U7857 ( .B1(n6936), .B2(keyinput49), .C1(n6935), .C2(keyinput37), 
        .A(n6934), .ZN(n6941) );
  INV_X1 U7858 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n6938) );
  AOI22_X1 U7859 ( .A1(n6939), .A2(keyinput100), .B1(keyinput65), .B2(n6938), 
        .ZN(n6937) );
  OAI221_X1 U7860 ( .B1(n6939), .B2(keyinput100), .C1(n6938), .C2(keyinput65), 
        .A(n6937), .ZN(n6940) );
  NOR4_X1 U7861 ( .A1(n6943), .A2(n6942), .A3(n6941), .A4(n6940), .ZN(n6991)
         );
  INV_X1 U7862 ( .A(UWORD_REG_8__SCAN_IN), .ZN(n6945) );
  AOI22_X1 U7863 ( .A1(n6946), .A2(keyinput6), .B1(keyinput47), .B2(n6945), 
        .ZN(n6944) );
  OAI221_X1 U7864 ( .B1(n6946), .B2(keyinput6), .C1(n6945), .C2(keyinput47), 
        .A(n6944), .ZN(n6957) );
  AOI22_X1 U7865 ( .A1(n6949), .A2(keyinput30), .B1(n6948), .B2(keyinput113), 
        .ZN(n6947) );
  OAI221_X1 U7866 ( .B1(n6949), .B2(keyinput30), .C1(n6948), .C2(keyinput113), 
        .A(n6947), .ZN(n6956) );
  AOI22_X1 U7867 ( .A1(n6951), .A2(keyinput33), .B1(n5806), .B2(keyinput54), 
        .ZN(n6950) );
  OAI221_X1 U7868 ( .B1(n6951), .B2(keyinput33), .C1(n5806), .C2(keyinput54), 
        .A(n6950), .ZN(n6955) );
  INV_X1 U7869 ( .A(DATAI_20_), .ZN(n6953) );
  AOI22_X1 U7870 ( .A1(n6953), .A2(keyinput53), .B1(n5849), .B2(keyinput127), 
        .ZN(n6952) );
  OAI221_X1 U7871 ( .B1(n6953), .B2(keyinput53), .C1(n5849), .C2(keyinput127), 
        .A(n6952), .ZN(n6954) );
  NOR4_X1 U7872 ( .A1(n6957), .A2(n6956), .A3(n6955), .A4(n6954), .ZN(n6990)
         );
  INV_X1 U7873 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6960) );
  AOI22_X1 U7874 ( .A1(n6960), .A2(keyinput31), .B1(keyinput102), .B2(n6959), 
        .ZN(n6958) );
  OAI221_X1 U7875 ( .B1(n6960), .B2(keyinput31), .C1(n6959), .C2(keyinput102), 
        .A(n6958), .ZN(n6972) );
  INV_X1 U7876 ( .A(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n6963) );
  AOI22_X1 U7877 ( .A1(n6963), .A2(keyinput8), .B1(keyinput114), .B2(n6962), 
        .ZN(n6961) );
  OAI221_X1 U7878 ( .B1(n6963), .B2(keyinput8), .C1(n6962), .C2(keyinput114), 
        .A(n6961), .ZN(n6971) );
  INV_X1 U7879 ( .A(keyinput15), .ZN(n6965) );
  AOI22_X1 U7880 ( .A1(n5280), .A2(keyinput60), .B1(DATAWIDTH_REG_4__SCAN_IN), 
        .B2(n6965), .ZN(n6964) );
  OAI221_X1 U7881 ( .B1(n5280), .B2(keyinput60), .C1(n6965), .C2(
        DATAWIDTH_REG_4__SCAN_IN), .A(n6964), .ZN(n6970) );
  INV_X1 U7882 ( .A(keyinput81), .ZN(n6966) );
  XOR2_X1 U7883 ( .A(DATAO_REG_31__SCAN_IN), .B(n6966), .Z(n6968) );
  XNOR2_X1 U7884 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .B(keyinput87), .ZN(n6967)
         );
  NAND2_X1 U7885 ( .A1(n6968), .A2(n6967), .ZN(n6969) );
  NOR4_X1 U7886 ( .A1(n6972), .A2(n6971), .A3(n6970), .A4(n6969), .ZN(n6989)
         );
  INV_X1 U7887 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n6975) );
  INV_X1 U7888 ( .A(keyinput120), .ZN(n6974) );
  AOI22_X1 U7889 ( .A1(n6975), .A2(keyinput75), .B1(BYTEENABLE_REG_0__SCAN_IN), 
        .B2(n6974), .ZN(n6973) );
  OAI221_X1 U7890 ( .B1(n6975), .B2(keyinput75), .C1(n6974), .C2(
        BYTEENABLE_REG_0__SCAN_IN), .A(n6973), .ZN(n6987) );
  INV_X1 U7891 ( .A(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n6980) );
  AOI22_X1 U7892 ( .A1(n6980), .A2(keyinput106), .B1(keyinput17), .B2(n6979), 
        .ZN(n6978) );
  OAI221_X1 U7893 ( .B1(n6980), .B2(keyinput106), .C1(n6979), .C2(keyinput17), 
        .A(n6978), .ZN(n6985) );
  INV_X1 U7894 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n6983) );
  AOI22_X1 U7895 ( .A1(n6983), .A2(keyinput50), .B1(n6982), .B2(keyinput36), 
        .ZN(n6981) );
  OAI221_X1 U7896 ( .B1(n6983), .B2(keyinput50), .C1(n6982), .C2(keyinput36), 
        .A(n6981), .ZN(n6984) );
  NOR4_X1 U7897 ( .A1(n6987), .A2(n6986), .A3(n6985), .A4(n6984), .ZN(n6988)
         );
  NAND4_X1 U7898 ( .A1(n6991), .A2(n6990), .A3(n6989), .A4(n6988), .ZN(n6992)
         );
  NOR4_X1 U7899 ( .A1(n6995), .A2(n6994), .A3(n6993), .A4(n6992), .ZN(n6996)
         );
  NAND4_X1 U7900 ( .A1(n6999), .A2(n6998), .A3(n6997), .A4(n6996), .ZN(n7000)
         );
  AOI211_X1 U7901 ( .C1(DATAO_REG_21__SCAN_IN), .C2(n7002), .A(n7001), .B(
        n7000), .ZN(n7006) );
  AOI222_X1 U7902 ( .A1(n6682), .A2(ADDRESS_REG_0__SCAN_IN), .B1(
        REIP_REG_2__SCAN_IN), .B2(n7004), .C1(REIP_REG_1__SCAN_IN), .C2(n7003), 
        .ZN(n7005) );
  XNOR2_X1 U7903 ( .A(n7006), .B(n7005), .ZN(U3184) );
  AND4_X1 U4045 ( .A1(n3176), .A2(n3175), .A3(n3174), .A4(n3173), .ZN(n3181)
         );
  AOI211_X2 U3568 ( .C1(n6477), .C2(n5786), .A(n5785), .B(n6476), .ZN(n5829)
         );
  CLKBUF_X1 U3594 ( .A(n3299), .Z(n4087) );
  CLKBUF_X1 U3599 ( .A(n3355), .Z(n3397) );
  CLKBUF_X1 U3747 ( .A(n3383), .Z(n3384) );
  CLKBUF_X1 U3756 ( .A(n3286), .Z(n4381) );
  CLKBUF_X1 U3823 ( .A(n3336), .Z(n4478) );
  CLKBUF_X1 U3896 ( .A(n5498), .Z(n5990) );
  CLKBUF_X1 U3940 ( .A(n4200), .Z(n5323) );
  CLKBUF_X1 U4166 ( .A(n5360), .Z(n5380) );
  CLKBUF_X1 U4248 ( .A(n3663), .Z(n4717) );
  CLKBUF_X1 U6671 ( .A(n5082), .Z(n6674) );
endmodule

