

module b17_C_AntiSAT_k_128_10 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9674,
         n9675, n9676, n9677, n9678, n9679, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727,
         n20728, n20729, n20730, n20731, n20732, n20733, n20734, n20735,
         n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743,
         n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751,
         n20752, n20753, n20754, n20755, n20756, n20757, n20758, n20759,
         n20760, n20761, n20762, n20763, n20764, n20765, n20766, n20767,
         n20768, n20769, n20770, n20771, n20772, n20773, n20774, n20775,
         n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
         n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791,
         n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799,
         n20800, n20801, n20802, n20803, n20804, n20805, n20806, n20807,
         n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815,
         n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823,
         n20824, n20825, n20826, n20827, n20828, n20829, n20830, n20831,
         n20832, n20833, n20834, n20835, n20836, n20837, n20838, n20839,
         n20840, n20841, n20842, n20843, n20844, n20845, n20846, n20847,
         n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
         n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863,
         n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871,
         n20872, n20873, n20874, n20875, n20876, n20877, n20878, n20879,
         n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887,
         n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895,
         n20896, n20897, n20898, n20899, n20900, n20901, n20902, n20903,
         n20904, n20905, n20906, n20907, n20908, n20909, n20910, n20911,
         n20912, n20913, n20914, n20915, n20916, n20917, n20918, n20919,
         n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
         n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935,
         n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943,
         n20944, n20945, n20946, n20947, n20948, n20949, n20950, n20951,
         n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959,
         n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967,
         n20968, n20969, n20970, n20971, n20972, n20973, n20974, n20975,
         n20976, n20977, n20978, n20979, n20980, n20981, n20982, n20983,
         n20984, n20985, n20986, n20987, n20988, n20989, n20990, n20991,
         n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
         n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007,
         n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015,
         n21016, n21017, n21018, n21019, n21020, n21021, n21022, n21023,
         n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031,
         n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039,
         n21040, n21041, n21042, n21043, n21044, n21045, n21046, n21047,
         n21048, n21049, n21050, n21051, n21052, n21053, n21054, n21055,
         n21056, n21057, n21058, n21059, n21060, n21061, n21062, n21063,
         n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
         n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079,
         n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087,
         n21088, n21089, n21090, n21091, n21092, n21093, n21094, n21095,
         n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103,
         n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111,
         n21112;

  AND2_X1 U11076 ( .A1(n14234), .A2(n10086), .ZN(n14221) );
  NAND2_X1 U11077 ( .A1(n14093), .A2(n14094), .ZN(n14222) );
  NAND2_X1 U11078 ( .A1(n9724), .A2(n10169), .ZN(n10745) );
  INV_X1 U11079 ( .A(n17546), .ZN(n17770) );
  NOR2_X1 U11080 ( .A1(n19819), .A2(n19407), .ZN(n19457) );
  NAND2_X1 U11081 ( .A1(n13732), .A2(n10078), .ZN(n13960) );
  NOR2_X1 U11082 ( .A1(n16043), .A2(n13612), .ZN(n13737) );
  OR2_X1 U11083 ( .A1(n10809), .A2(n10808), .ZN(n10812) );
  XNOR2_X1 U11084 ( .A(n13357), .B(n13387), .ZN(n13382) );
  NAND2_X1 U11085 ( .A1(n9941), .A2(n13352), .ZN(n13357) );
  BUF_X1 U11086 ( .A(n17438), .Z(n9681) );
  OR2_X1 U11087 ( .A1(n10379), .A2(n10358), .ZN(n19466) );
  CLKBUF_X1 U11088 ( .A(n19065), .Z(n9647) );
  INV_X1 U11089 ( .A(n9682), .ZN(n9685) );
  AOI21_X1 U11090 ( .B1(n11919), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11920), .ZN(n11925) );
  CLKBUF_X1 U11091 ( .A(n11497), .Z(n17159) );
  NAND2_X1 U11092 ( .A1(n10392), .A2(n9846), .ZN(n11114) );
  INV_X1 U11093 ( .A(n9717), .ZN(n14682) );
  AND2_X1 U11094 ( .A1(n10386), .A2(n14749), .ZN(n14767) );
  NOR2_X1 U11095 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14749) );
  CLKBUF_X2 U11096 ( .A(n12115), .Z(n9679) );
  CLKBUF_X2 U11097 ( .A(n11530), .Z(n17176) );
  CLKBUF_X2 U11098 ( .A(n11497), .Z(n17138) );
  INV_X1 U11099 ( .A(n15530), .ZN(n17161) );
  CLKBUF_X1 U11100 ( .A(n11530), .Z(n17069) );
  OR2_X1 U11101 ( .A1(n13132), .A2(n14096), .ZN(n13245) );
  NAND2_X2 U11102 ( .A1(n11892), .A2(n20104), .ZN(n9972) );
  INV_X2 U11103 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18796) );
  NAND4_X2 U11104 ( .A1(n11875), .A2(n11874), .A3(n11873), .A4(n11872), .ZN(
        n20114) );
  NOR2_X1 U11105 ( .A1(n11771), .A2(n11770), .ZN(n11772) );
  NAND2_X2 U11106 ( .A1(n10210), .A2(n10209), .ZN(n10265) );
  AND2_X1 U11107 ( .A1(n11762), .A2(n14599), .ZN(n11928) );
  AND2_X1 U11108 ( .A1(n11761), .A2(n11756), .ZN(n11800) );
  AND2_X1 U11109 ( .A1(n11761), .A2(n11764), .ZN(n11929) );
  AND2_X1 U11110 ( .A1(n13149), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11927) );
  AND2_X2 U11111 ( .A1(n11762), .A2(n13161), .ZN(n12028) );
  AND2_X2 U11112 ( .A1(n11761), .A2(n13161), .ZN(n12560) );
  AND2_X1 U11113 ( .A1(n9964), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11756) );
  AND2_X2 U11114 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10399) );
  CLKBUF_X1 U11115 ( .A(n20179), .Z(n9632) );
  NOR2_X1 U11116 ( .A1(n20101), .A2(n20102), .ZN(n20179) );
  INV_X1 U11117 ( .A(n9633), .ZN(n20795) );
  NAND2_X1 U11118 ( .A1(DATAI_22_), .A2(n9632), .ZN(n9634) );
  NAND2_X1 U11119 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n9636), .ZN(n9635) );
  NAND2_X1 U11120 ( .A1(n9634), .A2(n9635), .ZN(n9633) );
  CLKBUF_X1 U11121 ( .A(n20180), .Z(n9636) );
  NOR2_X1 U11122 ( .A1(n20101), .A2(n20100), .ZN(n20180) );
  INV_X4 U11123 ( .A(n18077), .ZN(n9654) );
  CLKBUF_X2 U11124 ( .A(n12560), .Z(n9666) );
  INV_X1 U11125 ( .A(n14738), .ZN(n14771) );
  AND2_X1 U11126 ( .A1(n10399), .A2(n10400), .ZN(n14782) );
  INV_X1 U11127 ( .A(n10158), .ZN(n14783) );
  INV_X2 U11128 ( .A(n9639), .ZN(n9644) );
  AND2_X1 U11129 ( .A1(n11763), .A2(n14599), .ZN(n12017) );
  AND2_X1 U11130 ( .A1(n11756), .A2(n11762), .ZN(n12115) );
  AND2_X2 U11131 ( .A1(n13462), .A2(n10387), .ZN(n10397) );
  NAND2_X1 U11132 ( .A1(n14757), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10472) );
  NAND2_X1 U11133 ( .A1(n10397), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10463) );
  NAND2_X1 U11134 ( .A1(n14748), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10467) );
  AND4_X1 U11135 ( .A1(n11783), .A2(n11782), .A3(n11781), .A4(n11780), .ZN(
        n11794) );
  NAND2_X1 U11136 ( .A1(n14505), .A2(n10097), .ZN(n10100) );
  AND2_X1 U11137 ( .A1(n15871), .A2(n15875), .ZN(n14053) );
  NAND2_X1 U11138 ( .A1(n13678), .A2(n13677), .ZN(n13680) );
  AND2_X1 U11139 ( .A1(n11761), .A2(n14599), .ZN(n12026) );
  OR2_X1 U11140 ( .A1(n11808), .A2(n11807), .ZN(n20119) );
  CLKBUF_X2 U11141 ( .A(n10328), .Z(n10873) );
  NAND2_X1 U11142 ( .A1(n18820), .A2(n18814), .ZN(n16905) );
  AND2_X1 U11143 ( .A1(n9818), .A2(n15836), .ZN(n14447) );
  INV_X1 U11144 ( .A(n20114), .ZN(n13219) );
  NAND2_X1 U11145 ( .A1(n12978), .A2(n10294), .ZN(n10269) );
  NAND2_X1 U11146 ( .A1(n9911), .A2(n10631), .ZN(n10632) );
  INV_X1 U11147 ( .A(n10984), .ZN(n10983) );
  INV_X1 U11148 ( .A(n13522), .ZN(n10022) );
  AND2_X1 U11149 ( .A1(n10376), .A2(n10373), .ZN(n13783) );
  NOR4_X2 U11150 ( .A1(n17369), .A2(n17371), .A3(n17340), .A4(n17225), .ZN(
        n17310) );
  INV_X1 U11151 ( .A(n18192), .ZN(n18840) );
  INV_X1 U11152 ( .A(n12649), .ZN(n9648) );
  INV_X1 U11153 ( .A(n19987), .ZN(n19932) );
  NAND2_X1 U11154 ( .A1(n14146), .A2(n13983), .ZN(n15853) );
  NAND2_X1 U11155 ( .A1(n13214), .A2(n13213), .ZN(n13260) );
  NOR2_X1 U11156 ( .A1(n10876), .A2(n11354), .ZN(n11353) );
  NOR2_X1 U11157 ( .A1(n16296), .A2(n15411), .ZN(n15399) );
  NOR2_X1 U11158 ( .A1(n11411), .A2(n11410), .ZN(n11435) );
  OR2_X1 U11159 ( .A1(n15098), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15263) );
  OAI21_X1 U11160 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18837), .A(n16524), 
        .ZN(n17858) );
  INV_X1 U11161 ( .A(n17858), .ZN(n17845) );
  NOR2_X1 U11162 ( .A1(n18840), .A2(n16524), .ZN(n17850) );
  INV_X1 U11163 ( .A(n19916), .ZN(n19923) );
  INV_X1 U11164 ( .A(n20074), .ZN(n19877) );
  INV_X2 U11165 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14130) );
  AND2_X1 U11166 ( .A1(n9805), .A2(n9804), .ZN(n9637) );
  OR3_X1 U11167 ( .A1(n15037), .A2(n10028), .A3(n10031), .ZN(n9638) );
  NAND2_X1 U11168 ( .A1(n13161), .A2(n11763), .ZN(n9639) );
  INV_X1 U11169 ( .A(n10265), .ZN(n11029) );
  NAND2_X2 U11171 ( .A1(n17835), .A2(n11539), .ZN(n11542) );
  NAND2_X2 U11172 ( .A1(n9949), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10291) );
  INV_X2 U11173 ( .A(n10391), .ZN(n10184) );
  NAND2_X1 U11174 ( .A1(n13231), .A2(n13230), .ZN(n13351) );
  NOR2_X2 U11175 ( .A1(n14255), .A2(n9774), .ZN(n14334) );
  OAI222_X1 U11176 ( .A1(n14350), .A2(n14431), .B1(n14100), .B2(n20016), .C1(
        n14567), .C2(n20005), .ZN(P1_U2844) );
  NAND2_X1 U11177 ( .A1(n10096), .A2(n12069), .ZN(n12076) );
  OAI211_X1 U11178 ( .C1(n9824), .C2(n9821), .A(n9741), .B(n9819), .ZN(n10096)
         );
  AND2_X4 U11179 ( .A1(n14234), .A2(n12513), .ZN(n14093) );
  AND2_X2 U11180 ( .A1(n13462), .A2(n10387), .ZN(n9640) );
  NOR2_X2 U11181 ( .A1(n17388), .A2(n17254), .ZN(n17249) );
  INV_X8 U11182 ( .A(n10156), .ZN(n17154) );
  AOI22_X1 U11183 ( .A1(n18838), .A2(n15713), .B1(n15712), .B2(n15711), .ZN(
        n17369) );
  INV_X2 U11184 ( .A(n9639), .ZN(n9642) );
  INV_X2 U11185 ( .A(n9639), .ZN(n9643) );
  OR2_X1 U11186 ( .A1(n20424), .A2(n13701), .ZN(n13241) );
  NAND2_X2 U11187 ( .A1(n10149), .A2(n10151), .ZN(n10829) );
  OR2_X2 U11188 ( .A1(n17541), .A2(n17645), .ZN(n9733) );
  NOR2_X2 U11189 ( .A1(n11757), .A2(n12579), .ZN(n13149) );
  INV_X1 U11190 ( .A(n10364), .ZN(n13068) );
  OR2_X4 U11191 ( .A1(n11854), .A2(n11853), .ZN(n20104) );
  INV_X4 U11192 ( .A(n10157), .ZN(n17171) );
  XNOR2_X2 U11193 ( .A(n10722), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15129) );
  AND2_X4 U11194 ( .A1(n10386), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9645) );
  NOR2_X4 U11195 ( .A1(n19231), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11075) );
  NOR2_X2 U11196 ( .A1(n18840), .A2(n17990), .ZN(n17923) );
  INV_X1 U11197 ( .A(n11800), .ZN(n9682) );
  AND2_X2 U11198 ( .A1(n13481), .A2(n13462), .ZN(n9646) );
  NAND2_X1 U11199 ( .A1(n14447), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14572) );
  NAND2_X1 U11200 ( .A1(n15211), .A2(n9873), .ZN(n15157) );
  OR2_X1 U11201 ( .A1(n14470), .A2(n13929), .ZN(n14051) );
  OR2_X1 U11203 ( .A1(n10588), .A2(n10587), .ZN(n10589) );
  AND2_X1 U11204 ( .A1(n13552), .A2(n10043), .ZN(n14024) );
  NAND2_X1 U11205 ( .A1(n10718), .A2(n10735), .ZN(n10716) );
  NAND2_X1 U11206 ( .A1(n13068), .A2(n10368), .ZN(n10571) );
  NAND2_X1 U11207 ( .A1(n13068), .A2(n10366), .ZN(n19677) );
  AND2_X1 U11208 ( .A1(n10376), .A2(n10374), .ZN(n19295) );
  NAND2_X1 U11209 ( .A1(n13068), .A2(n10365), .ZN(n13423) );
  NAND2_X1 U11210 ( .A1(n13068), .A2(n10367), .ZN(n10417) );
  NAND2_X1 U11211 ( .A1(n12976), .A2(n12975), .ZN(n15453) );
  BUF_X1 U11212 ( .A(n11360), .Z(n9690) );
  CLKBUF_X2 U11213 ( .A(n10353), .Z(n10360) );
  AND2_X1 U11214 ( .A1(n10979), .A2(n10252), .ZN(n11299) );
  NAND2_X1 U11215 ( .A1(n17311), .A2(n18188), .ZN(n11663) );
  INV_X2 U11216 ( .A(n9649), .ZN(n13441) );
  INV_X4 U11217 ( .A(n10640), .ZN(n10962) );
  NAND2_X1 U11218 ( .A1(n9729), .A2(n9990), .ZN(n17364) );
  INV_X1 U11219 ( .A(n10294), .ZN(n12971) );
  NAND2_X1 U11220 ( .A1(n10197), .A2(n10196), .ZN(n13434) );
  CLKBUF_X2 U11221 ( .A(n12026), .Z(n12027) );
  CLKBUF_X2 U11222 ( .A(n11928), .Z(n12471) );
  BUF_X2 U11223 ( .A(n12011), .Z(n12561) );
  BUF_X2 U11224 ( .A(n11485), .Z(n17149) );
  CLKBUF_X2 U11225 ( .A(n11930), .Z(n12360) );
  INV_X1 U11226 ( .A(n11443), .ZN(n15530) );
  CLKBUF_X2 U11227 ( .A(n11927), .Z(n12470) );
  BUF_X2 U11228 ( .A(n11929), .Z(n12033) );
  CLKBUF_X2 U11229 ( .A(n12017), .Z(n12555) );
  NOR2_X1 U11230 ( .A1(n11442), .A2(n11447), .ZN(n11443) );
  NOR2_X2 U11231 ( .A1(n16905), .A2(n11445), .ZN(n11446) );
  CLKBUF_X2 U11232 ( .A(n10257), .Z(n14826) );
  AND2_X1 U11233 ( .A1(n14130), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11764) );
  NOR2_X4 U11234 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13454) );
  AOI21_X1 U11236 ( .B1(n15276), .B2(n16314), .A(n15275), .ZN(n15277) );
  AOI21_X1 U11237 ( .B1(n14995), .B2(n16312), .A(n10036), .ZN(n11307) );
  NAND2_X1 U11238 ( .A1(n9871), .A2(n15104), .ZN(n15290) );
  AOI21_X1 U11239 ( .B1(n16197), .B2(n16269), .A(n9959), .ZN(n16200) );
  OAI22_X1 U11240 ( .A1(n14410), .A2(n9948), .B1(n14156), .B2(n9767), .ZN(
        n9947) );
  NAND2_X1 U11241 ( .A1(n9831), .A2(n9763), .ZN(n9830) );
  OR2_X1 U11242 ( .A1(n11394), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11395) );
  OR2_X1 U11243 ( .A1(n10747), .A2(n10746), .ZN(n10163) );
  OR2_X1 U11244 ( .A1(n11436), .A2(n19221), .ZN(n11437) );
  AND2_X1 U11245 ( .A1(n9963), .A2(n9962), .ZN(n16197) );
  OR2_X1 U11246 ( .A1(n11436), .A2(n16326), .ZN(n11427) );
  OR2_X1 U11247 ( .A1(n16202), .A2(n15389), .ZN(n9963) );
  NAND2_X1 U11248 ( .A1(n15410), .A2(n15385), .ZN(n16202) );
  NOR2_X1 U11249 ( .A1(n15217), .A2(n15151), .ZN(n15201) );
  CLKBUF_X1 U11250 ( .A(n15121), .Z(n15135) );
  AND2_X1 U11251 ( .A1(n15838), .A2(n15837), .ZN(n15944) );
  NAND2_X1 U11252 ( .A1(n10123), .A2(n15138), .ZN(n15130) );
  INV_X1 U11253 ( .A(n16231), .ZN(n15410) );
  OR2_X1 U11254 ( .A1(n15228), .A2(n15219), .ZN(n16231) );
  AOI21_X1 U11255 ( .B1(n14209), .B2(n15909), .A(n14165), .ZN(n14166) );
  NAND2_X1 U11256 ( .A1(n14152), .A2(n9834), .ZN(n15836) );
  XNOR2_X1 U11257 ( .A(n14162), .B(n14161), .ZN(n14209) );
  AOI21_X1 U11258 ( .B1(n10811), .B2(n9956), .A(n9955), .ZN(n9953) );
  OR2_X1 U11259 ( .A1(n14961), .A2(n9928), .ZN(n14879) );
  OR3_X1 U11260 ( .A1(n15853), .A2(n9834), .A3(n14518), .ZN(n15666) );
  OAI21_X1 U11261 ( .B1(n14963), .B2(n10047), .A(n10046), .ZN(n14948) );
  NAND2_X1 U11262 ( .A1(n9862), .A2(n10807), .ZN(n10811) );
  NAND2_X1 U11263 ( .A1(n14147), .A2(n9834), .ZN(n14460) );
  AND2_X1 U11264 ( .A1(n10806), .A2(n9863), .ZN(n9862) );
  XNOR2_X1 U11265 ( .A(n14857), .B(n10167), .ZN(n14963) );
  NAND2_X1 U11266 ( .A1(n14966), .A2(n14841), .ZN(n14857) );
  OR2_X1 U11267 ( .A1(n14840), .A2(n14839), .ZN(n14841) );
  XNOR2_X1 U11268 ( .A(n10813), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16246) );
  AND2_X1 U11269 ( .A1(n10099), .A2(n9799), .ZN(n10098) );
  NOR3_X1 U11270 ( .A1(n11401), .A2(n10109), .A3(n10108), .ZN(n11416) );
  NAND2_X1 U11271 ( .A1(n9924), .A2(n9923), .ZN(n14838) );
  AOI21_X1 U11272 ( .B1(n10091), .B2(n10090), .A(n9737), .ZN(n9826) );
  NAND3_X1 U11273 ( .A1(n9814), .A2(n9813), .A3(n9734), .ZN(n15908) );
  NAND2_X1 U11274 ( .A1(n10592), .A2(n19030), .ZN(n10593) );
  AOI21_X1 U11275 ( .B1(n9696), .B2(n10092), .A(n9739), .ZN(n10091) );
  AOI211_X1 U11276 ( .C1(n19110), .C2(BUF1_REG_28__SCAN_IN), .A(n15011), .B(
        n15010), .ZN(n15012) );
  NOR2_X1 U11277 ( .A1(n15064), .A2(n14792), .ZN(n14794) );
  NOR2_X2 U11278 ( .A1(n15055), .A2(n15057), .ZN(n15056) );
  AND2_X1 U11279 ( .A1(n9742), .A2(n13699), .ZN(n9696) );
  AND2_X1 U11280 ( .A1(n14056), .A2(n15874), .ZN(n9969) );
  OAI21_X1 U11281 ( .B1(n15014), .B2(n15009), .A(n15008), .ZN(n16097) );
  AOI211_X1 U11282 ( .C1(n17706), .C2(n16872), .A(n16412), .B(n16373), .ZN(
        n16378) );
  AND2_X1 U11283 ( .A1(n13976), .A2(n13975), .ZN(n15871) );
  OR2_X1 U11284 ( .A1(n13512), .A2(n13611), .ZN(n9806) );
  NAND2_X1 U11285 ( .A1(n10630), .A2(n10629), .ZN(n10808) );
  INV_X1 U11286 ( .A(n10138), .ZN(n10137) );
  INV_X2 U11287 ( .A(n15855), .ZN(n15831) );
  NOR2_X1 U11288 ( .A1(n9722), .A2(n15015), .ZN(n15014) );
  INV_X1 U11289 ( .A(n13705), .ZN(n15855) );
  NAND2_X1 U11290 ( .A1(n14024), .A2(n16178), .ZN(n14046) );
  OR2_X1 U11291 ( .A1(n13705), .A2(n15993), .ZN(n13976) );
  NOR2_X1 U11292 ( .A1(n19626), .A2(n19597), .ZN(n19614) );
  OR2_X1 U11293 ( .A1(n10613), .A2(n10612), .ZN(n10630) );
  XNOR2_X1 U11294 ( .A(n13704), .B(n12136), .ZN(n13691) );
  NOR2_X1 U11295 ( .A1(n19497), .A2(n19407), .ZN(n19286) );
  AND2_X1 U11296 ( .A1(n13408), .A2(n13343), .ZN(n13446) );
  OAI21_X1 U11297 ( .B1(n19466), .B2(n11178), .A(n9906), .ZN(n10359) );
  XNOR2_X1 U11298 ( .A(n13351), .B(n13244), .ZN(n13350) );
  AND2_X1 U11299 ( .A1(n10372), .A2(n10371), .ZN(n9662) );
  AND2_X1 U11300 ( .A1(n9909), .A2(n9910), .ZN(n10420) );
  NOR2_X2 U11301 ( .A1(n17861), .A2(n17341), .ZN(n17768) );
  AND2_X1 U11302 ( .A1(n13529), .A2(n13057), .ZN(n13065) );
  OR2_X1 U11303 ( .A1(n13192), .A2(n13056), .ZN(n13529) );
  AND2_X1 U11304 ( .A1(n10164), .A2(n13190), .ZN(n10042) );
  OR2_X1 U11305 ( .A1(n9715), .A2(n14307), .ZN(n14309) );
  OR2_X1 U11306 ( .A1(n13072), .A2(n13071), .ZN(n13074) );
  NAND2_X1 U11307 ( .A1(n13016), .A2(n13015), .ZN(n13061) );
  XNOR2_X1 U11308 ( .A(n15453), .B(n13010), .ZN(n13011) );
  CLKBUF_X1 U11309 ( .A(n16018), .Z(n16062) );
  NAND2_X2 U11310 ( .A1(n20016), .A2(n20172), .ZN(n14350) );
  AND2_X1 U11311 ( .A1(n9647), .A2(n10360), .ZN(n10375) );
  NAND2_X1 U11312 ( .A1(n12054), .A2(n12053), .ZN(n13227) );
  INV_X2 U11313 ( .A(n13182), .ZN(n20066) );
  AND2_X1 U11314 ( .A1(n9647), .A2(n10361), .ZN(n10377) );
  NOR2_X2 U11315 ( .A1(n16191), .A2(n19442), .ZN(n13433) );
  CLKBUF_X1 U11316 ( .A(n12056), .Z(n20225) );
  NAND2_X1 U11317 ( .A1(n10735), .A2(n10663), .ZN(n10662) );
  AND2_X1 U11318 ( .A1(n9802), .A2(n11959), .ZN(n11943) );
  NAND2_X1 U11319 ( .A1(n14078), .A2(n18658), .ZN(n18661) );
  OAI21_X2 U11320 ( .B1(n19743), .B2(n12792), .A(n12901), .ZN(n12793) );
  NOR2_X1 U11321 ( .A1(n11090), .A2(n10019), .ZN(n10021) );
  INV_X2 U11322 ( .A(n19071), .ZN(n19028) );
  NAND3_X1 U11323 ( .A1(n10161), .A2(n10306), .A3(n10305), .ZN(n9858) );
  AND2_X1 U11324 ( .A1(n10550), .A2(n10551), .ZN(n10591) );
  NAND2_X1 U11325 ( .A1(n11338), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11337) );
  INV_X2 U11326 ( .A(n17221), .ZN(n17214) );
  INV_X1 U11327 ( .A(n10013), .ZN(n11089) );
  OAI21_X1 U11328 ( .B1(n11881), .B2(n12953), .A(n13245), .ZN(n11882) );
  NAND2_X1 U11329 ( .A1(n11353), .A2(n10006), .ZN(n11358) );
  NAND2_X1 U11330 ( .A1(n9723), .A2(n12973), .ZN(n11019) );
  NAND3_X1 U11331 ( .A1(n13131), .A2(n11855), .A3(n13219), .ZN(n13075) );
  NOR2_X1 U11332 ( .A1(n11912), .A2(n11911), .ZN(n13254) );
  NOR4_X1 U11333 ( .A1(n18188), .A2(n11668), .A3(n17229), .A4(n11659), .ZN(
        n17438) );
  AND2_X1 U11334 ( .A1(n11888), .A2(n11887), .ZN(n13133) );
  NAND2_X1 U11335 ( .A1(n18188), .A2(n18840), .ZN(n11661) );
  INV_X1 U11336 ( .A(n11658), .ZN(n11668) );
  AND2_X1 U11337 ( .A1(n12626), .A2(n13690), .ZN(n12632) );
  OR2_X1 U11338 ( .A1(n11884), .A2(n11886), .ZN(n14594) );
  AND2_X1 U11339 ( .A1(n11351), .A2(n10002), .ZN(n11340) );
  INV_X1 U11340 ( .A(n13123), .ZN(n13148) );
  NOR2_X2 U11341 ( .A1(n11973), .A2(n20804), .ZN(n12626) );
  AND2_X1 U11342 ( .A1(n11973), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12631) );
  AND2_X1 U11343 ( .A1(n19257), .A2(n10265), .ZN(n9841) );
  NOR2_X1 U11344 ( .A1(n20124), .A2(n20119), .ZN(n13123) );
  NOR2_X2 U11345 ( .A1(n11611), .A2(n11610), .ZN(n18204) );
  NOR2_X2 U11346 ( .A1(n11571), .A2(n11570), .ZN(n18212) );
  OR2_X2 U11347 ( .A1(n11830), .A2(n11829), .ZN(n20124) );
  BUF_X4 U11348 ( .A(n12971), .Z(n9649) );
  NAND3_X2 U11349 ( .A1(n9725), .A2(n11816), .A3(n9692), .ZN(n20136) );
  NAND2_X2 U11350 ( .A1(n10222), .A2(n10221), .ZN(n19257) );
  AND4_X1 U11351 ( .A1(n11751), .A2(n11750), .A3(n11749), .A4(n11748), .ZN(
        n11775) );
  AND4_X1 U11352 ( .A1(n11863), .A2(n11862), .A3(n11861), .A4(n11860), .ZN(
        n11874) );
  AND2_X1 U11353 ( .A1(n11844), .A2(n11843), .ZN(n11848) );
  INV_X2 U11354 ( .A(U214), .ZN(n16464) );
  AND4_X1 U11355 ( .A1(n11779), .A2(n11778), .A3(n11777), .A4(n11776), .ZN(
        n11795) );
  AND4_X1 U11356 ( .A1(n11859), .A2(n11858), .A3(n11857), .A4(n11856), .ZN(
        n11875) );
  BUF_X4 U11357 ( .A(n11488), .Z(n9667) );
  AND4_X1 U11358 ( .A1(n11871), .A2(n11870), .A3(n11869), .A4(n11868), .ZN(
        n11872) );
  CLKBUF_X1 U11359 ( .A(n11820), .Z(n12514) );
  INV_X1 U11360 ( .A(n9682), .ZN(n9686) );
  AND4_X1 U11361 ( .A1(n11787), .A2(n11786), .A3(n11785), .A4(n11784), .ZN(
        n11793) );
  AND4_X1 U11362 ( .A1(n11791), .A2(n11790), .A3(n11789), .A4(n11788), .ZN(
        n11792) );
  INV_X2 U11363 ( .A(n15996), .ZN(n13376) );
  BUF_X2 U11364 ( .A(n11524), .Z(n17152) );
  BUF_X2 U11365 ( .A(n11485), .Z(n15557) );
  AND2_X1 U11366 ( .A1(n10244), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10015) );
  NAND2_X2 U11367 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19866), .ZN(n19805) );
  INV_X1 U11368 ( .A(n11446), .ZN(n15541) );
  NAND2_X2 U11369 ( .A1(n19866), .A2(n19752), .ZN(n19809) );
  AND2_X1 U11370 ( .A1(n10248), .A2(n9846), .ZN(n10017) );
  INV_X2 U11371 ( .A(n16511), .ZN(U215) );
  NAND2_X2 U11372 ( .A1(n18778), .A2(n18718), .ZN(n18770) );
  INV_X2 U11373 ( .A(n18717), .ZN(n18781) );
  CLKBUF_X2 U11374 ( .A(n11820), .Z(n12554) );
  CLKBUF_X1 U11375 ( .A(n13481), .Z(n9658) );
  AND2_X2 U11376 ( .A1(n10398), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9714) );
  BUF_X4 U11377 ( .A(n11477), .Z(n9651) );
  OR2_X1 U11378 ( .A1(n16905), .A2(n11444), .ZN(n9713) );
  OR2_X1 U11379 ( .A1(n11439), .A2(n18665), .ZN(n10155) );
  BUF_X4 U11380 ( .A(n11523), .Z(n9652) );
  AND2_X2 U11381 ( .A1(n9846), .A2(n10398), .ZN(n14784) );
  BUF_X4 U11382 ( .A(n11486), .Z(n9653) );
  INV_X2 U11383 ( .A(n16514), .ZN(n16516) );
  CLKBUF_X1 U11384 ( .A(n11359), .Z(n19036) );
  AND2_X2 U11385 ( .A1(n13161), .A2(n11765), .ZN(n12034) );
  NAND2_X1 U11386 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18814), .ZN(
        n11441) );
  BUF_X4 U11387 ( .A(n11525), .Z(n9655) );
  NAND2_X1 U11388 ( .A1(n18807), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11439) );
  OR2_X1 U11389 ( .A1(n11444), .A2(n18665), .ZN(n10157) );
  NOR2_X1 U11390 ( .A1(n11341), .A2(n10343), .ZN(n11343) );
  INV_X1 U11391 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12579) );
  NAND2_X2 U11392 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18665) );
  INV_X2 U11393 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18807) );
  INV_X1 U11394 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13150) );
  AND2_X1 U11395 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14599) );
  INV_X1 U11396 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10343) );
  INV_X1 U11397 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9664) );
  NOR2_X1 U11398 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10403) );
  NAND2_X1 U11399 ( .A1(n11021), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10304) );
  NAND2_X1 U11400 ( .A1(n9805), .A2(n9804), .ZN(n9656) );
  INV_X1 U11401 ( .A(n11877), .ZN(n9657) );
  AND2_X2 U11402 ( .A1(n10172), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13481) );
  NAND2_X1 U11404 ( .A1(n10304), .A2(n10303), .ZN(n10328) );
  NAND3_X1 U11405 ( .A1(n12971), .A2(n10271), .A3(n10268), .ZN(n9659) );
  CLKBUF_X1 U11406 ( .A(n11039), .Z(n9660) );
  NAND3_X1 U11407 ( .A1(n12971), .A2(n10271), .A3(n10268), .ZN(n11043) );
  NAND2_X2 U11408 ( .A1(n13359), .A2(n13358), .ZN(n13670) );
  AOI21_X1 U11409 ( .B1(n10124), .B2(n10265), .A(n11034), .ZN(n11039) );
  INV_X1 U11410 ( .A(n10173), .ZN(n9661) );
  AND2_X1 U11411 ( .A1(n10289), .A2(n10288), .ZN(n10161) );
  INV_X2 U11412 ( .A(n10311), .ZN(n10330) );
  INV_X2 U11413 ( .A(n18059), .ZN(n18656) );
  OAI222_X1 U11414 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n18219), .B1(
        P3_EBX_REG_17__SCAN_IN), .B2(n17063), .C1(n17076), .C2(n17062), .ZN(
        n17064) );
  BUF_X1 U11415 ( .A(n10777), .Z(n9663) );
  NOR3_X2 U11416 ( .A1(n17449), .A2(n17302), .A3(n17275), .ZN(n17265) );
  NAND2_X2 U11417 ( .A1(n9851), .A2(n10407), .ZN(n10484) );
  NAND2_X2 U11418 ( .A1(n10291), .A2(n10272), .ZN(n10340) );
  BUF_X4 U11419 ( .A(n12560), .Z(n9665) );
  AND2_X1 U11421 ( .A1(n10387), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9668) );
  AND2_X1 U11422 ( .A1(n10387), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9669) );
  NOR2_X4 U11423 ( .A1(n11591), .A2(n11590), .ZN(n18192) );
  AOI21_X1 U11424 ( .B1(n10330), .B2(P2_EBX_REG_0__SCAN_IN), .A(n10287), .ZN(
        n10288) );
  NAND2_X1 U11425 ( .A1(n10304), .A2(n10303), .ZN(n9670) );
  INV_X1 U11426 ( .A(n10873), .ZN(n9671) );
  AND2_X1 U11427 ( .A1(n14749), .A2(n10387), .ZN(n14766) );
  INV_X1 U11428 ( .A(n10410), .ZN(n19267) );
  AND2_X1 U11429 ( .A1(n13161), .A2(n11765), .ZN(n9672) );
  NAND2_X1 U11430 ( .A1(n11946), .A2(n20634), .ZN(n13724) );
  NAND2_X2 U11431 ( .A1(n11945), .A2(n11944), .ZN(n20634) );
  AND2_X2 U11432 ( .A1(n13474), .A2(n10293), .ZN(n9723) );
  INV_X1 U11433 ( .A(n10347), .ZN(n10337) );
  AND2_X1 U11434 ( .A1(n10014), .A2(n10016), .ZN(n9674) );
  NAND2_X2 U11435 ( .A1(n10298), .A2(n12978), .ZN(n10979) );
  AND2_X1 U11436 ( .A1(n11765), .A2(n11756), .ZN(n9675) );
  AND2_X1 U11437 ( .A1(n11765), .A2(n11756), .ZN(n11930) );
  BUF_X1 U11438 ( .A(n13472), .Z(n9676) );
  BUF_X2 U11439 ( .A(n13472), .Z(n9677) );
  NAND2_X1 U11441 ( .A1(n9845), .A2(n9842), .ZN(n13472) );
  NOR2_X2 U11442 ( .A1(n14046), .A2(n10038), .ZN(n14982) );
  AND2_X2 U11443 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10387) );
  XNOR2_X2 U11444 ( .A(n13680), .B(n13679), .ZN(n15913) );
  AND2_X2 U11445 ( .A1(n11300), .A2(n11033), .ZN(n11021) );
  NOR2_X2 U11446 ( .A1(n10280), .A2(n10279), .ZN(n11300) );
  NOR2_X2 U11447 ( .A1(n13960), .A2(n9773), .ZN(n14267) );
  OAI21_X1 U11448 ( .B1(n11396), .B2(n10136), .A(n10137), .ZN(n10135) );
  OR2_X2 U11449 ( .A1(n11396), .A2(n10134), .ZN(n9724) );
  XNOR2_X2 U11450 ( .A(n10593), .B(n10796), .ZN(n13743) );
  AOI21_X1 U11451 ( .B1(n15148), .B2(n15395), .A(n15149), .ZN(n16206) );
  NAND2_X2 U11452 ( .A1(n10128), .A2(n9768), .ZN(n15420) );
  NAND2_X2 U11453 ( .A1(n20114), .A2(n20124), .ZN(n12649) );
  AND2_X1 U11454 ( .A1(n10364), .A2(n10380), .ZN(n10376) );
  AND2_X1 U11455 ( .A1(n10364), .A2(n14657), .ZN(n10378) );
  INV_X1 U11456 ( .A(n11800), .ZN(n9683) );
  INV_X1 U11457 ( .A(n9682), .ZN(n9684) );
  INV_X1 U11458 ( .A(n9683), .ZN(n9687) );
  INV_X1 U11459 ( .A(n9683), .ZN(n9688) );
  INV_X1 U11460 ( .A(n9683), .ZN(n9689) );
  INV_X4 U11461 ( .A(n11027), .ZN(n19231) );
  NAND2_X1 U11462 ( .A1(n9674), .A2(n9676), .ZN(n10984) );
  AND2_X4 U11463 ( .A1(n10014), .A2(n10016), .ZN(n11027) );
  XNOR2_X2 U11464 ( .A(n10809), .B(n10808), .ZN(n10798) );
  OAI21_X1 U11465 ( .B1(n14673), .B2(n13049), .A(n13001), .ZN(n9922) );
  AOI22_X2 U11466 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n11323), .B1(n11377), 
        .B2(n16342), .ZN(n11360) );
  OAI21_X2 U11467 ( .B1(n14093), .B2(n14094), .A(n14222), .ZN(n14431) );
  NAND4_X4 U11468 ( .A1(n11775), .A2(n11774), .A3(n11773), .A4(n11772), .ZN(
        n11878) );
  NAND2_X1 U11469 ( .A1(n9637), .A2(n11998), .ZN(n12107) );
  NAND2_X1 U11470 ( .A1(n10319), .A2(n10318), .ZN(n10323) );
  INV_X1 U11471 ( .A(n10317), .ZN(n10318) );
  AND2_X1 U11472 ( .A1(n10798), .A2(n13866), .ZN(n10802) );
  AND2_X1 U11473 ( .A1(n19257), .A2(n19825), .ZN(n11078) );
  AND3_X1 U11474 ( .A1(n16085), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n10962), .ZN(n11423) );
  OAI21_X1 U11475 ( .B1(n19466), .B2(n11227), .A(n9908), .ZN(n10601) );
  OAI21_X1 U11476 ( .B1(n19466), .B2(n11214), .A(n9907), .ZN(n10574) );
  NAND2_X1 U11477 ( .A1(n10420), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n9867) );
  NAND2_X1 U11478 ( .A1(n10298), .A2(n10299), .ZN(n10300) );
  INV_X1 U11479 ( .A(n10359), .ZN(n9850) );
  NOR2_X1 U11480 ( .A1(n18219), .A2(n18200), .ZN(n11658) );
  AND2_X1 U11481 ( .A1(n10084), .A2(n9788), .ZN(n9803) );
  AND2_X1 U11482 ( .A1(n12270), .A2(n12248), .ZN(n10074) );
  INV_X1 U11483 ( .A(n13733), .ZN(n12172) );
  NAND2_X1 U11484 ( .A1(n9637), .A2(n9709), .ZN(n12131) );
  NAND2_X1 U11485 ( .A1(n9656), .A2(n11999), .ZN(n12000) );
  NAND2_X1 U11486 ( .A1(n14453), .A2(n14460), .ZN(n14152) );
  AND2_X1 U11487 ( .A1(n13980), .A2(n10102), .ZN(n10099) );
  NOR2_X1 U11488 ( .A1(n13981), .A2(n10101), .ZN(n10097) );
  INV_X1 U11489 ( .A(n13928), .ZN(n10101) );
  NOR2_X1 U11490 ( .A1(n10025), .A2(n15589), .ZN(n10024) );
  INV_X1 U11491 ( .A(n15384), .ZN(n10025) );
  NOR2_X1 U11492 ( .A1(n14049), .A2(n10114), .ZN(n10113) );
  INV_X1 U11493 ( .A(n15193), .ZN(n10114) );
  OR2_X1 U11494 ( .A1(n16250), .A2(n16247), .ZN(n10643) );
  NAND3_X1 U11495 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19830), .A3(n19679), 
        .ZN(n13429) );
  NOR2_X1 U11496 ( .A1(n16905), .A2(n11447), .ZN(n11486) );
  NOR2_X1 U11497 ( .A1(n11441), .A2(n11445), .ZN(n11477) );
  NOR2_X1 U11498 ( .A1(n11664), .A2(n11657), .ZN(n15472) );
  NAND2_X1 U11499 ( .A1(n17767), .A2(n11643), .ZN(n11561) );
  INV_X1 U11500 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9932) );
  NOR2_X1 U11501 ( .A1(n16523), .A2(n11661), .ZN(n14079) );
  OAI21_X1 U11502 ( .B1(n18200), .B2(n11656), .A(n11677), .ZN(n11666) );
  AOI21_X1 U11503 ( .B1(n11695), .B2(n11699), .A(n11694), .ZN(n11703) );
  NAND3_X1 U11504 ( .A1(n11658), .A2(n11706), .A3(n18640), .ZN(n15474) );
  INV_X1 U11505 ( .A(n12652), .ZN(n14167) );
  AND2_X1 U11506 ( .A1(n13268), .A2(n12952), .ZN(n13032) );
  INV_X1 U11507 ( .A(n13698), .ZN(n10092) );
  NAND2_X1 U11508 ( .A1(n15900), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13699) );
  NAND2_X1 U11509 ( .A1(n9824), .A2(n9820), .ZN(n9819) );
  INV_X1 U11510 ( .A(n10926), .ZN(n10109) );
  OR2_X1 U11511 ( .A1(n11402), .A2(n14954), .ZN(n10108) );
  AND4_X1 U11512 ( .A1(n10495), .A2(n10494), .A3(n10493), .A4(n10492), .ZN(
        n10501) );
  AND2_X1 U11513 ( .A1(n19231), .A2(n9649), .ZN(n11064) );
  NOR2_X1 U11514 ( .A1(n10145), .A2(n14133), .ZN(n10144) );
  INV_X1 U11515 ( .A(n10146), .ZN(n10145) );
  INV_X1 U11516 ( .A(n15051), .ZN(n10032) );
  INV_X1 U11517 ( .A(n10811), .ZN(n9957) );
  NAND2_X1 U11518 ( .A1(n14657), .A2(n13012), .ZN(n13016) );
  NAND2_X1 U11519 ( .A1(n11009), .A2(n11008), .ZN(n13467) );
  NAND2_X1 U11520 ( .A1(n19822), .A2(n19073), .ZN(n19592) );
  OR2_X1 U11521 ( .A1(n16163), .A2(n19011), .ZN(n10001) );
  INV_X1 U11522 ( .A(n10054), .ZN(n10959) );
  INV_X1 U11523 ( .A(n11063), .ZN(n11305) );
  INV_X1 U11524 ( .A(n16330), .ZN(n16312) );
  NAND2_X1 U11525 ( .A1(n20419), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12585) );
  INV_X1 U11526 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9964) );
  NAND2_X1 U11527 ( .A1(n10579), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n9866) );
  OR2_X1 U11528 ( .A1(n12590), .A2(n12595), .ZN(n12592) );
  AND2_X1 U11529 ( .A1(n12592), .A2(n12581), .ZN(n12610) );
  AND2_X1 U11530 ( .A1(n12470), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n9837) );
  CLKBUF_X1 U11531 ( .A(n12028), .Z(n12495) );
  CLKBUF_X1 U11532 ( .A(n12034), .Z(n12256) );
  AND2_X1 U11533 ( .A1(n12123), .A2(n12122), .ZN(n12132) );
  NAND2_X1 U11534 ( .A1(n11842), .A2(n20119), .ZN(n11819) );
  NAND2_X1 U11535 ( .A1(n11916), .A2(n11898), .ZN(n9809) );
  OAI21_X1 U11536 ( .B1(n10509), .B2(n10508), .A(n10507), .ZN(n10546) );
  NOR2_X1 U11537 ( .A1(n10685), .A2(n10064), .ZN(n10063) );
  INV_X1 U11538 ( .A(n10661), .ZN(n10064) );
  INV_X1 U11539 ( .A(n14973), .ZN(n9925) );
  NAND2_X1 U11540 ( .A1(n10598), .A2(n10597), .ZN(n10809) );
  INV_X1 U11541 ( .A(n10793), .ZN(n10598) );
  AND2_X1 U11542 ( .A1(n19251), .A2(n12986), .ZN(n10268) );
  NOR2_X1 U11543 ( .A1(n19244), .A2(n13434), .ZN(n10223) );
  AOI21_X1 U11544 ( .B1(n10971), .B2(n9841), .A(n13434), .ZN(n10972) );
  NOR2_X1 U11545 ( .A1(n11439), .A2(n11441), .ZN(n11494) );
  NOR2_X1 U11546 ( .A1(n17350), .A2(n11521), .ZN(n11519) );
  NAND2_X1 U11547 ( .A1(n19976), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13718) );
  AND2_X1 U11548 ( .A1(n9765), .A2(n14305), .ZN(n10084) );
  INV_X1 U11549 ( .A(n9797), .ZN(n10075) );
  INV_X1 U11550 ( .A(n13960), .ZN(n12249) );
  INV_X1 U11551 ( .A(n13763), .ZN(n10083) );
  NOR2_X1 U11552 ( .A1(n13887), .A2(n13951), .ZN(n10082) );
  OR2_X1 U11553 ( .A1(n20136), .A2(n20383), .ZN(n12264) );
  NAND2_X1 U11554 ( .A1(n9985), .A2(n14099), .ZN(n9984) );
  INV_X1 U11555 ( .A(n14247), .ZN(n9985) );
  OR2_X1 U11556 ( .A1(n12719), .A2(n9976), .ZN(n9975) );
  INV_X1 U11557 ( .A(n14328), .ZN(n9976) );
  NAND2_X1 U11558 ( .A1(n14459), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14453) );
  NOR2_X1 U11559 ( .A1(n9978), .A2(n13890), .ZN(n9977) );
  INV_X1 U11560 ( .A(n9979), .ZN(n9978) );
  NAND2_X1 U11561 ( .A1(n9942), .A2(n9731), .ZN(n13229) );
  NAND2_X1 U11562 ( .A1(n13724), .A2(n9944), .ZN(n9942) );
  NAND2_X1 U11563 ( .A1(n9944), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n9943) );
  OR2_X1 U11564 ( .A1(n11842), .A2(n12649), .ZN(n11888) );
  CLKBUF_X1 U11565 ( .A(n13036), .Z(n13201) );
  NOR2_X1 U11566 ( .A1(n10067), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10066) );
  INV_X1 U11567 ( .A(n10068), .ZN(n10067) );
  NAND2_X1 U11568 ( .A1(n10662), .A2(n9702), .ZN(n10702) );
  AND2_X1 U11569 ( .A1(n10591), .A2(n9727), .ZN(n10647) );
  OR2_X1 U11570 ( .A1(n10391), .A2(n9846), .ZN(n14738) );
  INV_X1 U11571 ( .A(n14858), .ZN(n9929) );
  INV_X1 U11572 ( .A(n13280), .ZN(n14876) );
  NAND2_X1 U11573 ( .A1(n14982), .A2(n15065), .ZN(n14793) );
  NAND2_X1 U11574 ( .A1(n10041), .A2(n10168), .ZN(n10040) );
  INV_X1 U11575 ( .A(n16171), .ZN(n10041) );
  AND2_X1 U11576 ( .A1(n10045), .A2(n10044), .ZN(n10043) );
  INV_X1 U11577 ( .A(n13861), .ZN(n10044) );
  NAND2_X1 U11578 ( .A1(n13000), .A2(n11027), .ZN(n13280) );
  NOR2_X1 U11579 ( .A1(n15105), .A2(n10012), .ZN(n10011) );
  INV_X1 U11580 ( .A(n14633), .ZN(n10112) );
  NOR2_X1 U11581 ( .A1(n10930), .A2(n10008), .ZN(n10007) );
  INV_X1 U11582 ( .A(n15024), .ZN(n10030) );
  INV_X1 U11583 ( .A(n15015), .ZN(n10029) );
  AND2_X1 U11584 ( .A1(n10118), .A2(n9917), .ZN(n9916) );
  NAND2_X1 U11585 ( .A1(n9726), .A2(n10715), .ZN(n9917) );
  NOR2_X1 U11586 ( .A1(n10122), .A2(n10119), .ZN(n10118) );
  INV_X1 U11587 ( .A(n15137), .ZN(n10119) );
  INV_X1 U11588 ( .A(n10120), .ZN(n9913) );
  AOI21_X1 U11589 ( .B1(n15129), .B2(n10121), .A(n9738), .ZN(n10120) );
  INV_X1 U11590 ( .A(n15138), .ZN(n10121) );
  AND2_X1 U11591 ( .A1(n14631), .A2(n15075), .ZN(n10035) );
  NOR2_X1 U11592 ( .A1(n13556), .A2(n10117), .ZN(n10116) );
  INV_X1 U11593 ( .A(n13445), .ZN(n10117) );
  NAND2_X1 U11594 ( .A1(n15211), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15228) );
  NOR2_X1 U11595 ( .A1(n10105), .A2(n13310), .ZN(n10104) );
  NAND3_X1 U11596 ( .A1(n9857), .A2(n9958), .A3(n13746), .ZN(n10799) );
  OR2_X1 U11597 ( .A1(n10440), .A2(n10439), .ZN(n10782) );
  NAND2_X1 U11598 ( .A1(n11071), .A2(n19231), .ZN(n11242) );
  AND2_X1 U11599 ( .A1(n13441), .A2(n19825), .ZN(n11071) );
  INV_X1 U11600 ( .A(n11242), .ZN(n11265) );
  AND2_X1 U11601 ( .A1(n14876), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n13010) );
  AND2_X1 U11602 ( .A1(n10356), .A2(n14673), .ZN(n9909) );
  AOI22_X1 U11603 ( .A1(n9645), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14826), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10186) );
  NAND2_X1 U11604 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11444) );
  NAND2_X1 U11605 ( .A1(n9904), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9903) );
  INV_X1 U11606 ( .A(n17536), .ZN(n9904) );
  AND2_X1 U11607 ( .A1(n17780), .A2(n11555), .ZN(n11556) );
  NAND2_X1 U11608 ( .A1(n11519), .A2(n17344), .ZN(n11552) );
  NOR2_X1 U11609 ( .A1(n17776), .A2(n18106), .ZN(n11734) );
  NOR2_X1 U11610 ( .A1(n18208), .A2(n18212), .ZN(n11651) );
  XNOR2_X1 U11611 ( .A(n17364), .B(n11726), .ZN(n11538) );
  INV_X1 U11612 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19899) );
  OR3_X1 U11613 ( .A1(n9981), .A2(n12703), .A3(n13984), .ZN(n9980) );
  INV_X1 U11614 ( .A(n13180), .ZN(n20054) );
  INV_X1 U11615 ( .A(n12078), .ZN(n14159) );
  AND2_X1 U11616 ( .A1(n20383), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14158) );
  AND2_X1 U11617 ( .A1(n14411), .A2(n13616), .ZN(n12575) );
  OR2_X1 U11618 ( .A1(n12533), .A2(n14226), .ZN(n13624) );
  AND2_X1 U11619 ( .A1(n10087), .A2(n12513), .ZN(n10086) );
  NOR2_X1 U11620 ( .A1(n10088), .A2(n14223), .ZN(n10087) );
  INV_X1 U11621 ( .A(n14094), .ZN(n10088) );
  NOR2_X1 U11622 ( .A1(n12464), .A2(n15728), .ZN(n12465) );
  NAND2_X1 U11623 ( .A1(n9970), .A2(n14470), .ZN(n14459) );
  NAND2_X1 U11624 ( .A1(n14146), .A2(n9971), .ZN(n9970) );
  AND2_X1 U11625 ( .A1(n13983), .A2(n14533), .ZN(n9971) );
  NAND2_X1 U11626 ( .A1(n10100), .A2(n10098), .ZN(n14147) );
  AND2_X1 U11627 ( .A1(n13616), .A2(n15764), .ZN(n12357) );
  INV_X1 U11628 ( .A(n14349), .ZN(n10073) );
  NAND2_X1 U11629 ( .A1(n12250), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12251) );
  NOR2_X1 U11630 ( .A1(n20934), .A2(n12251), .ZN(n12289) );
  INV_X1 U11631 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12127) );
  AND2_X1 U11632 ( .A1(n13209), .A2(n13213), .ZN(n13268) );
  NAND2_X1 U11633 ( .A1(n9831), .A2(n14563), .ZN(n14410) );
  NAND2_X1 U11634 ( .A1(n14470), .A2(n9829), .ZN(n9828) );
  INV_X1 U11635 ( .A(n9696), .ZN(n10090) );
  NAND2_X1 U11636 ( .A1(n13697), .A2(n13696), .ZN(n15900) );
  NAND2_X2 U11637 ( .A1(n9812), .A2(n15905), .ZN(n15902) );
  NAND2_X1 U11638 ( .A1(n15908), .A2(n15906), .ZN(n9812) );
  INV_X1 U11639 ( .A(n12076), .ZN(n9805) );
  NAND2_X1 U11640 ( .A1(n11919), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11972) );
  AND2_X1 U11641 ( .A1(n13121), .A2(n13120), .ZN(n15634) );
  AND2_X1 U11642 ( .A1(n20592), .A2(n20273), .ZN(n20504) );
  OR2_X1 U11643 ( .A1(n13020), .A2(n20185), .ZN(n20631) );
  INV_X1 U11644 ( .A(n20175), .ZN(n20273) );
  INV_X1 U11645 ( .A(n20744), .ZN(n20741) );
  AOI21_X1 U11646 ( .B1(n10755), .B2(n10754), .A(n10753), .ZN(n11007) );
  OR2_X1 U11647 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n10736), .ZN(n10741) );
  NOR2_X1 U11648 ( .A1(n10723), .A2(n10069), .ZN(n10068) );
  OR2_X1 U11649 ( .A1(n10670), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10718) );
  NAND2_X1 U11650 ( .A1(n10647), .A2(n13441), .ZN(n10735) );
  NAND2_X1 U11651 ( .A1(n10049), .A2(n10048), .ZN(n10047) );
  INV_X1 U11652 ( .A(n14962), .ZN(n10048) );
  NAND2_X1 U11653 ( .A1(n13516), .A2(n10020), .ZN(n10019) );
  INV_X1 U11654 ( .A(n13524), .ZN(n10020) );
  INV_X1 U11655 ( .A(n10269), .ZN(n12985) );
  INV_X1 U11656 ( .A(n11358), .ZN(n10931) );
  AND2_X1 U11657 ( .A1(n10880), .A2(n10879), .ZN(n15220) );
  NAND2_X1 U11658 ( .A1(n11351), .A2(n9698), .ZN(n11352) );
  AND2_X1 U11659 ( .A1(n15284), .A2(n11058), .ZN(n15259) );
  AND2_X1 U11660 ( .A1(n10035), .A2(n10034), .ZN(n10033) );
  INV_X1 U11661 ( .A(n15067), .ZN(n10034) );
  NAND2_X1 U11662 ( .A1(n9853), .A2(n15154), .ZN(n9852) );
  INV_X1 U11663 ( .A(n15153), .ZN(n9853) );
  AND2_X1 U11664 ( .A1(n11275), .A2(n11274), .ZN(n14645) );
  NAND2_X1 U11665 ( .A1(n16279), .A2(n9790), .ZN(n15365) );
  INV_X1 U11666 ( .A(n15363), .ZN(n10023) );
  INV_X1 U11667 ( .A(n15152), .ZN(n9855) );
  OAI21_X2 U11668 ( .B1(n15420), .B2(n15418), .A(n15416), .ZN(n15148) );
  INV_X1 U11669 ( .A(n15437), .ZN(n10132) );
  OR2_X1 U11670 ( .A1(n13896), .A2(n10643), .ZN(n10133) );
  NAND2_X1 U11671 ( .A1(n10805), .A2(n9863), .ZN(n9859) );
  AND2_X1 U11672 ( .A1(n10806), .A2(n10810), .ZN(n9861) );
  XNOR2_X1 U11673 ( .A(n11089), .B(n11088), .ZN(n13521) );
  INV_X1 U11674 ( .A(n11090), .ZN(n10018) );
  NAND2_X1 U11675 ( .A1(n12974), .A2(n19825), .ZN(n13054) );
  NOR2_X2 U11676 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19830) );
  NAND2_X1 U11677 ( .A1(n19831), .A2(n19832), .ZN(n19497) );
  OR2_X1 U11678 ( .A1(n19831), .A2(n19842), .ZN(n19597) );
  NAND2_X1 U11679 ( .A1(n19822), .A2(n19850), .ZN(n19626) );
  NOR2_X2 U11680 ( .A1(n13809), .A2(n13429), .ZN(n19261) );
  OR2_X1 U11681 ( .A1(n19831), .A2(n19832), .ZN(n19819) );
  NAND2_X1 U11682 ( .A1(n13426), .A2(n13425), .ZN(n19679) );
  INV_X1 U11683 ( .A(n19679), .ZN(n19442) );
  OAI21_X1 U11684 ( .B1(n9844), .B2(n9843), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9842) );
  OAI21_X1 U11685 ( .B1(n9848), .B2(n9847), .A(n9846), .ZN(n9845) );
  INV_X1 U11686 ( .A(n10261), .ZN(n9844) );
  AND2_X1 U11687 ( .A1(n15457), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11361) );
  NOR2_X1 U11688 ( .A1(n11703), .A2(n11702), .ZN(n18623) );
  AND2_X1 U11689 ( .A1(n9881), .A2(n9898), .ZN(n16606) );
  INV_X1 U11690 ( .A(n9883), .ZN(n9882) );
  AOI21_X1 U11691 ( .B1(n9898), .B2(n17547), .A(n16614), .ZN(n9883) );
  OR2_X1 U11692 ( .A1(n16628), .A2(n17547), .ZN(n9884) );
  NOR2_X1 U11693 ( .A1(n11444), .A2(n11441), .ZN(n11488) );
  INV_X1 U11694 ( .A(n11478), .ZN(n9994) );
  AOI21_X1 U11695 ( .B1(n17161), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A(n9993), .ZN(n9992) );
  AOI221_X1 U11696 ( .B1(n15474), .B2(n15473), .C1(n18620), .C2(n15473), .A(
        n18690), .ZN(n15712) );
  NOR2_X1 U11697 ( .A1(n18208), .A2(n11644), .ZN(n18645) );
  NOR2_X1 U11698 ( .A1(n16580), .A2(n16552), .ZN(n16392) );
  NAND3_X1 U11699 ( .A1(n9900), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16552) );
  AND2_X1 U11700 ( .A1(n18012), .A2(n18050), .ZN(n17679) );
  NOR2_X1 U11701 ( .A1(n17514), .A2(n17645), .ZN(n15686) );
  AND2_X1 U11702 ( .A1(n9933), .A2(n9699), .ZN(n11742) );
  OAI21_X1 U11703 ( .B1(n9699), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n9930), .ZN(n17513) );
  AND2_X1 U11704 ( .A1(n17540), .A2(n9793), .ZN(n9934) );
  NAND2_X1 U11705 ( .A1(n9936), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9935) );
  INV_X1 U11706 ( .A(n17541), .ZN(n9936) );
  NAND2_X1 U11707 ( .A1(n9728), .A2(n9935), .ZN(n9933) );
  OR2_X1 U11708 ( .A1(n17767), .A2(n17737), .ZN(n9997) );
  NOR2_X1 U11709 ( .A1(n17645), .A2(n17766), .ZN(n17744) );
  NAND2_X1 U11710 ( .A1(n11556), .A2(n18088), .ZN(n17765) );
  NAND2_X1 U11711 ( .A1(n11710), .A2(n11678), .ZN(n16356) );
  NOR2_X2 U11712 ( .A1(n11601), .A2(n11600), .ZN(n18188) );
  AND2_X1 U11713 ( .A1(n12639), .A2(n13213), .ZN(n20016) );
  NAND2_X1 U11714 ( .A1(n13180), .A2(n13080), .ZN(n14402) );
  INV_X1 U11715 ( .A(n13227), .ZN(n20185) );
  NAND2_X1 U11716 ( .A1(n19104), .A2(n19061), .ZN(n11375) );
  INV_X1 U11717 ( .A(n9858), .ZN(n10349) );
  NOR2_X1 U11718 ( .A1(n15453), .A2(n12980), .ZN(n19073) );
  OR2_X1 U11719 ( .A1(n10927), .A2(n11416), .ZN(n16098) );
  AND2_X1 U11720 ( .A1(n9720), .A2(n11403), .ZN(n16120) );
  NAND2_X1 U11721 ( .A1(n16199), .A2(n11389), .ZN(n9961) );
  NAND2_X1 U11722 ( .A1(n16198), .A2(n19225), .ZN(n9960) );
  AND2_X1 U11723 ( .A1(n16278), .A2(n12855), .ZN(n16268) );
  XNOR2_X1 U11724 ( .A(n11319), .B(n11318), .ZN(n16163) );
  NOR2_X1 U11725 ( .A1(n11414), .A2(n11312), .ZN(n11319) );
  XNOR2_X1 U11726 ( .A(n11376), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14142) );
  XNOR2_X1 U11727 ( .A(n9920), .B(n10965), .ZN(n11306) );
  NAND2_X1 U11728 ( .A1(n16202), .A2(n15389), .ZN(n9962) );
  INV_X1 U11729 ( .A(n16339), .ZN(n16314) );
  OR2_X1 U11730 ( .A1(n11304), .A2(n19862), .ZN(n16339) );
  OR2_X1 U11731 ( .A1(n11304), .A2(n11022), .ZN(n16327) );
  OR2_X1 U11732 ( .A1(n11304), .A2(n11303), .ZN(n16330) );
  INV_X1 U11733 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19855) );
  NOR2_X1 U11734 ( .A1(n19592), .A2(n19497), .ZN(n19555) );
  NOR2_X1 U11735 ( .A1(n18693), .A2(n18851), .ZN(n18838) );
  INV_X1 U11736 ( .A(n16569), .ZN(n9875) );
  NOR2_X1 U11737 ( .A1(n16571), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9876) );
  INV_X1 U11738 ( .A(n15581), .ZN(n17341) );
  NOR2_X1 U11739 ( .A1(n18219), .A2(n17369), .ZN(n17347) );
  INV_X1 U11740 ( .A(n18091), .ZN(n18031) );
  NOR2_X1 U11741 ( .A1(n9654), .A2(n18158), .ZN(n18153) );
  NAND2_X1 U11742 ( .A1(n12636), .A2(n20172), .ZN(n11906) );
  NAND2_X1 U11743 ( .A1(n12470), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12109) );
  NAND2_X1 U11744 ( .A1(n13113), .A2(n14594), .ZN(n11905) );
  NOR2_X1 U11745 ( .A1(n11916), .A2(n11898), .ZN(n9808) );
  AND2_X1 U11746 ( .A1(n13000), .A2(n9677), .ZN(n10299) );
  NAND2_X1 U11747 ( .A1(n10398), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14759) );
  NAND2_X1 U11748 ( .A1(n10398), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n14752) );
  OAI21_X1 U11749 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18807), .A(
        n11682), .ZN(n11683) );
  NAND2_X1 U11750 ( .A1(n20635), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12595) );
  INV_X1 U11751 ( .A(n12610), .ZN(n12584) );
  NAND2_X1 U11752 ( .A1(n12611), .A2(n12585), .ZN(n12587) );
  AND2_X1 U11753 ( .A1(n12587), .A2(n12586), .ZN(n12589) );
  NOR2_X1 U11754 ( .A1(n12631), .A2(n12602), .ZN(n12624) );
  NAND2_X1 U11755 ( .A1(n12470), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n12343) );
  NAND2_X1 U11756 ( .A1(n12470), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n12311) );
  NAND2_X1 U11757 ( .A1(n12470), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12277) );
  OR2_X1 U11758 ( .A1(n12100), .A2(n12099), .ZN(n13682) );
  NAND2_X1 U11759 ( .A1(n9972), .A2(n12643), .ZN(n12645) );
  INV_X1 U11760 ( .A(n11941), .ZN(n13234) );
  INV_X1 U11761 ( .A(n11958), .ZN(n9945) );
  OR2_X1 U11762 ( .A1(n11956), .A2(n11955), .ZN(n13233) );
  INV_X1 U11763 ( .A(n20136), .ZN(n13111) );
  NAND2_X1 U11764 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11757) );
  NAND2_X1 U11765 ( .A1(n11884), .A2(n20124), .ZN(n11904) );
  NAND2_X1 U11766 ( .A1(n12958), .A2(n14168), .ZN(n13128) );
  NAND3_X1 U11767 ( .A1(n9664), .A2(n10140), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10391) );
  NAND2_X1 U11768 ( .A1(n10050), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n14901) );
  NAND2_X1 U11769 ( .A1(n10050), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n14908) );
  NAND2_X1 U11770 ( .A1(n10050), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n14883) );
  NAND2_X1 U11771 ( .A1(n10050), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n14889) );
  NAND2_X1 U11772 ( .A1(n10050), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n14863) );
  NAND2_X1 U11773 ( .A1(n10050), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14869) );
  NAND2_X1 U11774 ( .A1(n10050), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n14843) );
  NAND2_X1 U11775 ( .A1(n10050), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14849) );
  NAND2_X1 U11776 ( .A1(n10050), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n14821) );
  NAND2_X1 U11777 ( .A1(n10050), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14828) );
  NAND2_X1 U11778 ( .A1(n10050), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14802) );
  NAND2_X1 U11779 ( .A1(n10398), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n14796) );
  INV_X1 U11780 ( .A(n10354), .ZN(n10150) );
  INV_X1 U11781 ( .A(n10141), .ZN(n10315) );
  INV_X1 U11782 ( .A(n15129), .ZN(n10122) );
  OAI21_X1 U11783 ( .B1(n11099), .B2(n11027), .A(n10589), .ZN(n10596) );
  NOR2_X1 U11784 ( .A1(n10415), .A2(n10414), .ZN(n10480) );
  NOR2_X1 U11785 ( .A1(n9865), .A2(n9864), .ZN(n9919) );
  INV_X1 U11786 ( .A(n10423), .ZN(n9864) );
  NOR2_X1 U11787 ( .A1(n10402), .A2(n10057), .ZN(n10510) );
  NAND2_X1 U11788 ( .A1(n10376), .A2(n10375), .ZN(n10410) );
  NAND2_X1 U11789 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18820), .ZN(
        n11442) );
  NOR2_X1 U11790 ( .A1(n11442), .A2(n11445), .ZN(n11523) );
  NOR2_X1 U11791 ( .A1(n14319), .A2(n14326), .ZN(n10085) );
  AOI21_X1 U11792 ( .B1(n11820), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A(n9837), .ZN(n12241) );
  INV_X1 U11793 ( .A(n13963), .ZN(n12248) );
  NOR2_X1 U11794 ( .A1(n10083), .A2(n10081), .ZN(n10080) );
  INV_X1 U11795 ( .A(n13887), .ZN(n10081) );
  NAND2_X1 U11796 ( .A1(n12068), .A2(n12067), .ZN(n13024) );
  OR2_X1 U11797 ( .A1(n14073), .A2(n9982), .ZN(n9981) );
  INV_X1 U11798 ( .A(n14057), .ZN(n9982) );
  NAND2_X1 U11799 ( .A1(n9968), .A2(n9967), .ZN(n14052) );
  NOR2_X1 U11800 ( .A1(n13764), .A2(n13740), .ZN(n9979) );
  INV_X1 U11801 ( .A(n12132), .ZN(n12133) );
  OR2_X1 U11802 ( .A1(n12023), .A2(n12022), .ZN(n13708) );
  INV_X1 U11803 ( .A(n13672), .ZN(n10094) );
  NAND2_X1 U11804 ( .A1(n12652), .A2(n12649), .ZN(n12735) );
  NAND2_X1 U11805 ( .A1(n13350), .A2(n10089), .ZN(n9941) );
  OR2_X1 U11806 ( .A1(n11878), .A2(n20804), .ZN(n11963) );
  INV_X1 U11807 ( .A(n12626), .ZN(n12621) );
  NAND2_X1 U11808 ( .A1(n12056), .A2(n20804), .ZN(n12048) );
  NOR2_X1 U11809 ( .A1(n9823), .A2(n11942), .ZN(n9820) );
  INV_X1 U11810 ( .A(n11942), .ZN(n9821) );
  OR2_X1 U11811 ( .A1(n11983), .A2(n11982), .ZN(n13361) );
  NAND2_X1 U11812 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11844) );
  NAND2_X1 U11813 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11859) );
  NAND2_X1 U11814 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11758) );
  NAND2_X1 U11815 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11779) );
  OAI21_X1 U11816 ( .B1(n20899), .B2(n13172), .A(n14614), .ZN(n20103) );
  AND2_X1 U11817 ( .A1(n12960), .A2(n12959), .ZN(n13114) );
  INV_X1 U11818 ( .A(n10515), .ZN(n10756) );
  NAND2_X1 U11819 ( .A1(n10056), .A2(n10055), .ZN(n10770) );
  NAND2_X1 U11820 ( .A1(n10984), .A2(n10750), .ZN(n10055) );
  NAND2_X1 U11821 ( .A1(n10510), .A2(n10983), .ZN(n10056) );
  AND2_X1 U11822 ( .A1(n10548), .A2(n10547), .ZN(n10755) );
  OR2_X1 U11823 ( .A1(n10546), .A2(n10545), .ZN(n10548) );
  OR2_X1 U11824 ( .A1(n10702), .A2(n10700), .ZN(n10699) );
  NOR2_X1 U11825 ( .A1(n10062), .A2(n10668), .ZN(n10061) );
  INV_X1 U11826 ( .A(n10063), .ZN(n10062) );
  NAND2_X1 U11827 ( .A1(n10662), .A2(n10063), .ZN(n10688) );
  OR2_X1 U11828 ( .A1(n10646), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10649) );
  NOR2_X1 U11829 ( .A1(n10649), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10653) );
  NOR2_X1 U11830 ( .A1(n10636), .A2(n10059), .ZN(n10058) );
  INV_X1 U11831 ( .A(n10590), .ZN(n10059) );
  NOR2_X1 U11832 ( .A1(n10512), .A2(n10511), .ZN(n10550) );
  CLKBUF_X1 U11833 ( .A(n10184), .Z(n14928) );
  NAND2_X1 U11834 ( .A1(n14902), .A2(n10052), .ZN(n10051) );
  NAND2_X1 U11835 ( .A1(n10050), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10052) );
  AOI21_X1 U11836 ( .B1(n14794), .B2(n9925), .A(n9789), .ZN(n9923) );
  AND2_X1 U11837 ( .A1(n13551), .A2(n10170), .ZN(n10045) );
  OR2_X1 U11838 ( .A1(n13280), .A2(n19243), .ZN(n13056) );
  NOR2_X1 U11839 ( .A1(n16216), .A2(n10004), .ZN(n10003) );
  AND2_X1 U11840 ( .A1(n10130), .A2(n10131), .ZN(n10129) );
  INV_X1 U11841 ( .A(n16226), .ZN(n10130) );
  NAND2_X1 U11842 ( .A1(n10129), .A2(n10643), .ZN(n10127) );
  OR2_X1 U11843 ( .A1(n18957), .A2(n10640), .ZN(n10666) );
  NAND2_X1 U11844 ( .A1(n10106), .A2(n13194), .ZN(n10105) );
  INV_X1 U11845 ( .A(n13571), .ZN(n10106) );
  NAND2_X1 U11846 ( .A1(n10342), .A2(n10341), .ZN(n10830) );
  XNOR2_X1 U11847 ( .A(n10830), .B(n10831), .ZN(n10832) );
  NAND3_X1 U11848 ( .A1(n10347), .A2(n10324), .A3(n10338), .ZN(n10325) );
  AND3_X1 U11849 ( .A1(n10479), .A2(n10478), .A3(n10477), .ZN(n10780) );
  NAND2_X1 U11850 ( .A1(n10054), .A2(n10053), .ZN(n11362) );
  INV_X1 U11851 ( .A(n10958), .ZN(n10053) );
  OAI21_X1 U11852 ( .B1(n10952), .B2(n10139), .A(n10169), .ZN(n10138) );
  NOR2_X1 U11853 ( .A1(n10147), .A2(n15270), .ZN(n10146) );
  INV_X1 U11854 ( .A(n10148), .ZN(n10147) );
  NOR2_X1 U11855 ( .A1(n21079), .A2(n15297), .ZN(n10148) );
  INV_X1 U11856 ( .A(n15157), .ZN(n10143) );
  AND2_X1 U11857 ( .A1(n10152), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9873) );
  AND2_X1 U11858 ( .A1(n10890), .A2(n10889), .ZN(n14049) );
  AND2_X1 U11859 ( .A1(n10153), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10152) );
  AND2_X1 U11860 ( .A1(n15370), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10153) );
  AND2_X1 U11861 ( .A1(n15230), .A2(n9762), .ZN(n10131) );
  INV_X1 U11862 ( .A(n16246), .ZN(n9955) );
  INV_X1 U11863 ( .A(n13904), .ZN(n10026) );
  INV_X1 U11864 ( .A(n13572), .ZN(n10103) );
  OR2_X1 U11865 ( .A1(n10544), .A2(n10543), .ZN(n11095) );
  AND3_X1 U11866 ( .A1(n10457), .A2(n10456), .A3(n10455), .ZN(n11081) );
  INV_X1 U11867 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10173) );
  INV_X1 U11868 ( .A(n11027), .ZN(n10274) );
  NAND2_X1 U11869 ( .A1(n14673), .A2(n10357), .ZN(n10358) );
  INV_X1 U11870 ( .A(n10255), .ZN(n9848) );
  NOR2_X1 U11871 ( .A1(n9898), .A2(n17511), .ZN(n9888) );
  NAND2_X1 U11872 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18796), .ZN(
        n11447) );
  INV_X1 U11873 ( .A(n11494), .ZN(n16938) );
  OR2_X1 U11874 ( .A1(n11442), .A2(n11439), .ZN(n10156) );
  NOR2_X1 U11875 ( .A1(n16938), .A2(n15529), .ZN(n9993) );
  NAND2_X1 U11876 ( .A1(n11494), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n9989) );
  INV_X1 U11877 ( .A(n18212), .ZN(n11644) );
  NOR2_X1 U11878 ( .A1(n15685), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16357) );
  NAND2_X1 U11879 ( .A1(n17606), .A2(n17592), .ZN(n17593) );
  OR2_X1 U11880 ( .A1(n9997), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9996) );
  NAND2_X1 U11881 ( .A1(n17788), .A2(n11551), .ZN(n11553) );
  NAND2_X1 U11882 ( .A1(n17817), .A2(n11546), .ZN(n11549) );
  INV_X1 U11883 ( .A(n11488), .ZN(n14087) );
  NAND2_X1 U11884 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18659) );
  OAI21_X1 U11885 ( .B1(n11663), .B2(n11662), .A(n18621), .ZN(n11665) );
  NOR2_X1 U11886 ( .A1(n11660), .A2(n11666), .ZN(n14078) );
  INV_X1 U11887 ( .A(n13076), .ZN(n9838) );
  AND2_X1 U11888 ( .A1(n14126), .A2(n12635), .ZN(n13242) );
  NOR2_X1 U11889 ( .A1(n15675), .A2(n9975), .ZN(n14330) );
  AND2_X1 U11890 ( .A1(n13737), .A2(n9777), .ZN(n13997) );
  AOI21_X1 U11891 ( .B1(n13673), .B2(n13021), .A(n12106), .ZN(n13393) );
  INV_X1 U11892 ( .A(n19871), .ZN(n13213) );
  AND2_X1 U11893 ( .A1(n12506), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12507) );
  NAND2_X1 U11894 ( .A1(n12512), .A2(n12511), .ZN(n14235) );
  AND2_X1 U11895 ( .A1(n12467), .A2(n12466), .ZN(n14305) );
  AND2_X1 U11896 ( .A1(n12446), .A2(n12445), .ZN(n14313) );
  NOR2_X1 U11897 ( .A1(n12426), .A2(n14464), .ZN(n12427) );
  INV_X1 U11898 ( .A(n14335), .ZN(n10077) );
  AND2_X1 U11899 ( .A1(n12339), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12340) );
  NAND2_X1 U11900 ( .A1(n12340), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12374) );
  NAND2_X1 U11901 ( .A1(n12289), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12306) );
  AND2_X1 U11902 ( .A1(n12269), .A2(n12268), .ZN(n14070) );
  AND2_X1 U11903 ( .A1(n12233), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12250) );
  NOR2_X1 U11904 ( .A1(n12229), .A2(n15805), .ZN(n12233) );
  NOR2_X1 U11905 ( .A1(n9712), .A2(n9792), .ZN(n10078) );
  AND2_X1 U11906 ( .A1(n12190), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12191) );
  NOR2_X1 U11907 ( .A1(n12173), .A2(n19899), .ZN(n12190) );
  AOI21_X1 U11908 ( .B1(n12171), .B2(n13616), .A(n12170), .ZN(n13733) );
  CLKBUF_X1 U11909 ( .A(n13609), .Z(n13610) );
  NOR2_X1 U11910 ( .A1(n12124), .A2(n12127), .ZN(n12137) );
  NAND2_X1 U11911 ( .A1(n12103), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12124) );
  NAND2_X1 U11912 ( .A1(n12130), .A2(n12129), .ZN(n13416) );
  AND2_X1 U11913 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12080), .ZN(
        n12103) );
  INV_X1 U11914 ( .A(n13398), .ZN(n12089) );
  NAND2_X1 U11915 ( .A1(n13087), .A2(n12075), .ZN(n13103) );
  AOI21_X1 U11916 ( .B1(n12073), .B2(n12264), .A(n10072), .ZN(n10071) );
  INV_X1 U11917 ( .A(n12075), .ZN(n10072) );
  INV_X1 U11918 ( .A(n12264), .ZN(n13021) );
  NOR2_X1 U11919 ( .A1(n14155), .A2(n9829), .ZN(n9833) );
  NOR2_X1 U11920 ( .A1(n14309), .A2(n9983), .ZN(n14224) );
  OR3_X1 U11921 ( .A1(n12737), .A2(n9984), .A3(n14225), .ZN(n9983) );
  INV_X1 U11922 ( .A(n9972), .ZN(n12738) );
  NOR3_X1 U11923 ( .A1(n14309), .A2(n12737), .A3(n14247), .ZN(n14241) );
  NAND2_X1 U11924 ( .A1(n15836), .A2(n9811), .ZN(n14427) );
  NAND2_X1 U11925 ( .A1(n14152), .A2(n14148), .ZN(n9811) );
  INV_X1 U11926 ( .A(n9817), .ZN(n9816) );
  OAI21_X1 U11927 ( .B1(n14460), .B2(n14534), .A(n14151), .ZN(n9817) );
  NOR2_X1 U11928 ( .A1(n14309), .A2(n14247), .ZN(n14246) );
  INV_X1 U11929 ( .A(n9975), .ZN(n9974) );
  NOR3_X1 U11930 ( .A1(n15675), .A2(n9975), .A3(n12725), .ZN(n14323) );
  OR2_X1 U11931 ( .A1(n9716), .A2(n14341), .ZN(n15675) );
  NOR2_X1 U11932 ( .A1(n15675), .A2(n12719), .ZN(n15679) );
  NAND2_X1 U11933 ( .A1(n10100), .A2(n10099), .ZN(n14471) );
  AND2_X1 U11934 ( .A1(n9966), .A2(n9969), .ZN(n15861) );
  NOR2_X1 U11935 ( .A1(n14072), .A2(n9981), .ZN(n14272) );
  XNOR2_X1 U11936 ( .A(n14470), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14056) );
  NOR2_X1 U11937 ( .A1(n14072), .A2(n14073), .ZN(n14071) );
  NAND2_X1 U11938 ( .A1(n13997), .A2(n13996), .ZN(n13995) );
  OR2_X1 U11939 ( .A1(n13995), .A2(n13939), .ZN(n14072) );
  NAND2_X1 U11940 ( .A1(n13737), .A2(n9979), .ZN(n13889) );
  NAND2_X1 U11941 ( .A1(n13737), .A2(n12680), .ZN(n13765) );
  AND2_X1 U11942 ( .A1(n12678), .A2(n12677), .ZN(n13612) );
  OR2_X1 U11943 ( .A1(n16060), .A2(n12674), .ZN(n16043) );
  INV_X1 U11944 ( .A(n14517), .ZN(n16032) );
  NOR2_X1 U11945 ( .A1(n13386), .A2(n13372), .ZN(n16058) );
  OR2_X1 U11946 ( .A1(n13384), .A2(n13383), .ZN(n13386) );
  OR2_X1 U11947 ( .A1(n13252), .A2(n13251), .ZN(n13384) );
  NOR2_X1 U11948 ( .A1(n13260), .A2(n14593), .ZN(n15668) );
  NAND2_X1 U11949 ( .A1(n9825), .A2(n11958), .ZN(n13220) );
  NAND2_X1 U11950 ( .A1(n9946), .A2(n20804), .ZN(n9825) );
  INV_X1 U11951 ( .A(n14594), .ZN(n14126) );
  INV_X1 U11952 ( .A(n15628), .ZN(n14593) );
  OR2_X1 U11953 ( .A1(n13353), .A2(n20425), .ZN(n20552) );
  OR2_X1 U11954 ( .A1(n13020), .A2(n13227), .ZN(n20582) );
  AND2_X1 U11955 ( .A1(n20507), .A2(n20273), .ZN(n20686) );
  NAND4_X1 U11956 ( .A1(n11806), .A2(n11805), .A3(n11804), .A4(n11803), .ZN(
        n11807) );
  AND2_X1 U11957 ( .A1(n11802), .A2(n11801), .ZN(n11804) );
  NAND2_X1 U11958 ( .A1(n13020), .A2(n20185), .ZN(n20681) );
  INV_X1 U11959 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20746) );
  INV_X1 U11960 ( .A(n13209), .ZN(n15656) );
  NAND2_X1 U11961 ( .A1(n21068), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15652) );
  OR2_X1 U11962 ( .A1(n19859), .A2(n10765), .ZN(n10776) );
  NOR2_X1 U11963 ( .A1(n10957), .A2(n10956), .ZN(n10054) );
  AND2_X1 U11964 ( .A1(n9707), .A2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10010) );
  NAND2_X1 U11965 ( .A1(n11365), .A2(n10743), .ZN(n10957) );
  NAND2_X1 U11966 ( .A1(n11336), .A2(n9707), .ZN(n11330) );
  NAND2_X1 U11967 ( .A1(n10716), .A2(n9710), .ZN(n10736) );
  NAND2_X1 U11968 ( .A1(n10741), .A2(n10735), .ZN(n11365) );
  NOR2_X1 U11969 ( .A1(n10699), .A2(n10697), .ZN(n10695) );
  NAND2_X1 U11970 ( .A1(n10662), .A2(n10661), .ZN(n10686) );
  NAND2_X1 U11971 ( .A1(n10591), .A2(n10590), .ZN(n10637) );
  AND3_X1 U11972 ( .A1(n14703), .A2(n14702), .A3(n14701), .ZN(n16171) );
  NAND2_X1 U11973 ( .A1(n15194), .A2(n15193), .ZN(n15196) );
  AND2_X1 U11974 ( .A1(n10883), .A2(n10882), .ZN(n13881) );
  AND2_X1 U11975 ( .A1(n10864), .A2(n10863), .ZN(n13407) );
  NOR2_X1 U11976 ( .A1(n9927), .A2(n13345), .ZN(n9926) );
  INV_X1 U11977 ( .A(n13281), .ZN(n9927) );
  NAND2_X1 U11978 ( .A1(n10050), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14920) );
  NAND2_X1 U11979 ( .A1(n9929), .A2(n14878), .ZN(n9928) );
  NOR2_X1 U11980 ( .A1(n14963), .A2(n14962), .ZN(n14961) );
  XNOR2_X1 U11981 ( .A(n14838), .B(n14839), .ZN(n14968) );
  NAND2_X1 U11982 ( .A1(n10039), .A2(n14984), .ZN(n10038) );
  INV_X1 U11983 ( .A(n10040), .ZN(n10039) );
  AND3_X1 U11984 ( .A1(n13836), .A2(n13835), .A3(n13834), .ZN(n13861) );
  INV_X1 U11985 ( .A(n11006), .ZN(n12872) );
  NOR2_X1 U11986 ( .A1(n11369), .A2(n10979), .ZN(n13657) );
  OAI21_X1 U11987 ( .B1(n12773), .B2(n12772), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12843) );
  INV_X1 U11988 ( .A(n12843), .ZN(n13809) );
  AND2_X1 U11989 ( .A1(n10920), .A2(n10919), .ZN(n14954) );
  NOR2_X1 U11990 ( .A1(n9720), .A2(n14954), .ZN(n14953) );
  NAND2_X1 U11991 ( .A1(n11336), .A2(n10011), .ZN(n11331) );
  NAND2_X1 U11992 ( .A1(n11336), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11334) );
  AND2_X1 U11993 ( .A1(n10910), .A2(n10909), .ZN(n14977) );
  NOR2_X1 U11994 ( .A1(n15125), .A2(n14977), .ZN(n14979) );
  OR2_X1 U11995 ( .A1(n15143), .A2(n15123), .ZN(n15125) );
  AND2_X1 U11996 ( .A1(n15194), .A2(n10110), .ZN(n15141) );
  AND2_X1 U11997 ( .A1(n9758), .A2(n10111), .ZN(n10110) );
  INV_X1 U11998 ( .A(n14986), .ZN(n10111) );
  AND2_X1 U11999 ( .A1(n10893), .A2(n10892), .ZN(n14633) );
  NAND2_X1 U12000 ( .A1(n15194), .A2(n10113), .ZN(n14634) );
  NAND2_X1 U12001 ( .A1(n15194), .A2(n9758), .ZN(n14987) );
  AND2_X1 U12002 ( .A1(n9711), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10006) );
  NAND2_X1 U12003 ( .A1(n11353), .A2(n10007), .ZN(n11356) );
  NAND2_X1 U12004 ( .A1(n11353), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11355) );
  INV_X1 U12005 ( .A(n15220), .ZN(n10115) );
  NAND2_X1 U12006 ( .A1(n13446), .A2(n9755), .ZN(n15221) );
  NAND2_X1 U12007 ( .A1(n11351), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11350) );
  NOR2_X1 U12008 ( .A1(n10861), .A2(n11348), .ZN(n11351) );
  NAND2_X1 U12009 ( .A1(n11349), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11348) );
  NOR2_X1 U12010 ( .A1(n11346), .A2(n10825), .ZN(n11349) );
  NOR2_X1 U12011 ( .A1(n11344), .A2(n10847), .ZN(n11347) );
  NAND2_X1 U12012 ( .A1(n11347), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11346) );
  AND2_X1 U12013 ( .A1(n10856), .A2(n10855), .ZN(n16241) );
  NOR2_X1 U12014 ( .A1(n13303), .A2(n16241), .ZN(n16242) );
  AND2_X1 U12015 ( .A1(n10846), .A2(n10845), .ZN(n13310) );
  NOR2_X1 U12016 ( .A1(n11342), .A2(n10838), .ZN(n11345) );
  OR2_X1 U12017 ( .A1(n13572), .A2(n10105), .ZN(n13309) );
  NOR2_X1 U12018 ( .A1(n13572), .A2(n13571), .ZN(n13193) );
  NAND2_X1 U12019 ( .A1(n11343), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11342) );
  NAND2_X1 U12020 ( .A1(n11416), .A2(n11415), .ZN(n11414) );
  INV_X1 U12021 ( .A(n11424), .ZN(n9921) );
  NAND2_X1 U12022 ( .A1(n10030), .A2(n10029), .ZN(n10027) );
  OR3_X1 U12023 ( .A1(n16129), .A2(n10640), .A3(n21079), .ZN(n15101) );
  AOI21_X1 U12024 ( .B1(n9916), .B2(n9914), .A(n9913), .ZN(n9912) );
  INV_X1 U12025 ( .A(n9916), .ZN(n9915) );
  INV_X1 U12026 ( .A(n10715), .ZN(n9914) );
  NAND2_X1 U12027 ( .A1(n15136), .A2(n15137), .ZN(n10123) );
  OR2_X1 U12028 ( .A1(n15356), .A2(n11045), .ZN(n15296) );
  OR2_X1 U12029 ( .A1(n10720), .A2(n15320), .ZN(n15138) );
  AND2_X1 U12030 ( .A1(n11052), .A2(n13569), .ZN(n15400) );
  AND2_X1 U12031 ( .A1(n15211), .A2(n10152), .ZN(n15179) );
  AND2_X1 U12032 ( .A1(n11273), .A2(n11272), .ZN(n15363) );
  NAND2_X1 U12033 ( .A1(n16279), .A2(n15384), .ZN(n15590) );
  AND2_X1 U12034 ( .A1(n13446), .A2(n10116), .ZN(n13649) );
  NAND2_X1 U12035 ( .A1(n13446), .A2(n13445), .ZN(n13555) );
  AND2_X1 U12036 ( .A1(n13406), .A2(n10865), .ZN(n13408) );
  INV_X1 U12037 ( .A(n13407), .ZN(n10865) );
  NAND2_X1 U12038 ( .A1(n10133), .A2(n10131), .ZN(n16225) );
  AND2_X1 U12039 ( .A1(n13905), .A2(n9705), .ZN(n16309) );
  NAND2_X1 U12040 ( .A1(n13895), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9954) );
  NAND2_X1 U12041 ( .A1(n13905), .A2(n13904), .ZN(n16310) );
  NAND2_X1 U12042 ( .A1(n10801), .A2(n10800), .ZN(n13867) );
  NAND2_X1 U12043 ( .A1(n13752), .A2(n11103), .ZN(n13870) );
  NAND2_X1 U12044 ( .A1(n10526), .A2(n13579), .ZN(n13564) );
  NAND2_X1 U12045 ( .A1(n10484), .A2(n10483), .ZN(n10791) );
  NAND2_X1 U12046 ( .A1(n10485), .A2(n10791), .ZN(n10514) );
  OAI211_X1 U12047 ( .C1(n11074), .C2(n11242), .A(n11085), .B(n11073), .ZN(
        n12982) );
  AND2_X1 U12048 ( .A1(n12981), .A2(n12982), .ZN(n12984) );
  OR2_X1 U12049 ( .A1(n11304), .A2(n11044), .ZN(n15598) );
  OR2_X1 U12050 ( .A1(n11304), .A2(n13295), .ZN(n14192) );
  OR3_X1 U12051 ( .A1(n19267), .A2(n19289), .A3(n19593), .ZN(n19271) );
  NAND2_X1 U12052 ( .A1(n19269), .A2(n19850), .ZN(n19407) );
  NAND2_X1 U12053 ( .A1(n19269), .A2(n19073), .ZN(n19435) );
  NAND2_X1 U12054 ( .A1(n9905), .A2(n13597), .ZN(n13602) );
  OAI21_X1 U12055 ( .B1(n10190), .B2(n10189), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10197) );
  INV_X1 U12056 ( .A(n10774), .ZN(n13473) );
  NOR2_X1 U12057 ( .A1(n18196), .A2(n11660), .ZN(n11676) );
  NOR2_X1 U12058 ( .A1(n9681), .A2(n14079), .ZN(n18621) );
  INV_X1 U12059 ( .A(n17511), .ZN(n9889) );
  INV_X1 U12060 ( .A(n9890), .ZN(n16581) );
  OAI21_X1 U12061 ( .B1(n16605), .B2(n9756), .A(n9886), .ZN(n9890) );
  NOR2_X1 U12062 ( .A1(n9887), .A2(n16582), .ZN(n9886) );
  NOR3_X1 U12063 ( .A1(n16835), .A2(n9888), .A3(n9889), .ZN(n9887) );
  OR2_X1 U12064 ( .A1(n9898), .A2(n17575), .ZN(n9897) );
  OR2_X1 U12065 ( .A1(n16657), .A2(n9743), .ZN(n9896) );
  OR2_X1 U12066 ( .A1(n16657), .A2(n16658), .ZN(n9899) );
  NOR2_X1 U12067 ( .A1(n17378), .A2(n17377), .ZN(n17380) );
  NOR2_X1 U12068 ( .A1(n18690), .A2(n18623), .ZN(n17440) );
  NAND2_X1 U12069 ( .A1(n9902), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9901) );
  INV_X1 U12070 ( .A(n9903), .ZN(n9902) );
  NOR2_X1 U12071 ( .A1(n17535), .A2(n9903), .ZN(n17493) );
  NOR2_X1 U12072 ( .A1(n17535), .A2(n17536), .ZN(n17524) );
  NAND2_X1 U12073 ( .A1(n17636), .A2(n9708), .ZN(n17582) );
  NOR2_X1 U12074 ( .A1(n17613), .A2(n9894), .ZN(n9893) );
  INV_X1 U12075 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9894) );
  NAND2_X1 U12076 ( .A1(n17636), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17612) );
  NOR2_X1 U12077 ( .A1(n17650), .A2(n17651), .ZN(n17636) );
  NAND2_X1 U12078 ( .A1(n17674), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17650) );
  NOR2_X1 U12079 ( .A1(n17721), .A2(n17692), .ZN(n17674) );
  AOI21_X1 U12080 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16366), .A(
        n18566), .ZN(n17691) );
  NAND2_X1 U12081 ( .A1(n17775), .A2(n17690), .ZN(n17721) );
  INV_X1 U12082 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17761) );
  XNOR2_X1 U12083 ( .A(n11549), .B(n11548), .ZN(n17802) );
  INV_X1 U12084 ( .A(n11547), .ZN(n11548) );
  INV_X1 U12085 ( .A(n16738), .ZN(n17794) );
  NAND2_X1 U12086 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17809) );
  NOR2_X1 U12087 ( .A1(n17845), .A2(n17810), .ZN(n17793) );
  NOR2_X1 U12088 ( .A1(n18192), .A2(n16524), .ZN(n16375) );
  NAND2_X1 U12089 ( .A1(n9939), .A2(n16359), .ZN(n15688) );
  NAND2_X1 U12090 ( .A1(n16357), .A2(n17645), .ZN(n9939) );
  NAND2_X1 U12091 ( .A1(n15688), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16358) );
  NOR3_X1 U12092 ( .A1(n17552), .A2(n17566), .A3(n17918), .ZN(n17541) );
  NAND2_X1 U12093 ( .A1(n17606), .A2(n9986), .ZN(n17553) );
  NAND2_X1 U12094 ( .A1(n9987), .A2(n9757), .ZN(n9986) );
  NAND2_X1 U12095 ( .A1(n17577), .A2(n17898), .ZN(n9987) );
  NAND2_X1 U12096 ( .A1(n17593), .A2(n9937), .ZN(n17566) );
  AND2_X1 U12097 ( .A1(n11560), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9937) );
  NAND2_X1 U12098 ( .A1(n17634), .A2(n17645), .ZN(n17606) );
  AND2_X1 U12099 ( .A1(n11559), .A2(n11558), .ZN(n17635) );
  AOI21_X1 U12100 ( .B1(n17920), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n9704), .ZN(n11558) );
  NAND2_X1 U12101 ( .A1(n17635), .A2(n17979), .ZN(n17634) );
  NOR2_X1 U12102 ( .A1(n17647), .A2(n17728), .ZN(n17897) );
  OR2_X1 U12103 ( .A1(n17765), .A2(n9995), .ZN(n17666) );
  OR2_X1 U12104 ( .A1(n9996), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9995) );
  NAND2_X1 U12105 ( .A1(n11670), .A2(n11669), .ZN(n18638) );
  NAND2_X1 U12106 ( .A1(n11739), .A2(n17756), .ZN(n18049) );
  NOR2_X1 U12107 ( .A1(n17765), .A2(n17767), .ZN(n17743) );
  XNOR2_X1 U12108 ( .A(n11553), .B(n9988), .ZN(n17781) );
  INV_X1 U12109 ( .A(n11554), .ZN(n9988) );
  NAND2_X1 U12110 ( .A1(n17781), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17780) );
  NOR2_X1 U12111 ( .A1(n17778), .A2(n17777), .ZN(n17776) );
  XNOR2_X1 U12112 ( .A(n11542), .B(n11541), .ZN(n17826) );
  INV_X1 U12113 ( .A(n11540), .ZN(n11541) );
  NAND2_X1 U12114 ( .A1(n17826), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n17825) );
  XNOR2_X1 U12115 ( .A(n11538), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17837) );
  INV_X1 U12116 ( .A(n11665), .ZN(n18658) );
  NOR2_X1 U12117 ( .A1(n18853), .A2(n15474), .ZN(n18635) );
  INV_X1 U12118 ( .A(n18659), .ZN(n18641) );
  NOR2_X1 U12119 ( .A1(n11641), .A2(n11640), .ZN(n18200) );
  NOR2_X1 U12120 ( .A1(n18288), .A2(n18334), .ZN(n18215) );
  NOR2_X1 U12121 ( .A1(n11621), .A2(n11620), .ZN(n18208) );
  OAI22_X1 U12122 ( .A1(n18625), .A2(n16356), .B1(n18620), .B2(n18627), .ZN(
        n18680) );
  INV_X1 U12123 ( .A(n19979), .ZN(n19935) );
  OR2_X1 U12124 ( .A1(n20894), .A2(n13618), .ZN(n19976) );
  INV_X1 U12125 ( .A(n19985), .ZN(n19940) );
  INV_X1 U12126 ( .A(n19965), .ZN(n19961) );
  INV_X1 U12127 ( .A(n19937), .ZN(n19991) );
  INV_X1 U12128 ( .A(n20005), .ZN(n20012) );
  INV_X1 U12129 ( .A(n14415), .ZN(n14355) );
  INV_X1 U12130 ( .A(n14404), .ZN(n14398) );
  INV_X1 U12131 ( .A(n14402), .ZN(n14397) );
  OR2_X1 U12132 ( .A1(n14397), .A2(n13081), .ZN(n14076) );
  NAND2_X1 U12133 ( .A1(n13032), .A2(n13031), .ZN(n13180) );
  XNOR2_X1 U12134 ( .A(n13625), .B(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14163) );
  NAND2_X1 U12135 ( .A1(n14221), .A2(n14157), .ZN(n14162) );
  INV_X1 U12136 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n14464) );
  INV_X1 U12137 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15774) );
  NAND2_X1 U12138 ( .A1(n19877), .A2(n13271), .ZN(n15918) );
  AND2_X1 U12139 ( .A1(n13269), .A2(n20741), .ZN(n15909) );
  INV_X1 U12140 ( .A(n15918), .ZN(n20076) );
  AND2_X1 U12141 ( .A1(n13268), .A2(n15642), .ZN(n20074) );
  XNOR2_X1 U12142 ( .A(n9965), .B(n14598), .ZN(n14541) );
  NAND2_X1 U12143 ( .A1(n9836), .A2(n9835), .ZN(n9965) );
  NAND2_X1 U12144 ( .A1(n9832), .A2(n9766), .ZN(n9835) );
  NAND2_X1 U12145 ( .A1(n9830), .A2(n9769), .ZN(n9836) );
  XNOR2_X1 U12146 ( .A(n9947), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14550) );
  NAND2_X1 U12147 ( .A1(n9834), .A2(n14535), .ZN(n9948) );
  NAND2_X1 U12148 ( .A1(n9830), .A2(n9828), .ZN(n14417) );
  NOR2_X1 U12149 ( .A1(n13260), .A2(n13250), .ZN(n16018) );
  OAI21_X1 U12150 ( .B1(n15902), .B2(n10090), .A(n10091), .ZN(n13927) );
  NAND2_X1 U12151 ( .A1(n10093), .A2(n13699), .ZN(n13789) );
  NAND2_X1 U12152 ( .A1(n15902), .A2(n13698), .ZN(n10093) );
  NAND2_X1 U12153 ( .A1(n10095), .A2(n13672), .ZN(n15912) );
  AND2_X1 U12154 ( .A1(n14526), .A2(n16003), .ZN(n14517) );
  OR2_X1 U12155 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20744) );
  INV_X1 U12156 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20419) );
  INV_X1 U12157 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20882) );
  NOR2_X1 U12158 ( .A1(n13116), .A2(n13219), .ZN(n15628) );
  CLKBUF_X1 U12159 ( .A(n13161), .Z(n14600) );
  INV_X1 U12160 ( .A(n14608), .ZN(n14614) );
  NAND2_X1 U12161 ( .A1(n9815), .A2(n20263), .ZN(n13163) );
  INV_X1 U12162 ( .A(n11967), .ZN(n9815) );
  INV_X1 U12163 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16074) );
  OR2_X1 U12164 ( .A1(n20390), .A2(n20681), .ZN(n20368) );
  OAI211_X1 U12165 ( .C1(n20509), .C2(n20506), .A(n20505), .B(n20504), .ZN(
        n20533) );
  OR2_X1 U12166 ( .A1(n20743), .A2(n20582), .ZN(n20645) );
  OAI22_X1 U12167 ( .A1(n20595), .A2(n20594), .B1(n20593), .B2(n20592), .ZN(
        n20625) );
  NAND2_X1 U12168 ( .A1(n20633), .A2(n20632), .ZN(n20730) );
  NAND2_X1 U12169 ( .A1(n20099), .A2(n20273), .ZN(n20739) );
  NAND2_X1 U12170 ( .A1(n20118), .A2(n20273), .ZN(n20762) );
  NAND2_X1 U12171 ( .A1(n20123), .A2(n20273), .ZN(n20769) );
  NAND2_X1 U12172 ( .A1(n20129), .A2(n20273), .ZN(n20776) );
  NAND2_X1 U12173 ( .A1(n20133), .A2(n20273), .ZN(n20783) );
  INV_X1 U12174 ( .A(n20626), .ZN(n20913) );
  OR2_X1 U12175 ( .A1(n15652), .A2(n20804), .ZN(n19871) );
  INV_X1 U12176 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n21068) );
  NAND2_X1 U12177 ( .A1(n10716), .A2(n10068), .ZN(n10725) );
  NAND2_X1 U12178 ( .A1(n9998), .A2(n15610), .ZN(n15609) );
  INV_X1 U12179 ( .A(n19064), .ZN(n19011) );
  OR2_X1 U12180 ( .A1(n11201), .A2(n11200), .ZN(n13346) );
  INV_X1 U12181 ( .A(n19095), .ZN(n19100) );
  AND2_X2 U12182 ( .A1(n13005), .A2(n16351), .ZN(n19103) );
  INV_X1 U12183 ( .A(n19111), .ZN(n15086) );
  NOR2_X1 U12184 ( .A1(n15056), .A2(n14794), .ZN(n14974) );
  AND2_X1 U12185 ( .A1(n13812), .A2(n13809), .ZN(n19110) );
  AND2_X1 U12186 ( .A1(n19169), .A2(n12972), .ZN(n19109) );
  AND2_X1 U12187 ( .A1(n12970), .A2(n16351), .ZN(n19169) );
  AND2_X1 U12188 ( .A1(n19169), .A2(n12986), .ZN(n19171) );
  INV_X1 U12189 ( .A(n19145), .ZN(n19175) );
  AND2_X1 U12190 ( .A1(n12871), .A2(n19737), .ZN(n19186) );
  AND2_X1 U12191 ( .A1(n13657), .A2(n19231), .ZN(n12840) );
  XNOR2_X1 U12192 ( .A(n11414), .B(n11312), .ZN(n14938) );
  INV_X1 U12193 ( .A(n9963), .ZN(n15377) );
  NAND2_X1 U12194 ( .A1(n15211), .A2(n15212), .ZN(n15594) );
  INV_X1 U12195 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10838) );
  INV_X1 U12196 ( .A(n16268), .ZN(n19229) );
  INV_X1 U12197 ( .A(n16278), .ZN(n19218) );
  INV_X1 U12198 ( .A(n10135), .ZN(n11425) );
  AOI211_X1 U12199 ( .C1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n15245), .A(
        n15244), .B(n15243), .ZN(n15250) );
  NAND2_X1 U12200 ( .A1(n15262), .A2(n10163), .ZN(n10749) );
  NAND2_X1 U12201 ( .A1(n15098), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15262) );
  NAND2_X1 U12202 ( .A1(n9872), .A2(n15297), .ZN(n9871) );
  NAND2_X1 U12203 ( .A1(n14630), .A2(n10033), .ZN(n15052) );
  XNOR2_X1 U12204 ( .A(n9856), .B(n9761), .ZN(n15339) );
  OAI21_X1 U12205 ( .B1(n15189), .B2(n9854), .A(n9775), .ZN(n9856) );
  INV_X1 U12206 ( .A(n15154), .ZN(n9854) );
  NAND2_X1 U12207 ( .A1(n15189), .A2(n15153), .ZN(n15164) );
  XNOR2_X1 U12208 ( .A(n9839), .B(n15177), .ZN(n15362) );
  NAND2_X1 U12209 ( .A1(n9840), .A2(n15187), .ZN(n9839) );
  NAND2_X1 U12210 ( .A1(n15189), .A2(n15186), .ZN(n9840) );
  NOR2_X1 U12211 ( .A1(n11047), .A2(n13899), .ZN(n15444) );
  INV_X1 U12212 ( .A(n16327), .ZN(n16316) );
  XNOR2_X1 U12213 ( .A(n15148), .B(n15397), .ZN(n16211) );
  AND2_X1 U12214 ( .A1(n10133), .A2(n9762), .ZN(n15232) );
  INV_X1 U12215 ( .A(n15211), .ZN(n15435) );
  NAND2_X1 U12216 ( .A1(n10133), .A2(n10642), .ZN(n15439) );
  NAND2_X1 U12217 ( .A1(n14192), .A2(n15598), .ZN(n16334) );
  INV_X1 U12218 ( .A(n19073), .ZN(n19850) );
  INV_X1 U12219 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19846) );
  INV_X1 U12220 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19837) );
  XNOR2_X1 U12221 ( .A(n13060), .B(n13018), .ZN(n19831) );
  INV_X1 U12222 ( .A(n19842), .ZN(n19832) );
  NOR2_X1 U12223 ( .A1(n13522), .A2(n11090), .ZN(n13517) );
  AOI22_X1 U12224 ( .A1(n13054), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19830), .B2(n19855), .ZN(n12975) );
  NAND2_X1 U12225 ( .A1(n19065), .A2(n13012), .ZN(n12976) );
  AND2_X1 U12226 ( .A1(n13467), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15467) );
  INV_X1 U12227 ( .A(n19269), .ZN(n19822) );
  INV_X1 U12228 ( .A(n10292), .ZN(n13474) );
  AOI21_X1 U12229 ( .B1(n13490), .B2(n16351), .A(n12922), .ZN(n15470) );
  INV_X1 U12230 ( .A(n19358), .ZN(n19350) );
  OAI21_X1 U12231 ( .B1(n13540), .B2(n19372), .A(n13539), .ZN(n19375) );
  NOR2_X1 U12232 ( .A1(n19435), .A2(n19597), .ZN(n19422) );
  INV_X1 U12233 ( .A(n19489), .ZN(n19491) );
  OAI21_X1 U12234 ( .B1(n19534), .B2(n19553), .A(n19679), .ZN(n19556) );
  NOR2_X1 U12235 ( .A1(n19626), .A2(n19329), .ZN(n19559) );
  INV_X1 U12236 ( .A(n19695), .ZN(n19539) );
  INV_X1 U12237 ( .A(n19701), .ZN(n19579) );
  INV_X1 U12238 ( .A(n19729), .ZN(n19643) );
  OR2_X1 U12239 ( .A1(n19592), .A2(n19597), .ZN(n19646) );
  INV_X1 U12240 ( .A(n19707), .ZN(n19647) );
  INV_X1 U12241 ( .A(n19713), .ZN(n19651) );
  INV_X1 U12242 ( .A(n19646), .ZN(n19661) );
  INV_X1 U12243 ( .A(n19607), .ZN(n19681) );
  INV_X1 U12244 ( .A(n19233), .ZN(n19687) );
  INV_X1 U12245 ( .A(n19542), .ZN(n19692) );
  INV_X1 U12246 ( .A(n19545), .ZN(n19698) );
  AND2_X1 U12247 ( .A1(n10265), .A2(n19256), .ZN(n19696) );
  AND2_X1 U12248 ( .A1(n19244), .A2(n19256), .ZN(n19702) );
  INV_X1 U12249 ( .A(n19654), .ZN(n19710) );
  AND2_X1 U12250 ( .A1(n13441), .A2(n19256), .ZN(n19708) );
  NOR2_X2 U12251 ( .A1(n19592), .A2(n19819), .ZN(n19725) );
  INV_X1 U12252 ( .A(n19666), .ZN(n19724) );
  AND2_X1 U12253 ( .A1(n19257), .A2(n19256), .ZN(n19720) );
  INV_X1 U12254 ( .A(n19036), .ZN(n19077) );
  AND2_X1 U12255 ( .A1(n11361), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16351) );
  NOR2_X1 U12256 ( .A1(n9681), .A2(n11676), .ZN(n16523) );
  INV_X1 U12257 ( .A(n17440), .ZN(n17378) );
  NOR2_X1 U12258 ( .A1(n16593), .A2(n17511), .ZN(n16592) );
  NOR2_X1 U12259 ( .A1(n16605), .A2(n16835), .ZN(n16593) );
  AND2_X1 U12260 ( .A1(n9884), .A2(n9898), .ZN(n16613) );
  NAND2_X1 U12261 ( .A1(n16628), .A2(n9898), .ZN(n9880) );
  NOR2_X1 U12262 ( .A1(n18682), .A2(n16543), .ZN(n16873) );
  NOR2_X1 U12263 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16663), .ZN(n16643) );
  AND2_X1 U12264 ( .A1(n9899), .A2(n9898), .ZN(n16645) );
  NAND2_X1 U12265 ( .A1(n9896), .A2(n9897), .ZN(n16644) );
  NOR2_X1 U12266 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16852), .ZN(n16841) );
  NOR2_X2 U12267 ( .A1(n18790), .A2(n16912), .ZN(n16902) );
  NOR2_X1 U12268 ( .A1(n16639), .A2(n16977), .ZN(n16982) );
  NOR2_X1 U12269 ( .A1(n17311), .A2(n17035), .ZN(n17022) );
  AND2_X1 U12270 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17063), .ZN(n17037) );
  NOR2_X1 U12271 ( .A1(n16723), .A2(n17089), .ZN(n17063) );
  NOR3_X1 U12272 ( .A1(n17106), .A2(n17211), .A3(n17102), .ZN(n17090) );
  INV_X1 U12273 ( .A(n17235), .ZN(n17231) );
  NOR2_X1 U12274 ( .A1(n17384), .A2(n17245), .ZN(n17241) );
  INV_X1 U12275 ( .A(n17259), .ZN(n17255) );
  NOR2_X1 U12276 ( .A1(n17311), .A2(n17264), .ZN(n17260) );
  NAND2_X1 U12277 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17306), .ZN(n17302) );
  NOR2_X1 U12278 ( .A1(n17489), .A2(n17314), .ZN(n17306) );
  NOR2_X1 U12279 ( .A1(n11466), .A2(n11465), .ZN(n17350) );
  NOR2_X1 U12280 ( .A1(n11476), .A2(n11475), .ZN(n17358) );
  NOR2_X1 U12281 ( .A1(n9994), .A2(n9991), .ZN(n9990) );
  INV_X1 U12282 ( .A(n17347), .ZN(n17363) );
  INV_X1 U12283 ( .A(n17345), .ZN(n17375) );
  INV_X1 U12284 ( .A(n17372), .ZN(n17361) );
  AND2_X1 U12285 ( .A1(n18645), .A2(n15717), .ZN(n17345) );
  INV_X1 U12286 ( .A(n17368), .ZN(n17370) );
  CLKBUF_X1 U12287 ( .A(n17485), .Z(n17476) );
  INV_X1 U12288 ( .A(n17488), .ZN(n17477) );
  OAI211_X1 U12289 ( .C1(n18834), .C2(n18192), .A(n9681), .B(n17440), .ZN(
        n17485) );
  NOR2_X1 U12290 ( .A1(n17476), .A2(n18192), .ZN(n17486) );
  AND2_X1 U12291 ( .A1(n17636), .A2(n9891), .ZN(n17562) );
  AND2_X1 U12292 ( .A1(n9708), .A2(n9892), .ZN(n9891) );
  INV_X1 U12293 ( .A(n17583), .ZN(n9892) );
  AND2_X1 U12294 ( .A1(n17794), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17775) );
  NOR2_X1 U12295 ( .A1(n17809), .A2(n17824), .ZN(n17806) );
  INV_X1 U12296 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17824) );
  INV_X1 U12297 ( .A(n18215), .ZN(n17816) );
  INV_X2 U12298 ( .A(n17816), .ZN(n18566) );
  NAND2_X1 U12299 ( .A1(n17600), .A2(n17696), .ZN(n17852) );
  INV_X1 U12300 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18800) );
  INV_X1 U12301 ( .A(n17850), .ZN(n17862) );
  INV_X1 U12302 ( .A(n11714), .ZN(n11741) );
  OAI21_X1 U12303 ( .B1(n17502), .B2(n11713), .A(n11712), .ZN(n11714) );
  OR2_X1 U12304 ( .A1(n15686), .A2(n9796), .ZN(n11713) );
  XNOR2_X1 U12305 ( .A(n17516), .B(n17767), .ZN(n17876) );
  NAND2_X1 U12306 ( .A1(n17515), .A2(n17514), .ZN(n17516) );
  NAND2_X1 U12307 ( .A1(n9935), .A2(n9934), .ZN(n17523) );
  INV_X1 U12308 ( .A(n9933), .ZN(n17522) );
  INV_X1 U12309 ( .A(n17897), .ZN(n18008) );
  OR2_X1 U12310 ( .A1(n17765), .A2(n9997), .ZN(n17717) );
  INV_X1 U12311 ( .A(n17923), .ZN(n18627) );
  AOI21_X2 U12312 ( .B1(n14083), .B2(n11711), .A(n18690), .ZN(n18158) );
  INV_X1 U12313 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18674) );
  INV_X2 U12314 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18820) );
  AOI211_X1 U12315 ( .C1(n18838), .C2(n18667), .A(n18187), .B(n14085), .ZN(
        n18821) );
  AND2_X1 U12316 ( .A1(n12762), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20102)
         );
  NAND2_X1 U12318 ( .A1(n14415), .A2(n12640), .ZN(n12750) );
  OAI22_X1 U12319 ( .A1(n12747), .A2(n20005), .B1(n14218), .B2(n20016), .ZN(
        n12748) );
  INV_X1 U12320 ( .A(n9999), .ZN(P2_U2824) );
  AOI21_X1 U12321 ( .B1(n14620), .B2(n9787), .A(n10000), .ZN(n9999) );
  OAI21_X1 U12322 ( .B1(n15278), .B2(n19221), .A(n11407), .ZN(n11408) );
  AOI21_X1 U12323 ( .B1(n16120), .B2(n19225), .A(n11406), .ZN(n11407) );
  OAI21_X1 U12324 ( .B1(n15290), .B2(n19219), .A(n9868), .ZN(P2_U2990) );
  INV_X1 U12325 ( .A(n9869), .ZN(n9868) );
  OAI21_X1 U12326 ( .B1(n15303), .B2(n19221), .A(n9870), .ZN(n9869) );
  AOI21_X1 U12327 ( .B1(n15295), .B2(n19225), .A(n15120), .ZN(n9870) );
  NAND2_X1 U12328 ( .A1(n9961), .A2(n9960), .ZN(n9959) );
  AOI21_X1 U12329 ( .B1(n19104), .B2(n16312), .A(n14141), .ZN(n14144) );
  OAI21_X1 U12330 ( .B1(n16163), .B2(n16327), .A(n10159), .ZN(n14141) );
  OAI21_X1 U12331 ( .B1(n11306), .B2(n16326), .A(n11305), .ZN(n10036) );
  NOR4_X1 U12332 ( .A1(n9876), .A2(n16567), .A3(n16566), .A4(n9875), .ZN(n9874) );
  INV_X1 U12333 ( .A(n16563), .ZN(n9878) );
  NAND2_X1 U12334 ( .A1(n13131), .A2(n11855), .ZN(n13116) );
  INV_X2 U12335 ( .A(n14470), .ZN(n9834) );
  NAND2_X1 U12336 ( .A1(n12249), .A2(n10074), .ZN(n14068) );
  NAND2_X1 U12337 ( .A1(n12400), .A2(n9765), .ZN(n9691) );
  NAND2_X1 U12338 ( .A1(n10076), .A2(n9797), .ZN(n14256) );
  NAND2_X1 U12339 ( .A1(n11967), .A2(n11926), .ZN(n13122) );
  AND3_X1 U12340 ( .A1(n11813), .A2(n11814), .A3(n11815), .ZN(n9692) );
  NAND2_X1 U12341 ( .A1(n14630), .A2(n10035), .ZN(n15066) );
  NOR2_X1 U12342 ( .A1(n14255), .A2(n9759), .ZN(n9693) );
  NAND2_X1 U12343 ( .A1(n12249), .A2(n12248), .ZN(n13961) );
  AND2_X1 U12344 ( .A1(n10143), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9694) );
  OR3_X1 U12345 ( .A1(n14309), .A2(n12737), .A3(n9984), .ZN(n9695) );
  AND3_X1 U12346 ( .A1(n11490), .A2(n11495), .A3(n9989), .ZN(n9697) );
  AND2_X1 U12347 ( .A1(n10003), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9698) );
  AND2_X1 U12348 ( .A1(n9733), .A2(n11561), .ZN(n9699) );
  NAND2_X1 U12349 ( .A1(n16279), .A2(n9786), .ZN(n13807) );
  AND2_X1 U12350 ( .A1(n9896), .A2(n9735), .ZN(n9700) );
  AND2_X1 U12351 ( .A1(n10384), .A2(n10362), .ZN(n9701) );
  AND2_X1 U12352 ( .A1(n10061), .A2(n9771), .ZN(n9702) );
  NAND2_X1 U12353 ( .A1(n14267), .A2(n14266), .ZN(n14255) );
  INV_X1 U12354 ( .A(n14255), .ZN(n10076) );
  NOR2_X1 U12355 ( .A1(n14974), .A2(n14973), .ZN(n9703) );
  NOR2_X1 U12356 ( .A1(n17645), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9704) );
  NOR2_X1 U12357 ( .A1(n16311), .A2(n10026), .ZN(n9705) );
  INV_X1 U12358 ( .A(n10079), .ZN(n13762) );
  AND2_X1 U12359 ( .A1(n11819), .A2(n11818), .ZN(n9706) );
  NAND2_X1 U12360 ( .A1(n10022), .A2(n9791), .ZN(n13518) );
  NAND2_X1 U12361 ( .A1(n14047), .A2(n10168), .ZN(n14704) );
  AND2_X1 U12362 ( .A1(n10011), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9707) );
  AND2_X1 U12363 ( .A1(n9893), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9708) );
  INV_X1 U12364 ( .A(n10639), .ZN(n10060) );
  AND2_X1 U12365 ( .A1(n11998), .A2(n12108), .ZN(n9709) );
  AND2_X1 U12366 ( .A1(n10066), .A2(n10730), .ZN(n9710) );
  AND2_X1 U12367 ( .A1(n10007), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9711) );
  INV_X2 U12368 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20804) );
  OR2_X1 U12369 ( .A1(n10083), .A2(n10082), .ZN(n9712) );
  INV_X2 U12370 ( .A(n15541), .ZN(n15558) );
  NOR3_X2 U12371 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18796), .A3(
        n18659), .ZN(n11525) );
  OR2_X1 U12372 ( .A1(n15675), .A2(n9973), .ZN(n9715) );
  NAND2_X1 U12373 ( .A1(n13246), .A2(n11877), .ZN(n11842) );
  INV_X4 U12374 ( .A(n16938), .ZN(n17160) );
  OR2_X1 U12375 ( .A1(n14072), .A2(n9980), .ZN(n9716) );
  NAND2_X1 U12376 ( .A1(n10403), .A2(n14749), .ZN(n9717) );
  NAND2_X1 U12377 ( .A1(n14505), .A2(n13928), .ZN(n13982) );
  NAND2_X1 U12378 ( .A1(n15211), .A2(n10153), .ZN(n15178) );
  NAND2_X1 U12379 ( .A1(n15211), .A2(n15370), .ZN(n15190) );
  AND2_X1 U12380 ( .A1(n10716), .A2(n10066), .ZN(n9718) );
  NAND2_X1 U12381 ( .A1(n13732), .A2(n10080), .ZN(n13886) );
  AND2_X1 U12382 ( .A1(n15130), .A2(n15129), .ZN(n9719) );
  INV_X1 U12383 ( .A(n10356), .ZN(n10380) );
  OR2_X1 U12384 ( .A1(n11401), .A2(n11402), .ZN(n9720) );
  AND2_X1 U12385 ( .A1(n12400), .A2(n10084), .ZN(n9721) );
  OR2_X1 U12386 ( .A1(n15037), .A2(n15024), .ZN(n9722) );
  NAND2_X1 U12387 ( .A1(n10662), .A2(n10061), .ZN(n10065) );
  AND2_X1 U12388 ( .A1(n15119), .A2(n10144), .ZN(n11410) );
  AND4_X1 U12389 ( .A1(n11812), .A2(n11811), .A3(n11810), .A4(n11809), .ZN(
        n9725) );
  NAND4_X1 U12390 ( .A1(n15156), .A2(n15218), .A3(n10704), .A4(n15154), .ZN(
        n9726) );
  AND2_X1 U12391 ( .A1(n12400), .A2(n10085), .ZN(n14312) );
  AOI21_X1 U12392 ( .B1(n10804), .B2(n10803), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10805) );
  INV_X1 U12393 ( .A(n14673), .ZN(n10363) );
  OAI21_X1 U12394 ( .B1(n15148), .B2(n9726), .A(n10715), .ZN(n15136) );
  NAND2_X1 U12395 ( .A1(n9954), .A2(n10811), .ZN(n16245) );
  AND2_X1 U12396 ( .A1(n10058), .A2(n10639), .ZN(n9727) );
  AND2_X1 U12397 ( .A1(n9934), .A2(n9932), .ZN(n9728) );
  INV_X1 U12398 ( .A(n9900), .ZN(n16554) );
  NOR2_X1 U12399 ( .A1(n17535), .A2(n9901), .ZN(n9900) );
  AND4_X1 U12400 ( .A1(n11482), .A2(n11481), .A3(n11480), .A4(n11479), .ZN(
        n9729) );
  NOR3_X1 U12401 ( .A1(n15037), .A2(n10031), .A3(n10027), .ZN(n11412) );
  AND3_X1 U12402 ( .A1(n11491), .A2(n11489), .A3(n11492), .ZN(n9730) );
  NAND2_X1 U12403 ( .A1(n13065), .A2(n13066), .ZN(n13191) );
  AND2_X1 U12404 ( .A1(n13225), .A2(n9943), .ZN(n9731) );
  AND2_X1 U12405 ( .A1(n15831), .A2(n14059), .ZN(n9732) );
  AND2_X1 U12406 ( .A1(n10347), .A2(n10351), .ZN(n19065) );
  INV_X1 U12407 ( .A(n9647), .ZN(n16328) );
  NOR2_X1 U12408 ( .A1(n9945), .A2(n13219), .ZN(n9944) );
  NAND2_X1 U12409 ( .A1(n13680), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9734) );
  AND2_X1 U12410 ( .A1(n9897), .A2(n9898), .ZN(n9735) );
  INV_X1 U12411 ( .A(n9823), .ZN(n9822) );
  NOR2_X1 U12412 ( .A1(n13234), .A2(n11963), .ZN(n9823) );
  INV_X1 U12413 ( .A(n11916), .ZN(n9810) );
  AND3_X1 U12414 ( .A1(n10385), .A2(n10382), .A3(n10383), .ZN(n9736) );
  NOR2_X1 U12415 ( .A1(n13705), .A2(n16022), .ZN(n9737) );
  NOR2_X1 U12416 ( .A1(n10722), .A2(n15307), .ZN(n9738) );
  INV_X1 U12417 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9940) );
  NOR2_X1 U12418 ( .A1(n13790), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9739) );
  INV_X1 U12419 ( .A(n10037), .ZN(n13192) );
  OAI21_X1 U12420 ( .B1(n10364), .B2(n13049), .A(n13055), .ZN(n10037) );
  AND4_X1 U12421 ( .A1(n10396), .A2(n10395), .A3(n10394), .A4(n10393), .ZN(
        n9740) );
  OR2_X1 U12422 ( .A1(n9822), .A2(n9821), .ZN(n9741) );
  INV_X1 U12423 ( .A(n15119), .ZN(n9872) );
  NAND2_X1 U12424 ( .A1(n13790), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9742) );
  OR2_X1 U12425 ( .A1(n17575), .A2(n16658), .ZN(n9743) );
  NAND2_X1 U12426 ( .A1(n12400), .A2(n12399), .ZN(n14318) );
  OR2_X1 U12427 ( .A1(n12984), .A2(n11082), .ZN(n9744) );
  AND2_X1 U12428 ( .A1(n11374), .A2(n11373), .ZN(n9745) );
  AND2_X1 U12429 ( .A1(n11904), .A2(n11841), .ZN(n9746) );
  AND2_X1 U12430 ( .A1(n9727), .A2(n10644), .ZN(n9747) );
  OR2_X1 U12431 ( .A1(n9834), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9748) );
  OR2_X1 U12432 ( .A1(n11409), .A2(n11408), .ZN(P2_U2988) );
  OR2_X1 U12433 ( .A1(n19257), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n9750) );
  INV_X1 U12434 ( .A(n13724), .ZN(n9946) );
  NAND2_X1 U12435 ( .A1(n13191), .A2(n10042), .ZN(n13282) );
  AND2_X1 U12436 ( .A1(n13282), .A2(n13281), .ZN(n9751) );
  NAND2_X1 U12437 ( .A1(n13552), .A2(n13551), .ZN(n13837) );
  AND2_X1 U12438 ( .A1(n13282), .A2(n9926), .ZN(n9752) );
  NOR2_X1 U12439 ( .A1(n15365), .A2(n14645), .ZN(n14630) );
  NOR2_X1 U12440 ( .A1(n14046), .A2(n10040), .ZN(n14983) );
  NOR2_X1 U12441 ( .A1(n17765), .A2(n9996), .ZN(n17698) );
  AND2_X1 U12442 ( .A1(n11351), .A2(n10003), .ZN(n9753) );
  AND2_X1 U12443 ( .A1(n11353), .A2(n9711), .ZN(n9754) );
  INV_X1 U12444 ( .A(n16872), .ZN(n16835) );
  AND2_X1 U12445 ( .A1(n10116), .A2(n13650), .ZN(n9755) );
  OR2_X1 U12446 ( .A1(n16835), .A2(n9888), .ZN(n9756) );
  AND2_X1 U12447 ( .A1(n14630), .A2(n14631), .ZN(n14629) );
  OR2_X1 U12448 ( .A1(n13415), .A2(n13512), .ZN(n13511) );
  AND2_X1 U12449 ( .A1(n16279), .A2(n10024), .ZN(n13806) );
  OR3_X1 U12450 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17576), .ZN(n9757) );
  NOR2_X1 U12451 ( .A1(n15236), .A2(n15235), .ZN(n13406) );
  AND2_X1 U12452 ( .A1(n10113), .A2(n10112), .ZN(n9758) );
  OAI211_X1 U12453 ( .C1(n10807), .C2(n10810), .A(n9860), .B(n9859), .ZN(
        n13895) );
  OR2_X1 U12454 ( .A1(n14339), .A2(n10075), .ZN(n9759) );
  NAND2_X1 U12455 ( .A1(n13591), .A2(n10789), .ZN(n13565) );
  OAI22_X1 U12456 ( .A1(n13011), .A2(n9922), .B1(n13010), .B2(n15453), .ZN(
        n13060) );
  NOR2_X1 U12457 ( .A1(n13392), .A2(n13393), .ZN(n13394) );
  AND2_X1 U12458 ( .A1(n10591), .A2(n10058), .ZN(n9760) );
  NAND2_X1 U12459 ( .A1(n17679), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17920) );
  AND2_X1 U12460 ( .A1(n15156), .A2(n15155), .ZN(n9761) );
  XNOR2_X1 U12461 ( .A(n14793), .B(n14792), .ZN(n15055) );
  AND2_X1 U12462 ( .A1(n10642), .A2(n10132), .ZN(n9762) );
  OR2_X1 U12463 ( .A1(n14470), .A2(n14563), .ZN(n9763) );
  OR3_X1 U12464 ( .A1(n14072), .A2(n9981), .A3(n12703), .ZN(n9764) );
  NAND2_X1 U12465 ( .A1(n14968), .A2(n14967), .ZN(n14966) );
  AND2_X1 U12466 ( .A1(n14313), .A2(n10085), .ZN(n9765) );
  OR2_X1 U12467 ( .A1(n14155), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9766) );
  NAND2_X1 U12468 ( .A1(n13732), .A2(n13763), .ZN(n10079) );
  OR2_X1 U12469 ( .A1(n9834), .A2(n14535), .ZN(n9767) );
  AND2_X1 U12470 ( .A1(n10127), .A2(n10660), .ZN(n9768) );
  AND2_X1 U12471 ( .A1(n9828), .A2(n14545), .ZN(n9769) );
  AND2_X1 U12472 ( .A1(n9880), .A2(n9883), .ZN(n9770) );
  NAND2_X1 U12473 ( .A1(n9649), .A2(n10669), .ZN(n9771) );
  AND2_X1 U12474 ( .A1(n13346), .A2(n13405), .ZN(n9772) );
  INV_X1 U12475 ( .A(n14326), .ZN(n12399) );
  NAND2_X1 U12476 ( .A1(n10074), .A2(n10073), .ZN(n9773) );
  OR2_X1 U12477 ( .A1(n10077), .A2(n9759), .ZN(n9774) );
  AND2_X1 U12478 ( .A1(n9852), .A2(n15165), .ZN(n9775) );
  NOR2_X1 U12479 ( .A1(n13933), .A2(n14497), .ZN(n9776) );
  AND2_X1 U12480 ( .A1(n9977), .A2(n13957), .ZN(n9777) );
  AND2_X1 U12481 ( .A1(n9926), .A2(n9772), .ZN(n9778) );
  AND2_X1 U12482 ( .A1(n11985), .A2(n11984), .ZN(n20269) );
  INV_X1 U12483 ( .A(n20269), .ZN(n9804) );
  NAND2_X1 U12484 ( .A1(n10779), .A2(n10780), .ZN(n9779) );
  AOI21_X1 U12485 ( .B1(n16605), .B2(n9889), .A(n9756), .ZN(n9885) );
  AND2_X1 U12486 ( .A1(n9705), .A2(n15441), .ZN(n9780) );
  AND2_X1 U12487 ( .A1(n9709), .A2(n12133), .ZN(n9781) );
  AND2_X1 U12488 ( .A1(n9755), .A2(n10115), .ZN(n9782) );
  AND4_X2 U12489 ( .A1(n10503), .A2(n10502), .A3(n10501), .A4(n10500), .ZN(
        n10640) );
  INV_X1 U12490 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9895) );
  NOR2_X1 U12491 ( .A1(n13997), .A2(n13958), .ZN(n9783) );
  NAND2_X1 U12492 ( .A1(n11107), .A2(n11106), .ZN(n13905) );
  AND2_X1 U12493 ( .A1(n13282), .A2(n9778), .ZN(n13552) );
  NAND2_X1 U12494 ( .A1(n13552), .A2(n10045), .ZN(n13860) );
  AND2_X1 U12495 ( .A1(n13737), .A2(n9977), .ZN(n9784) );
  AND2_X2 U12496 ( .A1(n11064), .A2(n11078), .ZN(n9785) );
  AND2_X1 U12497 ( .A1(n10024), .A2(n13808), .ZN(n9786) );
  INV_X1 U12498 ( .A(n14878), .ZN(n10049) );
  AND2_X1 U12499 ( .A1(n18910), .A2(n14619), .ZN(n9787) );
  NAND2_X1 U12500 ( .A1(n13191), .A2(n13190), .ZN(n13526) );
  XNOR2_X1 U12501 ( .A(n10294), .B(n19251), .ZN(n10976) );
  INV_X1 U12502 ( .A(n10717), .ZN(n10069) );
  AND2_X1 U12503 ( .A1(n12488), .A2(n12487), .ZN(n9788) );
  AND2_X1 U12504 ( .A1(n14816), .A2(n14815), .ZN(n9789) );
  AND2_X1 U12505 ( .A1(n9786), .A2(n10023), .ZN(n9790) );
  AND2_X1 U12506 ( .A1(n10018), .A2(n13516), .ZN(n9791) );
  NAND2_X1 U12507 ( .A1(n13991), .A2(n13954), .ZN(n9792) );
  OR2_X1 U12508 ( .A1(n17645), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9793) );
  NAND2_X1 U12509 ( .A1(n10103), .A2(n10104), .ZN(n10107) );
  AND2_X1 U12510 ( .A1(n10022), .A2(n10021), .ZN(n9794) );
  AND2_X1 U12511 ( .A1(n10033), .A2(n10032), .ZN(n9795) );
  OR2_X1 U12512 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n12152) );
  INV_X1 U12513 ( .A(n17767), .ZN(n17645) );
  INV_X1 U12514 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10008) );
  OR2_X1 U12515 ( .A1(n16356), .A2(n17341), .ZN(n9796) );
  AND2_X1 U12516 ( .A1(n12323), .A2(n12322), .ZN(n9797) );
  INV_X1 U12517 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10004) );
  INV_X1 U12518 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10005) );
  INV_X1 U12519 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10009) );
  INV_X1 U12520 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10012) );
  INV_X1 U12521 ( .A(n18698), .ZN(n16881) );
  AND2_X1 U12522 ( .A1(n17636), .A2(n9893), .ZN(n9798) );
  AND2_X1 U12523 ( .A1(n15682), .A2(n15674), .ZN(n9799) );
  AND2_X1 U12524 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n9800) );
  NOR2_X1 U12525 ( .A1(n14925), .A2(n10051), .ZN(n9801) );
  INV_X1 U12526 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n9931) );
  INV_X1 U12527 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n9956) );
  INV_X1 U12528 ( .A(n14561), .ZN(n9829) );
  INV_X1 U12529 ( .A(n15909), .ZN(n20101) );
  AOI22_X2 U12530 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n9636), .B1(DATAI_18_), 
        .B2(n9632), .ZN(n20767) );
  AOI22_X2 U12531 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n9636), .B1(DATAI_30_), 
        .B2(n9632), .ZN(n20722) );
  AOI22_X2 U12532 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n9636), .B1(DATAI_31_), 
        .B2(n9632), .ZN(n20910) );
  AOI22_X2 U12533 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n9636), .B1(DATAI_25_), 
        .B2(n9632), .ZN(n20697) );
  NOR3_X2 U12534 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18694), .A3(
        n18310), .ZN(n18238) );
  NOR3_X2 U12535 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18694), .A3(
        n18448), .ZN(n18419) );
  NOR3_X2 U12536 ( .A1(n18694), .A2(n18649), .A3(n18310), .ZN(n18281) );
  NOR3_X2 U12537 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18694), .A3(
        n18401), .ZN(n18375) );
  AOI22_X2 U12538 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n9636), .B1(DATAI_29_), 
        .B2(n9632), .ZN(n20717) );
  NOR3_X2 U12539 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18694), .A3(
        n18359), .ZN(n18327) );
  NOR2_X4 U12540 ( .A1(n20824), .A2(n20905), .ZN(n20864) );
  XNOR2_X1 U12541 ( .A(n9802), .B(n11960), .ZN(n12056) );
  NAND2_X1 U12542 ( .A1(n11902), .A2(n11901), .ZN(n9802) );
  NAND2_X2 U12543 ( .A1(n13111), .A2(n11877), .ZN(n11884) );
  AND2_X2 U12544 ( .A1(n12400), .A2(n9803), .ZN(n14234) );
  NOR2_X2 U12545 ( .A1(n13415), .A2(n9806), .ZN(n13609) );
  AND2_X2 U12546 ( .A1(n13609), .A2(n12172), .ZN(n13732) );
  NAND2_X1 U12547 ( .A1(n11899), .A2(n9808), .ZN(n9807) );
  OAI211_X2 U12548 ( .C1(n11899), .C2(n9810), .A(n9809), .B(n9807), .ZN(n20226) );
  NAND2_X1 U12549 ( .A1(n11946), .A2(n11924), .ZN(n11922) );
  NAND2_X2 U12550 ( .A1(n20226), .A2(n11943), .ZN(n11946) );
  NAND2_X1 U12551 ( .A1(n15913), .A2(n10094), .ZN(n9813) );
  NAND3_X1 U12552 ( .A1(n15913), .A2(n13670), .A3(n13669), .ZN(n9814) );
  XNOR2_X2 U12553 ( .A(n11967), .B(n20263), .ZN(n13145) );
  NAND2_X2 U12554 ( .A1(n10100), .A2(n13980), .ZN(n14146) );
  NAND2_X2 U12555 ( .A1(n9827), .A2(n9826), .ZN(n14505) );
  AND2_X2 U12556 ( .A1(n9746), .A2(n9706), .ZN(n13131) );
  MUX2_X1 U12557 ( .A(n13205), .B(n13206), .S(n13222), .Z(n13212) );
  OAI21_X1 U12558 ( .B1(n14453), .B2(n14534), .A(n9816), .ZN(n9818) );
  AND2_X2 U12559 ( .A1(n13220), .A2(n12008), .ZN(n12069) );
  NAND3_X1 U12560 ( .A1(n11967), .A2(n11926), .A3(n20804), .ZN(n9824) );
  NAND2_X1 U12561 ( .A1(n15902), .A2(n10091), .ZN(n9827) );
  INV_X1 U12562 ( .A(n14154), .ZN(n9831) );
  NAND2_X1 U12563 ( .A1(n14154), .A2(n14561), .ZN(n14156) );
  NAND2_X1 U12564 ( .A1(n14154), .A2(n9833), .ZN(n9832) );
  NAND2_X1 U12565 ( .A1(n11927), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11801) );
  NOR2_X1 U12566 ( .A1(n9838), .A2(n13116), .ZN(n12951) );
  NAND2_X1 U12567 ( .A1(n9637), .A2(n9781), .ZN(n13704) );
  OAI21_X2 U12568 ( .B1(n15201), .B2(n9855), .A(n15205), .ZN(n15189) );
  XNOR2_X2 U12569 ( .A(n10360), .B(n10347), .ZN(n14673) );
  XNOR2_X2 U12570 ( .A(n10355), .B(n10354), .ZN(n10356) );
  AND2_X2 U12571 ( .A1(n9841), .A2(n10223), .ZN(n10142) );
  NAND3_X1 U12572 ( .A1(n10260), .A2(n10258), .A3(n10259), .ZN(n9843) );
  NAND3_X1 U12573 ( .A1(n10254), .A2(n10253), .A3(n10256), .ZN(n9847) );
  NAND2_X1 U12574 ( .A1(n9849), .A2(n11027), .ZN(n9851) );
  NAND4_X1 U12575 ( .A1(n9736), .A2(n9850), .A3(n9662), .A4(n9701), .ZN(n9849)
         );
  OR2_X2 U12576 ( .A1(n10525), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13579) );
  OAI21_X2 U12577 ( .B1(n10514), .B2(n10962), .A(n13661), .ZN(n10525) );
  NAND2_X1 U12578 ( .A1(n10794), .A2(n13566), .ZN(n9857) );
  AND2_X1 U12579 ( .A1(n9958), .A2(n9857), .ZN(n13745) );
  NAND2_X2 U12580 ( .A1(n9858), .A2(n10348), .ZN(n10347) );
  NAND2_X1 U12581 ( .A1(n10807), .A2(n9861), .ZN(n9860) );
  INV_X1 U12582 ( .A(n10810), .ZN(n9863) );
  NAND3_X1 U12583 ( .A1(n10421), .A2(n9867), .A3(n9866), .ZN(n9865) );
  NAND2_X2 U12584 ( .A1(n10817), .A2(n10816), .ZN(n15211) );
  AND2_X2 U12585 ( .A1(n9918), .A2(n9779), .ZN(n10483) );
  OAI21_X1 U12586 ( .B1(n9877), .B2(n18698), .A(n9874), .ZN(P3_U2641) );
  XNOR2_X1 U12587 ( .A(n9879), .B(n9878), .ZN(n9877) );
  NOR2_X1 U12588 ( .A1(n16572), .A2(n16835), .ZN(n9879) );
  OR2_X1 U12589 ( .A1(n16628), .A2(n9882), .ZN(n9881) );
  INV_X1 U12590 ( .A(n9884), .ZN(n16627) );
  INV_X1 U12591 ( .A(n9899), .ZN(n16656) );
  INV_X1 U12592 ( .A(n16835), .ZN(n9898) );
  INV_X1 U12593 ( .A(n10420), .ZN(n9905) );
  NAND2_X1 U12594 ( .A1(n10420), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n9906) );
  NAND2_X1 U12595 ( .A1(n10420), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n9907) );
  NAND2_X1 U12596 ( .A1(n10420), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n9908) );
  INV_X1 U12597 ( .A(n10379), .ZN(n9910) );
  OR2_X2 U12598 ( .A1(n10798), .A2(n10962), .ZN(n9911) );
  OAI21_X2 U12599 ( .B1(n15148), .B2(n9915), .A(n9912), .ZN(n15115) );
  OAI21_X2 U12600 ( .B1(n15115), .B2(n15113), .A(n15111), .ZN(n11396) );
  NAND3_X1 U12601 ( .A1(n10484), .A2(n10483), .A3(n11095), .ZN(n10793) );
  NAND3_X1 U12602 ( .A1(n10480), .A2(n10422), .A3(n9919), .ZN(n9918) );
  NOR2_X2 U12603 ( .A1(n11384), .A2(n11423), .ZN(n9920) );
  AND2_X2 U12604 ( .A1(n10135), .A2(n9921), .ZN(n11384) );
  XNOR2_X1 U12605 ( .A(n13011), .B(n9922), .ZN(n19842) );
  NAND2_X1 U12606 ( .A1(n15056), .A2(n9925), .ZN(n9924) );
  NAND2_X1 U12607 ( .A1(n17836), .A2(n17837), .ZN(n17835) );
  NAND3_X1 U12608 ( .A1(n9728), .A2(n9935), .A3(n9931), .ZN(n9930) );
  NOR2_X2 U12609 ( .A1(n11556), .A2(n18088), .ZN(n18050) );
  NAND2_X1 U12610 ( .A1(n17856), .A2(n17848), .ZN(n17847) );
  XNOR2_X2 U12611 ( .A(n11726), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17848) );
  NAND4_X2 U12612 ( .A1(n9697), .A2(n9730), .A3(n9938), .A4(n11496), .ZN(
        n11726) );
  INV_X1 U12613 ( .A(n11493), .ZN(n9938) );
  AND2_X2 U12614 ( .A1(n9940), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11762) );
  XNOR2_X1 U12615 ( .A(n13228), .B(n13229), .ZN(n13267) );
  NAND2_X1 U12616 ( .A1(n9950), .A2(n9951), .ZN(n9949) );
  NAND2_X1 U12617 ( .A1(n11299), .A2(n9678), .ZN(n9950) );
  NAND2_X1 U12618 ( .A1(n9952), .A2(n10273), .ZN(n9951) );
  NAND2_X1 U12619 ( .A1(n11031), .A2(n10165), .ZN(n9952) );
  OAI21_X1 U12620 ( .B1(n9957), .B2(n13895), .A(n9953), .ZN(n10817) );
  NAND2_X1 U12621 ( .A1(n10795), .A2(n13750), .ZN(n9958) );
  NAND2_X1 U12622 ( .A1(n10799), .A2(n13747), .ZN(n10804) );
  AND2_X2 U12623 ( .A1(n13150), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11761) );
  NAND3_X1 U12624 ( .A1(n9966), .A2(n9748), .A3(n9969), .ZN(n13981) );
  NAND2_X1 U12625 ( .A1(n14052), .A2(n14053), .ZN(n9966) );
  INV_X1 U12626 ( .A(n13933), .ZN(n9967) );
  NOR2_X1 U12627 ( .A1(n14497), .A2(n9732), .ZN(n9968) );
  NAND3_X1 U12628 ( .A1(n11895), .A2(n11894), .A3(n13128), .ZN(n11896) );
  NAND2_X2 U12629 ( .A1(n12649), .A2(n9972), .ZN(n14168) );
  NAND2_X2 U12630 ( .A1(n13704), .A2(n13703), .ZN(n13705) );
  NAND2_X1 U12631 ( .A1(n9972), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n12651) );
  NAND2_X1 U12632 ( .A1(n9972), .A2(n13244), .ZN(n12655) );
  NAND2_X1 U12633 ( .A1(n9972), .A2(n16036), .ZN(n12671) );
  NAND2_X1 U12634 ( .A1(n9972), .A2(n16039), .ZN(n12676) );
  NAND2_X1 U12635 ( .A1(n9972), .A2(n14508), .ZN(n12682) );
  NAND2_X1 U12636 ( .A1(n9972), .A2(n13931), .ZN(n12687) );
  NAND2_X1 U12637 ( .A1(n9972), .A2(n14059), .ZN(n12694) );
  NAND2_X1 U12638 ( .A1(n9972), .A2(n15863), .ZN(n12699) );
  NAND2_X1 U12639 ( .A1(n9972), .A2(n15852), .ZN(n12705) );
  NAND2_X1 U12640 ( .A1(n9972), .A2(n14461), .ZN(n12721) );
  NAND2_X1 U12641 ( .A1(n9972), .A2(n14149), .ZN(n12727) );
  NAND2_X1 U12642 ( .A1(n9972), .A2(n14448), .ZN(n12732) );
  NAND2_X1 U12643 ( .A1(n12659), .A2(n9972), .ZN(n12661) );
  NAND2_X1 U12644 ( .A1(n12714), .A2(n9972), .ZN(n12716) );
  NAND3_X1 U12645 ( .A1(n12662), .A2(n12663), .A3(n9972), .ZN(n12664) );
  NAND3_X1 U12646 ( .A1(n12666), .A2(n12667), .A3(n9972), .ZN(n12668) );
  NAND3_X1 U12647 ( .A1(n12710), .A2(n12711), .A3(n9972), .ZN(n12712) );
  NAND3_X1 U12648 ( .A1(n9974), .A2(n14314), .A3(n14321), .ZN(n9973) );
  NAND3_X1 U12649 ( .A1(n11484), .A2(n11483), .A3(n9992), .ZN(n9991) );
  NAND2_X1 U12650 ( .A1(n11742), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17514) );
  INV_X2 U12651 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18814) );
  OAI211_X1 U12652 ( .C1(n9998), .C2(n15610), .A(n15609), .B(n19036), .ZN(
        n15611) );
  NAND2_X1 U12653 ( .A1(n18885), .A2(n11360), .ZN(n9998) );
  NAND2_X1 U12654 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11341) );
  NAND3_X1 U12655 ( .A1(n11375), .A2(n10001), .A3(n9745), .ZN(n10000) );
  AND2_X1 U12656 ( .A1(n9698), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10002) );
  AND2_X2 U12657 ( .A1(n11336), .A2(n10010), .ZN(n11327) );
  XNOR2_X1 U12658 ( .A(n12984), .B(n11082), .ZN(n12990) );
  OAI21_X1 U12659 ( .B1(n12990), .B2(n12989), .A(n9744), .ZN(n10013) );
  NAND4_X1 U12660 ( .A1(n10245), .A2(n10246), .A3(n10247), .A4(n10015), .ZN(
        n10014) );
  NAND4_X1 U12661 ( .A1(n10249), .A2(n10251), .A3(n10250), .A4(n10017), .ZN(
        n10016) );
  NAND3_X1 U12662 ( .A1(n10022), .A2(n10021), .A3(n13753), .ZN(n13752) );
  NAND2_X1 U12663 ( .A1(n13905), .A2(n9780), .ZN(n15440) );
  NAND3_X1 U12664 ( .A1(n10030), .A2(n10029), .A3(n11413), .ZN(n10028) );
  INV_X1 U12665 ( .A(n15009), .ZN(n10031) );
  NAND2_X1 U12666 ( .A1(n14630), .A2(n9795), .ZN(n15054) );
  XNOR2_X2 U12667 ( .A(n10829), .B(n10832), .ZN(n10364) );
  NAND2_X1 U12668 ( .A1(n14858), .A2(n10049), .ZN(n10046) );
  CLKBUF_X1 U12669 ( .A(n10398), .Z(n10050) );
  NAND4_X1 U12670 ( .A1(n9740), .A2(n10404), .A3(n10405), .A4(n10406), .ZN(
        n10057) );
  NAND2_X1 U12671 ( .A1(n9747), .A2(n10591), .ZN(n10646) );
  INV_X1 U12672 ( .A(n10065), .ZN(n10673) );
  NAND2_X1 U12673 ( .A1(n10716), .A2(n10717), .ZN(n10724) );
  NAND2_X1 U12674 ( .A1(n20424), .A2(n12073), .ZN(n10070) );
  XNOR2_X2 U12675 ( .A(n10096), .B(n12069), .ZN(n20424) );
  NAND2_X1 U12676 ( .A1(n10070), .A2(n10071), .ZN(n13085) );
  INV_X1 U12677 ( .A(n13085), .ZN(n12074) );
  NAND2_X1 U12678 ( .A1(n13241), .A2(n13240), .ZN(n10089) );
  XNOR2_X1 U12679 ( .A(n13350), .B(n10089), .ZN(n14122) );
  NAND2_X1 U12680 ( .A1(n13670), .A2(n13669), .ZN(n10095) );
  NOR2_X1 U12681 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10102) );
  NAND3_X1 U12682 ( .A1(n10103), .A2(n10104), .A3(n13302), .ZN(n13303) );
  INV_X1 U12683 ( .A(n10107), .ZN(n13311) );
  NAND2_X1 U12684 ( .A1(n13446), .A2(n9782), .ZN(n15223) );
  INV_X1 U12685 ( .A(n11028), .ZN(n10124) );
  NAND2_X1 U12686 ( .A1(n10126), .A2(n10125), .ZN(n11028) );
  AOI21_X1 U12687 ( .B1(n19244), .B2(n10269), .A(n12986), .ZN(n10125) );
  NAND2_X1 U12688 ( .A1(n10270), .A2(n10271), .ZN(n10126) );
  NAND2_X1 U12689 ( .A1(n13896), .A2(n10129), .ZN(n10128) );
  INV_X1 U12690 ( .A(n10166), .ZN(n10134) );
  NAND2_X1 U12691 ( .A1(n10954), .A2(n10166), .ZN(n10136) );
  INV_X1 U12692 ( .A(n15246), .ZN(n10139) );
  INV_X1 U12693 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10140) );
  AND2_X4 U12694 ( .A1(n10399), .A2(n10172), .ZN(n14929) );
  INV_X2 U12695 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10172) );
  NAND2_X1 U12696 ( .A1(n10335), .A2(n10141), .ZN(n10324) );
  NAND2_X1 U12697 ( .A1(n10320), .A2(n10141), .ZN(n10322) );
  XNOR2_X1 U12698 ( .A(n10335), .B(n10141), .ZN(n10353) );
  NAND2_X2 U12699 ( .A1(n10313), .A2(n10314), .ZN(n10141) );
  NAND2_X1 U12700 ( .A1(n10142), .A2(n10262), .ZN(n10774) );
  AND2_X2 U12701 ( .A1(n10142), .A2(n12971), .ZN(n10298) );
  NAND2_X1 U12702 ( .A1(n10143), .A2(n9800), .ZN(n15121) );
  NAND2_X1 U12703 ( .A1(n15119), .A2(n10146), .ZN(n11393) );
  AND2_X1 U12704 ( .A1(n15119), .A2(n10148), .ZN(n11394) );
  NAND2_X1 U12705 ( .A1(n15119), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15104) );
  NAND2_X1 U12706 ( .A1(n10339), .A2(n10338), .ZN(n10151) );
  NAND3_X1 U12707 ( .A1(n10327), .A2(n10326), .A3(n10325), .ZN(n10355) );
  NAND4_X1 U12708 ( .A1(n10327), .A2(n10326), .A3(n10325), .A4(n10150), .ZN(
        n10149) );
  NAND3_X1 U12709 ( .A1(n10485), .A2(n10791), .A3(n13590), .ZN(n13591) );
  NAND2_X1 U12710 ( .A1(n10514), .A2(n10154), .ZN(n16270) );
  INV_X1 U12711 ( .A(n13590), .ZN(n10154) );
  CLKBUF_X1 U12712 ( .A(n14024), .Z(n16179) );
  INV_X1 U12713 ( .A(n11340), .ZN(n11354) );
  XNOR2_X1 U12714 ( .A(n11322), .B(n11321), .ZN(n11377) );
  NAND2_X1 U12715 ( .A1(n11325), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11322) );
  NAND2_X1 U12716 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n11345), .ZN(
        n11344) );
  NOR2_X2 U12717 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11763) );
  NAND2_X1 U12718 ( .A1(n13145), .A2(n20804), .ZN(n11985) );
  NAND2_X1 U12719 ( .A1(n13075), .A2(n11879), .ZN(n13216) );
  CLKBUF_X1 U12720 ( .A(n13724), .Z(n20673) );
  NAND2_X1 U12721 ( .A1(n15141), .A2(n15140), .ZN(n15143) );
  INV_X1 U12722 ( .A(n14447), .ZN(n14449) );
  OR2_X1 U12724 ( .A1(n11306), .A2(n19221), .ZN(n10966) );
  NOR2_X1 U12725 ( .A1(n10951), .A2(n10950), .ZN(n10967) );
  INV_X2 U12726 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13462) );
  NAND2_X1 U12727 ( .A1(n13353), .A2(n20424), .ZN(n20229) );
  OR2_X1 U12728 ( .A1(n20424), .A2(n20269), .ZN(n20743) );
  NOR2_X2 U12729 ( .A1(n15121), .A2(n15307), .ZN(n15119) );
  AND2_X1 U12730 ( .A1(n10291), .A2(n10290), .ZN(n10306) );
  AOI22_X1 U12731 ( .A1(n14748), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10184), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10256) );
  NAND2_X1 U12732 ( .A1(n10186), .A2(n10185), .ZN(n10190) );
  NAND2_X1 U12733 ( .A1(n10188), .A2(n10187), .ZN(n10189) );
  NAND2_X1 U12734 ( .A1(n19169), .A2(n12985), .ZN(n19145) );
  NOR2_X2 U12735 ( .A1(n11043), .A2(n10265), .ZN(n11034) );
  INV_X1 U12736 ( .A(n14325), .ZN(n12400) );
  NAND2_X1 U12737 ( .A1(n10634), .A2(n10633), .ZN(n13896) );
  AND2_X4 U12738 ( .A1(n13454), .A2(n10172), .ZN(n10257) );
  INV_X1 U12739 ( .A(n9690), .ZN(n19041) );
  NAND2_X1 U12740 ( .A1(n9657), .A2(n20136), .ZN(n12636) );
  NAND2_X1 U12741 ( .A1(n10799), .A2(n10798), .ZN(n10800) );
  INV_X1 U12742 ( .A(n10798), .ZN(n10803) );
  CLKBUF_X1 U12743 ( .A(n12908), .Z(n12952) );
  NAND2_X1 U12744 ( .A1(n12908), .A2(n20114), .ZN(n11879) );
  NOR2_X1 U12745 ( .A1(n16905), .A2(n11439), .ZN(n11530) );
  INV_X1 U12746 ( .A(n14816), .ZN(n14792) );
  INV_X1 U12747 ( .A(n10836), .ZN(n10329) );
  NAND2_X1 U12748 ( .A1(n9658), .A2(n14749), .ZN(n10158) );
  NAND2_X2 U12749 ( .A1(n14402), .A2(n13081), .ZN(n14370) );
  AND2_X2 U12750 ( .A1(n11762), .A2(n11764), .ZN(n12016) );
  NOR2_X1 U12751 ( .A1(n14140), .A2(n14139), .ZN(n10159) );
  OR2_X1 U12752 ( .A1(n11018), .A2(n16339), .ZN(n10160) );
  NAND2_X1 U12753 ( .A1(n14979), .A2(n14969), .ZN(n11401) );
  NOR2_X1 U12754 ( .A1(n20746), .A2(n20745), .ZN(n10162) );
  NAND2_X1 U12755 ( .A1(n10037), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10164) );
  AND3_X1 U12756 ( .A1(n10269), .A2(n9659), .A3(n19231), .ZN(n10165) );
  NAND2_X1 U12757 ( .A1(n20808), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20863) );
  AND2_X1 U12758 ( .A1(n15102), .A2(n11398), .ZN(n10166) );
  AND2_X1 U12759 ( .A1(n14856), .A2(n14876), .ZN(n10167) );
  NAND3_X1 U12760 ( .A1(n14045), .A2(n14044), .A3(n14043), .ZN(n10168) );
  INV_X1 U12761 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19829) );
  AND2_X1 U12762 ( .A1(n15101), .A2(n10740), .ZN(n10169) );
  INV_X1 U12763 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12305) );
  INV_X1 U12764 ( .A(n13059), .ZN(n13017) );
  INV_X1 U12765 ( .A(n13610), .ZN(n13734) );
  INV_X2 U12766 ( .A(n20028), .ZN(n20038) );
  NOR2_X1 U12767 ( .A1(n19079), .A2(n19078), .ZN(n10170) );
  OR2_X1 U12768 ( .A1(n11743), .A2(n18166), .ZN(n10171) );
  INV_X1 U12769 ( .A(n18050), .ZN(n17766) );
  NAND2_X1 U12770 ( .A1(n19103), .A2(n19257), .ZN(n19095) );
  AND2_X1 U12771 ( .A1(n16278), .A2(n19838), .ZN(n19225) );
  INV_X1 U12772 ( .A(n19225), .ZN(n16273) );
  INV_X1 U12773 ( .A(n14350), .ZN(n12640) );
  NAND2_X1 U12774 ( .A1(n20746), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12581) );
  NAND2_X1 U12775 ( .A1(n11896), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11897) );
  INV_X1 U12776 ( .A(n12609), .ZN(n12583) );
  OR2_X1 U12777 ( .A1(n12121), .A2(n12120), .ZN(n13692) );
  NAND2_X1 U12778 ( .A1(n11885), .A2(n11884), .ZN(n13113) );
  NAND2_X1 U12779 ( .A1(n12584), .A2(n12583), .ZN(n12611) );
  NAND2_X1 U12780 ( .A1(n11919), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11902) );
  OR2_X1 U12781 ( .A1(n11940), .A2(n11939), .ZN(n11941) );
  INV_X1 U12782 ( .A(n19244), .ZN(n10271) );
  INV_X1 U12783 ( .A(n14657), .ZN(n10357) );
  AOI21_X1 U12784 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20882), .A(
        n12589), .ZN(n12622) );
  INV_X1 U12785 ( .A(n11757), .ZN(n11765) );
  NOR2_X1 U12786 ( .A1(n11877), .A2(n11878), .ZN(n12956) );
  AND2_X1 U12787 ( .A1(n11997), .A2(n11996), .ZN(n11999) );
  OR2_X1 U12788 ( .A1(n11995), .A2(n11994), .ZN(n13674) );
  AND4_X1 U12789 ( .A1(n11755), .A2(n11754), .A3(n11753), .A4(n11752), .ZN(
        n11774) );
  NAND2_X1 U12790 ( .A1(n11878), .A2(n20104), .ZN(n11973) );
  INV_X1 U12791 ( .A(n10635), .ZN(n10636) );
  INV_X1 U12792 ( .A(n14838), .ZN(n14840) );
  AND4_X1 U12793 ( .A1(n10499), .A2(n10498), .A3(n10497), .A4(n10496), .ZN(
        n10500) );
  INV_X1 U12794 ( .A(n10323), .ZN(n10338) );
  AND2_X1 U12795 ( .A1(n10752), .A2(n10751), .ZN(n10999) );
  OAI21_X1 U12796 ( .B1(n11002), .B2(n10983), .A(n11001), .ZN(n11004) );
  NAND2_X1 U12797 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12623), .ZN(
        n12905) );
  OR2_X1 U12798 ( .A1(n13624), .A2(n14413), .ZN(n13625) );
  OR2_X1 U12799 ( .A1(n20172), .A2(n20383), .ZN(n12078) );
  INV_X1 U12800 ( .A(n14158), .ZN(n12300) );
  OR2_X1 U12801 ( .A1(n12040), .A2(n12039), .ZN(n13232) );
  INV_X1 U12802 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20383) );
  INV_X1 U12803 ( .A(n12008), .ZN(n12009) );
  AND2_X1 U12804 ( .A1(n14857), .A2(n10167), .ZN(n14858) );
  NAND2_X1 U12805 ( .A1(n10969), .A2(n10285), .ZN(n10836) );
  AND2_X1 U12806 ( .A1(n11285), .A2(n11284), .ZN(n15044) );
  AND2_X1 U12807 ( .A1(n10860), .A2(n10859), .ZN(n15235) );
  AOI21_X1 U12808 ( .B1(n11313), .B2(P2_REIP_REG_2__SCAN_IN), .A(n10332), .ZN(
        n10333) );
  INV_X1 U12809 ( .A(n13434), .ZN(n11041) );
  AND2_X1 U12810 ( .A1(n10363), .A2(n16328), .ZN(n10374) );
  AND2_X1 U12811 ( .A1(n14657), .A2(n10377), .ZN(n10366) );
  INV_X1 U12812 ( .A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n21092) );
  INV_X1 U12813 ( .A(n11647), .ZN(n11706) );
  NOR2_X1 U12814 ( .A1(n11447), .A2(n18665), .ZN(n11497) );
  NOR2_X1 U12815 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18820), .ZN(
        n11687) );
  NOR2_X1 U12816 ( .A1(n12079), .A2(n14115), .ZN(n12080) );
  NAND2_X1 U12817 ( .A1(n14126), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12549) );
  AND2_X1 U12818 ( .A1(n12531), .A2(n12510), .ZN(n14438) );
  NOR2_X1 U12819 ( .A1(n12374), .A2(n15774), .ZN(n12375) );
  AND2_X1 U12820 ( .A1(n12001), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12085) );
  AND2_X1 U12821 ( .A1(n12684), .A2(n12683), .ZN(n13764) );
  AND2_X1 U12822 ( .A1(n20114), .A2(n11877), .ZN(n13690) );
  AND4_X1 U12823 ( .A1(n11867), .A2(n11866), .A3(n11865), .A4(n11864), .ZN(
        n11873) );
  AND2_X1 U12824 ( .A1(n20230), .A2(n20741), .ZN(n20232) );
  NAND2_X1 U12825 ( .A1(n11972), .A2(n11971), .ZN(n20263) );
  NAND2_X1 U12826 ( .A1(n9656), .A2(n12077), .ZN(n13353) );
  AND3_X1 U12827 ( .A1(n20804), .A2(n20103), .A3(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20173) );
  AND2_X1 U12828 ( .A1(n10655), .A2(n10654), .ZN(n18966) );
  AND2_X1 U12829 ( .A1(n10897), .A2(n10896), .ZN(n14986) );
  OR2_X1 U12830 ( .A1(n13280), .A2(n19239), .ZN(n13059) );
  AND2_X1 U12831 ( .A1(n11269), .A2(n11268), .ZN(n15589) );
  AND2_X1 U12832 ( .A1(n11281), .A2(n11280), .ZN(n15067) );
  INV_X1 U12833 ( .A(n13406), .ZN(n15238) );
  AND2_X1 U12834 ( .A1(n19009), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16247) );
  NAND2_X1 U12835 ( .A1(n10334), .A2(n10333), .ZN(n10354) );
  INV_X1 U12836 ( .A(n19440), .ZN(n19378) );
  INV_X2 U12838 ( .A(n9713), .ZN(n17017) );
  NOR2_X1 U12839 ( .A1(n18702), .A2(n17845), .ZN(n16366) );
  AOI21_X1 U12840 ( .B1(n16398), .B2(n18031), .A(n15584), .ZN(n11712) );
  NOR2_X1 U12841 ( .A1(n17358), .A2(n11522), .ZN(n11544) );
  NOR2_X1 U12842 ( .A1(n11649), .A2(n11642), .ZN(n11678) );
  OR2_X1 U12843 ( .A1(n12634), .A2(n12633), .ZN(n13209) );
  INV_X1 U12844 ( .A(n20104), .ZN(n13619) );
  NAND2_X1 U12845 ( .A1(n12156), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12173) );
  AND2_X1 U12846 ( .A1(n14163), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13626) );
  NAND2_X1 U12847 ( .A1(n13638), .A2(n13628), .ZN(n19987) );
  OR2_X1 U12848 ( .A1(n13078), .A2(n14167), .ZN(n12638) );
  NAND2_X1 U12850 ( .A1(n12507), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12531) );
  NAND2_X1 U12851 ( .A1(n12375), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12426) );
  NOR2_X1 U12852 ( .A1(n12306), .A2(n12305), .ZN(n12339) );
  INV_X1 U12853 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n20934) );
  INV_X1 U12854 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15805) );
  INV_X1 U12855 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14115) );
  AND2_X1 U12856 ( .A1(n13114), .A2(n12961), .ZN(n15642) );
  OR2_X1 U12857 ( .A1(n14470), .A2(n13977), .ZN(n15875) );
  NOR2_X1 U12858 ( .A1(n15668), .A2(n15669), .ZN(n16003) );
  NAND2_X1 U12859 ( .A1(n13243), .A2(n13242), .ZN(n14526) );
  NOR2_X1 U12860 ( .A1(n20589), .A2(n15656), .ZN(n14608) );
  AND2_X1 U12861 ( .A1(n20145), .A2(n20144), .ZN(n20176) );
  AND2_X1 U12862 ( .A1(n20267), .A2(n20266), .ZN(n20297) );
  OR2_X1 U12863 ( .A1(n20390), .A2(n20631), .ZN(n20374) );
  AND2_X1 U12864 ( .A1(n20422), .A2(n20421), .ZN(n20451) );
  AND2_X1 U12865 ( .A1(n20542), .A2(n20541), .ZN(n20574) );
  AOI21_X1 U12866 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20635), .A(n20175), 
        .ZN(n20748) );
  INV_X1 U12867 ( .A(n13465), .ZN(n11368) );
  AND2_X1 U12868 ( .A1(n10772), .A2(n10771), .ZN(n11002) );
  INV_X1 U12869 ( .A(n19057), .ZN(n19043) );
  NAND4_X1 U12870 ( .A1(n19046), .A2(n18861), .A3(n19077), .A4(n16352), .ZN(
        n19068) );
  AND2_X1 U12871 ( .A1(n10906), .A2(n10905), .ZN(n15123) );
  NAND2_X1 U12872 ( .A1(n10215), .A2(n9846), .ZN(n10222) );
  NOR2_X1 U12873 ( .A1(n14943), .A2(n14942), .ZN(n14941) );
  NOR2_X1 U12874 ( .A1(n14957), .A2(n14956), .ZN(n14955) );
  AND3_X1 U12875 ( .A1(n11098), .A2(n11097), .A3(n11096), .ZN(n13524) );
  OR2_X1 U12876 ( .A1(n18914), .A2(n10640), .ZN(n10677) );
  OR3_X1 U12877 ( .A1(n14636), .A2(n10640), .A3(n15344), .ZN(n15165) );
  OR2_X1 U12878 ( .A1(n18948), .A2(n10712), .ZN(n15395) );
  NAND2_X1 U12879 ( .A1(n15467), .A2(n16342), .ZN(n13426) );
  INV_X1 U12880 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19593) );
  NAND2_X1 U12881 ( .A1(n19831), .A2(n19842), .ZN(n19329) );
  INV_X1 U12882 ( .A(n19230), .ZN(n19256) );
  NOR2_X1 U12883 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16679), .ZN(n16667) );
  NOR2_X1 U12884 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16708), .ZN(n16688) );
  NOR2_X1 U12885 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16807), .ZN(n16788) );
  INV_X1 U12886 ( .A(n16917), .ZN(n16823) );
  NAND2_X1 U12887 ( .A1(n18854), .A2(n16540), .ZN(n16543) );
  INV_X1 U12888 ( .A(n16873), .ZN(n16904) );
  INV_X1 U12889 ( .A(n18188), .ZN(n16540) );
  INV_X1 U12890 ( .A(n18208), .ZN(n17229) );
  AND4_X1 U12891 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16774), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17690) );
  INV_X1 U12892 ( .A(n16366), .ZN(n17600) );
  NOR2_X1 U12893 ( .A1(n11680), .A2(n11679), .ZN(n14083) );
  INV_X1 U12894 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18649) );
  NAND2_X1 U12895 ( .A1(n11700), .A2(n11703), .ZN(n18620) );
  NOR2_X1 U12896 ( .A1(n13718), .A2(n13619), .ZN(n13638) );
  AND2_X1 U12897 ( .A1(n19976), .A2(n13629), .ZN(n19946) );
  AND2_X1 U12898 ( .A1(n19976), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19978) );
  NAND2_X1 U12899 ( .A1(n13638), .A2(n13621), .ZN(n19965) );
  AND2_X1 U12900 ( .A1(n19976), .A2(n13626), .ZN(n19916) );
  AND2_X1 U12901 ( .A1(n19976), .A2(n13632), .ZN(n19979) );
  INV_X1 U12902 ( .A(n19976), .ZN(n19960) );
  INV_X1 U12903 ( .A(n20016), .ZN(n14310) );
  AND2_X1 U12904 ( .A1(n13268), .A2(n13038), .ZN(n20026) );
  NAND2_X1 U12905 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n12465), .ZN(
        n12505) );
  NAND2_X1 U12906 ( .A1(n12427), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12464) );
  NAND2_X1 U12907 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n12191), .ZN(
        n12229) );
  AND2_X1 U12908 ( .A1(n12137), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12156) );
  AND2_X1 U12909 ( .A1(n15918), .A2(n20075), .ZN(n15889) );
  NAND2_X1 U12910 ( .A1(n16071), .A2(n20804), .ZN(n13270) );
  NOR2_X1 U12911 ( .A1(n16003), .A2(n13336), .ZN(n16005) );
  INV_X1 U12912 ( .A(n14526), .ZN(n15999) );
  NOR2_X2 U12913 ( .A1(n13260), .A2(n13218), .ZN(n20087) );
  NAND2_X1 U12914 ( .A1(n20804), .A2(n20103), .ZN(n20175) );
  NOR2_X1 U12915 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n16071) );
  INV_X1 U12916 ( .A(n20911), .ZN(n20181) );
  INV_X1 U12917 ( .A(n20340), .ZN(n20300) );
  OAI21_X1 U12918 ( .B1(n20275), .B2(n20274), .A(n20686), .ZN(n20301) );
  OR2_X1 U12919 ( .A1(n20424), .A2(n9804), .ZN(n20390) );
  INV_X1 U12920 ( .A(n20374), .ZN(n20370) );
  INV_X1 U12921 ( .A(n20368), .ZN(n20415) );
  OAI211_X1 U12922 ( .C1(n20430), .C2(n20589), .A(n20504), .B(n20429), .ZN(
        n20454) );
  INV_X1 U12923 ( .A(n20536), .ZN(n20499) );
  INV_X1 U12924 ( .A(n20480), .ZN(n20493) );
  OAI22_X1 U12925 ( .A1(n20509), .A2(n20508), .B1(n20507), .B2(n20675), .ZN(
        n20532) );
  INV_X1 U12926 ( .A(n20581), .ZN(n20565) );
  INV_X1 U12927 ( .A(n20776), .ZN(n20612) );
  INV_X1 U12928 ( .A(n20790), .ZN(n20620) );
  INV_X1 U12929 ( .A(n20645), .ZN(n20669) );
  OAI211_X1 U12930 ( .C1(n20688), .C2(n20687), .A(n20686), .B(n20685), .ZN(
        n20727) );
  INV_X1 U12931 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20808) );
  INV_X1 U12932 ( .A(n20866), .ZN(n20859) );
  AND2_X1 U12933 ( .A1(n13660), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n19057) );
  INV_X1 U12934 ( .A(n19068), .ZN(n19045) );
  INV_X1 U12935 ( .A(n11317), .ZN(n11318) );
  AND3_X1 U12936 ( .A1(n11263), .A2(n11262), .A3(n11261), .ZN(n19078) );
  OR2_X1 U12937 ( .A1(n13065), .A2(n13066), .ZN(n13067) );
  AND2_X1 U12938 ( .A1(n13812), .A2(n13811), .ZN(n19111) );
  INV_X1 U12939 ( .A(n19169), .ZN(n19170) );
  OR2_X1 U12940 ( .A1(n19109), .A2(n13812), .ZN(n19161) );
  INV_X1 U12941 ( .A(n12793), .ZN(n12898) );
  INV_X1 U12942 ( .A(n19221), .ZN(n11389) );
  AND2_X1 U12943 ( .A1(n10819), .A2(n19231), .ZN(n16269) );
  AOI211_X1 U12944 ( .C1(n11384), .C2(n11383), .A(n11382), .B(n11423), .ZN(
        n11388) );
  INV_X1 U12945 ( .A(n16326), .ZN(n16317) );
  NAND2_X1 U12946 ( .A1(n11016), .A2(n16351), .ZN(n11304) );
  INV_X1 U12947 ( .A(n13498), .ZN(n13490) );
  OAI21_X1 U12948 ( .B1(n13786), .B2(n13785), .A(n13784), .ZN(n19262) );
  AND2_X1 U12949 ( .A1(n19271), .A2(n19268), .ZN(n19290) );
  NOR2_X1 U12950 ( .A1(n19497), .A2(n19435), .ZN(n19324) );
  NOR2_X1 U12951 ( .A1(n19435), .A2(n19329), .ZN(n19374) );
  NOR2_X1 U12952 ( .A1(n19407), .A2(n19597), .ZN(n19395) );
  OR3_X1 U12953 ( .A1(n19413), .A2(n19442), .A3(n19412), .ZN(n19431) );
  NAND2_X1 U12954 ( .A1(n19474), .A2(n19473), .ZN(n19492) );
  INV_X1 U12955 ( .A(n19515), .ZN(n19520) );
  AND2_X1 U12956 ( .A1(n13432), .A2(n13431), .ZN(n19571) );
  INV_X1 U12957 ( .A(n19684), .ZN(n19604) );
  OAI21_X1 U12958 ( .B1(n19636), .B2(n19635), .A(n19634), .ZN(n19662) );
  INV_X1 U12959 ( .A(n19658), .ZN(n19716) );
  NOR2_X2 U12960 ( .A1(n13811), .A2(n13429), .ZN(n19260) );
  INV_X1 U12961 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19752) );
  INV_X1 U12962 ( .A(n18635), .ZN(n18662) );
  OR2_X1 U12963 ( .A1(n16584), .A2(P3_EBX_REG_29__SCAN_IN), .ZN(n16562) );
  NOR2_X1 U12964 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16638), .ZN(n16626) );
  INV_X1 U12965 ( .A(n16883), .ZN(n16913) );
  NOR2_X1 U12966 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16730), .ZN(n16712) );
  NOR2_X1 U12967 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16755), .ZN(n16735) );
  NOR2_X1 U12968 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16777), .ZN(n16761) );
  NOR2_X1 U12969 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16829), .ZN(n16811) );
  INV_X1 U12970 ( .A(n16914), .ZN(n16875) );
  NOR2_X1 U12971 ( .A1(n16661), .A2(n17009), .ZN(n16983) );
  NAND2_X1 U12972 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17049), .ZN(n17035) );
  INV_X1 U12973 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16853) );
  NAND3_X1 U12974 ( .A1(n15712), .A2(n18840), .A3(n16540), .ZN(n17211) );
  NAND2_X1 U12975 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17255), .ZN(n17254) );
  AND2_X1 U12976 ( .A1(n17270), .A2(n17296), .ZN(n17290) );
  NOR2_X1 U12977 ( .A1(n17311), .A2(n17302), .ZN(n17296) );
  INV_X2 U12978 ( .A(n18219), .ZN(n17311) );
  INV_X1 U12979 ( .A(n17696), .ZN(n17706) );
  INV_X1 U12980 ( .A(n18049), .ZN(n17728) );
  AOI21_X1 U12981 ( .B1(n17936), .B2(n17507), .A(n17496), .ZN(n11744) );
  AND2_X1 U12982 ( .A1(n17931), .A2(n18158), .ZN(n17936) );
  NAND2_X1 U12983 ( .A1(n18662), .A2(n18143), .ZN(n17990) );
  NOR2_X1 U12984 ( .A1(n18040), .A2(n18173), .ZN(n18074) );
  INV_X1 U12985 ( .A(n18646), .ZN(n18633) );
  NAND2_X1 U12986 ( .A1(n18843), .A2(n18186), .ZN(n18288) );
  NOR2_X1 U12987 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18790), .ZN(
        n18815) );
  INV_X1 U12988 ( .A(n18418), .ZN(n18420) );
  INV_X1 U12989 ( .A(n18608), .ZN(n18550) );
  INV_X1 U12990 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18851) );
  INV_X1 U12991 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18710) );
  INV_X1 U12992 ( .A(n13809), .ZN(n13811) );
  NOR2_X1 U12993 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12774), .ZN(n16499)
         );
  INV_X1 U12994 ( .A(U212), .ZN(n16475) );
  INV_X1 U12995 ( .A(n13032), .ZN(n12948) );
  NAND2_X1 U12996 ( .A1(n12948), .A2(n12947), .ZN(n20894) );
  NAND2_X1 U12997 ( .A1(n13638), .A2(n13637), .ZN(n19985) );
  INV_X1 U12998 ( .A(n19978), .ZN(n19898) );
  AND2_X1 U12999 ( .A1(n19923), .A2(n13720), .ZN(n19937) );
  NAND2_X1 U13000 ( .A1(n20016), .A2(n14208), .ZN(n20005) );
  OR2_X1 U13001 ( .A1(n13992), .A2(n13956), .ZN(n15886) );
  NAND2_X1 U13002 ( .A1(n20041), .A2(n20019), .ZN(n20028) );
  INV_X1 U13003 ( .A(n20026), .ZN(n20041) );
  AND2_X1 U13004 ( .A1(n13032), .A2(n13030), .ZN(n13182) );
  INV_X1 U13005 ( .A(n15889), .ZN(n15914) );
  OR2_X1 U13006 ( .A1(n13270), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15996) );
  INV_X1 U13007 ( .A(n20087), .ZN(n16008) );
  INV_X1 U13008 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20635) );
  AND2_X1 U13009 ( .A1(n20098), .A2(n20097), .ZN(n20914) );
  OR2_X1 U13010 ( .A1(n20229), .A2(n20582), .ZN(n20911) );
  OR2_X1 U13011 ( .A1(n20229), .A2(n20631), .ZN(n20221) );
  OR2_X1 U13012 ( .A1(n20229), .A2(n20681), .ZN(n20257) );
  OR2_X1 U13013 ( .A1(n20229), .A2(n20551), .ZN(n20304) );
  OR2_X1 U13014 ( .A1(n20390), .A2(n20582), .ZN(n20340) );
  NAND2_X1 U13015 ( .A1(n20113), .A2(n20273), .ZN(n20755) );
  NAND2_X1 U13016 ( .A1(n20138), .A2(n20273), .ZN(n20790) );
  NAND2_X1 U13017 ( .A1(n20381), .A2(n20380), .ZN(n20457) );
  OR2_X1 U13018 ( .A1(n20552), .A2(n20582), .ZN(n20480) );
  OR2_X1 U13019 ( .A1(n20552), .A2(n20631), .ZN(n20536) );
  OR2_X1 U13020 ( .A1(n20552), .A2(n20681), .ZN(n20581) );
  OR2_X1 U13021 ( .A1(n20552), .A2(n20551), .ZN(n20630) );
  OR2_X1 U13022 ( .A1(n20743), .A2(n20551), .ZN(n20909) );
  INV_X1 U13023 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20589) );
  INV_X1 U13024 ( .A(n20807), .ZN(n20874) );
  INV_X1 U13025 ( .A(n20863), .ZN(n20904) );
  OR2_X1 U13026 ( .A1(n20905), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20866) );
  OR2_X1 U13027 ( .A1(n12916), .A2(n12868), .ZN(n18861) );
  NAND2_X1 U13028 ( .A1(n10968), .A2(n11367), .ZN(n12780) );
  INV_X1 U13029 ( .A(n19061), .ZN(n19049) );
  NAND2_X1 U13030 ( .A1(n13191), .A2(n13067), .ZN(n19269) );
  INV_X1 U13031 ( .A(n19171), .ZN(n19153) );
  AND2_X1 U13032 ( .A1(n19153), .A2(n19145), .ZN(n19151) );
  INV_X1 U13033 ( .A(n19161), .ZN(n19179) );
  OR2_X1 U13034 ( .A1(n19186), .A2(n19214), .ZN(n19183) );
  INV_X1 U13035 ( .A(n19186), .ZN(n19216) );
  INV_X1 U13036 ( .A(n12840), .ZN(n12901) );
  OR2_X1 U13037 ( .A1(n12780), .A2(n19231), .ZN(n19221) );
  INV_X1 U13038 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16216) );
  INV_X1 U13039 ( .A(n16269), .ZN(n19219) );
  NAND2_X1 U13040 ( .A1(n12780), .A2(n10928), .ZN(n16278) );
  OR2_X1 U13041 ( .A1(n11304), .A2(n19857), .ZN(n16326) );
  INV_X1 U13042 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15710) );
  AOI211_X2 U13043 ( .C1(n13779), .C2(n13785), .A(n19442), .B(n13778), .ZN(
        n19266) );
  INV_X1 U13044 ( .A(n19286), .ZN(n19294) );
  INV_X1 U13045 ( .A(n19324), .ZN(n19321) );
  NAND2_X1 U13046 ( .A1(n19301), .A2(n19300), .ZN(n19358) );
  INV_X1 U13047 ( .A(n19374), .ZN(n19365) );
  INV_X1 U13048 ( .A(n19395), .ZN(n19406) );
  INV_X1 U13049 ( .A(n19422), .ZN(n19434) );
  INV_X1 U13050 ( .A(n19457), .ZN(n19464) );
  NAND2_X1 U13051 ( .A1(n19436), .A2(n19439), .ZN(n19489) );
  OR2_X1 U13052 ( .A1(n19626), .A2(n19497), .ZN(n19515) );
  INV_X1 U13053 ( .A(n19555), .ZN(n19552) );
  INV_X1 U13054 ( .A(n19559), .ZN(n19575) );
  AOI21_X1 U13055 ( .B1(n13599), .B2(n13600), .A(n13598), .ZN(n19591) );
  INV_X1 U13056 ( .A(n19614), .ZN(n19625) );
  OR2_X1 U13057 ( .A1(n19626), .A2(n19819), .ZN(n19729) );
  INV_X1 U13058 ( .A(n19816), .ZN(n19731) );
  AOI21_X1 U13059 ( .B1(n18621), .B2(n18661), .A(n17378), .ZN(n18854) );
  NAND2_X1 U13060 ( .A1(n18838), .A2(n18680), .ZN(n16524) );
  INV_X1 U13061 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n21064) );
  INV_X1 U13062 ( .A(n16902), .ZN(n16894) );
  NOR2_X1 U13063 ( .A1(n16620), .A2(n16968), .ZN(n16973) );
  AND2_X1 U13064 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17037), .ZN(n17049) );
  AND3_X1 U13065 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(n17343), .ZN(n17335) );
  NOR2_X1 U13066 ( .A1(n17311), .A2(n17336), .ZN(n17343) );
  NOR3_X1 U13067 ( .A1(n17431), .A2(n17371), .A3(n17361), .ZN(n17367) );
  OR2_X1 U13068 ( .A1(n18835), .A2(n17380), .ZN(n17404) );
  INV_X1 U13069 ( .A(n17393), .ZN(n17407) );
  INV_X1 U13070 ( .A(n17380), .ZN(n17436) );
  INV_X1 U13071 ( .A(n17486), .ZN(n17479) );
  NAND2_X1 U13072 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17793), .ZN(n17696) );
  INV_X1 U13073 ( .A(n17852), .ZN(n17842) );
  INV_X1 U13074 ( .A(n17768), .ZN(n17742) );
  AOI22_X1 U13075 ( .A1(n18049), .A2(n17850), .B1(n17770), .B2(n18050), .ZN(
        n17755) );
  INV_X1 U13076 ( .A(n16375), .ZN(n17861) );
  INV_X1 U13077 ( .A(n18158), .ZN(n18173) );
  INV_X1 U13078 ( .A(n18093), .ZN(n18070) );
  INV_X1 U13079 ( .A(n18153), .ZN(n18159) );
  INV_X1 U13080 ( .A(n18172), .ZN(n18166) );
  INV_X1 U13081 ( .A(n18614), .ZN(n18263) );
  INV_X1 U13082 ( .A(n18353), .ZN(n18351) );
  INV_X1 U13083 ( .A(n18398), .ZN(n18393) );
  INV_X1 U13084 ( .A(n18435), .ZN(n18446) );
  INV_X1 U13085 ( .A(n18511), .ZN(n18519) );
  INV_X1 U13086 ( .A(n18838), .ZN(n18690) );
  INV_X1 U13087 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18790) );
  INV_X1 U13088 ( .A(n18787), .ZN(n18703) );
  INV_X1 U13089 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18718) );
  INV_X1 U13090 ( .A(n16473), .ZN(n16477) );
  NAND2_X1 U13091 ( .A1(n12750), .A2(n12749), .ZN(P1_U2842) );
  OR2_X1 U13092 ( .A1(n11747), .A2(n11746), .ZN(P3_U2834) );
  INV_X1 U13093 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14037) );
  AOI22_X1 U13094 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14929), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10177) );
  AND2_X4 U13095 ( .A1(n10403), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10398) );
  AOI22_X1 U13096 ( .A1(n10257), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10398), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10176) );
  AND2_X4 U13097 ( .A1(n13481), .A2(n13462), .ZN(n14757) );
  NOR2_X2 U13098 ( .A1(n10173), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10386) );
  AND2_X4 U13099 ( .A1(n10386), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14748) );
  AOI22_X1 U13100 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n14748), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10175) );
  AND2_X4 U13101 ( .A1(n10387), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10392) );
  AOI22_X1 U13102 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9668), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10174) );
  NAND4_X1 U13103 ( .A1(n10177), .A2(n10176), .A3(n10175), .A4(n10174), .ZN(
        n10183) );
  AOI22_X1 U13104 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14929), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10181) );
  AOI22_X1 U13105 ( .A1(n10257), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n10398), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10180) );
  AOI22_X1 U13106 ( .A1(n14757), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10179) );
  AOI22_X1 U13107 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9668), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10178) );
  NAND4_X1 U13108 ( .A1(n10181), .A2(n10180), .A3(n10179), .A4(n10178), .ZN(
        n10182) );
  MUX2_X2 U13109 ( .A(n10183), .B(n10182), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19244) );
  AOI22_X1 U13110 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14929), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10185) );
  AOI22_X1 U13111 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10188) );
  AOI22_X1 U13112 ( .A1(n14757), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10398), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10187) );
  AOI22_X1 U13113 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14929), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10194) );
  BUF_X4 U13114 ( .A(n10257), .Z(n14927) );
  AOI22_X1 U13115 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10398), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10193) );
  AOI22_X1 U13116 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n9645), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10192) );
  AOI22_X1 U13117 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10191) );
  NAND4_X1 U13118 ( .A1(n10194), .A2(n10193), .A3(n10192), .A4(n10191), .ZN(
        n10195) );
  NAND2_X1 U13119 ( .A1(n10195), .A2(n9846), .ZN(n10196) );
  AOI22_X1 U13120 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14929), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U13121 ( .A1(n14757), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14748), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10200) );
  AOI22_X1 U13122 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10199) );
  AOI22_X1 U13123 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10398), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10198) );
  NAND4_X1 U13124 ( .A1(n10201), .A2(n10200), .A3(n10199), .A4(n10198), .ZN(
        n10202) );
  NAND2_X1 U13125 ( .A1(n10202), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10210) );
  AOI22_X1 U13126 ( .A1(n10257), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10398), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10205) );
  AOI22_X1 U13127 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n9645), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10204) );
  AOI22_X1 U13128 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(n9668), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10203) );
  NAND3_X1 U13129 ( .A1(n10205), .A2(n10204), .A3(n10203), .ZN(n10208) );
  AOI22_X1 U13130 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14929), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10206) );
  INV_X1 U13131 ( .A(n10206), .ZN(n10207) );
  OAI21_X1 U13132 ( .B1(n10208), .B2(n10207), .A(n9846), .ZN(n10209) );
  AOI22_X1 U13133 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14929), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10214) );
  AOI22_X1 U13134 ( .A1(n10257), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10398), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U13135 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(n9669), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U13136 ( .A1(n14757), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10211) );
  NAND4_X1 U13137 ( .A1(n10214), .A2(n10213), .A3(n10212), .A4(n10211), .ZN(
        n10215) );
  AOI22_X1 U13138 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14929), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10219) );
  AOI22_X1 U13139 ( .A1(n10257), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n10398), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10218) );
  AOI22_X1 U13140 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10217) );
  AOI22_X1 U13141 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9669), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10216) );
  NAND4_X1 U13142 ( .A1(n10219), .A2(n10218), .A3(n10217), .A4(n10216), .ZN(
        n10220) );
  NAND2_X1 U13143 ( .A1(n10220), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10221) );
  AOI22_X1 U13144 ( .A1(n14929), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10227) );
  AOI22_X1 U13145 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10184), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10226) );
  AOI22_X1 U13146 ( .A1(n14748), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9668), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10225) );
  AOI22_X1 U13147 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10398), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10224) );
  NAND4_X1 U13148 ( .A1(n10227), .A2(n10226), .A3(n10225), .A4(n10224), .ZN(
        n10233) );
  AOI22_X1 U13149 ( .A1(n14748), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14826), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10231) );
  AOI22_X1 U13150 ( .A1(n14757), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10398), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10230) );
  AOI22_X1 U13151 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14929), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10229) );
  AOI22_X1 U13152 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9669), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10228) );
  NAND4_X1 U13153 ( .A1(n10231), .A2(n10230), .A3(n10229), .A4(n10228), .ZN(
        n10232) );
  MUX2_X2 U13154 ( .A(n10233), .B(n10232), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10294) );
  AOI22_X1 U13155 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n14929), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10237) );
  AOI22_X1 U13156 ( .A1(n10257), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10398), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10236) );
  AOI22_X1 U13157 ( .A1(n14757), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n14748), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10235) );
  AOI22_X1 U13158 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(n9669), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10234) );
  NAND4_X1 U13159 ( .A1(n10237), .A2(n10236), .A3(n10235), .A4(n10234), .ZN(
        n10243) );
  AOI22_X1 U13160 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14929), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10241) );
  AOI22_X1 U13161 ( .A1(n10257), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10398), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10240) );
  AOI22_X1 U13162 ( .A1(n14757), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10239) );
  AOI22_X1 U13163 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9669), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10238) );
  NAND4_X1 U13164 ( .A1(n10241), .A2(n10240), .A3(n10239), .A4(n10238), .ZN(
        n10242) );
  MUX2_X2 U13165 ( .A(n10243), .B(n10242), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19251) );
  INV_X2 U13166 ( .A(n19251), .ZN(n12978) );
  AND2_X1 U13167 ( .A1(n19251), .A2(n10294), .ZN(n10262) );
  AOI22_X1 U13168 ( .A1(n14757), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14748), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10247) );
  AOI22_X1 U13169 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10398), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10246) );
  AOI22_X1 U13170 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14929), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10245) );
  AOI22_X1 U13171 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9669), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10244) );
  AOI22_X1 U13172 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10398), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10251) );
  AOI22_X1 U13173 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14748), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10250) );
  AOI22_X1 U13174 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14929), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10249) );
  AOI22_X1 U13175 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9668), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10248) );
  NAND3_X1 U13176 ( .A1(n10774), .A2(n11041), .A3(n11027), .ZN(n10252) );
  AOI22_X1 U13177 ( .A1(n14927), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n14929), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U13178 ( .A1(n14757), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10398), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U13179 ( .A1(n10397), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9669), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10253) );
  AOI22_X1 U13180 ( .A1(n10184), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14929), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10261) );
  AOI22_X1 U13181 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10398), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10260) );
  AOI22_X1 U13182 ( .A1(n14748), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10257), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10259) );
  AOI22_X1 U13183 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9668), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10258) );
  NAND2_X1 U13184 ( .A1(n10269), .A2(n10265), .ZN(n10277) );
  MUX2_X1 U13185 ( .A(n19251), .B(n19257), .S(n19244), .Z(n10264) );
  INV_X1 U13186 ( .A(n10262), .ZN(n10263) );
  NAND4_X1 U13187 ( .A1(n10277), .A2(n10264), .A3(n10263), .A4(n11041), .ZN(
        n10267) );
  NOR2_X1 U13188 ( .A1(n12971), .A2(n19244), .ZN(n10266) );
  AND2_X1 U13189 ( .A1(n11029), .A2(n13434), .ZN(n10297) );
  AND2_X1 U13190 ( .A1(n19257), .A2(n19251), .ZN(n12973) );
  NAND3_X1 U13191 ( .A1(n10266), .A2(n10297), .A3(n12973), .ZN(n12924) );
  NAND2_X1 U13192 ( .A1(n10267), .A2(n12924), .ZN(n11031) );
  INV_X1 U13193 ( .A(n19257), .ZN(n12986) );
  INV_X1 U13194 ( .A(n10976), .ZN(n10270) );
  AND2_X2 U13195 ( .A1(n10983), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10285) );
  NAND2_X1 U13196 ( .A1(n11039), .A2(n10285), .ZN(n10272) );
  NAND2_X1 U13197 ( .A1(n10340), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10284) );
  NOR2_X1 U13198 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12783) );
  INV_X1 U13199 ( .A(n12783), .ZN(n10281) );
  INV_X2 U13200 ( .A(n9677), .ZN(n10273) );
  NAND2_X1 U13201 ( .A1(n10273), .A2(n10274), .ZN(n10292) );
  NAND2_X1 U13202 ( .A1(n10292), .A2(n10984), .ZN(n11032) );
  NAND3_X1 U13203 ( .A1(n11032), .A2(n19257), .A3(n19244), .ZN(n10280) );
  NOR2_X1 U13204 ( .A1(n19251), .A2(n10294), .ZN(n10275) );
  NAND2_X1 U13205 ( .A1(n10275), .A2(n10274), .ZN(n10276) );
  NAND2_X1 U13206 ( .A1(n10276), .A2(n11029), .ZN(n10278) );
  NAND2_X1 U13207 ( .A1(n10278), .A2(n10277), .ZN(n10279) );
  NOR2_X1 U13208 ( .A1(n10265), .A2(n13434), .ZN(n11033) );
  NAND3_X2 U13209 ( .A1(n10285), .A2(n11034), .A3(n11041), .ZN(n10311) );
  OAI211_X1 U13210 ( .C1(n10281), .C2(n19855), .A(n10304), .B(n10311), .ZN(
        n10282) );
  INV_X1 U13211 ( .A(n10282), .ZN(n10283) );
  NAND2_X1 U13212 ( .A1(n10284), .A2(n10283), .ZN(n10348) );
  INV_X1 U13213 ( .A(n10979), .ZN(n10969) );
  INV_X1 U13214 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n12852) );
  NAND2_X1 U13215 ( .A1(n10329), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10289) );
  INV_X2 U13216 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15457) );
  NOR2_X1 U13217 ( .A1(n15457), .A2(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10286) );
  NOR2_X1 U13218 ( .A1(n11361), .A2(n10286), .ZN(n10287) );
  INV_X1 U13219 ( .A(n10165), .ZN(n11040) );
  NAND3_X1 U13220 ( .A1(n11039), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n11040), 
        .ZN(n10290) );
  NOR2_X1 U13221 ( .A1(n13434), .A2(n10294), .ZN(n10293) );
  NAND2_X1 U13222 ( .A1(n11029), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10302) );
  AND2_X1 U13223 ( .A1(n10294), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10296) );
  NOR2_X1 U13224 ( .A1(n19244), .A2(n9678), .ZN(n10295) );
  NAND4_X1 U13225 ( .A1(n10297), .A2(n12973), .A3(n10296), .A4(n10295), .ZN(
        n10301) );
  NOR2_X1 U13226 ( .A1(n19251), .A2(n16342), .ZN(n13000) );
  OAI211_X2 U13227 ( .C1(n11019), .C2(n10302), .A(n10301), .B(n10300), .ZN(
        n10308) );
  NAND2_X1 U13228 ( .A1(n10308), .A2(n19231), .ZN(n10303) );
  NAND2_X1 U13229 ( .A1(n9670), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10305) );
  NAND2_X1 U13230 ( .A1(n10340), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10310) );
  AND2_X1 U13231 ( .A1(n12783), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n10307) );
  NOR2_X1 U13232 ( .A1(n10308), .A2(n10307), .ZN(n10309) );
  NAND2_X2 U13233 ( .A1(n10310), .A2(n10309), .ZN(n10335) );
  INV_X1 U13234 ( .A(n10335), .ZN(n10316) );
  NAND2_X1 U13235 ( .A1(n9670), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10314) );
  INV_X1 U13236 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13006) );
  OAI22_X1 U13237 ( .A1(n10311), .A2(n13006), .B1(n15457), .B2(n12863), .ZN(
        n10312) );
  AOI21_X1 U13238 ( .B1(n10329), .B2(P2_REIP_REG_1__SCAN_IN), .A(n10312), .ZN(
        n10313) );
  NAND2_X1 U13239 ( .A1(n10316), .A2(n10315), .ZN(n10336) );
  NAND2_X1 U13240 ( .A1(n10340), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10319) );
  OAI21_X1 U13241 ( .B1(n19837), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n15457), 
        .ZN(n10317) );
  NAND3_X1 U13242 ( .A1(n10337), .A2(n10336), .A3(n10323), .ZN(n10327) );
  NAND2_X1 U13243 ( .A1(n10323), .A2(n10335), .ZN(n10320) );
  OAI21_X1 U13244 ( .B1(n10335), .B2(n10323), .A(n10315), .ZN(n10321) );
  NAND2_X1 U13245 ( .A1(n10322), .A2(n10321), .ZN(n10326) );
  NAND2_X1 U13246 ( .A1(n10328), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10334) );
  INV_X1 U13247 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10331) );
  INV_X1 U13248 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n14201) );
  OAI22_X1 U13249 ( .A1(n10311), .A2(n10331), .B1(n15457), .B2(n14201), .ZN(
        n10332) );
  OAI21_X1 U13250 ( .B1(n10353), .B2(n10337), .A(n10336), .ZN(n10339) );
  NAND2_X1 U13251 ( .A1(n10340), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10342) );
  NAND2_X1 U13252 ( .A1(n12783), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10341) );
  NAND2_X1 U13253 ( .A1(n10328), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10346) );
  INV_X1 U13254 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13069) );
  OAI22_X1 U13255 ( .A1(n10311), .A2(n13069), .B1(n15457), .B2(n10343), .ZN(
        n10344) );
  AOI21_X1 U13256 ( .B1(n11313), .B2(P2_REIP_REG_3__SCAN_IN), .A(n10344), .ZN(
        n10345) );
  NAND2_X1 U13257 ( .A1(n10346), .A2(n10345), .ZN(n10831) );
  INV_X1 U13258 ( .A(n10364), .ZN(n10352) );
  INV_X1 U13259 ( .A(n10348), .ZN(n10350) );
  NAND2_X1 U13260 ( .A1(n10350), .A2(n10349), .ZN(n10351) );
  NAND2_X1 U13261 ( .A1(n10352), .A2(n16328), .ZN(n10379) );
  BUF_X4 U13262 ( .A(n10356), .Z(n14657) );
  INV_X1 U13263 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11178) );
  AND2_X2 U13264 ( .A1(n10378), .A2(n10375), .ZN(n19383) );
  INV_X1 U13265 ( .A(n10360), .ZN(n10361) );
  AND2_X2 U13266 ( .A1(n10376), .A2(n10377), .ZN(n10579) );
  AOI22_X1 U13267 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19383), .B1(
        n10579), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10362) );
  AND2_X1 U13268 ( .A1(n14673), .A2(n16328), .ZN(n10373) );
  AND2_X2 U13269 ( .A1(n10378), .A2(n10373), .ZN(n13541) );
  AND2_X2 U13270 ( .A1(n10378), .A2(n10374), .ZN(n10580) );
  AOI22_X1 U13271 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n13541), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10372) );
  INV_X1 U13272 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11177) );
  AND2_X1 U13273 ( .A1(n10380), .A2(n10377), .ZN(n10365) );
  INV_X1 U13274 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11175) );
  OAI22_X1 U13275 ( .A1(n11177), .A2(n13423), .B1(n19677), .B2(n11175), .ZN(
        n10370) );
  INV_X1 U13276 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14038) );
  AND2_X1 U13277 ( .A1(n14657), .A2(n10375), .ZN(n10367) );
  AND2_X1 U13278 ( .A1(n10380), .A2(n10375), .ZN(n10368) );
  INV_X1 U13279 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14039) );
  OAI22_X1 U13280 ( .A1(n14038), .A2(n10417), .B1(n10571), .B2(n14039), .ZN(
        n10369) );
  NOR2_X1 U13281 ( .A1(n10370), .A2(n10369), .ZN(n10371) );
  AOI22_X1 U13282 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n13783), .B1(
        n19295), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10385) );
  AND2_X2 U13283 ( .A1(n10378), .A2(n10377), .ZN(n10416) );
  AOI22_X1 U13284 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19267), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10384) );
  OR2_X2 U13285 ( .A1(n10379), .A2(n14673), .ZN(n10381) );
  NOR2_X2 U13286 ( .A1(n10381), .A2(n14657), .ZN(n10582) );
  NAND2_X1 U13287 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10383) );
  NOR2_X2 U13288 ( .A1(n10381), .A2(n10357), .ZN(n10581) );
  NAND2_X1 U13289 ( .A1(n10581), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10382) );
  INV_X1 U13290 ( .A(n10467), .ZN(n11236) );
  INV_X1 U13291 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10389) );
  INV_X1 U13292 ( .A(n14767), .ZN(n10529) );
  INV_X1 U13293 ( .A(n14766), .ZN(n10528) );
  INV_X1 U13294 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10388) );
  OAI22_X1 U13295 ( .A1(n10389), .A2(n10529), .B1(n10528), .B2(n10388), .ZN(
        n10390) );
  AOI21_X1 U13296 ( .B1(n11236), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n10390), .ZN(n10396) );
  AND2_X2 U13297 ( .A1(n14748), .A2(n9846), .ZN(n10426) );
  AND2_X2 U13298 ( .A1(n14826), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10447) );
  AOI22_X1 U13299 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10447), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10395) );
  INV_X1 U13300 ( .A(n10472), .ZN(n14770) );
  AOI22_X1 U13301 ( .A1(n14770), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14771), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10394) );
  NAND2_X1 U13302 ( .A1(n14929), .A2(n9846), .ZN(n10473) );
  INV_X1 U13303 ( .A(n10473), .ZN(n10533) );
  INV_X1 U13304 ( .A(n10392), .ZN(n13290) );
  INV_X1 U13305 ( .A(n11114), .ZN(n10532) );
  AOI22_X1 U13306 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n10533), .B1(
        n10532), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10393) );
  INV_X1 U13307 ( .A(n10463), .ZN(n14733) );
  NAND2_X1 U13308 ( .A1(n14929), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10464) );
  INV_X1 U13309 ( .A(n10464), .ZN(n14734) );
  AOI22_X1 U13310 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n14733), .B1(
        n14734), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10406) );
  INV_X1 U13311 ( .A(n14784), .ZN(n14730) );
  INV_X1 U13312 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10401) );
  INV_X1 U13313 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19243) );
  AND2_X1 U13314 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10400) );
  INV_X1 U13315 ( .A(n14782), .ZN(n14727) );
  OAI22_X1 U13316 ( .A1(n14730), .A2(n10401), .B1(n19243), .B2(n14727), .ZN(
        n10402) );
  AOI22_X1 U13317 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10405) );
  NAND2_X1 U13318 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10404) );
  INV_X1 U13319 ( .A(n10510), .ZN(n11091) );
  NAND2_X1 U13320 ( .A1(n11091), .A2(n19231), .ZN(n10407) );
  INV_X1 U13321 ( .A(n10484), .ZN(n10482) );
  INV_X1 U13322 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13821) );
  INV_X1 U13323 ( .A(n10571), .ZN(n19501) );
  AOI21_X1 U13324 ( .B1(n19501), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n19231), .ZN(n10409) );
  INV_X1 U13325 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11138) );
  OR2_X1 U13326 ( .A1(n19677), .A2(n11138), .ZN(n10408) );
  OAI211_X1 U13327 ( .C1(n10410), .C2(n13821), .A(n10409), .B(n10408), .ZN(
        n10415) );
  AOI22_X1 U13328 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n13541), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10413) );
  NAND2_X1 U13329 ( .A1(n10581), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10412) );
  NAND2_X1 U13330 ( .A1(n10582), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n10411) );
  NAND3_X1 U13331 ( .A1(n10413), .A2(n10412), .A3(n10411), .ZN(n10414) );
  AOI22_X1 U13332 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n13783), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10423) );
  INV_X1 U13333 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11140) );
  NOR2_X1 U13334 ( .A1(n19466), .A2(n11140), .ZN(n10419) );
  INV_X1 U13335 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13829) );
  INV_X1 U13336 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n19562) );
  OAI22_X1 U13337 ( .A1(n13829), .A2(n10417), .B1(n13423), .B2(n19562), .ZN(
        n10418) );
  NOR2_X1 U13338 ( .A1(n10419), .A2(n10418), .ZN(n10422) );
  AOI22_X1 U13339 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19295), .B1(
        n19383), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10421) );
  INV_X1 U13340 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13843) );
  AOI22_X1 U13341 ( .A1(n14767), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10424) );
  OAI21_X1 U13342 ( .B1(n10467), .B2(n13843), .A(n10424), .ZN(n10425) );
  INV_X1 U13343 ( .A(n10425), .ZN(n10433) );
  AOI22_X1 U13344 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10447), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10432) );
  INV_X1 U13345 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13440) );
  INV_X1 U13346 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13853) );
  OAI22_X1 U13347 ( .A1(n10472), .A2(n13440), .B1(n14738), .B2(n13853), .ZN(
        n10427) );
  INV_X1 U13348 ( .A(n10427), .ZN(n10431) );
  INV_X1 U13349 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10428) );
  INV_X1 U13350 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11118) );
  OAI22_X1 U13351 ( .A1(n10473), .A2(n10428), .B1(n11114), .B2(n11118), .ZN(
        n10429) );
  INV_X1 U13352 ( .A(n10429), .ZN(n10430) );
  NAND4_X1 U13353 ( .A1(n10433), .A2(n10432), .A3(n10431), .A4(n10430), .ZN(
        n10440) );
  INV_X1 U13354 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13851) );
  INV_X1 U13355 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11122) );
  OAI22_X1 U13356 ( .A1(n10463), .A2(n13851), .B1(n10464), .B2(n11122), .ZN(
        n10434) );
  INV_X1 U13357 ( .A(n10434), .ZN(n10438) );
  AOI22_X1 U13358 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14782), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10437) );
  AOI22_X1 U13359 ( .A1(n14783), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10436) );
  NAND2_X1 U13360 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10435) );
  NAND4_X1 U13361 ( .A1(n10438), .A2(n10437), .A3(n10436), .A4(n10435), .ZN(
        n10439) );
  AND2_X1 U13362 ( .A1(n19231), .A2(n10782), .ZN(n12849) );
  AOI22_X1 U13363 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10444) );
  NAND2_X1 U13364 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10443) );
  NAND2_X1 U13365 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10442) );
  INV_X1 U13366 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19236) );
  NAND2_X1 U13367 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10441) );
  NAND4_X1 U13368 ( .A1(n10444), .A2(n10443), .A3(n10442), .A4(n10441), .ZN(
        n10446) );
  INV_X1 U13369 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13828) );
  OAI22_X1 U13370 ( .A1(n13828), .A2(n10463), .B1(n10464), .B2(n11138), .ZN(
        n10445) );
  NOR2_X1 U13371 ( .A1(n10446), .A2(n10445), .ZN(n10457) );
  INV_X1 U13372 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13820) );
  OR2_X1 U13373 ( .A1(n10467), .A2(n13820), .ZN(n10451) );
  AOI22_X1 U13374 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10450) );
  NAND2_X1 U13375 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10449) );
  NAND2_X1 U13376 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10448) );
  AND4_X1 U13377 ( .A1(n10451), .A2(n10450), .A3(n10449), .A4(n10448), .ZN(
        n10456) );
  INV_X1 U13378 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13831) );
  OAI22_X1 U13379 ( .A1(n10472), .A2(n19562), .B1(n14738), .B2(n13831), .ZN(
        n10454) );
  INV_X1 U13380 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10452) );
  OAI22_X1 U13381 ( .A1(n10452), .A2(n10473), .B1(n11114), .B2(n11140), .ZN(
        n10453) );
  NOR2_X1 U13382 ( .A1(n10454), .A2(n10453), .ZN(n10455) );
  INV_X1 U13383 ( .A(n11081), .ZN(n10458) );
  NAND2_X1 U13384 ( .A1(n12849), .A2(n10458), .ZN(n10779) );
  AOI22_X1 U13385 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U13386 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10461) );
  NAND2_X1 U13387 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10460) );
  NAND2_X1 U13388 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n10459) );
  NAND4_X1 U13389 ( .A1(n10462), .A2(n10461), .A3(n10460), .A4(n10459), .ZN(
        n10466) );
  INV_X1 U13390 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14014) );
  INV_X1 U13391 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11157) );
  OAI22_X1 U13392 ( .A1(n14014), .A2(n10463), .B1(n10464), .B2(n11157), .ZN(
        n10465) );
  NOR2_X1 U13393 ( .A1(n10466), .A2(n10465), .ZN(n10479) );
  INV_X1 U13394 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14008) );
  OR2_X1 U13395 ( .A1(n10467), .A2(n14008), .ZN(n10471) );
  AOI22_X1 U13396 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10470) );
  NAND2_X1 U13397 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10469) );
  NAND2_X1 U13398 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10468) );
  AND4_X1 U13399 ( .A1(n10471), .A2(n10470), .A3(n10469), .A4(n10468), .ZN(
        n10478) );
  INV_X1 U13400 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13437) );
  INV_X1 U13401 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14017) );
  OAI22_X1 U13402 ( .A1(n10472), .A2(n13437), .B1(n14738), .B2(n14017), .ZN(
        n10476) );
  INV_X1 U13403 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10474) );
  INV_X1 U13404 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11153) );
  OAI22_X1 U13405 ( .A1(n10474), .A2(n10473), .B1(n11114), .B2(n11153), .ZN(
        n10475) );
  NOR2_X1 U13406 ( .A1(n10476), .A2(n10475), .ZN(n10477) );
  INV_X1 U13407 ( .A(n10483), .ZN(n10481) );
  NAND2_X1 U13408 ( .A1(n10482), .A2(n10481), .ZN(n10485) );
  INV_X1 U13409 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14779) );
  NAND2_X1 U13410 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10486) );
  OAI21_X1 U13411 ( .B1(n10467), .B2(n14779), .A(n10486), .ZN(n10490) );
  INV_X1 U13412 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14924) );
  NAND2_X1 U13413 ( .A1(n14766), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10488) );
  NAND2_X1 U13414 ( .A1(n14767), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10487) );
  OAI211_X1 U13415 ( .C1(n10472), .C2(n14924), .A(n10488), .B(n10487), .ZN(
        n10489) );
  NOR2_X1 U13416 ( .A1(n10490), .A2(n10489), .ZN(n10503) );
  INV_X1 U13417 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11257) );
  INV_X1 U13418 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11252) );
  OAI22_X1 U13419 ( .A1(n11257), .A2(n10463), .B1(n10464), .B2(n11252), .ZN(
        n10491) );
  INV_X1 U13420 ( .A(n10491), .ZN(n10502) );
  AOI22_X1 U13421 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10495) );
  NAND2_X1 U13422 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10494) );
  NAND2_X1 U13423 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10493) );
  NAND2_X1 U13424 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10492) );
  NAND2_X1 U13425 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10499) );
  NAND2_X1 U13426 ( .A1(n14771), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10498) );
  NAND2_X1 U13427 ( .A1(n10533), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10497) );
  NAND2_X1 U13428 ( .A1(n10532), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10496) );
  INV_X1 U13429 ( .A(n10780), .ZN(n11083) );
  MUX2_X1 U13430 ( .A(n19846), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10988) );
  NAND2_X1 U13431 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19855), .ZN(
        n10515) );
  NAND2_X1 U13432 ( .A1(n10988), .A2(n10756), .ZN(n10757) );
  NAND2_X1 U13433 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n19846), .ZN(
        n10504) );
  NAND2_X1 U13434 ( .A1(n10757), .A2(n10504), .ZN(n10509) );
  NAND2_X1 U13435 ( .A1(n13462), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10507) );
  OAI21_X1 U13436 ( .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n13462), .A(
        n10507), .ZN(n10505) );
  XNOR2_X1 U13437 ( .A(n10509), .B(n10505), .ZN(n10986) );
  MUX2_X1 U13438 ( .A(n11083), .B(n10986), .S(n10984), .Z(n10766) );
  MUX2_X1 U13439 ( .A(n10331), .B(n10766), .S(n13441), .Z(n10522) );
  MUX2_X1 U13440 ( .A(n11081), .B(P2_EBX_REG_1__SCAN_IN), .S(n9649), .Z(n10506) );
  INV_X1 U13441 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n19058) );
  NOR2_X1 U13442 ( .A1(n13441), .A2(n19058), .ZN(n10517) );
  NOR2_X1 U13443 ( .A1(n10506), .A2(n10517), .ZN(n10520) );
  NAND2_X1 U13444 ( .A1(n10522), .A2(n10520), .ZN(n10512) );
  AND2_X1 U13445 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n19837), .ZN(
        n10508) );
  MUX2_X1 U13446 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n19829), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n10545) );
  XNOR2_X1 U13447 ( .A(n10546), .B(n10545), .ZN(n10750) );
  MUX2_X1 U13448 ( .A(n10770), .B(P2_EBX_REG_3__SCAN_IN), .S(n9649), .Z(n10511) );
  INV_X1 U13449 ( .A(n10550), .ZN(n10553) );
  NAND2_X1 U13450 ( .A1(n10512), .A2(n10511), .ZN(n10513) );
  NAND2_X1 U13451 ( .A1(n10553), .A2(n10513), .ZN(n13661) );
  NAND2_X1 U13452 ( .A1(n10525), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13578) );
  INV_X1 U13453 ( .A(n10782), .ZN(n11074) );
  OAI21_X1 U13454 ( .B1(n19855), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n10515), .ZN(n10990) );
  MUX2_X1 U13455 ( .A(n11074), .B(n10990), .S(n10984), .Z(n10769) );
  INV_X1 U13456 ( .A(n10517), .ZN(n10516) );
  OAI21_X1 U13457 ( .B1(n10769), .B2(n9649), .A(n10516), .ZN(n19056) );
  NAND2_X1 U13458 ( .A1(n19056), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12859) );
  AND2_X1 U13459 ( .A1(n10517), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10518) );
  OR2_X1 U13460 ( .A1(n10520), .A2(n10518), .ZN(n14669) );
  NOR2_X1 U13461 ( .A1(n12859), .A2(n14669), .ZN(n10519) );
  NAND2_X1 U13462 ( .A1(n12859), .A2(n14669), .ZN(n12858) );
  OAI21_X1 U13463 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10519), .A(
        n12858), .ZN(n14184) );
  INV_X1 U13464 ( .A(n10520), .ZN(n10521) );
  XNOR2_X1 U13465 ( .A(n10522), .B(n10521), .ZN(n14656) );
  XNOR2_X1 U13466 ( .A(n14656), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14183) );
  OR2_X1 U13467 ( .A1(n14184), .A2(n14183), .ZN(n14205) );
  NAND2_X1 U13468 ( .A1(n14656), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10523) );
  NAND2_X1 U13469 ( .A1(n14205), .A2(n10523), .ZN(n13580) );
  INV_X1 U13470 ( .A(n13580), .ZN(n10524) );
  NAND2_X1 U13471 ( .A1(n13578), .A2(n10524), .ZN(n10526) );
  INV_X1 U13472 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n10549) );
  INV_X1 U13473 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10530) );
  INV_X1 U13474 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10527) );
  OAI22_X1 U13475 ( .A1(n10530), .A2(n10529), .B1(n10528), .B2(n10527), .ZN(
        n10531) );
  AOI21_X1 U13476 ( .B1(n11236), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n10531), .ZN(n10537) );
  AOI22_X1 U13477 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10447), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10536) );
  AOI22_X1 U13478 ( .A1(n14770), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n14771), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10535) );
  AOI22_X1 U13479 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10533), .B1(
        n10532), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10534) );
  NAND4_X1 U13480 ( .A1(n10537), .A2(n10536), .A3(n10535), .A4(n10534), .ZN(
        n10544) );
  AOI22_X1 U13481 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n14733), .B1(
        n14734), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10542) );
  INV_X1 U13482 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19248) );
  NOR2_X1 U13483 ( .A1(n14727), .A2(n19248), .ZN(n10538) );
  AOI21_X1 U13484 ( .B1(n14784), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n10538), .ZN(n10541) );
  AOI22_X1 U13485 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10540) );
  NAND2_X1 U13486 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10539) );
  NAND4_X1 U13487 ( .A1(n10542), .A2(n10541), .A3(n10540), .A4(n10539), .ZN(
        n10543) );
  NAND2_X1 U13488 ( .A1(n19829), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10547) );
  NOR2_X1 U13489 ( .A1(n15710), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10753) );
  NAND2_X1 U13490 ( .A1(n10755), .A2(n10753), .ZN(n10752) );
  MUX2_X1 U13491 ( .A(n11095), .B(n10752), .S(n10984), .Z(n10772) );
  MUX2_X1 U13492 ( .A(n10549), .B(n10772), .S(n13441), .Z(n10551) );
  INV_X1 U13493 ( .A(n10591), .ZN(n10555) );
  INV_X1 U13494 ( .A(n10551), .ZN(n10552) );
  NAND2_X1 U13495 ( .A1(n10553), .A2(n10552), .ZN(n10554) );
  NAND2_X1 U13496 ( .A1(n10555), .A2(n10554), .ZN(n19044) );
  INV_X1 U13497 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13750) );
  XNOR2_X1 U13498 ( .A(n19044), .B(n13750), .ZN(n13563) );
  OAI22_X2 U13499 ( .A1(n13564), .A2(n13563), .B1(n19044), .B2(n13750), .ZN(
        n13744) );
  AOI22_X1 U13500 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10559) );
  NAND2_X1 U13501 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n10558) );
  NAND2_X1 U13502 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10557) );
  NAND2_X1 U13503 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10556) );
  NAND4_X1 U13504 ( .A1(n10559), .A2(n10558), .A3(n10557), .A4(n10556), .ZN(
        n10562) );
  INV_X1 U13505 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10560) );
  INV_X1 U13506 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14715) );
  OAI22_X1 U13507 ( .A1(n10560), .A2(n10473), .B1(n10463), .B2(n14715), .ZN(
        n10561) );
  NOR2_X1 U13508 ( .A1(n10562), .A2(n10561), .ZN(n10570) );
  INV_X1 U13509 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14709) );
  AOI22_X1 U13510 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10563) );
  OAI21_X1 U13511 ( .B1(n10467), .B2(n14709), .A(n10563), .ZN(n10564) );
  INV_X1 U13512 ( .A(n10564), .ZN(n10569) );
  INV_X1 U13513 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13444) );
  INV_X1 U13514 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14718) );
  OAI22_X1 U13515 ( .A1(n10472), .A2(n13444), .B1(n14738), .B2(n14718), .ZN(
        n10566) );
  INV_X1 U13516 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11214) );
  INV_X1 U13517 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11212) );
  OAI22_X1 U13518 ( .A1(n11214), .A2(n11114), .B1(n10464), .B2(n11212), .ZN(
        n10565) );
  NOR2_X1 U13519 ( .A1(n10566), .A2(n10565), .ZN(n10568) );
  AOI22_X1 U13520 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10447), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10567) );
  NAND4_X1 U13521 ( .A1(n10570), .A2(n10569), .A3(n10568), .A4(n10567), .ZN(
        n11099) );
  AOI22_X1 U13522 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n13541), .B1(
        n19267), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10578) );
  AOI22_X1 U13523 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n10416), .B1(
        n19383), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10577) );
  OAI22_X1 U13524 ( .A1(n11212), .A2(n19677), .B1(n13423), .B2(n13444), .ZN(
        n10573) );
  INV_X1 U13525 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14716) );
  INV_X1 U13526 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14717) );
  OAI22_X1 U13527 ( .A1(n14716), .A2(n10417), .B1(n10571), .B2(n14717), .ZN(
        n10572) );
  NOR2_X1 U13528 ( .A1(n10573), .A2(n10572), .ZN(n10576) );
  INV_X1 U13529 ( .A(n10574), .ZN(n10575) );
  NAND4_X1 U13530 ( .A1(n10578), .A2(n10577), .A3(n10576), .A4(n10575), .ZN(
        n10588) );
  AOI22_X1 U13531 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19295), .B1(
        n13783), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10586) );
  AOI22_X1 U13532 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n10579), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10585) );
  NAND2_X1 U13533 ( .A1(n19633), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10584) );
  NAND2_X1 U13534 ( .A1(n19530), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n10583) );
  NAND4_X1 U13535 ( .A1(n10583), .A2(n10585), .A3(n10584), .A4(n10586), .ZN(
        n10587) );
  XNOR2_X1 U13536 ( .A(n10793), .B(n10596), .ZN(n10797) );
  INV_X1 U13537 ( .A(n10797), .ZN(n10777) );
  NAND2_X1 U13538 ( .A1(n10777), .A2(n10640), .ZN(n10592) );
  INV_X1 U13539 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n10839) );
  MUX2_X1 U13540 ( .A(n10839), .B(n11099), .S(n13441), .Z(n10590) );
  OAI21_X1 U13541 ( .B1(n10591), .B2(n10590), .A(n10637), .ZN(n19030) );
  INV_X1 U13542 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10796) );
  NAND2_X1 U13543 ( .A1(n13744), .A2(n13743), .ZN(n10595) );
  NAND2_X1 U13544 ( .A1(n10593), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10594) );
  NAND2_X1 U13545 ( .A1(n10595), .A2(n10594), .ZN(n13864) );
  INV_X1 U13546 ( .A(n10596), .ZN(n10597) );
  AOI22_X1 U13547 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19267), .B1(
        n10579), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U13548 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19383), .B1(
        n10580), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10604) );
  INV_X1 U13549 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11231) );
  OAI22_X1 U13550 ( .A1(n11231), .A2(n13423), .B1(n19677), .B2(n20919), .ZN(
        n10600) );
  INV_X1 U13551 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14739) );
  INV_X1 U13552 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14740) );
  OAI22_X1 U13553 ( .A1(n14739), .A2(n10417), .B1(n10571), .B2(n14740), .ZN(
        n10599) );
  NOR2_X1 U13554 ( .A1(n10600), .A2(n10599), .ZN(n10603) );
  INV_X1 U13555 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11227) );
  INV_X1 U13556 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14737) );
  INV_X1 U13557 ( .A(n10601), .ZN(n10602) );
  NAND4_X1 U13558 ( .A1(n10605), .A2(n10604), .A3(n10603), .A4(n10602), .ZN(
        n10613) );
  AOI22_X1 U13559 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n13541), .B1(
        n10416), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10611) );
  INV_X1 U13560 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19255) );
  INV_X1 U13561 ( .A(n13783), .ZN(n10606) );
  INV_X1 U13562 ( .A(n19295), .ZN(n19299) );
  INV_X1 U13563 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14728) );
  OAI22_X1 U13564 ( .A1(n19255), .A2(n10606), .B1(n19299), .B2(n14728), .ZN(
        n10607) );
  INV_X1 U13565 ( .A(n10607), .ZN(n10610) );
  NAND2_X1 U13566 ( .A1(n19633), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10609) );
  NAND2_X1 U13567 ( .A1(n19530), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10608) );
  NAND4_X1 U13568 ( .A1(n10611), .A2(n10610), .A3(n10609), .A4(n10608), .ZN(
        n10612) );
  AOI22_X1 U13569 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10617) );
  NAND2_X1 U13570 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n10616) );
  NAND2_X1 U13571 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10615) );
  NAND2_X1 U13572 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10614) );
  NAND4_X1 U13573 ( .A1(n10617), .A2(n10616), .A3(n10615), .A4(n10614), .ZN(
        n10619) );
  OAI22_X1 U13574 ( .A1(n14737), .A2(n10463), .B1(n10464), .B2(n20919), .ZN(
        n10618) );
  NOR2_X1 U13575 ( .A1(n10619), .A2(n10618), .ZN(n10627) );
  INV_X1 U13576 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14899) );
  AOI22_X1 U13577 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10620) );
  OAI21_X1 U13578 ( .B1(n14899), .B2(n10467), .A(n10620), .ZN(n10621) );
  INV_X1 U13579 ( .A(n10621), .ZN(n10626) );
  INV_X1 U13580 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n14741) );
  OAI22_X1 U13581 ( .A1(n10472), .A2(n11231), .B1(n14738), .B2(n14741), .ZN(
        n10623) );
  INV_X1 U13582 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14729) );
  OAI22_X1 U13583 ( .A1(n14729), .A2(n10473), .B1(n11114), .B2(n11227), .ZN(
        n10622) );
  NOR2_X1 U13584 ( .A1(n10623), .A2(n10622), .ZN(n10625) );
  AOI22_X1 U13585 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10447), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10624) );
  NAND4_X1 U13586 ( .A1(n10627), .A2(n10626), .A3(n10625), .A4(n10624), .ZN(
        n11102) );
  INV_X1 U13587 ( .A(n11102), .ZN(n10628) );
  NAND2_X1 U13588 ( .A1(n19231), .A2(n10628), .ZN(n10629) );
  INV_X1 U13589 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13315) );
  MUX2_X1 U13590 ( .A(n13315), .B(n11102), .S(n13441), .Z(n10635) );
  XNOR2_X1 U13591 ( .A(n10637), .B(n10635), .ZN(n19017) );
  INV_X1 U13592 ( .A(n19017), .ZN(n10631) );
  INV_X1 U13593 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13901) );
  XNOR2_X1 U13594 ( .A(n10632), .B(n13901), .ZN(n13865) );
  NAND2_X1 U13595 ( .A1(n13864), .A2(n13865), .ZN(n10634) );
  NAND2_X1 U13596 ( .A1(n10632), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10633) );
  INV_X1 U13597 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10848) );
  MUX2_X1 U13598 ( .A(n10848), .B(n10962), .S(n13441), .Z(n10639) );
  NAND2_X1 U13599 ( .A1(n9649), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10644) );
  INV_X1 U13600 ( .A(n10644), .ZN(n10638) );
  XNOR2_X1 U13601 ( .A(n10647), .B(n10638), .ZN(n18999) );
  AND2_X1 U13602 ( .A1(n10962), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10814) );
  AND2_X1 U13603 ( .A1(n18999), .A2(n10814), .ZN(n16250) );
  XNOR2_X1 U13604 ( .A(n9760), .B(n10060), .ZN(n19009) );
  NAND2_X1 U13605 ( .A1(n18999), .A2(n10962), .ZN(n10641) );
  INV_X1 U13606 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16320) );
  NAND2_X1 U13607 ( .A1(n10641), .A2(n16320), .ZN(n16249) );
  OR2_X1 U13608 ( .A1(n19009), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16248) );
  AND2_X1 U13609 ( .A1(n16249), .A2(n16248), .ZN(n10642) );
  NAND2_X1 U13610 ( .A1(n9649), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10645) );
  XNOR2_X1 U13611 ( .A(n10646), .B(n10645), .ZN(n18989) );
  AOI21_X1 U13612 ( .B1(n18989), .B2(n10962), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15437) );
  NAND3_X1 U13613 ( .A1(n10649), .A2(n9649), .A3(P2_EBX_REG_10__SCAN_IN), .ZN(
        n10648) );
  NAND2_X1 U13614 ( .A1(n10648), .A2(n10735), .ZN(n10650) );
  OR2_X1 U13615 ( .A1(n10650), .A2(n10653), .ZN(n18979) );
  INV_X1 U13616 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10651) );
  OAI21_X1 U13617 ( .B1(n18979), .B2(n10640), .A(n10651), .ZN(n15230) );
  NAND2_X1 U13618 ( .A1(n9649), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10652) );
  OR2_X1 U13619 ( .A1(n10653), .A2(n10652), .ZN(n10655) );
  INV_X1 U13620 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13410) );
  NAND2_X1 U13621 ( .A1(n13410), .A2(n10653), .ZN(n10663) );
  INV_X1 U13622 ( .A(n10662), .ZN(n10654) );
  AOI21_X1 U13623 ( .B1(n18966), .B2(n10962), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16226) );
  INV_X1 U13624 ( .A(n18979), .ZN(n10657) );
  AND2_X1 U13625 ( .A1(n10962), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10656) );
  NAND2_X1 U13626 ( .A1(n10657), .A2(n10656), .ZN(n15229) );
  AND2_X1 U13627 ( .A1(n10962), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10658) );
  NAND2_X1 U13628 ( .A1(n18989), .A2(n10658), .ZN(n15231) );
  NAND2_X1 U13629 ( .A1(n15229), .A2(n15231), .ZN(n16223) );
  AND2_X1 U13630 ( .A1(n10962), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10659) );
  AND2_X1 U13631 ( .A1(n18966), .A2(n10659), .ZN(n16227) );
  NOR2_X1 U13632 ( .A1(n16223), .A2(n16227), .ZN(n10660) );
  NAND2_X1 U13633 ( .A1(n9649), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10661) );
  NAND3_X1 U13634 ( .A1(n9649), .A2(n10663), .A3(P2_EBX_REG_12__SCAN_IN), .ZN(
        n10664) );
  NAND2_X1 U13635 ( .A1(n10686), .A2(n10664), .ZN(n18957) );
  INV_X1 U13636 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10665) );
  NOR2_X1 U13637 ( .A1(n10666), .A2(n10665), .ZN(n15418) );
  NAND2_X1 U13638 ( .A1(n10666), .A2(n10665), .ZN(n15416) );
  INV_X1 U13639 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n13448) );
  NOR2_X1 U13640 ( .A1(n13441), .A2(n13448), .ZN(n10685) );
  NOR2_X1 U13641 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(P2_EBX_REG_14__SCAN_IN), 
        .ZN(n10667) );
  NOR2_X1 U13642 ( .A1(n13441), .A2(n10667), .ZN(n10668) );
  INV_X1 U13643 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n10877) );
  INV_X1 U13644 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n13920) );
  NAND2_X1 U13645 ( .A1(n10877), .A2(n13920), .ZN(n10669) );
  INV_X1 U13646 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n16181) );
  NOR2_X1 U13647 ( .A1(n13441), .A2(n16181), .ZN(n10700) );
  INV_X1 U13648 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10887) );
  NOR2_X1 U13649 ( .A1(n13441), .A2(n10887), .ZN(n10697) );
  INV_X1 U13650 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n16177) );
  NAND2_X1 U13651 ( .A1(n10695), .A2(n16177), .ZN(n10670) );
  AND3_X1 U13652 ( .A1(n10670), .A2(n9649), .A3(P2_EBX_REG_21__SCAN_IN), .ZN(
        n10671) );
  OR2_X1 U13653 ( .A1(n10716), .A2(n10671), .ZN(n18892) );
  OR2_X1 U13654 ( .A1(n18892), .A2(n10640), .ZN(n10672) );
  INV_X1 U13655 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15334) );
  NAND2_X1 U13656 ( .A1(n10672), .A2(n15334), .ZN(n15156) );
  NAND2_X1 U13657 ( .A1(n10673), .A2(n10877), .ZN(n10679) );
  NOR2_X1 U13658 ( .A1(n13441), .A2(n10877), .ZN(n10675) );
  INV_X1 U13659 ( .A(n10735), .ZN(n10674) );
  AOI21_X1 U13660 ( .B1(n10065), .B2(n10675), .A(n10674), .ZN(n10676) );
  NAND2_X1 U13661 ( .A1(n10679), .A2(n10676), .ZN(n18914) );
  XNOR2_X1 U13662 ( .A(n10677), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15218) );
  NOR2_X1 U13663 ( .A1(n13441), .A2(n13920), .ZN(n10678) );
  NAND2_X1 U13664 ( .A1(n10679), .A2(n10678), .ZN(n10680) );
  NAND2_X1 U13665 ( .A1(n10680), .A2(n10702), .ZN(n13919) );
  OR2_X1 U13666 ( .A1(n13919), .A2(n10640), .ZN(n10681) );
  INV_X1 U13667 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15626) );
  NAND2_X1 U13668 ( .A1(n10681), .A2(n15626), .ZN(n15205) );
  NAND2_X1 U13669 ( .A1(n10688), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10682) );
  MUX2_X1 U13670 ( .A(n10688), .B(n10682), .S(n9649), .Z(n10683) );
  OR2_X1 U13671 ( .A1(n10688), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10691) );
  NAND2_X1 U13672 ( .A1(n10683), .A2(n10691), .ZN(n18935) );
  INV_X1 U13673 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10684) );
  OAI21_X1 U13674 ( .B1(n18935), .B2(n10640), .A(n10684), .ZN(n16205) );
  NAND2_X1 U13675 ( .A1(n10686), .A2(n10685), .ZN(n10687) );
  NAND2_X1 U13676 ( .A1(n10688), .A2(n10687), .ZN(n18948) );
  OR2_X1 U13677 ( .A1(n18948), .A2(n10640), .ZN(n10690) );
  INV_X1 U13678 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10689) );
  AND2_X1 U13679 ( .A1(n10690), .A2(n10689), .ZN(n15149) );
  INV_X1 U13680 ( .A(n15149), .ZN(n15396) );
  NAND3_X1 U13681 ( .A1(n10691), .A2(n9649), .A3(P2_EBX_REG_15__SCAN_IN), .ZN(
        n10692) );
  NAND2_X1 U13682 ( .A1(n10065), .A2(n10692), .ZN(n18923) );
  OR2_X1 U13683 ( .A1(n18923), .A2(n10640), .ZN(n10693) );
  INV_X1 U13684 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15389) );
  NAND2_X1 U13685 ( .A1(n10693), .A2(n15389), .ZN(n15381) );
  AND4_X1 U13686 ( .A1(n15205), .A2(n16205), .A3(n15396), .A4(n15381), .ZN(
        n10704) );
  NAND2_X1 U13687 ( .A1(n9649), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10694) );
  XNOR2_X1 U13688 ( .A(n10695), .B(n10694), .ZN(n14636) );
  OR2_X1 U13689 ( .A1(n14636), .A2(n10640), .ZN(n10696) );
  INV_X1 U13690 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15344) );
  NAND2_X1 U13691 ( .A1(n10696), .A2(n15344), .ZN(n15166) );
  INV_X1 U13692 ( .A(n10697), .ZN(n10698) );
  XNOR2_X1 U13693 ( .A(n10699), .B(n10698), .ZN(n14648) );
  NAND2_X1 U13694 ( .A1(n14648), .A2(n10962), .ZN(n10706) );
  INV_X1 U13695 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15343) );
  NAND2_X1 U13696 ( .A1(n10706), .A2(n15343), .ZN(n15175) );
  INV_X1 U13697 ( .A(n10700), .ZN(n10701) );
  XNOR2_X1 U13698 ( .A(n10702), .B(n10701), .ZN(n18900) );
  NAND2_X1 U13699 ( .A1(n18900), .A2(n10962), .ZN(n10703) );
  INV_X1 U13700 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15369) );
  NAND2_X1 U13701 ( .A1(n10703), .A2(n15369), .ZN(n15187) );
  AND2_X1 U13702 ( .A1(n15175), .A2(n15187), .ZN(n15163) );
  AND2_X1 U13703 ( .A1(n15166), .A2(n15163), .ZN(n15154) );
  NAND2_X1 U13704 ( .A1(n10962), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10705) );
  OR2_X1 U13705 ( .A1(n18892), .A2(n10705), .ZN(n15155) );
  OR2_X1 U13706 ( .A1(n10706), .A2(n15343), .ZN(n15176) );
  AND2_X1 U13707 ( .A1(n10962), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10707) );
  NAND2_X1 U13708 ( .A1(n18900), .A2(n10707), .ZN(n15186) );
  AND2_X1 U13709 ( .A1(n15176), .A2(n15186), .ZN(n15153) );
  OR3_X1 U13710 ( .A1(n13919), .A2(n10640), .A3(n15626), .ZN(n15204) );
  NAND2_X1 U13711 ( .A1(n10962), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10708) );
  OR2_X1 U13712 ( .A1(n18914), .A2(n10708), .ZN(n15202) );
  AND2_X1 U13713 ( .A1(n15204), .A2(n15202), .ZN(n15152) );
  INV_X1 U13714 ( .A(n18935), .ZN(n10710) );
  AND2_X1 U13715 ( .A1(n10962), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10709) );
  NAND2_X1 U13716 ( .A1(n10710), .A2(n10709), .ZN(n16204) );
  NAND2_X1 U13717 ( .A1(n10962), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10711) );
  OR2_X1 U13718 ( .A1(n18923), .A2(n10711), .ZN(n15380) );
  NAND2_X1 U13719 ( .A1(n16204), .A2(n15380), .ZN(n15150) );
  INV_X1 U13720 ( .A(n15150), .ZN(n10713) );
  NAND2_X1 U13721 ( .A1(n10962), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10712) );
  AND3_X1 U13722 ( .A1(n15152), .A2(n10713), .A3(n15395), .ZN(n10714) );
  AND4_X1 U13723 ( .A1(n15155), .A2(n15153), .A3(n10714), .A4(n15165), .ZN(
        n10715) );
  NAND2_X1 U13724 ( .A1(n9649), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10717) );
  NAND2_X1 U13725 ( .A1(n10718), .A2(n10069), .ZN(n10719) );
  AND2_X1 U13726 ( .A1(n10724), .A2(n10719), .ZN(n15605) );
  NAND2_X1 U13727 ( .A1(n15605), .A2(n10962), .ZN(n10720) );
  INV_X1 U13728 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15320) );
  NAND2_X1 U13729 ( .A1(n10720), .A2(n15320), .ZN(n15137) );
  INV_X1 U13730 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10903) );
  NOR2_X1 U13731 ( .A1(n13441), .A2(n10903), .ZN(n10723) );
  INV_X1 U13732 ( .A(n10723), .ZN(n10721) );
  XNOR2_X1 U13733 ( .A(n10724), .B(n10721), .ZN(n16152) );
  NAND2_X1 U13734 ( .A1(n16152), .A2(n10962), .ZN(n10722) );
  INV_X1 U13735 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15307) );
  NAND3_X1 U13736 ( .A1(n10725), .A2(n9649), .A3(P2_EBX_REG_24__SCAN_IN), .ZN(
        n10726) );
  NAND2_X1 U13737 ( .A1(n10726), .A2(n10735), .ZN(n10727) );
  NOR2_X1 U13738 ( .A1(n9718), .A2(n10727), .ZN(n16141) );
  AND2_X1 U13739 ( .A1(n16141), .A2(n10962), .ZN(n10728) );
  AND2_X1 U13740 ( .A1(n10728), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15113) );
  INV_X1 U13741 ( .A(n10728), .ZN(n10729) );
  INV_X1 U13742 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15297) );
  NAND2_X1 U13743 ( .A1(n10729), .A2(n15297), .ZN(n15111) );
  INV_X1 U13744 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n10730) );
  NOR2_X1 U13745 ( .A1(n9718), .A2(n10730), .ZN(n10731) );
  NAND2_X1 U13746 ( .A1(n9649), .A2(n10731), .ZN(n10732) );
  AND2_X1 U13747 ( .A1(n10735), .A2(n10732), .ZN(n10733) );
  NAND2_X1 U13748 ( .A1(n10736), .A2(n10733), .ZN(n16129) );
  OR2_X1 U13749 ( .A1(n16129), .A2(n10640), .ZN(n10734) );
  INV_X1 U13750 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21079) );
  NAND2_X1 U13751 ( .A1(n10734), .A2(n21079), .ZN(n15102) );
  NAND2_X1 U13752 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n10736), .ZN(n10737) );
  NOR2_X1 U13753 ( .A1(n13441), .A2(n10737), .ZN(n10738) );
  NOR2_X1 U13754 ( .A1(n11365), .A2(n10738), .ZN(n16118) );
  NAND2_X1 U13755 ( .A1(n16118), .A2(n10962), .ZN(n10739) );
  XNOR2_X1 U13756 ( .A(n10739), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11398) );
  INV_X1 U13757 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15270) );
  OR2_X1 U13758 ( .A1(n10739), .A2(n15270), .ZN(n10740) );
  NAND2_X1 U13759 ( .A1(n9649), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10743) );
  INV_X1 U13760 ( .A(n10741), .ZN(n10742) );
  OR2_X1 U13761 ( .A1(n10743), .A2(n10742), .ZN(n10744) );
  AND2_X1 U13762 ( .A1(n10957), .A2(n10744), .ZN(n16108) );
  NAND2_X1 U13763 ( .A1(n16108), .A2(n10962), .ZN(n10746) );
  XNOR2_X1 U13764 ( .A(n10745), .B(n10746), .ZN(n15098) );
  INV_X1 U13765 ( .A(n10745), .ZN(n10747) );
  INV_X1 U13766 ( .A(P2_EBX_REG_28__SCAN_IN), .ZN(n10922) );
  NOR2_X1 U13767 ( .A1(n13441), .A2(n10922), .ZN(n10956) );
  XOR2_X1 U13768 ( .A(n10956), .B(n10957), .Z(n16096) );
  NAND2_X1 U13769 ( .A1(n16096), .A2(n10962), .ZN(n10952) );
  XNOR2_X1 U13770 ( .A(n10952), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10748) );
  XNOR2_X1 U13771 ( .A(n10749), .B(n10748), .ZN(n15254) );
  INV_X1 U13772 ( .A(n10750), .ZN(n10751) );
  NAND2_X1 U13773 ( .A1(n10999), .A2(n10986), .ZN(n10760) );
  NAND2_X1 U13774 ( .A1(n15710), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n10754) );
  NOR2_X1 U13775 ( .A1(n10988), .A2(n10756), .ZN(n10768) );
  INV_X1 U13776 ( .A(n10768), .ZN(n10758) );
  NAND2_X1 U13777 ( .A1(n10758), .A2(n10757), .ZN(n10991) );
  NOR2_X1 U13778 ( .A1(n10991), .A2(n10760), .ZN(n10759) );
  OR2_X1 U13779 ( .A1(n11007), .A2(n10759), .ZN(n13465) );
  OAI211_X1 U13780 ( .C1(n10990), .C2(n10760), .A(n15457), .B(n11368), .ZN(
        n10761) );
  INV_X1 U13781 ( .A(n10761), .ZN(n10764) );
  INV_X1 U13782 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12927) );
  NAND3_X1 U13783 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10762) );
  AND2_X1 U13784 ( .A1(n12927), .A2(n10762), .ZN(n12923) );
  NAND2_X1 U13785 ( .A1(n10467), .A2(n12923), .ZN(n10763) );
  INV_X1 U13786 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n12921) );
  AOI21_X1 U13787 ( .B1(n10763), .B2(n12921), .A(n15457), .ZN(n16346) );
  NOR2_X1 U13788 ( .A1(n10764), .A2(n16346), .ZN(n19859) );
  NAND2_X1 U13789 ( .A1(n13473), .A2(n11027), .ZN(n10765) );
  INV_X1 U13790 ( .A(n10766), .ZN(n10767) );
  OAI21_X1 U13791 ( .B1(n10769), .B2(n10768), .A(n10767), .ZN(n10773) );
  INV_X1 U13792 ( .A(n10770), .ZN(n10771) );
  AOI21_X1 U13793 ( .B1(n10773), .B2(n11002), .A(n11007), .ZN(n19863) );
  NAND2_X1 U13794 ( .A1(n19231), .A2(n9677), .ZN(n11311) );
  NOR2_X1 U13795 ( .A1(n10774), .A2(n11311), .ZN(n11017) );
  NAND2_X1 U13796 ( .A1(n19863), .A2(n11017), .ZN(n10775) );
  NAND2_X1 U13797 ( .A1(n10776), .A2(n10775), .ZN(n10968) );
  AND2_X1 U13798 ( .A1(n9677), .A2(n16351), .ZN(n11367) );
  NAND2_X1 U13799 ( .A1(n9663), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13747) );
  INV_X1 U13800 ( .A(n13747), .ZN(n10778) );
  NAND2_X1 U13801 ( .A1(n10778), .A2(n10808), .ZN(n13866) );
  XOR2_X1 U13802 ( .A(n10780), .B(n10779), .Z(n14182) );
  INV_X1 U13803 ( .A(n12849), .ZN(n10781) );
  NAND2_X1 U13804 ( .A1(n10781), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12851) );
  XOR2_X1 U13805 ( .A(n10782), .B(n11081), .Z(n10783) );
  NOR2_X1 U13806 ( .A1(n12851), .A2(n10783), .ZN(n10784) );
  INV_X1 U13807 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15456) );
  XNOR2_X1 U13808 ( .A(n12851), .B(n10783), .ZN(n12862) );
  NOR2_X1 U13809 ( .A1(n15456), .A2(n12862), .ZN(n12861) );
  NOR2_X1 U13810 ( .A1(n10784), .A2(n12861), .ZN(n10786) );
  XOR2_X1 U13811 ( .A(n10786), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(
        n14181) );
  NOR2_X1 U13812 ( .A1(n14182), .A2(n14181), .ZN(n14180) );
  INV_X1 U13813 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10785) );
  NOR2_X1 U13814 ( .A1(n10786), .A2(n10785), .ZN(n10787) );
  OR2_X1 U13815 ( .A1(n14180), .A2(n10787), .ZN(n10788) );
  INV_X1 U13816 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13582) );
  XNOR2_X1 U13817 ( .A(n10788), .B(n13582), .ZN(n13590) );
  NAND2_X1 U13818 ( .A1(n10788), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10789) );
  NAND2_X1 U13819 ( .A1(n13565), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10794) );
  INV_X1 U13820 ( .A(n11095), .ZN(n10790) );
  NAND2_X1 U13821 ( .A1(n10791), .A2(n10790), .ZN(n10792) );
  NAND2_X1 U13822 ( .A1(n10793), .A2(n10792), .ZN(n13566) );
  INV_X1 U13823 ( .A(n13565), .ZN(n10795) );
  NAND2_X1 U13824 ( .A1(n10797), .A2(n10796), .ZN(n13746) );
  NAND2_X1 U13825 ( .A1(n10804), .A2(n10803), .ZN(n10801) );
  NAND2_X1 U13826 ( .A1(n10802), .A2(n13867), .ZN(n10807) );
  INV_X1 U13827 ( .A(n10805), .ZN(n10806) );
  XNOR2_X1 U13828 ( .A(n10812), .B(n10640), .ZN(n10810) );
  INV_X1 U13829 ( .A(n10812), .ZN(n10815) );
  NAND2_X1 U13830 ( .A1(n10815), .A2(n10962), .ZN(n10813) );
  NAND2_X1 U13831 ( .A1(n10815), .A2(n10814), .ZN(n10816) );
  NAND2_X1 U13832 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16283) );
  NOR2_X1 U13833 ( .A1(n10684), .A2(n16283), .ZN(n15385) );
  INV_X1 U13834 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21061) );
  INV_X1 U13835 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16300) );
  NOR2_X1 U13836 ( .A1(n10651), .A2(n16300), .ZN(n16295) );
  INV_X1 U13837 ( .A(n16295), .ZN(n15219) );
  NOR2_X1 U13838 ( .A1(n21061), .A2(n15219), .ZN(n15402) );
  AND2_X1 U13839 ( .A1(n15385), .A2(n15402), .ZN(n15386) );
  AND2_X1 U13840 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10818) );
  AND2_X1 U13841 ( .A1(n15386), .A2(n10818), .ZN(n15212) );
  AND2_X1 U13842 ( .A1(n15212), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15370) );
  INV_X1 U13843 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15258) );
  NOR2_X2 U13844 ( .A1(n11393), .A2(n15258), .ZN(n15092) );
  INV_X1 U13845 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10953) );
  XNOR2_X1 U13846 ( .A(n15092), .B(n10953), .ZN(n15252) );
  INV_X1 U13847 ( .A(n12780), .ZN(n10819) );
  NAND2_X1 U13848 ( .A1(n15252), .A2(n16269), .ZN(n10937) );
  NAND2_X1 U13849 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10824) );
  INV_X4 U13850 ( .A(n10836), .ZN(n11313) );
  INV_X2 U13851 ( .A(n10330), .ZN(n10943) );
  INV_X1 U13852 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10821) );
  INV_X1 U13853 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10820) );
  OAI22_X1 U13854 ( .A1(n10943), .A2(n10821), .B1(n15457), .B2(n10820), .ZN(
        n10822) );
  AOI21_X1 U13855 ( .B1(n11313), .B2(P2_REIP_REG_15__SCAN_IN), .A(n10822), 
        .ZN(n10823) );
  NAND2_X1 U13856 ( .A1(n10824), .A2(n10823), .ZN(n13650) );
  NAND2_X1 U13857 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10828) );
  INV_X1 U13858 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10825) );
  OAI22_X1 U13859 ( .A1(n10943), .A2(n13285), .B1(n15457), .B2(n10825), .ZN(
        n10826) );
  AOI21_X1 U13860 ( .B1(n11313), .B2(P2_REIP_REG_9__SCAN_IN), .A(n10826), .ZN(
        n10827) );
  NAND2_X1 U13861 ( .A1(n10828), .A2(n10827), .ZN(n13283) );
  INV_X1 U13862 ( .A(n10829), .ZN(n10833) );
  OAI22_X1 U13863 ( .A1(n10833), .A2(n10832), .B1(n10831), .B2(n10830), .ZN(
        n13572) );
  INV_X1 U13864 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10835) );
  AOI22_X1 U13865 ( .A1(n10330), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10834) );
  OAI21_X1 U13866 ( .B1(n10836), .B2(n10835), .A(n10834), .ZN(n10837) );
  AOI21_X1 U13867 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n10873), .A(
        n10837), .ZN(n13571) );
  NAND2_X1 U13868 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10842) );
  OAI22_X1 U13869 ( .A1(n10943), .A2(n10839), .B1(n15457), .B2(n10838), .ZN(
        n10840) );
  AOI21_X1 U13870 ( .B1(n11313), .B2(P2_REIP_REG_5__SCAN_IN), .A(n10840), .ZN(
        n10841) );
  NAND2_X1 U13871 ( .A1(n10842), .A2(n10841), .ZN(n13194) );
  NAND2_X1 U13872 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10846) );
  INV_X1 U13873 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10843) );
  OAI22_X1 U13874 ( .A1(n10943), .A2(n13315), .B1(n15457), .B2(n10843), .ZN(
        n10844) );
  AOI21_X1 U13875 ( .B1(n11313), .B2(P2_REIP_REG_6__SCAN_IN), .A(n10844), .ZN(
        n10845) );
  NAND2_X1 U13876 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10851) );
  INV_X1 U13877 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10847) );
  OAI22_X1 U13878 ( .A1(n10943), .A2(n10848), .B1(n15457), .B2(n10847), .ZN(
        n10849) );
  AOI21_X1 U13879 ( .B1(n11313), .B2(P2_REIP_REG_7__SCAN_IN), .A(n10849), .ZN(
        n10850) );
  NAND2_X1 U13880 ( .A1(n10851), .A2(n10850), .ZN(n13302) );
  NAND2_X1 U13881 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10856) );
  INV_X1 U13882 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n10853) );
  INV_X1 U13883 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10852) );
  OAI22_X1 U13884 ( .A1(n10943), .A2(n10853), .B1(n15457), .B2(n10852), .ZN(
        n10854) );
  AOI21_X1 U13885 ( .B1(n11313), .B2(P2_REIP_REG_8__SCAN_IN), .A(n10854), .ZN(
        n10855) );
  NAND2_X1 U13886 ( .A1(n13283), .A2(n16242), .ZN(n15236) );
  NAND2_X1 U13887 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10860) );
  INV_X1 U13888 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10857) );
  INV_X1 U13889 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15239) );
  OAI22_X1 U13890 ( .A1(n10943), .A2(n10857), .B1(n15457), .B2(n15239), .ZN(
        n10858) );
  AOI21_X1 U13891 ( .B1(n11313), .B2(P2_REIP_REG_10__SCAN_IN), .A(n10858), 
        .ZN(n10859) );
  NAND2_X1 U13892 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10864) );
  INV_X1 U13893 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10861) );
  OAI22_X1 U13894 ( .A1(n10943), .A2(n13410), .B1(n15457), .B2(n10861), .ZN(
        n10862) );
  AOI21_X1 U13895 ( .B1(n11313), .B2(P2_REIP_REG_11__SCAN_IN), .A(n10862), 
        .ZN(n10863) );
  NAND2_X1 U13896 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10869) );
  INV_X1 U13897 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n10866) );
  OAI22_X1 U13898 ( .A1(n10943), .A2(n10866), .B1(n15457), .B2(n10004), .ZN(
        n10867) );
  AOI21_X1 U13899 ( .B1(n11313), .B2(P2_REIP_REG_12__SCAN_IN), .A(n10867), 
        .ZN(n10868) );
  NAND2_X1 U13900 ( .A1(n10869), .A2(n10868), .ZN(n13343) );
  NAND2_X1 U13901 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10872) );
  OAI22_X1 U13902 ( .A1(n10943), .A2(n13448), .B1(n15457), .B2(n16216), .ZN(
        n10870) );
  AOI21_X1 U13903 ( .B1(n11313), .B2(P2_REIP_REG_13__SCAN_IN), .A(n10870), 
        .ZN(n10871) );
  NAND2_X1 U13904 ( .A1(n10872), .A2(n10871), .ZN(n13445) );
  INV_X1 U13905 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13559) );
  OAI22_X1 U13906 ( .A1(n10943), .A2(n13559), .B1(n15457), .B2(n10005), .ZN(
        n10875) );
  NOR2_X1 U13907 ( .A1(n9671), .A2(n10684), .ZN(n10874) );
  AOI211_X1 U13908 ( .C1(n11313), .C2(P2_REIP_REG_14__SCAN_IN), .A(n10875), 
        .B(n10874), .ZN(n13556) );
  NAND2_X1 U13909 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10880) );
  INV_X1 U13910 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10876) );
  OAI22_X1 U13911 ( .A1(n10943), .A2(n10877), .B1(n15457), .B2(n10876), .ZN(
        n10878) );
  AOI21_X1 U13912 ( .B1(n11313), .B2(P2_REIP_REG_16__SCAN_IN), .A(n10878), 
        .ZN(n10879) );
  NAND2_X1 U13913 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10883) );
  OAI22_X1 U13914 ( .A1(n10943), .A2(n13920), .B1(n15457), .B2(n10008), .ZN(
        n10881) );
  AOI21_X1 U13915 ( .B1(n11313), .B2(P2_REIP_REG_17__SCAN_IN), .A(n10881), 
        .ZN(n10882) );
  NOR2_X2 U13916 ( .A1(n15223), .A2(n13881), .ZN(n15194) );
  NAND2_X1 U13917 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10886) );
  INV_X1 U13918 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10930) );
  OAI22_X1 U13919 ( .A1(n10943), .A2(n16181), .B1(n15457), .B2(n10930), .ZN(
        n10884) );
  AOI21_X1 U13920 ( .B1(n11313), .B2(P2_REIP_REG_18__SCAN_IN), .A(n10884), 
        .ZN(n10885) );
  NAND2_X1 U13921 ( .A1(n10886), .A2(n10885), .ZN(n15193) );
  NAND2_X1 U13922 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10890) );
  INV_X1 U13923 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n11339) );
  OAI22_X1 U13924 ( .A1(n10943), .A2(n10887), .B1(n15457), .B2(n11339), .ZN(
        n10888) );
  AOI21_X1 U13925 ( .B1(n11313), .B2(P2_REIP_REG_19__SCAN_IN), .A(n10888), 
        .ZN(n10889) );
  NAND2_X1 U13926 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10893) );
  OAI22_X1 U13927 ( .A1(n10943), .A2(n16177), .B1(n15457), .B2(n10009), .ZN(
        n10891) );
  AOI21_X1 U13928 ( .B1(n11313), .B2(P2_REIP_REG_20__SCAN_IN), .A(n10891), 
        .ZN(n10892) );
  NAND2_X1 U13929 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10897) );
  INV_X1 U13930 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10894) );
  INV_X1 U13931 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18890) );
  OAI22_X1 U13932 ( .A1(n10943), .A2(n10894), .B1(n15457), .B2(n18890), .ZN(
        n10895) );
  AOI21_X1 U13933 ( .B1(n11313), .B2(P2_REIP_REG_21__SCAN_IN), .A(n10895), 
        .ZN(n10896) );
  NAND2_X1 U13934 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10902) );
  INV_X1 U13935 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n10899) );
  INV_X1 U13936 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10898) );
  OAI22_X1 U13937 ( .A1(n10943), .A2(n10899), .B1(n15457), .B2(n10898), .ZN(
        n10900) );
  AOI21_X1 U13938 ( .B1(n11313), .B2(P2_REIP_REG_22__SCAN_IN), .A(n10900), 
        .ZN(n10901) );
  NAND2_X1 U13939 ( .A1(n10902), .A2(n10901), .ZN(n15140) );
  NAND2_X1 U13940 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10906) );
  INV_X1 U13941 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15128) );
  OAI22_X1 U13942 ( .A1(n10943), .A2(n10903), .B1(n15457), .B2(n15128), .ZN(
        n10904) );
  AOI21_X1 U13943 ( .B1(n11313), .B2(P2_REIP_REG_23__SCAN_IN), .A(n10904), 
        .ZN(n10905) );
  NAND2_X1 U13944 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10910) );
  INV_X1 U13945 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n10907) );
  OAI22_X1 U13946 ( .A1(n10943), .A2(n10907), .B1(n15457), .B2(n10012), .ZN(
        n10908) );
  AOI21_X1 U13947 ( .B1(n11313), .B2(P2_REIP_REG_24__SCAN_IN), .A(n10908), 
        .ZN(n10909) );
  NAND2_X1 U13948 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10913) );
  INV_X1 U13949 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15105) );
  OAI22_X1 U13950 ( .A1(n10943), .A2(n10730), .B1(n15457), .B2(n15105), .ZN(
        n10911) );
  AOI21_X1 U13951 ( .B1(n11313), .B2(P2_REIP_REG_25__SCAN_IN), .A(n10911), 
        .ZN(n10912) );
  NAND2_X1 U13952 ( .A1(n10913), .A2(n10912), .ZN(n14969) );
  NAND2_X1 U13953 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10916) );
  INV_X1 U13954 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n21077) );
  INV_X1 U13955 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11328) );
  OAI22_X1 U13956 ( .A1(n10943), .A2(n21077), .B1(n15457), .B2(n11328), .ZN(
        n10914) );
  AOI21_X1 U13957 ( .B1(n11313), .B2(P2_REIP_REG_26__SCAN_IN), .A(n10914), 
        .ZN(n10915) );
  AND2_X1 U13958 ( .A1(n10916), .A2(n10915), .ZN(n11402) );
  NAND2_X1 U13959 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10920) );
  INV_X1 U13960 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n10917) );
  INV_X1 U13961 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n20923) );
  OAI22_X1 U13962 ( .A1(n10943), .A2(n10917), .B1(n15457), .B2(n20923), .ZN(
        n10918) );
  AOI21_X1 U13963 ( .B1(n11313), .B2(P2_REIP_REG_27__SCAN_IN), .A(n10918), 
        .ZN(n10919) );
  NAND2_X1 U13964 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10925) );
  INV_X1 U13965 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10921) );
  OAI22_X1 U13966 ( .A1(n10943), .A2(n10922), .B1(n15457), .B2(n10921), .ZN(
        n10923) );
  AOI21_X1 U13967 ( .B1(n11313), .B2(P2_REIP_REG_28__SCAN_IN), .A(n10923), 
        .ZN(n10924) );
  NAND2_X1 U13968 ( .A1(n10925), .A2(n10924), .ZN(n10926) );
  NOR2_X1 U13969 ( .A1(n14953), .A2(n10926), .ZN(n10927) );
  NAND2_X1 U13970 ( .A1(n15457), .A2(n19825), .ZN(n19820) );
  INV_X1 U13971 ( .A(n19820), .ZN(n15463) );
  OR2_X1 U13972 ( .A1(n19830), .A2(n15463), .ZN(n19847) );
  INV_X1 U13973 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n16342) );
  NAND2_X1 U13974 ( .A1(n19847), .A2(n16342), .ZN(n10928) );
  AND2_X1 U13975 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19838) );
  NAND2_X1 U13976 ( .A1(n19830), .A2(n15457), .ZN(n18862) );
  OR2_X2 U13977 ( .A1(n18862), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19046) );
  INV_X1 U13978 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n11294) );
  NOR2_X1 U13979 ( .A1(n19046), .A2(n11294), .ZN(n15244) );
  NAND2_X1 U13980 ( .A1(n16342), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13049) );
  INV_X1 U13981 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19818) );
  NAND2_X1 U13982 ( .A1(n19818), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10929) );
  NAND2_X1 U13983 ( .A1(n13049), .A2(n10929), .ZN(n12855) );
  AND2_X2 U13984 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n10931), .ZN(
        n11338) );
  NOR2_X4 U13985 ( .A1(n11337), .A2(n15128), .ZN(n11336) );
  AND2_X2 U13986 ( .A1(n11327), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11324) );
  NOR2_X1 U13987 ( .A1(n11327), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10932) );
  OR2_X1 U13988 ( .A1(n11324), .A2(n10932), .ZN(n16103) );
  NOR2_X1 U13989 ( .A1(n19229), .A2(n16103), .ZN(n10933) );
  AOI211_X1 U13990 ( .C1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n19218), .A(
        n15244), .B(n10933), .ZN(n10934) );
  OAI21_X1 U13991 ( .B1(n16098), .B2(n16273), .A(n10934), .ZN(n10935) );
  INV_X1 U13992 ( .A(n10935), .ZN(n10936) );
  OAI211_X1 U13993 ( .C1(n15254), .C2(n19221), .A(n10937), .B(n10936), .ZN(
        P2_U2986) );
  NAND2_X1 U13994 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15247) );
  INV_X1 U13995 ( .A(n15247), .ZN(n10938) );
  NAND2_X1 U13996 ( .A1(n10938), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14133) );
  XNOR2_X1 U13997 ( .A(n11410), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11018) );
  NOR2_X1 U13998 ( .A1(n11018), .A2(n19219), .ZN(n10951) );
  NAND2_X1 U13999 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10941) );
  INV_X1 U14000 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n10955) );
  INV_X1 U14001 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11430) );
  OAI22_X1 U14002 ( .A1(n10943), .A2(n10955), .B1(n15457), .B2(n11430), .ZN(
        n10939) );
  AOI21_X1 U14003 ( .B1(n11313), .B2(P2_REIP_REG_29__SCAN_IN), .A(n10939), 
        .ZN(n10940) );
  NAND2_X1 U14004 ( .A1(n10941), .A2(n10940), .ZN(n11415) );
  NAND2_X1 U14005 ( .A1(n10873), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10946) );
  INV_X1 U14006 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n10960) );
  INV_X1 U14007 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10942) );
  OAI22_X1 U14008 ( .A1(n10943), .A2(n10960), .B1(n15457), .B2(n10942), .ZN(
        n10944) );
  AOI21_X1 U14009 ( .B1(n11313), .B2(P2_REIP_REG_30__SCAN_IN), .A(n10944), 
        .ZN(n10945) );
  AND2_X1 U14010 ( .A1(n10946), .A2(n10945), .ZN(n11312) );
  AND2_X2 U14011 ( .A1(n11324), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11325) );
  XNOR2_X1 U14012 ( .A(n11325), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14619) );
  INV_X2 U14013 ( .A(n19046), .ZN(n19217) );
  NAND2_X1 U14014 ( .A1(n19217), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11061) );
  NAND2_X1 U14015 ( .A1(n19218), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10947) );
  OAI211_X1 U14016 ( .C1(n19229), .C2(n14619), .A(n11061), .B(n10947), .ZN(
        n10948) );
  INV_X1 U14017 ( .A(n10948), .ZN(n10949) );
  OAI21_X1 U14018 ( .B1(n14938), .B2(n16273), .A(n10949), .ZN(n10950) );
  NAND2_X1 U14019 ( .A1(n10952), .A2(n15247), .ZN(n10954) );
  NAND2_X1 U14020 ( .A1(n15258), .A2(n10953), .ZN(n15246) );
  NOR2_X1 U14021 ( .A1(n13441), .A2(n10955), .ZN(n10958) );
  XOR2_X1 U14022 ( .A(n10958), .B(n10959), .Z(n16085) );
  AOI21_X1 U14023 ( .B1(n16085), .B2(n10962), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11424) );
  NOR2_X1 U14024 ( .A1(n13441), .A2(n10960), .ZN(n10961) );
  XNOR2_X1 U14025 ( .A(n11362), .B(n10961), .ZN(n14621) );
  NAND2_X1 U14026 ( .A1(n10962), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10963) );
  NOR2_X1 U14027 ( .A1(n14621), .A2(n10963), .ZN(n11382) );
  INV_X1 U14028 ( .A(n11382), .ZN(n10964) );
  INV_X1 U14029 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14134) );
  OAI21_X1 U14030 ( .B1(n14621), .B2(n10640), .A(n14134), .ZN(n11383) );
  NAND2_X1 U14031 ( .A1(n10964), .A2(n11383), .ZN(n10965) );
  NAND2_X1 U14032 ( .A1(n10967), .A2(n10966), .ZN(P2_U2984) );
  INV_X1 U14033 ( .A(n10968), .ZN(n11015) );
  NAND2_X1 U14034 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n16355) );
  INV_X1 U14035 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n18859) );
  NOR2_X1 U14036 ( .A1(n18859), .A2(n19752), .ZN(n19744) );
  NOR2_X1 U14037 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19745) );
  NOR3_X1 U14038 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19744), .A3(n19745), 
        .ZN(n19737) );
  NAND2_X1 U14039 ( .A1(n16355), .A2(n19737), .ZN(n12911) );
  INV_X1 U14040 ( .A(n12911), .ZN(n12778) );
  NAND3_X1 U14041 ( .A1(n10969), .A2(n11368), .A3(n12778), .ZN(n10978) );
  OR2_X1 U14042 ( .A1(n12924), .A2(n9678), .ZN(n12912) );
  NAND2_X1 U14043 ( .A1(n10269), .A2(n19244), .ZN(n10970) );
  NAND2_X1 U14044 ( .A1(n10970), .A2(n11041), .ZN(n10973) );
  NAND2_X1 U14045 ( .A1(n19231), .A2(n19244), .ZN(n11023) );
  NAND2_X1 U14046 ( .A1(n11023), .A2(n10273), .ZN(n10971) );
  AOI21_X1 U14047 ( .B1(n12912), .B2(n10973), .A(n10972), .ZN(n11025) );
  NAND2_X1 U14048 ( .A1(n10976), .A2(n19257), .ZN(n10975) );
  INV_X1 U14049 ( .A(n11311), .ZN(n10974) );
  NAND2_X1 U14050 ( .A1(n10975), .A2(n10974), .ZN(n11030) );
  NAND2_X1 U14051 ( .A1(n10270), .A2(n10271), .ZN(n10977) );
  NAND4_X1 U14052 ( .A1(n10978), .A2(n11025), .A3(n11030), .A4(n10977), .ZN(
        n12918) );
  MUX2_X1 U14053 ( .A(n10979), .B(n11041), .S(n19231), .Z(n10981) );
  NAND2_X1 U14054 ( .A1(n11368), .A2(n16355), .ZN(n10980) );
  NOR2_X1 U14055 ( .A1(n10981), .A2(n10980), .ZN(n10982) );
  NOR2_X1 U14056 ( .A1(n12918), .A2(n10982), .ZN(n11014) );
  NAND2_X1 U14057 ( .A1(n9677), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11006) );
  NAND2_X1 U14058 ( .A1(n11027), .A2(n11006), .ZN(n10985) );
  MUX2_X1 U14059 ( .A(n10985), .B(n10984), .S(n10986), .Z(n10998) );
  NAND2_X1 U14060 ( .A1(n13474), .A2(n10986), .ZN(n10996) );
  INV_X1 U14061 ( .A(n10990), .ZN(n10987) );
  NAND2_X1 U14062 ( .A1(n10988), .A2(n10987), .ZN(n10989) );
  NAND2_X1 U14063 ( .A1(n10983), .A2(n10989), .ZN(n10995) );
  NAND2_X1 U14064 ( .A1(n19231), .A2(n10990), .ZN(n10993) );
  INV_X1 U14065 ( .A(n10991), .ZN(n10992) );
  NAND3_X1 U14066 ( .A1(n10993), .A2(n10273), .A3(n10992), .ZN(n10994) );
  NAND3_X1 U14067 ( .A1(n10996), .A2(n10995), .A3(n10994), .ZN(n10997) );
  NAND2_X1 U14068 ( .A1(n10998), .A2(n10997), .ZN(n11000) );
  NAND2_X1 U14069 ( .A1(n11000), .A2(n10999), .ZN(n11001) );
  INV_X1 U14070 ( .A(n11007), .ZN(n11003) );
  NAND2_X1 U14071 ( .A1(n11004), .A2(n11003), .ZN(n11005) );
  MUX2_X1 U14072 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n11005), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n11009) );
  NAND2_X1 U14073 ( .A1(n11007), .A2(n12872), .ZN(n11008) );
  AND2_X1 U14074 ( .A1(n13467), .A2(n11027), .ZN(n12914) );
  INV_X1 U14075 ( .A(n12914), .ZN(n11011) );
  AOI21_X1 U14076 ( .B1(n11009), .B2(n10273), .A(n10271), .ZN(n11010) );
  NAND2_X1 U14077 ( .A1(n11011), .A2(n11010), .ZN(n11013) );
  NAND3_X1 U14078 ( .A1(n12914), .A2(n13434), .A3(n12778), .ZN(n11012) );
  NAND4_X1 U14079 ( .A1(n11015), .A2(n11014), .A3(n11013), .A4(n11012), .ZN(
        n11016) );
  INV_X1 U14080 ( .A(n11017), .ZN(n19862) );
  NAND2_X1 U14081 ( .A1(n13473), .A2(n10983), .ZN(n19857) );
  OAI21_X1 U14082 ( .B1(n10979), .B2(n10273), .A(n12912), .ZN(n13464) );
  NOR2_X1 U14083 ( .A1(n11019), .A2(n10265), .ZN(n11020) );
  OR2_X1 U14084 ( .A1(n13464), .A2(n11020), .ZN(n13485) );
  AOI21_X1 U14085 ( .B1(n13485), .B2(n19231), .A(n11021), .ZN(n11022) );
  NAND3_X1 U14086 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13900) );
  NOR2_X1 U14087 ( .A1(n13901), .A2(n13900), .ZN(n13872) );
  NAND3_X1 U14088 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(n13872), .ZN(n11047) );
  INV_X1 U14089 ( .A(n11023), .ZN(n11024) );
  NAND3_X1 U14090 ( .A1(n11025), .A2(n11024), .A3(n11030), .ZN(n13295) );
  NAND2_X1 U14091 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14193) );
  INV_X1 U14092 ( .A(n14193), .ZN(n14189) );
  NAND2_X1 U14093 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14189), .ZN(
        n11026) );
  NOR2_X1 U14094 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14189), .ZN(
        n13568) );
  AOI21_X1 U14095 ( .B1(n14192), .B2(n11026), .A(n13568), .ZN(n13588) );
  NAND2_X1 U14096 ( .A1(n11028), .A2(n11027), .ZN(n13479) );
  AOI21_X1 U14097 ( .B1(n13479), .B2(n11030), .A(n11029), .ZN(n11038) );
  MUX2_X1 U14098 ( .A(n11031), .B(n11041), .S(n9678), .Z(n11036) );
  INV_X1 U14099 ( .A(n11032), .ZN(n12786) );
  OAI21_X1 U14100 ( .B1(n11033), .B2(n19244), .A(n12786), .ZN(n11035) );
  NAND2_X1 U14101 ( .A1(n11034), .A2(n9723), .ZN(n12968) );
  NAND3_X1 U14102 ( .A1(n11036), .A2(n11035), .A3(n12968), .ZN(n11037) );
  NOR2_X1 U14103 ( .A1(n11038), .A2(n11037), .ZN(n13003) );
  NAND3_X1 U14104 ( .A1(n9660), .A2(n11041), .A3(n11040), .ZN(n11042) );
  NAND2_X1 U14105 ( .A1(n13003), .A2(n11042), .ZN(n13488) );
  INV_X1 U14106 ( .A(n9659), .ZN(n13002) );
  NOR2_X1 U14107 ( .A1(n13488), .A2(n13002), .ZN(n11044) );
  NAND2_X1 U14108 ( .A1(n13588), .A2(n16334), .ZN(n13899) );
  AND2_X1 U14109 ( .A1(n15370), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15340) );
  NAND2_X1 U14110 ( .A1(n15444), .A2(n15340), .ZN(n15356) );
  NOR2_X1 U14111 ( .A1(n15343), .A2(n15344), .ZN(n15342) );
  NAND2_X1 U14112 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15342), .ZN(
        n11045) );
  NOR2_X1 U14113 ( .A1(n15320), .A2(n15307), .ZN(n15305) );
  NAND2_X1 U14114 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15305), .ZN(
        n11046) );
  NOR2_X1 U14115 ( .A1(n15296), .A2(n11046), .ZN(n15279) );
  AND2_X1 U14116 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11056) );
  NAND2_X1 U14117 ( .A1(n15279), .A2(n11056), .ZN(n15255) );
  OAI21_X1 U14118 ( .B1(n15255), .B2(n14133), .A(n14134), .ZN(n11060) );
  INV_X1 U14119 ( .A(n16334), .ZN(n15401) );
  AND2_X1 U14120 ( .A1(n11304), .A2(n19046), .ZN(n12991) );
  INV_X1 U14121 ( .A(n12991), .ZN(n16331) );
  NAND2_X1 U14122 ( .A1(n15401), .A2(n16331), .ZN(n15426) );
  INV_X1 U14123 ( .A(n13568), .ZN(n11049) );
  INV_X1 U14124 ( .A(n11047), .ZN(n11048) );
  NAND2_X1 U14125 ( .A1(n11049), .A2(n11048), .ZN(n11050) );
  NAND2_X1 U14126 ( .A1(n16334), .A2(n11050), .ZN(n11052) );
  AOI21_X1 U14127 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n14189), .A(
        n15598), .ZN(n11051) );
  NOR2_X1 U14128 ( .A1(n12991), .A2(n11051), .ZN(n13569) );
  NAND4_X1 U14129 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15400), .A3(
        n15340), .A4(n15342), .ZN(n15306) );
  INV_X1 U14130 ( .A(n15306), .ZN(n11053) );
  NAND2_X1 U14131 ( .A1(n11053), .A2(n15305), .ZN(n11054) );
  NAND2_X1 U14132 ( .A1(n15426), .A2(n11054), .ZN(n15292) );
  NAND2_X1 U14133 ( .A1(n16334), .A2(n15297), .ZN(n11055) );
  AND2_X1 U14134 ( .A1(n15292), .A2(n11055), .ZN(n15284) );
  INV_X1 U14135 ( .A(n11056), .ZN(n11057) );
  NAND2_X1 U14136 ( .A1(n16334), .A2(n11057), .ZN(n11058) );
  AOI21_X1 U14137 ( .B1(n16334), .B2(n14133), .A(n14134), .ZN(n11059) );
  NAND2_X1 U14138 ( .A1(n15259), .A2(n11059), .ZN(n14135) );
  NAND2_X1 U14139 ( .A1(n11060), .A2(n14135), .ZN(n11062) );
  OAI211_X1 U14140 ( .C1(n14938), .C2(n16327), .A(n11062), .B(n11061), .ZN(
        n11063) );
  INV_X2 U14141 ( .A(n9750), .ZN(n11308) );
  AOI22_X1 U14142 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n11066) );
  NAND2_X1 U14143 ( .A1(n9785), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n11065) );
  AND2_X1 U14144 ( .A1(n11066), .A2(n11065), .ZN(n11298) );
  NAND2_X1 U14145 ( .A1(n9785), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n11070) );
  INV_X1 U14146 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16335) );
  NAND2_X1 U14147 ( .A1(n12986), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n11067) );
  OAI211_X1 U14148 ( .C1(n19231), .C2(n16335), .A(n11067), .B(n19825), .ZN(
        n11068) );
  INV_X1 U14149 ( .A(n11068), .ZN(n11069) );
  NAND2_X1 U14150 ( .A1(n11070), .A2(n11069), .ZN(n12981) );
  NAND2_X1 U14151 ( .A1(n11075), .A2(n12985), .ZN(n11085) );
  INV_X1 U14152 ( .A(n11078), .ZN(n11072) );
  OAI21_X1 U14153 ( .B1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19825), .A(
        n11072), .ZN(n11073) );
  INV_X1 U14154 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19212) );
  NAND2_X1 U14155 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11077) );
  INV_X1 U14156 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19753) );
  NAND2_X1 U14157 ( .A1(n9785), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11076) );
  OAI211_X1 U14158 ( .C1(n9750), .C2(n19212), .A(n11077), .B(n11076), .ZN(
        n11082) );
  NAND2_X1 U14159 ( .A1(n10269), .A2(n11078), .ZN(n11080) );
  NAND2_X1 U14160 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11079) );
  OAI211_X1 U14161 ( .C1(n11242), .C2(n11081), .A(n11080), .B(n11079), .ZN(
        n12989) );
  NAND2_X1 U14162 ( .A1(n11265), .A2(n11083), .ZN(n11084) );
  OAI211_X1 U14163 ( .C1(n19825), .C2(n19837), .A(n11085), .B(n11084), .ZN(
        n11088) );
  INV_X1 U14164 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19209) );
  NAND2_X1 U14165 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11087) );
  NAND2_X1 U14166 ( .A1(n9785), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n11086) );
  OAI211_X1 U14167 ( .C1(n9750), .C2(n19209), .A(n11087), .B(n11086), .ZN(
        n13520) );
  NOR2_X1 U14168 ( .A1(n13521), .A2(n13520), .ZN(n13522) );
  NOR2_X1 U14169 ( .A1(n11089), .A2(n11088), .ZN(n11090) );
  AOI22_X1 U14170 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n11094) );
  AOI22_X1 U14171 ( .A1(n11265), .A2(n11091), .B1(n11308), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n11093) );
  NAND2_X1 U14172 ( .A1(n9785), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n11092) );
  NAND3_X1 U14173 ( .A1(n11094), .A2(n11093), .A3(n11092), .ZN(n13516) );
  AOI22_X1 U14174 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n11098) );
  NAND2_X1 U14175 ( .A1(n9785), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n11097) );
  NAND2_X1 U14176 ( .A1(n11265), .A2(n11095), .ZN(n11096) );
  AOI22_X1 U14177 ( .A1(n9785), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n11265), .B2(
        n11099), .ZN(n11101) );
  AOI22_X1 U14178 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n11100) );
  NAND2_X1 U14179 ( .A1(n11101), .A2(n11100), .ZN(n13753) );
  NAND2_X1 U14180 ( .A1(n11265), .A2(n11102), .ZN(n11103) );
  INV_X1 U14181 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19203) );
  NAND2_X1 U14182 ( .A1(n9785), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n11105) );
  NAND2_X1 U14183 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11104) );
  OAI211_X1 U14184 ( .C1(n9750), .C2(n19203), .A(n11105), .B(n11104), .ZN(
        n13869) );
  NAND2_X1 U14185 ( .A1(n13870), .A2(n13869), .ZN(n11107) );
  NAND2_X1 U14186 ( .A1(n11265), .A2(n10962), .ZN(n11106) );
  INV_X1 U14187 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19201) );
  NAND2_X1 U14188 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11109) );
  NAND2_X1 U14189 ( .A1(n9785), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n11108) );
  OAI211_X1 U14190 ( .C1(n9750), .C2(n19201), .A(n11109), .B(n11108), .ZN(
        n13904) );
  AOI22_X1 U14191 ( .A1(n14783), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11113) );
  NAND2_X1 U14192 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11112) );
  NAND2_X1 U14193 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11111) );
  NAND2_X1 U14194 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11110) );
  NAND4_X1 U14195 ( .A1(n11113), .A2(n11112), .A3(n11111), .A4(n11110), .ZN(
        n11116) );
  INV_X1 U14196 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13846) );
  INV_X1 U14197 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13854) );
  OAI22_X1 U14198 ( .A1(n10464), .A2(n13846), .B1(n11114), .B2(n13854), .ZN(
        n11115) );
  NOR2_X1 U14199 ( .A1(n11116), .A2(n11115), .ZN(n11127) );
  NAND2_X1 U14200 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11117) );
  OAI21_X1 U14201 ( .B1(n10472), .B2(n13851), .A(n11117), .ZN(n11120) );
  INV_X1 U14202 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13852) );
  OAI22_X1 U14203 ( .A1(n10463), .A2(n13852), .B1(n10473), .B2(n11118), .ZN(
        n11119) );
  NOR2_X1 U14204 ( .A1(n11120), .A2(n11119), .ZN(n11126) );
  AOI22_X1 U14205 ( .A1(n14767), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11121) );
  OAI21_X1 U14206 ( .B1(n10467), .B2(n11122), .A(n11121), .ZN(n11123) );
  INV_X1 U14207 ( .A(n11123), .ZN(n11125) );
  AOI22_X1 U14208 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14771), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11124) );
  NAND4_X1 U14209 ( .A1(n11127), .A2(n11126), .A3(n11125), .A4(n11124), .ZN(
        n19093) );
  INV_X1 U14210 ( .A(n19093), .ZN(n11129) );
  AOI22_X1 U14211 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n11128) );
  OAI21_X1 U14212 ( .B1(n11129), .B2(n11242), .A(n11128), .ZN(n11130) );
  AOI21_X1 U14213 ( .B1(n9785), .B2(P2_REIP_REG_8__SCAN_IN), .A(n11130), .ZN(
        n16311) );
  AOI22_X1 U14214 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11134) );
  NAND2_X1 U14215 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11133) );
  NAND2_X1 U14216 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11132) );
  NAND2_X1 U14217 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11131) );
  NAND4_X1 U14218 ( .A1(n11134), .A2(n11133), .A3(n11132), .A4(n11131), .ZN(
        n11136) );
  OAI22_X1 U14219 ( .A1(n19236), .A2(n10464), .B1(n10463), .B2(n13829), .ZN(
        n11135) );
  NOR2_X1 U14220 ( .A1(n11136), .A2(n11135), .ZN(n11146) );
  AOI22_X1 U14221 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11137) );
  OAI21_X1 U14222 ( .B1(n11138), .B2(n10467), .A(n11137), .ZN(n11139) );
  INV_X1 U14223 ( .A(n11139), .ZN(n11145) );
  OAI22_X1 U14224 ( .A1(n10472), .A2(n13828), .B1(n14738), .B2(n19562), .ZN(
        n11142) );
  INV_X1 U14225 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13830) );
  OAI22_X1 U14226 ( .A1(n11140), .A2(n10473), .B1(n11114), .B2(n13830), .ZN(
        n11141) );
  NOR2_X1 U14227 ( .A1(n11142), .A2(n11141), .ZN(n11144) );
  AOI22_X1 U14228 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10447), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11143) );
  NAND4_X1 U14229 ( .A1(n11146), .A2(n11145), .A3(n11144), .A4(n11143), .ZN(
        n19086) );
  AOI22_X1 U14230 ( .A1(n9785), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n11265), .B2(
        n19086), .ZN(n11148) );
  AOI22_X1 U14231 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n11147) );
  NAND2_X1 U14232 ( .A1(n11148), .A2(n11147), .ZN(n15441) );
  AOI22_X1 U14233 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11152) );
  NAND2_X1 U14234 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11151) );
  NAND2_X1 U14235 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11150) );
  NAND2_X1 U14236 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n11149) );
  NAND4_X1 U14237 ( .A1(n11152), .A2(n11151), .A3(n11150), .A4(n11149), .ZN(
        n11155) );
  OAI22_X1 U14238 ( .A1(n19239), .A2(n10464), .B1(n10473), .B2(n11153), .ZN(
        n11154) );
  NOR2_X1 U14239 ( .A1(n11155), .A2(n11154), .ZN(n11164) );
  AOI22_X1 U14240 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11156) );
  OAI21_X1 U14241 ( .B1(n10467), .B2(n11157), .A(n11156), .ZN(n11158) );
  INV_X1 U14242 ( .A(n11158), .ZN(n11163) );
  OAI22_X1 U14243 ( .A1(n10472), .A2(n14014), .B1(n14738), .B2(n13437), .ZN(
        n11160) );
  INV_X1 U14244 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14015) );
  INV_X1 U14245 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14016) );
  OAI22_X1 U14246 ( .A1(n14015), .A2(n10463), .B1(n11114), .B2(n14016), .ZN(
        n11159) );
  NOR2_X1 U14247 ( .A1(n11160), .A2(n11159), .ZN(n11162) );
  AOI22_X1 U14248 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n10447), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11161) );
  NAND4_X1 U14249 ( .A1(n11164), .A2(n11163), .A3(n11162), .A4(n11161), .ZN(
        n19085) );
  INV_X1 U14250 ( .A(n19085), .ZN(n11166) );
  AOI22_X1 U14251 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n11165) );
  OAI21_X1 U14252 ( .B1(n11166), .B2(n11242), .A(n11165), .ZN(n11167) );
  AOI21_X1 U14253 ( .B1(n9785), .B2(P2_REIP_REG_10__SCAN_IN), .A(n11167), .ZN(
        n15425) );
  NOR2_X2 U14254 ( .A1(n15440), .A2(n15425), .ZN(n16298) );
  AOI22_X1 U14255 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11171) );
  NAND2_X1 U14256 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11170) );
  NAND2_X1 U14257 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11169) );
  NAND2_X1 U14258 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n11168) );
  NAND4_X1 U14259 ( .A1(n11171), .A2(n11170), .A3(n11169), .A4(n11168), .ZN(
        n11173) );
  OAI22_X1 U14260 ( .A1(n19243), .A2(n10464), .B1(n10463), .B2(n14038), .ZN(
        n11172) );
  NOR2_X1 U14261 ( .A1(n11173), .A2(n11172), .ZN(n11184) );
  AOI22_X1 U14262 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11174) );
  OAI21_X1 U14263 ( .B1(n10467), .B2(n11175), .A(n11174), .ZN(n11176) );
  INV_X1 U14264 ( .A(n11176), .ZN(n11183) );
  OAI22_X1 U14265 ( .A1(n10472), .A2(n14037), .B1(n14738), .B2(n11177), .ZN(
        n11180) );
  OAI22_X1 U14266 ( .A1(n11178), .A2(n10473), .B1(n11114), .B2(n14039), .ZN(
        n11179) );
  NOR2_X1 U14267 ( .A1(n11180), .A2(n11179), .ZN(n11182) );
  AOI22_X1 U14268 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10447), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11181) );
  NAND4_X1 U14269 ( .A1(n11184), .A2(n11183), .A3(n11182), .A4(n11181), .ZN(
        n13405) );
  AOI22_X1 U14270 ( .A1(n9785), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n11265), 
        .B2(n13405), .ZN(n11186) );
  AOI22_X1 U14271 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n11185) );
  NAND2_X1 U14272 ( .A1(n11186), .A2(n11185), .ZN(n16297) );
  NAND2_X1 U14273 ( .A1(n16298), .A2(n16297), .ZN(n16296) );
  AOI22_X1 U14274 ( .A1(n11236), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11193) );
  INV_X1 U14275 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14695) );
  AOI22_X1 U14276 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11187) );
  OAI21_X1 U14277 ( .B1(n14695), .B2(n10472), .A(n11187), .ZN(n11188) );
  INV_X1 U14278 ( .A(n11188), .ZN(n11192) );
  AOI22_X1 U14279 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n14771), .B1(
        n10447), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11191) );
  INV_X1 U14280 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14697) );
  OAI22_X1 U14281 ( .A1(n19248), .A2(n10464), .B1(n11114), .B2(n14697), .ZN(
        n11189) );
  INV_X1 U14282 ( .A(n11189), .ZN(n11190) );
  NAND4_X1 U14283 ( .A1(n11193), .A2(n11192), .A3(n11191), .A4(n11190), .ZN(
        n11201) );
  INV_X1 U14284 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11194) );
  INV_X1 U14285 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14696) );
  OAI22_X1 U14286 ( .A1(n11194), .A2(n10473), .B1(n10463), .B2(n14696), .ZN(
        n11195) );
  INV_X1 U14287 ( .A(n11195), .ZN(n11199) );
  AOI22_X1 U14288 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n14782), .ZN(n11198) );
  AOI22_X1 U14289 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11197) );
  NAND2_X1 U14290 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11196) );
  NAND4_X1 U14291 ( .A1(n11199), .A2(n11198), .A3(n11197), .A4(n11196), .ZN(
        n11200) );
  INV_X1 U14292 ( .A(n13346), .ZN(n11203) );
  AOI22_X1 U14293 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n11202) );
  OAI21_X1 U14294 ( .B1(n11203), .B2(n11242), .A(n11202), .ZN(n11204) );
  AOI21_X1 U14295 ( .B1(n9785), .B2(P2_REIP_REG_12__SCAN_IN), .A(n11204), .ZN(
        n15411) );
  AOI22_X1 U14296 ( .A1(n9785), .A2(P2_REIP_REG_13__SCAN_IN), .B1(n11308), 
        .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n11222) );
  AOI22_X1 U14297 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11208) );
  NAND2_X1 U14298 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11207) );
  NAND2_X1 U14299 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11206) );
  NAND2_X1 U14300 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11205) );
  NAND4_X1 U14301 ( .A1(n11208), .A2(n11207), .A3(n11206), .A4(n11205), .ZN(
        n11210) );
  INV_X1 U14302 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n21045) );
  OAI22_X1 U14303 ( .A1(n21045), .A2(n10464), .B1(n10463), .B2(n14716), .ZN(
        n11209) );
  NOR2_X1 U14304 ( .A1(n11210), .A2(n11209), .ZN(n11220) );
  AOI22_X1 U14305 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11211) );
  OAI21_X1 U14306 ( .B1(n10467), .B2(n11212), .A(n11211), .ZN(n11213) );
  INV_X1 U14307 ( .A(n11213), .ZN(n11219) );
  OAI22_X1 U14308 ( .A1(n10472), .A2(n14715), .B1(n14738), .B2(n13444), .ZN(
        n11216) );
  OAI22_X1 U14309 ( .A1(n11214), .A2(n10473), .B1(n11114), .B2(n14717), .ZN(
        n11215) );
  NOR2_X1 U14310 ( .A1(n11216), .A2(n11215), .ZN(n11218) );
  AOI22_X1 U14311 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10447), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11217) );
  NAND4_X1 U14312 ( .A1(n11220), .A2(n11219), .A3(n11218), .A4(n11217), .ZN(
        n13550) );
  AOI22_X1 U14313 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n11075), .B1(
        n11265), .B2(n13550), .ZN(n11221) );
  NAND2_X1 U14314 ( .A1(n11222), .A2(n11221), .ZN(n15398) );
  NAND2_X1 U14315 ( .A1(n15399), .A2(n15398), .ZN(n16281) );
  AOI22_X1 U14316 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11226) );
  NAND2_X1 U14317 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11225) );
  NAND2_X1 U14318 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11224) );
  NAND2_X1 U14319 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11223) );
  NAND4_X1 U14320 ( .A1(n11226), .A2(n11225), .A3(n11224), .A4(n11223), .ZN(
        n11229) );
  OAI22_X1 U14321 ( .A1(n19255), .A2(n10464), .B1(n10473), .B2(n11227), .ZN(
        n11228) );
  NOR2_X1 U14322 ( .A1(n11229), .A2(n11228), .ZN(n11240) );
  NAND2_X1 U14323 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11230) );
  OAI21_X1 U14324 ( .B1(n14738), .B2(n11231), .A(n11230), .ZN(n11233) );
  OAI22_X1 U14325 ( .A1(n14739), .A2(n10463), .B1(n11114), .B2(n14740), .ZN(
        n11232) );
  NOR2_X1 U14326 ( .A1(n11233), .A2(n11232), .ZN(n11239) );
  AOI22_X1 U14327 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11234) );
  OAI21_X1 U14328 ( .B1(n14737), .B2(n10472), .A(n11234), .ZN(n11235) );
  INV_X1 U14329 ( .A(n11235), .ZN(n11238) );
  AOI22_X1 U14330 ( .A1(n11236), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10426), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11237) );
  NAND4_X1 U14331 ( .A1(n11240), .A2(n11239), .A3(n11238), .A4(n11237), .ZN(
        n13553) );
  INV_X1 U14332 ( .A(n13553), .ZN(n11243) );
  AOI22_X1 U14333 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n11241) );
  OAI21_X1 U14334 ( .B1(n11243), .B2(n11242), .A(n11241), .ZN(n11244) );
  AOI21_X1 U14335 ( .B1(n9785), .B2(P2_REIP_REG_14__SCAN_IN), .A(n11244), .ZN(
        n16280) );
  NOR2_X2 U14336 ( .A1(n16281), .A2(n16280), .ZN(n16279) );
  AOI22_X1 U14337 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11248) );
  NAND2_X1 U14338 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11247) );
  NAND2_X1 U14339 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11246) );
  NAND2_X1 U14340 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11245) );
  NAND4_X1 U14341 ( .A1(n11248), .A2(n11247), .A3(n11246), .A4(n11245), .ZN(
        n11251) );
  INV_X1 U14342 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19265) );
  INV_X1 U14343 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11249) );
  OAI22_X1 U14344 ( .A1(n19265), .A2(n10464), .B1(n10463), .B2(n11249), .ZN(
        n11250) );
  NOR2_X1 U14345 ( .A1(n11251), .A2(n11250), .ZN(n11263) );
  OR2_X1 U14346 ( .A1(n10467), .A2(n11252), .ZN(n11256) );
  AOI22_X1 U14347 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11255) );
  NAND2_X1 U14348 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11254) );
  NAND2_X1 U14349 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11253) );
  AND4_X1 U14350 ( .A1(n11256), .A2(n11255), .A3(n11254), .A4(n11253), .ZN(
        n11262) );
  OAI22_X1 U14351 ( .A1(n10472), .A2(n11257), .B1(n14738), .B2(n14924), .ZN(
        n11260) );
  INV_X1 U14352 ( .A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11258) );
  INV_X1 U14353 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14772) );
  OAI22_X1 U14354 ( .A1(n11258), .A2(n10473), .B1(n11114), .B2(n14772), .ZN(
        n11259) );
  NOR2_X1 U14355 ( .A1(n11260), .A2(n11259), .ZN(n11261) );
  INV_X1 U14356 ( .A(n19078), .ZN(n11264) );
  AOI22_X1 U14357 ( .A1(n9785), .A2(P2_REIP_REG_15__SCAN_IN), .B1(n11265), 
        .B2(n11264), .ZN(n11267) );
  AOI22_X1 U14358 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n11266) );
  NAND2_X1 U14359 ( .A1(n11267), .A2(n11266), .ZN(n15384) );
  AOI22_X1 U14360 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n11269) );
  NAND2_X1 U14361 ( .A1(n9785), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11268) );
  INV_X1 U14362 ( .A(n9785), .ZN(n11297) );
  INV_X1 U14363 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19784) );
  NAND2_X1 U14364 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11271) );
  NAND2_X1 U14365 ( .A1(n11308), .A2(P2_EAX_REG_17__SCAN_IN), .ZN(n11270) );
  OAI211_X1 U14366 ( .C1(n11297), .C2(n19784), .A(n11271), .B(n11270), .ZN(
        n13808) );
  AOI22_X1 U14367 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n11273) );
  NAND2_X1 U14368 ( .A1(n9785), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11272) );
  AOI22_X1 U14369 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n11275) );
  NAND2_X1 U14370 ( .A1(n9785), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11274) );
  INV_X1 U14371 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19789) );
  NAND2_X1 U14372 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11277) );
  NAND2_X1 U14373 ( .A1(n11308), .A2(P2_EAX_REG_20__SCAN_IN), .ZN(n11276) );
  OAI211_X1 U14374 ( .C1(n11297), .C2(n19789), .A(n11277), .B(n11276), .ZN(
        n14631) );
  INV_X1 U14375 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19790) );
  NAND2_X1 U14376 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11279) );
  NAND2_X1 U14377 ( .A1(n11308), .A2(P2_EAX_REG_21__SCAN_IN), .ZN(n11278) );
  OAI211_X1 U14378 ( .C1(n11297), .C2(n19790), .A(n11279), .B(n11278), .ZN(
        n15075) );
  AOI22_X1 U14379 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n11281) );
  NAND2_X1 U14380 ( .A1(n9785), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U14381 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n11283) );
  NAND2_X1 U14382 ( .A1(n9785), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11282) );
  AND2_X1 U14383 ( .A1(n11283), .A2(n11282), .ZN(n15051) );
  AOI22_X1 U14384 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n11285) );
  NAND2_X1 U14385 ( .A1(n9785), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11284) );
  NOR2_X2 U14386 ( .A1(n15054), .A2(n15044), .ZN(n15045) );
  INV_X1 U14387 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19797) );
  NAND2_X1 U14388 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11287) );
  NAND2_X1 U14389 ( .A1(n11308), .A2(P2_EAX_REG_25__SCAN_IN), .ZN(n11286) );
  OAI211_X1 U14390 ( .C1(n11297), .C2(n19797), .A(n11287), .B(n11286), .ZN(
        n15035) );
  NAND2_X1 U14391 ( .A1(n15045), .A2(n15035), .ZN(n15037) );
  AOI22_X1 U14392 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n11289) );
  NAND2_X1 U14393 ( .A1(n9785), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11288) );
  AND2_X1 U14394 ( .A1(n11289), .A2(n11288), .ZN(n15024) );
  AOI22_X1 U14395 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n11308), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n11291) );
  NAND2_X1 U14396 ( .A1(n9785), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11290) );
  AND2_X1 U14397 ( .A1(n11291), .A2(n11290), .ZN(n15015) );
  NAND2_X1 U14398 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11293) );
  NAND2_X1 U14399 ( .A1(n11308), .A2(P2_EAX_REG_28__SCAN_IN), .ZN(n11292) );
  OAI211_X1 U14400 ( .C1(n11297), .C2(n11294), .A(n11293), .B(n11292), .ZN(
        n15009) );
  INV_X1 U14401 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19803) );
  NAND2_X1 U14402 ( .A1(n11075), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11296) );
  NAND2_X1 U14403 ( .A1(n11308), .A2(P2_EAX_REG_29__SCAN_IN), .ZN(n11295) );
  OAI211_X1 U14404 ( .C1(n11297), .C2(n19803), .A(n11296), .B(n11295), .ZN(
        n11413) );
  NOR2_X2 U14405 ( .A1(n9638), .A2(n11298), .ZN(n11310) );
  AOI21_X1 U14406 ( .B1(n11298), .B2(n9638), .A(n11310), .ZN(n14995) );
  INV_X1 U14407 ( .A(n11299), .ZN(n11301) );
  NAND2_X1 U14408 ( .A1(n11301), .A2(n11300), .ZN(n13296) );
  NAND2_X1 U14409 ( .A1(n13464), .A2(n11027), .ZN(n11302) );
  AND2_X1 U14410 ( .A1(n13296), .A2(n11302), .ZN(n11303) );
  NAND2_X1 U14411 ( .A1(n10160), .A2(n11307), .ZN(P2_U3016) );
  AOI222_X1 U14412 ( .A1(n9785), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n11075), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C1(n11308), .C2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n11309) );
  XNOR2_X1 U14413 ( .A(n11310), .B(n11309), .ZN(n19104) );
  NAND2_X1 U14414 ( .A1(n13464), .A2(n11368), .ZN(n12916) );
  INV_X1 U14415 ( .A(n16351), .ZN(n12868) );
  NAND2_X1 U14416 ( .A1(n19818), .A2(n12778), .ZN(n11370) );
  OR2_X1 U14417 ( .A1(n11311), .A2(n11370), .ZN(n13503) );
  NOR2_X2 U14418 ( .A1(n18861), .A2(n13503), .ZN(n19061) );
  AOI22_X1 U14419 ( .A1(n10330), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11315) );
  NAND2_X1 U14420 ( .A1(n11313), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n11314) );
  NAND2_X1 U14421 ( .A1(n11315), .A2(n11314), .ZN(n11316) );
  AOI21_X1 U14422 ( .B1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n10873), .A(
        n11316), .ZN(n11317) );
  INV_X1 U14423 ( .A(n16355), .ZN(n19743) );
  NOR2_X1 U14424 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19743), .ZN(n13655) );
  NAND2_X1 U14425 ( .A1(n10983), .A2(n13655), .ZN(n11320) );
  NOR2_X2 U14426 ( .A1(n18861), .A2(n11320), .ZN(n19064) );
  INV_X1 U14427 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11323) );
  INV_X1 U14428 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11321) );
  INV_X1 U14429 ( .A(n11324), .ZN(n11326) );
  AOI21_X1 U14430 ( .B1(n11326), .B2(n11430), .A(n11325), .ZN(n11432) );
  INV_X1 U14431 ( .A(n11432), .ZN(n16091) );
  AOI21_X1 U14432 ( .B1(n20923), .B2(n11330), .A(n11327), .ZN(n15095) );
  INV_X1 U14433 ( .A(n15095), .ZN(n16113) );
  NAND2_X1 U14434 ( .A1(n11331), .A2(n11328), .ZN(n11329) );
  NAND2_X1 U14435 ( .A1(n11330), .A2(n11329), .ZN(n16124) );
  INV_X1 U14436 ( .A(n11331), .ZN(n11332) );
  AOI21_X1 U14437 ( .B1(n15105), .B2(n11334), .A(n11332), .ZN(n15107) );
  INV_X1 U14438 ( .A(n15107), .ZN(n16136) );
  OR2_X1 U14439 ( .A1(n11336), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11333) );
  NAND2_X1 U14440 ( .A1(n11334), .A2(n11333), .ZN(n16147) );
  AND2_X1 U14441 ( .A1(n11337), .A2(n15128), .ZN(n11335) );
  NOR2_X1 U14442 ( .A1(n11336), .A2(n11335), .ZN(n15126) );
  INV_X1 U14443 ( .A(n15126), .ZN(n16157) );
  OAI21_X1 U14444 ( .B1(n11338), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n11337), .ZN(n15610) );
  AOI21_X1 U14445 ( .B1(n11358), .B2(n18890), .A(n11338), .ZN(n15159) );
  INV_X1 U14446 ( .A(n15159), .ZN(n18887) );
  AOI21_X1 U14447 ( .B1(n11339), .B2(n11356), .A(n9754), .ZN(n15180) );
  OAI21_X1 U14448 ( .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n11353), .A(
        n11355), .ZN(n13918) );
  INV_X1 U14449 ( .A(n13918), .ZN(n15210) );
  AOI21_X1 U14450 ( .B1(n10820), .B2(n11352), .A(n11340), .ZN(n18930) );
  AOI21_X1 U14451 ( .B1(n16216), .B2(n11350), .A(n9753), .ZN(n18941) );
  AOI21_X1 U14452 ( .B1(n10861), .B2(n11348), .A(n11351), .ZN(n18971) );
  AOI21_X1 U14453 ( .B1(n10825), .B2(n11346), .A(n11349), .ZN(n18987) );
  AOI21_X1 U14454 ( .B1(n10847), .B2(n11344), .A(n11347), .ZN(n19007) );
  AOI21_X1 U14455 ( .B1(n10838), .B2(n11342), .A(n11345), .ZN(n19034) );
  AOI21_X1 U14456 ( .B1(n10343), .B2(n11341), .A(n11343), .ZN(n16267) );
  OAI22_X1 U14457 ( .A1(n16342), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n15450) );
  INV_X1 U14458 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n12863) );
  OAI22_X1 U14459 ( .A1(n16342), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n12863), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14678) );
  AND2_X1 U14460 ( .A1(n15450), .A2(n14678), .ZN(n14662) );
  OAI21_X1 U14461 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n11341), .ZN(n14664) );
  NAND2_X1 U14462 ( .A1(n14662), .A2(n14664), .ZN(n13653) );
  NOR2_X1 U14463 ( .A1(n16267), .A2(n13653), .ZN(n19040) );
  OAI21_X1 U14464 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n11343), .A(
        n11342), .ZN(n19228) );
  NAND2_X1 U14465 ( .A1(n19040), .A2(n19228), .ZN(n19032) );
  NOR2_X1 U14466 ( .A1(n19034), .A2(n19032), .ZN(n19021) );
  OAI21_X1 U14467 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n11345), .A(
        n11344), .ZN(n19022) );
  NAND2_X1 U14468 ( .A1(n19021), .A2(n19022), .ZN(n19006) );
  NOR2_X1 U14469 ( .A1(n19007), .A2(n19006), .ZN(n18996) );
  OAI21_X1 U14470 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n11347), .A(
        n11346), .ZN(n18997) );
  NAND2_X1 U14471 ( .A1(n18996), .A2(n18997), .ZN(n18986) );
  NOR2_X1 U14472 ( .A1(n18987), .A2(n18986), .ZN(n18976) );
  OAI21_X1 U14473 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n11349), .A(
        n11348), .ZN(n18977) );
  NAND2_X1 U14474 ( .A1(n18976), .A2(n18977), .ZN(n18969) );
  NOR2_X1 U14475 ( .A1(n18971), .A2(n18969), .ZN(n18959) );
  OAI21_X1 U14476 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n11351), .A(
        n11350), .ZN(n18960) );
  NAND2_X1 U14477 ( .A1(n18959), .A2(n18960), .ZN(n18950) );
  NOR2_X1 U14478 ( .A1(n18941), .A2(n18950), .ZN(n18932) );
  OAI21_X1 U14479 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n9753), .A(
        n11352), .ZN(n18933) );
  NAND2_X1 U14480 ( .A1(n18932), .A2(n18933), .ZN(n18929) );
  NOR2_X1 U14481 ( .A1(n18930), .A2(n18929), .ZN(n18909) );
  AOI21_X1 U14482 ( .B1(n10876), .B2(n11354), .A(n11353), .ZN(n18920) );
  INV_X1 U14483 ( .A(n18920), .ZN(n18911) );
  NAND2_X1 U14484 ( .A1(n18909), .A2(n18911), .ZN(n13916) );
  NOR2_X1 U14485 ( .A1(n15210), .A2(n13916), .ZN(n18897) );
  INV_X1 U14486 ( .A(n11355), .ZN(n11357) );
  OAI21_X1 U14487 ( .B1(n11357), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n11356), .ZN(n18898) );
  NAND2_X1 U14488 ( .A1(n18897), .A2(n18898), .ZN(n14646) );
  NOR2_X1 U14489 ( .A1(n15180), .A2(n14646), .ZN(n14638) );
  OAI21_X1 U14490 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n9754), .A(
        n11358), .ZN(n15171) );
  NAND2_X1 U14491 ( .A1(n14638), .A2(n15171), .ZN(n14637) );
  NAND2_X1 U14492 ( .A1(n11360), .A2(n14637), .ZN(n18886) );
  NAND2_X1 U14493 ( .A1(n18887), .A2(n18886), .ZN(n18885) );
  NAND2_X1 U14494 ( .A1(n9690), .A2(n15609), .ZN(n16156) );
  NAND2_X1 U14495 ( .A1(n16157), .A2(n16156), .ZN(n16155) );
  NAND2_X1 U14496 ( .A1(n9690), .A2(n16155), .ZN(n16146) );
  NAND2_X1 U14497 ( .A1(n16147), .A2(n16146), .ZN(n16145) );
  NAND2_X1 U14498 ( .A1(n9690), .A2(n16145), .ZN(n16135) );
  NAND2_X1 U14499 ( .A1(n16136), .A2(n16135), .ZN(n16134) );
  NAND2_X1 U14500 ( .A1(n9690), .A2(n16134), .ZN(n16123) );
  NAND2_X1 U14501 ( .A1(n16124), .A2(n16123), .ZN(n16122) );
  NAND2_X1 U14502 ( .A1(n9690), .A2(n16122), .ZN(n16112) );
  NAND2_X1 U14503 ( .A1(n16113), .A2(n16112), .ZN(n16111) );
  NAND2_X1 U14504 ( .A1(n9690), .A2(n16111), .ZN(n16102) );
  NAND2_X1 U14505 ( .A1(n16103), .A2(n16102), .ZN(n16101) );
  NAND2_X1 U14506 ( .A1(n11360), .A2(n16101), .ZN(n16090) );
  NAND2_X1 U14507 ( .A1(n16091), .A2(n16090), .ZN(n16089) );
  NAND2_X1 U14508 ( .A1(n9690), .A2(n16089), .ZN(n14620) );
  NOR4_X1 U14509 ( .A1(n15457), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(
        P2_STATE2_REG_0__SCAN_IN), .A4(P2_STATEBS16_REG_SCAN_IN), .ZN(n11359)
         );
  NOR2_X1 U14510 ( .A1(n19077), .A2(n19041), .ZN(n18910) );
  NOR2_X1 U14511 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19825), .ZN(n19437) );
  NAND2_X1 U14512 ( .A1(n11361), .A2(n19437), .ZN(n16352) );
  NAND2_X1 U14513 ( .A1(n19068), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19071) );
  INV_X1 U14514 ( .A(n11362), .ZN(n11363) );
  NAND2_X1 U14515 ( .A1(n11363), .A2(n10960), .ZN(n11364) );
  MUX2_X1 U14516 ( .A(n11365), .B(n11364), .S(n9649), .Z(n11385) );
  OAI21_X1 U14517 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n19743), .A(n10983), 
        .ZN(n11366) );
  NOR2_X1 U14518 ( .A1(n18861), .A2(n11366), .ZN(n13660) );
  INV_X1 U14519 ( .A(n13660), .ZN(n11371) );
  NAND2_X1 U14520 ( .A1(n11368), .A2(n11367), .ZN(n11369) );
  NAND2_X1 U14521 ( .A1(n12840), .A2(n11370), .ZN(n13659) );
  OAI21_X1 U14522 ( .B1(n11385), .B2(n11371), .A(n13659), .ZN(n11372) );
  AOI22_X1 U14523 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n19028), .B1(
        P2_EBX_REG_31__SCAN_IN), .B2(n11372), .ZN(n11374) );
  INV_X1 U14524 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19808) );
  OR2_X1 U14525 ( .A1(n19068), .A2(n19808), .ZN(n11373) );
  NAND2_X1 U14526 ( .A1(n11410), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11376) );
  NOR2_X1 U14527 ( .A1(n19046), .A2(n19808), .ZN(n14136) );
  AOI21_X1 U14528 ( .B1(n19218), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14136), .ZN(n11380) );
  INV_X1 U14529 ( .A(n11377), .ZN(n11378) );
  NAND2_X1 U14530 ( .A1(n16268), .A2(n11378), .ZN(n11379) );
  OAI211_X1 U14531 ( .C1(n16163), .C2(n16273), .A(n11380), .B(n11379), .ZN(
        n11381) );
  AOI21_X1 U14532 ( .B1(n14142), .B2(n16269), .A(n11381), .ZN(n11392) );
  NOR2_X1 U14533 ( .A1(n11385), .A2(n10640), .ZN(n11386) );
  XNOR2_X1 U14534 ( .A(n11386), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11387) );
  XNOR2_X1 U14535 ( .A(n11388), .B(n11387), .ZN(n14145) );
  INV_X1 U14536 ( .A(n14145), .ZN(n11390) );
  NAND2_X1 U14537 ( .A1(n11390), .A2(n11389), .ZN(n11391) );
  NAND2_X1 U14538 ( .A1(n11392), .A2(n11391), .ZN(P2_U2983) );
  NAND2_X1 U14539 ( .A1(n11393), .A2(n11395), .ZN(n15267) );
  NOR2_X1 U14540 ( .A1(n15267), .A2(n19219), .ZN(n11409) );
  INV_X1 U14541 ( .A(n15102), .ZN(n11397) );
  AOI21_X1 U14542 ( .B1(n11396), .B2(n15101), .A(n11397), .ZN(n11399) );
  MUX2_X1 U14543 ( .A(n11399), .B(n15101), .S(n11398), .Z(n11400) );
  NAND2_X1 U14544 ( .A1(n11400), .A2(n9724), .ZN(n15278) );
  NAND2_X1 U14545 ( .A1(n11401), .A2(n11402), .ZN(n11403) );
  INV_X1 U14546 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n11404) );
  NOR2_X1 U14547 ( .A1(n19046), .A2(n11404), .ZN(n15268) );
  AOI21_X1 U14548 ( .B1(n19218), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15268), .ZN(n11405) );
  OAI21_X1 U14549 ( .B1(n19229), .B2(n16124), .A(n11405), .ZN(n11406) );
  AOI21_X1 U14550 ( .B1(n15092), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11411) );
  OAI21_X1 U14551 ( .B1(n11412), .B2(n11413), .A(n9638), .ZN(n16086) );
  OAI21_X1 U14552 ( .B1(n11416), .B2(n11415), .A(n11414), .ZN(n14946) );
  INV_X1 U14553 ( .A(n14946), .ZN(n16087) );
  INV_X1 U14554 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11418) );
  NAND2_X1 U14555 ( .A1(n19217), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11429) );
  OAI21_X1 U14556 ( .B1(n15259), .B2(n11418), .A(n11429), .ZN(n11420) );
  INV_X1 U14557 ( .A(n14133), .ZN(n11417) );
  AOI211_X1 U14558 ( .C1(n15247), .C2(n11418), .A(n11417), .B(n15255), .ZN(
        n11419) );
  AOI211_X1 U14559 ( .C1(n16087), .C2(n16316), .A(n11420), .B(n11419), .ZN(
        n11421) );
  OAI21_X1 U14560 ( .B1(n16086), .B2(n16330), .A(n11421), .ZN(n11422) );
  AOI21_X1 U14561 ( .B1(n11435), .B2(n16314), .A(n11422), .ZN(n11428) );
  NOR2_X1 U14562 ( .A1(n11424), .A2(n11423), .ZN(n11426) );
  XOR2_X1 U14563 ( .A(n11426), .B(n11425), .Z(n11436) );
  NAND2_X1 U14564 ( .A1(n11428), .A2(n11427), .ZN(P2_U3017) );
  OAI21_X1 U14565 ( .B1(n16278), .B2(n11430), .A(n11429), .ZN(n11431) );
  AOI21_X1 U14566 ( .B1(n16268), .B2(n11432), .A(n11431), .ZN(n11433) );
  OAI21_X1 U14567 ( .B1(n14946), .B2(n16273), .A(n11433), .ZN(n11434) );
  AOI21_X1 U14568 ( .B1(n11435), .B2(n16269), .A(n11434), .ZN(n11438) );
  NAND2_X1 U14569 ( .A1(n11438), .A2(n11437), .ZN(P2_U2985) );
  AOI22_X1 U14570 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11456) );
  NAND2_X2 U14571 ( .A1(n18796), .A2(n18807), .ZN(n11445) );
  AOI22_X1 U14572 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11455) );
  INV_X1 U14573 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n20953) );
  INV_X2 U14574 ( .A(n10155), .ZN(n15559) );
  AOI22_X1 U14575 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11440) );
  OAI21_X1 U14576 ( .B1(n14087), .B2(n20953), .A(n11440), .ZN(n11453) );
  NOR2_X2 U14577 ( .A1(n11441), .A2(n11447), .ZN(n11485) );
  AOI22_X1 U14578 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11451) );
  INV_X2 U14579 ( .A(n15530), .ZN(n17050) );
  NOR2_X2 U14580 ( .A1(n11445), .A2(n18665), .ZN(n11524) );
  AOI22_X1 U14581 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U14582 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11449) );
  AOI22_X1 U14583 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11448) );
  NAND4_X1 U14584 ( .A1(n11451), .A2(n11450), .A3(n11449), .A4(n11448), .ZN(
        n11452) );
  AOI211_X1 U14585 ( .C1(n9651), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n11453), .B(n11452), .ZN(n11454) );
  NAND3_X1 U14586 ( .A1(n11456), .A2(n11455), .A3(n11454), .ZN(n15581) );
  AOI22_X1 U14587 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14588 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11459) );
  AOI22_X1 U14589 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11458) );
  AOI22_X1 U14590 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11457) );
  NAND4_X1 U14591 ( .A1(n11460), .A2(n11459), .A3(n11458), .A4(n11457), .ZN(
        n11466) );
  AOI22_X1 U14592 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U14593 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U14594 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U14595 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11461) );
  NAND4_X1 U14596 ( .A1(n11464), .A2(n11463), .A3(n11462), .A4(n11461), .ZN(
        n11465) );
  AOI22_X1 U14597 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11470) );
  AOI22_X1 U14598 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n9667), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11469) );
  AOI22_X1 U14599 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11468) );
  AOI22_X1 U14600 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11467) );
  NAND4_X1 U14601 ( .A1(n11470), .A2(n11469), .A3(n11468), .A4(n11467), .ZN(
        n11476) );
  AOI22_X1 U14602 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14603 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U14604 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11472) );
  INV_X2 U14605 ( .A(n10155), .ZN(n17124) );
  AOI22_X1 U14606 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11471) );
  NAND4_X1 U14607 ( .A1(n11474), .A2(n11473), .A3(n11472), .A4(n11471), .ZN(
        n11475) );
  AOI22_X1 U14608 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(n9653), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14609 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11483) );
  INV_X1 U14610 ( .A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n15529) );
  AOI22_X1 U14611 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11478) );
  AOI22_X1 U14612 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U14613 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14614 ( .A1(n11488), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11480) );
  AOI22_X1 U14615 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11525), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11479) );
  INV_X2 U14616 ( .A(n15541), .ZN(n17151) );
  AOI22_X1 U14617 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17151), .B1(
        n17138), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11496) );
  AOI22_X1 U14618 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17149), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n9653), .ZN(n11495) );
  INV_X1 U14619 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17216) );
  AOI22_X1 U14620 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11487) );
  OAI21_X1 U14621 ( .B1(n10157), .B2(n17216), .A(n11487), .ZN(n11493) );
  AOI22_X1 U14622 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11443), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11492) );
  AOI22_X1 U14623 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n9652), .ZN(n11491) );
  AOI22_X1 U14624 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11488), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U14625 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17124), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n11525), .ZN(n11489) );
  NAND2_X1 U14626 ( .A1(n17364), .A2(n11726), .ZN(n11522) );
  AOI22_X1 U14627 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U14628 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11506) );
  INV_X1 U14629 ( .A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n21097) );
  AOI22_X1 U14630 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11498) );
  OAI21_X1 U14631 ( .B1(n14087), .B2(n21097), .A(n11498), .ZN(n11504) );
  AOI22_X1 U14632 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11502) );
  AOI22_X1 U14633 ( .A1(n15559), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11501) );
  AOI22_X1 U14634 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U14635 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11525), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11499) );
  NAND4_X1 U14636 ( .A1(n11502), .A2(n11501), .A3(n11500), .A4(n11499), .ZN(
        n11503) );
  AOI211_X1 U14637 ( .C1(n17050), .C2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n11504), .B(n11503), .ZN(n11505) );
  NAND3_X1 U14638 ( .A1(n11507), .A2(n11506), .A3(n11505), .ZN(n17354) );
  NAND2_X1 U14639 ( .A1(n11544), .A2(n17354), .ZN(n11521) );
  AOI22_X1 U14640 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U14641 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11516) );
  AOI22_X1 U14642 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(n9655), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11508) );
  OAI21_X1 U14643 ( .B1(n9713), .B2(n21092), .A(n11508), .ZN(n11514) );
  AOI22_X1 U14644 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11485), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11512) );
  AOI22_X1 U14645 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n9667), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11511) );
  AOI22_X1 U14646 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11510) );
  AOI22_X1 U14647 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11509) );
  NAND4_X1 U14648 ( .A1(n11512), .A2(n11511), .A3(n11510), .A4(n11509), .ZN(
        n11513) );
  AOI211_X1 U14649 ( .C1(n17050), .C2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A(
        n11514), .B(n11513), .ZN(n11515) );
  NAND3_X1 U14650 ( .A1(n11517), .A2(n11516), .A3(n11515), .ZN(n17344) );
  NOR2_X4 U14651 ( .A1(n17341), .A2(n11552), .ZN(n17767) );
  INV_X1 U14652 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17500) );
  AOI22_X1 U14653 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17645), .B1(
        n17767), .B2(n17500), .ZN(n17504) );
  INV_X1 U14654 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17892) );
  NOR2_X1 U14655 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17767), .ZN(
        n17629) );
  INV_X1 U14656 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17964) );
  NAND2_X1 U14657 ( .A1(n17629), .A2(n17964), .ZN(n11518) );
  NOR2_X1 U14658 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11518), .ZN(
        n17594) );
  INV_X1 U14659 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17596) );
  NAND2_X1 U14660 ( .A1(n17594), .A2(n17596), .ZN(n17576) );
  INV_X1 U14661 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17995) );
  INV_X1 U14662 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17979) );
  NOR2_X1 U14663 ( .A1(n17995), .A2(n17979), .ZN(n17971) );
  INV_X1 U14664 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17608) );
  NOR2_X1 U14665 ( .A1(n17964), .A2(n17608), .ZN(n17942) );
  AND3_X1 U14666 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n17942), .ZN(n11560) );
  AND2_X1 U14667 ( .A1(n17971), .A2(n11560), .ZN(n17932) );
  AND2_X1 U14668 ( .A1(n17932), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n17913) );
  NAND2_X1 U14669 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17913), .ZN(
        n17551) );
  INV_X1 U14670 ( .A(n17551), .ZN(n17898) );
  NAND2_X1 U14671 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17720) );
  INV_X1 U14672 ( .A(n17720), .ZN(n18056) );
  NAND2_X1 U14673 ( .A1(n18056), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18038) );
  INV_X1 U14674 ( .A(n18038), .ZN(n18027) );
  NAND2_X1 U14675 ( .A1(n18027), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18013) );
  INV_X1 U14676 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18015) );
  INV_X1 U14677 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18026) );
  NOR3_X1 U14678 ( .A1(n18013), .A2(n18015), .A3(n18026), .ZN(n18012) );
  INV_X1 U14679 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18088) );
  XOR2_X1 U14680 ( .A(n17344), .B(n11519), .Z(n11520) );
  NAND2_X1 U14681 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11520), .ZN(
        n11551) );
  XOR2_X1 U14682 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n11520), .Z(
        n17790) );
  XOR2_X1 U14683 ( .A(n17350), .B(n11521), .Z(n11547) );
  XOR2_X1 U14684 ( .A(n17358), .B(n11522), .Z(n11540) );
  INV_X1 U14685 ( .A(n11726), .ZN(n17376) );
  NAND2_X1 U14686 ( .A1(n17376), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11537) );
  AOI22_X1 U14687 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11529) );
  AOI22_X1 U14688 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11528) );
  BUF_X2 U14689 ( .A(n11524), .Z(n17055) );
  AOI22_X1 U14690 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14691 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11525), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11526) );
  NAND4_X1 U14692 ( .A1(n11529), .A2(n11528), .A3(n11527), .A4(n11526), .ZN(
        n11536) );
  AOI22_X1 U14693 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11534) );
  AOI22_X1 U14694 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14695 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14696 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11531) );
  NAND4_X1 U14697 ( .A1(n11534), .A2(n11533), .A3(n11532), .A4(n11531), .ZN(
        n11535) );
  NOR2_X1 U14698 ( .A1(n11536), .A2(n11535), .ZN(n17857) );
  INV_X1 U14699 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18817) );
  NOR2_X1 U14700 ( .A1(n17857), .A2(n18817), .ZN(n17856) );
  NAND2_X1 U14701 ( .A1(n11537), .A2(n17847), .ZN(n17836) );
  INV_X1 U14702 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18147) );
  OR2_X1 U14703 ( .A1(n18147), .A2(n11538), .ZN(n11539) );
  NAND2_X1 U14704 ( .A1(n11540), .A2(n11542), .ZN(n11543) );
  NAND2_X1 U14705 ( .A1(n11543), .A2(n17825), .ZN(n17818) );
  XOR2_X1 U14706 ( .A(n17354), .B(n11544), .Z(n11545) );
  XOR2_X1 U14707 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n11545), .Z(
        n17819) );
  NAND2_X1 U14708 ( .A1(n17818), .A2(n17819), .ZN(n17817) );
  NAND2_X1 U14709 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11545), .ZN(
        n11546) );
  NAND2_X1 U14710 ( .A1(n11547), .A2(n11549), .ZN(n11550) );
  NAND2_X1 U14711 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n17802), .ZN(
        n17801) );
  NAND2_X1 U14712 ( .A1(n11550), .A2(n17801), .ZN(n17789) );
  NAND2_X1 U14713 ( .A1(n17790), .A2(n17789), .ZN(n17788) );
  AOI21_X1 U14714 ( .B1(n17341), .B2(n11552), .A(n17767), .ZN(n11554) );
  NAND2_X1 U14715 ( .A1(n11554), .A2(n11553), .ZN(n11555) );
  INV_X1 U14716 ( .A(n17920), .ZN(n17577) );
  INV_X1 U14717 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18073) );
  INV_X1 U14718 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18067) );
  NOR2_X1 U14719 ( .A1(n17666), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17681) );
  INV_X1 U14720 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18004) );
  AND2_X1 U14721 ( .A1(n18026), .A2(n18004), .ZN(n11557) );
  NAND2_X1 U14722 ( .A1(n17681), .A2(n11557), .ZN(n17646) );
  NAND2_X1 U14723 ( .A1(n17645), .A2(n17646), .ZN(n11559) );
  NOR2_X2 U14724 ( .A1(n17553), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17552) );
  NAND2_X1 U14725 ( .A1(n17971), .A2(n17577), .ZN(n17592) );
  INV_X1 U14726 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17918) );
  OR2_X1 U14727 ( .A1(n17767), .A2(n17552), .ZN(n17540) );
  NAND2_X1 U14728 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11643) );
  AOI21_X1 U14729 ( .B1(n17767), .B2(n17514), .A(n17513), .ZN(n17503) );
  NOR2_X1 U14730 ( .A1(n17504), .A2(n17503), .ZN(n17502) );
  AOI22_X1 U14731 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U14732 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14733 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11563) );
  AOI22_X1 U14734 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11562) );
  NAND4_X1 U14735 ( .A1(n11565), .A2(n11564), .A3(n11563), .A4(n11562), .ZN(
        n11571) );
  AOI22_X1 U14736 ( .A1(n15559), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U14737 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11568) );
  AOI22_X1 U14738 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U14739 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11566) );
  NAND4_X1 U14740 ( .A1(n11569), .A2(n11568), .A3(n11567), .A4(n11566), .ZN(
        n11570) );
  AOI22_X1 U14741 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n9652), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11575) );
  AOI22_X1 U14742 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11574) );
  AOI22_X1 U14743 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11573) );
  AOI22_X1 U14744 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11572) );
  NAND4_X1 U14745 ( .A1(n11575), .A2(n11574), .A3(n11573), .A4(n11572), .ZN(
        n11581) );
  AOI22_X1 U14746 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14747 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14748 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11577) );
  AOI22_X1 U14749 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11576) );
  NAND4_X1 U14750 ( .A1(n11579), .A2(n11578), .A3(n11577), .A4(n11576), .ZN(
        n11580) );
  NOR2_X4 U14751 ( .A1(n11581), .A2(n11580), .ZN(n18196) );
  AOI22_X1 U14752 ( .A1(n15559), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11585) );
  AOI22_X1 U14753 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14754 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14755 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11582) );
  NAND4_X1 U14756 ( .A1(n11585), .A2(n11584), .A3(n11583), .A4(n11582), .ZN(
        n11591) );
  AOI22_X1 U14757 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n9667), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11589) );
  AOI22_X1 U14758 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U14759 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U14760 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11586) );
  NAND4_X1 U14761 ( .A1(n11589), .A2(n11588), .A3(n11587), .A4(n11586), .ZN(
        n11590) );
  NAND2_X1 U14762 ( .A1(n18196), .A2(n18840), .ZN(n11704) );
  NOR2_X1 U14763 ( .A1(n18212), .A2(n11704), .ZN(n11710) );
  AOI22_X1 U14764 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U14765 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11594) );
  AOI22_X1 U14766 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U14767 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11592) );
  NAND4_X1 U14768 ( .A1(n11595), .A2(n11594), .A3(n11593), .A4(n11592), .ZN(
        n11601) );
  AOI22_X1 U14769 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U14770 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11598) );
  AOI22_X1 U14771 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U14772 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11596) );
  NAND4_X1 U14773 ( .A1(n11599), .A2(n11598), .A3(n11597), .A4(n11596), .ZN(
        n11600) );
  NAND2_X1 U14774 ( .A1(n18196), .A2(n11661), .ZN(n11649) );
  AOI22_X1 U14775 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14776 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14777 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14778 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11602) );
  NAND4_X1 U14779 ( .A1(n11605), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n11611) );
  AOI22_X1 U14780 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11609) );
  AOI22_X1 U14781 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11608) );
  AOI22_X1 U14782 ( .A1(n15559), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11607) );
  AOI22_X1 U14783 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11606) );
  NAND4_X1 U14784 ( .A1(n11609), .A2(n11608), .A3(n11607), .A4(n11606), .ZN(
        n11610) );
  AOI22_X1 U14785 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U14786 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11614) );
  AOI22_X1 U14787 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11613) );
  AOI22_X1 U14788 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11612) );
  NAND4_X1 U14789 ( .A1(n11615), .A2(n11614), .A3(n11613), .A4(n11612), .ZN(
        n11621) );
  AOI22_X1 U14790 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14791 ( .A1(n15559), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14792 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11617) );
  AOI22_X1 U14793 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11616) );
  NAND4_X1 U14794 ( .A1(n11619), .A2(n11618), .A3(n11617), .A4(n11616), .ZN(
        n11620) );
  AOI22_X1 U14795 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U14796 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14797 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U14798 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11622) );
  NAND4_X1 U14799 ( .A1(n11625), .A2(n11624), .A3(n11623), .A4(n11622), .ZN(
        n11631) );
  AOI22_X1 U14800 ( .A1(n11488), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U14801 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11628) );
  INV_X2 U14802 ( .A(n9713), .ZN(n17153) );
  AOI22_X1 U14803 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11627) );
  AOI22_X1 U14804 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11626) );
  NAND4_X1 U14805 ( .A1(n11629), .A2(n11628), .A3(n11627), .A4(n11626), .ZN(
        n11630) );
  NOR2_X4 U14806 ( .A1(n11631), .A2(n11630), .ZN(n18219) );
  AOI22_X1 U14807 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U14808 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11634) );
  AOI22_X1 U14809 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11633) );
  AOI22_X1 U14810 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11632) );
  NAND4_X1 U14811 ( .A1(n11635), .A2(n11634), .A3(n11633), .A4(n11632), .ZN(
        n11641) );
  AOI22_X1 U14812 ( .A1(n11488), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11639) );
  AOI22_X1 U14813 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11638) );
  AOI22_X1 U14814 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U14815 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11636) );
  NAND4_X1 U14816 ( .A1(n11639), .A2(n11638), .A3(n11637), .A4(n11636), .ZN(
        n11640) );
  NAND2_X1 U14817 ( .A1(n18208), .A2(n11644), .ZN(n11657) );
  OAI211_X1 U14818 ( .C1(n18204), .C2(n18645), .A(n11658), .B(n11657), .ZN(
        n11642) );
  NAND2_X1 U14819 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16403) );
  INV_X1 U14820 ( .A(n11643), .ZN(n17866) );
  INV_X1 U14821 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17906) );
  NOR2_X1 U14822 ( .A1(n17551), .A2(n17906), .ZN(n11671) );
  INV_X1 U14823 ( .A(n11671), .ZN(n17884) );
  NOR2_X1 U14824 ( .A1(n17884), .A2(n17920), .ZN(n17532) );
  NAND2_X1 U14825 ( .A1(n17866), .A2(n17532), .ZN(n17499) );
  OR2_X1 U14826 ( .A1(n16403), .A2(n17499), .ZN(n16398) );
  INV_X1 U14827 ( .A(n16356), .ZN(n18624) );
  NAND2_X1 U14828 ( .A1(n18624), .A2(n17341), .ZN(n18091) );
  NAND2_X1 U14829 ( .A1(n18192), .A2(n16540), .ZN(n11646) );
  NAND2_X1 U14830 ( .A1(n11661), .A2(n11646), .ZN(n18853) );
  NAND2_X1 U14831 ( .A1(n17229), .A2(n18196), .ZN(n11647) );
  NOR2_X1 U14832 ( .A1(n18204), .A2(n11644), .ZN(n18640) );
  INV_X1 U14833 ( .A(n11663), .ZN(n11645) );
  NAND4_X1 U14834 ( .A1(n18200), .A2(n18204), .A3(n11645), .A4(n11651), .ZN(
        n11660) );
  NAND3_X1 U14835 ( .A1(n18196), .A2(n18204), .A3(n18212), .ZN(n11659) );
  NOR2_X1 U14836 ( .A1(n18219), .A2(n18645), .ZN(n15714) );
  NOR2_X1 U14837 ( .A1(n15714), .A2(n11646), .ZN(n11680) );
  AOI21_X1 U14838 ( .B1(n11647), .B2(n11659), .A(n11680), .ZN(n11656) );
  NAND2_X1 U14839 ( .A1(n18196), .A2(n11651), .ZN(n11701) );
  NAND2_X1 U14840 ( .A1(n11659), .A2(n11701), .ZN(n11655) );
  AOI22_X1 U14841 ( .A1(n11663), .A2(n18200), .B1(n18204), .B2(n18645), .ZN(
        n11648) );
  INV_X1 U14842 ( .A(n11648), .ZN(n11654) );
  NOR2_X1 U14843 ( .A1(n18219), .A2(n11651), .ZN(n11652) );
  INV_X1 U14844 ( .A(n11649), .ZN(n11650) );
  OAI22_X1 U14845 ( .A1(n18204), .A2(n11652), .B1(n11651), .B2(n11650), .ZN(
        n11653) );
  NAND2_X1 U14847 ( .A1(n18200), .A2(n18196), .ZN(n11664) );
  NAND2_X1 U14848 ( .A1(n18192), .A2(n15472), .ZN(n11662) );
  NOR2_X2 U14849 ( .A1(n14078), .A2(n11665), .ZN(n18646) );
  NOR2_X1 U14850 ( .A1(n18635), .A2(n18633), .ZN(n18064) );
  INV_X1 U14851 ( .A(n11664), .ZN(n18639) );
  INV_X1 U14852 ( .A(n11666), .ZN(n11670) );
  INV_X1 U14853 ( .A(n14079), .ZN(n11667) );
  NAND3_X1 U14854 ( .A1(n11668), .A2(n18840), .A3(n11667), .ZN(n11669) );
  AOI21_X4 U14855 ( .B1(n18639), .B2(n18658), .A(n18638), .ZN(n18059) );
  NAND2_X1 U14856 ( .A1(n11671), .A2(n17866), .ZN(n16379) );
  INV_X1 U14857 ( .A(n16379), .ZN(n11673) );
  NAND2_X1 U14858 ( .A1(n18012), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17647) );
  INV_X1 U14859 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18801) );
  NOR2_X1 U14860 ( .A1(n18147), .A2(n18801), .ZN(n18079) );
  INV_X1 U14861 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18117) );
  INV_X1 U14862 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18132) );
  INV_X1 U14863 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20931) );
  NOR3_X1 U14864 ( .A1(n18117), .A2(n18132), .A3(n20931), .ZN(n18087) );
  NAND4_X1 U14865 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A4(n18087), .ZN(n17965) );
  INV_X1 U14866 ( .A(n17965), .ZN(n11672) );
  NAND2_X1 U14867 ( .A1(n18079), .A2(n11672), .ZN(n17985) );
  OR2_X1 U14868 ( .A1(n18817), .A2(n17985), .ZN(n18052) );
  NOR2_X1 U14869 ( .A1(n17647), .A2(n18052), .ZN(n17987) );
  NAND3_X1 U14870 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n11673), .A3(
        n17987), .ZN(n11675) );
  NOR2_X1 U14871 ( .A1(n17647), .A2(n17985), .ZN(n17968) );
  AOI21_X1 U14872 ( .B1(n17968), .B2(n11673), .A(n18646), .ZN(n11674) );
  OAI21_X1 U14873 ( .B1(n18817), .B2(n18801), .A(n18147), .ZN(n18144) );
  NAND2_X1 U14874 ( .A1(n11672), .A2(n18144), .ZN(n17986) );
  NOR2_X1 U14875 ( .A1(n17647), .A2(n17986), .ZN(n17903) );
  AOI21_X1 U14876 ( .B1(n17903), .B2(n11673), .A(n18662), .ZN(n17871) );
  AOI211_X1 U14877 ( .C1(n18656), .C2(n11675), .A(n11674), .B(n17871), .ZN(
        n15689) );
  NAND2_X1 U14878 ( .A1(n18800), .A2(n18790), .ZN(n18794) );
  OR3_X2 U14879 ( .A1(n18794), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18077) );
  AOI21_X1 U14880 ( .B1(n11678), .B2(n11677), .A(n11676), .ZN(n11679) );
  OAI22_X1 U14881 ( .A1(n18814), .A2(n18649), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11697) );
  INV_X1 U14882 ( .A(n11697), .ZN(n11686) );
  INV_X1 U14883 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18670) );
  AOI22_X1 U14884 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18670), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18807), .ZN(n11689) );
  NAND2_X1 U14885 ( .A1(n11697), .A2(n11687), .ZN(n11681) );
  OAI21_X1 U14886 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18814), .A(
        n11681), .ZN(n11688) );
  NAND2_X1 U14887 ( .A1(n11689), .A2(n11688), .ZN(n11682) );
  NAND2_X1 U14888 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11683), .ZN(
        n11690) );
  OAI22_X1 U14889 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18674), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11683), .ZN(n11692) );
  AOI21_X1 U14890 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n11690), .A(
        n11692), .ZN(n11684) );
  AOI21_X1 U14891 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18674), .A(
        n11684), .ZN(n11693) );
  OAI21_X1 U14892 ( .B1(n11687), .B2(n11686), .A(n11693), .ZN(n11685) );
  AOI21_X1 U14893 ( .B1(n11687), .B2(n11686), .A(n11685), .ZN(n11702) );
  AOI21_X1 U14894 ( .B1(n18820), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n11687), .ZN(n11698) );
  INV_X1 U14895 ( .A(n11698), .ZN(n11696) );
  XOR2_X1 U14896 ( .A(n11689), .B(n11688), .Z(n11695) );
  NOR2_X1 U14897 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18674), .ZN(
        n11691) );
  AOI22_X1 U14898 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11692), .B1(
        n11691), .B2(n11690), .ZN(n11699) );
  INV_X1 U14899 ( .A(n11693), .ZN(n11694) );
  AOI21_X1 U14900 ( .B1(n11702), .B2(n11696), .A(n11703), .ZN(n18625) );
  INV_X1 U14901 ( .A(n18625), .ZN(n11709) );
  NAND3_X1 U14902 ( .A1(n11699), .A2(n11698), .A3(n11697), .ZN(n11700) );
  AOI21_X1 U14903 ( .B1(n18204), .B2(n11701), .A(n18620), .ZN(n11708) );
  NAND2_X1 U14904 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18710), .ZN(n18849) );
  NOR2_X1 U14905 ( .A1(n18849), .A2(n18718), .ZN(n18717) );
  NOR2_X1 U14906 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18704) );
  NOR3_X1 U14907 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18717), .A3(n18704), 
        .ZN(n18839) );
  OAI21_X1 U14908 ( .B1(n18196), .B2(n18840), .A(n11704), .ZN(n11705) );
  NAND2_X1 U14909 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18834) );
  OAI21_X1 U14910 ( .B1(n18839), .B2(n11705), .A(n18834), .ZN(n16521) );
  NOR3_X1 U14911 ( .A1(n11706), .A2(n18623), .A3(n16521), .ZN(n11707) );
  AOI211_X1 U14912 ( .C1(n11710), .C2(n11709), .A(n11708), .B(n11707), .ZN(
        n11711) );
  NAND2_X1 U14913 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18800), .ZN(n18693) );
  OAI211_X1 U14914 ( .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n18064), .A(
        n15689), .B(n18159), .ZN(n15584) );
  NOR2_X1 U14915 ( .A1(n17857), .A2(n17376), .ZN(n11722) );
  NOR2_X1 U14916 ( .A1(n11722), .A2(n17364), .ZN(n11720) );
  NOR2_X1 U14917 ( .A1(n11720), .A2(n17358), .ZN(n11719) );
  NAND2_X1 U14918 ( .A1(n11719), .A2(n17354), .ZN(n11717) );
  NOR2_X1 U14919 ( .A1(n17350), .A2(n11717), .ZN(n11716) );
  NAND2_X1 U14920 ( .A1(n11716), .A2(n17344), .ZN(n11715) );
  NOR2_X1 U14921 ( .A1(n17341), .A2(n11715), .ZN(n11738) );
  XOR2_X1 U14922 ( .A(n11715), .B(n17341), .Z(n17778) );
  XOR2_X1 U14923 ( .A(n11716), .B(n17344), .Z(n11731) );
  XOR2_X1 U14924 ( .A(n11717), .B(n17350), .Z(n11718) );
  NAND2_X1 U14925 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11718), .ZN(
        n11730) );
  XOR2_X1 U14926 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B(n11718), .Z(
        n17800) );
  XOR2_X1 U14927 ( .A(n11719), .B(n17354), .Z(n17812) );
  XOR2_X1 U14928 ( .A(n17358), .B(n11720), .Z(n11721) );
  NAND2_X1 U14929 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11721), .ZN(
        n11728) );
  XOR2_X1 U14930 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n11721), .Z(
        n17829) );
  XOR2_X1 U14931 ( .A(n17364), .B(n11722), .Z(n11723) );
  OR2_X1 U14932 ( .A1(n18147), .A2(n11723), .ZN(n11727) );
  XOR2_X1 U14933 ( .A(n18147), .B(n11723), .Z(n17840) );
  INV_X1 U14934 ( .A(n17857), .ZN(n15715) );
  AOI21_X1 U14935 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n11726), .A(
        n15715), .ZN(n11725) );
  NOR2_X1 U14936 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n11726), .ZN(
        n11724) );
  AOI221_X1 U14937 ( .B1(n15715), .B2(n11726), .C1(n11725), .C2(n18817), .A(
        n11724), .ZN(n17839) );
  NAND2_X1 U14938 ( .A1(n17840), .A2(n17839), .ZN(n17838) );
  NAND2_X1 U14939 ( .A1(n11727), .A2(n17838), .ZN(n17828) );
  NAND2_X1 U14940 ( .A1(n17829), .A2(n17828), .ZN(n17827) );
  NAND2_X1 U14941 ( .A1(n11728), .A2(n17827), .ZN(n17813) );
  NAND2_X1 U14942 ( .A1(n17812), .A2(n17813), .ZN(n17811) );
  NOR2_X1 U14943 ( .A1(n17812), .A2(n17813), .ZN(n11729) );
  AOI21_X1 U14944 ( .B1(n20931), .B2(n17811), .A(n11729), .ZN(n17799) );
  NAND2_X1 U14945 ( .A1(n17800), .A2(n17799), .ZN(n17798) );
  NAND2_X1 U14946 ( .A1(n11730), .A2(n17798), .ZN(n11732) );
  NAND2_X1 U14947 ( .A1(n11731), .A2(n11732), .ZN(n11733) );
  XOR2_X1 U14948 ( .A(n11732), .B(n11731), .Z(n17787) );
  NAND2_X1 U14949 ( .A1(n17787), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17786) );
  NAND2_X1 U14950 ( .A1(n11733), .A2(n17786), .ZN(n17777) );
  INV_X1 U14951 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18106) );
  NAND2_X1 U14952 ( .A1(n11738), .A2(n11734), .ZN(n11739) );
  INV_X1 U14953 ( .A(n11734), .ZN(n11737) );
  NAND2_X1 U14954 ( .A1(n17778), .A2(n17777), .ZN(n11736) );
  NAND2_X1 U14955 ( .A1(n11738), .A2(n11737), .ZN(n11735) );
  OAI211_X1 U14956 ( .C1(n11738), .C2(n11737), .A(n11736), .B(n11735), .ZN(
        n17757) );
  NAND2_X1 U14957 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17757), .ZN(
        n17756) );
  NOR2_X1 U14958 ( .A1(n18008), .A2(n17884), .ZN(n17539) );
  NAND2_X1 U14959 ( .A1(n17539), .A2(n17866), .ZN(n17498) );
  NOR2_X4 U14960 ( .A1(n18633), .A2(n18656), .ZN(n18143) );
  OAI21_X1 U14961 ( .B1(n17498), .B2(n16403), .A(n17923), .ZN(n11740) );
  AOI211_X1 U14962 ( .C1(n11741), .C2(n11740), .A(n9654), .B(n17500), .ZN(
        n11747) );
  NOR3_X4 U14963 ( .A1(n16356), .A2(n18173), .A3(n17341), .ZN(n18093) );
  NAND3_X1 U14964 ( .A1(n17513), .A2(n18093), .A3(n17504), .ZN(n11745) );
  NAND4_X1 U14965 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17767), .A3(
        n11742), .A4(n17500), .ZN(n11743) );
  NOR2_X1 U14966 ( .A1(n16356), .A2(n18173), .ZN(n18172) );
  OAI22_X1 U14967 ( .A1(n18627), .A2(n17728), .B1(n17766), .B2(n18091), .ZN(
        n17966) );
  INV_X1 U14968 ( .A(n17647), .ZN(n17967) );
  NAND2_X1 U14969 ( .A1(n17966), .A2(n17967), .ZN(n15576) );
  OAI21_X1 U14970 ( .B1(n18059), .B2(n18817), .A(n18646), .ZN(n18148) );
  AOI22_X1 U14971 ( .A1(n18635), .A2(n17903), .B1(n18148), .B2(n17968), .ZN(
        n15575) );
  NAND2_X1 U14972 ( .A1(n15576), .A2(n15575), .ZN(n17931) );
  NOR3_X1 U14973 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n9931), .A3(
        n16379), .ZN(n17507) );
  INV_X1 U14974 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18774) );
  NOR2_X1 U14975 ( .A1(n18077), .A2(n18774), .ZN(n17496) );
  NAND3_X1 U14976 ( .A1(n11745), .A2(n10171), .A3(n11744), .ZN(n11746) );
  NAND2_X1 U14977 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11751) );
  NAND2_X1 U14978 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11750) );
  AND2_X2 U14979 ( .A1(n11756), .A2(n11763), .ZN(n12025) );
  NAND2_X1 U14980 ( .A1(n12025), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11749) );
  NOR2_X4 U14981 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13161) );
  NAND2_X1 U14982 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11748) );
  NAND2_X1 U14983 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11755) );
  NAND2_X1 U14984 ( .A1(n12016), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11754) );
  NAND2_X1 U14985 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11753) );
  NAND2_X1 U14986 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11752) );
  NAND2_X1 U14987 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11773) );
  NAND2_X1 U14988 ( .A1(n9675), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11760) );
  AND2_X2 U14989 ( .A1(n13149), .A2(n14130), .ZN(n11820) );
  NAND2_X1 U14990 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11759) );
  NAND3_X1 U14991 ( .A1(n11760), .A2(n11759), .A3(n11758), .ZN(n11771) );
  NAND2_X1 U14992 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11769) );
  NAND2_X1 U14993 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11768) );
  AND2_X2 U14994 ( .A1(n11764), .A2(n11763), .ZN(n12011) );
  NAND2_X1 U14995 ( .A1(n12011), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11767) );
  NAND2_X1 U14996 ( .A1(n9672), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11766) );
  NAND4_X1 U14997 ( .A1(n11769), .A2(n11768), .A3(n11767), .A4(n11766), .ZN(
        n11770) );
  INV_X2 U14998 ( .A(n11878), .ZN(n13246) );
  NAND2_X1 U14999 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11778) );
  NAND2_X1 U15000 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11777) );
  NAND2_X1 U15001 ( .A1(n12560), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11776) );
  NAND2_X1 U15002 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11783) );
  NAND2_X1 U15003 ( .A1(n12025), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11782) );
  NAND2_X1 U15004 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11781) );
  NAND2_X1 U15005 ( .A1(n9642), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11780) );
  NAND2_X1 U15006 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11787) );
  NAND2_X1 U15007 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11786) );
  NAND2_X1 U15008 ( .A1(n12011), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11785) );
  NAND2_X1 U15009 ( .A1(n12034), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11784) );
  NAND2_X1 U15010 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11791) );
  NAND2_X1 U15011 ( .A1(n12016), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11790) );
  NAND2_X1 U15012 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11789) );
  NAND2_X1 U15013 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11788) );
  NAND4_X4 U15014 ( .A1(n11795), .A2(n11794), .A3(n11793), .A4(n11792), .ZN(
        n11877) );
  AOI22_X1 U15015 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12016), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U15016 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11929), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U15017 ( .A1(n12025), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12011), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U15018 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11796) );
  NAND4_X1 U15019 ( .A1(n11799), .A2(n11798), .A3(n11797), .A4(n11796), .ZN(
        n11808) );
  AOI22_X1 U15020 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11806) );
  AOI22_X1 U15021 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12026), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11805) );
  NAND2_X1 U15022 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11802) );
  AOI22_X1 U15023 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12017), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11803) );
  INV_X2 U15024 ( .A(n20119), .ZN(n13222) );
  AOI22_X1 U15025 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U15026 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12011), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U15027 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U15028 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U15029 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n12554), .B1(
        n11927), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U15030 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12016), .B1(
        n11928), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U15031 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n11929), .B1(
        n12017), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U15032 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n11930), .B1(
        n12560), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11813) );
  AND2_X1 U15033 ( .A1(n11877), .A2(n20136), .ZN(n11817) );
  NAND2_X1 U15034 ( .A1(n11817), .A2(n13222), .ZN(n11818) );
  AOI22_X1 U15035 ( .A1(n12554), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11927), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11824) );
  AOI22_X1 U15036 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12016), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11823) );
  AOI22_X1 U15037 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12017), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11822) );
  AOI22_X1 U15038 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11821) );
  NAND4_X1 U15039 ( .A1(n11824), .A2(n11823), .A3(n11822), .A4(n11821), .ZN(
        n11830) );
  AOI22_X1 U15040 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U15041 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12011), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U15042 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11826) );
  AOI22_X1 U15043 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11825) );
  NAND4_X1 U15044 ( .A1(n11828), .A2(n11827), .A3(n11826), .A4(n11825), .ZN(
        n11829) );
  AOI22_X1 U15045 ( .A1(n12554), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11927), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11834) );
  AOI22_X1 U15046 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U15047 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12026), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U15048 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12011), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11831) );
  NAND4_X1 U15049 ( .A1(n11834), .A2(n11833), .A3(n11832), .A4(n11831), .ZN(
        n11840) );
  AOI22_X1 U15050 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12016), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U15051 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11929), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U15052 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U15053 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12017), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11835) );
  NAND4_X1 U15054 ( .A1(n11838), .A2(n11837), .A3(n11836), .A4(n11835), .ZN(
        n11839) );
  OR2_X2 U15055 ( .A1(n11840), .A2(n11839), .ZN(n20172) );
  NAND2_X1 U15056 ( .A1(n20172), .A2(n11878), .ZN(n11886) );
  NAND2_X1 U15057 ( .A1(n20136), .A2(n20172), .ZN(n11880) );
  NAND2_X1 U15058 ( .A1(n11886), .A2(n11880), .ZN(n11841) );
  NAND2_X1 U15059 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11843) );
  AOI22_X1 U15060 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U15061 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11846) );
  AOI22_X1 U15062 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11845) );
  NAND4_X1 U15063 ( .A1(n11848), .A2(n11847), .A3(n11846), .A4(n11845), .ZN(
        n11854) );
  AOI22_X1 U15064 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12016), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11852) );
  AOI22_X1 U15065 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11851) );
  AOI22_X1 U15066 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12011), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11850) );
  AOI22_X1 U15067 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12017), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11849) );
  NAND4_X1 U15068 ( .A1(n11852), .A2(n11851), .A3(n11850), .A4(n11849), .ZN(
        n11853) );
  NOR2_X1 U15069 ( .A1(n11842), .A2(n20104), .ZN(n11855) );
  NAND2_X1 U15070 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11858) );
  NAND2_X1 U15071 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11857) );
  NAND2_X1 U15072 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11856) );
  NAND2_X1 U15073 ( .A1(n12115), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11863) );
  NAND2_X1 U15074 ( .A1(n11800), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11862) );
  NAND2_X1 U15075 ( .A1(n12025), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11861) );
  NAND2_X1 U15076 ( .A1(n9643), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11860) );
  NAND2_X1 U15077 ( .A1(n12026), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11867) );
  NAND2_X1 U15078 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11866) );
  NAND2_X1 U15079 ( .A1(n12011), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11865) );
  NAND2_X1 U15080 ( .A1(n12034), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11864) );
  NAND2_X1 U15081 ( .A1(n11928), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11871) );
  NAND2_X1 U15082 ( .A1(n12016), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11870) );
  NAND2_X1 U15083 ( .A1(n11929), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11869) );
  NAND2_X1 U15084 ( .A1(n12017), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11868) );
  NAND2_X1 U15085 ( .A1(n13222), .A2(n20124), .ZN(n11876) );
  NOR2_X2 U15086 ( .A1(n11906), .A2(n11876), .ZN(n11891) );
  NAND2_X1 U15087 ( .A1(n11891), .A2(n12956), .ZN(n13036) );
  NOR2_X2 U15088 ( .A1(n13036), .A2(n13619), .ZN(n12908) );
  INV_X1 U15089 ( .A(n12908), .ZN(n11881) );
  XNOR2_X1 U15090 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12953) );
  NOR2_X4 U15091 ( .A1(n20114), .A2(n20104), .ZN(n13719) );
  NAND3_X1 U15092 ( .A1(n13123), .A2(n13719), .A3(n9657), .ZN(n13132) );
  OR2_X2 U15093 ( .A1(n13216), .A2(n11882), .ZN(n11883) );
  NAND2_X2 U15094 ( .A1(n11883), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11916) );
  NAND2_X1 U15095 ( .A1(n13219), .A2(n20104), .ZN(n20898) );
  NOR2_X1 U15096 ( .A1(n11906), .A2(n11878), .ZN(n11885) );
  NAND2_X1 U15097 ( .A1(n20104), .A2(n20119), .ZN(n11887) );
  OAI211_X1 U15098 ( .C1(n13246), .C2(n20898), .A(n11905), .B(n13133), .ZN(
        n11889) );
  INV_X1 U15099 ( .A(n11889), .ZN(n11895) );
  OR2_X1 U15100 ( .A1(n11884), .A2(n11878), .ZN(n11890) );
  NAND2_X1 U15101 ( .A1(n11891), .A2(n11890), .ZN(n12958) );
  INV_X1 U15102 ( .A(n20124), .ZN(n11892) );
  INV_X1 U15103 ( .A(n13131), .ZN(n11903) );
  NAND2_X1 U15104 ( .A1(n13148), .A2(n13219), .ZN(n11893) );
  OAI21_X1 U15105 ( .B1(n11903), .B2(n11893), .A(n13619), .ZN(n11894) );
  NAND2_X2 U15106 ( .A1(n11916), .A2(n11897), .ZN(n11919) );
  NAND2_X1 U15107 ( .A1(n11919), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11899) );
  NAND2_X1 U15108 ( .A1(n20746), .A2(n20635), .ZN(n20583) );
  NAND2_X1 U15109 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20538) );
  NAND2_X1 U15110 ( .A1(n20583), .A2(n20538), .ZN(n20501) );
  NAND2_X1 U15111 ( .A1(n15652), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11917) );
  OAI21_X1 U15112 ( .B1(n13270), .B2(n20501), .A(n11917), .ZN(n11898) );
  INV_X1 U15113 ( .A(n15652), .ZN(n11900) );
  MUX2_X1 U15114 ( .A(n11900), .B(n13270), .S(n20635), .Z(n11901) );
  OAI21_X1 U15115 ( .B1(n13719), .B2(n11904), .A(n11903), .ZN(n11915) );
  AND2_X2 U15116 ( .A1(n20104), .A2(n20114), .ZN(n12652) );
  NAND2_X1 U15117 ( .A1(n11905), .A2(n12652), .ZN(n11910) );
  INV_X1 U15118 ( .A(n11906), .ZN(n11908) );
  NOR2_X1 U15119 ( .A1(n11878), .A2(n20114), .ZN(n11907) );
  AOI21_X1 U15120 ( .B1(n11908), .B2(n11907), .A(n13719), .ZN(n11909) );
  NAND2_X1 U15121 ( .A1(n11910), .A2(n11909), .ZN(n11914) );
  INV_X1 U15122 ( .A(n13133), .ZN(n11912) );
  NOR2_X1 U15123 ( .A1(n13148), .A2(n20136), .ZN(n11911) );
  INV_X1 U15124 ( .A(n16071), .ZN(n14616) );
  NOR2_X1 U15125 ( .A1(n14616), .A2(n20804), .ZN(n11913) );
  NAND4_X1 U15126 ( .A1(n11915), .A2(n11914), .A3(n13254), .A4(n11913), .ZN(
        n11959) );
  NAND2_X1 U15127 ( .A1(n11917), .A2(n12579), .ZN(n11918) );
  NAND2_X1 U15128 ( .A1(n9810), .A2(n11918), .ZN(n11924) );
  XNOR2_X1 U15129 ( .A(n20538), .B(n20419), .ZN(n20106) );
  NOR2_X1 U15130 ( .A1(n20106), .A2(n13270), .ZN(n11920) );
  NAND2_X1 U15131 ( .A1(n15652), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11923) );
  NAND2_X1 U15132 ( .A1(n11925), .A2(n11923), .ZN(n11921) );
  NAND2_X1 U15133 ( .A1(n11922), .A2(n11921), .ZN(n11967) );
  NAND4_X1 U15134 ( .A1(n11946), .A2(n11925), .A3(n11924), .A4(n11923), .ZN(
        n11926) );
  AOI22_X1 U15135 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U15136 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12090), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U15137 ( .A1(n12033), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11932) );
  AOI22_X1 U15138 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11931) );
  NAND4_X1 U15139 ( .A1(n11934), .A2(n11933), .A3(n11932), .A4(n11931), .ZN(
        n11940) );
  AOI22_X1 U15140 ( .A1(n9686), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U15141 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U15142 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11936) );
  AOI22_X1 U15143 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11935) );
  NAND4_X1 U15144 ( .A1(n11938), .A2(n11937), .A3(n11936), .A4(n11935), .ZN(
        n11939) );
  NOR2_X1 U15145 ( .A1(n20104), .A2(n20804), .ZN(n11961) );
  AOI22_X1 U15146 ( .A1(n12626), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11961), .B2(n11941), .ZN(n11942) );
  INV_X1 U15147 ( .A(n20226), .ZN(n11945) );
  INV_X1 U15148 ( .A(n11943), .ZN(n11944) );
  INV_X1 U15149 ( .A(n11963), .ZN(n11957) );
  AOI22_X1 U15150 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U15151 ( .A1(n9687), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U15152 ( .A1(n12090), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U15153 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11947) );
  NAND4_X1 U15154 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n11956) );
  AOI22_X1 U15155 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U15156 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11953) );
  AOI22_X1 U15157 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U15158 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11951) );
  NAND4_X1 U15159 ( .A1(n11954), .A2(n11953), .A3(n11952), .A4(n11951), .ZN(
        n11955) );
  NAND2_X1 U15160 ( .A1(n11957), .A2(n13233), .ZN(n11958) );
  INV_X1 U15161 ( .A(n11959), .ZN(n11960) );
  INV_X1 U15162 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11964) );
  NAND2_X1 U15163 ( .A1(n11961), .A2(n13233), .ZN(n11962) );
  OAI211_X1 U15164 ( .C1(n12621), .C2(n11964), .A(n11963), .B(n11962), .ZN(
        n11965) );
  INV_X1 U15165 ( .A(n11965), .ZN(n11966) );
  NAND2_X1 U15166 ( .A1(n12048), .A2(n11966), .ZN(n12008) );
  OAI21_X1 U15167 ( .B1(n20538), .B2(n20419), .A(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11969) );
  INV_X1 U15168 ( .A(n20538), .ZN(n20734) );
  NAND2_X1 U15169 ( .A1(n20882), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20344) );
  INV_X1 U15170 ( .A(n20344), .ZN(n11968) );
  NAND2_X1 U15171 ( .A1(n20734), .A2(n11968), .ZN(n20413) );
  NAND2_X1 U15172 ( .A1(n11969), .A2(n20413), .ZN(n20420) );
  INV_X1 U15173 ( .A(n13270), .ZN(n11970) );
  AOI22_X1 U15174 ( .A1(n20420), .A2(n11970), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n15652), .ZN(n11971) );
  AOI22_X1 U15175 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11977) );
  AOI22_X1 U15176 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12090), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11976) );
  AOI22_X1 U15177 ( .A1(n12033), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11975) );
  AOI22_X1 U15178 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11974) );
  NAND4_X1 U15179 ( .A1(n11977), .A2(n11976), .A3(n11975), .A4(n11974), .ZN(
        n11983) );
  AOI22_X1 U15180 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11981) );
  AOI22_X1 U15181 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11980) );
  AOI22_X1 U15182 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11979) );
  AOI22_X1 U15183 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11978) );
  NAND4_X1 U15184 ( .A1(n11981), .A2(n11980), .A3(n11979), .A4(n11978), .ZN(
        n11982) );
  AOI22_X1 U15185 ( .A1(n12626), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12631), .B2(n13361), .ZN(n11984) );
  NAND2_X1 U15186 ( .A1(n12626), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11997) );
  AOI22_X1 U15187 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11989) );
  AOI22_X1 U15188 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12090), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11988) );
  AOI22_X1 U15189 ( .A1(n12033), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11987) );
  AOI22_X1 U15190 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11986) );
  NAND4_X1 U15191 ( .A1(n11989), .A2(n11988), .A3(n11987), .A4(n11986), .ZN(
        n11995) );
  AOI22_X1 U15192 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11993) );
  AOI22_X1 U15193 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U15194 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U15195 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11990) );
  NAND4_X1 U15196 ( .A1(n11993), .A2(n11992), .A3(n11991), .A4(n11990), .ZN(
        n11994) );
  NAND2_X1 U15197 ( .A1(n12631), .A2(n13674), .ZN(n11996) );
  INV_X1 U15198 ( .A(n11999), .ZN(n11998) );
  AND2_X1 U15199 ( .A1(n12107), .A2(n12000), .ZN(n13360) );
  INV_X1 U15200 ( .A(n14096), .ZN(n12001) );
  INV_X1 U15201 ( .A(n12085), .ZN(n12059) );
  INV_X1 U15202 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20466) );
  OAI21_X1 U15203 ( .B1(n20466), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20383), .ZN(n12003) );
  NAND2_X1 U15204 ( .A1(n14159), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12002) );
  OAI211_X1 U15205 ( .C1(n12059), .C2(n16074), .A(n12003), .B(n12002), .ZN(
        n12006) );
  NAND2_X1 U15206 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12079) );
  NOR2_X1 U15207 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n12080), .ZN(
        n12004) );
  NOR2_X1 U15208 ( .A1(n12103), .A2(n12004), .ZN(n19954) );
  NAND2_X1 U15209 ( .A1(n19954), .A2(n13616), .ZN(n12005) );
  AND2_X1 U15210 ( .A1(n12006), .A2(n12005), .ZN(n12007) );
  AOI21_X1 U15211 ( .B1(n13360), .B2(n13021), .A(n12007), .ZN(n13398) );
  XNOR2_X1 U15212 ( .A(n13220), .B(n12009), .ZN(n13020) );
  AOI22_X1 U15213 ( .A1(n12554), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12015) );
  BUF_X1 U15214 ( .A(n12025), .Z(n12010) );
  AOI22_X1 U15215 ( .A1(n9689), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U15216 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U15217 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12012) );
  NAND4_X1 U15218 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(
        n12023) );
  AOI22_X1 U15219 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12021) );
  AOI22_X1 U15220 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12020) );
  BUF_X1 U15221 ( .A(n12016), .Z(n12090) );
  AOI22_X1 U15222 ( .A1(n12090), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U15223 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12018) );
  NAND4_X1 U15224 ( .A1(n12021), .A2(n12020), .A3(n12019), .A4(n12018), .ZN(
        n12022) );
  NAND2_X1 U15225 ( .A1(n13246), .A2(n13708), .ZN(n13700) );
  INV_X1 U15226 ( .A(n13708), .ZN(n12024) );
  NAND2_X1 U15227 ( .A1(n12024), .A2(n13246), .ZN(n12041) );
  AOI22_X1 U15228 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U15229 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12031) );
  AOI22_X1 U15230 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12030) );
  AOI22_X1 U15231 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12029) );
  NAND4_X1 U15232 ( .A1(n12032), .A2(n12031), .A3(n12030), .A4(n12029), .ZN(
        n12040) );
  AOI22_X1 U15233 ( .A1(n11930), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U15234 ( .A1(n12090), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15235 ( .A1(n9688), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U15236 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12035) );
  NAND4_X1 U15237 ( .A1(n12038), .A2(n12037), .A3(n12036), .A4(n12035), .ZN(
        n12039) );
  MUX2_X1 U15238 ( .A(n13700), .B(n12041), .S(n13232), .Z(n12042) );
  INV_X1 U15239 ( .A(n12042), .ZN(n12043) );
  NAND2_X1 U15240 ( .A1(n12043), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12050) );
  NAND2_X1 U15241 ( .A1(n12626), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12046) );
  AOI21_X1 U15242 ( .B1(n13619), .B2(n13232), .A(n20804), .ZN(n12044) );
  AND2_X1 U15243 ( .A1(n12044), .A2(n13700), .ZN(n12045) );
  NAND2_X1 U15244 ( .A1(n12046), .A2(n12045), .ZN(n12049) );
  AND2_X1 U15245 ( .A1(n12050), .A2(n12049), .ZN(n12047) );
  NAND2_X1 U15246 ( .A1(n12048), .A2(n12047), .ZN(n12054) );
  INV_X1 U15247 ( .A(n12049), .ZN(n12052) );
  INV_X1 U15248 ( .A(n12050), .ZN(n12051) );
  NAND2_X1 U15249 ( .A1(n12052), .A2(n12051), .ZN(n12053) );
  OR2_X1 U15250 ( .A1(n13227), .A2(n20136), .ZN(n12055) );
  NAND2_X1 U15251 ( .A1(n12055), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13072) );
  NAND2_X1 U15252 ( .A1(n14159), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12058) );
  NAND2_X1 U15253 ( .A1(n20383), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12057) );
  OAI211_X1 U15254 ( .C1(n12059), .C2(n14130), .A(n12058), .B(n12057), .ZN(
        n12060) );
  AOI21_X1 U15255 ( .B1(n20225), .B2(n13021), .A(n12060), .ZN(n13071) );
  INV_X1 U15256 ( .A(n13071), .ZN(n12061) );
  OR2_X1 U15257 ( .A1(n12061), .A2(n12152), .ZN(n12062) );
  NAND2_X1 U15258 ( .A1(n13074), .A2(n12062), .ZN(n13025) );
  AND2_X1 U15259 ( .A1(n13021), .A2(n13025), .ZN(n12063) );
  NAND2_X1 U15260 ( .A1(n13020), .A2(n12063), .ZN(n12068) );
  INV_X1 U15261 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n12064) );
  INV_X1 U15262 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13725) );
  OAI22_X1 U15263 ( .A1(n12078), .A2(n12064), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n13725), .ZN(n12065) );
  AOI21_X1 U15264 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n12085), .A(
        n12065), .ZN(n13022) );
  INV_X1 U15265 ( .A(n13022), .ZN(n12066) );
  NAND2_X1 U15266 ( .A1(n13025), .A2(n12066), .ZN(n12067) );
  INV_X1 U15267 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n12071) );
  INV_X2 U15268 ( .A(n12152), .ZN(n13616) );
  XNOR2_X1 U15269 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19977) );
  AOI21_X1 U15270 ( .B1(n13616), .B2(n19977), .A(n14158), .ZN(n12070) );
  OAI21_X1 U15271 ( .B1(n12078), .B2(n12071), .A(n12070), .ZN(n12072) );
  AOI21_X1 U15272 ( .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n12085), .A(
        n12072), .ZN(n12073) );
  NAND2_X1 U15273 ( .A1(n14158), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12075) );
  NAND2_X1 U15274 ( .A1(n13024), .A2(n12074), .ZN(n13087) );
  NAND2_X1 U15275 ( .A1(n12076), .A2(n20269), .ZN(n12077) );
  OR2_X1 U15276 ( .A1(n13353), .A2(n12264), .ZN(n12087) );
  INV_X1 U15277 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n13104) );
  INV_X1 U15278 ( .A(n12079), .ZN(n12082) );
  INV_X1 U15279 ( .A(n12080), .ZN(n12081) );
  OAI21_X1 U15280 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12082), .A(
        n12081), .ZN(n14113) );
  AOI22_X1 U15281 ( .A1(n13616), .A2(n14113), .B1(n14158), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12083) );
  OAI21_X1 U15282 ( .B1(n12078), .B2(n13104), .A(n12083), .ZN(n12084) );
  AOI21_X1 U15283 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12085), .A(
        n12084), .ZN(n12086) );
  NAND2_X1 U15284 ( .A1(n12087), .A2(n12086), .ZN(n13102) );
  NAND2_X1 U15285 ( .A1(n13103), .A2(n13102), .ZN(n13101) );
  INV_X1 U15286 ( .A(n13101), .ZN(n12088) );
  NAND2_X1 U15287 ( .A1(n12089), .A2(n12088), .ZN(n13392) );
  NAND2_X1 U15288 ( .A1(n12626), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12102) );
  AOI22_X1 U15289 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12094) );
  AOI22_X1 U15290 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12090), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U15291 ( .A1(n12033), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15292 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12091) );
  NAND4_X1 U15293 ( .A1(n12094), .A2(n12093), .A3(n12092), .A4(n12091), .ZN(
        n12100) );
  AOI22_X1 U15294 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U15295 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15296 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15297 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12095) );
  NAND4_X1 U15298 ( .A1(n12098), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n12099) );
  NAND2_X1 U15299 ( .A1(n12631), .A2(n13682), .ZN(n12101) );
  NAND2_X1 U15300 ( .A1(n12102), .A2(n12101), .ZN(n12108) );
  INV_X1 U15302 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n12105) );
  OAI21_X1 U15303 ( .B1(n12103), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n12124), .ZN(n19936) );
  AOI22_X1 U15304 ( .A1(n19936), .A2(n13616), .B1(n14158), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12104) );
  OAI21_X1 U15305 ( .B1(n12078), .B2(n12105), .A(n12104), .ZN(n12106) );
  NAND2_X1 U15306 ( .A1(n12626), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12123) );
  NAND2_X1 U15307 ( .A1(n11820), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12110) );
  AND2_X1 U15308 ( .A1(n12110), .A2(n12109), .ZN(n12114) );
  AOI22_X1 U15309 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12113) );
  AOI22_X1 U15310 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U15311 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12111) );
  NAND4_X1 U15312 ( .A1(n12114), .A2(n12113), .A3(n12112), .A4(n12111), .ZN(
        n12121) );
  AOI22_X1 U15313 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n9679), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12119) );
  AOI22_X1 U15314 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12090), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12118) );
  AOI22_X1 U15315 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12117) );
  AOI22_X1 U15316 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12116) );
  NAND4_X1 U15317 ( .A1(n12119), .A2(n12118), .A3(n12117), .A4(n12116), .ZN(
        n12120) );
  NAND2_X1 U15318 ( .A1(n12631), .A2(n13692), .ZN(n12122) );
  NAND2_X1 U15319 ( .A1(n12131), .A2(n12132), .ZN(n13681) );
  NAND2_X1 U15320 ( .A1(n13681), .A2(n13021), .ZN(n12130) );
  AND2_X1 U15321 ( .A1(n12124), .A2(n12127), .ZN(n12125) );
  OR2_X1 U15322 ( .A1(n12125), .A2(n12137), .ZN(n19922) );
  NAND2_X1 U15323 ( .A1(n19922), .A2(n13616), .ZN(n12126) );
  OAI21_X1 U15324 ( .B1(n12127), .B2(n12300), .A(n12126), .ZN(n12128) );
  AOI21_X1 U15325 ( .B1(n14159), .B2(P1_EAX_REG_6__SCAN_IN), .A(n12128), .ZN(
        n12129) );
  NAND2_X1 U15326 ( .A1(n13394), .A2(n13416), .ZN(n13415) );
  INV_X1 U15327 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12135) );
  NAND2_X1 U15328 ( .A1(n12631), .A2(n13708), .ZN(n12134) );
  OAI21_X1 U15329 ( .B1(n12621), .B2(n12135), .A(n12134), .ZN(n12136) );
  INV_X1 U15330 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13514) );
  NOR2_X1 U15331 ( .A1(n12137), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12138) );
  OR2_X1 U15332 ( .A1(n12156), .A2(n12138), .ZN(n19909) );
  AOI22_X1 U15333 ( .A1(n19909), .A2(n13616), .B1(n14158), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12139) );
  OAI21_X1 U15334 ( .B1(n12078), .B2(n13514), .A(n12139), .ZN(n12140) );
  AOI21_X1 U15335 ( .B1(n13691), .B2(n13021), .A(n12140), .ZN(n13512) );
  INV_X1 U15336 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13646) );
  INV_X1 U15337 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12151) );
  OAI22_X1 U15338 ( .A1(n12078), .A2(n13646), .B1(n12300), .B2(n12151), .ZN(
        n12155) );
  AOI22_X1 U15339 ( .A1(n12554), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U15340 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n9643), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U15341 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12142) );
  AOI22_X1 U15342 ( .A1(n12090), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12141) );
  NAND4_X1 U15343 ( .A1(n12144), .A2(n12143), .A3(n12142), .A4(n12141), .ZN(
        n12150) );
  AOI22_X1 U15344 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12148) );
  AOI22_X1 U15345 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12147) );
  AOI22_X1 U15346 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15347 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12145) );
  NAND4_X1 U15348 ( .A1(n12148), .A2(n12147), .A3(n12146), .A4(n12145), .ZN(
        n12149) );
  NOR2_X1 U15349 ( .A1(n12150), .A2(n12149), .ZN(n12153) );
  XNOR2_X1 U15350 ( .A(n12156), .B(n12151), .ZN(n13712) );
  OAI22_X1 U15351 ( .A1(n12264), .A2(n12153), .B1(n13712), .B2(n12152), .ZN(
        n12154) );
  NOR2_X1 U15352 ( .A1(n12155), .A2(n12154), .ZN(n13611) );
  XOR2_X1 U15353 ( .A(n19899), .B(n12173), .Z(n19902) );
  INV_X1 U15354 ( .A(n19902), .ZN(n12171) );
  NAND2_X1 U15355 ( .A1(n14159), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15356 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12360), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U15357 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15358 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12158) );
  AOI22_X1 U15359 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12157) );
  NAND4_X1 U15360 ( .A1(n12160), .A2(n12159), .A3(n12158), .A4(n12157), .ZN(
        n12166) );
  AOI22_X1 U15361 ( .A1(n12554), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15362 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15363 ( .A1(n12090), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12162) );
  AOI22_X1 U15364 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12161) );
  NAND4_X1 U15365 ( .A1(n12164), .A2(n12163), .A3(n12162), .A4(n12161), .ZN(
        n12165) );
  OAI21_X1 U15366 ( .B1(n12166), .B2(n12165), .A(n13021), .ZN(n12168) );
  NAND2_X1 U15367 ( .A1(n14158), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12167) );
  NAND3_X1 U15368 ( .A1(n12169), .A2(n12168), .A3(n12167), .ZN(n12170) );
  XNOR2_X1 U15369 ( .A(n12190), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14512) );
  NAND2_X1 U15370 ( .A1(n14512), .A2(n13616), .ZN(n12189) );
  INV_X1 U15371 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13804) );
  INV_X1 U15372 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12174) );
  OAI22_X1 U15373 ( .A1(n12078), .A2(n13804), .B1(n12300), .B2(n12174), .ZN(
        n12187) );
  AOI22_X1 U15374 ( .A1(n12554), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15375 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U15376 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12471), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U15377 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12175) );
  NAND4_X1 U15378 ( .A1(n12178), .A2(n12177), .A3(n12176), .A4(n12175), .ZN(
        n12184) );
  AOI22_X1 U15379 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12182) );
  AOI22_X1 U15380 ( .A1(n12090), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12181) );
  AOI22_X1 U15381 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15382 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12179) );
  NAND4_X1 U15383 ( .A1(n12182), .A2(n12181), .A3(n12180), .A4(n12179), .ZN(
        n12183) );
  NOR2_X1 U15384 ( .A1(n12184), .A2(n12183), .ZN(n12185) );
  NOR2_X1 U15385 ( .A1(n12264), .A2(n12185), .ZN(n12186) );
  NOR2_X1 U15386 ( .A1(n12187), .A2(n12186), .ZN(n12188) );
  NAND2_X1 U15387 ( .A1(n12189), .A2(n12188), .ZN(n13763) );
  INV_X1 U15388 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n13892) );
  OAI21_X1 U15389 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12191), .A(
        n12229), .ZN(n15899) );
  AOI22_X1 U15390 ( .A1(n13616), .A2(n15899), .B1(n14158), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12192) );
  OAI21_X1 U15391 ( .B1(n12078), .B2(n13892), .A(n12192), .ZN(n13887) );
  AOI22_X1 U15392 ( .A1(n12554), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12196) );
  AOI22_X1 U15393 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15394 ( .A1(n12090), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15395 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12193) );
  NAND4_X1 U15396 ( .A1(n12196), .A2(n12195), .A3(n12194), .A4(n12193), .ZN(
        n12202) );
  AOI22_X1 U15397 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12200) );
  AOI22_X1 U15398 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15399 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15400 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12197) );
  NAND4_X1 U15401 ( .A1(n12200), .A2(n12199), .A3(n12198), .A4(n12197), .ZN(
        n12201) );
  NOR2_X1 U15402 ( .A1(n12202), .A2(n12201), .ZN(n12203) );
  NOR2_X1 U15403 ( .A1(n12264), .A2(n12203), .ZN(n13951) );
  XOR2_X1 U15404 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12233), .Z(
        n14501) );
  AOI22_X1 U15405 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15406 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15407 ( .A1(n12090), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U15408 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12204) );
  NAND4_X1 U15409 ( .A1(n12207), .A2(n12206), .A3(n12205), .A4(n12204), .ZN(
        n12213) );
  AOI22_X1 U15410 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n9679), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U15411 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15412 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12034), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12209) );
  AOI22_X1 U15413 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12208) );
  NAND4_X1 U15414 ( .A1(n12211), .A2(n12210), .A3(n12209), .A4(n12208), .ZN(
        n12212) );
  NOR2_X1 U15415 ( .A1(n12213), .A2(n12212), .ZN(n12214) );
  INV_X1 U15416 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14499) );
  OAI22_X1 U15417 ( .A1(n12264), .A2(n12214), .B1(n12300), .B2(n14499), .ZN(
        n12216) );
  INV_X1 U15418 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14065) );
  NOR2_X1 U15419 ( .A1(n12078), .A2(n14065), .ZN(n12215) );
  NOR2_X1 U15420 ( .A1(n12216), .A2(n12215), .ZN(n12217) );
  OAI21_X1 U15421 ( .B1(n14501), .B2(n12152), .A(n12217), .ZN(n13991) );
  INV_X1 U15422 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n13967) );
  AOI22_X1 U15423 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12221) );
  AOI22_X1 U15424 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(n9643), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12220) );
  AOI22_X1 U15425 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12219) );
  AOI22_X1 U15426 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12218) );
  NAND4_X1 U15427 ( .A1(n12221), .A2(n12220), .A3(n12219), .A4(n12218), .ZN(
        n12227) );
  AOI22_X1 U15428 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12225) );
  AOI22_X1 U15429 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12090), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15430 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15431 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12222) );
  NAND4_X1 U15432 ( .A1(n12225), .A2(n12224), .A3(n12223), .A4(n12222), .ZN(
        n12226) );
  OR2_X1 U15433 ( .A1(n12227), .A2(n12226), .ZN(n12228) );
  NAND2_X1 U15434 ( .A1(n13021), .A2(n12228), .ZN(n12232) );
  XOR2_X1 U15435 ( .A(n15805), .B(n12229), .Z(n15888) );
  INV_X1 U15436 ( .A(n15888), .ZN(n12230) );
  AOI22_X1 U15437 ( .A1(n14158), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13616), .B2(n12230), .ZN(n12231) );
  OAI211_X1 U15438 ( .C1(n13967), .C2(n12078), .A(n12232), .B(n12231), .ZN(
        n13954) );
  XNOR2_X1 U15439 ( .A(n12250), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14280) );
  INV_X1 U15440 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15441 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U15442 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n12090), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12236) );
  AOI22_X1 U15443 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n9666), .B1(
        n12360), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U15444 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n12561), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12234) );
  NAND4_X1 U15445 ( .A1(n12237), .A2(n12236), .A3(n12235), .A4(n12234), .ZN(
        n12243) );
  AOI22_X1 U15446 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(n9644), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12240) );
  AOI22_X1 U15447 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12495), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U15448 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n12471), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12238) );
  NAND4_X1 U15449 ( .A1(n12241), .A2(n12240), .A3(n12239), .A4(n12238), .ZN(
        n12242) );
  OAI21_X1 U15450 ( .B1(n12243), .B2(n12242), .A(n13021), .ZN(n12245) );
  NAND2_X1 U15451 ( .A1(n14159), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12244) );
  OAI211_X1 U15452 ( .C1(n12300), .C2(n12246), .A(n12245), .B(n12244), .ZN(
        n12247) );
  AOI21_X1 U15453 ( .B1(n14280), .B2(n13616), .A(n12247), .ZN(n13963) );
  AOI21_X1 U15454 ( .B1(n20934), .B2(n12251), .A(n12289), .ZN(n15878) );
  OR2_X1 U15455 ( .A1(n15878), .A2(n12152), .ZN(n12269) );
  AOI22_X1 U15456 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U15457 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U15458 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15459 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12252) );
  NAND4_X1 U15460 ( .A1(n12255), .A2(n12254), .A3(n12253), .A4(n12252), .ZN(
        n12262) );
  AOI22_X1 U15461 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12260) );
  AOI22_X1 U15462 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(n9644), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12259) );
  AOI22_X1 U15463 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12258) );
  AOI22_X1 U15464 ( .A1(n12016), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12257) );
  NAND4_X1 U15465 ( .A1(n12260), .A2(n12259), .A3(n12258), .A4(n12257), .ZN(
        n12261) );
  NOR2_X1 U15466 ( .A1(n12262), .A2(n12261), .ZN(n12263) );
  OAI22_X1 U15467 ( .A1(n12264), .A2(n12263), .B1(n12300), .B2(n20934), .ZN(
        n12267) );
  INV_X1 U15468 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n12265) );
  NOR2_X1 U15469 ( .A1(n12078), .A2(n12265), .ZN(n12266) );
  NOR2_X1 U15470 ( .A1(n12267), .A2(n12266), .ZN(n12268) );
  INV_X1 U15471 ( .A(n14070), .ZN(n12270) );
  INV_X1 U15472 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12271) );
  XNOR2_X1 U15473 ( .A(n12289), .B(n12271), .ZN(n15792) );
  NAND2_X1 U15474 ( .A1(n15792), .A2(n13616), .ZN(n12288) );
  AOI22_X1 U15475 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12495), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U15476 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12471), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12274) );
  AOI22_X1 U15477 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15478 ( .A1(n12256), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12272) );
  NAND4_X1 U15479 ( .A1(n12275), .A2(n12274), .A3(n12273), .A4(n12272), .ZN(
        n12283) );
  AOI22_X1 U15480 ( .A1(n12025), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12281) );
  AOI21_X1 U15481 ( .B1(n9644), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A(n13616), .ZN(n12276) );
  AND2_X1 U15482 ( .A1(n12277), .A2(n12276), .ZN(n12280) );
  AOI22_X1 U15483 ( .A1(n12016), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12279) );
  AOI22_X1 U15484 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12278) );
  NAND4_X1 U15485 ( .A1(n12281), .A2(n12280), .A3(n12279), .A4(n12278), .ZN(
        n12282) );
  NAND2_X1 U15486 ( .A1(n12549), .A2(n12152), .ZN(n12392) );
  OAI21_X1 U15487 ( .B1(n12283), .B2(n12282), .A(n12392), .ZN(n12286) );
  NAND2_X1 U15488 ( .A1(n14159), .A2(P1_EAX_REG_16__SCAN_IN), .ZN(n12285) );
  NAND2_X1 U15489 ( .A1(n20383), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12284) );
  NAND3_X1 U15490 ( .A1(n12286), .A2(n12285), .A3(n12284), .ZN(n12287) );
  NAND2_X1 U15491 ( .A1(n12288), .A2(n12287), .ZN(n14349) );
  XOR2_X1 U15492 ( .A(n12305), .B(n12306), .Z(n15867) );
  INV_X1 U15493 ( .A(n12549), .ZN(n12570) );
  AOI22_X1 U15494 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12293) );
  AOI22_X1 U15495 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12292) );
  AOI22_X1 U15496 ( .A1(n12090), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U15497 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12290) );
  NAND4_X1 U15498 ( .A1(n12293), .A2(n12292), .A3(n12291), .A4(n12290), .ZN(
        n12299) );
  AOI22_X1 U15499 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(n9679), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15500 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12296) );
  AOI22_X1 U15501 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U15502 ( .A1(n12561), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12294) );
  NAND4_X1 U15503 ( .A1(n12297), .A2(n12296), .A3(n12295), .A4(n12294), .ZN(
        n12298) );
  OR2_X1 U15504 ( .A1(n12299), .A2(n12298), .ZN(n12303) );
  INV_X1 U15505 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n12301) );
  OAI22_X1 U15506 ( .A1(n12078), .A2(n12301), .B1(n12300), .B2(n12305), .ZN(
        n12302) );
  AOI21_X1 U15507 ( .B1(n12570), .B2(n12303), .A(n12302), .ZN(n12304) );
  OAI21_X1 U15508 ( .B1(n15867), .B2(n12152), .A(n12304), .ZN(n14266) );
  INV_X1 U15509 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14478) );
  XNOR2_X1 U15510 ( .A(n12339), .B(n14478), .ZN(n14480) );
  NAND2_X1 U15511 ( .A1(n14480), .A2(n13616), .ZN(n12323) );
  AOI22_X1 U15512 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12016), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U15513 ( .A1(n9666), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15514 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U15515 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12307) );
  NAND4_X1 U15516 ( .A1(n12310), .A2(n12309), .A3(n12308), .A4(n12307), .ZN(
        n12318) );
  AOI21_X1 U15517 ( .B1(n12010), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n13616), .ZN(n12312) );
  AND2_X1 U15518 ( .A1(n12312), .A2(n12311), .ZN(n12316) );
  AOI22_X1 U15519 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12315) );
  AOI22_X1 U15520 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12360), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U15521 ( .A1(n12033), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12313) );
  NAND4_X1 U15522 ( .A1(n12316), .A2(n12315), .A3(n12314), .A4(n12313), .ZN(
        n12317) );
  OAI21_X1 U15523 ( .B1(n12318), .B2(n12317), .A(n12392), .ZN(n12321) );
  NAND2_X1 U15524 ( .A1(n14159), .A2(P1_EAX_REG_18__SCAN_IN), .ZN(n12320) );
  NAND2_X1 U15525 ( .A1(n20383), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12319) );
  NAND3_X1 U15526 ( .A1(n12321), .A2(n12320), .A3(n12319), .ZN(n12322) );
  AOI22_X1 U15527 ( .A1(n12554), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15528 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12326) );
  AOI22_X1 U15529 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12325) );
  AOI22_X1 U15530 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12324) );
  NAND4_X1 U15531 ( .A1(n12327), .A2(n12326), .A3(n12325), .A4(n12324), .ZN(
        n12333) );
  AOI22_X1 U15532 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12331) );
  AOI22_X1 U15533 ( .A1(n12090), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12330) );
  AOI22_X1 U15534 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U15535 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12328) );
  NAND4_X1 U15536 ( .A1(n12331), .A2(n12330), .A3(n12329), .A4(n12328), .ZN(
        n12332) );
  NOR2_X1 U15537 ( .A1(n12333), .A2(n12332), .ZN(n12338) );
  INV_X1 U15538 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n12335) );
  NAND2_X1 U15539 ( .A1(n20383), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12334) );
  OAI211_X1 U15540 ( .C1(n12078), .C2(n12335), .A(n12152), .B(n12334), .ZN(
        n12336) );
  INV_X1 U15541 ( .A(n12336), .ZN(n12337) );
  OAI21_X1 U15542 ( .B1(n12549), .B2(n12338), .A(n12337), .ZN(n12342) );
  OAI21_X1 U15543 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n12340), .A(
        n12374), .ZN(n15860) );
  OR2_X1 U15544 ( .A1(n12152), .A2(n15860), .ZN(n12341) );
  NAND2_X1 U15545 ( .A1(n12342), .A2(n12341), .ZN(n14339) );
  AOI21_X1 U15546 ( .B1(n12025), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n13616), .ZN(n12344) );
  AND2_X1 U15547 ( .A1(n12344), .A2(n12343), .ZN(n12348) );
  AOI22_X1 U15548 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U15549 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U15550 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12345) );
  NAND4_X1 U15551 ( .A1(n12348), .A2(n12347), .A3(n12346), .A4(n12345), .ZN(
        n12354) );
  AOI22_X1 U15552 ( .A1(n12090), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12360), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U15553 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U15554 ( .A1(n12561), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12350) );
  AOI22_X1 U15555 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12349) );
  NAND4_X1 U15556 ( .A1(n12352), .A2(n12351), .A3(n12350), .A4(n12349), .ZN(
        n12353) );
  OR2_X1 U15557 ( .A1(n12354), .A2(n12353), .ZN(n12355) );
  NAND2_X1 U15558 ( .A1(n12392), .A2(n12355), .ZN(n12359) );
  INV_X1 U15559 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n14384) );
  OAI22_X1 U15560 ( .A1(n12078), .A2(n14384), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n15774), .ZN(n12356) );
  INV_X1 U15561 ( .A(n12356), .ZN(n12358) );
  XNOR2_X1 U15562 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n12374), .ZN(
        n15764) );
  AOI21_X1 U15563 ( .B1(n12359), .B2(n12358), .A(n12357), .ZN(n14335) );
  AOI22_X1 U15564 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12364) );
  AOI22_X1 U15565 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12363) );
  AOI22_X1 U15566 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12471), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U15567 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12361) );
  NAND4_X1 U15568 ( .A1(n12364), .A2(n12363), .A3(n12362), .A4(n12361), .ZN(
        n12370) );
  AOI22_X1 U15569 ( .A1(n12010), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12368) );
  AOI22_X1 U15570 ( .A1(n12016), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12367) );
  AOI22_X1 U15571 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12366) );
  AOI22_X1 U15572 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12365) );
  NAND4_X1 U15573 ( .A1(n12368), .A2(n12367), .A3(n12366), .A4(n12365), .ZN(
        n12369) );
  NOR2_X1 U15574 ( .A1(n12370), .A2(n12369), .ZN(n12371) );
  OR2_X1 U15575 ( .A1(n12549), .A2(n12371), .ZN(n12378) );
  INV_X1 U15576 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n14379) );
  NAND2_X1 U15577 ( .A1(n20383), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12372) );
  OAI211_X1 U15578 ( .C1(n12078), .C2(n14379), .A(n12152), .B(n12372), .ZN(
        n12373) );
  INV_X1 U15579 ( .A(n12373), .ZN(n12377) );
  OAI21_X1 U15580 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n12375), .A(
        n12426), .ZN(n15845) );
  NOR2_X1 U15581 ( .A1(n15845), .A2(n12152), .ZN(n12376) );
  AOI21_X1 U15582 ( .B1(n12378), .B2(n12377), .A(n12376), .ZN(n14377) );
  NAND2_X1 U15583 ( .A1(n14334), .A2(n14377), .ZN(n14325) );
  AOI22_X1 U15584 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9679), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12382) );
  AOI22_X1 U15585 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15586 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12027), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12380) );
  AOI22_X1 U15587 ( .A1(n9665), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12379) );
  NAND4_X1 U15588 ( .A1(n12382), .A2(n12381), .A3(n12380), .A4(n12379), .ZN(
        n12390) );
  NAND2_X1 U15589 ( .A1(n12470), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n12384) );
  AOI21_X1 U15590 ( .B1(n9643), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A(n13616), .ZN(n12383) );
  AND2_X1 U15591 ( .A1(n12384), .A2(n12383), .ZN(n12388) );
  AOI22_X1 U15592 ( .A1(n12554), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12360), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12387) );
  AOI22_X1 U15593 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12386) );
  AOI22_X1 U15594 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n12090), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12385) );
  NAND4_X1 U15595 ( .A1(n12388), .A2(n12387), .A3(n12386), .A4(n12385), .ZN(
        n12389) );
  OR2_X1 U15596 ( .A1(n12390), .A2(n12389), .ZN(n12391) );
  NAND2_X1 U15597 ( .A1(n12392), .A2(n12391), .ZN(n12396) );
  INV_X1 U15598 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n12393) );
  OAI22_X1 U15599 ( .A1(n12078), .A2(n12393), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n14464), .ZN(n12394) );
  INV_X1 U15600 ( .A(n12394), .ZN(n12395) );
  NAND2_X1 U15601 ( .A1(n12396), .A2(n12395), .ZN(n12398) );
  XNOR2_X1 U15602 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n12426), .ZN(
        n15747) );
  NAND2_X1 U15603 ( .A1(n15747), .A2(n13616), .ZN(n12397) );
  NAND2_X1 U15604 ( .A1(n12398), .A2(n12397), .ZN(n14326) );
  AOI22_X1 U15605 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12404) );
  AOI22_X1 U15606 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12403) );
  AOI22_X1 U15607 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12402) );
  AOI22_X1 U15608 ( .A1(n12090), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12401) );
  NAND4_X1 U15609 ( .A1(n12404), .A2(n12403), .A3(n12402), .A4(n12401), .ZN(
        n12410) );
  AOI22_X1 U15610 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12033), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12408) );
  AOI22_X1 U15611 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12407) );
  AOI22_X1 U15612 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12406) );
  AOI22_X1 U15613 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9643), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12405) );
  NAND4_X1 U15614 ( .A1(n12408), .A2(n12407), .A3(n12406), .A4(n12405), .ZN(
        n12409) );
  NOR2_X1 U15615 ( .A1(n12410), .A2(n12409), .ZN(n12430) );
  AOI22_X1 U15616 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U15617 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U15618 ( .A1(n12090), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12412) );
  AOI22_X1 U15619 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12411) );
  NAND4_X1 U15620 ( .A1(n12414), .A2(n12413), .A3(n12412), .A4(n12411), .ZN(
        n12420) );
  AOI22_X1 U15621 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9642), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12418) );
  AOI22_X1 U15622 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U15623 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9672), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U15624 ( .A1(n12033), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12415) );
  NAND4_X1 U15625 ( .A1(n12418), .A2(n12417), .A3(n12416), .A4(n12415), .ZN(
        n12419) );
  NOR2_X1 U15626 ( .A1(n12420), .A2(n12419), .ZN(n12431) );
  XNOR2_X1 U15627 ( .A(n12430), .B(n12431), .ZN(n12425) );
  INV_X1 U15628 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n12422) );
  NAND2_X1 U15629 ( .A1(n20383), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12421) );
  OAI211_X1 U15630 ( .C1(n12078), .C2(n12422), .A(n12152), .B(n12421), .ZN(
        n12423) );
  INV_X1 U15631 ( .A(n12423), .ZN(n12424) );
  OAI21_X1 U15632 ( .B1(n12549), .B2(n12425), .A(n12424), .ZN(n12429) );
  OAI21_X1 U15633 ( .B1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n12427), .A(
        n12464), .ZN(n15843) );
  OR2_X1 U15634 ( .A1(n12152), .A2(n15843), .ZN(n12428) );
  NAND2_X1 U15635 ( .A1(n12429), .A2(n12428), .ZN(n14319) );
  NOR2_X1 U15636 ( .A1(n12431), .A2(n12430), .ZN(n12448) );
  AOI22_X1 U15637 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12435) );
  AOI22_X1 U15638 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12016), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12434) );
  AOI22_X1 U15639 ( .A1(n12033), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12433) );
  AOI22_X1 U15640 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12432) );
  NAND4_X1 U15641 ( .A1(n12435), .A2(n12434), .A3(n12433), .A4(n12432), .ZN(
        n12441) );
  AOI22_X1 U15642 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12439) );
  AOI22_X1 U15643 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15644 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U15645 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12436) );
  NAND4_X1 U15646 ( .A1(n12439), .A2(n12438), .A3(n12437), .A4(n12436), .ZN(
        n12440) );
  OR2_X1 U15647 ( .A1(n12441), .A2(n12440), .ZN(n12447) );
  XNOR2_X1 U15648 ( .A(n12448), .B(n12447), .ZN(n12444) );
  NAND2_X1 U15649 ( .A1(n14159), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n12443) );
  OAI21_X1 U15650 ( .B1(n20466), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n20383), .ZN(n12442) );
  OAI211_X1 U15651 ( .C1(n12444), .C2(n12549), .A(n12443), .B(n12442), .ZN(
        n12446) );
  XNOR2_X1 U15652 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B(n12464), .ZN(
        n15726) );
  NAND2_X1 U15653 ( .A1(n15726), .A2(n13616), .ZN(n12445) );
  NAND2_X1 U15654 ( .A1(n12448), .A2(n12447), .ZN(n12468) );
  AOI22_X1 U15655 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12452) );
  AOI22_X1 U15656 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12451) );
  AOI22_X1 U15657 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12450) );
  AOI22_X1 U15658 ( .A1(n12033), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12449) );
  NAND4_X1 U15659 ( .A1(n12452), .A2(n12451), .A3(n12450), .A4(n12449), .ZN(
        n12458) );
  AOI22_X1 U15660 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12090), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12456) );
  AOI22_X1 U15661 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U15662 ( .A1(n12025), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12454) );
  AOI22_X1 U15663 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12453) );
  NAND4_X1 U15664 ( .A1(n12456), .A2(n12455), .A3(n12454), .A4(n12453), .ZN(
        n12457) );
  NOR2_X1 U15665 ( .A1(n12458), .A2(n12457), .ZN(n12469) );
  XNOR2_X1 U15666 ( .A(n12468), .B(n12469), .ZN(n12463) );
  INV_X1 U15667 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12460) );
  NAND2_X1 U15668 ( .A1(n20383), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12459) );
  OAI211_X1 U15669 ( .C1(n12078), .C2(n12460), .A(n12152), .B(n12459), .ZN(
        n12461) );
  INV_X1 U15670 ( .A(n12461), .ZN(n12462) );
  OAI21_X1 U15671 ( .B1(n12463), .B2(n12549), .A(n12462), .ZN(n12467) );
  INV_X1 U15672 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15728) );
  OAI21_X1 U15673 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n12465), .A(
        n12505), .ZN(n15830) );
  OR2_X1 U15674 ( .A1(n15830), .A2(n12152), .ZN(n12466) );
  NOR2_X1 U15675 ( .A1(n12469), .A2(n12468), .ZN(n12490) );
  AOI22_X1 U15676 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U15677 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12090), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12474) );
  AOI22_X1 U15678 ( .A1(n12033), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12473) );
  AOI22_X1 U15679 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12472) );
  NAND4_X1 U15680 ( .A1(n12475), .A2(n12474), .A3(n12473), .A4(n12472), .ZN(
        n12481) );
  AOI22_X1 U15681 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12479) );
  AOI22_X1 U15682 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12478) );
  AOI22_X1 U15683 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U15684 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12476) );
  NAND4_X1 U15685 ( .A1(n12479), .A2(n12478), .A3(n12477), .A4(n12476), .ZN(
        n12480) );
  OR2_X1 U15686 ( .A1(n12481), .A2(n12480), .ZN(n12489) );
  XNOR2_X1 U15687 ( .A(n12490), .B(n12489), .ZN(n12486) );
  INV_X1 U15688 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n12483) );
  NAND2_X1 U15689 ( .A1(n20383), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12482) );
  OAI211_X1 U15690 ( .C1(n12078), .C2(n12483), .A(n12152), .B(n12482), .ZN(
        n12484) );
  INV_X1 U15691 ( .A(n12484), .ZN(n12485) );
  OAI21_X1 U15692 ( .B1(n12486), .B2(n12549), .A(n12485), .ZN(n12488) );
  XNOR2_X1 U15693 ( .A(n12505), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14446) );
  NAND2_X1 U15694 ( .A1(n14446), .A2(n13616), .ZN(n12487) );
  NAND2_X1 U15695 ( .A1(n12490), .A2(n12489), .ZN(n12525) );
  AOI22_X1 U15696 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12494) );
  AOI22_X1 U15697 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12493) );
  AOI22_X1 U15698 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12492) );
  AOI22_X1 U15699 ( .A1(n12033), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12491) );
  NAND4_X1 U15700 ( .A1(n12494), .A2(n12493), .A3(n12492), .A4(n12491), .ZN(
        n12501) );
  AOI22_X1 U15701 ( .A1(n12495), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12016), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12499) );
  AOI22_X1 U15702 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12498) );
  AOI22_X1 U15703 ( .A1(n9644), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12497) );
  AOI22_X1 U15704 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12496) );
  NAND4_X1 U15705 ( .A1(n12499), .A2(n12498), .A3(n12497), .A4(n12496), .ZN(
        n12500) );
  NOR2_X1 U15706 ( .A1(n12501), .A2(n12500), .ZN(n12526) );
  XNOR2_X1 U15707 ( .A(n12525), .B(n12526), .ZN(n12504) );
  OAI21_X1 U15708 ( .B1(n20466), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n20383), .ZN(n12503) );
  NAND2_X1 U15709 ( .A1(n14159), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n12502) );
  OAI211_X1 U15710 ( .C1(n12504), .C2(n12549), .A(n12503), .B(n12502), .ZN(
        n12512) );
  INV_X1 U15711 ( .A(n12505), .ZN(n12506) );
  INV_X1 U15712 ( .A(n12507), .ZN(n12509) );
  INV_X1 U15713 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12508) );
  NAND2_X1 U15714 ( .A1(n12509), .A2(n12508), .ZN(n12510) );
  NAND2_X1 U15715 ( .A1(n14438), .A2(n13616), .ZN(n12511) );
  INV_X1 U15716 ( .A(n14235), .ZN(n12513) );
  AOI22_X1 U15717 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12518) );
  AOI22_X1 U15718 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12090), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12517) );
  AOI22_X1 U15719 ( .A1(n12033), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12516) );
  AOI22_X1 U15720 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9666), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12515) );
  NAND4_X1 U15721 ( .A1(n12518), .A2(n12517), .A3(n12516), .A4(n12515), .ZN(
        n12524) );
  AOI22_X1 U15722 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12010), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12522) );
  AOI22_X1 U15723 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12521) );
  AOI22_X1 U15724 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12520) );
  AOI22_X1 U15725 ( .A1(n12027), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12519) );
  NAND4_X1 U15726 ( .A1(n12522), .A2(n12521), .A3(n12520), .A4(n12519), .ZN(
        n12523) );
  OR2_X1 U15727 ( .A1(n12524), .A2(n12523), .ZN(n12535) );
  NOR2_X1 U15728 ( .A1(n12526), .A2(n12525), .ZN(n12536) );
  XOR2_X1 U15729 ( .A(n12535), .B(n12536), .Z(n12527) );
  NAND2_X1 U15730 ( .A1(n12527), .A2(n12570), .ZN(n12530) );
  INV_X1 U15731 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14430) );
  NOR2_X1 U15732 ( .A1(n14430), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12528) );
  AOI211_X1 U15733 ( .C1(n14159), .C2(P1_EAX_REG_28__SCAN_IN), .A(n13616), .B(
        n12528), .ZN(n12529) );
  XNOR2_X1 U15734 ( .A(n12531), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14434) );
  AOI22_X1 U15735 ( .A1(n12530), .A2(n12529), .B1(n13616), .B2(n14434), .ZN(
        n14094) );
  INV_X1 U15736 ( .A(n12531), .ZN(n12532) );
  NAND2_X1 U15737 ( .A1(n12532), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12533) );
  INV_X1 U15738 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14226) );
  NAND2_X1 U15739 ( .A1(n12533), .A2(n14226), .ZN(n12534) );
  NAND2_X1 U15740 ( .A1(n13624), .A2(n12534), .ZN(n14420) );
  NAND2_X1 U15741 ( .A1(n12536), .A2(n12535), .ZN(n12552) );
  AOI22_X1 U15742 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12514), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12540) );
  AOI22_X1 U15743 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9643), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12539) );
  AOI22_X1 U15744 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n12027), .B1(
        n12025), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12538) );
  AOI22_X1 U15745 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n9666), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12537) );
  NAND4_X1 U15746 ( .A1(n12540), .A2(n12539), .A3(n12538), .A4(n12537), .ZN(
        n12546) );
  AOI22_X1 U15747 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12016), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12544) );
  AOI22_X1 U15748 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n12033), .B1(
        n12360), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U15749 ( .A1(n9684), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12542) );
  AOI22_X1 U15750 ( .A1(n12471), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12541) );
  NAND4_X1 U15751 ( .A1(n12544), .A2(n12543), .A3(n12542), .A4(n12541), .ZN(
        n12545) );
  NOR2_X1 U15752 ( .A1(n12546), .A2(n12545), .ZN(n12553) );
  XNOR2_X1 U15753 ( .A(n12552), .B(n12553), .ZN(n12550) );
  AOI21_X1 U15754 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20383), .A(
        n13616), .ZN(n12548) );
  NAND2_X1 U15755 ( .A1(n14159), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12547) );
  OAI211_X1 U15756 ( .C1(n12550), .C2(n12549), .A(n12548), .B(n12547), .ZN(
        n12551) );
  OAI21_X1 U15757 ( .B1(n12152), .B2(n14420), .A(n12551), .ZN(n14223) );
  NOR2_X1 U15758 ( .A1(n12553), .A2(n12552), .ZN(n12569) );
  AOI22_X1 U15759 ( .A1(n12554), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12470), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12559) );
  AOI22_X1 U15760 ( .A1(n9679), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12027), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12558) );
  AOI22_X1 U15761 ( .A1(n12028), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12471), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U15762 ( .A1(n12033), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12555), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12556) );
  NAND4_X1 U15763 ( .A1(n12559), .A2(n12558), .A3(n12557), .A4(n12556), .ZN(
        n12567) );
  AOI22_X1 U15764 ( .A1(n12360), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9665), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12565) );
  AOI22_X1 U15765 ( .A1(n12016), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12561), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U15766 ( .A1(n12025), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9644), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12563) );
  AOI22_X1 U15767 ( .A1(n9685), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12256), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12562) );
  NAND4_X1 U15768 ( .A1(n12565), .A2(n12564), .A3(n12563), .A4(n12562), .ZN(
        n12566) );
  NOR2_X1 U15769 ( .A1(n12567), .A2(n12566), .ZN(n12568) );
  XNOR2_X1 U15770 ( .A(n12569), .B(n12568), .ZN(n12571) );
  NAND2_X1 U15771 ( .A1(n12571), .A2(n12570), .ZN(n12577) );
  INV_X1 U15772 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n12573) );
  NAND2_X1 U15773 ( .A1(n20383), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12572) );
  OAI211_X1 U15774 ( .C1(n12078), .C2(n12573), .A(n12572), .B(n12152), .ZN(
        n12574) );
  INV_X1 U15775 ( .A(n12574), .ZN(n12576) );
  XNOR2_X1 U15776 ( .A(n13624), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14411) );
  AOI21_X1 U15777 ( .B1(n12577), .B2(n12576), .A(n12575), .ZN(n14157) );
  INV_X1 U15778 ( .A(n14157), .ZN(n12578) );
  XNOR2_X1 U15779 ( .A(n14221), .B(n12578), .ZN(n14415) );
  NAND2_X1 U15780 ( .A1(n12579), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12580) );
  NAND2_X1 U15781 ( .A1(n12581), .A2(n12580), .ZN(n12590) );
  NAND2_X1 U15782 ( .A1(n9940), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n12582) );
  NAND2_X1 U15783 ( .A1(n12585), .A2(n12582), .ZN(n12609) );
  XNOR2_X1 U15784 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12586) );
  AOI222_X1 U15785 ( .A1(n12622), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .B1(n12622), .B2(n16074), .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .C2(n16074), .ZN(n12906) );
  NOR2_X1 U15786 ( .A1(n12587), .A2(n12586), .ZN(n12588) );
  OR2_X1 U15787 ( .A1(n12589), .A2(n12588), .ZN(n12904) );
  INV_X1 U15788 ( .A(n12631), .ZN(n12594) );
  NAND2_X1 U15789 ( .A1(n12590), .A2(n12595), .ZN(n12591) );
  NAND2_X1 U15790 ( .A1(n12592), .A2(n12591), .ZN(n12903) );
  NOR2_X1 U15791 ( .A1(n11877), .A2(n20804), .ZN(n12600) );
  AOI21_X1 U15792 ( .B1(n12626), .B2(n12903), .A(n12600), .ZN(n12593) );
  OAI21_X1 U15793 ( .B1(n12594), .B2(n13219), .A(n12593), .ZN(n12604) );
  INV_X1 U15794 ( .A(n12604), .ZN(n12608) );
  AND2_X1 U15795 ( .A1(n13246), .A2(n11877), .ZN(n12961) );
  OAI21_X1 U15796 ( .B1(n20635), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n12595), .ZN(n12596) );
  AOI21_X1 U15797 ( .B1(n9657), .B2(n20104), .A(n20114), .ZN(n12616) );
  AOI211_X1 U15798 ( .C1(n12961), .C2(n20104), .A(n12596), .B(n12616), .ZN(
        n12599) );
  INV_X1 U15799 ( .A(n12596), .ZN(n12597) );
  AOI21_X1 U15800 ( .B1(n12631), .B2(n12597), .A(n12632), .ZN(n12598) );
  NOR2_X1 U15801 ( .A1(n12599), .A2(n12598), .ZN(n12605) );
  INV_X1 U15802 ( .A(n12605), .ZN(n12607) );
  INV_X1 U15803 ( .A(n12600), .ZN(n12601) );
  NAND2_X1 U15804 ( .A1(n12601), .A2(n20114), .ZN(n12602) );
  INV_X1 U15805 ( .A(n12903), .ZN(n12603) );
  OAI22_X1 U15806 ( .A1(n12605), .A2(n12604), .B1(n12624), .B2(n12603), .ZN(
        n12606) );
  OAI21_X1 U15807 ( .B1(n12608), .B2(n12607), .A(n12606), .ZN(n12619) );
  NAND2_X1 U15808 ( .A1(n12610), .A2(n12609), .ZN(n12612) );
  NAND2_X1 U15809 ( .A1(n12612), .A2(n12611), .ZN(n12902) );
  INV_X1 U15810 ( .A(n12902), .ZN(n12614) );
  NAND2_X1 U15811 ( .A1(n12631), .A2(n12614), .ZN(n12615) );
  INV_X1 U15812 ( .A(n12616), .ZN(n12613) );
  OAI211_X1 U15813 ( .C1(n12621), .C2(n12614), .A(n12615), .B(n12613), .ZN(
        n12618) );
  INV_X1 U15814 ( .A(n12615), .ZN(n12617) );
  AOI222_X1 U15815 ( .A1(n12619), .A2(n12618), .B1(n12617), .B2(n12616), .C1(
        n12904), .C2(n13690), .ZN(n12620) );
  AOI21_X1 U15816 ( .B1(n12621), .B2(n12904), .A(n12620), .ZN(n12628) );
  AND2_X1 U15817 ( .A1(n16074), .A2(n12622), .ZN(n12623) );
  INV_X1 U15818 ( .A(n12624), .ZN(n12625) );
  NOR2_X1 U15819 ( .A1(n12905), .A2(n12625), .ZN(n12627) );
  OAI22_X1 U15820 ( .A1(n12628), .A2(n12627), .B1(n12626), .B2(n12905), .ZN(
        n12629) );
  OAI21_X1 U15821 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n16074), .A(n12629), 
        .ZN(n12630) );
  AOI21_X1 U15822 ( .B1(n12631), .B2(n12906), .A(n12630), .ZN(n12634) );
  AND2_X1 U15823 ( .A1(n12906), .A2(n12632), .ZN(n12633) );
  NAND3_X1 U15824 ( .A1(n13222), .A2(n20104), .A3(n20124), .ZN(n13256) );
  NOR2_X1 U15825 ( .A1(n13256), .A2(n13219), .ZN(n12635) );
  NAND2_X1 U15826 ( .A1(n15656), .A2(n13242), .ZN(n13121) );
  INV_X1 U15827 ( .A(n12636), .ZN(n12637) );
  INV_X1 U15828 ( .A(n20172), .ZN(n14208) );
  NAND4_X1 U15829 ( .A1(n12637), .A2(n13123), .A3(n13246), .A4(n14208), .ZN(
        n13078) );
  NAND2_X1 U15830 ( .A1(n13121), .A2(n12638), .ZN(n12639) );
  NAND2_X1 U15831 ( .A1(n14168), .A2(P1_EBX_REG_30__SCAN_IN), .ZN(n12642) );
  NAND2_X1 U15832 ( .A1(n14167), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12641) );
  NAND2_X1 U15833 ( .A1(n12642), .A2(n12641), .ZN(n14169) );
  INV_X1 U15834 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12643) );
  INV_X1 U15835 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n12646) );
  NAND2_X1 U15836 ( .A1(n12652), .A2(n12646), .ZN(n12644) );
  NAND3_X1 U15837 ( .A1(n12645), .A2(n12649), .A3(n12644), .ZN(n12648) );
  NAND2_X1 U15838 ( .A1(n9648), .A2(n12646), .ZN(n12647) );
  NAND2_X1 U15839 ( .A1(n12648), .A2(n12647), .ZN(n12653) );
  INV_X1 U15840 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n14293) );
  NAND2_X1 U15841 ( .A1(n12649), .A2(n14293), .ZN(n12650) );
  NAND2_X1 U15842 ( .A1(n12651), .A2(n12650), .ZN(n13096) );
  XNOR2_X1 U15843 ( .A(n12653), .B(n13096), .ZN(n13028) );
  NAND2_X1 U15844 ( .A1(n13028), .A2(n12652), .ZN(n13027) );
  NAND2_X1 U15845 ( .A1(n13027), .A2(n12653), .ZN(n13252) );
  INV_X1 U15846 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13244) );
  INV_X1 U15847 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n19986) );
  NAND2_X1 U15848 ( .A1(n12652), .A2(n19986), .ZN(n12654) );
  NAND3_X1 U15849 ( .A1(n12655), .A2(n12649), .A3(n12654), .ZN(n12657) );
  NAND2_X1 U15850 ( .A1(n9648), .A2(n19986), .ZN(n12656) );
  AND2_X1 U15851 ( .A1(n12657), .A2(n12656), .ZN(n13251) );
  MUX2_X1 U15852 ( .A(n12735), .B(n12649), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n12658) );
  OAI21_X1 U15853 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14168), .A(
        n12658), .ZN(n13383) );
  NAND2_X1 U15854 ( .A1(n12649), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12659) );
  INV_X1 U15855 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n19951) );
  NAND2_X1 U15856 ( .A1(n12652), .A2(n19951), .ZN(n12660) );
  AOI22_X1 U15857 ( .A1(n12661), .A2(n12660), .B1(n9648), .B2(n19951), .ZN(
        n13372) );
  INV_X1 U15858 ( .A(n12735), .ZN(n12709) );
  INV_X1 U15859 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n20009) );
  NAND2_X1 U15860 ( .A1(n12709), .A2(n20009), .ZN(n12665) );
  NAND2_X1 U15861 ( .A1(n12652), .A2(n20009), .ZN(n12663) );
  NAND2_X1 U15862 ( .A1(n12745), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12662) );
  AND2_X1 U15863 ( .A1(n12665), .A2(n12664), .ZN(n16057) );
  NAND2_X1 U15864 ( .A1(n16058), .A2(n16057), .ZN(n16060) );
  INV_X1 U15865 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19999) );
  NAND2_X1 U15866 ( .A1(n12709), .A2(n19999), .ZN(n12669) );
  NAND2_X1 U15867 ( .A1(n12652), .A2(n19999), .ZN(n12667) );
  INV_X1 U15868 ( .A(n9648), .ZN(n12745) );
  NAND2_X1 U15869 ( .A1(n12745), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12666) );
  AND2_X1 U15870 ( .A1(n12669), .A2(n12668), .ZN(n16040) );
  INV_X1 U15871 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16036) );
  INV_X1 U15872 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20003) );
  NAND2_X1 U15873 ( .A1(n12652), .A2(n20003), .ZN(n12670) );
  NAND3_X1 U15874 ( .A1(n12671), .A2(n12745), .A3(n12670), .ZN(n12673) );
  NAND2_X1 U15875 ( .A1(n9648), .A2(n20003), .ZN(n12672) );
  NAND2_X1 U15876 ( .A1(n12673), .A2(n12672), .ZN(n16051) );
  NAND2_X1 U15877 ( .A1(n16040), .A2(n16051), .ZN(n12674) );
  INV_X1 U15878 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16039) );
  INV_X1 U15879 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13635) );
  NAND2_X1 U15880 ( .A1(n12652), .A2(n13635), .ZN(n12675) );
  NAND3_X1 U15881 ( .A1(n12676), .A2(n12745), .A3(n12675), .ZN(n12678) );
  NAND2_X1 U15882 ( .A1(n9648), .A2(n13635), .ZN(n12677) );
  MUX2_X1 U15883 ( .A(n12735), .B(n12745), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n12679) );
  OAI21_X1 U15884 ( .B1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n14168), .A(
        n12679), .ZN(n13740) );
  INV_X1 U15885 ( .A(n13740), .ZN(n12680) );
  INV_X1 U15886 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14508) );
  INV_X1 U15887 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13771) );
  NAND2_X1 U15888 ( .A1(n12652), .A2(n13771), .ZN(n12681) );
  NAND3_X1 U15889 ( .A1(n12682), .A2(n12745), .A3(n12681), .ZN(n12684) );
  NAND2_X1 U15890 ( .A1(n9648), .A2(n13771), .ZN(n12683) );
  MUX2_X1 U15891 ( .A(n12735), .B(n12649), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n12685) );
  OAI21_X1 U15892 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n14168), .A(
        n12685), .ZN(n13890) );
  INV_X1 U15893 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n13931) );
  INV_X1 U15894 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n12688) );
  NAND2_X1 U15895 ( .A1(n12652), .A2(n12688), .ZN(n12686) );
  NAND3_X1 U15896 ( .A1(n12687), .A2(n12745), .A3(n12686), .ZN(n12690) );
  NAND2_X1 U15897 ( .A1(n9648), .A2(n12688), .ZN(n12689) );
  NAND2_X1 U15898 ( .A1(n12690), .A2(n12689), .ZN(n13957) );
  MUX2_X1 U15899 ( .A(n12735), .B(n12745), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n12691) );
  OAI21_X1 U15900 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14168), .A(
        n12691), .ZN(n12692) );
  INV_X1 U15901 ( .A(n12692), .ZN(n13996) );
  INV_X1 U15902 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14059) );
  INV_X1 U15903 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14285) );
  NAND2_X1 U15904 ( .A1(n12652), .A2(n14285), .ZN(n12693) );
  NAND3_X1 U15905 ( .A1(n12694), .A2(n12745), .A3(n12693), .ZN(n12696) );
  NAND2_X1 U15906 ( .A1(n9648), .A2(n14285), .ZN(n12695) );
  AND2_X1 U15907 ( .A1(n12696), .A2(n12695), .ZN(n13939) );
  MUX2_X1 U15908 ( .A(n12735), .B(n12745), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n12697) );
  OAI21_X1 U15909 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n14168), .A(
        n12697), .ZN(n14073) );
  INV_X1 U15910 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15863) );
  INV_X1 U15911 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15787) );
  NAND2_X1 U15912 ( .A1(n12652), .A2(n15787), .ZN(n12698) );
  NAND3_X1 U15913 ( .A1(n12699), .A2(n12745), .A3(n12698), .ZN(n12701) );
  NAND2_X1 U15914 ( .A1(n9648), .A2(n15787), .ZN(n12700) );
  NAND2_X1 U15915 ( .A1(n12701), .A2(n12700), .ZN(n14057) );
  MUX2_X1 U15916 ( .A(n12735), .B(n12745), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n12702) );
  OAI21_X1 U15917 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n14168), .A(
        n12702), .ZN(n12703) );
  INV_X1 U15918 ( .A(n12703), .ZN(n14271) );
  INV_X1 U15919 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15852) );
  INV_X1 U15920 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14344) );
  NAND2_X1 U15921 ( .A1(n12652), .A2(n14344), .ZN(n12704) );
  NAND3_X1 U15922 ( .A1(n12705), .A2(n12745), .A3(n12704), .ZN(n12707) );
  NAND2_X1 U15923 ( .A1(n9648), .A2(n14344), .ZN(n12706) );
  AND2_X1 U15924 ( .A1(n12707), .A2(n12706), .ZN(n13984) );
  MUX2_X1 U15925 ( .A(n12735), .B(n12745), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n12708) );
  OAI21_X1 U15926 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n14168), .A(
        n12708), .ZN(n14341) );
  INV_X1 U15927 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15823) );
  NAND2_X1 U15928 ( .A1(n12709), .A2(n15823), .ZN(n12713) );
  NAND2_X1 U15929 ( .A1(n12652), .A2(n15823), .ZN(n12711) );
  NAND2_X1 U15930 ( .A1(n12745), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12710) );
  AND2_X1 U15931 ( .A1(n12713), .A2(n12712), .ZN(n15676) );
  NAND2_X1 U15932 ( .A1(n12745), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12714) );
  INV_X1 U15933 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14338) );
  NAND2_X1 U15934 ( .A1(n12652), .A2(n14338), .ZN(n12715) );
  NAND2_X1 U15935 ( .A1(n12716), .A2(n12715), .ZN(n12718) );
  OR2_X1 U15936 ( .A1(n12745), .A2(P1_EBX_REG_20__SCAN_IN), .ZN(n12717) );
  NAND2_X1 U15937 ( .A1(n12718), .A2(n12717), .ZN(n15677) );
  NAND2_X1 U15938 ( .A1(n15676), .A2(n15677), .ZN(n12719) );
  INV_X1 U15939 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14461) );
  INV_X1 U15940 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14331) );
  NAND2_X1 U15941 ( .A1(n12652), .A2(n14331), .ZN(n12720) );
  NAND3_X1 U15942 ( .A1(n12721), .A2(n12745), .A3(n12720), .ZN(n12723) );
  NAND2_X1 U15943 ( .A1(n9648), .A2(n14331), .ZN(n12722) );
  NAND2_X1 U15944 ( .A1(n12723), .A2(n12722), .ZN(n14328) );
  MUX2_X1 U15945 ( .A(n12735), .B(n12649), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n12724) );
  OAI21_X1 U15946 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14168), .A(
        n12724), .ZN(n12725) );
  INV_X1 U15947 ( .A(n12725), .ZN(n14321) );
  INV_X1 U15948 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14149) );
  INV_X1 U15949 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15729) );
  NAND2_X1 U15950 ( .A1(n12652), .A2(n15729), .ZN(n12726) );
  NAND3_X1 U15951 ( .A1(n12727), .A2(n12745), .A3(n12726), .ZN(n12729) );
  NAND2_X1 U15952 ( .A1(n9648), .A2(n15729), .ZN(n12728) );
  NAND2_X1 U15953 ( .A1(n12729), .A2(n12728), .ZN(n14314) );
  MUX2_X1 U15954 ( .A(n12735), .B(n12745), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n12730) );
  OAI21_X1 U15955 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14168), .A(
        n12730), .ZN(n14307) );
  INV_X1 U15956 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14448) );
  INV_X1 U15957 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14304) );
  NAND2_X1 U15958 ( .A1(n12652), .A2(n14304), .ZN(n12731) );
  NAND3_X1 U15959 ( .A1(n12732), .A2(n12745), .A3(n12731), .ZN(n12734) );
  OR2_X1 U15960 ( .A1(n12745), .A2(P1_EBX_REG_26__SCAN_IN), .ZN(n12733) );
  AND2_X1 U15961 ( .A1(n12734), .A2(n12733), .ZN(n14247) );
  MUX2_X1 U15962 ( .A(n12735), .B(n12745), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n12736) );
  OAI21_X1 U15963 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14168), .A(
        n12736), .ZN(n12737) );
  INV_X1 U15964 ( .A(n12737), .ZN(n14239) );
  AOI21_X1 U15965 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n12745), .A(
        n12738), .ZN(n12740) );
  NOR2_X1 U15966 ( .A1(n14167), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n12739) );
  OAI22_X1 U15967 ( .A1(n12740), .A2(n12739), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n12745), .ZN(n14099) );
  OR2_X1 U15968 ( .A1(n14168), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12743) );
  INV_X1 U15969 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n12741) );
  NAND2_X1 U15970 ( .A1(n12652), .A2(n12741), .ZN(n12742) );
  NAND2_X1 U15971 ( .A1(n12743), .A2(n12742), .ZN(n12744) );
  MUX2_X1 U15972 ( .A(P1_EBX_REG_29__SCAN_IN), .B(n12744), .S(n12745), .Z(
        n14225) );
  OAI22_X1 U15973 ( .A1(n14224), .A2(n12745), .B1(n12744), .B2(n9695), .ZN(
        n12746) );
  XOR2_X1 U15974 ( .A(n14169), .B(n12746), .Z(n14548) );
  INV_X1 U15975 ( .A(n14548), .ZN(n12747) );
  INV_X1 U15976 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14218) );
  INV_X1 U15977 ( .A(n12748), .ZN(n12749) );
  NOR2_X1 U15978 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n12752) );
  NOR4_X1 U15979 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12751) );
  NAND4_X1 U15980 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n12752), .A4(n12751), .ZN(n12774) );
  NOR4_X1 U15981 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n12756) );
  NOR4_X1 U15982 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_15__SCAN_IN), .A4(
        P1_ADDRESS_REG_17__SCAN_IN), .ZN(n12755) );
  NOR4_X1 U15983 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12754) );
  NOR4_X1 U15984 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n12753) );
  AND4_X1 U15985 ( .A1(n12756), .A2(n12755), .A3(n12754), .A4(n12753), .ZN(
        n12761) );
  NOR4_X1 U15986 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n12759) );
  NOR4_X1 U15987 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n12758) );
  NOR4_X1 U15988 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n12757) );
  INV_X1 U15989 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20826) );
  AND4_X1 U15990 ( .A1(n12759), .A2(n12758), .A3(n12757), .A4(n20826), .ZN(
        n12760) );
  NAND2_X1 U15991 ( .A1(n12761), .A2(n12760), .ZN(n12762) );
  INV_X1 U15992 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20893) );
  NOR3_X1 U15993 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20893), .ZN(n12764) );
  NOR4_X1 U15994 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12763) );
  NAND4_X1 U15995 ( .A1(n20102), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12764), .A4(
        n12763), .ZN(U214) );
  NOR4_X1 U15996 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n12768) );
  NOR4_X1 U15997 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_16__SCAN_IN), .A4(
        P2_ADDRESS_REG_15__SCAN_IN), .ZN(n12767) );
  NOR4_X1 U15998 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n12766) );
  NOR4_X1 U15999 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_9__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_7__SCAN_IN), .ZN(n12765) );
  NAND4_X1 U16000 ( .A1(n12768), .A2(n12767), .A3(n12766), .A4(n12765), .ZN(
        n12773) );
  NOR4_X1 U16001 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_19__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n12771) );
  NOR4_X1 U16002 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n12770) );
  NOR4_X1 U16003 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n12769) );
  INV_X1 U16004 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19757) );
  NAND4_X1 U16005 ( .A1(n12771), .A2(n12770), .A3(n12769), .A4(n19757), .ZN(
        n12772) );
  NOR2_X1 U16006 ( .A1(n13811), .A2(n12774), .ZN(n16424) );
  NAND2_X1 U16007 ( .A1(n16424), .A2(U214), .ZN(U212) );
  INV_X1 U16008 ( .A(n12912), .ZN(n12776) );
  NOR2_X1 U16009 ( .A1(n13465), .A2(n12868), .ZN(n12775) );
  AND2_X1 U16010 ( .A1(n12776), .A2(n12775), .ZN(n19074) );
  INV_X1 U16011 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12777) );
  INV_X1 U16012 ( .A(n13657), .ZN(n12792) );
  OAI211_X1 U16013 ( .C1(n19074), .C2(n12777), .A(n12792), .B(n18862), .ZN(
        P2_U2814) );
  NAND2_X1 U16014 ( .A1(n11032), .A2(n16355), .ZN(n12915) );
  INV_X1 U16015 ( .A(n12915), .ZN(n12779) );
  NOR3_X1 U16016 ( .A1(n12916), .A2(n12779), .A3(n12778), .ZN(n13476) );
  NOR2_X1 U16017 ( .A1(n13476), .A2(n12868), .ZN(n19864) );
  OAI21_X1 U16018 ( .B1(n12921), .B2(n19864), .A(n12780), .ZN(P2_U2819) );
  INV_X1 U16019 ( .A(n18862), .ZN(n12781) );
  OAI21_X1 U16020 ( .B1(n12781), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n18861), 
        .ZN(n12782) );
  OAI21_X1 U16021 ( .B1(n12786), .B2(n18861), .A(n12782), .ZN(P2_U3612) );
  OR2_X1 U16022 ( .A1(n12783), .A2(n19593), .ZN(n13504) );
  NAND2_X1 U16023 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n13424) );
  NOR2_X1 U16024 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13424), .ZN(n19210) );
  INV_X1 U16025 ( .A(n19210), .ZN(n19188) );
  OAI21_X1 U16026 ( .B1(n19743), .B2(n19188), .A(n18861), .ZN(n12784) );
  AOI21_X1 U16027 ( .B1(n19825), .B2(n13504), .A(n12784), .ZN(n12791) );
  INV_X1 U16028 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19736) );
  AOI21_X1 U16029 ( .B1(n19593), .B2(n15457), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n16341) );
  AOI21_X1 U16030 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n16355), .A(n16341), 
        .ZN(n12785) );
  NOR2_X1 U16031 ( .A1(n12791), .A2(n12785), .ZN(n12790) );
  NOR2_X1 U16032 ( .A1(n11027), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n12788) );
  INV_X1 U16033 ( .A(n19737), .ZN(n12787) );
  OAI211_X1 U16034 ( .C1(n12788), .C2(n12787), .A(n12786), .B(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n12789) );
  AOI22_X1 U16035 ( .A1(n12791), .A2(n19736), .B1(n12790), .B2(n12789), .ZN(
        P2_U3610) );
  INV_X1 U16036 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n12795) );
  NAND3_X1 U16037 ( .A1(n13657), .A2(n11027), .A3(n16355), .ZN(n12848) );
  AOI22_X1 U16038 ( .A1(n13809), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13811), .ZN(n19143) );
  NOR2_X1 U16039 ( .A1(n12848), .A2(n19143), .ZN(n12812) );
  AOI21_X1 U16040 ( .B1(n12840), .B2(P2_EAX_REG_5__SCAN_IN), .A(n12812), .ZN(
        n12794) );
  OAI21_X1 U16041 ( .B1(n12793), .B2(n12795), .A(n12794), .ZN(P2_U2972) );
  INV_X1 U16042 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n12797) );
  AOI22_X1 U16043 ( .A1(n13809), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n12843), .ZN(n19240) );
  NOR2_X1 U16044 ( .A1(n12848), .A2(n19240), .ZN(n12809) );
  AOI21_X1 U16045 ( .B1(n12840), .B2(P2_EAX_REG_3__SCAN_IN), .A(n12809), .ZN(
        n12796) );
  OAI21_X1 U16046 ( .B1(n12793), .B2(n12797), .A(n12796), .ZN(P2_U2970) );
  INV_X1 U16047 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n12799) );
  AOI22_X1 U16048 ( .A1(n13809), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13811), .ZN(n19232) );
  NOR2_X1 U16049 ( .A1(n12848), .A2(n19232), .ZN(n12806) );
  AOI21_X1 U16050 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n12840), .A(n12806), .ZN(
        n12798) );
  OAI21_X1 U16051 ( .B1(n12793), .B2(n12799), .A(n12798), .ZN(P2_U2968) );
  INV_X1 U16052 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n12801) );
  AOI22_X1 U16053 ( .A1(n13809), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n12843), .ZN(n19252) );
  NOR2_X1 U16054 ( .A1(n12848), .A2(n19252), .ZN(n12815) );
  AOI21_X1 U16055 ( .B1(n12840), .B2(P2_EAX_REG_6__SCAN_IN), .A(n12815), .ZN(
        n12800) );
  OAI21_X1 U16056 ( .B1(n12793), .B2(n12801), .A(n12800), .ZN(P2_U2973) );
  INV_X1 U16057 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U16058 ( .A1(n13809), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n12843), .ZN(n19259) );
  NOR2_X1 U16059 ( .A1(n12848), .A2(n19259), .ZN(n12821) );
  AOI21_X1 U16060 ( .B1(n12840), .B2(P2_EAX_REG_7__SCAN_IN), .A(n12821), .ZN(
        n12802) );
  OAI21_X1 U16061 ( .B1(n12793), .B2(n12803), .A(n12802), .ZN(P2_U2974) );
  INV_X1 U16062 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n12805) );
  OAI22_X1 U16063 ( .A1(n13811), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13809), .ZN(n16191) );
  NOR2_X1 U16064 ( .A1(n12848), .A2(n16191), .ZN(n12818) );
  AOI21_X1 U16065 ( .B1(n12840), .B2(P2_EAX_REG_2__SCAN_IN), .A(n12818), .ZN(
        n12804) );
  OAI21_X1 U16066 ( .B1(n12793), .B2(n12805), .A(n12804), .ZN(P2_U2969) );
  INV_X1 U16067 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n12808) );
  AOI21_X1 U16068 ( .B1(n12840), .B2(P2_EAX_REG_17__SCAN_IN), .A(n12806), .ZN(
        n12807) );
  OAI21_X1 U16069 ( .B1(n12793), .B2(n12808), .A(n12807), .ZN(P2_U2953) );
  INV_X1 U16070 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n12811) );
  AOI21_X1 U16071 ( .B1(n12840), .B2(P2_EAX_REG_19__SCAN_IN), .A(n12809), .ZN(
        n12810) );
  OAI21_X1 U16072 ( .B1(n12793), .B2(n12811), .A(n12810), .ZN(P2_U2955) );
  INV_X1 U16073 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n12814) );
  AOI21_X1 U16074 ( .B1(n12840), .B2(P2_EAX_REG_21__SCAN_IN), .A(n12812), .ZN(
        n12813) );
  OAI21_X1 U16075 ( .B1(n12793), .B2(n12814), .A(n12813), .ZN(P2_U2957) );
  INV_X1 U16076 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n12817) );
  AOI21_X1 U16077 ( .B1(n12840), .B2(P2_EAX_REG_22__SCAN_IN), .A(n12815), .ZN(
        n12816) );
  OAI21_X1 U16078 ( .B1(n12793), .B2(n12817), .A(n12816), .ZN(P2_U2958) );
  INV_X1 U16079 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n12820) );
  AOI21_X1 U16080 ( .B1(n12840), .B2(P2_EAX_REG_18__SCAN_IN), .A(n12818), .ZN(
        n12819) );
  OAI21_X1 U16081 ( .B1(n12793), .B2(n12820), .A(n12819), .ZN(P2_U2954) );
  INV_X1 U16082 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n12823) );
  AOI21_X1 U16083 ( .B1(n12840), .B2(P2_EAX_REG_23__SCAN_IN), .A(n12821), .ZN(
        n12822) );
  OAI21_X1 U16084 ( .B1(n12793), .B2(n12823), .A(n12822), .ZN(P2_U2959) );
  INV_X1 U16085 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n12828) );
  INV_X1 U16086 ( .A(n12848), .ZN(n12891) );
  INV_X1 U16087 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n12824) );
  OR2_X1 U16088 ( .A1(n13811), .A2(n12824), .ZN(n12826) );
  NAND2_X1 U16089 ( .A1(n13811), .A2(BUF2_REG_9__SCAN_IN), .ZN(n12825) );
  AND2_X1 U16090 ( .A1(n12826), .A2(n12825), .ZN(n19135) );
  INV_X1 U16091 ( .A(n19135), .ZN(n15032) );
  NAND2_X1 U16092 ( .A1(n12891), .A2(n15032), .ZN(n12878) );
  NAND2_X1 U16093 ( .A1(n12840), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n12827) );
  OAI211_X1 U16094 ( .C1(n12793), .C2(n12828), .A(n12878), .B(n12827), .ZN(
        P2_U2976) );
  INV_X1 U16095 ( .A(P2_LWORD_REG_14__SCAN_IN), .ZN(n20924) );
  MUX2_X1 U16096 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n13811), .Z(n19121) );
  NAND2_X1 U16097 ( .A1(n12891), .A2(n19121), .ZN(n12882) );
  NAND2_X1 U16098 ( .A1(n12840), .A2(P2_EAX_REG_14__SCAN_IN), .ZN(n12829) );
  OAI211_X1 U16099 ( .C1(n12793), .C2(n20924), .A(n12882), .B(n12829), .ZN(
        P2_U2981) );
  INV_X1 U16100 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n12835) );
  INV_X1 U16101 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n12830) );
  OR2_X1 U16102 ( .A1(n13811), .A2(n12830), .ZN(n12832) );
  NAND2_X1 U16103 ( .A1(n13811), .A2(BUF2_REG_13__SCAN_IN), .ZN(n12831) );
  AND2_X1 U16104 ( .A1(n12832), .A2(n12831), .ZN(n19124) );
  INV_X1 U16105 ( .A(n19124), .ZN(n12833) );
  NAND2_X1 U16106 ( .A1(n12891), .A2(n12833), .ZN(n12884) );
  NAND2_X1 U16107 ( .A1(n12840), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n12834) );
  OAI211_X1 U16108 ( .C1(n12793), .C2(n12835), .A(n12884), .B(n12834), .ZN(
        P2_U2980) );
  INV_X1 U16109 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n12842) );
  INV_X1 U16110 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n12836) );
  OR2_X1 U16111 ( .A1(n13811), .A2(n12836), .ZN(n12838) );
  NAND2_X1 U16112 ( .A1(n13811), .A2(BUF2_REG_11__SCAN_IN), .ZN(n12837) );
  AND2_X1 U16113 ( .A1(n12838), .A2(n12837), .ZN(n19129) );
  INV_X1 U16114 ( .A(n19129), .ZN(n12839) );
  NAND2_X1 U16115 ( .A1(n12891), .A2(n12839), .ZN(n12876) );
  NAND2_X1 U16116 ( .A1(n12840), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n12841) );
  OAI211_X1 U16117 ( .C1(n12793), .C2(n12842), .A(n12876), .B(n12841), .ZN(
        P2_U2978) );
  INV_X1 U16118 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12844) );
  AOI22_X1 U16119 ( .A1(n13809), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n12843), .ZN(n19118) );
  INV_X1 U16120 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19185) );
  OAI222_X1 U16121 ( .A1(n12793), .A2(n12844), .B1(n12848), .B2(n19118), .C1(
        n12901), .C2(n19185), .ZN(P2_U2982) );
  INV_X1 U16122 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n12846) );
  OAI22_X1 U16123 ( .A1(n13811), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13809), .ZN(n19107) );
  INV_X1 U16124 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12845) );
  OAI222_X1 U16125 ( .A1(n12846), .A2(n12793), .B1(n12848), .B2(n19107), .C1(
        n12845), .C2(n12901), .ZN(P2_U2967) );
  INV_X1 U16126 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n21052) );
  INV_X1 U16127 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n12847) );
  OAI222_X1 U16128 ( .A1(n12848), .A2(n19107), .B1(n12793), .B2(n21052), .C1(
        n12847), .C2(n12901), .ZN(P2_U2952) );
  OAI21_X1 U16129 ( .B1(n19056), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12859), .ZN(n16325) );
  INV_X1 U16130 ( .A(n16325), .ZN(n12854) );
  NAND2_X1 U16131 ( .A1(n12849), .A2(n16335), .ZN(n12850) );
  NAND2_X1 U16132 ( .A1(n12851), .A2(n12850), .ZN(n16338) );
  OR2_X1 U16133 ( .A1(n19046), .A2(n12852), .ZN(n16336) );
  OAI21_X1 U16134 ( .B1(n19219), .B2(n16338), .A(n16336), .ZN(n12853) );
  AOI21_X1 U16135 ( .B1(n11389), .B2(n12854), .A(n12853), .ZN(n12857) );
  OAI21_X1 U16136 ( .B1(n19218), .B2(n12855), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12856) );
  OAI211_X1 U16137 ( .C1(n16273), .C2(n16328), .A(n12857), .B(n12856), .ZN(
        P2_U3014) );
  OAI21_X1 U16138 ( .B1(n14669), .B2(n12859), .A(n12858), .ZN(n12860) );
  XOR2_X1 U16139 ( .A(n12860), .B(n15456), .Z(n12993) );
  AOI21_X1 U16140 ( .B1(n15456), .B2(n12862), .A(n12861), .ZN(n12994) );
  NOR2_X1 U16141 ( .A1(n19046), .A2(n19753), .ZN(n12992) );
  AOI21_X1 U16142 ( .B1(n16269), .B2(n12994), .A(n12992), .ZN(n12865) );
  NAND2_X1 U16143 ( .A1(n16268), .A2(n12863), .ZN(n12864) );
  OAI211_X1 U16144 ( .C1(n16278), .C2(n12863), .A(n12865), .B(n12864), .ZN(
        n12866) );
  AOI21_X1 U16145 ( .B1(n11389), .B2(n12993), .A(n12866), .ZN(n12867) );
  OAI21_X1 U16146 ( .B1(n14673), .B2(n16273), .A(n12867), .ZN(P2_U3013) );
  NOR2_X1 U16147 ( .A1(n12912), .A2(n12868), .ZN(n12869) );
  NAND2_X1 U16148 ( .A1(n12914), .A2(n12869), .ZN(n12870) );
  NAND2_X1 U16149 ( .A1(n12870), .A2(n12901), .ZN(n12871) );
  INV_X1 U16150 ( .A(n19188), .ZN(n19214) );
  INV_X1 U16151 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n12874) );
  NAND2_X1 U16152 ( .A1(n19186), .A2(n12872), .ZN(n12946) );
  INV_X1 U16153 ( .A(n12946), .ZN(n19181) );
  AOI22_X1 U16154 ( .A1(n19181), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n19214), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n12873) );
  OAI21_X1 U16155 ( .B1(n19183), .B2(n12874), .A(n12873), .ZN(P2_U2935) );
  INV_X1 U16156 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19191) );
  NAND2_X1 U16157 ( .A1(n12898), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12875) );
  MUX2_X1 U16158 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n13811), .Z(n19126) );
  NAND2_X1 U16159 ( .A1(n12891), .A2(n19126), .ZN(n12880) );
  OAI211_X1 U16160 ( .C1(n19191), .C2(n12901), .A(n12875), .B(n12880), .ZN(
        P2_U2979) );
  INV_X1 U16161 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15017) );
  NAND2_X1 U16162 ( .A1(n12898), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n12877) );
  OAI211_X1 U16163 ( .C1(n12901), .C2(n15017), .A(n12877), .B(n12876), .ZN(
        P2_U2963) );
  INV_X1 U16164 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n12935) );
  NAND2_X1 U16165 ( .A1(n12898), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n12879) );
  OAI211_X1 U16166 ( .C1(n12901), .C2(n12935), .A(n12879), .B(n12878), .ZN(
        P2_U2961) );
  INV_X1 U16167 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n12939) );
  NAND2_X1 U16168 ( .A1(n12898), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12881) );
  OAI211_X1 U16169 ( .C1(n12939), .C2(n12901), .A(n12881), .B(n12880), .ZN(
        P2_U2964) );
  INV_X1 U16170 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12942) );
  NAND2_X1 U16171 ( .A1(n12898), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n12883) );
  OAI211_X1 U16172 ( .C1(n12942), .C2(n12901), .A(n12883), .B(n12882), .ZN(
        P2_U2966) );
  INV_X1 U16173 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n15000) );
  NAND2_X1 U16174 ( .A1(n12898), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n12885) );
  OAI211_X1 U16175 ( .C1(n12901), .C2(n15000), .A(n12885), .B(n12884), .ZN(
        P2_U2965) );
  INV_X1 U16176 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19195) );
  NAND2_X1 U16177 ( .A1(n12898), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12886) );
  MUX2_X1 U16178 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n13811), .Z(n19132) );
  NAND2_X1 U16179 ( .A1(n12891), .A2(n19132), .ZN(n12893) );
  OAI211_X1 U16180 ( .C1(n19195), .C2(n12901), .A(n12886), .B(n12893), .ZN(
        P2_U2977) );
  INV_X1 U16181 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n12888) );
  NAND2_X1 U16182 ( .A1(n12898), .A2(P2_UWORD_REG_4__SCAN_IN), .ZN(n12887) );
  OAI22_X1 U16183 ( .A1(n13811), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13809), .ZN(n19245) );
  INV_X1 U16184 ( .A(n19245), .ZN(n16184) );
  NAND2_X1 U16185 ( .A1(n12891), .A2(n16184), .ZN(n12895) );
  OAI211_X1 U16186 ( .C1(n12901), .C2(n12888), .A(n12887), .B(n12895), .ZN(
        P2_U2956) );
  INV_X1 U16187 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19199) );
  NAND2_X1 U16188 ( .A1(n12898), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12892) );
  NAND2_X1 U16189 ( .A1(n13811), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12890) );
  INV_X1 U16190 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16463) );
  OR2_X1 U16191 ( .A1(n13811), .A2(n16463), .ZN(n12889) );
  NAND2_X1 U16192 ( .A1(n12890), .A2(n12889), .ZN(n19138) );
  NAND2_X1 U16193 ( .A1(n12891), .A2(n19138), .ZN(n12899) );
  OAI211_X1 U16194 ( .C1(n19199), .C2(n12901), .A(n12892), .B(n12899), .ZN(
        P2_U2975) );
  INV_X1 U16195 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n21081) );
  NAND2_X1 U16196 ( .A1(n12898), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12894) );
  OAI211_X1 U16197 ( .C1(n21081), .C2(n12901), .A(n12894), .B(n12893), .ZN(
        P2_U2962) );
  INV_X1 U16198 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n12897) );
  NAND2_X1 U16199 ( .A1(n12898), .A2(P2_LWORD_REG_4__SCAN_IN), .ZN(n12896) );
  OAI211_X1 U16200 ( .C1(n12901), .C2(n12897), .A(n12896), .B(n12895), .ZN(
        P2_U2971) );
  INV_X1 U16201 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n12933) );
  NAND2_X1 U16202 ( .A1(n12898), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12900) );
  OAI211_X1 U16203 ( .C1(n12933), .C2(n12901), .A(n12900), .B(n12899), .ZN(
        P2_U2960) );
  NOR3_X1 U16204 ( .A1(n12904), .A2(n12903), .A3(n12902), .ZN(n12907) );
  OAI21_X1 U16205 ( .B1(n12907), .B2(n12906), .A(n12905), .ZN(n13076) );
  NAND2_X1 U16206 ( .A1(n12951), .A2(n13213), .ZN(n12947) );
  INV_X1 U16207 ( .A(n12947), .ZN(n12910) );
  INV_X1 U16208 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n12909) );
  NAND2_X1 U16209 ( .A1(n20741), .A2(n21068), .ZN(n19874) );
  OAI211_X1 U16210 ( .C1(n12910), .C2(n12909), .A(n12948), .B(n19874), .ZN(
        P1_U2801) );
  NOR2_X1 U16211 ( .A1(n12912), .A2(n12911), .ZN(n12913) );
  NAND2_X1 U16212 ( .A1(n12914), .A2(n12913), .ZN(n12920) );
  INV_X1 U16213 ( .A(n13295), .ZN(n13468) );
  NOR2_X1 U16214 ( .A1(n12916), .A2(n12915), .ZN(n12917) );
  AOI21_X1 U16215 ( .B1(n13467), .B2(n13468), .A(n12917), .ZN(n12969) );
  INV_X1 U16216 ( .A(n12918), .ZN(n12919) );
  INV_X1 U16217 ( .A(n13467), .ZN(n13469) );
  INV_X1 U16218 ( .A(n13296), .ZN(n13466) );
  NAND2_X1 U16219 ( .A1(n13469), .A2(n13466), .ZN(n13004) );
  AND4_X1 U16220 ( .A1(n12920), .A2(n12969), .A3(n12919), .A4(n13004), .ZN(
        n13498) );
  NOR2_X1 U16221 ( .A1(n16342), .A2(n13424), .ZN(n15709) );
  INV_X1 U16222 ( .A(n15709), .ZN(n13509) );
  OAI22_X1 U16223 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19825), .B1(n13509), 
        .B2(n12921), .ZN(n12922) );
  INV_X1 U16224 ( .A(n15470), .ZN(n12926) );
  NOR2_X1 U16225 ( .A1(n12924), .A2(n12923), .ZN(n13475) );
  NAND4_X1 U16226 ( .A1(n12926), .A2(n13474), .A3(n13475), .A4(n15463), .ZN(
        n12925) );
  OAI21_X1 U16227 ( .B1(n12927), .B2(n12926), .A(n12925), .ZN(P2_U3595) );
  INV_X1 U16228 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n15083) );
  INV_X2 U16229 ( .A(n19183), .ZN(n19213) );
  AOI22_X1 U16230 ( .A1(n19210), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12928) );
  OAI21_X1 U16231 ( .B1(n15083), .B2(n12946), .A(n12928), .ZN(P2_U2932) );
  INV_X1 U16232 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n15076) );
  AOI22_X1 U16233 ( .A1(n19210), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12929) );
  OAI21_X1 U16234 ( .B1(n15076), .B2(n12946), .A(n12929), .ZN(P2_U2930) );
  INV_X1 U16235 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n15069) );
  AOI22_X1 U16236 ( .A1(n19210), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12930) );
  OAI21_X1 U16237 ( .B1(n15069), .B2(n12946), .A(n12930), .ZN(P2_U2929) );
  INV_X1 U16238 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15058) );
  AOI22_X1 U16239 ( .A1(n19210), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12931) );
  OAI21_X1 U16240 ( .B1(n15058), .B2(n12946), .A(n12931), .ZN(P2_U2928) );
  AOI22_X1 U16241 ( .A1(n19210), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12932) );
  OAI21_X1 U16242 ( .B1(n12933), .B2(n12946), .A(n12932), .ZN(P2_U2927) );
  AOI22_X1 U16243 ( .A1(n19210), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12934) );
  OAI21_X1 U16244 ( .B1(n12935), .B2(n12946), .A(n12934), .ZN(P2_U2926) );
  AOI22_X1 U16245 ( .A1(n19210), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12936) );
  OAI21_X1 U16246 ( .B1(n21081), .B2(n12946), .A(n12936), .ZN(P2_U2925) );
  AOI22_X1 U16247 ( .A1(n19214), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12937) );
  OAI21_X1 U16248 ( .B1(n15017), .B2(n12946), .A(n12937), .ZN(P2_U2924) );
  AOI22_X1 U16249 ( .A1(n19214), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12938) );
  OAI21_X1 U16250 ( .B1(n12939), .B2(n12946), .A(n12938), .ZN(P2_U2923) );
  AOI22_X1 U16251 ( .A1(n19214), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12940) );
  OAI21_X1 U16252 ( .B1(n15000), .B2(n12946), .A(n12940), .ZN(P2_U2922) );
  AOI22_X1 U16253 ( .A1(n19214), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n12941) );
  OAI21_X1 U16254 ( .B1(n12942), .B2(n12946), .A(n12941), .ZN(P2_U2921) );
  INV_X1 U16255 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n12944) );
  AOI22_X1 U16256 ( .A1(n19210), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12943) );
  OAI21_X1 U16257 ( .B1(n12944), .B2(n12946), .A(n12943), .ZN(P2_U2933) );
  INV_X1 U16258 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n13810) );
  AOI22_X1 U16259 ( .A1(n19210), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12945) );
  OAI21_X1 U16260 ( .B1(n13810), .B2(n12946), .A(n12945), .ZN(P2_U2934) );
  INV_X1 U16261 ( .A(n19874), .ZN(n13629) );
  NOR2_X1 U16262 ( .A1(n13629), .A2(P1_READREQUEST_REG_SCAN_IN), .ZN(n12950)
         );
  OAI21_X1 U16263 ( .B1(n13719), .B2(n9648), .A(n20894), .ZN(n12949) );
  OAI21_X1 U16264 ( .B1(n12950), .B2(n20894), .A(n12949), .ZN(P1_U3487) );
  INV_X1 U16265 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n12967) );
  OAI22_X1 U16266 ( .A1(n13209), .A2(n13719), .B1(n12952), .B2(n12951), .ZN(
        n19872) );
  INV_X1 U16267 ( .A(n13719), .ZN(n13130) );
  INV_X1 U16268 ( .A(n12953), .ZN(n12954) );
  NAND2_X1 U16269 ( .A1(n12954), .A2(n20808), .ZN(n15697) );
  NAND3_X1 U16270 ( .A1(n13130), .A2(n14167), .A3(n15697), .ZN(n12955) );
  NAND2_X1 U16271 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n20896) );
  AND2_X1 U16272 ( .A1(n12955), .A2(n20896), .ZN(n20897) );
  NOR2_X1 U16273 ( .A1(n19872), .A2(n20897), .ZN(n15644) );
  NOR2_X1 U16274 ( .A1(n15644), .A2(n19871), .ZN(n19879) );
  INV_X1 U16275 ( .A(n12956), .ZN(n12957) );
  NOR3_X1 U16276 ( .A1(n12957), .A2(n13256), .A3(n20136), .ZN(n12962) );
  INV_X1 U16277 ( .A(n12958), .ZN(n12960) );
  NAND2_X1 U16278 ( .A1(n14594), .A2(n13619), .ZN(n12959) );
  AND2_X1 U16279 ( .A1(n13114), .A2(n13719), .ZN(n13109) );
  OR2_X1 U16280 ( .A1(n13109), .A2(n15642), .ZN(n13217) );
  OAI21_X1 U16281 ( .B1(n12962), .B2(n13217), .A(n15656), .ZN(n12963) );
  OAI21_X1 U16282 ( .B1(n13076), .B2(n13116), .A(n12963), .ZN(n12964) );
  AOI21_X1 U16283 ( .B1(n13242), .B2(n13209), .A(n12964), .ZN(n12965) );
  NOR2_X1 U16284 ( .A1(n12965), .A2(n14208), .ZN(n15643) );
  NAND2_X1 U16285 ( .A1(n15643), .A2(n19879), .ZN(n12966) );
  OAI21_X1 U16286 ( .B1(n12967), .B2(n19879), .A(n12966), .ZN(P1_U3484) );
  NAND2_X1 U16287 ( .A1(n12969), .A2(n12968), .ZN(n12970) );
  AND2_X1 U16288 ( .A1(n9649), .A2(n19257), .ZN(n12972) );
  AND2_X1 U16289 ( .A1(n19169), .A2(n12973), .ZN(n13812) );
  INV_X1 U16290 ( .A(n13049), .ZN(n13012) );
  NAND2_X1 U16291 ( .A1(n19251), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12974) );
  AND2_X1 U16292 ( .A1(n19825), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12977) );
  OAI211_X1 U16293 ( .C1(n19231), .C2(n13846), .A(n12978), .B(n12977), .ZN(
        n12979) );
  INV_X1 U16294 ( .A(n12979), .ZN(n12980) );
  NOR2_X1 U16295 ( .A1(n12982), .A2(n12981), .ZN(n12983) );
  OR2_X1 U16296 ( .A1(n12984), .A2(n12983), .ZN(n16329) );
  INV_X1 U16297 ( .A(n16329), .ZN(n19060) );
  NAND2_X1 U16298 ( .A1(n19073), .A2(n19060), .ZN(n19173) );
  OAI211_X1 U16299 ( .C1(n19073), .C2(n19060), .A(n19173), .B(n19175), .ZN(
        n12988) );
  AOI22_X1 U16300 ( .A1(n19171), .A2(n19060), .B1(n19170), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n12987) );
  OAI211_X1 U16301 ( .C1(n19179), .C2(n19107), .A(n12988), .B(n12987), .ZN(
        P2_U2919) );
  XNOR2_X1 U16302 ( .A(n12990), .B(n12989), .ZN(n19844) );
  AOI22_X1 U16303 ( .A1(n16312), .A2(n19844), .B1(n12991), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12998) );
  AOI21_X1 U16304 ( .B1(n16317), .B2(n12993), .A(n12992), .ZN(n12997) );
  NAND2_X1 U16305 ( .A1(n16314), .A2(n12994), .ZN(n12996) );
  OAI211_X1 U16306 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(n16334), .B(n14193), .ZN(n12995) );
  AND4_X1 U16307 ( .A1(n12998), .A2(n12997), .A3(n12996), .A4(n12995), .ZN(
        n12999) );
  OAI21_X1 U16308 ( .B1(n14673), .B2(n16327), .A(n12999), .ZN(P2_U3045) );
  NAND2_X1 U16309 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19846), .ZN(
        n19496) );
  NAND2_X1 U16310 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19855), .ZN(
        n19526) );
  NAND2_X1 U16311 ( .A1(n19496), .A2(n19526), .ZN(n13536) );
  AND2_X1 U16312 ( .A1(n19830), .A2(n13536), .ZN(n19525) );
  AOI21_X1 U16313 ( .B1(n13054), .B2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n19525), .ZN(n13001) );
  NAND2_X1 U16314 ( .A1(n13003), .A2(n13002), .ZN(n13289) );
  NAND2_X1 U16315 ( .A1(n13004), .A2(n13289), .ZN(n13005) );
  INV_X2 U16316 ( .A(n19103), .ZN(n19089) );
  MUX2_X1 U16317 ( .A(n14673), .B(n13006), .S(n19089), .Z(n13007) );
  OAI21_X1 U16318 ( .B1(n19832), .B2(n19095), .A(n13007), .ZN(P2_U2886) );
  NAND2_X1 U16319 ( .A1(n19073), .A2(n19100), .ZN(n13009) );
  NAND2_X1 U16320 ( .A1(n19103), .A2(n9647), .ZN(n13008) );
  OAI211_X1 U16321 ( .C1(n19058), .C2(n19103), .A(n13009), .B(n13008), .ZN(
        P2_U2887) );
  INV_X1 U16322 ( .A(n19830), .ZN(n19676) );
  NAND2_X1 U16323 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19328) );
  NAND2_X1 U16324 ( .A1(n19328), .A2(n19837), .ZN(n13013) );
  NOR2_X1 U16325 ( .A1(n19837), .A2(n19846), .ZN(n19667) );
  NAND2_X1 U16326 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19667), .ZN(
        n13051) );
  NAND2_X1 U16327 ( .A1(n13013), .A2(n13051), .ZN(n13537) );
  NOR2_X1 U16328 ( .A1(n19676), .A2(n13537), .ZN(n13014) );
  AOI21_X1 U16329 ( .B1(n13054), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n13014), .ZN(n13015) );
  XNOR2_X1 U16330 ( .A(n13061), .B(n13017), .ZN(n13018) );
  MUX2_X1 U16331 ( .A(n10380), .B(n10331), .S(n19089), .Z(n13019) );
  OAI21_X1 U16332 ( .B1(n19831), .B2(n19095), .A(n13019), .ZN(P2_U2885) );
  NAND2_X1 U16333 ( .A1(n13020), .A2(n13021), .ZN(n13023) );
  NAND2_X1 U16334 ( .A1(n13023), .A2(n13022), .ZN(n13026) );
  INV_X1 U16335 ( .A(n13024), .ZN(n13084) );
  OAI21_X1 U16336 ( .B1(n13026), .B2(n13025), .A(n13084), .ZN(n13731) );
  OAI21_X1 U16337 ( .B1(n13028), .B2(n12652), .A(n13027), .ZN(n13721) );
  AOI22_X1 U16338 ( .A1(n20012), .A2(n13721), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14310), .ZN(n13029) );
  OAI21_X1 U16339 ( .B1(n14350), .B2(n13731), .A(n13029), .ZN(P1_U2871) );
  INV_X1 U16340 ( .A(n20896), .ZN(n20814) );
  NAND2_X1 U16341 ( .A1(n20898), .A2(n20814), .ZN(n13030) );
  AND2_X2 U16342 ( .A1(n13182), .A2(n13219), .ZN(n20069) );
  INV_X1 U16343 ( .A(n20069), .ZN(n13181) );
  AND2_X1 U16344 ( .A1(n20114), .A2(n20896), .ZN(n13031) );
  INV_X1 U16345 ( .A(n20102), .ZN(n20100) );
  INV_X1 U16346 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13033) );
  NOR2_X1 U16347 ( .A1(n20100), .A2(n13033), .ZN(n13034) );
  AOI21_X1 U16348 ( .B1(DATAI_15_), .B2(n20100), .A(n13034), .ZN(n14075) );
  INV_X1 U16349 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13035) );
  OAI222_X1 U16350 ( .A1(n13181), .A2(n12265), .B1(n13180), .B2(n14075), .C1(
        n13182), .C2(n13035), .ZN(P1_U2967) );
  INV_X1 U16351 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13040) );
  OR2_X1 U16352 ( .A1(n13201), .A2(n20898), .ZN(n13249) );
  NOR2_X1 U16353 ( .A1(n13249), .A2(n15697), .ZN(n15654) );
  INV_X1 U16354 ( .A(n15654), .ZN(n13037) );
  INV_X1 U16355 ( .A(n15697), .ZN(n13199) );
  NAND2_X1 U16356 ( .A1(n15628), .A2(n13199), .ZN(n13106) );
  NAND2_X1 U16357 ( .A1(n13037), .A2(n13106), .ZN(n13038) );
  NAND2_X1 U16358 ( .A1(n20026), .A2(n20104), .ZN(n13100) );
  NAND2_X1 U16359 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16079) );
  INV_X1 U16360 ( .A(n16079), .ZN(n13172) );
  NAND2_X1 U16361 ( .A1(n20804), .A2(n13172), .ZN(n20019) );
  INV_X2 U16362 ( .A(n20019), .ZN(n20039) );
  AOI22_X1 U16363 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20038), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20039), .ZN(n13039) );
  OAI21_X1 U16364 ( .B1(n13040), .B2(n13100), .A(n13039), .ZN(P1_U2920) );
  AOI22_X1 U16365 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13041) );
  OAI21_X1 U16366 ( .B1(n12335), .B2(n13100), .A(n13041), .ZN(P1_U2917) );
  AOI22_X1 U16367 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13042) );
  OAI21_X1 U16368 ( .B1(n12422), .B2(n13100), .A(n13042), .ZN(P1_U2913) );
  AOI22_X1 U16369 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13043) );
  OAI21_X1 U16370 ( .B1(n14384), .B2(n13100), .A(n13043), .ZN(P1_U2916) );
  AOI22_X1 U16371 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13044) );
  OAI21_X1 U16372 ( .B1(n14379), .B2(n13100), .A(n13044), .ZN(P1_U2915) );
  AOI22_X1 U16373 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13045) );
  OAI21_X1 U16374 ( .B1(n12301), .B2(n13100), .A(n13045), .ZN(P1_U2919) );
  AOI22_X1 U16375 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13046) );
  OAI21_X1 U16376 ( .B1(n12573), .B2(n13100), .A(n13046), .ZN(P1_U2906) );
  AOI22_X1 U16377 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13047) );
  OAI21_X1 U16378 ( .B1(n12393), .B2(n13100), .A(n13047), .ZN(P1_U2914) );
  AOI22_X1 U16379 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13048) );
  OAI21_X1 U16380 ( .B1(n14392), .B2(n13100), .A(n13048), .ZN(P1_U2918) );
  INV_X1 U16381 ( .A(n13051), .ZN(n13050) );
  NAND2_X1 U16382 ( .A1(n13050), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19675) );
  NAND2_X1 U16383 ( .A1(n19829), .A2(n13051), .ZN(n13052) );
  AND3_X1 U16384 ( .A1(n19675), .A2(n19830), .A3(n13052), .ZN(n13053) );
  AOI21_X1 U16385 ( .B1(n13054), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n13053), .ZN(n13055) );
  NAND2_X1 U16386 ( .A1(n13192), .A2(n13056), .ZN(n13057) );
  INV_X1 U16387 ( .A(n13060), .ZN(n13058) );
  NAND2_X1 U16388 ( .A1(n13058), .A2(n13017), .ZN(n13064) );
  NAND2_X1 U16389 ( .A1(n13060), .A2(n13059), .ZN(n13062) );
  NAND2_X1 U16390 ( .A1(n13062), .A2(n13061), .ZN(n13063) );
  NAND2_X1 U16391 ( .A1(n13064), .A2(n13063), .ZN(n13066) );
  INV_X1 U16392 ( .A(n13068), .ZN(n16272) );
  MUX2_X1 U16393 ( .A(n16272), .B(n13069), .S(n19089), .Z(n13070) );
  OAI21_X1 U16394 ( .B1(n19269), .B2(n19095), .A(n13070), .ZN(P2_U2884) );
  NAND2_X1 U16395 ( .A1(n13072), .A2(n13071), .ZN(n13073) );
  NAND2_X1 U16396 ( .A1(n13074), .A2(n13073), .ZN(n20079) );
  NAND2_X1 U16397 ( .A1(n13209), .A2(n13109), .ZN(n13077) );
  INV_X1 U16398 ( .A(n13075), .ZN(n16070) );
  AND2_X1 U16399 ( .A1(n20896), .A2(n13076), .ZN(n13203) );
  NAND2_X1 U16400 ( .A1(n16070), .A2(n13203), .ZN(n13117) );
  OAI211_X1 U16401 ( .C1(n13130), .C2(n13078), .A(n13077), .B(n13117), .ZN(
        n13079) );
  NAND2_X1 U16402 ( .A1(n13079), .A2(n13213), .ZN(n13080) );
  NAND2_X1 U16403 ( .A1(n11884), .A2(n20172), .ZN(n13081) );
  MUX2_X1 U16404 ( .A(DATAI_0_), .B(BUF1_REG_0__SCAN_IN), .S(n20102), .Z(
        n20099) );
  INV_X1 U16405 ( .A(n20099), .ZN(n13082) );
  INV_X1 U16406 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20042) );
  OAI222_X1 U16407 ( .A1(n20079), .A2(n14370), .B1(n14076), .B2(n13082), .C1(
        n14402), .C2(n20042), .ZN(P1_U2904) );
  MUX2_X1 U16408 ( .A(DATAI_1_), .B(BUF1_REG_1__SCAN_IN), .S(n20102), .Z(
        n20113) );
  INV_X1 U16409 ( .A(n20113), .ZN(n13083) );
  OAI222_X1 U16410 ( .A1(n13731), .A2(n14370), .B1(n14076), .B2(n13083), .C1(
        n14402), .C2(n12064), .ZN(P1_U2903) );
  NAND2_X1 U16411 ( .A1(n13085), .A2(n13084), .ZN(n13086) );
  AND2_X1 U16412 ( .A1(n13087), .A2(n13086), .ZN(n19990) );
  INV_X1 U16413 ( .A(n19990), .ZN(n14125) );
  MUX2_X1 U16414 ( .A(DATAI_2_), .B(BUF1_REG_2__SCAN_IN), .S(n20102), .Z(
        n20118) );
  INV_X1 U16415 ( .A(n20118), .ZN(n13088) );
  OAI222_X1 U16416 ( .A1(n14125), .A2(n14370), .B1(n14076), .B2(n13088), .C1(
        n14402), .C2(n12071), .ZN(P1_U2902) );
  INV_X1 U16417 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13090) );
  AOI22_X1 U16418 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13089) );
  OAI21_X1 U16419 ( .B1(n13090), .B2(n13100), .A(n13089), .ZN(P1_U2909) );
  INV_X1 U16420 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n13092) );
  AOI22_X1 U16421 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13091) );
  OAI21_X1 U16422 ( .B1(n13092), .B2(n13100), .A(n13091), .ZN(P1_U2908) );
  AOI22_X1 U16423 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13093) );
  OAI21_X1 U16424 ( .B1(n12460), .B2(n13100), .A(n13093), .ZN(P1_U2911) );
  INV_X1 U16425 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n13095) );
  AOI22_X1 U16426 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13094) );
  OAI21_X1 U16427 ( .B1(n13095), .B2(n13100), .A(n13094), .ZN(P1_U2912) );
  OAI21_X1 U16428 ( .B1(n14168), .B2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13096), .ZN(n20083) );
  OAI222_X1 U16429 ( .A1(n20083), .A2(n20005), .B1(n14293), .B2(n20016), .C1(
        n20079), .C2(n14350), .ZN(P1_U2872) );
  INV_X1 U16430 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13098) );
  AOI22_X1 U16431 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13097) );
  OAI21_X1 U16432 ( .B1(n13098), .B2(n13100), .A(n13097), .ZN(P1_U2907) );
  AOI22_X1 U16433 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13099) );
  OAI21_X1 U16434 ( .B1(n12483), .B2(n13100), .A(n13099), .ZN(P1_U2910) );
  OAI21_X1 U16435 ( .B1(n13103), .B2(n13102), .A(n13101), .ZN(n19971) );
  MUX2_X1 U16436 ( .A(DATAI_3_), .B(BUF1_REG_3__SCAN_IN), .S(n20102), .Z(
        n20123) );
  INV_X1 U16437 ( .A(n20123), .ZN(n13105) );
  OAI222_X1 U16438 ( .A1(n19971), .A2(n14370), .B1(n14076), .B2(n13105), .C1(
        n13104), .C2(n14402), .ZN(P1_U2901) );
  INV_X1 U16439 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19878) );
  AND2_X1 U16440 ( .A1(n19878), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13166) );
  NOR2_X1 U16441 ( .A1(n12652), .A2(n13199), .ZN(n13107) );
  OAI21_X1 U16442 ( .B1(n13107), .B2(n13201), .A(n13106), .ZN(n13108) );
  NAND2_X1 U16443 ( .A1(n13108), .A2(n20896), .ZN(n13110) );
  INV_X1 U16444 ( .A(n13109), .ZN(n13138) );
  NAND2_X1 U16445 ( .A1(n13110), .A2(n13138), .ZN(n13119) );
  NAND2_X1 U16446 ( .A1(n13619), .A2(n20114), .ZN(n13124) );
  AOI21_X1 U16447 ( .B1(n13690), .B2(n13111), .A(n13619), .ZN(n13112) );
  NAND2_X1 U16448 ( .A1(n13113), .A2(n13112), .ZN(n13127) );
  NAND2_X1 U16449 ( .A1(n13114), .A2(n13127), .ZN(n13115) );
  NAND2_X1 U16450 ( .A1(n13116), .A2(n13115), .ZN(n13207) );
  OAI211_X1 U16451 ( .C1(n20119), .C2(n13124), .A(n13117), .B(n13207), .ZN(
        n13118) );
  AOI21_X1 U16452 ( .B1(n13209), .B2(n13119), .A(n13118), .ZN(n13120) );
  INV_X1 U16453 ( .A(n13122), .ZN(n20094) );
  OR2_X1 U16454 ( .A1(n13123), .A2(n11842), .ZN(n13125) );
  INV_X1 U16455 ( .A(n13124), .ZN(n13722) );
  AOI22_X1 U16456 ( .A1(n13125), .A2(n13722), .B1(n20119), .B2(n14096), .ZN(
        n13126) );
  AND2_X1 U16457 ( .A1(n13127), .A2(n13126), .ZN(n13129) );
  OAI211_X1 U16458 ( .C1(n13131), .C2(n13130), .A(n13129), .B(n13128), .ZN(
        n13255) );
  NAND3_X1 U16459 ( .A1(n13201), .A2(n13133), .A3(n13132), .ZN(n13134) );
  NOR2_X1 U16460 ( .A1(n13255), .A2(n13134), .ZN(n13135) );
  NAND2_X1 U16461 ( .A1(n13135), .A2(n13075), .ZN(n14597) );
  NAND2_X1 U16462 ( .A1(n14599), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13147) );
  INV_X1 U16463 ( .A(n13147), .ZN(n13136) );
  NOR2_X1 U16464 ( .A1(n14599), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13146) );
  OR2_X1 U16465 ( .A1(n13136), .A2(n13146), .ZN(n13139) );
  NOR3_X1 U16466 ( .A1(n14597), .A2(n13148), .A3(n13139), .ZN(n13143) );
  INV_X1 U16467 ( .A(n13242), .ZN(n13137) );
  NAND2_X1 U16468 ( .A1(n13138), .A2(n13137), .ZN(n13155) );
  INV_X1 U16469 ( .A(n13155), .ZN(n13141) );
  INV_X1 U16470 ( .A(n13139), .ZN(n14609) );
  XNOR2_X1 U16471 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13140) );
  OAI22_X1 U16472 ( .A1(n13141), .A2(n14609), .B1(n14593), .B2(n13140), .ZN(
        n13142) );
  AOI211_X1 U16473 ( .C1(n20094), .C2(n14597), .A(n13143), .B(n13142), .ZN(
        n14611) );
  NAND2_X1 U16474 ( .A1(n15634), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13144) );
  OAI21_X1 U16475 ( .B1(n15634), .B2(n14611), .A(n13144), .ZN(n15637) );
  AOI22_X1 U16476 ( .A1(n13166), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15637), .B2(n21068), .ZN(n13160) );
  INV_X1 U16477 ( .A(n13145), .ZN(n13158) );
  INV_X1 U16478 ( .A(n14597), .ZN(n13157) );
  XNOR2_X1 U16479 ( .A(n13146), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13154) );
  AOI21_X1 U16480 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13147), .A(
        n12027), .ZN(n14615) );
  NOR3_X1 U16481 ( .A1(n14597), .A2(n14615), .A3(n13148), .ZN(n13153) );
  NAND2_X1 U16482 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13151) );
  AOI211_X1 U16483 ( .C1(n13151), .C2(n13150), .A(n13149), .B(n14593), .ZN(
        n13152) );
  AOI211_X1 U16484 ( .C1(n13155), .C2(n13154), .A(n13153), .B(n13152), .ZN(
        n13156) );
  OAI21_X1 U16485 ( .B1(n13158), .B2(n13157), .A(n13156), .ZN(n14613) );
  MUX2_X1 U16486 ( .A(n14613), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15634), .Z(n15641) );
  AOI22_X1 U16487 ( .A1(n13166), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n21068), .B2(n15641), .ZN(n13159) );
  NOR2_X1 U16488 ( .A1(n13160), .A2(n13159), .ZN(n15650) );
  INV_X1 U16489 ( .A(n14600), .ZN(n13162) );
  NAND2_X1 U16490 ( .A1(n15650), .A2(n13162), .ZN(n13170) );
  INV_X1 U16491 ( .A(n20263), .ZN(n20587) );
  XNOR2_X1 U16492 ( .A(n13163), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19947) );
  AND2_X1 U16493 ( .A1(n19947), .A2(n16070), .ZN(n13165) );
  NAND2_X1 U16494 ( .A1(n15634), .A2(n16074), .ZN(n13164) );
  OAI211_X1 U16495 ( .C1(n15634), .C2(n13165), .A(n13164), .B(n21068), .ZN(
        n13168) );
  NAND2_X1 U16496 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13166), .ZN(
        n13167) );
  NAND2_X1 U16497 ( .A1(n13168), .A2(n13167), .ZN(n15649) );
  INV_X1 U16498 ( .A(n15649), .ZN(n13169) );
  NAND2_X1 U16499 ( .A1(n13170), .A2(n13169), .ZN(n13177) );
  NAND2_X1 U16500 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13172), .ZN(n16083) );
  INV_X1 U16501 ( .A(n16083), .ZN(n13171) );
  OAI21_X1 U16502 ( .B1(n13177), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13171), .ZN(
        n13173) );
  NOR2_X1 U16503 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20899) );
  NAND2_X1 U16504 ( .A1(n13173), .A2(n20175), .ZN(n20883) );
  NAND2_X1 U16505 ( .A1(n20589), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20877) );
  INV_X1 U16506 ( .A(n20877), .ZN(n14591) );
  NOR2_X1 U16507 ( .A1(n13122), .A2(n14591), .ZN(n13175) );
  NAND2_X1 U16508 ( .A1(n13020), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20742) );
  AND2_X1 U16509 ( .A1(n20742), .A2(n20741), .ZN(n20548) );
  NOR2_X1 U16510 ( .A1(n20742), .A2(n20744), .ZN(n20388) );
  MUX2_X1 U16511 ( .A(n20548), .B(n20388), .S(n20424), .Z(n13174) );
  OAI21_X1 U16512 ( .B1(n13175), .B2(n13174), .A(n20883), .ZN(n13176) );
  OAI21_X1 U16513 ( .B1(n20883), .B2(n20419), .A(n13176), .ZN(P1_U3476) );
  NOR2_X1 U16514 ( .A1(n13177), .A2(n16079), .ZN(n15659) );
  INV_X1 U16515 ( .A(n20225), .ZN(n14292) );
  OAI22_X1 U16516 ( .A1(n20185), .A2(n20744), .B1(n14292), .B2(n14591), .ZN(
        n13178) );
  OAI21_X1 U16517 ( .B1(n15659), .B2(n13178), .A(n20883), .ZN(n13179) );
  OAI21_X1 U16518 ( .B1(n20883), .B2(n20635), .A(n13179), .ZN(P1_U3478) );
  MUX2_X1 U16519 ( .A(DATAI_5_), .B(BUF1_REG_5__SCAN_IN), .S(n20102), .Z(
        n20133) );
  NAND2_X1 U16520 ( .A1(n20054), .A2(n20133), .ZN(n13333) );
  AOI22_X1 U16521 ( .A1(n20069), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20066), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13183) );
  NAND2_X1 U16522 ( .A1(n13333), .A2(n13183), .ZN(P1_U2957) );
  NAND2_X1 U16523 ( .A1(n20100), .A2(DATAI_7_), .ZN(n13185) );
  NAND2_X1 U16524 ( .A1(n20102), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13184) );
  AND2_X1 U16525 ( .A1(n13185), .A2(n13184), .ZN(n20174) );
  INV_X1 U16526 ( .A(n20174), .ZN(n14371) );
  NAND2_X1 U16527 ( .A1(n20054), .A2(n14371), .ZN(n13319) );
  AOI22_X1 U16528 ( .A1(n20069), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20066), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13186) );
  NAND2_X1 U16529 ( .A1(n13319), .A2(n13186), .ZN(P1_U2959) );
  MUX2_X1 U16530 ( .A(DATAI_4_), .B(BUF1_REG_4__SCAN_IN), .S(n20102), .Z(
        n20129) );
  NAND2_X1 U16531 ( .A1(n20054), .A2(n20129), .ZN(n13317) );
  AOI22_X1 U16532 ( .A1(n20069), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20066), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13187) );
  NAND2_X1 U16533 ( .A1(n13317), .A2(n13187), .ZN(P1_U2956) );
  MUX2_X1 U16534 ( .A(DATAI_6_), .B(BUF1_REG_6__SCAN_IN), .S(n20102), .Z(
        n20138) );
  NAND2_X1 U16535 ( .A1(n20054), .A2(n20138), .ZN(n13323) );
  AOI22_X1 U16536 ( .A1(n20069), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20066), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13188) );
  NAND2_X1 U16537 ( .A1(n13323), .A2(n13188), .ZN(P1_U2958) );
  NAND2_X1 U16538 ( .A1(n20054), .A2(n20123), .ZN(n13325) );
  AOI22_X1 U16539 ( .A1(n20069), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20066), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13189) );
  NAND2_X1 U16540 ( .A1(n13325), .A2(n13189), .ZN(P1_U2955) );
  NAND2_X1 U16541 ( .A1(n19251), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13190) );
  NOR2_X1 U16542 ( .A1(n13280), .A2(n19248), .ZN(n13527) );
  NAND2_X1 U16543 ( .A1(n13282), .A2(n13527), .ZN(n13530) );
  XOR2_X1 U16544 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13530), .Z(n13198)
         );
  OR2_X1 U16545 ( .A1(n13194), .A2(n13193), .ZN(n13195) );
  AND2_X1 U16546 ( .A1(n13195), .A2(n13309), .ZN(n19035) );
  NOR2_X1 U16547 ( .A1(n19103), .A2(n10839), .ZN(n13196) );
  AOI21_X1 U16548 ( .B1(n19035), .B2(n19103), .A(n13196), .ZN(n13197) );
  OAI21_X1 U16549 ( .B1(n13198), .B2(n19095), .A(n13197), .ZN(P2_U2882) );
  OR2_X1 U16550 ( .A1(n20114), .A2(n13199), .ZN(n13620) );
  NAND2_X1 U16551 ( .A1(n13620), .A2(n20896), .ZN(n13200) );
  OAI211_X1 U16552 ( .C1(n13201), .C2(n13200), .A(n20104), .B(n14096), .ZN(
        n13202) );
  NAND2_X1 U16553 ( .A1(n13209), .A2(n13202), .ZN(n13206) );
  NAND2_X1 U16554 ( .A1(n20114), .A2(n15697), .ZN(n13204) );
  NAND2_X1 U16555 ( .A1(n13204), .A2(n13203), .ZN(n13205) );
  NAND2_X1 U16556 ( .A1(n14126), .A2(n20114), .ZN(n13208) );
  OAI21_X1 U16557 ( .B1(n13209), .B2(n13208), .A(n13207), .ZN(n13210) );
  INV_X1 U16558 ( .A(n13210), .ZN(n13211) );
  NAND2_X1 U16559 ( .A1(n13212), .A2(n13211), .ZN(n13214) );
  NOR2_X1 U16560 ( .A1(n13245), .A2(n13246), .ZN(n13215) );
  NOR3_X1 U16561 ( .A1(n13217), .A2(n13216), .A3(n13215), .ZN(n13218) );
  INV_X1 U16562 ( .A(n13232), .ZN(n13221) );
  XNOR2_X1 U16563 ( .A(n13221), .B(n13233), .ZN(n13224) );
  INV_X1 U16564 ( .A(n20898), .ZN(n13695) );
  NAND3_X1 U16565 ( .A1(n13222), .A2(n11877), .A3(n20124), .ZN(n13223) );
  AOI21_X1 U16566 ( .B1(n13224), .B2(n13695), .A(n13223), .ZN(n13225) );
  NAND2_X1 U16567 ( .A1(n13619), .A2(n20124), .ZN(n13237) );
  OAI21_X1 U16568 ( .B1(n20898), .B2(n13232), .A(n13237), .ZN(n13226) );
  AOI21_X1 U16569 ( .B1(n13227), .B2(n13690), .A(n13226), .ZN(n20073) );
  INV_X1 U16570 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20091) );
  OR2_X1 U16571 ( .A1(n20073), .A2(n20091), .ZN(n13228) );
  NAND2_X1 U16572 ( .A1(n13267), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13231) );
  INV_X1 U16573 ( .A(n13228), .ZN(n20072) );
  NAND2_X1 U16574 ( .A1(n20072), .A2(n13229), .ZN(n13230) );
  INV_X1 U16575 ( .A(n13690), .ZN(n13701) );
  NAND2_X1 U16576 ( .A1(n13233), .A2(n13232), .ZN(n13235) );
  AND2_X1 U16577 ( .A1(n13235), .A2(n13234), .ZN(n13362) );
  NOR2_X1 U16578 ( .A1(n13235), .A2(n13234), .ZN(n13236) );
  OR2_X1 U16579 ( .A1(n13362), .A2(n13236), .ZN(n13239) );
  INV_X1 U16580 ( .A(n13237), .ZN(n13238) );
  AOI21_X1 U16581 ( .B1(n13239), .B2(n13695), .A(n13238), .ZN(n13240) );
  INV_X1 U16582 ( .A(n13260), .ZN(n13243) );
  NAND2_X1 U16583 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13369) );
  NAND2_X1 U16584 ( .A1(n13244), .A2(n13369), .ZN(n13796) );
  OAI21_X1 U16585 ( .B1(n13369), .B2(n13244), .A(n13796), .ZN(n13265) );
  INV_X1 U16586 ( .A(n13245), .ZN(n13247) );
  NAND2_X1 U16587 ( .A1(n13247), .A2(n13246), .ZN(n13248) );
  AND2_X1 U16588 ( .A1(n13249), .A2(n13248), .ZN(n13250) );
  INV_X1 U16589 ( .A(n16018), .ZN(n20084) );
  NAND2_X1 U16590 ( .A1(n13252), .A2(n13251), .ZN(n13253) );
  NAND2_X1 U16591 ( .A1(n13384), .A2(n13253), .ZN(n19984) );
  INV_X1 U16592 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20827) );
  OAI22_X1 U16593 ( .A1(n20084), .A2(n19984), .B1(n20827), .B2(n15996), .ZN(
        n13264) );
  INV_X1 U16594 ( .A(n13254), .ZN(n13257) );
  AOI21_X1 U16595 ( .B1(n13257), .B2(n13256), .A(n13255), .ZN(n13258) );
  NOR2_X1 U16596 ( .A1(n13260), .A2(n13258), .ZN(n15669) );
  NOR2_X1 U16597 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15668), .ZN(
        n13336) );
  INV_X1 U16598 ( .A(n16005), .ZN(n13259) );
  NOR2_X1 U16599 ( .A1(n12643), .A2(n13259), .ZN(n13262) );
  INV_X1 U16600 ( .A(n16003), .ZN(n16029) );
  NAND2_X1 U16601 ( .A1(n15996), .A2(n13260), .ZN(n20089) );
  NAND2_X1 U16602 ( .A1(n15669), .A2(n20091), .ZN(n20081) );
  NAND2_X1 U16603 ( .A1(n20089), .A2(n20081), .ZN(n14522) );
  AOI21_X1 U16604 ( .B1(n12643), .B2(n16029), .A(n14522), .ZN(n13370) );
  INV_X1 U16605 ( .A(n13370), .ZN(n13261) );
  MUX2_X1 U16606 ( .A(n13262), .B(n13261), .S(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n13263) );
  AOI211_X1 U16607 ( .C1(n15999), .C2(n13265), .A(n13264), .B(n13263), .ZN(
        n13266) );
  OAI21_X1 U16608 ( .B1(n16008), .B2(n14122), .A(n13266), .ZN(P1_U3029) );
  XNOR2_X1 U16609 ( .A(n13267), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13340) );
  NAND3_X1 U16610 ( .A1(n20804), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16077) );
  INV_X1 U16611 ( .A(n16077), .ZN(n13269) );
  INV_X1 U16612 ( .A(n13731), .ZN(n13276) );
  NAND2_X1 U16613 ( .A1(n20744), .A2(n13270), .ZN(n20895) );
  NAND2_X1 U16614 ( .A1(n20895), .A2(n20804), .ZN(n13271) );
  NAND2_X1 U16615 ( .A1(n20804), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13273) );
  NAND2_X1 U16616 ( .A1(n20466), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13272) );
  NAND2_X1 U16617 ( .A1(n13273), .A2(n13272), .ZN(n20075) );
  INV_X1 U16618 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20825) );
  NOR2_X1 U16619 ( .A1(n15996), .A2(n20825), .ZN(n13337) );
  AOI21_X1 U16620 ( .B1(n20076), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13337), .ZN(n13274) );
  OAI21_X1 U16621 ( .B1(n15914), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13274), .ZN(n13275) );
  AOI21_X1 U16622 ( .B1(n15909), .B2(n13276), .A(n13275), .ZN(n13277) );
  OAI21_X1 U16623 ( .B1(n13340), .B2(n19877), .A(n13277), .ZN(P1_U2998) );
  AND4_X1 U16624 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .A3(P2_INSTQUEUE_REG_0__6__SCAN_IN), 
        .A4(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13278) );
  NAND2_X1 U16625 ( .A1(n19093), .A2(n13278), .ZN(n13279) );
  NOR2_X1 U16626 ( .A1(n13280), .A2(n13279), .ZN(n13281) );
  XNOR2_X1 U16627 ( .A(n9751), .B(n19086), .ZN(n13287) );
  INV_X1 U16628 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13285) );
  OR2_X1 U16629 ( .A1(n13283), .A2(n16242), .ZN(n13284) );
  AND2_X1 U16630 ( .A1(n15236), .A2(n13284), .ZN(n16236) );
  INV_X1 U16631 ( .A(n16236), .ZN(n18991) );
  MUX2_X1 U16632 ( .A(n13285), .B(n18991), .S(n19103), .Z(n13286) );
  OAI21_X1 U16633 ( .B1(n13287), .B2(n19095), .A(n13286), .ZN(P2_U2878) );
  INV_X1 U16634 ( .A(n13488), .ZN(n13484) );
  INV_X1 U16635 ( .A(n11021), .ZN(n13288) );
  NAND2_X1 U16636 ( .A1(n13289), .A2(n13288), .ZN(n13459) );
  INV_X1 U16637 ( .A(n10399), .ZN(n13291) );
  NAND2_X1 U16638 ( .A1(n13485), .A2(n13291), .ZN(n13293) );
  INV_X1 U16639 ( .A(n10387), .ZN(n13292) );
  NAND2_X1 U16640 ( .A1(n13292), .A2(n13462), .ZN(n13453) );
  NAND2_X1 U16641 ( .A1(n13293), .A2(n13453), .ZN(n13294) );
  AOI21_X1 U16642 ( .B1(n13459), .B2(n13290), .A(n13294), .ZN(n13298) );
  NAND2_X1 U16643 ( .A1(n13296), .A2(n13295), .ZN(n13457) );
  AOI22_X1 U16644 ( .A1(n13457), .A2(n13453), .B1(n13485), .B2(n10399), .ZN(
        n13297) );
  MUX2_X1 U16645 ( .A(n13298), .B(n13297), .S(n9846), .Z(n13299) );
  OAI211_X1 U16646 ( .C1(n16272), .C2(n13484), .A(n11114), .B(n13299), .ZN(
        n13452) );
  AOI22_X1 U16647 ( .A1(n19822), .A2(n15467), .B1(n15463), .B2(n13452), .ZN(
        n13301) );
  NAND2_X1 U16648 ( .A1(n15470), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13300) );
  OAI21_X1 U16649 ( .B1(n13301), .B2(n15470), .A(n13300), .ZN(P2_U3596) );
  NOR3_X1 U16650 ( .A1(n13530), .A2(n19255), .A3(n21045), .ZN(n19094) );
  XNOR2_X1 U16651 ( .A(n19094), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13306) );
  OR2_X1 U16652 ( .A1(n13302), .A2(n13311), .ZN(n13304) );
  NAND2_X1 U16653 ( .A1(n13304), .A2(n13303), .ZN(n19012) );
  MUX2_X1 U16654 ( .A(n10848), .B(n19012), .S(n19103), .Z(n13305) );
  OAI21_X1 U16655 ( .B1(n13306), .B2(n19095), .A(n13305), .ZN(P2_U2880) );
  NOR2_X1 U16656 ( .A1(n13530), .A2(n21045), .ZN(n13308) );
  INV_X1 U16657 ( .A(n19094), .ZN(n13307) );
  OAI211_X1 U16658 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13308), .A(
        n13307), .B(n19100), .ZN(n13314) );
  NAND2_X1 U16659 ( .A1(n13310), .A2(n13309), .ZN(n13312) );
  AND2_X1 U16660 ( .A1(n13312), .A2(n10107), .ZN(n19024) );
  NAND2_X1 U16661 ( .A1(n19103), .A2(n19024), .ZN(n13313) );
  OAI211_X1 U16662 ( .C1(n19103), .C2(n13315), .A(n13314), .B(n13313), .ZN(
        P2_U2881) );
  AOI22_X1 U16663 ( .A1(n20069), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20066), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13316) );
  NAND2_X1 U16664 ( .A1(n13317), .A2(n13316), .ZN(P1_U2941) );
  AOI22_X1 U16665 ( .A1(n20069), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20066), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13318) );
  NAND2_X1 U16666 ( .A1(n13319), .A2(n13318), .ZN(P1_U2944) );
  NAND2_X1 U16667 ( .A1(n20054), .A2(n20113), .ZN(n13329) );
  AOI22_X1 U16668 ( .A1(n20069), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20066), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13320) );
  NAND2_X1 U16669 ( .A1(n13329), .A2(n13320), .ZN(P1_U2938) );
  NAND2_X1 U16670 ( .A1(n20054), .A2(n20099), .ZN(n13331) );
  AOI22_X1 U16671 ( .A1(n20069), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20066), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13321) );
  NAND2_X1 U16672 ( .A1(n13331), .A2(n13321), .ZN(P1_U2952) );
  AOI22_X1 U16673 ( .A1(n20069), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20066), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13322) );
  NAND2_X1 U16674 ( .A1(n13323), .A2(n13322), .ZN(P1_U2943) );
  AOI22_X1 U16675 ( .A1(n20069), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20066), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13324) );
  NAND2_X1 U16676 ( .A1(n13325), .A2(n13324), .ZN(P1_U2940) );
  NAND2_X1 U16677 ( .A1(n20054), .A2(n20118), .ZN(n13335) );
  AOI22_X1 U16678 ( .A1(n20069), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20066), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13326) );
  NAND2_X1 U16679 ( .A1(n13335), .A2(n13326), .ZN(P1_U2954) );
  MUX2_X1 U16680 ( .A(DATAI_11_), .B(BUF1_REG_11__SCAN_IN), .S(n20102), .Z(
        n14359) );
  NAND2_X1 U16681 ( .A1(n20054), .A2(n14359), .ZN(n20062) );
  AOI22_X1 U16682 ( .A1(n20069), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20066), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n13327) );
  NAND2_X1 U16683 ( .A1(n20062), .A2(n13327), .ZN(P1_U2948) );
  AOI22_X1 U16684 ( .A1(n20069), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20066), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13328) );
  NAND2_X1 U16685 ( .A1(n13329), .A2(n13328), .ZN(P1_U2953) );
  AOI22_X1 U16686 ( .A1(n20069), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20066), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13330) );
  NAND2_X1 U16687 ( .A1(n13331), .A2(n13330), .ZN(P1_U2937) );
  AOI22_X1 U16688 ( .A1(n20069), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20066), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13332) );
  NAND2_X1 U16689 ( .A1(n13333), .A2(n13332), .ZN(P1_U2942) );
  AOI22_X1 U16690 ( .A1(n20069), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20066), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13334) );
  NAND2_X1 U16691 ( .A1(n13335), .A2(n13334), .ZN(P1_U2939) );
  NOR3_X1 U16692 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14517), .A3(
        n13336), .ZN(n13342) );
  AOI21_X1 U16693 ( .B1(n16062), .B2(n13721), .A(n13337), .ZN(n13339) );
  NOR2_X1 U16694 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n14526), .ZN(
        n20080) );
  OAI21_X1 U16695 ( .B1(n20080), .B2(n14522), .A(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13338) );
  OAI211_X1 U16696 ( .C1(n13340), .C2(n16008), .A(n13339), .B(n13338), .ZN(
        n13341) );
  OR2_X1 U16697 ( .A1(n13342), .A2(n13341), .ZN(P1_U3030) );
  NOR2_X1 U16698 ( .A1(n13408), .A2(n13343), .ZN(n13344) );
  OR2_X1 U16699 ( .A1(n13446), .A2(n13344), .ZN(n16217) );
  NAND2_X1 U16700 ( .A1(n19086), .A2(n19085), .ZN(n13345) );
  AOI21_X1 U16701 ( .B1(n9752), .B2(n13405), .A(n13346), .ZN(n13347) );
  OR3_X1 U16702 ( .A1(n13552), .A2(n13347), .A3(n19095), .ZN(n13349) );
  NAND2_X1 U16703 ( .A1(n19089), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13348) );
  OAI211_X1 U16704 ( .C1(n16217), .C2(n19089), .A(n13349), .B(n13348), .ZN(
        P2_U2875) );
  NAND2_X1 U16705 ( .A1(n13351), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13352) );
  INV_X1 U16706 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13387) );
  OR2_X1 U16707 ( .A1(n13353), .A2(n13701), .ZN(n13356) );
  XNOR2_X1 U16708 ( .A(n13362), .B(n13361), .ZN(n13354) );
  NAND2_X1 U16709 ( .A1(n13354), .A2(n13695), .ZN(n13355) );
  NAND2_X1 U16710 ( .A1(n13356), .A2(n13355), .ZN(n13381) );
  NAND2_X1 U16711 ( .A1(n13382), .A2(n13381), .ZN(n13359) );
  NAND2_X1 U16712 ( .A1(n13357), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13358) );
  NAND2_X1 U16713 ( .A1(n13360), .A2(n13690), .ZN(n13367) );
  INV_X1 U16714 ( .A(n13361), .ZN(n13363) );
  NOR2_X1 U16715 ( .A1(n13363), .A2(n13362), .ZN(n13675) );
  INV_X1 U16716 ( .A(n13675), .ZN(n13364) );
  XNOR2_X1 U16717 ( .A(n13674), .B(n13364), .ZN(n13365) );
  NAND2_X1 U16718 ( .A1(n13695), .A2(n13365), .ZN(n13366) );
  NAND2_X1 U16719 ( .A1(n13367), .A2(n13366), .ZN(n13671) );
  INV_X1 U16720 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13368) );
  XNOR2_X1 U16721 ( .A(n13671), .B(n13368), .ZN(n13669) );
  XNOR2_X1 U16722 ( .A(n13670), .B(n13669), .ZN(n13404) );
  AOI21_X1 U16723 ( .B1(n15999), .B2(n13369), .A(n16029), .ZN(n13371) );
  OAI21_X1 U16724 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n13371), .A(
        n13370), .ZN(n13388) );
  INV_X1 U16725 ( .A(n16058), .ZN(n13374) );
  NAND2_X1 U16726 ( .A1(n13386), .A2(n13372), .ZN(n13373) );
  NAND2_X1 U16727 ( .A1(n13374), .A2(n13373), .ZN(n19950) );
  NAND3_X1 U16728 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n16005), .ZN(n16031) );
  INV_X1 U16729 ( .A(n16031), .ZN(n13375) );
  AOI21_X1 U16730 ( .B1(n15999), .B2(n13796), .A(n13375), .ZN(n16065) );
  INV_X1 U16731 ( .A(n16065), .ZN(n13798) );
  NAND2_X1 U16732 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16028) );
  OAI211_X1 U16733 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n13798), .B(n16028), .ZN(n13378) );
  AND2_X1 U16734 ( .A1(n13376), .A2(P1_REIP_REG_4__SCAN_IN), .ZN(n13399) );
  INV_X1 U16735 ( .A(n13399), .ZN(n13377) );
  OAI211_X1 U16736 ( .C1(n20084), .C2(n19950), .A(n13378), .B(n13377), .ZN(
        n13379) );
  AOI21_X1 U16737 ( .B1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13388), .A(
        n13379), .ZN(n13380) );
  OAI21_X1 U16738 ( .B1(n16008), .B2(n13404), .A(n13380), .ZN(P1_U3027) );
  XOR2_X1 U16739 ( .A(n13382), .B(n13381), .Z(n14112) );
  NAND2_X1 U16740 ( .A1(n13384), .A2(n13383), .ZN(n13385) );
  NAND2_X1 U16741 ( .A1(n13386), .A2(n13385), .ZN(n20010) );
  AOI22_X1 U16742 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13388), .B1(
        n13798), .B2(n13387), .ZN(n13389) );
  NAND2_X1 U16743 ( .A1(n13376), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n14114) );
  OAI211_X1 U16744 ( .C1(n20084), .C2(n20010), .A(n13389), .B(n14114), .ZN(
        n13390) );
  AOI21_X1 U16745 ( .B1(n14112), .B2(n20087), .A(n13390), .ZN(n13391) );
  INV_X1 U16746 ( .A(n13391), .ZN(P1_U3028) );
  AND2_X1 U16747 ( .A1(n13392), .A2(n13393), .ZN(n13395) );
  OR2_X1 U16748 ( .A1(n13395), .A2(n13394), .ZN(n20006) );
  INV_X1 U16749 ( .A(n20133), .ZN(n13396) );
  OAI222_X1 U16750 ( .A1(n20006), .A2(n14370), .B1(n14076), .B2(n13396), .C1(
        n14402), .C2(n12105), .ZN(P1_U2899) );
  INV_X1 U16751 ( .A(n13392), .ZN(n13397) );
  AOI21_X1 U16752 ( .B1(n13398), .B2(n13101), .A(n13397), .ZN(n19955) );
  INV_X1 U16753 ( .A(n19954), .ZN(n13401) );
  AOI21_X1 U16754 ( .B1(n20076), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n13399), .ZN(n13400) );
  OAI21_X1 U16755 ( .B1(n15914), .B2(n13401), .A(n13400), .ZN(n13402) );
  AOI21_X1 U16756 ( .B1(n19955), .B2(n15909), .A(n13402), .ZN(n13403) );
  OAI21_X1 U16757 ( .B1(n19877), .B2(n13404), .A(n13403), .ZN(P1_U2995) );
  XNOR2_X1 U16758 ( .A(n9752), .B(n13405), .ZN(n13412) );
  AND2_X1 U16759 ( .A1(n15238), .A2(n13407), .ZN(n13409) );
  OR2_X1 U16760 ( .A1(n13409), .A2(n13408), .ZN(n16303) );
  MUX2_X1 U16761 ( .A(n16303), .B(n13410), .S(n19089), .Z(n13411) );
  OAI21_X1 U16762 ( .B1(n13412), .B2(n19095), .A(n13411), .ZN(P2_U2876) );
  INV_X1 U16763 ( .A(n19955), .ZN(n13414) );
  INV_X1 U16764 ( .A(n20129), .ZN(n13413) );
  INV_X1 U16765 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20034) );
  OAI222_X1 U16766 ( .A1(n13414), .A2(n14370), .B1(n14076), .B2(n13413), .C1(
        n20034), .C2(n14402), .ZN(P1_U2900) );
  OAI222_X1 U16767 ( .A1(n13414), .A2(n14350), .B1(n20016), .B2(n19951), .C1(
        n19950), .C2(n20005), .ZN(P1_U2868) );
  OR2_X1 U16768 ( .A1(n13394), .A2(n13416), .ZN(n13417) );
  AND2_X1 U16769 ( .A1(n13415), .A2(n13417), .ZN(n20001) );
  INV_X1 U16770 ( .A(n20001), .ZN(n19924) );
  INV_X1 U16771 ( .A(n20138), .ZN(n13418) );
  INV_X1 U16772 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n20031) );
  OAI222_X1 U16773 ( .A1(n19924), .A2(n14370), .B1(n14076), .B2(n13418), .C1(
        n14402), .C2(n20031), .ZN(P1_U2898) );
  NOR2_X1 U16774 ( .A1(n19269), .A2(n19818), .ZN(n19599) );
  INV_X1 U16775 ( .A(n19329), .ZN(n19300) );
  NAND2_X1 U16776 ( .A1(n19599), .A2(n19300), .ZN(n13428) );
  NAND2_X1 U16777 ( .A1(n19837), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19529) );
  OR2_X1 U16778 ( .A1(n19846), .A2(n19529), .ZN(n13430) );
  INV_X1 U16779 ( .A(n19328), .ZN(n13420) );
  INV_X1 U16780 ( .A(n19529), .ZN(n13419) );
  NAND2_X1 U16781 ( .A1(n13420), .A2(n13419), .ZN(n13421) );
  INV_X1 U16782 ( .A(n13421), .ZN(n19570) );
  AND2_X1 U16783 ( .A1(n13421), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13422) );
  NAND2_X1 U16784 ( .A1(n13423), .A2(n13422), .ZN(n13432) );
  NAND2_X1 U16785 ( .A1(n16341), .A2(n13424), .ZN(n13425) );
  OAI211_X1 U16786 ( .C1(n19570), .C2(n19825), .A(n13432), .B(n19679), .ZN(
        n13427) );
  AOI21_X1 U16787 ( .B1(n13428), .B2(n13430), .A(n13427), .ZN(n19563) );
  AOI22_X1 U16788 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19260), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19261), .ZN(n19695) );
  NOR2_X2 U16789 ( .A1(n19592), .A2(n19329), .ZN(n19588) );
  AOI22_X1 U16790 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19260), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19261), .ZN(n19542) );
  AOI22_X1 U16791 ( .A1(n19559), .A2(n19539), .B1(n19588), .B2(n19692), .ZN(
        n13436) );
  OAI21_X1 U16792 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n13430), .A(n19593), 
        .ZN(n13431) );
  NAND2_X1 U16793 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19679), .ZN(n19230) );
  AND2_X1 U16794 ( .A1(n13434), .A2(n19256), .ZN(n19691) );
  AOI22_X1 U16795 ( .A1(n19571), .A2(n13433), .B1(n19691), .B2(n19570), .ZN(
        n13435) );
  OAI211_X1 U16796 ( .C1(n19563), .C2(n13437), .A(n13436), .B(n13435), .ZN(
        P2_U3138) );
  AOI22_X1 U16797 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19260), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19261), .ZN(n19607) );
  AOI22_X1 U16798 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19260), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19261), .ZN(n19684) );
  AOI22_X1 U16799 ( .A1(n19588), .A2(n19681), .B1(n19559), .B2(n19604), .ZN(
        n13439) );
  NOR2_X2 U16800 ( .A1(n19107), .A2(n19442), .ZN(n19672) );
  AND2_X1 U16801 ( .A1(n9677), .A2(n19256), .ZN(n19671) );
  AOI22_X1 U16802 ( .A1(n19571), .A2(n19672), .B1(n19671), .B2(n19570), .ZN(
        n13438) );
  OAI211_X1 U16803 ( .C1(n19563), .C2(n13440), .A(n13439), .B(n13438), .ZN(
        P2_U3136) );
  AOI22_X1 U16804 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19260), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19261), .ZN(n19654) );
  AOI22_X1 U16805 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19261), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19260), .ZN(n19713) );
  AOI22_X1 U16806 ( .A1(n19588), .A2(n19710), .B1(n19559), .B2(n19651), .ZN(
        n13443) );
  NOR2_X2 U16807 ( .A1(n19143), .A2(n19442), .ZN(n19709) );
  AOI22_X1 U16808 ( .A1(n19571), .A2(n19709), .B1(n19708), .B2(n19570), .ZN(
        n13442) );
  OAI211_X1 U16809 ( .C1(n19563), .C2(n13444), .A(n13443), .B(n13442), .ZN(
        P2_U3141) );
  XNOR2_X1 U16810 ( .A(n13552), .B(n13550), .ZN(n13451) );
  OR2_X1 U16811 ( .A1(n13446), .A2(n13445), .ZN(n13447) );
  AND2_X1 U16812 ( .A1(n13447), .A2(n13555), .ZN(n18945) );
  NOR2_X1 U16813 ( .A1(n19103), .A2(n13448), .ZN(n13449) );
  AOI21_X1 U16814 ( .B1(n18945), .B2(n19103), .A(n13449), .ZN(n13450) );
  OAI21_X1 U16815 ( .B1(n13451), .B2(n19095), .A(n13450), .ZN(P2_U2874) );
  INV_X1 U16816 ( .A(n13452), .ZN(n13493) );
  MUX2_X1 U16817 ( .A(n9846), .B(n13493), .S(n13490), .Z(n13502) );
  AND2_X1 U16818 ( .A1(n13290), .A2(n13453), .ZN(n13458) );
  INV_X1 U16819 ( .A(n13458), .ZN(n13456) );
  NOR2_X1 U16820 ( .A1(n13454), .A2(n10399), .ZN(n13455) );
  AOI22_X1 U16821 ( .A1(n13457), .A2(n13456), .B1(n13485), .B2(n13455), .ZN(
        n13461) );
  NAND2_X1 U16822 ( .A1(n13459), .A2(n13458), .ZN(n13460) );
  OAI211_X1 U16823 ( .C1(n10380), .C2(n13484), .A(n13461), .B(n13460), .ZN(
        n15464) );
  NAND2_X1 U16824 ( .A1(n13498), .A2(n13462), .ZN(n13463) );
  OAI21_X1 U16825 ( .B1(n15464), .B2(n13498), .A(n13463), .ZN(n13501) );
  AOI22_X1 U16826 ( .A1(n13467), .A2(n13466), .B1(n13465), .B2(n13464), .ZN(
        n13471) );
  NAND2_X1 U16827 ( .A1(n13469), .A2(n13468), .ZN(n13470) );
  AND2_X1 U16828 ( .A1(n13471), .A2(n13470), .ZN(n19861) );
  AOI22_X1 U16829 ( .A1(n13475), .A2(n13474), .B1(n13473), .B2(n9678), .ZN(
        n13478) );
  OAI21_X1 U16830 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(P2_MORE_REG_SCAN_IN), .A(
        n13476), .ZN(n13477) );
  AND3_X1 U16831 ( .A1(n19861), .A2(n13478), .A3(n13477), .ZN(n13500) );
  NOR2_X1 U16832 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13501), .ZN(
        n13495) );
  NAND2_X1 U16833 ( .A1(n13485), .A2(n10140), .ZN(n13483) );
  INV_X1 U16834 ( .A(n11300), .ZN(n13480) );
  NAND2_X1 U16835 ( .A1(n13480), .A2(n13479), .ZN(n13486) );
  OAI21_X1 U16836 ( .B1(n9658), .B2(n10386), .A(n13486), .ZN(n13482) );
  OAI211_X1 U16837 ( .C1(n14673), .C2(n13484), .A(n13483), .B(n13482), .ZN(
        n15460) );
  MUX2_X1 U16838 ( .A(n13486), .B(n13485), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13487) );
  AOI21_X1 U16839 ( .B1(n9647), .B2(n13488), .A(n13487), .ZN(n15452) );
  INV_X1 U16840 ( .A(n15452), .ZN(n13489) );
  AOI211_X1 U16841 ( .C1(n15460), .C2(n19846), .A(n19855), .B(n13489), .ZN(
        n13492) );
  OAI21_X1 U16842 ( .B1(n15460), .B2(n19846), .A(n13490), .ZN(n13491) );
  AOI211_X1 U16843 ( .C1(n13493), .C2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n13492), .B(n13491), .ZN(n13494) );
  AOI222_X1 U16844 ( .A1(n13495), .A2(n13494), .B1(n13495), .B2(n19837), .C1(
        n13494), .C2(n19837), .ZN(n13496) );
  OAI21_X1 U16845 ( .B1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13502), .A(
        n13496), .ZN(n13497) );
  AOI22_X1 U16846 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13498), .B1(
        n15710), .B2(n13497), .ZN(n13499) );
  OAI211_X1 U16847 ( .C1(n13502), .C2(n13501), .A(n13500), .B(n13499), .ZN(
        n16350) );
  OAI21_X1 U16848 ( .B1(n16350), .B2(P2_STATE2_REG_1__SCAN_IN), .A(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n13507) );
  INV_X1 U16849 ( .A(n13503), .ZN(n13505) );
  AOI21_X1 U16850 ( .B1(n10969), .B2(n13505), .A(n13504), .ZN(n13506) );
  NAND2_X1 U16851 ( .A1(n13507), .A2(n13506), .ZN(n16347) );
  INV_X1 U16852 ( .A(n16347), .ZN(n13508) );
  OAI21_X1 U16853 ( .B1(n13508), .B2(n16342), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13510) );
  NAND2_X1 U16854 ( .A1(n13510), .A2(n13509), .ZN(P2_U3593) );
  NAND2_X1 U16855 ( .A1(n13415), .A2(n13512), .ZN(n13513) );
  AND2_X1 U16856 ( .A1(n13511), .A2(n13513), .ZN(n19997) );
  INV_X1 U16857 ( .A(n19997), .ZN(n13515) );
  OAI222_X1 U16858 ( .A1(n13515), .A2(n14370), .B1(n14076), .B2(n20174), .C1(
        n13514), .C2(n14402), .ZN(P1_U2897) );
  OR2_X1 U16859 ( .A1(n13517), .A2(n13516), .ZN(n13519) );
  NAND2_X1 U16860 ( .A1(n13519), .A2(n13518), .ZN(n19826) );
  INV_X1 U16861 ( .A(n19826), .ZN(n13585) );
  XNOR2_X1 U16862 ( .A(n19269), .B(n13585), .ZN(n19157) );
  NAND2_X1 U16863 ( .A1(n13521), .A2(n13520), .ZN(n13523) );
  NAND2_X1 U16864 ( .A1(n13523), .A2(n10022), .ZN(n19835) );
  INV_X1 U16865 ( .A(n19831), .ZN(n15468) );
  XNOR2_X1 U16866 ( .A(n19831), .B(n19835), .ZN(n19165) );
  XNOR2_X1 U16867 ( .A(n19832), .B(n19844), .ZN(n19174) );
  NAND2_X1 U16868 ( .A1(n19174), .A2(n19173), .ZN(n19172) );
  OAI21_X1 U16869 ( .B1(n19842), .B2(n19844), .A(n19172), .ZN(n19164) );
  NAND2_X1 U16870 ( .A1(n19165), .A2(n19164), .ZN(n19163) );
  OAI21_X1 U16871 ( .B1(n19835), .B2(n15468), .A(n19163), .ZN(n19156) );
  NAND2_X1 U16872 ( .A1(n19157), .A2(n19156), .ZN(n19155) );
  NAND2_X1 U16873 ( .A1(n19269), .A2(n19826), .ZN(n13525) );
  XNOR2_X1 U16874 ( .A(n13518), .B(n13524), .ZN(n19048) );
  INV_X1 U16875 ( .A(n19048), .ZN(n13573) );
  AOI21_X1 U16876 ( .B1(n19155), .B2(n13525), .A(n13573), .ZN(n19147) );
  INV_X1 U16877 ( .A(n13527), .ZN(n13528) );
  NAND2_X1 U16878 ( .A1(n13529), .A2(n13528), .ZN(n13531) );
  OAI21_X1 U16879 ( .B1(n13526), .B2(n13531), .A(n13530), .ZN(n19146) );
  XNOR2_X1 U16880 ( .A(n19147), .B(n19146), .ZN(n13534) );
  AOI22_X1 U16881 ( .A1(n19171), .A2(n13573), .B1(n19170), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n13533) );
  NAND2_X1 U16882 ( .A1(n19161), .A2(n16184), .ZN(n13532) );
  OAI211_X1 U16883 ( .C1(n13534), .C2(n19145), .A(n13533), .B(n13532), .ZN(
        P2_U2915) );
  INV_X1 U16884 ( .A(n13541), .ZN(n13535) );
  AOI21_X1 U16885 ( .B1(n13535), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n13540) );
  NOR3_X1 U16886 ( .A1(n19837), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19382) );
  INV_X1 U16887 ( .A(n19382), .ZN(n19385) );
  NOR2_X1 U16888 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19385), .ZN(
        n19372) );
  OAI21_X1 U16889 ( .B1(n19374), .B2(n19395), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13538) );
  NOR2_X1 U16890 ( .A1(n13537), .A2(n13536), .ZN(n13595) );
  NAND2_X1 U16891 ( .A1(n13595), .A2(n19829), .ZN(n13543) );
  AOI21_X1 U16892 ( .B1(n13538), .B2(n13543), .A(n19442), .ZN(n13539) );
  INV_X1 U16893 ( .A(n19375), .ZN(n13549) );
  INV_X1 U16894 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13548) );
  OAI21_X1 U16895 ( .B1(n13541), .B2(n19372), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13542) );
  OAI21_X1 U16896 ( .B1(n13543), .B2(n19676), .A(n13542), .ZN(n19373) );
  INV_X1 U16897 ( .A(n19671), .ZN(n13781) );
  INV_X1 U16898 ( .A(n19372), .ZN(n13545) );
  AOI22_X1 U16899 ( .A1(n19395), .A2(n19681), .B1(n19374), .B2(n19604), .ZN(
        n13544) );
  OAI21_X1 U16900 ( .B1(n13781), .B2(n13545), .A(n13544), .ZN(n13546) );
  AOI21_X1 U16901 ( .B1(n19373), .B2(n19672), .A(n13546), .ZN(n13547) );
  OAI21_X1 U16902 ( .B1(n13549), .B2(n13548), .A(n13547), .ZN(P2_U3080) );
  AND2_X1 U16903 ( .A1(n13552), .A2(n13550), .ZN(n13554) );
  AND2_X1 U16904 ( .A1(n13550), .A2(n13553), .ZN(n13551) );
  OAI211_X1 U16905 ( .C1(n13554), .C2(n13553), .A(n19100), .B(n13837), .ZN(
        n13558) );
  AOI21_X1 U16906 ( .B1(n13556), .B2(n13555), .A(n13649), .ZN(n18937) );
  NAND2_X1 U16907 ( .A1(n18937), .A2(n19103), .ZN(n13557) );
  OAI211_X1 U16908 ( .C1(n19103), .C2(n13559), .A(n13558), .B(n13557), .ZN(
        P2_U2873) );
  NOR2_X1 U16909 ( .A1(n16342), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16340) );
  NOR2_X1 U16910 ( .A1(n16347), .A2(n16355), .ZN(n16345) );
  AOI21_X1 U16911 ( .B1(n19743), .B2(n16340), .A(n16345), .ZN(n13562) );
  NOR2_X1 U16912 ( .A1(n19743), .A2(n16342), .ZN(n15706) );
  AND2_X1 U16913 ( .A1(n15463), .A2(n15706), .ZN(n13560) );
  OAI21_X1 U16914 ( .B1(n16351), .B2(n13560), .A(n16347), .ZN(n13561) );
  OAI211_X1 U16915 ( .C1(n13562), .C2(n15457), .A(n19077), .B(n13561), .ZN(
        P2_U3177) );
  XNOR2_X1 U16916 ( .A(n13564), .B(n13563), .ZN(n19222) );
  XNOR2_X1 U16917 ( .A(n13566), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13567) );
  XNOR2_X1 U16918 ( .A(n13565), .B(n13567), .ZN(n19220) );
  NOR2_X1 U16919 ( .A1(n13582), .A2(n13899), .ZN(n13749) );
  INV_X1 U16920 ( .A(n14192), .ZN(n15595) );
  NAND2_X1 U16921 ( .A1(n15595), .A2(n13568), .ZN(n14187) );
  AND2_X1 U16922 ( .A1(n14187), .A2(n13569), .ZN(n13871) );
  OAI21_X1 U16923 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15401), .A(
        n13871), .ZN(n13751) );
  NOR2_X1 U16924 ( .A1(n10835), .A2(n19046), .ZN(n13570) );
  AOI221_X1 U16925 ( .B1(n13749), .B2(n13750), .C1(n13751), .C2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n13570), .ZN(n13575) );
  AOI21_X1 U16926 ( .B1(n13572), .B2(n13571), .A(n13193), .ZN(n19224) );
  AOI22_X1 U16927 ( .A1(n19224), .A2(n16316), .B1(n16312), .B2(n13573), .ZN(
        n13574) );
  OAI211_X1 U16928 ( .C1(n19220), .C2(n16339), .A(n13575), .B(n13574), .ZN(
        n13576) );
  INV_X1 U16929 ( .A(n13576), .ZN(n13577) );
  OAI21_X1 U16930 ( .B1(n16326), .B2(n19222), .A(n13577), .ZN(P2_U3042) );
  NAND2_X1 U16931 ( .A1(n13579), .A2(n13578), .ZN(n13581) );
  XNOR2_X1 U16932 ( .A(n13581), .B(n13580), .ZN(n16275) );
  INV_X1 U16933 ( .A(n16275), .ZN(n13594) );
  NOR2_X1 U16934 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n15401), .ZN(
        n13589) );
  INV_X1 U16935 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19758) );
  NOR2_X1 U16936 ( .A1(n19758), .A2(n19046), .ZN(n13584) );
  NOR2_X1 U16937 ( .A1(n13871), .A2(n13582), .ZN(n13583) );
  AOI211_X1 U16938 ( .C1(n13585), .C2(n16312), .A(n13584), .B(n13583), .ZN(
        n13586) );
  OAI21_X1 U16939 ( .B1(n16272), .B2(n16327), .A(n13586), .ZN(n13587) );
  AOI21_X1 U16940 ( .B1(n13589), .B2(n13588), .A(n13587), .ZN(n13593) );
  NAND3_X1 U16941 ( .A1(n16270), .A2(n16314), .A3(n13591), .ZN(n13592) );
  OAI211_X1 U16942 ( .C1(n13594), .C2(n16326), .A(n13593), .B(n13592), .ZN(
        P2_U3043) );
  OAI21_X1 U16943 ( .B1(n19614), .B2(n19588), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13599) );
  NAND2_X1 U16944 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13595), .ZN(
        n13600) );
  NAND3_X1 U16945 ( .A1(n19846), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19601) );
  NOR2_X1 U16946 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19601), .ZN(
        n19586) );
  INV_X1 U16947 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19825) );
  INV_X1 U16948 ( .A(n19586), .ZN(n13596) );
  AND2_X1 U16949 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n13596), .ZN(n13597) );
  OAI211_X1 U16950 ( .C1(n19586), .C2(n19825), .A(n13602), .B(n19679), .ZN(
        n13598) );
  AOI22_X1 U16951 ( .A1(n19614), .A2(n19681), .B1(n19588), .B2(n19604), .ZN(
        n13604) );
  OAI21_X1 U16952 ( .B1(n13600), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19593), 
        .ZN(n13601) );
  AND2_X1 U16953 ( .A1(n13602), .A2(n13601), .ZN(n19587) );
  AOI22_X1 U16954 ( .A1(n19587), .A2(n19672), .B1(n19671), .B2(n19586), .ZN(
        n13603) );
  OAI211_X1 U16955 ( .C1(n19591), .C2(n13851), .A(n13604), .B(n13603), .ZN(
        P2_U3144) );
  AOI22_X1 U16956 ( .A1(n19614), .A2(n19710), .B1(n19588), .B2(n19651), .ZN(
        n13606) );
  AOI22_X1 U16957 ( .A1(n19587), .A2(n19709), .B1(n19586), .B2(n19708), .ZN(
        n13605) );
  OAI211_X1 U16958 ( .C1(n19591), .C2(n14715), .A(n13606), .B(n13605), .ZN(
        P2_U3149) );
  AOI22_X1 U16959 ( .A1(n19588), .A2(n19539), .B1(n19614), .B2(n19692), .ZN(
        n13608) );
  AOI22_X1 U16960 ( .A1(n19587), .A2(n13433), .B1(n19586), .B2(n19691), .ZN(
        n13607) );
  OAI211_X1 U16961 ( .C1(n19591), .C2(n14014), .A(n13608), .B(n13607), .ZN(
        P2_U3146) );
  AOI21_X1 U16962 ( .B1(n13611), .B2(n13511), .A(n13610), .ZN(n13716) );
  INV_X1 U16963 ( .A(n13716), .ZN(n13648) );
  AND2_X1 U16964 ( .A1(n16043), .A2(n13612), .ZN(n13613) );
  NOR2_X1 U16965 ( .A1(n13737), .A2(n13613), .ZN(n16035) );
  AOI22_X1 U16966 ( .A1(n20012), .A2(n16035), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n14310), .ZN(n13614) );
  OAI21_X1 U16967 ( .B1(n13648), .B2(n14350), .A(n13614), .ZN(P1_U2864) );
  INV_X1 U16968 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n19918) );
  NAND4_X1 U16969 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n19931)
         );
  NAND2_X1 U16970 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19913) );
  NOR3_X1 U16971 ( .A1(n19918), .A2(n19931), .A3(n19913), .ZN(n13622) );
  INV_X1 U16972 ( .A(n13622), .ZN(n13645) );
  AND2_X1 U16973 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20804), .ZN(n13615) );
  NAND2_X1 U16974 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20899), .ZN(n15655) );
  INV_X1 U16975 ( .A(n15655), .ZN(n15658) );
  AOI22_X1 U16976 ( .A1(n13616), .A2(n13615), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15658), .ZN(n13617) );
  NAND2_X1 U16977 ( .A1(n15996), .A2(n13617), .ZN(n13618) );
  AND2_X1 U16978 ( .A1(n20896), .A2(n20466), .ZN(n15653) );
  NAND2_X1 U16979 ( .A1(n13620), .A2(n15653), .ZN(n13627) );
  INV_X1 U16980 ( .A(n13627), .ZN(n13621) );
  NAND2_X1 U16981 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n13622), .ZN(n19895) );
  INV_X1 U16982 ( .A(n19895), .ZN(n13623) );
  OR2_X1 U16983 ( .A1(n19965), .A2(n13623), .ZN(n13644) );
  INV_X1 U16984 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14413) );
  NAND2_X1 U16985 ( .A1(n13716), .A2(n19916), .ZN(n13643) );
  NAND2_X1 U16986 ( .A1(n20114), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13636) );
  AND2_X1 U16987 ( .A1(n13627), .A2(n13636), .ZN(n13628) );
  NAND2_X1 U16988 ( .A1(n19976), .A2(n13644), .ZN(n13630) );
  AND2_X1 U16989 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n13630), .ZN(n13631) );
  NOR2_X1 U16990 ( .A1(n19946), .A2(n13631), .ZN(n13634) );
  NOR2_X1 U16991 ( .A1(n14163), .A2(n21068), .ZN(n13632) );
  AOI22_X1 U16992 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19978), .B1(
        n19979), .B2(n13712), .ZN(n13633) );
  OAI211_X1 U16993 ( .C1(n19987), .C2(n13635), .A(n13634), .B(n13633), .ZN(
        n13641) );
  NOR2_X1 U16994 ( .A1(n13636), .A2(n15653), .ZN(n13637) );
  INV_X1 U16995 ( .A(n16035), .ZN(n13639) );
  NOR2_X1 U16996 ( .A1(n19985), .A2(n13639), .ZN(n13640) );
  NOR2_X1 U16997 ( .A1(n13641), .A2(n13640), .ZN(n13642) );
  OAI211_X1 U16998 ( .C1(n13645), .C2(n13644), .A(n13643), .B(n13642), .ZN(
        P1_U2832) );
  MUX2_X1 U16999 ( .A(DATAI_8_), .B(BUF1_REG_8__SCAN_IN), .S(n20102), .Z(
        n20043) );
  INV_X1 U17000 ( .A(n20043), .ZN(n13647) );
  OAI222_X1 U17001 ( .A1(n13648), .A2(n14370), .B1(n14076), .B2(n13647), .C1(
        n13646), .C2(n14402), .ZN(P1_U2896) );
  XNOR2_X1 U17002 ( .A(n13837), .B(n19078), .ZN(n13652) );
  OAI21_X1 U17003 ( .B1(n13650), .B2(n13649), .A(n15221), .ZN(n18924) );
  MUX2_X1 U17004 ( .A(n10821), .B(n18924), .S(n19103), .Z(n13651) );
  OAI21_X1 U17005 ( .B1(n13652), .B2(n19095), .A(n13651), .ZN(P2_U2872) );
  NAND2_X1 U17006 ( .A1(n11360), .A2(n13653), .ZN(n13654) );
  XNOR2_X1 U17007 ( .A(n16267), .B(n13654), .ZN(n13667) );
  NOR2_X1 U17008 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13655), .ZN(n13656) );
  NAND2_X1 U17009 ( .A1(n13657), .A2(n13656), .ZN(n13658) );
  NAND2_X2 U17010 ( .A1(n13659), .A2(n13658), .ZN(n19059) );
  OAI22_X1 U17011 ( .A1(n19758), .A2(n19068), .B1(n10343), .B2(n19071), .ZN(
        n13663) );
  OAI22_X1 U17012 ( .A1(n13661), .A2(n19043), .B1(n19049), .B2(n19826), .ZN(
        n13662) );
  AOI211_X1 U17013 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n19059), .A(n13663), .B(
        n13662), .ZN(n13665) );
  NAND2_X1 U17014 ( .A1(n19822), .A2(n19074), .ZN(n13664) );
  OAI211_X1 U17015 ( .C1(n19011), .C2(n16272), .A(n13665), .B(n13664), .ZN(
        n13666) );
  AOI21_X1 U17016 ( .B1(n13667), .B2(n19036), .A(n13666), .ZN(n13668) );
  INV_X1 U17017 ( .A(n13668), .ZN(P2_U2852) );
  NAND2_X1 U17018 ( .A1(n13671), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13672) );
  NAND2_X1 U17019 ( .A1(n13673), .A2(n13690), .ZN(n13678) );
  NAND2_X1 U17020 ( .A1(n13675), .A2(n13674), .ZN(n13683) );
  XNOR2_X1 U17021 ( .A(n13682), .B(n13683), .ZN(n13676) );
  NAND2_X1 U17022 ( .A1(n13695), .A2(n13676), .ZN(n13677) );
  INV_X1 U17023 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13679) );
  NAND3_X1 U17024 ( .A1(n13704), .A2(n13681), .A3(n13690), .ZN(n13688) );
  INV_X1 U17025 ( .A(n13682), .ZN(n13684) );
  NOR2_X1 U17026 ( .A1(n13684), .A2(n13683), .ZN(n13693) );
  INV_X1 U17027 ( .A(n13693), .ZN(n13685) );
  XNOR2_X1 U17028 ( .A(n13692), .B(n13685), .ZN(n13686) );
  NAND2_X1 U17029 ( .A1(n13695), .A2(n13686), .ZN(n13687) );
  NAND2_X1 U17030 ( .A1(n13688), .A2(n13687), .ZN(n13689) );
  OR2_X1 U17031 ( .A1(n13689), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15906) );
  NAND2_X1 U17032 ( .A1(n13689), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15905) );
  NAND2_X1 U17033 ( .A1(n13691), .A2(n13690), .ZN(n13697) );
  NAND2_X1 U17034 ( .A1(n13693), .A2(n13692), .ZN(n13706) );
  XNOR2_X1 U17035 ( .A(n13708), .B(n13706), .ZN(n13694) );
  NAND2_X1 U17036 ( .A1(n13695), .A2(n13694), .ZN(n13696) );
  OR2_X1 U17037 ( .A1(n15900), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13698) );
  OR2_X1 U17038 ( .A1(n13700), .A2(n20804), .ZN(n13702) );
  NOR2_X1 U17039 ( .A1(n13702), .A2(n13701), .ZN(n13703) );
  INV_X1 U17040 ( .A(n13706), .ZN(n13707) );
  NAND2_X1 U17041 ( .A1(n13708), .A2(n13707), .ZN(n13709) );
  OR2_X1 U17042 ( .A1(n20898), .A2(n13709), .ZN(n13710) );
  NAND2_X1 U17043 ( .A1(n13705), .A2(n13710), .ZN(n13790) );
  XNOR2_X1 U17044 ( .A(n13790), .B(n16039), .ZN(n13711) );
  XNOR2_X1 U17045 ( .A(n13789), .B(n13711), .ZN(n16033) );
  INV_X1 U17046 ( .A(n13712), .ZN(n13714) );
  AOI22_X1 U17047 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n13376), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13713) );
  OAI21_X1 U17048 ( .B1(n15914), .B2(n13714), .A(n13713), .ZN(n13715) );
  AOI21_X1 U17049 ( .B1(n13716), .B2(n15909), .A(n13715), .ZN(n13717) );
  OAI21_X1 U17050 ( .B1(n16033), .B2(n19877), .A(n13717), .ZN(P1_U2991) );
  INV_X1 U17051 ( .A(n13718), .ZN(n13723) );
  NAND2_X1 U17052 ( .A1(n13723), .A2(n13719), .ZN(n13720) );
  AOI22_X1 U17053 ( .A1(n19940), .A2(n13721), .B1(n19932), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13730) );
  NAND2_X1 U17054 ( .A1(n13723), .A2(n13722), .ZN(n19981) );
  AOI22_X1 U17055 ( .A1(n19979), .A2(n13725), .B1(n19960), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n13727) );
  NAND2_X1 U17056 ( .A1(n19978), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13726) );
  OAI211_X1 U17057 ( .C1(n19981), .C2(n20673), .A(n13727), .B(n13726), .ZN(
        n13728) );
  AOI21_X1 U17058 ( .B1(n19961), .B2(n20825), .A(n13728), .ZN(n13729) );
  OAI211_X1 U17059 ( .C1(n19937), .C2(n13731), .A(n13730), .B(n13729), .ZN(
        P1_U2839) );
  AND2_X1 U17060 ( .A1(n13734), .A2(n13733), .ZN(n13735) );
  NOR2_X1 U17061 ( .A1(n13732), .A2(n13735), .ZN(n19903) );
  INV_X1 U17062 ( .A(n19903), .ZN(n13742) );
  INV_X1 U17063 ( .A(n14076), .ZN(n13964) );
  MUX2_X1 U17064 ( .A(DATAI_9_), .B(BUF1_REG_9__SCAN_IN), .S(n20102), .Z(
        n20045) );
  AOI22_X1 U17065 ( .A1(n13964), .A2(n20045), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n14397), .ZN(n13736) );
  OAI21_X1 U17066 ( .B1(n13742), .B2(n14370), .A(n13736), .ZN(P1_U2895) );
  INV_X1 U17067 ( .A(n13737), .ZN(n13739) );
  INV_X1 U17068 ( .A(n13765), .ZN(n13738) );
  AOI21_X1 U17069 ( .B1(n13740), .B2(n13739), .A(n13738), .ZN(n19901) );
  AOI22_X1 U17070 ( .A1(n20012), .A2(n19901), .B1(P1_EBX_REG_9__SCAN_IN), .B2(
        n14310), .ZN(n13741) );
  OAI21_X1 U17071 ( .B1(n13742), .B2(n14350), .A(n13741), .ZN(P1_U2863) );
  XOR2_X1 U17072 ( .A(n13744), .B(n13743), .Z(n16264) );
  INV_X1 U17073 ( .A(n16264), .ZN(n13761) );
  NAND2_X1 U17074 ( .A1(n13747), .A2(n13746), .ZN(n13748) );
  XNOR2_X1 U17075 ( .A(n13745), .B(n13748), .ZN(n16263) );
  OAI221_X1 U17076 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n13750), .C2(n10796), .A(
        n13749), .ZN(n13758) );
  AOI22_X1 U17077 ( .A1(n19217), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n13751), .ZN(n13757) );
  NAND2_X1 U17078 ( .A1(n16316), .A2(n19035), .ZN(n13756) );
  OAI21_X1 U17079 ( .B1(n9794), .B2(n13753), .A(n13752), .ZN(n19150) );
  INV_X1 U17080 ( .A(n19150), .ZN(n13754) );
  NAND2_X1 U17081 ( .A1(n13754), .A2(n16312), .ZN(n13755) );
  NAND4_X1 U17082 ( .A1(n13758), .A2(n13757), .A3(n13756), .A4(n13755), .ZN(
        n13759) );
  AOI21_X1 U17083 ( .B1(n16263), .B2(n16314), .A(n13759), .ZN(n13760) );
  OAI21_X1 U17084 ( .B1(n13761), .B2(n16326), .A(n13760), .ZN(P2_U3041) );
  OAI21_X1 U17085 ( .B1(n13732), .B2(n13763), .A(n10079), .ZN(n14516) );
  NAND2_X1 U17086 ( .A1(n13765), .A2(n13764), .ZN(n13766) );
  NAND2_X1 U17087 ( .A1(n13889), .A2(n13766), .ZN(n13772) );
  INV_X1 U17088 ( .A(n13772), .ZN(n16017) );
  AOI22_X1 U17089 ( .A1(n20012), .A2(n16017), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14310), .ZN(n13767) );
  OAI21_X1 U17090 ( .B1(n14516), .B2(n14350), .A(n13767), .ZN(P1_U2862) );
  INV_X1 U17091 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n20836) );
  AOI211_X1 U17092 ( .C1(n19961), .C2(n19895), .A(n19960), .B(n20836), .ZN(
        n19907) );
  NAND2_X1 U17093 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n15812) );
  NOR2_X1 U17094 ( .A1(n19895), .A2(n15812), .ZN(n13993) );
  OAI21_X1 U17095 ( .B1(n13993), .B2(n19965), .A(n19976), .ZN(n15817) );
  OAI21_X1 U17096 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n19907), .A(n15817), 
        .ZN(n13776) );
  AOI21_X1 U17097 ( .B1(n19978), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19946), .ZN(n13770) );
  INV_X1 U17098 ( .A(n14512), .ZN(n13768) );
  NAND2_X1 U17099 ( .A1(n19979), .A2(n13768), .ZN(n13769) );
  OAI211_X1 U17100 ( .C1(n19987), .C2(n13771), .A(n13770), .B(n13769), .ZN(
        n13774) );
  NOR2_X1 U17101 ( .A1(n19985), .A2(n13772), .ZN(n13773) );
  NOR2_X1 U17102 ( .A1(n13774), .A2(n13773), .ZN(n13775) );
  OAI211_X1 U17103 ( .C1(n14516), .C2(n19923), .A(n13776), .B(n13775), .ZN(
        P1_U2830) );
  OAI21_X1 U17104 ( .B1(n19725), .B2(n19286), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13777) );
  NAND2_X1 U17105 ( .A1(n13777), .A2(n19830), .ZN(n13786) );
  INV_X1 U17106 ( .A(n13786), .ZN(n13779) );
  NAND2_X1 U17107 ( .A1(n19829), .A2(n19837), .ZN(n19330) );
  OR2_X1 U17108 ( .A1(n19330), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19270) );
  NOR2_X1 U17109 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19270), .ZN(
        n19258) );
  INV_X1 U17110 ( .A(n19258), .ZN(n13780) );
  AND2_X1 U17111 ( .A1(n19675), .A2(n13780), .ZN(n13785) );
  AOI211_X1 U17112 ( .C1(n13783), .C2(n19825), .A(n19830), .B(n19258), .ZN(
        n13778) );
  OAI22_X1 U17113 ( .A1(n19607), .A2(n19294), .B1(n13781), .B2(n13780), .ZN(
        n13782) );
  AOI21_X1 U17114 ( .B1(n19725), .B2(n19604), .A(n13782), .ZN(n13788) );
  OAI21_X1 U17115 ( .B1(n13783), .B2(n19258), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13784) );
  NAND2_X1 U17116 ( .A1(n19262), .A2(n19672), .ZN(n13787) );
  OAI211_X1 U17117 ( .C1(n19266), .C2(n13846), .A(n13788), .B(n13787), .ZN(
        P2_U3048) );
  INV_X4 U17118 ( .A(n15855), .ZN(n14470) );
  INV_X1 U17119 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16022) );
  XNOR2_X1 U17120 ( .A(n14470), .B(n16022), .ZN(n13791) );
  XNOR2_X1 U17121 ( .A(n13927), .B(n13791), .ZN(n13803) );
  NOR2_X1 U17122 ( .A1(n15996), .A2(n20836), .ZN(n13800) );
  AOI21_X1 U17123 ( .B1(n20076), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n13800), .ZN(n13793) );
  NAND2_X1 U17124 ( .A1(n15889), .A2(n19902), .ZN(n13792) );
  NAND2_X1 U17125 ( .A1(n13793), .A2(n13792), .ZN(n13794) );
  AOI21_X1 U17126 ( .B1(n19903), .B2(n15909), .A(n13794), .ZN(n13795) );
  OAI21_X1 U17127 ( .B1(n13803), .B2(n19877), .A(n13795), .ZN(P1_U2990) );
  NOR2_X1 U17128 ( .A1(n13679), .A2(n16028), .ZN(n13799) );
  NAND2_X1 U17129 ( .A1(n13799), .A2(n13796), .ZN(n13942) );
  AOI21_X1 U17130 ( .B1(n15999), .B2(n13942), .A(n14522), .ZN(n16026) );
  NAND3_X1 U17131 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n13799), .ZN(n13943) );
  NAND3_X1 U17132 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13941) );
  AOI21_X1 U17133 ( .B1(n16029), .B2(n13943), .A(n13941), .ZN(n13797) );
  AND2_X1 U17134 ( .A1(n20089), .A2(n14517), .ZN(n14524) );
  AOI21_X1 U17135 ( .B1(n16026), .B2(n13797), .A(n14524), .ZN(n16020) );
  NAND2_X1 U17136 ( .A1(n13799), .A2(n13798), .ZN(n16056) );
  NOR2_X1 U17137 ( .A1(n13941), .A2(n16056), .ZN(n16021) );
  AOI22_X1 U17138 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n16020), .B1(
        n16021), .B2(n16022), .ZN(n13802) );
  AOI21_X1 U17139 ( .B1(n16018), .B2(n19901), .A(n13800), .ZN(n13801) );
  OAI211_X1 U17140 ( .C1(n13803), .C2(n16008), .A(n13802), .B(n13801), .ZN(
        P1_U3022) );
  MUX2_X1 U17141 ( .A(DATAI_10_), .B(BUF1_REG_10__SCAN_IN), .S(n20102), .Z(
        n20047) );
  INV_X1 U17142 ( .A(n20047), .ZN(n13805) );
  OAI222_X1 U17143 ( .A1(n14516), .A2(n14370), .B1(n14076), .B2(n13805), .C1(
        n13804), .C2(n14402), .ZN(P1_U2894) );
  OAI21_X1 U17144 ( .B1(n13806), .B2(n13808), .A(n13807), .ZN(n15618) );
  INV_X1 U17145 ( .A(n19109), .ZN(n15084) );
  OAI22_X1 U17146 ( .A1(n15084), .A2(n19232), .B1(n13810), .B2(n19169), .ZN(
        n13815) );
  INV_X1 U17147 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n13813) );
  NOR2_X1 U17148 ( .A1(n15086), .A2(n13813), .ZN(n13814) );
  AOI211_X1 U17149 ( .C1(BUF1_REG_17__SCAN_IN), .C2(n19110), .A(n13815), .B(
        n13814), .ZN(n13863) );
  AOI22_X1 U17150 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13819) );
  NAND2_X1 U17151 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n13818) );
  NAND2_X1 U17152 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n13817) );
  NAND2_X1 U17153 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n13816) );
  NAND4_X1 U17154 ( .A1(n13819), .A2(n13818), .A3(n13817), .A4(n13816), .ZN(
        n13823) );
  OAI22_X1 U17155 ( .A1(n13821), .A2(n10464), .B1(n10463), .B2(n13820), .ZN(
        n13822) );
  NOR2_X1 U17156 ( .A1(n13823), .A2(n13822), .ZN(n13836) );
  OR2_X1 U17157 ( .A1(n10467), .A2(n19236), .ZN(n13827) );
  AOI22_X1 U17158 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13826) );
  NAND2_X1 U17159 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n13825) );
  NAND2_X1 U17160 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n13824) );
  AND4_X1 U17161 ( .A1(n13827), .A2(n13826), .A3(n13825), .A4(n13824), .ZN(
        n13835) );
  OAI22_X1 U17162 ( .A1(n10472), .A2(n13829), .B1(n14738), .B2(n13828), .ZN(
        n13833) );
  OAI22_X1 U17163 ( .A1(n13831), .A2(n11114), .B1(n10473), .B2(n13830), .ZN(
        n13832) );
  NOR2_X1 U17164 ( .A1(n13833), .A2(n13832), .ZN(n13834) );
  AOI22_X1 U17165 ( .A1(n14783), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13841) );
  NAND2_X1 U17166 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n13840) );
  NAND2_X1 U17167 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n13839) );
  NAND2_X1 U17168 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n13838) );
  NAND4_X1 U17169 ( .A1(n13841), .A2(n13840), .A3(n13839), .A4(n13838), .ZN(
        n13845) );
  INV_X1 U17170 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13842) );
  OAI22_X1 U17171 ( .A1(n10463), .A2(n13843), .B1(n10464), .B2(n13842), .ZN(
        n13844) );
  NOR2_X1 U17172 ( .A1(n13845), .A2(n13844), .ZN(n13859) );
  OR2_X1 U17173 ( .A1(n10467), .A2(n13846), .ZN(n13850) );
  AOI22_X1 U17174 ( .A1(n14767), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13849) );
  NAND2_X1 U17175 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n13848) );
  NAND2_X1 U17176 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n13847) );
  AND4_X1 U17177 ( .A1(n13850), .A2(n13849), .A3(n13848), .A4(n13847), .ZN(
        n13858) );
  OAI22_X1 U17178 ( .A1(n10472), .A2(n13852), .B1(n14738), .B2(n13851), .ZN(
        n13856) );
  OAI22_X1 U17179 ( .A1(n10473), .A2(n13854), .B1(n11114), .B2(n13853), .ZN(
        n13855) );
  NOR2_X1 U17180 ( .A1(n13856), .A2(n13855), .ZN(n13857) );
  AND3_X1 U17181 ( .A1(n13859), .A2(n13858), .A3(n13857), .ZN(n19079) );
  AOI21_X1 U17182 ( .B1(n13861), .B2(n13860), .A(n16179), .ZN(n13880) );
  NAND2_X1 U17183 ( .A1(n13880), .A2(n19175), .ZN(n13862) );
  OAI211_X1 U17184 ( .C1(n15618), .C2(n19153), .A(n13863), .B(n13862), .ZN(
        P2_U2902) );
  XNOR2_X1 U17185 ( .A(n13864), .B(n13865), .ZN(n16258) );
  NAND2_X1 U17186 ( .A1(n13867), .A2(n13866), .ZN(n13868) );
  XNOR2_X1 U17187 ( .A(n13868), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16259) );
  INV_X1 U17188 ( .A(n16259), .ZN(n13878) );
  XNOR2_X1 U17189 ( .A(n13870), .B(n13869), .ZN(n19142) );
  NOR2_X1 U17190 ( .A1(n13900), .A2(n13899), .ZN(n13874) );
  OAI21_X1 U17191 ( .B1(n15401), .B2(n13872), .A(n13871), .ZN(n16313) );
  INV_X1 U17192 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19762) );
  NOR2_X1 U17193 ( .A1(n19762), .A2(n19046), .ZN(n13873) );
  AOI221_X1 U17194 ( .B1(n13874), .B2(n13901), .C1(n16313), .C2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n13873), .ZN(n13876) );
  NAND2_X1 U17195 ( .A1(n16316), .A2(n19024), .ZN(n13875) );
  OAI211_X1 U17196 ( .C1(n16330), .C2(n19142), .A(n13876), .B(n13875), .ZN(
        n13877) );
  AOI21_X1 U17197 ( .B1(n13878), .B2(n16314), .A(n13877), .ZN(n13879) );
  OAI21_X1 U17198 ( .B1(n16326), .B2(n16258), .A(n13879), .ZN(P2_U3040) );
  NAND2_X1 U17199 ( .A1(n13880), .A2(n19100), .ZN(n13885) );
  AND2_X1 U17200 ( .A1(n15223), .A2(n13881), .ZN(n13882) );
  OR2_X1 U17201 ( .A1(n13882), .A2(n15194), .ZN(n15620) );
  INV_X1 U17202 ( .A(n15620), .ZN(n13883) );
  NAND2_X1 U17203 ( .A1(n13883), .A2(n19103), .ZN(n13884) );
  OAI211_X1 U17204 ( .C1(n13920), .C2(n19103), .A(n13885), .B(n13884), .ZN(
        P2_U2870) );
  OR2_X1 U17205 ( .A1(n13762), .A2(n13887), .ZN(n13888) );
  NAND2_X1 U17206 ( .A1(n13886), .A2(n13888), .ZN(n13953) );
  XNOR2_X1 U17207 ( .A(n13953), .B(n13951), .ZN(n15896) );
  INV_X1 U17208 ( .A(n15896), .ZN(n13894) );
  AOI21_X1 U17209 ( .B1(n13890), .B2(n13889), .A(n9784), .ZN(n16010) );
  AOI22_X1 U17210 ( .A1(n20012), .A2(n16010), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n14310), .ZN(n13891) );
  OAI21_X1 U17211 ( .B1(n13894), .B2(n14350), .A(n13891), .ZN(P1_U2861) );
  INV_X1 U17212 ( .A(n14359), .ZN(n13893) );
  OAI222_X1 U17213 ( .A1(n13894), .A2(n14370), .B1(n14076), .B2(n13893), .C1(
        n13892), .C2(n14402), .ZN(P1_U2893) );
  XNOR2_X1 U17214 ( .A(n13895), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13915) );
  INV_X1 U17215 ( .A(n16247), .ZN(n13897) );
  NAND2_X1 U17216 ( .A1(n13897), .A2(n16248), .ZN(n13898) );
  XNOR2_X1 U17217 ( .A(n13896), .B(n13898), .ZN(n13913) );
  NOR3_X1 U17218 ( .A1(n13901), .A2(n13900), .A3(n13899), .ZN(n16319) );
  INV_X1 U17219 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19764) );
  NOR2_X1 U17220 ( .A1(n19764), .A2(n19046), .ZN(n13902) );
  AOI221_X1 U17221 ( .B1(n16319), .B2(n9956), .C1(n16313), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n13902), .ZN(n13903) );
  INV_X1 U17222 ( .A(n13903), .ZN(n13908) );
  OR2_X1 U17223 ( .A1(n13905), .A2(n13904), .ZN(n13906) );
  NAND2_X1 U17224 ( .A1(n13906), .A2(n16310), .ZN(n19141) );
  OAI22_X1 U17225 ( .A1(n19141), .A2(n16330), .B1(n16327), .B2(n19012), .ZN(
        n13907) );
  AOI211_X1 U17226 ( .C1(n13913), .C2(n16317), .A(n13908), .B(n13907), .ZN(
        n13909) );
  OAI21_X1 U17227 ( .B1(n13915), .B2(n16339), .A(n13909), .ZN(P2_U3039) );
  OAI22_X1 U17228 ( .A1(n10847), .A2(n16278), .B1(n19764), .B2(n19046), .ZN(
        n13912) );
  INV_X1 U17229 ( .A(n19007), .ZN(n13910) );
  OAI22_X1 U17230 ( .A1(n16273), .A2(n19012), .B1(n19229), .B2(n13910), .ZN(
        n13911) );
  AOI211_X1 U17231 ( .C1(n13913), .C2(n11389), .A(n13912), .B(n13911), .ZN(
        n13914) );
  OAI21_X1 U17232 ( .B1(n13915), .B2(n19219), .A(n13914), .ZN(P2_U3007) );
  NAND2_X1 U17233 ( .A1(n11360), .A2(n13916), .ZN(n13917) );
  XOR2_X1 U17234 ( .A(n13918), .B(n13917), .Z(n13925) );
  OAI21_X1 U17235 ( .B1(n19784), .B2(n19068), .A(n19046), .ZN(n13922) );
  INV_X1 U17236 ( .A(n19059), .ZN(n19001) );
  OAI22_X1 U17237 ( .A1(n19001), .A2(n13920), .B1(n13919), .B2(n19043), .ZN(
        n13921) );
  AOI211_X1 U17238 ( .C1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n19028), .A(
        n13922), .B(n13921), .ZN(n13923) );
  OAI21_X1 U17239 ( .B1(n15620), .B2(n19011), .A(n13923), .ZN(n13924) );
  AOI21_X1 U17240 ( .B1(n13925), .B2(n19036), .A(n13924), .ZN(n13926) );
  OAI21_X1 U17241 ( .B1(n15618), .B2(n19049), .A(n13926), .ZN(P2_U2838) );
  NAND2_X1 U17242 ( .A1(n15831), .A2(n16022), .ZN(n13928) );
  NOR2_X1 U17243 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14491) );
  AND2_X1 U17244 ( .A1(n14491), .A2(n13931), .ZN(n13929) );
  NAND2_X1 U17245 ( .A1(n13982), .A2(n14051), .ZN(n13935) );
  INV_X1 U17246 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15993) );
  NAND2_X1 U17247 ( .A1(n15831), .A2(n15993), .ZN(n13930) );
  NAND2_X1 U17248 ( .A1(n13976), .A2(n13930), .ZN(n14497) );
  NAND2_X1 U17249 ( .A1(n13705), .A2(n13931), .ZN(n14495) );
  NAND2_X1 U17250 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n13932) );
  NAND2_X1 U17251 ( .A1(n15831), .A2(n13932), .ZN(n14493) );
  NAND2_X1 U17252 ( .A1(n14495), .A2(n14493), .ZN(n13933) );
  INV_X1 U17253 ( .A(n13976), .ZN(n13934) );
  AOI21_X1 U17254 ( .B1(n13935), .B2(n9776), .A(n13934), .ZN(n13937) );
  XNOR2_X1 U17255 ( .A(n14470), .B(n14059), .ZN(n13936) );
  XNOR2_X1 U17256 ( .A(n13937), .B(n13936), .ZN(n13974) );
  INV_X1 U17257 ( .A(n14072), .ZN(n13938) );
  AOI21_X1 U17258 ( .B1(n13939), .B2(n13995), .A(n13938), .ZN(n14282) );
  INV_X1 U17259 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n13940) );
  NOR2_X1 U17260 ( .A1(n15996), .A2(n13940), .ZN(n13969) );
  OR3_X1 U17261 ( .A1(n14508), .A2(n16022), .A3(n13941), .ZN(n16000) );
  NOR2_X1 U17262 ( .A1(n16000), .A2(n13942), .ZN(n13944) );
  NAND4_X1 U17263 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n15999), .A4(n13944), .ZN(
        n15670) );
  NOR2_X1 U17264 ( .A1(n13943), .A2(n16000), .ZN(n16002) );
  NAND3_X1 U17265 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n16002), .ZN(n15985) );
  NOR2_X1 U17266 ( .A1(n15993), .A2(n15985), .ZN(n14520) );
  NAND2_X1 U17267 ( .A1(n14520), .A2(n16005), .ZN(n14583) );
  OAI21_X1 U17268 ( .B1(n15993), .B2(n15670), .A(n14583), .ZN(n14532) );
  INV_X1 U17269 ( .A(n13944), .ZN(n13946) );
  NAND3_X1 U17270 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n13945) );
  NOR2_X1 U17271 ( .A1(n13946), .A2(n13945), .ZN(n14521) );
  OAI22_X1 U17272 ( .A1(n16003), .A2(n14520), .B1(n14521), .B2(n14526), .ZN(
        n13947) );
  NOR2_X1 U17273 ( .A1(n14522), .A2(n13947), .ZN(n15994) );
  INV_X1 U17274 ( .A(n15994), .ZN(n13948) );
  MUX2_X1 U17275 ( .A(n14532), .B(n13948), .S(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n13949) );
  AOI211_X1 U17276 ( .C1(n16062), .C2(n14282), .A(n13969), .B(n13949), .ZN(
        n13950) );
  OAI21_X1 U17277 ( .B1(n13974), .B2(n16008), .A(n13950), .ZN(P1_U3017) );
  INV_X1 U17278 ( .A(n13951), .ZN(n13952) );
  OAI21_X1 U17279 ( .B1(n13953), .B2(n13952), .A(n13886), .ZN(n13955) );
  AND2_X1 U17280 ( .A1(n13955), .A2(n13954), .ZN(n13992) );
  NOR2_X1 U17281 ( .A1(n13955), .A2(n13954), .ZN(n13956) );
  NOR2_X1 U17282 ( .A1(n9784), .A2(n13957), .ZN(n13958) );
  AOI22_X1 U17283 ( .A1(n20012), .A2(n9783), .B1(P1_EBX_REG_12__SCAN_IN), .B2(
        n14310), .ZN(n13959) );
  OAI21_X1 U17284 ( .B1(n15886), .B2(n14350), .A(n13959), .ZN(P1_U2860) );
  INV_X1 U17285 ( .A(n13961), .ZN(n13962) );
  AOI21_X1 U17286 ( .B1(n13963), .B2(n13960), .A(n13962), .ZN(n13972) );
  INV_X1 U17287 ( .A(n13972), .ZN(n14290) );
  MUX2_X1 U17288 ( .A(DATAI_14_), .B(BUF1_REG_14__SCAN_IN), .S(n20102), .Z(
        n20053) );
  AOI22_X1 U17289 ( .A1(n13964), .A2(n20053), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14397), .ZN(n13965) );
  OAI21_X1 U17290 ( .B1(n14290), .B2(n14370), .A(n13965), .ZN(P1_U2890) );
  AOI22_X1 U17291 ( .A1(n14282), .A2(n20012), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n14310), .ZN(n13966) );
  OAI21_X1 U17292 ( .B1(n14290), .B2(n14350), .A(n13966), .ZN(P1_U2858) );
  MUX2_X1 U17293 ( .A(DATAI_12_), .B(BUF1_REG_12__SCAN_IN), .S(n20102), .Z(
        n20049) );
  INV_X1 U17294 ( .A(n20049), .ZN(n13968) );
  OAI222_X1 U17295 ( .A1(n15886), .A2(n14370), .B1(n14076), .B2(n13968), .C1(
        n13967), .C2(n14402), .ZN(P1_U2892) );
  AOI21_X1 U17296 ( .B1(n20076), .B2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n13969), .ZN(n13970) );
  OAI21_X1 U17297 ( .B1(n15914), .B2(n14280), .A(n13970), .ZN(n13971) );
  AOI21_X1 U17298 ( .B1(n13972), .B2(n15909), .A(n13971), .ZN(n13973) );
  OAI21_X1 U17299 ( .B1(n13974), .B2(n19877), .A(n13973), .ZN(P1_U2985) );
  OR2_X1 U17300 ( .A1(n13705), .A2(n14059), .ZN(n13975) );
  INV_X1 U17301 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n13977) );
  NAND2_X1 U17302 ( .A1(n15831), .A2(n13977), .ZN(n15874) );
  NAND2_X1 U17303 ( .A1(n14053), .A2(n14051), .ZN(n15862) );
  NOR2_X1 U17304 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13978) );
  NOR2_X1 U17305 ( .A1(n15831), .A2(n13978), .ZN(n13979) );
  NOR2_X1 U17306 ( .A1(n15862), .A2(n13979), .ZN(n13980) );
  XNOR2_X1 U17307 ( .A(n14470), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13983) );
  OR2_X1 U17308 ( .A1(n14146), .A2(n13983), .ZN(n14481) );
  NAND3_X1 U17309 ( .A1(n14481), .A2(n15853), .A3(n20087), .ZN(n13990) );
  INV_X1 U17310 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15969) );
  NOR4_X1 U17311 ( .A1(n13977), .A2(n14059), .A3(n15863), .A4(n15969), .ZN(
        n13986) );
  OAI21_X1 U17312 ( .B1(n14517), .B2(n13986), .A(n15994), .ZN(n15974) );
  NAND2_X1 U17313 ( .A1(n9764), .A2(n13984), .ZN(n13985) );
  AND2_X1 U17314 ( .A1(n9716), .A2(n13985), .ZN(n14346) );
  INV_X1 U17315 ( .A(n14346), .ZN(n14260) );
  NAND2_X1 U17316 ( .A1(n13376), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14477) );
  OAI21_X1 U17317 ( .B1(n14260), .B2(n20084), .A(n14477), .ZN(n13988) );
  INV_X1 U17318 ( .A(n14532), .ZN(n15971) );
  INV_X1 U17319 ( .A(n13986), .ZN(n14519) );
  NOR3_X1 U17320 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15971), .A3(
        n14519), .ZN(n13987) );
  AOI211_X1 U17321 ( .C1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n15974), .A(
        n13988), .B(n13987), .ZN(n13989) );
  NAND2_X1 U17322 ( .A1(n13990), .A2(n13989), .ZN(P1_U3013) );
  OAI21_X1 U17323 ( .B1(n13992), .B2(n13991), .A(n13960), .ZN(n14504) );
  INV_X1 U17324 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n20839) );
  NAND2_X1 U17325 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n13993), .ZN(n15807) );
  NOR2_X1 U17326 ( .A1(n20839), .A2(n15807), .ZN(n14101) );
  OAI21_X1 U17327 ( .B1(n14101), .B2(n19965), .A(n19976), .ZN(n15809) );
  AOI21_X1 U17328 ( .B1(n14501), .B2(n19979), .A(n19946), .ZN(n13994) );
  OAI21_X1 U17329 ( .B1(n14499), .B2(n19898), .A(n13994), .ZN(n14002) );
  NAND2_X1 U17330 ( .A1(n19961), .A2(n14101), .ZN(n14000) );
  OAI21_X1 U17331 ( .B1(n13997), .B2(n13996), .A(n13995), .ZN(n15986) );
  INV_X1 U17332 ( .A(n15986), .ZN(n13998) );
  AOI22_X1 U17333 ( .A1(n19940), .A2(n13998), .B1(n19932), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n13999) );
  OAI21_X1 U17334 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n14000), .A(n13999), 
        .ZN(n14001) );
  AOI211_X1 U17335 ( .C1(n15809), .C2(P1_REIP_REG_13__SCAN_IN), .A(n14002), 
        .B(n14001), .ZN(n14003) );
  OAI21_X1 U17336 ( .B1(n14504), .B2(n19923), .A(n14003), .ZN(P1_U2827) );
  AOI22_X1 U17337 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14007) );
  NAND2_X1 U17338 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n14006) );
  NAND2_X1 U17339 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n14005) );
  NAND2_X1 U17340 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n14004) );
  NAND4_X1 U17341 ( .A1(n14007), .A2(n14006), .A3(n14005), .A4(n14004), .ZN(
        n14011) );
  INV_X1 U17342 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14009) );
  OAI22_X1 U17343 ( .A1(n14009), .A2(n10464), .B1(n10463), .B2(n14008), .ZN(
        n14010) );
  NOR2_X1 U17344 ( .A1(n14011), .A2(n14010), .ZN(n14023) );
  AOI22_X1 U17345 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14012) );
  OAI21_X1 U17346 ( .B1(n10467), .B2(n19239), .A(n14012), .ZN(n14013) );
  INV_X1 U17347 ( .A(n14013), .ZN(n14022) );
  OAI22_X1 U17348 ( .A1(n10472), .A2(n14015), .B1(n14738), .B2(n14014), .ZN(
        n14019) );
  OAI22_X1 U17349 ( .A1(n14017), .A2(n11114), .B1(n10473), .B2(n14016), .ZN(
        n14018) );
  NOR2_X1 U17350 ( .A1(n14019), .A2(n14018), .ZN(n14021) );
  AOI22_X1 U17351 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n10447), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14020) );
  NAND4_X1 U17352 ( .A1(n14023), .A2(n14022), .A3(n14021), .A4(n14020), .ZN(
        n16178) );
  INV_X1 U17353 ( .A(n14046), .ZN(n14047) );
  AOI22_X1 U17354 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14028) );
  NAND2_X1 U17355 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n14027) );
  NAND2_X1 U17356 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n14026) );
  NAND2_X1 U17357 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n14025) );
  NAND4_X1 U17358 ( .A1(n14028), .A2(n14027), .A3(n14026), .A4(n14025), .ZN(
        n14032) );
  INV_X1 U17359 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14030) );
  INV_X1 U17360 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14029) );
  OAI22_X1 U17361 ( .A1(n14030), .A2(n10464), .B1(n10463), .B2(n14029), .ZN(
        n14031) );
  NOR2_X1 U17362 ( .A1(n14032), .A2(n14031), .ZN(n14045) );
  OR2_X1 U17363 ( .A1(n10467), .A2(n19243), .ZN(n14036) );
  AOI22_X1 U17364 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n14035) );
  NAND2_X1 U17365 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n14034) );
  NAND2_X1 U17366 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14033) );
  AND4_X1 U17367 ( .A1(n14036), .A2(n14035), .A3(n14034), .A4(n14033), .ZN(
        n14044) );
  OAI22_X1 U17368 ( .A1(n10472), .A2(n14038), .B1(n14738), .B2(n14037), .ZN(
        n14042) );
  INV_X1 U17369 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14040) );
  OAI22_X1 U17370 ( .A1(n14040), .A2(n11114), .B1(n10473), .B2(n14039), .ZN(
        n14041) );
  NOR2_X1 U17371 ( .A1(n14042), .A2(n14041), .ZN(n14043) );
  OAI21_X1 U17372 ( .B1(n14047), .B2(n10168), .A(n14704), .ZN(n15091) );
  INV_X1 U17373 ( .A(n14634), .ZN(n14048) );
  AOI21_X1 U17374 ( .B1(n14049), .B2(n15196), .A(n14048), .ZN(n15353) );
  INV_X1 U17375 ( .A(n15353), .ZN(n15183) );
  MUX2_X1 U17376 ( .A(n10887), .B(n15183), .S(n19103), .Z(n14050) );
  OAI21_X1 U17377 ( .B1(n15091), .B2(n19095), .A(n14050), .ZN(P2_U2868) );
  OAI21_X1 U17378 ( .B1(n13982), .B2(n14052), .A(n14051), .ZN(n15873) );
  INV_X1 U17379 ( .A(n14053), .ZN(n14054) );
  OAI21_X1 U17380 ( .B1(n15873), .B2(n14054), .A(n15874), .ZN(n14055) );
  XOR2_X1 U17381 ( .A(n14056), .B(n14055), .Z(n14490) );
  NOR4_X1 U17382 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n15971), .A3(
        n14059), .A4(n13977), .ZN(n14063) );
  NOR2_X1 U17383 ( .A1(n14071), .A2(n14057), .ZN(n14058) );
  OR2_X1 U17384 ( .A1(n14272), .A2(n14058), .ZN(n15788) );
  NOR3_X1 U17385 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15971), .A3(
        n14059), .ZN(n15980) );
  OAI21_X1 U17386 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14517), .A(
        n15994), .ZN(n15981) );
  OAI21_X1 U17387 ( .B1(n15980), .B2(n15981), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14061) );
  INV_X1 U17388 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n15795) );
  OR2_X1 U17389 ( .A1(n15996), .A2(n15795), .ZN(n14060) );
  OAI211_X1 U17390 ( .C1(n20084), .C2(n15788), .A(n14061), .B(n14060), .ZN(
        n14062) );
  NOR2_X1 U17391 ( .A1(n14063), .A2(n14062), .ZN(n14064) );
  OAI21_X1 U17392 ( .B1(n14490), .B2(n16008), .A(n14064), .ZN(P1_U3015) );
  MUX2_X1 U17393 ( .A(DATAI_13_), .B(BUF1_REG_13__SCAN_IN), .S(n20102), .Z(
        n20051) );
  INV_X1 U17394 ( .A(n20051), .ZN(n14066) );
  OAI222_X1 U17395 ( .A1(n14504), .A2(n14370), .B1(n14076), .B2(n14066), .C1(
        n14065), .C2(n14402), .ZN(P1_U2891) );
  INV_X1 U17396 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14067) );
  OAI222_X1 U17397 ( .A1(n15986), .A2(n20005), .B1(n14067), .B2(n20016), .C1(
        n14504), .C2(n14350), .ZN(P1_U2859) );
  INV_X1 U17398 ( .A(n14068), .ZN(n14069) );
  AOI21_X1 U17399 ( .B1(n14070), .B2(n13961), .A(n14069), .ZN(n15879) );
  INV_X1 U17400 ( .A(n15879), .ZN(n14077) );
  AOI21_X1 U17401 ( .B1(n14073), .B2(n14072), .A(n14071), .ZN(n15979) );
  AOI22_X1 U17402 ( .A1(n15979), .A2(n20012), .B1(P1_EBX_REG_15__SCAN_IN), 
        .B2(n14310), .ZN(n14074) );
  OAI21_X1 U17403 ( .B1(n14077), .B2(n14350), .A(n14074), .ZN(P1_U2857) );
  OAI222_X1 U17404 ( .A1(n14077), .A2(n14370), .B1(n14076), .B2(n14075), .C1(
        n14402), .C2(n12265), .ZN(P1_U2889) );
  AOI21_X1 U17405 ( .B1(n18641), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14088) );
  OR2_X1 U17406 ( .A1(n18661), .A2(n14088), .ZN(n18630) );
  NOR2_X1 U17407 ( .A1(n18794), .A2(n18630), .ZN(n14086) );
  NAND2_X1 U17408 ( .A1(n18192), .A2(n9681), .ZN(n18683) );
  INV_X1 U17409 ( .A(n18683), .ZN(n17439) );
  OAI21_X1 U17410 ( .B1(n14079), .B2(n17439), .A(n18839), .ZN(n17377) );
  INV_X1 U17411 ( .A(n18834), .ZN(n18841) );
  OR2_X1 U17412 ( .A1(n18623), .A2(n18841), .ZN(n14084) );
  INV_X1 U17413 ( .A(n9681), .ZN(n14080) );
  AOI221_X2 U17414 ( .B1(n18192), .B2(n18661), .C1(n14080), .C2(n18661), .A(
        n14084), .ZN(n15713) );
  NOR2_X1 U17415 ( .A1(n18620), .A2(n15474), .ZN(n14081) );
  NOR2_X1 U17416 ( .A1(n15713), .A2(n14081), .ZN(n14082) );
  OAI211_X1 U17417 ( .C1(n17377), .C2(n14084), .A(n14083), .B(n14082), .ZN(
        n18667) );
  NOR2_X1 U17418 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18790), .ZN(n18187) );
  INV_X1 U17419 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18178) );
  NAND3_X1 U17420 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18788)
         );
  NOR2_X1 U17421 ( .A1(n18178), .A2(n18788), .ZN(n14085) );
  MUX2_X1 U17422 ( .A(n14086), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18821), .Z(P3_U3284) );
  NAND2_X1 U17423 ( .A1(n14088), .A2(n14087), .ZN(n18177) );
  NOR2_X1 U17424 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18177), .ZN(n14089) );
  INV_X1 U17425 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18843) );
  NOR2_X1 U17426 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18846) );
  AOI21_X1 U17427 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n18846), .ZN(n18699) );
  OR2_X1 U17428 ( .A1(n18815), .A2(n18699), .ZN(n18186) );
  OAI21_X1 U17429 ( .B1(n14089), .B2(n18788), .A(n18288), .ZN(n18183) );
  INV_X1 U17430 ( .A(n18183), .ZN(n14090) );
  NAND2_X1 U17431 ( .A1(n18851), .A2(n18790), .ZN(n16519) );
  AND2_X1 U17432 ( .A1(n18794), .A2(n16519), .ZN(n18837) );
  INV_X1 U17433 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n16542) );
  NOR2_X1 U17434 ( .A1(n18800), .A2(n16542), .ZN(n17810) );
  NOR2_X1 U17435 ( .A1(n18837), .A2(n17810), .ZN(n15572) );
  AOI21_X1 U17436 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15572), .ZN(n15573) );
  NOR2_X1 U17437 ( .A1(n14090), .A2(n15573), .ZN(n14092) );
  NAND3_X1 U17438 ( .A1(n18851), .A2(n18790), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18334) );
  INV_X1 U17439 ( .A(n18334), .ZN(n18524) );
  NOR2_X1 U17440 ( .A1(n18790), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18223) );
  OR2_X1 U17441 ( .A1(n18223), .A2(n14090), .ZN(n15571) );
  OR2_X1 U17442 ( .A1(n18524), .A2(n15571), .ZN(n14091) );
  MUX2_X1 U17443 ( .A(n14092), .B(n14091), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NOR2_X1 U17444 ( .A1(n14096), .A2(n20100), .ZN(n14095) );
  NAND2_X1 U17445 ( .A1(n14402), .A2(n14095), .ZN(n14404) );
  AOI22_X1 U17446 ( .A1(n14398), .A2(BUF1_REG_28__SCAN_IN), .B1(
        P1_EAX_REG_28__SCAN_IN), .B2(n14397), .ZN(n14098) );
  NOR3_X4 U17447 ( .A1(n14397), .A2(n14208), .A3(n11877), .ZN(n14407) );
  NOR3_X4 U17448 ( .A1(n14397), .A2(n20102), .A3(n14096), .ZN(n14406) );
  AOI22_X1 U17449 ( .A1(n14407), .A2(n20049), .B1(n14406), .B2(DATAI_28_), 
        .ZN(n14097) );
  OAI211_X1 U17450 ( .C1(n14431), .C2(n14370), .A(n14098), .B(n14097), .ZN(
        P1_U2876) );
  INV_X1 U17451 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14100) );
  OAI21_X1 U17452 ( .B1(n14241), .B2(n14099), .A(n9695), .ZN(n14567) );
  INV_X1 U17453 ( .A(n14567), .ZN(n14110) );
  NOR2_X1 U17454 ( .A1(n19961), .A2(n19960), .ZN(n14299) );
  INV_X1 U17455 ( .A(n14299), .ZN(n15750) );
  NAND2_X1 U17456 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n14227) );
  INV_X1 U17457 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20849) );
  NAND2_X1 U17458 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n14101), .ZN(n14279) );
  NOR2_X1 U17459 ( .A1(n13940), .A2(n14279), .ZN(n14262) );
  INV_X1 U17460 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14270) );
  INV_X1 U17461 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n15803) );
  NOR3_X1 U17462 ( .A1(n14270), .A2(n15795), .A3(n15803), .ZN(n14261) );
  NAND2_X1 U17463 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n14261), .ZN(n15766) );
  INV_X1 U17464 ( .A(n15766), .ZN(n14102) );
  NAND4_X1 U17465 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_19__SCAN_IN), 
        .A3(n14262), .A4(n14102), .ZN(n15756) );
  NOR2_X1 U17466 ( .A1(n20849), .A2(n15756), .ZN(n15738) );
  NAND3_X1 U17467 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(n15738), .ZN(n15727) );
  INV_X1 U17468 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20853) );
  NOR2_X1 U17469 ( .A1(n15727), .A2(n20853), .ZN(n15718) );
  AND2_X1 U17470 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14103) );
  NAND2_X1 U17471 ( .A1(n15718), .A2(n14103), .ZN(n14173) );
  INV_X1 U17472 ( .A(n14173), .ZN(n14104) );
  AOI21_X1 U17473 ( .B1(n14104), .B2(n19976), .A(n14299), .ZN(n14249) );
  AOI21_X1 U17474 ( .B1(n15750), .B2(n14227), .A(n14249), .ZN(n14231) );
  NAND2_X1 U17475 ( .A1(n19961), .A2(n14104), .ZN(n14238) );
  INV_X1 U17476 ( .A(n14238), .ZN(n14105) );
  AOI21_X1 U17477 ( .B1(n14105), .B2(P1_REIP_REG_27__SCAN_IN), .A(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14108) );
  AOI22_X1 U17478 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19978), .B1(
        n19979), .B2(n14434), .ZN(n14107) );
  NAND2_X1 U17479 ( .A1(n19932), .A2(P1_EBX_REG_28__SCAN_IN), .ZN(n14106) );
  OAI211_X1 U17480 ( .C1(n14231), .C2(n14108), .A(n14107), .B(n14106), .ZN(
        n14109) );
  AOI21_X1 U17481 ( .B1(n14110), .B2(n19940), .A(n14109), .ZN(n14111) );
  OAI21_X1 U17482 ( .B1(n14431), .B2(n19923), .A(n14111), .ZN(P1_U2812) );
  NAND2_X1 U17483 ( .A1(n14112), .A2(n20074), .ZN(n14118) );
  INV_X1 U17484 ( .A(n14113), .ZN(n19972) );
  OAI21_X1 U17485 ( .B1(n15918), .B2(n14115), .A(n14114), .ZN(n14116) );
  AOI21_X1 U17486 ( .B1(n19972), .B2(n15889), .A(n14116), .ZN(n14117) );
  OAI211_X1 U17487 ( .C1(n20101), .C2(n19971), .A(n14118), .B(n14117), .ZN(
        P1_U2996) );
  AOI22_X1 U17488 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n13376), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n14119) );
  OAI21_X1 U17489 ( .B1(n15914), .B2(n19977), .A(n14119), .ZN(n14120) );
  AOI21_X1 U17490 ( .B1(n15909), .B2(n19990), .A(n14120), .ZN(n14121) );
  OAI21_X1 U17491 ( .B1(n19877), .B2(n14122), .A(n14121), .ZN(P1_U2997) );
  INV_X1 U17492 ( .A(n19984), .ZN(n14123) );
  AOI22_X1 U17493 ( .A1(n20012), .A2(n14123), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n14310), .ZN(n14124) );
  OAI21_X1 U17494 ( .B1(n14125), .B2(n14350), .A(n14124), .ZN(P1_U2870) );
  NAND2_X1 U17495 ( .A1(n20225), .A2(n14597), .ZN(n14128) );
  NAND2_X1 U17496 ( .A1(n14126), .A2(n14130), .ZN(n14127) );
  NAND2_X1 U17497 ( .A1(n14128), .A2(n14127), .ZN(n15631) );
  OAI22_X1 U17498 ( .A1(n21068), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14614), .ZN(n14129) );
  AOI21_X1 U17499 ( .B1(n15631), .B2(n16071), .A(n14129), .ZN(n14132) );
  OAI22_X1 U17500 ( .A1(n15634), .A2(n19871), .B1(n16083), .B2(n19878), .ZN(
        n16072) );
  AOI21_X1 U17501 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20804), .A(n16072), 
        .ZN(n14603) );
  AOI21_X1 U17502 ( .B1(n15628), .B2(n16071), .A(n14603), .ZN(n14131) );
  OAI22_X1 U17503 ( .A1(n14132), .A2(n14603), .B1(n14131), .B2(n14130), .ZN(
        P1_U3474) );
  NOR4_X1 U17504 ( .A1(n15255), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14134), .A4(n14133), .ZN(n14140) );
  NAND3_X1 U17505 ( .A1(n14135), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n15426), .ZN(n14138) );
  INV_X1 U17506 ( .A(n14136), .ZN(n14137) );
  NAND2_X1 U17507 ( .A1(n14138), .A2(n14137), .ZN(n14139) );
  NAND2_X1 U17508 ( .A1(n14142), .A2(n16314), .ZN(n14143) );
  OAI211_X1 U17509 ( .C1(n14145), .C2(n16326), .A(n14144), .B(n14143), .ZN(
        P2_U3015) );
  AND3_X1 U17510 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14533) );
  INV_X1 U17511 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15682) );
  INV_X1 U17512 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15674) );
  NAND3_X1 U17513 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14534) );
  INV_X1 U17514 ( .A(n14534), .ZN(n14148) );
  NOR2_X1 U17515 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14150) );
  NAND2_X1 U17516 ( .A1(n14150), .A2(n14149), .ZN(n14424) );
  OR2_X1 U17517 ( .A1(n13705), .A2(n14424), .ZN(n14151) );
  OAI21_X1 U17518 ( .B1(n15832), .B2(n14424), .A(n9834), .ZN(n14153) );
  NAND2_X1 U17519 ( .A1(n14572), .A2(n14153), .ZN(n14154) );
  AND2_X1 U17520 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14561) );
  NOR2_X1 U17521 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14563) );
  INV_X1 U17522 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14545) );
  XNOR2_X1 U17523 ( .A(n14470), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14418) );
  OAI21_X1 U17524 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n14545), .A(
        n14418), .ZN(n14155) );
  AOI22_X1 U17525 ( .A1(n14159), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n14158), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14160) );
  INV_X1 U17526 ( .A(n14160), .ZN(n14161) );
  INV_X1 U17527 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n21089) );
  NAND2_X1 U17528 ( .A1(n15889), .A2(n14163), .ZN(n14164) );
  NAND2_X1 U17529 ( .A1(n13376), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14531) );
  OAI211_X1 U17530 ( .C1(n15918), .C2(n21089), .A(n14164), .B(n14531), .ZN(
        n14165) );
  OAI21_X1 U17531 ( .B1(n19877), .B2(n14541), .A(n14166), .ZN(P1_U2968) );
  AOI22_X1 U17532 ( .A1(n14168), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14167), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14171) );
  MUX2_X1 U17533 ( .A(n9648), .B(n14169), .S(n14224), .Z(n14170) );
  XOR2_X1 U17534 ( .A(n14171), .B(n14170), .Z(n14530) );
  NAND2_X1 U17535 ( .A1(n14209), .A2(n19916), .ZN(n14179) );
  INV_X1 U17536 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14175) );
  NAND3_X1 U17537 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .A3(P1_REIP_REG_27__SCAN_IN), .ZN(n14172) );
  OR2_X1 U17538 ( .A1(n14173), .A2(n14172), .ZN(n14213) );
  NOR3_X1 U17539 ( .A1(n19960), .A2(n14175), .A3(n14213), .ZN(n14174) );
  NOR2_X1 U17540 ( .A1(n14299), .A2(n14174), .ZN(n14214) );
  NOR4_X1 U17541 ( .A1(n19965), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14175), 
        .A4(n14213), .ZN(n14177) );
  INV_X1 U17542 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14300) );
  OAI22_X1 U17543 ( .A1(n19987), .A2(n14300), .B1(n21089), .B2(n19898), .ZN(
        n14176) );
  AOI211_X1 U17544 ( .C1(n14214), .C2(P1_REIP_REG_31__SCAN_IN), .A(n14177), 
        .B(n14176), .ZN(n14178) );
  OAI211_X1 U17545 ( .C1(n14530), .C2(n19985), .A(n14179), .B(n14178), .ZN(
        P1_U2809) );
  NAND2_X1 U17546 ( .A1(n19217), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n14199) );
  AOI21_X1 U17547 ( .B1(n14182), .B2(n14181), .A(n14180), .ZN(n14203) );
  NAND2_X1 U17548 ( .A1(n16314), .A2(n14203), .ZN(n14186) );
  NAND2_X1 U17549 ( .A1(n14184), .A2(n14183), .ZN(n14204) );
  NAND3_X1 U17550 ( .A1(n16317), .A2(n14205), .A3(n14204), .ZN(n14185) );
  NAND4_X1 U17551 ( .A1(n14187), .A2(n14199), .A3(n14186), .A4(n14185), .ZN(
        n14188) );
  AOI21_X1 U17552 ( .B1(n19835), .B2(n16312), .A(n14188), .ZN(n14198) );
  INV_X1 U17553 ( .A(n15598), .ZN(n14190) );
  NAND2_X1 U17554 ( .A1(n14190), .A2(n14189), .ZN(n14196) );
  NAND2_X1 U17555 ( .A1(n14190), .A2(n14193), .ZN(n14191) );
  OAI211_X1 U17556 ( .C1(n14193), .C2(n14192), .A(n14191), .B(n16331), .ZN(
        n14194) );
  INV_X1 U17557 ( .A(n14194), .ZN(n14195) );
  MUX2_X1 U17558 ( .A(n14196), .B(n14195), .S(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n14197) );
  OAI211_X1 U17559 ( .C1(n10357), .C2(n16327), .A(n14198), .B(n14197), .ZN(
        P2_U3044) );
  INV_X1 U17560 ( .A(n14664), .ZN(n14665) );
  NAND2_X1 U17561 ( .A1(n16268), .A2(n14665), .ZN(n14200) );
  OAI211_X1 U17562 ( .C1(n16278), .C2(n14201), .A(n14200), .B(n14199), .ZN(
        n14202) );
  AOI21_X1 U17563 ( .B1(n16269), .B2(n14203), .A(n14202), .ZN(n14207) );
  NAND3_X1 U17564 ( .A1(n14205), .A2(n11389), .A3(n14204), .ZN(n14206) );
  OAI211_X1 U17565 ( .C1(n10380), .C2(n16273), .A(n14207), .B(n14206), .ZN(
        P2_U3012) );
  INV_X1 U17566 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16425) );
  AND2_X1 U17567 ( .A1(n14402), .A2(n14208), .ZN(n14210) );
  NAND2_X1 U17568 ( .A1(n14210), .A2(n14209), .ZN(n14212) );
  AOI22_X1 U17569 ( .A1(n14406), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14397), .ZN(n14211) );
  OAI211_X1 U17570 ( .C1(n14404), .C2(n16425), .A(n14212), .B(n14211), .ZN(
        P1_U2873) );
  NOR2_X1 U17571 ( .A1(n19965), .A2(n14213), .ZN(n14215) );
  OAI21_X1 U17572 ( .B1(P1_REIP_REG_30__SCAN_IN), .B2(n14215), .A(n14214), 
        .ZN(n14217) );
  AOI22_X1 U17573 ( .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19978), .B1(
        n19979), .B2(n14411), .ZN(n14216) );
  OAI211_X1 U17574 ( .C1(n19987), .C2(n14218), .A(n14217), .B(n14216), .ZN(
        n14219) );
  AOI21_X1 U17575 ( .B1(n14548), .B2(n19940), .A(n14219), .ZN(n14220) );
  OAI21_X1 U17576 ( .B1(n14355), .B2(n19923), .A(n14220), .ZN(P1_U2810) );
  AOI21_X1 U17577 ( .B1(n14223), .B2(n14222), .A(n14221), .ZN(n14422) );
  INV_X1 U17578 ( .A(n14422), .ZN(n14358) );
  AOI21_X1 U17579 ( .B1(n14225), .B2(n9695), .A(n14224), .ZN(n14552) );
  INV_X1 U17580 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20862) );
  OAI22_X1 U17581 ( .A1(n14226), .A2(n19898), .B1(n19935), .B2(n14420), .ZN(
        n14229) );
  NOR3_X1 U17582 ( .A1(n14238), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n14227), 
        .ZN(n14228) );
  AOI211_X1 U17583 ( .C1(P1_EBX_REG_29__SCAN_IN), .C2(n19932), .A(n14229), .B(
        n14228), .ZN(n14230) );
  OAI21_X1 U17584 ( .B1(n14231), .B2(n20862), .A(n14230), .ZN(n14232) );
  AOI21_X1 U17585 ( .B1(n14552), .B2(n19940), .A(n14232), .ZN(n14233) );
  OAI21_X1 U17586 ( .B1(n14358), .B2(n19923), .A(n14233), .ZN(P1_U2811) );
  INV_X1 U17587 ( .A(n14234), .ZN(n14245) );
  AOI21_X1 U17588 ( .B1(n14235), .B2(n14245), .A(n14093), .ZN(n14442) );
  INV_X1 U17589 ( .A(n14442), .ZN(n14362) );
  AOI22_X1 U17590 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19978), .B1(
        n19979), .B2(n14438), .ZN(n14237) );
  NAND2_X1 U17591 ( .A1(n19932), .A2(P1_EBX_REG_27__SCAN_IN), .ZN(n14236) );
  OAI211_X1 U17592 ( .C1(n14238), .C2(P1_REIP_REG_27__SCAN_IN), .A(n14237), 
        .B(n14236), .ZN(n14243) );
  NOR2_X1 U17593 ( .A1(n14246), .A2(n14239), .ZN(n14240) );
  OR2_X1 U17594 ( .A1(n14241), .A2(n14240), .ZN(n15921) );
  NOR2_X1 U17595 ( .A1(n15921), .A2(n19985), .ZN(n14242) );
  AOI211_X1 U17596 ( .C1(n14249), .C2(P1_REIP_REG_27__SCAN_IN), .A(n14243), 
        .B(n14242), .ZN(n14244) );
  OAI21_X1 U17597 ( .B1(n14362), .B2(n19923), .A(n14244), .ZN(P1_U2813) );
  OAI21_X1 U17598 ( .B1(n9721), .B2(n9788), .A(n14245), .ZN(n14452) );
  AOI21_X1 U17599 ( .B1(n14247), .B2(n14309), .A(n14246), .ZN(n14576) );
  NAND2_X1 U17600 ( .A1(n15718), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14248) );
  NOR2_X1 U17601 ( .A1(n19965), .A2(n14248), .ZN(n14250) );
  OAI21_X1 U17602 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(n14250), .A(n14249), 
        .ZN(n14252) );
  AOI22_X1 U17603 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19978), .B1(
        n19979), .B2(n14446), .ZN(n14251) );
  OAI211_X1 U17604 ( .C1(n19987), .C2(n14304), .A(n14252), .B(n14251), .ZN(
        n14253) );
  AOI21_X1 U17605 ( .B1(n14576), .B2(n19940), .A(n14253), .ZN(n14254) );
  OAI21_X1 U17606 ( .B1(n14452), .B2(n19923), .A(n14254), .ZN(P1_U2814) );
  OAI21_X1 U17607 ( .B1(n10076), .B2(n9797), .A(n14256), .ZN(n14484) );
  OAI21_X1 U17608 ( .B1(n19965), .B2(n14262), .A(n19976), .ZN(n14288) );
  INV_X1 U17609 ( .A(n14288), .ZN(n15802) );
  OAI21_X1 U17610 ( .B1(n14299), .B2(n14261), .A(n15802), .ZN(n15779) );
  NOR2_X1 U17611 ( .A1(n19898), .A2(n14478), .ZN(n14257) );
  AOI211_X1 U17612 ( .C1(n19979), .C2(n14480), .A(n19946), .B(n14257), .ZN(
        n14259) );
  NAND2_X1 U17613 ( .A1(n19932), .A2(P1_EBX_REG_18__SCAN_IN), .ZN(n14258) );
  OAI211_X1 U17614 ( .C1(n14260), .C2(n19985), .A(n14259), .B(n14258), .ZN(
        n14264) );
  INV_X1 U17615 ( .A(n14261), .ZN(n14263) );
  NAND2_X1 U17616 ( .A1(n19961), .A2(n14262), .ZN(n15798) );
  NOR3_X1 U17617 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n14263), .A3(n15798), 
        .ZN(n15780) );
  AOI211_X1 U17618 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n15779), .A(n14264), 
        .B(n15780), .ZN(n14265) );
  OAI21_X1 U17619 ( .B1(n14484), .B2(n19923), .A(n14265), .ZN(P1_U2822) );
  INV_X1 U17620 ( .A(n14266), .ZN(n14269) );
  INV_X1 U17621 ( .A(n14267), .ZN(n14268) );
  AOI21_X1 U17622 ( .B1(n14269), .B2(n14268), .A(n10076), .ZN(n15868) );
  INV_X1 U17623 ( .A(n15868), .ZN(n14401) );
  NAND2_X1 U17624 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15784) );
  OAI21_X1 U17625 ( .B1(n15784), .B2(n15798), .A(n14270), .ZN(n14277) );
  OAI21_X1 U17626 ( .B1(n14272), .B2(n14271), .A(n9764), .ZN(n15972) );
  NOR2_X1 U17627 ( .A1(n19898), .A2(n12305), .ZN(n14273) );
  AOI211_X1 U17628 ( .C1(n19979), .C2(n15867), .A(n19946), .B(n14273), .ZN(
        n14275) );
  NAND2_X1 U17629 ( .A1(n19932), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n14274) );
  OAI211_X1 U17630 ( .C1(n15972), .C2(n19985), .A(n14275), .B(n14274), .ZN(
        n14276) );
  AOI21_X1 U17631 ( .B1(n15779), .B2(n14277), .A(n14276), .ZN(n14278) );
  OAI21_X1 U17632 ( .B1(n14401), .B2(n19923), .A(n14278), .ZN(P1_U2823) );
  OAI21_X1 U17633 ( .B1(n19965), .B2(n14279), .A(n13940), .ZN(n14287) );
  NOR2_X1 U17634 ( .A1(n19935), .A2(n14280), .ZN(n14281) );
  AOI211_X1 U17635 ( .C1(n19978), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n19946), .B(n14281), .ZN(n14284) );
  NAND2_X1 U17636 ( .A1(n19940), .A2(n14282), .ZN(n14283) );
  OAI211_X1 U17637 ( .C1(n14285), .C2(n19987), .A(n14284), .B(n14283), .ZN(
        n14286) );
  AOI21_X1 U17638 ( .B1(n14288), .B2(n14287), .A(n14286), .ZN(n14289) );
  OAI21_X1 U17639 ( .B1(n14290), .B2(n19923), .A(n14289), .ZN(P1_U2826) );
  INV_X1 U17640 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n14298) );
  INV_X1 U17641 ( .A(n20079), .ZN(n14296) );
  OAI21_X1 U17642 ( .B1(n19978), .B2(n19979), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14291) );
  OAI21_X1 U17643 ( .B1(n19981), .B2(n14292), .A(n14291), .ZN(n14295) );
  OAI22_X1 U17644 ( .A1(n14293), .A2(n19987), .B1(n19985), .B2(n20083), .ZN(
        n14294) );
  AOI211_X1 U17645 ( .C1(n14296), .C2(n19991), .A(n14295), .B(n14294), .ZN(
        n14297) );
  OAI21_X1 U17646 ( .B1(n14299), .B2(n14298), .A(n14297), .ZN(P1_U2840) );
  OAI22_X1 U17647 ( .A1(n14530), .A2(n20005), .B1(n20016), .B2(n14300), .ZN(
        P1_U2841) );
  AOI22_X1 U17648 ( .A1(n14552), .A2(n20012), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14310), .ZN(n14301) );
  OAI21_X1 U17649 ( .B1(n14358), .B2(n14350), .A(n14301), .ZN(P1_U2843) );
  INV_X1 U17650 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14302) );
  OAI222_X1 U17651 ( .A1(n14350), .A2(n14362), .B1(n14302), .B2(n20016), .C1(
        n15921), .C2(n20005), .ZN(P1_U2845) );
  INV_X1 U17652 ( .A(n14576), .ZN(n14303) );
  OAI222_X1 U17653 ( .A1(n14452), .A2(n14350), .B1(n14304), .B2(n20016), .C1(
        n14303), .C2(n20005), .ZN(P1_U2846) );
  INV_X1 U17654 ( .A(n14305), .ZN(n14306) );
  AOI21_X1 U17655 ( .B1(n14306), .B2(n9691), .A(n9721), .ZN(n15827) );
  INV_X1 U17656 ( .A(n15827), .ZN(n14367) );
  NAND2_X1 U17657 ( .A1(n9715), .A2(n14307), .ZN(n14308) );
  AND2_X1 U17658 ( .A1(n14309), .A2(n14308), .ZN(n15937) );
  AOI22_X1 U17659 ( .A1(n15937), .A2(n20012), .B1(P1_EBX_REG_25__SCAN_IN), 
        .B2(n14310), .ZN(n14311) );
  OAI21_X1 U17660 ( .B1(n14367), .B2(n14350), .A(n14311), .ZN(P1_U2847) );
  OAI21_X1 U17661 ( .B1(n14313), .B2(n14312), .A(n9691), .ZN(n15731) );
  OR2_X1 U17662 ( .A1(n14323), .A2(n14314), .ZN(n14315) );
  NAND2_X1 U17663 ( .A1(n9715), .A2(n14315), .ZN(n15730) );
  OAI22_X1 U17664 ( .A1(n15730), .A2(n20005), .B1(n15729), .B2(n20016), .ZN(
        n14316) );
  INV_X1 U17665 ( .A(n14316), .ZN(n14317) );
  OAI21_X1 U17666 ( .B1(n15731), .B2(n14350), .A(n14317), .ZN(P1_U2848) );
  AND2_X1 U17667 ( .A1(n14318), .A2(n14319), .ZN(n14320) );
  OR2_X1 U17668 ( .A1(n14320), .A2(n14312), .ZN(n15839) );
  INV_X1 U17669 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14324) );
  NOR2_X1 U17670 ( .A1(n14330), .A2(n14321), .ZN(n14322) );
  OR2_X1 U17671 ( .A1(n14323), .A2(n14322), .ZN(n15945) );
  OAI222_X1 U17672 ( .A1(n15839), .A2(n14350), .B1(n14324), .B2(n20016), .C1(
        n15945), .C2(n20005), .ZN(P1_U2849) );
  NAND2_X1 U17673 ( .A1(n14325), .A2(n14326), .ZN(n14327) );
  AND2_X1 U17674 ( .A1(n14318), .A2(n14327), .ZN(n15749) );
  INV_X1 U17675 ( .A(n15749), .ZN(n14376) );
  NOR2_X1 U17676 ( .A1(n15679), .A2(n14328), .ZN(n14329) );
  OR2_X1 U17677 ( .A1(n14330), .A2(n14329), .ZN(n15953) );
  OAI22_X1 U17678 ( .A1(n15953), .A2(n20005), .B1(n14331), .B2(n20016), .ZN(
        n14332) );
  INV_X1 U17679 ( .A(n14332), .ZN(n14333) );
  OAI21_X1 U17680 ( .B1(n14376), .B2(n14350), .A(n14333), .ZN(P1_U2850) );
  NOR2_X1 U17681 ( .A1(n9693), .A2(n14335), .ZN(n14336) );
  OR2_X1 U17682 ( .A1(n14334), .A2(n14336), .ZN(n15765) );
  INV_X1 U17683 ( .A(n15677), .ZN(n14337) );
  XNOR2_X1 U17684 ( .A(n15675), .B(n14337), .ZN(n15767) );
  OAI222_X1 U17685 ( .A1(n15765), .A2(n14350), .B1(n14338), .B2(n20016), .C1(
        n20005), .C2(n15767), .ZN(P1_U2852) );
  AND2_X1 U17686 ( .A1(n14256), .A2(n14339), .ZN(n14340) );
  NOR2_X1 U17687 ( .A1(n9693), .A2(n14340), .ZN(n15857) );
  INV_X1 U17688 ( .A(n15857), .ZN(n14391) );
  INV_X1 U17689 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14343) );
  NAND2_X1 U17690 ( .A1(n9716), .A2(n14341), .ZN(n14342) );
  NAND2_X1 U17691 ( .A1(n15675), .A2(n14342), .ZN(n15961) );
  OAI222_X1 U17692 ( .A1(n14391), .A2(n14350), .B1(n14343), .B2(n20016), .C1(
        n15961), .C2(n20005), .ZN(P1_U2853) );
  NOR2_X1 U17693 ( .A1(n20016), .A2(n14344), .ZN(n14345) );
  AOI21_X1 U17694 ( .B1(n14346), .B2(n20012), .A(n14345), .ZN(n14347) );
  OAI21_X1 U17695 ( .B1(n14484), .B2(n14350), .A(n14347), .ZN(P1_U2854) );
  INV_X1 U17696 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14348) );
  OAI222_X1 U17697 ( .A1(n15972), .A2(n20005), .B1(n14348), .B2(n20016), .C1(
        n14401), .C2(n14350), .ZN(P1_U2855) );
  AOI21_X1 U17698 ( .B1(n14349), .B2(n14068), .A(n14267), .ZN(n14488) );
  OAI22_X1 U17699 ( .A1(n15788), .A2(n20005), .B1(n15787), .B2(n20016), .ZN(
        n14351) );
  AOI21_X1 U17700 ( .B1(n14488), .B2(n12640), .A(n14351), .ZN(n14352) );
  INV_X1 U17701 ( .A(n14352), .ZN(P1_U2856) );
  AOI22_X1 U17702 ( .A1(n14398), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14397), .ZN(n14354) );
  AOI22_X1 U17703 ( .A1(n14407), .A2(n20053), .B1(n14406), .B2(DATAI_30_), 
        .ZN(n14353) );
  OAI211_X1 U17704 ( .C1(n14355), .C2(n14370), .A(n14354), .B(n14353), .ZN(
        P1_U2874) );
  AOI22_X1 U17705 ( .A1(n14398), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14397), .ZN(n14357) );
  AOI22_X1 U17706 ( .A1(n14407), .A2(n20051), .B1(n14406), .B2(DATAI_29_), 
        .ZN(n14356) );
  OAI211_X1 U17707 ( .C1(n14358), .C2(n14370), .A(n14357), .B(n14356), .ZN(
        P1_U2875) );
  AOI22_X1 U17708 ( .A1(n14398), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14397), .ZN(n14361) );
  AOI22_X1 U17709 ( .A1(n14407), .A2(n14359), .B1(n14406), .B2(DATAI_27_), 
        .ZN(n14360) );
  OAI211_X1 U17710 ( .C1(n14362), .C2(n14370), .A(n14361), .B(n14360), .ZN(
        P1_U2877) );
  AOI22_X1 U17711 ( .A1(n14398), .A2(BUF1_REG_26__SCAN_IN), .B1(
        P1_EAX_REG_26__SCAN_IN), .B2(n14397), .ZN(n14364) );
  AOI22_X1 U17712 ( .A1(n14407), .A2(n20047), .B1(n14406), .B2(DATAI_26_), 
        .ZN(n14363) );
  OAI211_X1 U17713 ( .C1(n14452), .C2(n14370), .A(n14364), .B(n14363), .ZN(
        P1_U2878) );
  AOI22_X1 U17714 ( .A1(n14398), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14397), .ZN(n14366) );
  AOI22_X1 U17715 ( .A1(n14407), .A2(n20045), .B1(n14406), .B2(DATAI_25_), 
        .ZN(n14365) );
  OAI211_X1 U17716 ( .C1(n14367), .C2(n14370), .A(n14366), .B(n14365), .ZN(
        P1_U2879) );
  AOI22_X1 U17717 ( .A1(n14398), .A2(BUF1_REG_24__SCAN_IN), .B1(
        P1_EAX_REG_24__SCAN_IN), .B2(n14397), .ZN(n14369) );
  AOI22_X1 U17718 ( .A1(n14407), .A2(n20043), .B1(n14406), .B2(DATAI_24_), 
        .ZN(n14368) );
  OAI211_X1 U17719 ( .C1(n15731), .C2(n14370), .A(n14369), .B(n14368), .ZN(
        P1_U2880) );
  AOI22_X1 U17720 ( .A1(n14398), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n14397), .ZN(n14373) );
  AOI22_X1 U17721 ( .A1(n14407), .A2(n14371), .B1(n14406), .B2(DATAI_23_), 
        .ZN(n14372) );
  OAI211_X1 U17722 ( .C1(n15839), .C2(n14370), .A(n14373), .B(n14372), .ZN(
        P1_U2881) );
  AOI22_X1 U17723 ( .A1(n14398), .A2(BUF1_REG_22__SCAN_IN), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(n14397), .ZN(n14375) );
  AOI22_X1 U17724 ( .A1(n14407), .A2(n20138), .B1(n14406), .B2(DATAI_22_), 
        .ZN(n14374) );
  OAI211_X1 U17725 ( .C1(n14376), .C2(n14370), .A(n14375), .B(n14374), .ZN(
        P1_U2882) );
  OR2_X1 U17726 ( .A1(n14334), .A2(n14377), .ZN(n14378) );
  AND2_X1 U17727 ( .A1(n14325), .A2(n14378), .ZN(n15846) );
  INV_X1 U17728 ( .A(n15846), .ZN(n14383) );
  INV_X1 U17729 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16444) );
  OAI22_X1 U17730 ( .A1(n14404), .A2(n16444), .B1(n14379), .B2(n14402), .ZN(
        n14380) );
  INV_X1 U17731 ( .A(n14380), .ZN(n14382) );
  AOI22_X1 U17732 ( .A1(n14407), .A2(n20133), .B1(n14406), .B2(DATAI_21_), 
        .ZN(n14381) );
  OAI211_X1 U17733 ( .C1(n14383), .C2(n14370), .A(n14382), .B(n14381), .ZN(
        P1_U2883) );
  INV_X1 U17734 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n14385) );
  OAI22_X1 U17735 ( .A1(n14404), .A2(n14385), .B1(n14384), .B2(n14402), .ZN(
        n14386) );
  INV_X1 U17736 ( .A(n14386), .ZN(n14388) );
  AOI22_X1 U17737 ( .A1(n14407), .A2(n20129), .B1(n14406), .B2(DATAI_20_), 
        .ZN(n14387) );
  OAI211_X1 U17738 ( .C1(n15765), .C2(n14370), .A(n14388), .B(n14387), .ZN(
        P1_U2884) );
  AOI22_X1 U17739 ( .A1(n14398), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14397), .ZN(n14390) );
  AOI22_X1 U17740 ( .A1(n14407), .A2(n20123), .B1(n14406), .B2(DATAI_19_), 
        .ZN(n14389) );
  OAI211_X1 U17741 ( .C1(n14391), .C2(n14370), .A(n14390), .B(n14389), .ZN(
        P1_U2885) );
  INV_X1 U17742 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n14393) );
  INV_X1 U17743 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14392) );
  OAI22_X1 U17744 ( .A1(n14404), .A2(n14393), .B1(n14392), .B2(n14402), .ZN(
        n14394) );
  INV_X1 U17745 ( .A(n14394), .ZN(n14396) );
  AOI22_X1 U17746 ( .A1(n14407), .A2(n20118), .B1(n14406), .B2(DATAI_18_), 
        .ZN(n14395) );
  OAI211_X1 U17747 ( .C1(n14484), .C2(n14370), .A(n14396), .B(n14395), .ZN(
        P1_U2886) );
  AOI22_X1 U17748 ( .A1(n14398), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14397), .ZN(n14400) );
  AOI22_X1 U17749 ( .A1(n14407), .A2(n20113), .B1(n14406), .B2(DATAI_17_), 
        .ZN(n14399) );
  OAI211_X1 U17750 ( .C1(n14401), .C2(n14370), .A(n14400), .B(n14399), .ZN(
        P1_U2887) );
  INV_X1 U17751 ( .A(n14488), .ZN(n15789) );
  INV_X1 U17752 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n14403) );
  OAI22_X1 U17753 ( .A1(n14404), .A2(n14403), .B1(n13040), .B2(n14402), .ZN(
        n14405) );
  INV_X1 U17754 ( .A(n14405), .ZN(n14409) );
  AOI22_X1 U17755 ( .A1(n14407), .A2(n20099), .B1(n14406), .B2(DATAI_16_), 
        .ZN(n14408) );
  OAI211_X1 U17756 ( .C1(n15789), .C2(n14370), .A(n14409), .B(n14408), .ZN(
        P1_U2888) );
  NAND2_X1 U17757 ( .A1(n15889), .A2(n14411), .ZN(n14412) );
  NAND2_X1 U17758 ( .A1(n13376), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14542) );
  OAI211_X1 U17759 ( .C1(n14413), .C2(n15918), .A(n14412), .B(n14542), .ZN(
        n14414) );
  AOI21_X1 U17760 ( .B1(n14415), .B2(n15909), .A(n14414), .ZN(n14416) );
  OAI21_X1 U17761 ( .B1(n14550), .B2(n19877), .A(n14416), .ZN(P1_U2969) );
  XOR2_X1 U17762 ( .A(n14418), .B(n14417), .Z(n14560) );
  NOR2_X1 U17763 ( .A1(n15996), .A2(n20862), .ZN(n14551) );
  AOI21_X1 U17764 ( .B1(n20076), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14551), .ZN(n14419) );
  OAI21_X1 U17765 ( .B1(n15914), .B2(n14420), .A(n14419), .ZN(n14421) );
  AOI21_X1 U17766 ( .B1(n14422), .B2(n15909), .A(n14421), .ZN(n14423) );
  OAI21_X1 U17767 ( .B1(n19877), .B2(n14560), .A(n14423), .ZN(P1_U2970) );
  INV_X1 U17768 ( .A(n14424), .ZN(n14425) );
  AOI21_X1 U17769 ( .B1(n14425), .B2(n14448), .A(n14427), .ZN(n14426) );
  AOI21_X1 U17770 ( .B1(n14470), .B2(n14448), .A(n14426), .ZN(n14436) );
  INV_X1 U17771 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15926) );
  AOI22_X1 U17772 ( .A1(n14427), .A2(n15926), .B1(n9834), .B2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14428) );
  NAND2_X1 U17773 ( .A1(n14436), .A2(n14428), .ZN(n14429) );
  XOR2_X1 U17774 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14429), .Z(
        n14570) );
  NAND2_X1 U17775 ( .A1(n13376), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14566) );
  OAI21_X1 U17776 ( .B1(n15918), .B2(n14430), .A(n14566), .ZN(n14433) );
  NOR2_X1 U17777 ( .A1(n14431), .A2(n20101), .ZN(n14432) );
  OAI21_X1 U17779 ( .B1(n19877), .B2(n14570), .A(n14435), .ZN(P1_U2971) );
  NAND2_X1 U17780 ( .A1(n14436), .A2(n14447), .ZN(n14437) );
  XOR2_X1 U17781 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n14437), .Z(
        n15920) );
  INV_X1 U17782 ( .A(n14438), .ZN(n14440) );
  AOI22_X1 U17783 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n13376), .B2(P1_REIP_REG_27__SCAN_IN), .ZN(n14439) );
  OAI21_X1 U17784 ( .B1(n15914), .B2(n14440), .A(n14439), .ZN(n14441) );
  AOI21_X1 U17785 ( .B1(n14442), .B2(n15909), .A(n14441), .ZN(n14443) );
  OAI21_X1 U17786 ( .B1(n19877), .B2(n15920), .A(n14443), .ZN(P1_U2972) );
  INV_X1 U17787 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14444) );
  NAND2_X1 U17788 ( .A1(n13376), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14578) );
  OAI21_X1 U17789 ( .B1(n15918), .B2(n14444), .A(n14578), .ZN(n14445) );
  AOI21_X1 U17790 ( .B1(n14446), .B2(n15889), .A(n14445), .ZN(n14451) );
  NAND2_X1 U17791 ( .A1(n14449), .A2(n14448), .ZN(n14571) );
  NAND3_X1 U17792 ( .A1(n14572), .A2(n14571), .A3(n20074), .ZN(n14450) );
  OAI211_X1 U17793 ( .C1(n14452), .C2(n20101), .A(n14451), .B(n14450), .ZN(
        P1_U2973) );
  INV_X1 U17794 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15835) );
  AOI21_X1 U17795 ( .B1(n14453), .B2(n15831), .A(n15835), .ZN(n15824) );
  NOR2_X1 U17796 ( .A1(n15824), .A2(n15832), .ZN(n14454) );
  MUX2_X1 U17797 ( .A(n15824), .B(n14454), .S(n9834), .Z(n14455) );
  XNOR2_X1 U17798 ( .A(n14455), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14589) );
  NAND2_X1 U17799 ( .A1(n13376), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14584) );
  OAI21_X1 U17800 ( .B1(n15918), .B2(n15728), .A(n14584), .ZN(n14457) );
  NOR2_X1 U17801 ( .A1(n15731), .A2(n20101), .ZN(n14456) );
  AOI211_X1 U17802 ( .C1(n15889), .C2(n15726), .A(n14457), .B(n14456), .ZN(
        n14458) );
  OAI21_X1 U17803 ( .B1(n19877), .B2(n14589), .A(n14458), .ZN(P1_U2975) );
  NAND2_X1 U17804 ( .A1(n14460), .A2(n14459), .ZN(n14462) );
  XNOR2_X1 U17805 ( .A(n14462), .B(n14461), .ZN(n15952) );
  NAND2_X1 U17806 ( .A1(n15749), .A2(n15909), .ZN(n14467) );
  INV_X1 U17807 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14463) );
  OAI22_X1 U17808 ( .A1(n15918), .A2(n14464), .B1(n15996), .B2(n14463), .ZN(
        n14465) );
  AOI21_X1 U17809 ( .B1(n15889), .B2(n15747), .A(n14465), .ZN(n14466) );
  OAI211_X1 U17810 ( .C1(n15952), .C2(n19877), .A(n14467), .B(n14466), .ZN(
        P1_U2977) );
  INV_X1 U17811 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n14468) );
  OAI22_X1 U17812 ( .A1(n15918), .A2(n15774), .B1(n15996), .B2(n14468), .ZN(
        n14469) );
  AOI21_X1 U17813 ( .B1(n15889), .B2(n15764), .A(n14469), .ZN(n14476) );
  INV_X1 U17814 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14518) );
  NOR2_X1 U17815 ( .A1(n14471), .A2(n14470), .ZN(n14473) );
  INV_X1 U17816 ( .A(n14473), .ZN(n14472) );
  NAND3_X1 U17817 ( .A1(n14472), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n15666), .ZN(n14474) );
  NAND2_X1 U17818 ( .A1(n14473), .A2(n15674), .ZN(n15665) );
  OAI211_X1 U17819 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15666), .A(
        n14474), .B(n15665), .ZN(n15702) );
  NAND2_X1 U17820 ( .A1(n15702), .A2(n20074), .ZN(n14475) );
  OAI211_X1 U17821 ( .C1(n15765), .C2(n20101), .A(n14476), .B(n14475), .ZN(
        P1_U2979) );
  OAI21_X1 U17822 ( .B1(n15918), .B2(n14478), .A(n14477), .ZN(n14479) );
  AOI21_X1 U17823 ( .B1(n14480), .B2(n15889), .A(n14479), .ZN(n14483) );
  NAND3_X1 U17824 ( .A1(n14481), .A2(n15853), .A3(n20074), .ZN(n14482) );
  OAI211_X1 U17825 ( .C1(n14484), .C2(n20101), .A(n14483), .B(n14482), .ZN(
        P1_U2981) );
  INV_X1 U17826 ( .A(n15792), .ZN(n14486) );
  AOI22_X1 U17827 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n13376), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n14485) );
  OAI21_X1 U17828 ( .B1(n15914), .B2(n14486), .A(n14485), .ZN(n14487) );
  AOI21_X1 U17829 ( .B1(n14488), .B2(n15909), .A(n14487), .ZN(n14489) );
  OAI21_X1 U17830 ( .B1(n14490), .B2(n19877), .A(n14489), .ZN(P1_U2983) );
  INV_X1 U17831 ( .A(n13982), .ZN(n15892) );
  INV_X1 U17832 ( .A(n14491), .ZN(n14492) );
  AOI22_X1 U17833 ( .A1(n15892), .A2(n14493), .B1(n9834), .B2(n14492), .ZN(
        n15884) );
  INV_X1 U17834 ( .A(n14495), .ZN(n14494) );
  AOI21_X1 U17835 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n9834), .A(
        n14494), .ZN(n15883) );
  NAND2_X1 U17836 ( .A1(n15884), .A2(n15883), .ZN(n15882) );
  NAND2_X1 U17837 ( .A1(n15882), .A2(n14495), .ZN(n14496) );
  XOR2_X1 U17838 ( .A(n14497), .B(n14496), .Z(n15990) );
  NAND2_X1 U17839 ( .A1(n15990), .A2(n20074), .ZN(n14503) );
  INV_X1 U17840 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n14498) );
  OAI22_X1 U17841 ( .A1(n15918), .A2(n14499), .B1(n15996), .B2(n14498), .ZN(
        n14500) );
  AOI21_X1 U17842 ( .B1(n15889), .B2(n14501), .A(n14500), .ZN(n14502) );
  OAI211_X1 U17843 ( .C1(n20101), .C2(n14504), .A(n14503), .B(n14502), .ZN(
        P1_U2986) );
  NAND2_X1 U17844 ( .A1(n14505), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14507) );
  XNOR2_X1 U17845 ( .A(n13982), .B(n14508), .ZN(n14506) );
  MUX2_X1 U17846 ( .A(n14507), .B(n14506), .S(n13705), .Z(n14510) );
  INV_X1 U17847 ( .A(n14505), .ZN(n14509) );
  NAND3_X1 U17848 ( .A1(n14509), .A2(n15855), .A3(n14508), .ZN(n15893) );
  NAND2_X1 U17849 ( .A1(n14510), .A2(n15893), .ZN(n16019) );
  NAND2_X1 U17850 ( .A1(n16019), .A2(n20074), .ZN(n14515) );
  INV_X1 U17851 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14511) );
  NOR2_X1 U17852 ( .A1(n15996), .A2(n14511), .ZN(n16016) );
  NOR2_X1 U17853 ( .A1(n15914), .A2(n14512), .ZN(n14513) );
  AOI211_X1 U17854 ( .C1(n20076), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16016), .B(n14513), .ZN(n14514) );
  OAI211_X1 U17855 ( .C1(n20101), .C2(n14516), .A(n14515), .B(n14514), .ZN(
        P1_U2989) );
  NAND2_X1 U17856 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14573) );
  NAND2_X1 U17857 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15956) );
  NOR2_X1 U17858 ( .A1(n15674), .A2(n14518), .ZN(n14525) );
  NOR2_X1 U17859 ( .A1(n15852), .A2(n14519), .ZN(n15672) );
  NAND2_X1 U17860 ( .A1(n14520), .A2(n15672), .ZN(n15673) );
  AOI21_X1 U17861 ( .B1(n15672), .B2(n14521), .A(n14526), .ZN(n14523) );
  AOI211_X1 U17862 ( .C1(n16029), .C2(n15673), .A(n14523), .B(n14522), .ZN(
        n15964) );
  AOI21_X1 U17863 ( .B1(n14525), .B2(n15964), .A(n14524), .ZN(n15951) );
  AOI21_X1 U17864 ( .B1(n16032), .B2(n15956), .A(n15951), .ZN(n15950) );
  OAI21_X1 U17865 ( .B1(n14526), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15950), .ZN(n14581) );
  AOI21_X1 U17866 ( .B1(n14573), .B2(n16032), .A(n14581), .ZN(n15936) );
  NAND2_X1 U17867 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15936), .ZN(
        n14574) );
  INV_X1 U17868 ( .A(n14574), .ZN(n14528) );
  INV_X1 U17869 ( .A(n15950), .ZN(n14527) );
  NOR2_X1 U17870 ( .A1(n14527), .A2(n16032), .ZN(n14555) );
  AOI21_X1 U17871 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14528), .A(
        n14555), .ZN(n15928) );
  INV_X1 U17872 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14535) );
  NOR2_X1 U17873 ( .A1(n15928), .A2(n14535), .ZN(n14554) );
  AOI21_X1 U17874 ( .B1(n14554), .B2(n14561), .A(n14555), .ZN(n14529) );
  NOR2_X1 U17875 ( .A1(n14529), .A2(n14545), .ZN(n14543) );
  INV_X1 U17876 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14598) );
  NOR3_X1 U17877 ( .A1(n14543), .A2(n14555), .A3(n14598), .ZN(n14539) );
  NOR2_X1 U17878 ( .A1(n14530), .A2(n20084), .ZN(n14538) );
  INV_X1 U17879 ( .A(n14531), .ZN(n14537) );
  NAND4_X1 U17880 ( .A1(n14533), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n15672), .A4(n14532), .ZN(n15942) );
  NOR2_X1 U17881 ( .A1(n14534), .A2(n15942), .ZN(n14575) );
  NAND2_X1 U17882 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n14575), .ZN(
        n14562) );
  INV_X1 U17883 ( .A(n14562), .ZN(n15927) );
  NAND2_X1 U17884 ( .A1(n15927), .A2(n14561), .ZN(n14553) );
  NOR4_X1 U17885 ( .A1(n14553), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14545), .A4(n14535), .ZN(n14536) );
  NOR4_X1 U17886 ( .A1(n14539), .A2(n14538), .A3(n14537), .A4(n14536), .ZN(
        n14540) );
  OAI21_X1 U17887 ( .B1(n14541), .B2(n16008), .A(n14540), .ZN(P1_U3000) );
  INV_X1 U17888 ( .A(n14542), .ZN(n14547) );
  NAND3_X1 U17889 ( .A1(n15927), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14561), .ZN(n14544) );
  AOI21_X1 U17890 ( .B1(n14545), .B2(n14544), .A(n14543), .ZN(n14546) );
  AOI211_X1 U17891 ( .C1(n14548), .C2(n16018), .A(n14547), .B(n14546), .ZN(
        n14549) );
  OAI21_X1 U17892 ( .B1(n14550), .B2(n16008), .A(n14549), .ZN(P1_U3001) );
  AOI21_X1 U17893 ( .B1(n14552), .B2(n16018), .A(n14551), .ZN(n14559) );
  INV_X1 U17894 ( .A(n14553), .ZN(n14557) );
  OAI21_X1 U17895 ( .B1(n14561), .B2(n14555), .A(n14554), .ZN(n14556) );
  OAI21_X1 U17896 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n14557), .A(
        n14556), .ZN(n14558) );
  OAI211_X1 U17897 ( .C1(n14560), .C2(n16008), .A(n14559), .B(n14558), .ZN(
        P1_U3002) );
  NOR2_X1 U17898 ( .A1(n14563), .A2(n14562), .ZN(n14564) );
  NAND2_X1 U17899 ( .A1(n9829), .A2(n14564), .ZN(n14565) );
  OAI211_X1 U17900 ( .C1(n14567), .C2(n20084), .A(n14566), .B(n14565), .ZN(
        n14568) );
  AOI21_X1 U17901 ( .B1(n15928), .B2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14568), .ZN(n14569) );
  OAI21_X1 U17902 ( .B1(n14570), .B2(n16008), .A(n14569), .ZN(P1_U3003) );
  NAND3_X1 U17903 ( .A1(n14572), .A2(n14571), .A3(n20087), .ZN(n14580) );
  NOR3_X1 U17904 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n14573), .A3(
        n15942), .ZN(n15933) );
  OAI22_X1 U17905 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n14575), .B1(
        n15933), .B2(n14574), .ZN(n14579) );
  NAND2_X1 U17906 ( .A1(n14576), .A2(n16018), .ZN(n14577) );
  NAND4_X1 U17907 ( .A1(n14580), .A2(n14579), .A3(n14578), .A4(n14577), .ZN(
        P1_U3005) );
  INV_X1 U17908 ( .A(n14581), .ZN(n14582) );
  OAI21_X1 U17909 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14583), .A(
        n14582), .ZN(n14587) );
  NOR3_X1 U17910 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15835), .A3(
        n15942), .ZN(n14586) );
  OAI21_X1 U17911 ( .B1(n15730), .B2(n20084), .A(n14584), .ZN(n14585) );
  AOI211_X1 U17912 ( .C1(n14587), .C2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n14586), .B(n14585), .ZN(n14588) );
  OAI21_X1 U17913 ( .B1(n14589), .B2(n16008), .A(n14588), .ZN(P1_U3007) );
  OAI21_X1 U17914 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n13020), .A(n20548), 
        .ZN(n14590) );
  OAI21_X1 U17915 ( .B1(n20673), .B2(n14591), .A(n14590), .ZN(n14592) );
  MUX2_X1 U17916 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14592), .S(
        n20883), .Z(P1_U3477) );
  NOR2_X1 U17917 ( .A1(n14593), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14596) );
  NOR3_X1 U17918 ( .A1(n14594), .A2(n14600), .A3(n14599), .ZN(n14595) );
  AOI211_X1 U17919 ( .C1(n9946), .C2(n14597), .A(n14596), .B(n14595), .ZN(
        n15633) );
  OAI22_X1 U17920 ( .A1(n14598), .A2(n12643), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14605) );
  NOR2_X1 U17921 ( .A1(n21068), .A2(n20091), .ZN(n14607) );
  NOR3_X1 U17922 ( .A1(n14600), .A2(n14599), .A3(n14614), .ZN(n14601) );
  AOI21_X1 U17923 ( .B1(n14605), .B2(n14607), .A(n14601), .ZN(n14602) );
  OAI21_X1 U17924 ( .B1(n15633), .B2(n14616), .A(n14602), .ZN(n14604) );
  INV_X1 U17925 ( .A(n14603), .ZN(n16075) );
  MUX2_X1 U17926 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14604), .S(
        n16075), .Z(P1_U3473) );
  INV_X1 U17927 ( .A(n14605), .ZN(n14606) );
  AOI22_X1 U17928 ( .A1(n14609), .A2(n14608), .B1(n14607), .B2(n14606), .ZN(
        n14610) );
  OAI21_X1 U17929 ( .B1(n14611), .B2(n14616), .A(n14610), .ZN(n14612) );
  MUX2_X1 U17930 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14612), .S(
        n16075), .Z(P1_U3472) );
  INV_X1 U17931 ( .A(n14613), .ZN(n14617) );
  OAI22_X1 U17932 ( .A1(n14617), .A2(n14616), .B1(n14615), .B2(n14614), .ZN(
        n14618) );
  MUX2_X1 U17933 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14618), .S(
        n16075), .Z(P1_U3469) );
  XNOR2_X1 U17934 ( .A(n14620), .B(n14619), .ZN(n14628) );
  NAND2_X1 U17935 ( .A1(n14995), .A2(n19061), .ZN(n14627) );
  INV_X1 U17936 ( .A(n14938), .ZN(n14625) );
  OAI22_X1 U17937 ( .A1(n19001), .A2(n10960), .B1(n14621), .B2(n19043), .ZN(
        n14624) );
  AOI22_X1 U17938 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19045), .ZN(n14622) );
  INV_X1 U17939 ( .A(n14622), .ZN(n14623) );
  AOI211_X1 U17940 ( .C1(n14625), .C2(n19064), .A(n14624), .B(n14623), .ZN(
        n14626) );
  OAI211_X1 U17941 ( .C1(n14628), .C2(n19077), .A(n14627), .B(n14626), .ZN(
        P2_U2825) );
  NOR2_X1 U17942 ( .A1(n14630), .A2(n14631), .ZN(n14632) );
  OR2_X1 U17943 ( .A1(n14629), .A2(n14632), .ZN(n16186) );
  NAND2_X1 U17944 ( .A1(n14634), .A2(n14633), .ZN(n14635) );
  NAND2_X1 U17945 ( .A1(n14987), .A2(n14635), .ZN(n16174) );
  INV_X1 U17946 ( .A(n16174), .ZN(n14643) );
  NAND2_X1 U17947 ( .A1(n19041), .A2(n19036), .ZN(n18943) );
  OAI22_X1 U17948 ( .A1(n14636), .A2(n19043), .B1(n18943), .B2(n15171), .ZN(
        n14642) );
  AOI22_X1 U17949 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19028), .B1(
        P2_EBX_REG_20__SCAN_IN), .B2(n19059), .ZN(n14640) );
  OAI211_X1 U17950 ( .C1(n14638), .C2(n15171), .A(n18910), .B(n14637), .ZN(
        n14639) );
  OAI211_X1 U17951 ( .C1(n19068), .C2(n19789), .A(n14640), .B(n14639), .ZN(
        n14641) );
  AOI211_X1 U17952 ( .C1(n19064), .C2(n14643), .A(n14642), .B(n14641), .ZN(
        n14644) );
  OAI21_X1 U17953 ( .B1(n16186), .B2(n19049), .A(n14644), .ZN(P2_U2835) );
  AOI21_X1 U17954 ( .B1(n14645), .B2(n15365), .A(n14630), .ZN(n15358) );
  INV_X1 U17955 ( .A(n15358), .ZN(n14655) );
  NAND2_X1 U17956 ( .A1(n9690), .A2(n14646), .ZN(n14647) );
  XNOR2_X1 U17957 ( .A(n15180), .B(n14647), .ZN(n14653) );
  INV_X1 U17958 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19787) );
  AOI22_X1 U17959 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(n19059), .B1(n14648), 
        .B2(n19057), .ZN(n14649) );
  OAI211_X1 U17960 ( .C1(n19787), .C2(n19068), .A(n14649), .B(n19046), .ZN(
        n14650) );
  AOI21_X1 U17961 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n19028), .A(
        n14650), .ZN(n14651) );
  OAI21_X1 U17962 ( .B1(n15183), .B2(n19011), .A(n14651), .ZN(n14652) );
  AOI21_X1 U17963 ( .B1(n14653), .B2(n19036), .A(n14652), .ZN(n14654) );
  OAI21_X1 U17964 ( .B1(n14655), .B2(n19049), .A(n14654), .ZN(P2_U2836) );
  NAND2_X1 U17965 ( .A1(n19835), .A2(n19061), .ZN(n14661) );
  AOI22_X1 U17966 ( .A1(P2_EBX_REG_2__SCAN_IN), .A2(n19059), .B1(n14656), .B2(
        n19057), .ZN(n14660) );
  AOI22_X1 U17967 ( .A1(P2_REIP_REG_2__SCAN_IN), .A2(n19045), .B1(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19028), .ZN(n14659) );
  NAND2_X1 U17968 ( .A1(n14657), .A2(n19064), .ZN(n14658) );
  NAND4_X1 U17969 ( .A1(n14661), .A2(n14660), .A3(n14659), .A4(n14658), .ZN(
        n14667) );
  NOR2_X1 U17970 ( .A1(n19041), .A2(n14662), .ZN(n14677) );
  INV_X1 U17971 ( .A(n14677), .ZN(n14663) );
  AOI221_X1 U17972 ( .B1(n14665), .B2(n14677), .C1(n14664), .C2(n14663), .A(
        n19077), .ZN(n14666) );
  AOI211_X1 U17973 ( .C1(n19074), .C2(n15468), .A(n14667), .B(n14666), .ZN(
        n14668) );
  INV_X1 U17974 ( .A(n14668), .ZN(P2_U2853) );
  AOI22_X1 U17975 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_1__SCAN_IN), .B2(n19045), .ZN(n14676) );
  INV_X1 U17976 ( .A(n14669), .ZN(n14672) );
  AOI22_X1 U17977 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(n19059), .B1(n19061), .B2(
        n19844), .ZN(n14670) );
  OAI21_X1 U17978 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18943), .A(
        n14670), .ZN(n14671) );
  AOI21_X1 U17979 ( .B1(n19057), .B2(n14672), .A(n14671), .ZN(n14675) );
  OR2_X1 U17980 ( .A1(n14673), .A2(n19011), .ZN(n14674) );
  NAND3_X1 U17981 ( .A1(n14676), .A2(n14675), .A3(n14674), .ZN(n14680) );
  OAI21_X1 U17982 ( .B1(n15450), .B2(n14678), .A(n14677), .ZN(n15455) );
  NOR2_X1 U17983 ( .A1(n15455), .A2(n19077), .ZN(n14679) );
  AOI211_X1 U17984 ( .C1(n19074), .C2(n19842), .A(n14680), .B(n14679), .ZN(
        n14681) );
  INV_X1 U17985 ( .A(n14681), .ZN(P2_U2854) );
  AOI22_X1 U17986 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14686) );
  NAND2_X1 U17987 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n14685) );
  NAND2_X1 U17988 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n14684) );
  NAND2_X1 U17989 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14683) );
  NAND4_X1 U17990 ( .A1(n14686), .A2(n14685), .A3(n14684), .A4(n14683), .ZN(
        n14690) );
  INV_X1 U17991 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14688) );
  INV_X1 U17992 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14687) );
  OAI22_X1 U17993 ( .A1(n14688), .A2(n10464), .B1(n10463), .B2(n14687), .ZN(
        n14689) );
  NOR2_X1 U17994 ( .A1(n14690), .A2(n14689), .ZN(n14703) );
  OR2_X1 U17995 ( .A1(n10467), .A2(n19248), .ZN(n14694) );
  AOI22_X1 U17996 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14693) );
  NAND2_X1 U17997 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n14692) );
  NAND2_X1 U17998 ( .A1(n10447), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14691) );
  AND4_X1 U17999 ( .A1(n14694), .A2(n14693), .A3(n14692), .A4(n14691), .ZN(
        n14702) );
  OAI22_X1 U18000 ( .A1(n10472), .A2(n14696), .B1(n14738), .B2(n14695), .ZN(
        n14700) );
  INV_X1 U18001 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14698) );
  OAI22_X1 U18002 ( .A1(n14698), .A2(n11114), .B1(n10473), .B2(n14697), .ZN(
        n14699) );
  NOR2_X1 U18003 ( .A1(n14700), .A2(n14699), .ZN(n14701) );
  AOI22_X1 U18004 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14708) );
  NAND2_X1 U18005 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n14707) );
  NAND2_X1 U18006 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n14706) );
  NAND2_X1 U18007 ( .A1(n14782), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14705) );
  NAND4_X1 U18008 ( .A1(n14708), .A2(n14707), .A3(n14706), .A4(n14705), .ZN(
        n14712) );
  INV_X1 U18009 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14710) );
  OAI22_X1 U18010 ( .A1(n14710), .A2(n10464), .B1(n10463), .B2(n14709), .ZN(
        n14711) );
  NOR2_X1 U18011 ( .A1(n14712), .A2(n14711), .ZN(n14724) );
  AOI22_X1 U18012 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n14713) );
  OAI21_X1 U18013 ( .B1(n21045), .B2(n10467), .A(n14713), .ZN(n14714) );
  INV_X1 U18014 ( .A(n14714), .ZN(n14723) );
  OAI22_X1 U18015 ( .A1(n10472), .A2(n14716), .B1(n14738), .B2(n14715), .ZN(
        n14720) );
  OAI22_X1 U18016 ( .A1(n14718), .A2(n11114), .B1(n10473), .B2(n14717), .ZN(
        n14719) );
  NOR2_X1 U18017 ( .A1(n14720), .A2(n14719), .ZN(n14722) );
  AOI22_X1 U18018 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10447), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14721) );
  NAND4_X1 U18019 ( .A1(n14724), .A2(n14723), .A3(n14722), .A4(n14721), .ZN(
        n14984) );
  INV_X1 U18020 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14726) );
  INV_X1 U18021 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14725) );
  OAI22_X1 U18022 ( .A1(n14726), .A2(n10158), .B1(n9717), .B2(n14725), .ZN(
        n14732) );
  OAI22_X1 U18023 ( .A1(n14730), .A2(n14729), .B1(n14728), .B2(n14727), .ZN(
        n14731) );
  AOI211_X1 U18024 ( .C1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .C2(n9714), .A(
        n14732), .B(n14731), .ZN(n14747) );
  AOI22_X1 U18025 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n14734), .B1(
        n14733), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14746) );
  AOI22_X1 U18026 ( .A1(n10426), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n10447), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14736) );
  AOI22_X1 U18027 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n14735) );
  OAI211_X1 U18028 ( .C1(n10467), .C2(n19255), .A(n14736), .B(n14735), .ZN(
        n14744) );
  OAI22_X1 U18029 ( .A1(n10472), .A2(n14739), .B1(n14738), .B2(n14737), .ZN(
        n14743) );
  OAI22_X1 U18030 ( .A1(n14741), .A2(n11114), .B1(n10473), .B2(n14740), .ZN(
        n14742) );
  NOR3_X1 U18031 ( .A1(n14744), .A2(n14743), .A3(n14742), .ZN(n14745) );
  NAND3_X1 U18032 ( .A1(n14747), .A2(n14746), .A3(n14745), .ZN(n15065) );
  AOI22_X1 U18033 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14756) );
  AOI22_X1 U18034 ( .A1(n14928), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n14826), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14755) );
  AOI22_X1 U18035 ( .A1(n14929), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14754) );
  AND2_X1 U18036 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14750) );
  OR2_X1 U18037 ( .A1(n14750), .A2(n14749), .ZN(n14926) );
  INV_X1 U18038 ( .A(n14926), .ZN(n14902) );
  NAND2_X1 U18039 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14751) );
  AND3_X1 U18040 ( .A1(n14902), .A2(n14752), .A3(n14751), .ZN(n14753) );
  NAND4_X1 U18041 ( .A1(n14756), .A2(n14755), .A3(n14754), .A4(n14753), .ZN(
        n14765) );
  AOI22_X1 U18042 ( .A1(n14757), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n14763) );
  AOI22_X1 U18043 ( .A1(n14928), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14826), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14762) );
  AOI22_X1 U18044 ( .A1(n14929), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10397), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14761) );
  NAND2_X1 U18045 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n14758) );
  AND3_X1 U18046 ( .A1(n14759), .A2(n14926), .A3(n14758), .ZN(n14760) );
  NAND4_X1 U18047 ( .A1(n14763), .A2(n14762), .A3(n14761), .A4(n14760), .ZN(
        n14764) );
  NAND2_X1 U18048 ( .A1(n14765), .A2(n14764), .ZN(n14814) );
  NOR2_X1 U18049 ( .A1(n19231), .A2(n14814), .ZN(n14791) );
  AOI22_X1 U18050 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n14767), .B1(
        n14766), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14768) );
  OAI21_X1 U18051 ( .B1(n10467), .B2(n19265), .A(n14768), .ZN(n14769) );
  INV_X1 U18052 ( .A(n14769), .ZN(n14778) );
  AOI22_X1 U18053 ( .A1(n14770), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10447), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14777) );
  AOI22_X1 U18054 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10426), .B1(
        n14771), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14776) );
  INV_X1 U18055 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14773) );
  OAI22_X1 U18056 ( .A1(n14773), .A2(n11114), .B1(n10473), .B2(n14772), .ZN(
        n14774) );
  INV_X1 U18057 ( .A(n14774), .ZN(n14775) );
  NAND4_X1 U18058 ( .A1(n14778), .A2(n14777), .A3(n14776), .A4(n14775), .ZN(
        n14790) );
  INV_X1 U18059 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14780) );
  OAI22_X1 U18060 ( .A1(n14780), .A2(n10464), .B1(n10463), .B2(n14779), .ZN(
        n14781) );
  INV_X1 U18061 ( .A(n14781), .ZN(n14788) );
  AOI22_X1 U18062 ( .A1(n9714), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n14782), .ZN(n14787) );
  AOI22_X1 U18063 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n14783), .B1(
        n14682), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14786) );
  NAND2_X1 U18064 ( .A1(n14784), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n14785) );
  NAND4_X1 U18065 ( .A1(n14788), .A2(n14787), .A3(n14786), .A4(n14785), .ZN(
        n14789) );
  NOR2_X1 U18066 ( .A1(n14790), .A2(n14789), .ZN(n14809) );
  XNOR2_X1 U18067 ( .A(n14791), .B(n14809), .ZN(n14816) );
  INV_X1 U18068 ( .A(n14814), .ZN(n14810) );
  NAND2_X1 U18069 ( .A1(n19231), .A2(n14810), .ZN(n15057) );
  AOI22_X1 U18070 ( .A1(n14928), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14800) );
  AOI22_X1 U18071 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14826), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14799) );
  AOI22_X1 U18072 ( .A1(n14929), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14798) );
  NAND2_X1 U18073 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n14795) );
  AND3_X1 U18074 ( .A1(n14902), .A2(n14796), .A3(n14795), .ZN(n14797) );
  NAND4_X1 U18075 ( .A1(n14800), .A2(n14799), .A3(n14798), .A4(n14797), .ZN(
        n14808) );
  AOI22_X1 U18076 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n14928), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14806) );
  AOI22_X1 U18077 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14826), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14805) );
  AOI22_X1 U18078 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n14929), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14804) );
  NAND2_X1 U18079 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n14801) );
  AND3_X1 U18080 ( .A1(n14802), .A2(n14926), .A3(n14801), .ZN(n14803) );
  NAND4_X1 U18081 ( .A1(n14806), .A2(n14805), .A3(n14804), .A4(n14803), .ZN(
        n14807) );
  NAND2_X1 U18082 ( .A1(n14808), .A2(n14807), .ZN(n14813) );
  INV_X1 U18083 ( .A(n14809), .ZN(n14811) );
  NAND2_X1 U18084 ( .A1(n14811), .A2(n14810), .ZN(n14817) );
  XOR2_X1 U18085 ( .A(n14813), .B(n14817), .Z(n14812) );
  NAND2_X1 U18086 ( .A1(n14812), .A2(n14876), .ZN(n14973) );
  INV_X1 U18087 ( .A(n14813), .ZN(n14818) );
  NAND2_X1 U18088 ( .A1(n19231), .A2(n14818), .ZN(n14976) );
  NOR2_X1 U18089 ( .A1(n14976), .A2(n14814), .ZN(n14815) );
  INV_X1 U18090 ( .A(n14817), .ZN(n14819) );
  AND2_X1 U18091 ( .A1(n14819), .A2(n14818), .ZN(n14835) );
  AOI22_X1 U18092 ( .A1(n14928), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14825) );
  AOI22_X1 U18093 ( .A1(n14757), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14826), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14824) );
  AOI22_X1 U18094 ( .A1(n14929), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10397), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14823) );
  NAND2_X1 U18095 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14820) );
  AND3_X1 U18096 ( .A1(n14902), .A2(n14821), .A3(n14820), .ZN(n14822) );
  NAND4_X1 U18097 ( .A1(n14825), .A2(n14824), .A3(n14823), .A4(n14822), .ZN(
        n14834) );
  AOI22_X1 U18098 ( .A1(n14928), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14748), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14832) );
  AOI22_X1 U18099 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14826), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14831) );
  AOI22_X1 U18100 ( .A1(n14929), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14830) );
  NAND2_X1 U18101 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n14827) );
  AND3_X1 U18102 ( .A1(n14828), .A2(n14926), .A3(n14827), .ZN(n14829) );
  NAND4_X1 U18103 ( .A1(n14832), .A2(n14831), .A3(n14830), .A4(n14829), .ZN(
        n14833) );
  AND2_X1 U18104 ( .A1(n14834), .A2(n14833), .ZN(n14836) );
  NAND2_X1 U18105 ( .A1(n14835), .A2(n14836), .ZN(n14859) );
  OAI211_X1 U18106 ( .C1(n14835), .C2(n14836), .A(n14876), .B(n14859), .ZN(
        n14839) );
  INV_X1 U18107 ( .A(n14836), .ZN(n14837) );
  NOR2_X1 U18108 ( .A1(n11027), .A2(n14837), .ZN(n14967) );
  AOI22_X1 U18109 ( .A1(n14928), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14847) );
  AOI22_X1 U18110 ( .A1(n14757), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14927), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14846) );
  AOI22_X1 U18111 ( .A1(n14929), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10397), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14845) );
  NAND2_X1 U18112 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n14842) );
  AND3_X1 U18113 ( .A1(n14902), .A2(n14843), .A3(n14842), .ZN(n14844) );
  NAND4_X1 U18114 ( .A1(n14847), .A2(n14846), .A3(n14845), .A4(n14844), .ZN(
        n14855) );
  AOI22_X1 U18115 ( .A1(n14928), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14748), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n14853) );
  AOI22_X1 U18116 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14927), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14852) );
  AOI22_X1 U18117 ( .A1(n14929), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14851) );
  NAND2_X1 U18118 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n14848) );
  AND3_X1 U18119 ( .A1(n14849), .A2(n14926), .A3(n14848), .ZN(n14850) );
  NAND4_X1 U18120 ( .A1(n14853), .A2(n14852), .A3(n14851), .A4(n14850), .ZN(
        n14854) );
  AND2_X1 U18121 ( .A1(n14855), .A2(n14854), .ZN(n14860) );
  XNOR2_X1 U18122 ( .A(n14859), .B(n14860), .ZN(n14856) );
  NAND2_X1 U18123 ( .A1(n19231), .A2(n14860), .ZN(n14962) );
  INV_X1 U18124 ( .A(n14859), .ZN(n14861) );
  AND2_X1 U18125 ( .A1(n14861), .A2(n14860), .ZN(n14877) );
  AOI22_X1 U18126 ( .A1(n14928), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14867) );
  AOI22_X1 U18127 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14927), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14866) );
  AOI22_X1 U18128 ( .A1(n14929), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10397), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14865) );
  NAND2_X1 U18129 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n14862) );
  AND3_X1 U18130 ( .A1(n14902), .A2(n14863), .A3(n14862), .ZN(n14864) );
  NAND4_X1 U18131 ( .A1(n14867), .A2(n14866), .A3(n14865), .A4(n14864), .ZN(
        n14875) );
  AOI22_X1 U18132 ( .A1(n14928), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14748), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n14873) );
  AOI22_X1 U18133 ( .A1(n14757), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14927), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14872) );
  AOI22_X1 U18134 ( .A1(n14929), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14871) );
  NAND2_X1 U18135 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n14868) );
  AND3_X1 U18136 ( .A1(n14869), .A2(n14926), .A3(n14868), .ZN(n14870) );
  NAND4_X1 U18137 ( .A1(n14873), .A2(n14872), .A3(n14871), .A4(n14870), .ZN(
        n14874) );
  AND2_X1 U18138 ( .A1(n14875), .A2(n14874), .ZN(n14881) );
  NAND2_X1 U18139 ( .A1(n14877), .A2(n14881), .ZN(n14896) );
  OAI211_X1 U18140 ( .C1(n14877), .C2(n14881), .A(n14876), .B(n14896), .ZN(
        n14878) );
  INV_X1 U18141 ( .A(n14948), .ZN(n14880) );
  NAND2_X1 U18142 ( .A1(n14880), .A2(n14879), .ZN(n14957) );
  NAND2_X1 U18143 ( .A1(n19231), .A2(n14881), .ZN(n14956) );
  AOI22_X1 U18144 ( .A1(n14928), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14887) );
  AOI22_X1 U18145 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14927), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14886) );
  AOI22_X1 U18146 ( .A1(n14929), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14885) );
  NAND2_X1 U18147 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n14882) );
  AND3_X1 U18148 ( .A1(n14902), .A2(n14883), .A3(n14882), .ZN(n14884) );
  NAND4_X1 U18149 ( .A1(n14887), .A2(n14886), .A3(n14885), .A4(n14884), .ZN(
        n14895) );
  AOI22_X1 U18150 ( .A1(n14928), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14748), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n14893) );
  AOI22_X1 U18151 ( .A1(n14757), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14927), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14892) );
  AOI22_X1 U18152 ( .A1(n14929), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10397), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14891) );
  NAND2_X1 U18153 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n14888) );
  AND3_X1 U18154 ( .A1(n14889), .A2(n14926), .A3(n14888), .ZN(n14890) );
  NAND4_X1 U18155 ( .A1(n14893), .A2(n14892), .A3(n14891), .A4(n14890), .ZN(
        n14894) );
  AND2_X1 U18156 ( .A1(n14895), .A2(n14894), .ZN(n14897) );
  OAI21_X1 U18157 ( .B1(n14955), .B2(n14948), .A(n14897), .ZN(n14943) );
  INV_X1 U18158 ( .A(n14896), .ZN(n14947) );
  INV_X1 U18159 ( .A(n14897), .ZN(n14949) );
  NOR2_X1 U18160 ( .A1(n19231), .A2(n14949), .ZN(n14898) );
  AND2_X1 U18161 ( .A1(n14947), .A2(n14898), .ZN(n14916) );
  AOI22_X1 U18162 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14906) );
  AOI22_X1 U18163 ( .A1(n14928), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n14927), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14905) );
  AOI22_X1 U18164 ( .A1(n14929), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9640), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14904) );
  NAND2_X1 U18165 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n14900) );
  AND3_X1 U18166 ( .A1(n14902), .A2(n14901), .A3(n14900), .ZN(n14903) );
  NAND4_X1 U18167 ( .A1(n14906), .A2(n14905), .A3(n14904), .A4(n14903), .ZN(
        n14914) );
  AOI22_X1 U18168 ( .A1(n14928), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14748), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n14912) );
  AOI22_X1 U18169 ( .A1(n14757), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14927), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14911) );
  AOI22_X1 U18170 ( .A1(n14929), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10397), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14910) );
  NAND2_X1 U18171 ( .A1(n10392), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n14907) );
  AND3_X1 U18172 ( .A1(n14908), .A2(n14926), .A3(n14907), .ZN(n14909) );
  NAND4_X1 U18173 ( .A1(n14912), .A2(n14911), .A3(n14910), .A4(n14909), .ZN(
        n14913) );
  AND2_X1 U18174 ( .A1(n14914), .A2(n14913), .ZN(n14915) );
  NAND2_X1 U18175 ( .A1(n14916), .A2(n14915), .ZN(n14917) );
  OAI21_X1 U18176 ( .B1(n14916), .B2(n14915), .A(n14917), .ZN(n14942) );
  INV_X1 U18177 ( .A(n14917), .ZN(n14918) );
  NOR2_X1 U18178 ( .A1(n14941), .A2(n14918), .ZN(n14937) );
  AOI22_X1 U18179 ( .A1(n9640), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n10392), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14921) );
  NAND2_X1 U18180 ( .A1(n14929), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n14919) );
  NAND4_X1 U18181 ( .A1(n14921), .A2(n14920), .A3(n14919), .A4(n14926), .ZN(
        n14935) );
  AOI22_X1 U18182 ( .A1(n14928), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14748), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14923) );
  AOI22_X1 U18183 ( .A1(n14757), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14927), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14922) );
  NAND2_X1 U18184 ( .A1(n14923), .A2(n14922), .ZN(n14934) );
  NOR2_X1 U18185 ( .A1(n13290), .A2(n14924), .ZN(n14925) );
  AOI22_X1 U18186 ( .A1(n9646), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14927), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14932) );
  AOI22_X1 U18187 ( .A1(n14928), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9645), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n14931) );
  AOI22_X1 U18188 ( .A1(n14929), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10397), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14930) );
  NAND4_X1 U18189 ( .A1(n9801), .A2(n14932), .A3(n14931), .A4(n14930), .ZN(
        n14933) );
  OAI21_X1 U18190 ( .B1(n14935), .B2(n14934), .A(n14933), .ZN(n14936) );
  XNOR2_X1 U18191 ( .A(n14937), .B(n14936), .ZN(n14997) );
  NOR2_X1 U18192 ( .A1(n14938), .A2(n19089), .ZN(n14939) );
  AOI21_X1 U18193 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19089), .A(n14939), .ZN(
        n14940) );
  OAI21_X1 U18194 ( .B1(n14997), .B2(n19095), .A(n14940), .ZN(P2_U2857) );
  INV_X1 U18195 ( .A(n14941), .ZN(n14999) );
  NAND2_X1 U18196 ( .A1(n14943), .A2(n14942), .ZN(n14998) );
  NAND3_X1 U18197 ( .A1(n14999), .A2(n19100), .A3(n14998), .ZN(n14945) );
  NAND2_X1 U18198 ( .A1(n19089), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14944) );
  OAI211_X1 U18199 ( .C1(n14946), .C2(n19089), .A(n14945), .B(n14944), .ZN(
        P2_U2858) );
  NOR2_X1 U18200 ( .A1(n14948), .A2(n14947), .ZN(n14950) );
  XNOR2_X1 U18201 ( .A(n14950), .B(n14949), .ZN(n15013) );
  NOR2_X1 U18202 ( .A1(n16098), .A2(n19089), .ZN(n14951) );
  AOI21_X1 U18203 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n19089), .A(n14951), .ZN(
        n14952) );
  OAI21_X1 U18204 ( .B1(n15013), .B2(n19095), .A(n14952), .ZN(P2_U2859) );
  AOI21_X1 U18205 ( .B1(n14954), .B2(n9720), .A(n14953), .ZN(n16109) );
  INV_X1 U18206 ( .A(n16109), .ZN(n14960) );
  AOI21_X1 U18207 ( .B1(n14957), .B2(n14956), .A(n14955), .ZN(n15016) );
  NAND2_X1 U18208 ( .A1(n15016), .A2(n19100), .ZN(n14959) );
  NAND2_X1 U18209 ( .A1(n19089), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14958) );
  OAI211_X1 U18210 ( .C1(n14960), .C2(n19089), .A(n14959), .B(n14958), .ZN(
        P2_U2860) );
  AOI21_X1 U18211 ( .B1(n14963), .B2(n14962), .A(n14961), .ZN(n15026) );
  NAND2_X1 U18212 ( .A1(n15026), .A2(n19100), .ZN(n14965) );
  NAND2_X1 U18213 ( .A1(n16120), .A2(n19103), .ZN(n14964) );
  OAI211_X1 U18214 ( .C1(n19103), .C2(n21077), .A(n14965), .B(n14964), .ZN(
        P2_U2861) );
  OAI21_X1 U18215 ( .B1(n14968), .B2(n14967), .A(n14966), .ZN(n15041) );
  OR2_X1 U18216 ( .A1(n14979), .A2(n14969), .ZN(n14970) );
  NAND2_X1 U18217 ( .A1(n11401), .A2(n14970), .ZN(n16131) );
  NOR2_X1 U18218 ( .A1(n16131), .A2(n19089), .ZN(n14971) );
  AOI21_X1 U18219 ( .B1(P2_EBX_REG_25__SCAN_IN), .B2(n19089), .A(n14971), .ZN(
        n14972) );
  OAI21_X1 U18220 ( .B1(n15041), .B2(n19095), .A(n14972), .ZN(P2_U2862) );
  AOI21_X1 U18221 ( .B1(n14974), .B2(n14973), .A(n9703), .ZN(n14975) );
  XOR2_X1 U18222 ( .A(n14976), .B(n14975), .Z(n15050) );
  AND2_X1 U18223 ( .A1(n15125), .A2(n14977), .ZN(n14978) );
  NOR2_X1 U18224 ( .A1(n14979), .A2(n14978), .ZN(n15295) );
  INV_X1 U18225 ( .A(n15295), .ZN(n16142) );
  NOR2_X1 U18226 ( .A1(n16142), .A2(n19089), .ZN(n14980) );
  AOI21_X1 U18227 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n19089), .A(n14980), .ZN(
        n14981) );
  OAI21_X1 U18228 ( .B1(n15050), .B2(n19095), .A(n14981), .ZN(P2_U2863) );
  NOR2_X1 U18229 ( .A1(n14983), .A2(n14984), .ZN(n14985) );
  OR2_X1 U18230 ( .A1(n14982), .A2(n14985), .ZN(n15082) );
  INV_X1 U18231 ( .A(n15141), .ZN(n14989) );
  NAND2_X1 U18232 ( .A1(n14987), .A2(n14986), .ZN(n14988) );
  NAND2_X1 U18233 ( .A1(n14989), .A2(n14988), .ZN(n18891) );
  MUX2_X1 U18234 ( .A(n10894), .B(n18891), .S(n19103), .Z(n14990) );
  OAI21_X1 U18235 ( .B1(n15082), .B2(n19095), .A(n14990), .ZN(P2_U2866) );
  INV_X1 U18236 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n14993) );
  AOI22_X1 U18237 ( .A1(n19109), .A2(n19121), .B1(n19170), .B2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n14992) );
  NAND2_X1 U18238 ( .A1(n19110), .A2(BUF1_REG_30__SCAN_IN), .ZN(n14991) );
  OAI211_X1 U18239 ( .C1(n15086), .C2(n14993), .A(n14992), .B(n14991), .ZN(
        n14994) );
  AOI21_X1 U18240 ( .B1(n14995), .B2(n19171), .A(n14994), .ZN(n14996) );
  OAI21_X1 U18241 ( .B1(n14997), .B2(n19145), .A(n14996), .ZN(P2_U2889) );
  NAND3_X1 U18242 ( .A1(n14999), .A2(n19175), .A3(n14998), .ZN(n15005) );
  OAI22_X1 U18243 ( .A1(n15084), .A2(n19124), .B1(n19169), .B2(n15000), .ZN(
        n15003) );
  INV_X1 U18244 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n15001) );
  NOR2_X1 U18245 ( .A1(n15086), .A2(n15001), .ZN(n15002) );
  AOI211_X1 U18246 ( .C1(BUF1_REG_29__SCAN_IN), .C2(n19110), .A(n15003), .B(
        n15002), .ZN(n15004) );
  OAI211_X1 U18247 ( .C1(n16086), .C2(n19153), .A(n15005), .B(n15004), .ZN(
        P2_U2890) );
  INV_X1 U18248 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n15007) );
  AOI22_X1 U18249 ( .A1(n19109), .A2(n19126), .B1(n19170), .B2(
        P2_EAX_REG_28__SCAN_IN), .ZN(n15006) );
  OAI21_X1 U18250 ( .B1(n15086), .B2(n15007), .A(n15006), .ZN(n15011) );
  INV_X1 U18251 ( .A(n11412), .ZN(n15008) );
  NOR2_X1 U18252 ( .A1(n16097), .A2(n19153), .ZN(n15010) );
  OAI21_X1 U18253 ( .B1(n15013), .B2(n19145), .A(n15012), .ZN(P2_U2891) );
  AOI21_X1 U18254 ( .B1(n15015), .B2(n9722), .A(n15014), .ZN(n16110) );
  INV_X1 U18255 ( .A(n16110), .ZN(n15023) );
  NAND2_X1 U18256 ( .A1(n15016), .A2(n19175), .ZN(n15022) );
  OAI22_X1 U18257 ( .A1(n15084), .A2(n19129), .B1(n19169), .B2(n15017), .ZN(
        n15020) );
  INV_X1 U18258 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n15018) );
  NOR2_X1 U18259 ( .A1(n15086), .A2(n15018), .ZN(n15019) );
  AOI211_X1 U18260 ( .C1(BUF1_REG_27__SCAN_IN), .C2(n19110), .A(n15020), .B(
        n15019), .ZN(n15021) );
  OAI211_X1 U18261 ( .C1(n15023), .C2(n19153), .A(n15022), .B(n15021), .ZN(
        P2_U2892) );
  NAND2_X1 U18262 ( .A1(n15037), .A2(n15024), .ZN(n15025) );
  NAND2_X1 U18263 ( .A1(n9722), .A2(n15025), .ZN(n16119) );
  NAND2_X1 U18264 ( .A1(n15026), .A2(n19175), .ZN(n15031) );
  INV_X1 U18265 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n15028) );
  AOI22_X1 U18266 ( .A1(n19109), .A2(n19132), .B1(n19170), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15027) );
  OAI21_X1 U18267 ( .B1(n15086), .B2(n15028), .A(n15027), .ZN(n15029) );
  AOI21_X1 U18268 ( .B1(n19110), .B2(BUF1_REG_26__SCAN_IN), .A(n15029), .ZN(
        n15030) );
  OAI211_X1 U18269 ( .C1(n16119), .C2(n19153), .A(n15031), .B(n15030), .ZN(
        P2_U2893) );
  NAND2_X1 U18270 ( .A1(n19111), .A2(BUF2_REG_25__SCAN_IN), .ZN(n15034) );
  AOI22_X1 U18271 ( .A1(n19109), .A2(n15032), .B1(n19170), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15033) );
  NAND2_X1 U18272 ( .A1(n15034), .A2(n15033), .ZN(n15039) );
  OR2_X1 U18273 ( .A1(n15045), .A2(n15035), .ZN(n15036) );
  NAND2_X1 U18274 ( .A1(n15037), .A2(n15036), .ZN(n16132) );
  NOR2_X1 U18275 ( .A1(n16132), .A2(n19153), .ZN(n15038) );
  AOI211_X1 U18276 ( .C1(n19110), .C2(BUF1_REG_25__SCAN_IN), .A(n15039), .B(
        n15038), .ZN(n15040) );
  OAI21_X1 U18277 ( .B1(n19145), .B2(n15041), .A(n15040), .ZN(P2_U2894) );
  NAND2_X1 U18278 ( .A1(n19111), .A2(BUF2_REG_24__SCAN_IN), .ZN(n15043) );
  AOI22_X1 U18279 ( .A1(n19109), .A2(n19138), .B1(n19170), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n15042) );
  NAND2_X1 U18280 ( .A1(n15043), .A2(n15042), .ZN(n15048) );
  AND2_X1 U18281 ( .A1(n15054), .A2(n15044), .ZN(n15046) );
  OR2_X1 U18282 ( .A1(n15046), .A2(n15045), .ZN(n16143) );
  NOR2_X1 U18283 ( .A1(n16143), .A2(n19153), .ZN(n15047) );
  AOI211_X1 U18284 ( .C1(n19110), .C2(BUF1_REG_24__SCAN_IN), .A(n15048), .B(
        n15047), .ZN(n15049) );
  OAI21_X1 U18285 ( .B1(n15050), .B2(n19145), .A(n15049), .ZN(P2_U2895) );
  NAND2_X1 U18286 ( .A1(n15052), .A2(n15051), .ZN(n15053) );
  NAND2_X1 U18287 ( .A1(n15054), .A2(n15053), .ZN(n16153) );
  AOI21_X1 U18288 ( .B1(n15055), .B2(n15057), .A(n15056), .ZN(n16164) );
  NAND2_X1 U18289 ( .A1(n16164), .A2(n19175), .ZN(n15063) );
  OAI22_X1 U18290 ( .A1(n15084), .A2(n19259), .B1(n15058), .B2(n19169), .ZN(
        n15061) );
  INV_X1 U18291 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n15059) );
  NOR2_X1 U18292 ( .A1(n15086), .A2(n15059), .ZN(n15060) );
  AOI211_X1 U18293 ( .C1(BUF1_REG_23__SCAN_IN), .C2(n19110), .A(n15061), .B(
        n15060), .ZN(n15062) );
  OAI211_X1 U18294 ( .C1(n16153), .C2(n19153), .A(n15063), .B(n15062), .ZN(
        P2_U2896) );
  OAI21_X1 U18295 ( .B1(n14982), .B2(n15065), .A(n15064), .ZN(n16167) );
  XNOR2_X1 U18296 ( .A(n15066), .B(n15067), .ZN(n15607) );
  INV_X1 U18297 ( .A(n15607), .ZN(n15068) );
  NAND2_X1 U18298 ( .A1(n15068), .A2(n19171), .ZN(n15074) );
  OAI22_X1 U18299 ( .A1(n15084), .A2(n19252), .B1(n19169), .B2(n15069), .ZN(
        n15072) );
  INV_X1 U18300 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n15070) );
  NOR2_X1 U18301 ( .A1(n15086), .A2(n15070), .ZN(n15071) );
  AOI211_X1 U18302 ( .C1(BUF1_REG_22__SCAN_IN), .C2(n19110), .A(n15072), .B(
        n15071), .ZN(n15073) );
  OAI211_X1 U18303 ( .C1(n19145), .C2(n16167), .A(n15074), .B(n15073), .ZN(
        P2_U2897) );
  OAI21_X1 U18304 ( .B1(n14629), .B2(n15075), .A(n15066), .ZN(n15327) );
  INV_X1 U18305 ( .A(n15327), .ZN(n18895) );
  NAND2_X1 U18306 ( .A1(n18895), .A2(n19171), .ZN(n15081) );
  OAI22_X1 U18307 ( .A1(n15084), .A2(n19143), .B1(n15076), .B2(n19169), .ZN(
        n15079) );
  INV_X1 U18308 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15077) );
  NOR2_X1 U18309 ( .A1(n15086), .A2(n15077), .ZN(n15078) );
  AOI211_X1 U18310 ( .C1(BUF1_REG_21__SCAN_IN), .C2(n19110), .A(n15079), .B(
        n15078), .ZN(n15080) );
  OAI211_X1 U18311 ( .C1(n19145), .C2(n15082), .A(n15081), .B(n15080), .ZN(
        P2_U2898) );
  NAND2_X1 U18312 ( .A1(n15358), .A2(n19171), .ZN(n15090) );
  OAI22_X1 U18313 ( .A1(n15084), .A2(n19240), .B1(n15083), .B2(n19169), .ZN(
        n15088) );
  INV_X1 U18314 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15085) );
  NOR2_X1 U18315 ( .A1(n15086), .A2(n15085), .ZN(n15087) );
  AOI211_X1 U18316 ( .C1(BUF1_REG_19__SCAN_IN), .C2(n19110), .A(n15088), .B(
        n15087), .ZN(n15089) );
  OAI211_X1 U18317 ( .C1(n19145), .C2(n15091), .A(n15090), .B(n15089), .ZN(
        P2_U2900) );
  INV_X1 U18318 ( .A(n11393), .ZN(n15094) );
  INV_X1 U18319 ( .A(n15092), .ZN(n15093) );
  OAI21_X1 U18320 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n15094), .A(
        n15093), .ZN(n15266) );
  NAND2_X1 U18321 ( .A1(n16268), .A2(n15095), .ZN(n15096) );
  INV_X1 U18322 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19801) );
  OR2_X1 U18323 ( .A1(n19046), .A2(n19801), .ZN(n15256) );
  OAI211_X1 U18324 ( .C1(n20923), .C2(n16278), .A(n15096), .B(n15256), .ZN(
        n15097) );
  AOI21_X1 U18325 ( .B1(n16109), .B2(n19225), .A(n15097), .ZN(n15100) );
  NAND3_X1 U18326 ( .A1(n15263), .A2(n11389), .A3(n15262), .ZN(n15099) );
  OAI211_X1 U18327 ( .C1(n15266), .C2(n19219), .A(n15100), .B(n15099), .ZN(
        P2_U2987) );
  NAND2_X1 U18328 ( .A1(n15102), .A2(n15101), .ZN(n15103) );
  XNOR2_X1 U18329 ( .A(n11396), .B(n15103), .ZN(n15289) );
  AOI21_X1 U18330 ( .B1(n21079), .B2(n15104), .A(n11394), .ZN(n15287) );
  NOR2_X1 U18331 ( .A1(n19046), .A2(n19797), .ZN(n15280) );
  NOR2_X1 U18332 ( .A1(n16278), .A2(n15105), .ZN(n15106) );
  AOI211_X1 U18333 ( .C1(n15107), .C2(n16268), .A(n15280), .B(n15106), .ZN(
        n15108) );
  OAI21_X1 U18334 ( .B1(n16131), .B2(n16273), .A(n15108), .ZN(n15109) );
  AOI21_X1 U18335 ( .B1(n15287), .B2(n16269), .A(n15109), .ZN(n15110) );
  OAI21_X1 U18336 ( .B1(n19221), .B2(n15289), .A(n15110), .ZN(P2_U2989) );
  INV_X1 U18337 ( .A(n15111), .ZN(n15112) );
  NOR2_X1 U18338 ( .A1(n15113), .A2(n15112), .ZN(n15114) );
  XNOR2_X1 U18339 ( .A(n15115), .B(n15114), .ZN(n15303) );
  INV_X1 U18340 ( .A(n16147), .ZN(n15116) );
  NAND2_X1 U18341 ( .A1(n16268), .A2(n15116), .ZN(n15118) );
  INV_X1 U18342 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n15117) );
  OR2_X1 U18343 ( .A1(n19046), .A2(n15117), .ZN(n15291) );
  OAI211_X1 U18344 ( .C1(n10012), .C2(n16278), .A(n15118), .B(n15291), .ZN(
        n15120) );
  INV_X1 U18345 ( .A(n15135), .ZN(n15122) );
  OAI21_X1 U18346 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15122), .A(
        n9872), .ZN(n15316) );
  NAND2_X1 U18347 ( .A1(n15143), .A2(n15123), .ZN(n15124) );
  NAND2_X1 U18348 ( .A1(n15125), .A2(n15124), .ZN(n16166) );
  INV_X1 U18349 ( .A(n16166), .ZN(n15133) );
  NAND2_X1 U18350 ( .A1(n16268), .A2(n15126), .ZN(n15127) );
  INV_X1 U18351 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19794) );
  OR2_X1 U18352 ( .A1(n19046), .A2(n19794), .ZN(n15309) );
  OAI211_X1 U18353 ( .C1(n15128), .C2(n16278), .A(n15127), .B(n15309), .ZN(
        n15132) );
  NOR2_X1 U18354 ( .A1(n15130), .A2(n15129), .ZN(n15304) );
  NOR3_X1 U18355 ( .A1(n15304), .A2(n9719), .A3(n19221), .ZN(n15131) );
  AOI211_X1 U18356 ( .C1(n19225), .C2(n15133), .A(n15132), .B(n15131), .ZN(
        n15134) );
  OAI21_X1 U18357 ( .B1(n19219), .B2(n15316), .A(n15134), .ZN(P2_U2991) );
  OAI21_X1 U18358 ( .B1(n9694), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15135), .ZN(n15326) );
  NAND2_X1 U18359 ( .A1(n15138), .A2(n15137), .ZN(n15139) );
  XNOR2_X1 U18360 ( .A(n15136), .B(n15139), .ZN(n15324) );
  OR2_X1 U18361 ( .A1(n15141), .A2(n15140), .ZN(n15142) );
  NAND2_X1 U18362 ( .A1(n15143), .A2(n15142), .ZN(n15606) );
  INV_X1 U18363 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19792) );
  NOR2_X1 U18364 ( .A1(n19046), .A2(n19792), .ZN(n15317) );
  NOR2_X1 U18365 ( .A1(n19229), .A2(n15610), .ZN(n15144) );
  AOI211_X1 U18366 ( .C1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n19218), .A(
        n15317), .B(n15144), .ZN(n15145) );
  OAI21_X1 U18367 ( .B1(n16273), .B2(n15606), .A(n15145), .ZN(n15146) );
  AOI21_X1 U18368 ( .B1(n15324), .B2(n11389), .A(n15146), .ZN(n15147) );
  OAI21_X1 U18369 ( .B1(n15326), .B2(n19219), .A(n15147), .ZN(P2_U2992) );
  AND2_X1 U18370 ( .A1(n16206), .A2(n16205), .ZN(n15379) );
  OAI21_X1 U18371 ( .B1(n15379), .B2(n15150), .A(n15381), .ZN(n15217) );
  INV_X1 U18372 ( .A(n15218), .ZN(n15151) );
  AOI21_X1 U18373 ( .B1(n15334), .B2(n15157), .A(n9694), .ZN(n15337) );
  NOR2_X1 U18374 ( .A1(n19046), .A2(n19790), .ZN(n15329) );
  NOR2_X1 U18375 ( .A1(n16278), .A2(n18890), .ZN(n15158) );
  AOI211_X1 U18376 ( .C1(n15159), .C2(n16268), .A(n15329), .B(n15158), .ZN(
        n15160) );
  OAI21_X1 U18377 ( .B1(n18891), .B2(n16273), .A(n15160), .ZN(n15161) );
  AOI21_X1 U18378 ( .B1(n15337), .B2(n16269), .A(n15161), .ZN(n15162) );
  OAI21_X1 U18379 ( .B1(n15339), .B2(n19221), .A(n15162), .ZN(P2_U2993) );
  NAND2_X1 U18380 ( .A1(n15164), .A2(n15163), .ZN(n15168) );
  NAND2_X1 U18381 ( .A1(n15166), .A2(n15165), .ZN(n15167) );
  XNOR2_X1 U18382 ( .A(n15168), .B(n15167), .ZN(n15351) );
  OR2_X1 U18383 ( .A1(n15179), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15169) );
  AND2_X1 U18384 ( .A1(n15157), .A2(n15169), .ZN(n15349) );
  NOR2_X1 U18385 ( .A1(n16174), .A2(n16273), .ZN(n15173) );
  OR2_X1 U18386 ( .A1(n19046), .A2(n19789), .ZN(n15341) );
  NAND2_X1 U18387 ( .A1(n19218), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15170) );
  OAI211_X1 U18388 ( .C1(n19229), .C2(n15171), .A(n15341), .B(n15170), .ZN(
        n15172) );
  AOI211_X1 U18389 ( .C1(n15349), .C2(n16269), .A(n15173), .B(n15172), .ZN(
        n15174) );
  OAI21_X1 U18390 ( .B1(n15351), .B2(n19221), .A(n15174), .ZN(P2_U2994) );
  NAND2_X1 U18391 ( .A1(n15176), .A2(n15175), .ZN(n15177) );
  AOI21_X1 U18392 ( .B1(n15343), .B2(n15178), .A(n15179), .ZN(n15359) );
  NAND2_X1 U18393 ( .A1(n15180), .A2(n16268), .ZN(n15182) );
  NOR2_X1 U18394 ( .A1(n19046), .A2(n19787), .ZN(n15352) );
  AOI21_X1 U18395 ( .B1(n19218), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n15352), .ZN(n15181) );
  OAI211_X1 U18396 ( .C1(n16273), .C2(n15183), .A(n15182), .B(n15181), .ZN(
        n15184) );
  AOI21_X1 U18397 ( .B1(n15359), .B2(n16269), .A(n15184), .ZN(n15185) );
  OAI21_X1 U18398 ( .B1(n15362), .B2(n19221), .A(n15185), .ZN(P2_U2995) );
  NAND2_X1 U18399 ( .A1(n15187), .A2(n15186), .ZN(n15188) );
  XNOR2_X1 U18400 ( .A(n15189), .B(n15188), .ZN(n15376) );
  INV_X1 U18401 ( .A(n15178), .ZN(n15191) );
  AOI21_X1 U18402 ( .B1(n15369), .B2(n15190), .A(n15191), .ZN(n15374) );
  INV_X1 U18403 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n15192) );
  NOR2_X1 U18404 ( .A1(n19046), .A2(n15192), .ZN(n15367) );
  OR2_X1 U18405 ( .A1(n15194), .A2(n15193), .ZN(n15195) );
  NAND2_X1 U18406 ( .A1(n15196), .A2(n15195), .ZN(n18903) );
  NOR2_X1 U18407 ( .A1(n16273), .A2(n18903), .ZN(n15197) );
  AOI211_X1 U18408 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n19218), .A(
        n15367), .B(n15197), .ZN(n15198) );
  OAI21_X1 U18409 ( .B1(n19229), .B2(n18898), .A(n15198), .ZN(n15199) );
  AOI21_X1 U18410 ( .B1(n15374), .B2(n16269), .A(n15199), .ZN(n15200) );
  OAI21_X1 U18411 ( .B1(n15376), .B2(n19221), .A(n15200), .ZN(P2_U2996) );
  INV_X1 U18412 ( .A(n15201), .ZN(n15203) );
  NAND2_X1 U18413 ( .A1(n15203), .A2(n15202), .ZN(n15207) );
  NAND2_X1 U18414 ( .A1(n15205), .A2(n15204), .ZN(n15206) );
  XNOR2_X1 U18415 ( .A(n15207), .B(n15206), .ZN(n15623) );
  INV_X1 U18416 ( .A(n15623), .ZN(n15216) );
  OR2_X1 U18417 ( .A1(n19046), .A2(n19784), .ZN(n15619) );
  OAI21_X1 U18418 ( .B1(n16278), .B2(n10008), .A(n15619), .ZN(n15209) );
  NOR2_X1 U18419 ( .A1(n16273), .A2(n15620), .ZN(n15208) );
  AOI211_X1 U18420 ( .C1(n16268), .C2(n15210), .A(n15209), .B(n15208), .ZN(
        n15215) );
  INV_X1 U18421 ( .A(n15594), .ZN(n15213) );
  OAI211_X1 U18422 ( .C1(n15213), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16269), .B(n15190), .ZN(n15214) );
  OAI211_X1 U18423 ( .C1(n15216), .C2(n19221), .A(n15215), .B(n15214), .ZN(
        P2_U2997) );
  XOR2_X1 U18424 ( .A(n15218), .B(n15217), .Z(n15593) );
  OAI211_X1 U18425 ( .C1(n15377), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n16269), .B(n15594), .ZN(n15227) );
  NAND2_X1 U18426 ( .A1(n15221), .A2(n15220), .ZN(n15222) );
  NAND2_X1 U18427 ( .A1(n15223), .A2(n15222), .ZN(n19082) );
  NAND2_X1 U18428 ( .A1(n19217), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15601) );
  NAND2_X1 U18429 ( .A1(n19218), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15224) );
  OAI211_X1 U18430 ( .C1(n16273), .C2(n19082), .A(n15601), .B(n15224), .ZN(
        n15225) );
  AOI21_X1 U18431 ( .B1(n16268), .B2(n18920), .A(n15225), .ZN(n15226) );
  OAI211_X1 U18432 ( .C1(n19221), .C2(n15593), .A(n15227), .B(n15226), .ZN(
        P2_U2998) );
  INV_X1 U18433 ( .A(n15228), .ZN(n15434) );
  OR2_X1 U18434 ( .A1(n15228), .A2(n10651), .ZN(n16230) );
  OAI21_X1 U18435 ( .B1(n15434), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16230), .ZN(n15433) );
  NAND2_X1 U18436 ( .A1(n15230), .A2(n15229), .ZN(n15234) );
  INV_X1 U18437 ( .A(n15231), .ZN(n15436) );
  NOR2_X1 U18438 ( .A1(n15232), .A2(n15436), .ZN(n15233) );
  XOR2_X1 U18439 ( .A(n15234), .B(n15233), .Z(n15430) );
  INV_X1 U18440 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19770) );
  OAI22_X1 U18441 ( .A1(n19770), .A2(n19046), .B1(n19229), .B2(n18977), .ZN(
        n15241) );
  NAND2_X1 U18442 ( .A1(n15236), .A2(n15235), .ZN(n15237) );
  NAND2_X1 U18443 ( .A1(n15238), .A2(n15237), .ZN(n19090) );
  OAI22_X1 U18444 ( .A1(n16273), .A2(n19090), .B1(n16278), .B2(n15239), .ZN(
        n15240) );
  AOI211_X1 U18445 ( .C1(n15430), .C2(n11389), .A(n15241), .B(n15240), .ZN(
        n15242) );
  OAI21_X1 U18446 ( .B1(n15433), .B2(n19219), .A(n15242), .ZN(P2_U3004) );
  INV_X1 U18447 ( .A(n15259), .ZN(n15245) );
  NOR2_X1 U18448 ( .A1(n16098), .A2(n16327), .ZN(n15243) );
  INV_X1 U18449 ( .A(n15255), .ZN(n15248) );
  NAND3_X1 U18450 ( .A1(n15248), .A2(n15247), .A3(n15246), .ZN(n15249) );
  OAI211_X1 U18451 ( .C1(n16097), .C2(n16330), .A(n15250), .B(n15249), .ZN(
        n15251) );
  AOI21_X1 U18452 ( .B1(n15252), .B2(n16314), .A(n15251), .ZN(n15253) );
  OAI21_X1 U18453 ( .B1(n15254), .B2(n16326), .A(n15253), .ZN(P2_U3018) );
  NOR2_X1 U18454 ( .A1(n15255), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15261) );
  NAND2_X1 U18455 ( .A1(n16109), .A2(n16316), .ZN(n15257) );
  OAI211_X1 U18456 ( .C1(n15259), .C2(n15258), .A(n15257), .B(n15256), .ZN(
        n15260) );
  AOI211_X1 U18457 ( .C1(n16110), .C2(n16312), .A(n15261), .B(n15260), .ZN(
        n15265) );
  NAND3_X1 U18458 ( .A1(n15263), .A2(n16317), .A3(n15262), .ZN(n15264) );
  OAI211_X1 U18459 ( .C1(n15266), .C2(n16339), .A(n15265), .B(n15264), .ZN(
        P2_U3019) );
  INV_X1 U18460 ( .A(n15267), .ZN(n15276) );
  INV_X1 U18461 ( .A(n15268), .ZN(n15269) );
  OAI21_X1 U18462 ( .B1(n15284), .B2(n15270), .A(n15269), .ZN(n15271) );
  AOI21_X1 U18463 ( .B1(n16120), .B2(n16316), .A(n15271), .ZN(n15274) );
  XNOR2_X1 U18464 ( .A(n21079), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15272) );
  NAND2_X1 U18465 ( .A1(n15279), .A2(n15272), .ZN(n15273) );
  OAI211_X1 U18466 ( .C1(n16119), .C2(n16330), .A(n15274), .B(n15273), .ZN(
        n15275) );
  OAI21_X1 U18467 ( .B1(n16326), .B2(n15278), .A(n15277), .ZN(P2_U3020) );
  NOR2_X1 U18468 ( .A1(n16132), .A2(n16330), .ZN(n15286) );
  NAND2_X1 U18469 ( .A1(n15279), .A2(n21079), .ZN(n15283) );
  INV_X1 U18470 ( .A(n16131), .ZN(n15281) );
  AOI21_X1 U18471 ( .B1(n15281), .B2(n16316), .A(n15280), .ZN(n15282) );
  OAI211_X1 U18472 ( .C1(n15284), .C2(n21079), .A(n15283), .B(n15282), .ZN(
        n15285) );
  AOI211_X1 U18473 ( .C1(n15287), .C2(n16314), .A(n15286), .B(n15285), .ZN(
        n15288) );
  OAI21_X1 U18474 ( .B1(n16326), .B2(n15289), .A(n15288), .ZN(P2_U3021) );
  INV_X1 U18475 ( .A(n15290), .ZN(n15301) );
  INV_X1 U18476 ( .A(n15291), .ZN(n15294) );
  NOR2_X1 U18477 ( .A1(n15292), .A2(n15297), .ZN(n15293) );
  AOI211_X1 U18478 ( .C1(n15295), .C2(n16316), .A(n15294), .B(n15293), .ZN(
        n15299) );
  INV_X1 U18479 ( .A(n15296), .ZN(n15321) );
  NAND3_X1 U18480 ( .A1(n15321), .A2(n15305), .A3(n15297), .ZN(n15298) );
  OAI211_X1 U18481 ( .C1(n16143), .C2(n16330), .A(n15299), .B(n15298), .ZN(
        n15300) );
  AOI21_X1 U18482 ( .B1(n15301), .B2(n16314), .A(n15300), .ZN(n15302) );
  OAI21_X1 U18483 ( .B1(n15303), .B2(n16326), .A(n15302), .ZN(P2_U3022) );
  NOR3_X1 U18484 ( .A1(n15304), .A2(n9719), .A3(n16326), .ZN(n15314) );
  AOI21_X1 U18485 ( .B1(n15320), .B2(n15307), .A(n15305), .ZN(n15311) );
  NAND2_X1 U18486 ( .A1(n15426), .A2(n15306), .ZN(n15333) );
  OR2_X1 U18487 ( .A1(n15333), .A2(n15307), .ZN(n15308) );
  OAI211_X1 U18488 ( .C1(n16166), .C2(n16327), .A(n15309), .B(n15308), .ZN(
        n15310) );
  AOI21_X1 U18489 ( .B1(n15321), .B2(n15311), .A(n15310), .ZN(n15312) );
  OAI21_X1 U18490 ( .B1(n16153), .B2(n16330), .A(n15312), .ZN(n15313) );
  NOR2_X1 U18491 ( .A1(n15314), .A2(n15313), .ZN(n15315) );
  OAI21_X1 U18492 ( .B1(n15316), .B2(n16339), .A(n15315), .ZN(P2_U3023) );
  INV_X1 U18493 ( .A(n15606), .ZN(n16168) );
  AOI21_X1 U18494 ( .B1(n16168), .B2(n16316), .A(n15317), .ZN(n15318) );
  OAI21_X1 U18495 ( .B1(n15320), .B2(n15333), .A(n15318), .ZN(n15319) );
  AOI21_X1 U18496 ( .B1(n15321), .B2(n15320), .A(n15319), .ZN(n15322) );
  OAI21_X1 U18497 ( .B1(n15607), .B2(n16330), .A(n15322), .ZN(n15323) );
  AOI21_X1 U18498 ( .B1(n15324), .B2(n16317), .A(n15323), .ZN(n15325) );
  OAI21_X1 U18499 ( .B1(n15326), .B2(n16339), .A(n15325), .ZN(P2_U3024) );
  NOR2_X1 U18500 ( .A1(n15327), .A2(n16330), .ZN(n15336) );
  INV_X1 U18501 ( .A(n15356), .ZN(n15328) );
  NAND3_X1 U18502 ( .A1(n15328), .A2(n15342), .A3(n15334), .ZN(n15332) );
  INV_X1 U18503 ( .A(n18891), .ZN(n15330) );
  AOI21_X1 U18504 ( .B1(n15330), .B2(n16316), .A(n15329), .ZN(n15331) );
  OAI211_X1 U18505 ( .C1(n15334), .C2(n15333), .A(n15332), .B(n15331), .ZN(
        n15335) );
  AOI211_X1 U18506 ( .C1(n15337), .C2(n16314), .A(n15336), .B(n15335), .ZN(
        n15338) );
  OAI21_X1 U18507 ( .B1(n15339), .B2(n16326), .A(n15338), .ZN(P2_U3025) );
  OAI21_X1 U18508 ( .B1(n15401), .B2(n15340), .A(n15400), .ZN(n15368) );
  OAI21_X1 U18509 ( .B1(n16174), .B2(n16327), .A(n15341), .ZN(n15346) );
  AOI211_X1 U18510 ( .C1(n15344), .C2(n15343), .A(n15342), .B(n15356), .ZN(
        n15345) );
  AOI211_X1 U18511 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15368), .A(
        n15346), .B(n15345), .ZN(n15347) );
  OAI21_X1 U18512 ( .B1(n16186), .B2(n16330), .A(n15347), .ZN(n15348) );
  AOI21_X1 U18513 ( .B1(n15349), .B2(n16314), .A(n15348), .ZN(n15350) );
  OAI21_X1 U18514 ( .B1(n15351), .B2(n16326), .A(n15350), .ZN(P2_U3026) );
  AOI21_X1 U18515 ( .B1(n15353), .B2(n16316), .A(n15352), .ZN(n15355) );
  NAND2_X1 U18516 ( .A1(n15368), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15354) );
  OAI211_X1 U18517 ( .C1(n15356), .C2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n15355), .B(n15354), .ZN(n15357) );
  AOI21_X1 U18518 ( .B1(n15358), .B2(n16312), .A(n15357), .ZN(n15361) );
  NAND2_X1 U18519 ( .A1(n15359), .A2(n16314), .ZN(n15360) );
  OAI211_X1 U18520 ( .C1(n15362), .C2(n16326), .A(n15361), .B(n15360), .ZN(
        P2_U3027) );
  NAND2_X1 U18521 ( .A1(n13807), .A2(n15363), .ZN(n15364) );
  NAND2_X1 U18522 ( .A1(n15365), .A2(n15364), .ZN(n18904) );
  NOR2_X1 U18523 ( .A1(n16327), .A2(n18903), .ZN(n15366) );
  AOI211_X1 U18524 ( .C1(n15368), .C2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15367), .B(n15366), .ZN(n15372) );
  NAND3_X1 U18525 ( .A1(n15444), .A2(n15370), .A3(n15369), .ZN(n15371) );
  OAI211_X1 U18526 ( .C1(n18904), .C2(n16330), .A(n15372), .B(n15371), .ZN(
        n15373) );
  AOI21_X1 U18527 ( .B1(n15374), .B2(n16314), .A(n15373), .ZN(n15375) );
  OAI21_X1 U18528 ( .B1(n15376), .B2(n16326), .A(n15375), .ZN(P2_U3028) );
  INV_X1 U18529 ( .A(n16197), .ZN(n15394) );
  INV_X1 U18530 ( .A(n16204), .ZN(n15378) );
  OR2_X1 U18531 ( .A1(n15379), .A2(n15378), .ZN(n15383) );
  NAND2_X1 U18532 ( .A1(n15381), .A2(n15380), .ZN(n15382) );
  XNOR2_X1 U18533 ( .A(n15383), .B(n15382), .ZN(n16199) );
  XNOR2_X1 U18534 ( .A(n16279), .B(n15384), .ZN(n19119) );
  INV_X1 U18535 ( .A(n18924), .ZN(n16198) );
  NAND2_X1 U18536 ( .A1(n15402), .A2(n15444), .ZN(n16282) );
  INV_X1 U18537 ( .A(n16282), .ZN(n15414) );
  NAND2_X1 U18538 ( .A1(n15385), .A2(n15414), .ZN(n15600) );
  INV_X1 U18539 ( .A(n15386), .ZN(n15387) );
  INV_X1 U18540 ( .A(n15400), .ZN(n15443) );
  AOI21_X1 U18541 ( .B1(n15387), .B2(n16334), .A(n15443), .ZN(n15596) );
  NAND2_X1 U18542 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19217), .ZN(n15388) );
  OAI221_X1 U18543 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15600), 
        .C1(n15389), .C2(n15596), .A(n15388), .ZN(n15390) );
  AOI21_X1 U18544 ( .B1(n16198), .B2(n16316), .A(n15390), .ZN(n15391) );
  OAI21_X1 U18545 ( .B1(n19119), .B2(n16330), .A(n15391), .ZN(n15392) );
  AOI21_X1 U18546 ( .B1(n16199), .B2(n16317), .A(n15392), .ZN(n15393) );
  OAI21_X1 U18547 ( .B1(n15394), .B2(n16339), .A(n15393), .ZN(P2_U3031) );
  NAND2_X1 U18548 ( .A1(n15396), .A2(n15395), .ZN(n15397) );
  NAND2_X1 U18549 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15410), .ZN(
        n15409) );
  NOR2_X1 U18550 ( .A1(n16283), .A2(n16231), .ZN(n16203) );
  AOI21_X1 U18551 ( .B1(n10689), .B2(n15409), .A(n16203), .ZN(n16213) );
  NAND2_X1 U18552 ( .A1(n16213), .A2(n16314), .ZN(n15408) );
  OAI21_X1 U18553 ( .B1(n15399), .B2(n15398), .A(n16281), .ZN(n19125) );
  INV_X1 U18554 ( .A(n19125), .ZN(n15406) );
  OAI21_X1 U18555 ( .B1(n15402), .B2(n15401), .A(n15400), .ZN(n15413) );
  AOI21_X1 U18556 ( .B1(n15414), .B2(n16283), .A(n15413), .ZN(n16284) );
  AOI21_X1 U18557 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15414), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15404) );
  AOI22_X1 U18558 ( .A1(n16316), .A2(n18945), .B1(n19217), .B2(
        P2_REIP_REG_13__SCAN_IN), .ZN(n15403) );
  OAI21_X1 U18559 ( .B1(n16284), .B2(n15404), .A(n15403), .ZN(n15405) );
  AOI21_X1 U18560 ( .B1(n15406), .B2(n16312), .A(n15405), .ZN(n15407) );
  OAI211_X1 U18561 ( .C1(n16211), .C2(n16326), .A(n15408), .B(n15407), .ZN(
        P2_U3033) );
  OAI21_X1 U18562 ( .B1(n15410), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15409), .ZN(n16219) );
  XNOR2_X1 U18563 ( .A(n16296), .B(n15411), .ZN(n19128) );
  INV_X1 U18564 ( .A(n19128), .ZN(n15423) );
  INV_X1 U18565 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19774) );
  NOR2_X1 U18566 ( .A1(n19774), .A2(n19046), .ZN(n15412) );
  AOI221_X1 U18567 ( .B1(n15414), .B2(n10665), .C1(n15413), .C2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n15412), .ZN(n15415) );
  OAI21_X1 U18568 ( .B1(n16327), .B2(n16217), .A(n15415), .ZN(n15422) );
  INV_X1 U18569 ( .A(n15416), .ZN(n15417) );
  NOR2_X1 U18570 ( .A1(n15418), .A2(n15417), .ZN(n15419) );
  XNOR2_X1 U18571 ( .A(n15420), .B(n15419), .ZN(n16218) );
  NOR2_X1 U18572 ( .A1(n16218), .A2(n16326), .ZN(n15421) );
  AOI211_X1 U18573 ( .C1(n16312), .C2(n15423), .A(n15422), .B(n15421), .ZN(
        n15424) );
  OAI21_X1 U18574 ( .B1(n16339), .B2(n16219), .A(n15424), .ZN(P2_U3034) );
  AOI21_X1 U18575 ( .B1(n15440), .B2(n15425), .A(n16298), .ZN(n19131) );
  NOR2_X1 U18576 ( .A1(n16327), .A2(n19090), .ZN(n15429) );
  NAND2_X1 U18577 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15444), .ZN(
        n16294) );
  OAI21_X1 U18578 ( .B1(n15443), .B2(n21061), .A(n15426), .ZN(n16299) );
  NAND2_X1 U18579 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19217), .ZN(n15427) );
  OAI221_X1 U18580 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16294), 
        .C1(n10651), .C2(n16299), .A(n15427), .ZN(n15428) );
  AOI211_X1 U18581 ( .C1(n19131), .C2(n16312), .A(n15429), .B(n15428), .ZN(
        n15432) );
  NAND2_X1 U18582 ( .A1(n15430), .A2(n16317), .ZN(n15431) );
  OAI211_X1 U18583 ( .C1(n15433), .C2(n16339), .A(n15432), .B(n15431), .ZN(
        P2_U3036) );
  AOI21_X1 U18584 ( .B1(n15435), .B2(n21061), .A(n15434), .ZN(n16238) );
  INV_X1 U18585 ( .A(n16238), .ZN(n15449) );
  NOR2_X1 U18586 ( .A1(n15437), .A2(n15436), .ZN(n15438) );
  XNOR2_X1 U18587 ( .A(n15439), .B(n15438), .ZN(n16237) );
  OAI21_X1 U18588 ( .B1(n16309), .B2(n15441), .A(n15440), .ZN(n19136) );
  INV_X1 U18589 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19768) );
  NOR2_X1 U18590 ( .A1(n19768), .A2(n19046), .ZN(n15442) );
  AOI221_X1 U18591 ( .B1(n15444), .B2(n21061), .C1(n15443), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15442), .ZN(n15446) );
  NAND2_X1 U18592 ( .A1(n16316), .A2(n16236), .ZN(n15445) );
  OAI211_X1 U18593 ( .C1(n19136), .C2(n16330), .A(n15446), .B(n15445), .ZN(
        n15447) );
  AOI21_X1 U18594 ( .B1(n16237), .B2(n16317), .A(n15447), .ZN(n15448) );
  OAI21_X1 U18595 ( .B1(n15449), .B2(n16339), .A(n15448), .ZN(P2_U3037) );
  INV_X1 U18596 ( .A(n15467), .ZN(n16343) );
  INV_X1 U18597 ( .A(n15450), .ZN(n19055) );
  AOI22_X1 U18598 ( .A1(n19041), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19055), .B2(n9690), .ZN(n15458) );
  INV_X1 U18599 ( .A(n15458), .ZN(n15451) );
  OAI222_X1 U18600 ( .A1(n16343), .A2(n15453), .B1(n19820), .B2(n15452), .C1(
        n15457), .C2(n15451), .ZN(n15454) );
  MUX2_X1 U18601 ( .A(n15454), .B(n9661), .S(n15470), .Z(P2_U3601) );
  OAI21_X1 U18602 ( .B1(n9690), .B2(n15456), .A(n15455), .ZN(n15466) );
  INV_X1 U18603 ( .A(n15466), .ZN(n15459) );
  NOR2_X1 U18604 ( .A1(n15458), .A2(n15457), .ZN(n15465) );
  AOI222_X1 U18605 ( .A1(n15460), .A2(n15463), .B1(n15467), .B2(n19842), .C1(
        n15459), .C2(n15465), .ZN(n15462) );
  NAND2_X1 U18606 ( .A1(n15470), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15461) );
  OAI21_X1 U18607 ( .B1(n15462), .B2(n15470), .A(n15461), .ZN(P2_U3600) );
  AOI222_X1 U18608 ( .A1(n15468), .A2(n15467), .B1(n15466), .B2(n15465), .C1(
        n15464), .C2(n15463), .ZN(n15471) );
  NAND2_X1 U18609 ( .A1(n15470), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15469) );
  OAI21_X1 U18610 ( .B1(n15471), .B2(n15470), .A(n15469), .ZN(P2_U3599) );
  NAND3_X1 U18611 ( .A1(n18219), .A2(n18204), .A3(n15472), .ZN(n15473) );
  INV_X1 U18612 ( .A(n17211), .ZN(n17224) );
  NAND2_X1 U18613 ( .A1(n18219), .A2(n17224), .ZN(n17218) );
  INV_X1 U18614 ( .A(n17218), .ZN(n17220) );
  NAND2_X1 U18615 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16955) );
  NOR2_X2 U18616 ( .A1(n17211), .A2(n18219), .ZN(n17221) );
  INV_X1 U18617 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16620) );
  INV_X1 U18618 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16639) );
  INV_X1 U18619 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16661) );
  INV_X1 U18620 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n16723) );
  INV_X1 U18621 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17106) );
  INV_X1 U18622 ( .A(P3_EBX_REG_2__SCAN_IN), .ZN(n17212) );
  NAND2_X1 U18623 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17210) );
  NOR2_X1 U18624 ( .A1(n17212), .A2(n17210), .ZN(n17199) );
  NAND3_X1 U18625 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17199), .ZN(n17201) );
  NAND4_X1 U18626 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(P3_EBX_REG_6__SCAN_IN), .A4(P3_EBX_REG_5__SCAN_IN), .ZN(n15476) );
  NAND4_X1 U18627 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(P3_EBX_REG_10__SCAN_IN), .A4(P3_EBX_REG_7__SCAN_IN), .ZN(n15475)
         );
  NOR3_X1 U18628 ( .A1(n17201), .A2(n15476), .A3(n15475), .ZN(n15554) );
  NAND2_X1 U18629 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n15554), .ZN(n17102) );
  NAND2_X1 U18630 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(n17090), .ZN(n17089) );
  NAND2_X1 U18631 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17022), .ZN(n17009) );
  NAND2_X1 U18632 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16983), .ZN(n16977) );
  NAND2_X1 U18633 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16982), .ZN(n16968) );
  NAND2_X1 U18634 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16973), .ZN(n16964) );
  AOI22_X1 U18635 ( .A1(n17220), .A2(n16955), .B1(n17214), .B2(n16964), .ZN(
        n16954) );
  INV_X1 U18636 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16585) );
  AOI22_X1 U18637 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11524), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15480) );
  AOI22_X1 U18638 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15479) );
  AOI22_X1 U18639 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15478) );
  AOI22_X1 U18640 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15477) );
  NAND4_X1 U18641 ( .A1(n15480), .A2(n15479), .A3(n15478), .A4(n15477), .ZN(
        n15486) );
  AOI22_X1 U18642 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15484) );
  AOI22_X1 U18643 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15483) );
  AOI22_X1 U18644 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15482) );
  AOI22_X1 U18645 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n9653), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15481) );
  NAND4_X1 U18646 ( .A1(n15484), .A2(n15483), .A3(n15482), .A4(n15481), .ZN(
        n15485) );
  NOR2_X1 U18647 ( .A1(n15486), .A2(n15485), .ZN(n15551) );
  AOI22_X1 U18648 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n15490) );
  AOI22_X1 U18649 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15489) );
  AOI22_X1 U18650 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15488) );
  AOI22_X1 U18651 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15487) );
  NAND4_X1 U18652 ( .A1(n15490), .A2(n15489), .A3(n15488), .A4(n15487), .ZN(
        n15496) );
  AOI22_X1 U18653 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11524), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15494) );
  AOI22_X1 U18654 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15493) );
  AOI22_X1 U18655 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15492) );
  AOI22_X1 U18656 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n9667), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15491) );
  NAND4_X1 U18657 ( .A1(n15494), .A2(n15493), .A3(n15492), .A4(n15491), .ZN(
        n15495) );
  NOR2_X1 U18658 ( .A1(n15496), .A2(n15495), .ZN(n16965) );
  AOI22_X1 U18659 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17050), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n15500) );
  AOI22_X1 U18660 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17171), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15499) );
  AOI22_X1 U18661 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17124), .ZN(n15498) );
  AOI22_X1 U18662 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n9667), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n9655), .ZN(n15497) );
  NAND4_X1 U18663 ( .A1(n15500), .A2(n15499), .A3(n15498), .A4(n15497), .ZN(
        n15506) );
  AOI22_X1 U18664 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17160), .ZN(n15504) );
  AOI22_X1 U18665 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9652), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17149), .ZN(n15503) );
  AOI22_X1 U18666 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17176), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17055), .ZN(n15502) );
  AOI22_X1 U18667 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n9653), .ZN(n15501) );
  NAND4_X1 U18668 ( .A1(n15504), .A2(n15503), .A3(n15502), .A4(n15501), .ZN(
        n15505) );
  NOR2_X1 U18669 ( .A1(n15506), .A2(n15505), .ZN(n16974) );
  AOI22_X1 U18670 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15517) );
  AOI22_X1 U18671 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15516) );
  INV_X1 U18672 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15508) );
  AOI22_X1 U18673 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15507) );
  OAI21_X1 U18674 ( .B1(n9713), .B2(n15508), .A(n15507), .ZN(n15514) );
  AOI22_X1 U18675 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15512) );
  AOI22_X1 U18676 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15511) );
  AOI22_X1 U18677 ( .A1(n17159), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n15510) );
  AOI22_X1 U18678 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(n9655), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15509) );
  NAND4_X1 U18679 ( .A1(n15512), .A2(n15511), .A3(n15510), .A4(n15509), .ZN(
        n15513) );
  AOI211_X1 U18680 ( .C1(n17171), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n15514), .B(n15513), .ZN(n15515) );
  NAND3_X1 U18681 ( .A1(n15517), .A2(n15516), .A3(n15515), .ZN(n16979) );
  AOI22_X1 U18682 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15527) );
  AOI22_X1 U18683 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15526) );
  AOI22_X1 U18684 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15518) );
  OAI21_X1 U18685 ( .B1(n10155), .B2(n20953), .A(n15518), .ZN(n15524) );
  AOI22_X1 U18686 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n9653), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15522) );
  AOI22_X1 U18687 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n15521) );
  AOI22_X1 U18688 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11524), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15520) );
  AOI22_X1 U18689 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15519) );
  NAND4_X1 U18690 ( .A1(n15522), .A2(n15521), .A3(n15520), .A4(n15519), .ZN(
        n15523) );
  AOI211_X1 U18691 ( .C1(n17017), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n15524), .B(n15523), .ZN(n15525) );
  NAND3_X1 U18692 ( .A1(n15527), .A2(n15526), .A3(n15525), .ZN(n16980) );
  NAND2_X1 U18693 ( .A1(n16979), .A2(n16980), .ZN(n16978) );
  NOR2_X1 U18694 ( .A1(n16974), .A2(n16978), .ZN(n16971) );
  AOI22_X1 U18695 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n15539) );
  AOI22_X1 U18696 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15538) );
  AOI22_X1 U18697 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15528) );
  OAI21_X1 U18698 ( .B1(n15530), .B2(n15529), .A(n15528), .ZN(n15536) );
  AOI22_X1 U18699 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15534) );
  AOI22_X1 U18700 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n15533) );
  AOI22_X1 U18701 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15532) );
  AOI22_X1 U18702 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n9653), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15531) );
  NAND4_X1 U18703 ( .A1(n15534), .A2(n15533), .A3(n15532), .A4(n15531), .ZN(
        n15535) );
  AOI211_X1 U18704 ( .C1(n17017), .C2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A(
        n15536), .B(n15535), .ZN(n15537) );
  NAND3_X1 U18705 ( .A1(n15539), .A2(n15538), .A3(n15537), .ZN(n16970) );
  NAND2_X1 U18706 ( .A1(n16971), .A2(n16970), .ZN(n16969) );
  NOR2_X1 U18707 ( .A1(n16965), .A2(n16969), .ZN(n16962) );
  AOI22_X1 U18708 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n15550) );
  AOI22_X1 U18709 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15549) );
  INV_X1 U18710 ( .A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n21067) );
  AOI22_X1 U18711 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15540) );
  OAI21_X1 U18712 ( .B1(n15541), .B2(n21067), .A(n15540), .ZN(n15547) );
  AOI22_X1 U18713 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15545) );
  AOI22_X1 U18714 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15544) );
  AOI22_X1 U18715 ( .A1(n9652), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15543) );
  AOI22_X1 U18716 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15542) );
  NAND4_X1 U18717 ( .A1(n15545), .A2(n15544), .A3(n15543), .A4(n15542), .ZN(
        n15546) );
  AOI211_X1 U18718 ( .C1(n17154), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(
        n15547), .B(n15546), .ZN(n15548) );
  NAND3_X1 U18719 ( .A1(n15550), .A2(n15549), .A3(n15548), .ZN(n16961) );
  NAND2_X1 U18720 ( .A1(n16962), .A2(n16961), .ZN(n16960) );
  NOR2_X1 U18721 ( .A1(n15551), .A2(n16960), .ZN(n16953) );
  AOI21_X1 U18722 ( .B1(n15551), .B2(n16960), .A(n16953), .ZN(n17239) );
  INV_X1 U18723 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16598) );
  NOR3_X1 U18724 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16598), .A3(n16964), .ZN(
        n15552) );
  AOI21_X1 U18725 ( .B1(n17221), .B2(n17239), .A(n15552), .ZN(n15553) );
  OAI21_X1 U18726 ( .B1(n16954), .B2(n16585), .A(n15553), .ZN(P3_U2675) );
  INV_X1 U18727 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16756) );
  NAND2_X1 U18728 ( .A1(n17220), .A2(n16756), .ZN(n17105) );
  INV_X1 U18729 ( .A(n15554), .ZN(n15570) );
  AOI22_X1 U18730 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15568) );
  AOI22_X1 U18731 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15567) );
  INV_X1 U18732 ( .A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15556) );
  AOI22_X1 U18733 ( .A1(n17055), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15555) );
  OAI21_X1 U18734 ( .B1(n16938), .B2(n15556), .A(n15555), .ZN(n15565) );
  AOI22_X1 U18735 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15563) );
  AOI22_X1 U18736 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15562) );
  AOI22_X1 U18737 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15561) );
  AOI22_X1 U18738 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15560) );
  NAND4_X1 U18739 ( .A1(n15563), .A2(n15562), .A3(n15561), .A4(n15560), .ZN(
        n15564) );
  AOI211_X1 U18740 ( .C1(n17050), .C2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n15565), .B(n15564), .ZN(n15566) );
  NAND3_X1 U18741 ( .A1(n15568), .A2(n15567), .A3(n15566), .ZN(n17318) );
  INV_X1 U18742 ( .A(n17318), .ZN(n15569) );
  INV_X1 U18743 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17117) );
  INV_X1 U18744 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17146) );
  INV_X1 U18745 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16808) );
  INV_X1 U18746 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17184) );
  INV_X1 U18747 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17191) );
  NOR3_X1 U18748 ( .A1(n16853), .A2(n17211), .A3(n17201), .ZN(n17198) );
  NAND2_X1 U18749 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17198), .ZN(n17188) );
  NOR2_X1 U18750 ( .A1(n17191), .A2(n17188), .ZN(n17183) );
  INV_X1 U18751 ( .A(n17183), .ZN(n17185) );
  NOR3_X1 U18752 ( .A1(n16808), .A2(n17184), .A3(n17185), .ZN(n17145) );
  INV_X1 U18753 ( .A(n17145), .ZN(n17168) );
  NOR2_X1 U18754 ( .A1(n17146), .A2(n17168), .ZN(n17132) );
  NAND2_X1 U18755 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(n17132), .ZN(n17131) );
  OAI21_X1 U18756 ( .B1(n17117), .B2(n17131), .A(n17214), .ZN(n17118) );
  OAI222_X1 U18757 ( .A1(n17105), .A2(n15570), .B1(n17214), .B2(n15569), .C1(
        n16756), .C2(n17118), .ZN(P3_U2690) );
  NAND2_X1 U18758 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18401) );
  AOI221_X1 U18759 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18401), .C1(n15572), 
        .C2(n18401), .A(n15571), .ZN(n18182) );
  NOR2_X1 U18760 ( .A1(n15573), .A2(n18649), .ZN(n15574) );
  OAI21_X1 U18761 ( .B1(n15574), .B2(n18524), .A(n18183), .ZN(n18180) );
  AOI22_X1 U18762 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18182), .B1(
        n18180), .B2(n18670), .ZN(P3_U2865) );
  NOR2_X1 U18763 ( .A1(n15575), .A2(n17884), .ZN(n17890) );
  NAND2_X1 U18764 ( .A1(n17866), .A2(n17890), .ZN(n16414) );
  OAI21_X1 U18765 ( .B1(n16379), .B2(n15576), .A(n16414), .ZN(n15577) );
  INV_X1 U18766 ( .A(n15577), .ZN(n17863) );
  NOR2_X1 U18767 ( .A1(n17863), .A2(n18173), .ZN(n15694) );
  INV_X1 U18768 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16399) );
  NAND2_X1 U18769 ( .A1(n15694), .A2(n16399), .ZN(n15588) );
  INV_X1 U18770 ( .A(n15686), .ZN(n15579) );
  NAND2_X1 U18771 ( .A1(n17513), .A2(n17500), .ZN(n15685) );
  NOR2_X1 U18772 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17645), .ZN(
        n15578) );
  AOI21_X1 U18773 ( .B1(n15579), .B2(n15685), .A(n15578), .ZN(n15580) );
  XOR2_X1 U18774 ( .A(n15580), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n16402) );
  NOR2_X1 U18775 ( .A1(n16403), .A2(n16399), .ZN(n15687) );
  INV_X1 U18776 ( .A(n15687), .ZN(n16415) );
  NOR2_X1 U18777 ( .A1(n16415), .A2(n17499), .ZN(n16387) );
  NOR3_X1 U18778 ( .A1(n16387), .A2(n15581), .A3(n18166), .ZN(n15583) );
  NOR2_X1 U18779 ( .A1(n17498), .A2(n16415), .ZN(n16388) );
  NAND2_X1 U18780 ( .A1(n17923), .A2(n18158), .ZN(n18140) );
  NOR2_X1 U18781 ( .A1(n16388), .A2(n18140), .ZN(n15582) );
  NOR2_X1 U18782 ( .A1(n15583), .A2(n15582), .ZN(n15692) );
  NAND2_X1 U18783 ( .A1(n17990), .A2(n18158), .ZN(n18160) );
  INV_X1 U18784 ( .A(n18160), .ZN(n15691) );
  AOI22_X1 U18785 ( .A1(n15691), .A2(n17500), .B1(n18077), .B2(n15584), .ZN(
        n15585) );
  AOI21_X1 U18786 ( .B1(n15692), .B2(n15585), .A(n16399), .ZN(n15586) );
  AOI21_X1 U18787 ( .B1(n16402), .B2(n18093), .A(n15586), .ZN(n15587) );
  NAND2_X1 U18788 ( .A1(n9654), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16407) );
  OAI211_X1 U18789 ( .C1(n16403), .C2(n15588), .A(n15587), .B(n16407), .ZN(
        P3_U2833) );
  AND2_X1 U18790 ( .A1(n15590), .A2(n15589), .ZN(n15591) );
  OR2_X1 U18791 ( .A1(n15591), .A2(n13806), .ZN(n19113) );
  OAI22_X1 U18792 ( .A1(n19113), .A2(n16330), .B1(n16327), .B2(n19082), .ZN(
        n15592) );
  INV_X1 U18793 ( .A(n15592), .ZN(n15604) );
  INV_X1 U18794 ( .A(n15593), .ZN(n15599) );
  OAI21_X1 U18795 ( .B1(n16314), .B2(n15595), .A(n15594), .ZN(n15597) );
  OAI211_X1 U18796 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15598), .A(
        n15597), .B(n15596), .ZN(n15616) );
  AOI22_X1 U18797 ( .A1(n15599), .A2(n16317), .B1(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n15616), .ZN(n15603) );
  INV_X1 U18798 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15617) );
  OAI21_X1 U18799 ( .B1(n16339), .B2(n16202), .A(n15600), .ZN(n15615) );
  NAND3_X1 U18800 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n15617), .A3(
        n15615), .ZN(n15602) );
  NAND4_X1 U18801 ( .A1(n15604), .A2(n15603), .A3(n15602), .A4(n15601), .ZN(
        P2_U3030) );
  AOI22_X1 U18802 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19045), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19028), .ZN(n15614) );
  AOI22_X1 U18803 ( .A1(P2_EBX_REG_22__SCAN_IN), .A2(n19059), .B1(n15605), 
        .B2(n19057), .ZN(n15613) );
  OAI22_X1 U18804 ( .A1(n15607), .A2(n19049), .B1(n15606), .B2(n19011), .ZN(
        n15608) );
  INV_X1 U18805 ( .A(n15608), .ZN(n15612) );
  NAND4_X1 U18806 ( .A1(n15614), .A2(n15613), .A3(n15612), .A4(n15611), .ZN(
        P2_U2833) );
  NAND3_X1 U18807 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(n15615), .ZN(n15627) );
  AOI21_X1 U18808 ( .B1(n15617), .B2(n16334), .A(n15616), .ZN(n15625) );
  NOR2_X1 U18809 ( .A1(n15618), .A2(n16330), .ZN(n15622) );
  OAI21_X1 U18810 ( .B1(n16327), .B2(n15620), .A(n15619), .ZN(n15621) );
  AOI211_X1 U18811 ( .C1(n15623), .C2(n16317), .A(n15622), .B(n15621), .ZN(
        n15624) );
  OAI221_X1 U18812 ( .B1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n15627), 
        .C1(n15626), .C2(n15625), .A(n15624), .ZN(P2_U3029) );
  NAND2_X1 U18813 ( .A1(n15628), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15629) );
  NAND2_X1 U18814 ( .A1(n15629), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n15630) );
  OR2_X1 U18815 ( .A1(n15631), .A2(n15630), .ZN(n15636) );
  INV_X1 U18816 ( .A(n15636), .ZN(n15632) );
  OAI22_X1 U18817 ( .A1(n15634), .A2(n15633), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n15632), .ZN(n15635) );
  OAI21_X1 U18818 ( .B1(n15636), .B2(n20746), .A(n15635), .ZN(n15639) );
  INV_X1 U18819 ( .A(n15637), .ZN(n15638) );
  AOI222_X1 U18820 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n15639), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15638), .C1(n15639), 
        .C2(n15638), .ZN(n15640) );
  AOI222_X1 U18821 ( .A1(n20882), .A2(n15641), .B1(n20882), .B2(n15640), .C1(
        n15641), .C2(n15640), .ZN(n15647) );
  NOR2_X1 U18822 ( .A1(n15643), .A2(n15642), .ZN(n15646) );
  OAI21_X1 U18823 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15644), .ZN(n15645) );
  OAI211_X1 U18824 ( .C1(n15647), .C2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n15646), .B(n15645), .ZN(n15648) );
  NOR3_X1 U18825 ( .A1(n15650), .A2(n15649), .A3(n15648), .ZN(n15664) );
  NAND3_X1 U18826 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20814), .A3(n20804), 
        .ZN(n15651) );
  AOI22_X1 U18827 ( .A1(n15654), .A2(n15653), .B1(n15652), .B2(n15651), .ZN(
        n16078) );
  OAI221_X1 U18828 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n15664), 
        .A(n16078), .ZN(n16084) );
  NOR2_X1 U18829 ( .A1(n15656), .A2(n15655), .ZN(n15657) );
  NOR2_X1 U18830 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15657), .ZN(n15662) );
  AOI211_X1 U18831 ( .C1(n20814), .C2(n20383), .A(n15659), .B(n15658), .ZN(
        n15660) );
  NAND2_X1 U18832 ( .A1(n16084), .A2(n15660), .ZN(n15661) );
  AOI22_X1 U18833 ( .A1(n16084), .A2(n15662), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15661), .ZN(n15663) );
  OAI21_X1 U18834 ( .B1(n15664), .B2(n19871), .A(n15663), .ZN(P1_U3161) );
  OAI21_X1 U18835 ( .B1(n15674), .B2(n15666), .A(n15665), .ZN(n15667) );
  XNOR2_X1 U18836 ( .A(n15667), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15844) );
  AOI22_X1 U18837 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15951), .B1(
        n13376), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15684) );
  INV_X1 U18838 ( .A(n15668), .ZN(n20090) );
  NAND2_X1 U18839 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15669), .ZN(
        n15671) );
  OAI21_X1 U18840 ( .B1(n15985), .B2(n15671), .A(n15670), .ZN(n15989) );
  NAND3_X1 U18841 ( .A1(n15672), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n15989), .ZN(n15699) );
  OAI21_X1 U18842 ( .B1(n20090), .B2(n15673), .A(n15699), .ZN(n15966) );
  NAND2_X1 U18843 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15966), .ZN(
        n15705) );
  NOR2_X1 U18844 ( .A1(n15674), .A2(n15705), .ZN(n15957) );
  INV_X1 U18845 ( .A(n15675), .ZN(n15678) );
  AOI21_X1 U18846 ( .B1(n15678), .B2(n15677), .A(n15676), .ZN(n15680) );
  OR2_X1 U18847 ( .A1(n15680), .A2(n15679), .ZN(n15820) );
  INV_X1 U18848 ( .A(n15820), .ZN(n15681) );
  AOI22_X1 U18849 ( .A1(n15957), .A2(n15682), .B1(n15681), .B2(n16062), .ZN(
        n15683) );
  OAI211_X1 U18850 ( .C1(n15844), .C2(n16008), .A(n15684), .B(n15683), .ZN(
        P1_U3010) );
  NAND2_X1 U18851 ( .A1(n15687), .A2(n15686), .ZN(n16359) );
  OAI21_X1 U18852 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15688), .A(
        n16358), .ZN(n16391) );
  NOR2_X1 U18853 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16415), .ZN(
        n16386) );
  OAI21_X1 U18854 ( .B1(n15689), .B2(n18173), .A(n18159), .ZN(n15690) );
  AOI21_X1 U18855 ( .B1(n15691), .B2(n16415), .A(n15690), .ZN(n16410) );
  INV_X1 U18856 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16416) );
  AOI21_X1 U18857 ( .B1(n16410), .B2(n15692), .A(n16416), .ZN(n15693) );
  AOI21_X1 U18858 ( .B1(n16386), .B2(n15694), .A(n15693), .ZN(n15695) );
  NAND2_X1 U18859 ( .A1(n9654), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16383) );
  OAI211_X1 U18860 ( .C1(n18070), .C2(n16391), .A(n15695), .B(n16383), .ZN(
        P3_U2832) );
  INV_X1 U18861 ( .A(HOLD), .ZN(n20809) );
  INV_X1 U18862 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20824) );
  NAND2_X1 U18863 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20824), .ZN(n20813) );
  INV_X1 U18864 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20815) );
  NOR2_X1 U18865 ( .A1(n20808), .A2(n20815), .ZN(n15696) );
  AND2_X1 U18866 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20814), .ZN(n20819) );
  AOI221_X1 U18867 ( .B1(n20809), .B2(n15696), .C1(n20824), .C2(n15696), .A(
        n20819), .ZN(n15698) );
  OAI211_X1 U18868 ( .C1(n20809), .C2(n20813), .A(n15698), .B(n15697), .ZN(
        P1_U3195) );
  INV_X1 U18869 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16513) );
  NOR2_X1 U18870 ( .A1(n20028), .A2(n16513), .ZN(P1_U2905) );
  OAI221_X1 U18871 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n20090), 
        .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15699), .A(n15964), .ZN(
        n15700) );
  AOI22_X1 U18872 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15700), .B1(
        n13376), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n15704) );
  INV_X1 U18873 ( .A(n15767), .ZN(n15701) );
  AOI22_X1 U18874 ( .A1(n15702), .A2(n20087), .B1(n16018), .B2(n15701), .ZN(
        n15703) );
  OAI211_X1 U18875 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15705), .A(
        n15704), .B(n15703), .ZN(P1_U3011) );
  NAND2_X1 U18876 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15706), .ZN(n15708) );
  AOI21_X1 U18877 ( .B1(n19838), .B2(n16342), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15707) );
  AOI21_X1 U18878 ( .B1(n15708), .B2(n15707), .A(n15709), .ZN(P2_U3178) );
  AOI221_X1 U18879 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n15709), .C1(n19859), .C2(
        n15709), .A(n19679), .ZN(n19853) );
  INV_X1 U18880 ( .A(n19853), .ZN(n19854) );
  NOR2_X1 U18881 ( .A1(n15710), .A2(n19854), .ZN(P2_U3047) );
  NOR2_X1 U18882 ( .A1(n18840), .A2(n16540), .ZN(n15711) );
  NOR2_X1 U18883 ( .A1(n17311), .A2(n17369), .ZN(n17372) );
  INV_X1 U18884 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17437) );
  INV_X1 U18885 ( .A(n17369), .ZN(n15717) );
  NAND2_X1 U18886 ( .A1(n15714), .A2(n15717), .ZN(n17368) );
  AOI22_X1 U18887 ( .A1(n17370), .A2(BUF2_REG_0__SCAN_IN), .B1(n17345), .B2(
        n15715), .ZN(n15716) );
  OAI221_X1 U18888 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17361), .C1(n17437), 
        .C2(n15717), .A(n15716), .ZN(P3_U2735) );
  AOI22_X1 U18889 ( .A1(n19932), .A2(P1_EBX_REG_25__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19978), .ZN(n15724) );
  INV_X1 U18890 ( .A(n15830), .ZN(n15720) );
  AND2_X1 U18891 ( .A1(n19961), .A2(n15718), .ZN(n15719) );
  INV_X1 U18892 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n15931) );
  AOI22_X1 U18893 ( .A1(n15720), .A2(n19979), .B1(n15719), .B2(n15931), .ZN(
        n15723) );
  AOI22_X1 U18894 ( .A1(n15827), .A2(n19916), .B1(n19940), .B2(n15937), .ZN(
        n15722) );
  NOR2_X1 U18895 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n19965), .ZN(n15734) );
  AOI21_X1 U18896 ( .B1(n15727), .B2(n19961), .A(n19960), .ZN(n15745) );
  INV_X1 U18897 ( .A(n15745), .ZN(n15725) );
  OAI21_X1 U18898 ( .B1(n15734), .B2(n15725), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n15721) );
  NAND4_X1 U18899 ( .A1(n15724), .A2(n15723), .A3(n15722), .A4(n15721), .ZN(
        P1_U2815) );
  AOI22_X1 U18900 ( .A1(n15726), .A2(n19979), .B1(P1_REIP_REG_24__SCAN_IN), 
        .B2(n15725), .ZN(n15737) );
  INV_X1 U18901 ( .A(n15727), .ZN(n15735) );
  OAI22_X1 U18902 ( .A1(n19987), .A2(n15729), .B1(n19898), .B2(n15728), .ZN(
        n15733) );
  OAI22_X1 U18903 ( .A1(n15731), .A2(n19923), .B1(n15730), .B2(n19985), .ZN(
        n15732) );
  AOI211_X1 U18904 ( .C1(n15735), .C2(n15734), .A(n15733), .B(n15732), .ZN(
        n15736) );
  NAND2_X1 U18905 ( .A1(n15737), .A2(n15736), .ZN(P1_U2816) );
  AND2_X1 U18906 ( .A1(n19961), .A2(n15738), .ZN(n15746) );
  AOI21_X1 U18907 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n15746), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n15744) );
  INV_X1 U18908 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15739) );
  OAI22_X1 U18909 ( .A1(n15739), .A2(n19898), .B1(n19935), .B2(n15843), .ZN(
        n15740) );
  AOI21_X1 U18910 ( .B1(n19932), .B2(P1_EBX_REG_23__SCAN_IN), .A(n15740), .ZN(
        n15743) );
  OAI22_X1 U18911 ( .A1(n15839), .A2(n19923), .B1(n19985), .B2(n15945), .ZN(
        n15741) );
  INV_X1 U18912 ( .A(n15741), .ZN(n15742) );
  OAI211_X1 U18913 ( .C1(n15745), .C2(n15744), .A(n15743), .B(n15742), .ZN(
        P1_U2817) );
  AOI22_X1 U18914 ( .A1(n19932), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19978), .ZN(n15755) );
  AOI22_X1 U18915 ( .A1(n15747), .A2(n19979), .B1(n15746), .B2(n14463), .ZN(
        n15754) );
  NOR2_X1 U18916 ( .A1(n15953), .A2(n19985), .ZN(n15748) );
  AOI21_X1 U18917 ( .B1(n15749), .B2(n19916), .A(n15748), .ZN(n15753) );
  NOR2_X1 U18918 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n19965), .ZN(n15759) );
  OAI21_X1 U18919 ( .B1(n19960), .B2(n15756), .A(n15750), .ZN(n15768) );
  INV_X1 U18920 ( .A(n15768), .ZN(n15751) );
  OAI21_X1 U18921 ( .B1(n15759), .B2(n15751), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15752) );
  NAND4_X1 U18922 ( .A1(n15755), .A2(n15754), .A3(n15753), .A4(n15752), .ZN(
        P1_U2818) );
  INV_X1 U18923 ( .A(n15756), .ZN(n15760) );
  OAI22_X1 U18924 ( .A1(n15768), .A2(n20849), .B1(n15845), .B2(n19935), .ZN(
        n15758) );
  INV_X1 U18925 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15851) );
  OAI22_X1 U18926 ( .A1(n19987), .A2(n15823), .B1(n15851), .B2(n19898), .ZN(
        n15757) );
  AOI211_X1 U18927 ( .C1(n15760), .C2(n15759), .A(n15758), .B(n15757), .ZN(
        n15763) );
  NOR2_X1 U18928 ( .A1(n15820), .A2(n19985), .ZN(n15761) );
  AOI21_X1 U18929 ( .B1(n15846), .B2(n19916), .A(n15761), .ZN(n15762) );
  NAND2_X1 U18930 ( .A1(n15763), .A2(n15762), .ZN(P1_U2819) );
  AOI22_X1 U18931 ( .A1(n19932), .A2(P1_EBX_REG_20__SCAN_IN), .B1(n19979), 
        .B2(n15764), .ZN(n15773) );
  INV_X1 U18932 ( .A(n15765), .ZN(n15771) );
  NOR2_X1 U18933 ( .A1(n15766), .A2(n15798), .ZN(n15775) );
  AOI21_X1 U18934 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(n15775), .A(
        P1_REIP_REG_20__SCAN_IN), .ZN(n15769) );
  OAI22_X1 U18935 ( .A1(n15769), .A2(n15768), .B1(n15767), .B2(n19985), .ZN(
        n15770) );
  AOI21_X1 U18936 ( .B1(n15771), .B2(n19916), .A(n15770), .ZN(n15772) );
  OAI211_X1 U18937 ( .C1(n15774), .C2(n19898), .A(n15773), .B(n15772), .ZN(
        P1_U2820) );
  INV_X1 U18938 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n20847) );
  AOI22_X1 U18939 ( .A1(n15775), .A2(n20847), .B1(n19932), .B2(
        P1_EBX_REG_19__SCAN_IN), .ZN(n15776) );
  OAI21_X1 U18940 ( .B1(n15860), .B2(n19935), .A(n15776), .ZN(n15777) );
  AOI211_X1 U18941 ( .C1(n19978), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n19946), .B(n15777), .ZN(n15783) );
  NOR2_X1 U18942 ( .A1(n15961), .A2(n19985), .ZN(n15778) );
  AOI21_X1 U18943 ( .B1(n15857), .B2(n19916), .A(n15778), .ZN(n15782) );
  OAI21_X1 U18944 ( .B1(n15780), .B2(n15779), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15781) );
  NAND3_X1 U18945 ( .A1(n15783), .A2(n15782), .A3(n15781), .ZN(P1_U2821) );
  INV_X1 U18946 ( .A(n15798), .ZN(n15785) );
  OAI211_X1 U18947 ( .C1(P1_REIP_REG_16__SCAN_IN), .C2(P1_REIP_REG_15__SCAN_IN), .A(n15785), .B(n15784), .ZN(n15786) );
  INV_X1 U18948 ( .A(n19946), .ZN(n19921) );
  OAI211_X1 U18949 ( .C1(n15787), .C2(n19987), .A(n15786), .B(n19921), .ZN(
        n15791) );
  OAI22_X1 U18950 ( .A1(n15789), .A2(n19923), .B1(n19985), .B2(n15788), .ZN(
        n15790) );
  AOI211_X1 U18951 ( .C1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n19978), .A(
        n15791), .B(n15790), .ZN(n15794) );
  NAND2_X1 U18952 ( .A1(n15792), .A2(n19979), .ZN(n15793) );
  OAI211_X1 U18953 ( .C1(n15802), .C2(n15795), .A(n15794), .B(n15793), .ZN(
        P1_U2824) );
  AOI22_X1 U18954 ( .A1(n19940), .A2(n15979), .B1(n19979), .B2(n15878), .ZN(
        n15801) );
  NOR2_X1 U18955 ( .A1(n19898), .A2(n20934), .ZN(n15796) );
  AOI211_X1 U18956 ( .C1(n19932), .C2(P1_EBX_REG_15__SCAN_IN), .A(n19946), .B(
        n15796), .ZN(n15797) );
  OAI21_X1 U18957 ( .B1(n15798), .B2(P1_REIP_REG_15__SCAN_IN), .A(n15797), 
        .ZN(n15799) );
  AOI21_X1 U18958 ( .B1(n15879), .B2(n19916), .A(n15799), .ZN(n15800) );
  OAI211_X1 U18959 ( .C1(n15803), .C2(n15802), .A(n15801), .B(n15800), .ZN(
        P1_U2825) );
  NAND2_X1 U18960 ( .A1(n19940), .A2(n9783), .ZN(n15804) );
  OAI211_X1 U18961 ( .C1(n15805), .C2(n19898), .A(n15804), .B(n19921), .ZN(
        n15806) );
  AOI21_X1 U18962 ( .B1(n19932), .B2(P1_EBX_REG_12__SCAN_IN), .A(n15806), .ZN(
        n15811) );
  OAI21_X1 U18963 ( .B1(n19965), .B2(n15807), .A(n20839), .ZN(n15808) );
  AOI22_X1 U18964 ( .A1(n15888), .A2(n19979), .B1(n15809), .B2(n15808), .ZN(
        n15810) );
  OAI211_X1 U18965 ( .C1(n19923), .C2(n15886), .A(n15811), .B(n15810), .ZN(
        P1_U2828) );
  NOR4_X1 U18966 ( .A1(n19965), .A2(P1_REIP_REG_11__SCAN_IN), .A3(n19895), 
        .A4(n15812), .ZN(n15816) );
  NAND2_X1 U18967 ( .A1(n19940), .A2(n16010), .ZN(n15814) );
  AOI21_X1 U18968 ( .B1(n19978), .B2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n19946), .ZN(n15813) );
  OAI211_X1 U18969 ( .C1(n19935), .C2(n15899), .A(n15814), .B(n15813), .ZN(
        n15815) );
  AOI211_X1 U18970 ( .C1(P1_EBX_REG_11__SCAN_IN), .C2(n19932), .A(n15816), .B(
        n15815), .ZN(n15819) );
  AOI22_X1 U18971 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15817), .B1(n19916), 
        .B2(n15896), .ZN(n15818) );
  NAND2_X1 U18972 ( .A1(n15819), .A2(n15818), .ZN(P1_U2829) );
  NOR2_X1 U18973 ( .A1(n15820), .A2(n20005), .ZN(n15821) );
  AOI21_X1 U18974 ( .B1(n15846), .B2(n12640), .A(n15821), .ZN(n15822) );
  OAI21_X1 U18975 ( .B1(n20016), .B2(n15823), .A(n15822), .ZN(P1_U2851) );
  AOI22_X1 U18976 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(
        n13376), .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n15829) );
  MUX2_X1 U18977 ( .A(n15855), .B(n15824), .S(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .Z(n15825) );
  OAI211_X1 U18978 ( .C1(n15835), .C2(n15831), .A(n15825), .B(n15836), .ZN(
        n15826) );
  XNOR2_X1 U18979 ( .A(n15826), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15934) );
  AOI22_X1 U18980 ( .A1(n15827), .A2(n15909), .B1(n20074), .B2(n15934), .ZN(
        n15828) );
  OAI211_X1 U18981 ( .C1(n15914), .C2(n15830), .A(n15829), .B(n15828), .ZN(
        P1_U2974) );
  AOI22_X1 U18982 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(
        n13376), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n15842) );
  MUX2_X1 U18983 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n15835), .S(
        n13705), .Z(n15834) );
  NAND2_X1 U18984 ( .A1(n15831), .A2(n15835), .ZN(n15833) );
  MUX2_X1 U18985 ( .A(n15834), .B(n15833), .S(n15832), .Z(n15838) );
  OR2_X1 U18986 ( .A1(n15836), .A2(n15835), .ZN(n15837) );
  OAI22_X1 U18987 ( .A1(n15839), .A2(n20101), .B1(n15944), .B2(n19877), .ZN(
        n15840) );
  INV_X1 U18988 ( .A(n15840), .ZN(n15841) );
  OAI211_X1 U18989 ( .C1(n15914), .C2(n15843), .A(n15842), .B(n15841), .ZN(
        P1_U2976) );
  INV_X1 U18990 ( .A(n15844), .ZN(n15848) );
  INV_X1 U18991 ( .A(n15845), .ZN(n15847) );
  AOI222_X1 U18992 ( .A1(n15848), .A2(n20074), .B1(n15847), .B2(n15889), .C1(
        n15909), .C2(n15846), .ZN(n15850) );
  NAND2_X1 U18993 ( .A1(n13376), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15849) );
  OAI211_X1 U18994 ( .C1(n15851), .C2(n15918), .A(n15850), .B(n15849), .ZN(
        P1_U2978) );
  AOI22_X1 U18995 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n13376), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15859) );
  NAND2_X1 U18996 ( .A1(n9834), .A2(n15852), .ZN(n15854) );
  MUX2_X1 U18997 ( .A(n15855), .B(n15854), .S(n15853), .Z(n15856) );
  XNOR2_X1 U18998 ( .A(n15856), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15963) );
  AOI22_X1 U18999 ( .A1(n15857), .A2(n15909), .B1(n20074), .B2(n15963), .ZN(
        n15858) );
  OAI211_X1 U19000 ( .C1(n15914), .C2(n15860), .A(n15859), .B(n15858), .ZN(
        P1_U2980) );
  OAI21_X1 U19001 ( .B1(n15892), .B2(n15862), .A(n15861), .ZN(n15865) );
  NAND2_X1 U19002 ( .A1(n15865), .A2(n15863), .ZN(n15864) );
  MUX2_X1 U19003 ( .A(n15865), .B(n15864), .S(n9834), .Z(n15866) );
  XNOR2_X1 U19004 ( .A(n15866), .B(n15969), .ZN(n15978) );
  AOI22_X1 U19005 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n13376), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15870) );
  AOI22_X1 U19006 ( .A1(n15868), .A2(n15909), .B1(n15889), .B2(n15867), .ZN(
        n15869) );
  OAI211_X1 U19007 ( .C1(n19877), .C2(n15978), .A(n15870), .B(n15869), .ZN(
        P1_U2982) );
  INV_X1 U19008 ( .A(n15871), .ZN(n15872) );
  NOR2_X1 U19009 ( .A1(n15873), .A2(n15872), .ZN(n15877) );
  NAND2_X1 U19010 ( .A1(n15875), .A2(n15874), .ZN(n15876) );
  XNOR2_X1 U19011 ( .A(n15877), .B(n15876), .ZN(n15984) );
  AOI22_X1 U19012 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n13376), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15881) );
  AOI22_X1 U19013 ( .A1(n15879), .A2(n15909), .B1(n15889), .B2(n15878), .ZN(
        n15880) );
  OAI211_X1 U19014 ( .C1(n15984), .C2(n19877), .A(n15881), .B(n15880), .ZN(
        P1_U2984) );
  OAI21_X1 U19015 ( .B1(n15884), .B2(n15883), .A(n15882), .ZN(n15885) );
  INV_X1 U19016 ( .A(n15885), .ZN(n16009) );
  AOI22_X1 U19017 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13376), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15891) );
  INV_X1 U19018 ( .A(n15886), .ZN(n15887) );
  AOI22_X1 U19019 ( .A1(n15889), .A2(n15888), .B1(n15909), .B2(n15887), .ZN(
        n15890) );
  OAI211_X1 U19020 ( .C1(n16009), .C2(n19877), .A(n15891), .B(n15890), .ZN(
        P1_U2987) );
  AOI22_X1 U19021 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n13376), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15898) );
  NAND3_X1 U19022 ( .A1(n15892), .A2(n13705), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15894) );
  NAND2_X1 U19023 ( .A1(n15894), .A2(n15893), .ZN(n15895) );
  XOR2_X1 U19024 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n15895), .Z(
        n16011) );
  AOI22_X1 U19025 ( .A1(n20074), .A2(n16011), .B1(n15909), .B2(n15896), .ZN(
        n15897) );
  OAI211_X1 U19026 ( .C1(n15914), .C2(n15899), .A(n15898), .B(n15897), .ZN(
        P1_U2988) );
  AOI22_X1 U19027 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n13376), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15904) );
  XNOR2_X1 U19028 ( .A(n15900), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15901) );
  XNOR2_X1 U19029 ( .A(n15902), .B(n15901), .ZN(n16046) );
  AOI22_X1 U19030 ( .A1(n16046), .A2(n20074), .B1(n15909), .B2(n19997), .ZN(
        n15903) );
  OAI211_X1 U19031 ( .C1(n15914), .C2(n19909), .A(n15904), .B(n15903), .ZN(
        P1_U2992) );
  AOI22_X1 U19032 ( .A1(n20076), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n13376), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15911) );
  NAND2_X1 U19033 ( .A1(n15906), .A2(n15905), .ZN(n15907) );
  XNOR2_X1 U19034 ( .A(n15908), .B(n15907), .ZN(n16052) );
  AOI22_X1 U19035 ( .A1(n16052), .A2(n20074), .B1(n15909), .B2(n20001), .ZN(
        n15910) );
  OAI211_X1 U19036 ( .C1(n15914), .C2(n19922), .A(n15911), .B(n15910), .ZN(
        P1_U2993) );
  INV_X1 U19037 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n15919) );
  XOR2_X1 U19038 ( .A(n15913), .B(n15912), .Z(n16067) );
  OAI22_X1 U19039 ( .A1(n20006), .A2(n20101), .B1(n19936), .B2(n15914), .ZN(
        n15915) );
  AOI21_X1 U19040 ( .B1(n16067), .B2(n20074), .A(n15915), .ZN(n15917) );
  INV_X1 U19041 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n19944) );
  NOR2_X1 U19042 ( .A1(n15996), .A2(n19944), .ZN(n16061) );
  INV_X1 U19043 ( .A(n16061), .ZN(n15916) );
  OAI211_X1 U19044 ( .C1(n15919), .C2(n15918), .A(n15917), .B(n15916), .ZN(
        P1_U2994) );
  INV_X1 U19045 ( .A(n15920), .ZN(n15923) );
  INV_X1 U19046 ( .A(n15921), .ZN(n15922) );
  AOI22_X1 U19047 ( .A1(n15923), .A2(n20087), .B1(n16018), .B2(n15922), .ZN(
        n15930) );
  INV_X1 U19048 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n15924) );
  NOR2_X1 U19049 ( .A1(n15996), .A2(n15924), .ZN(n15925) );
  AOI221_X1 U19050 ( .B1(n15928), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), 
        .C1(n15927), .C2(n15926), .A(n15925), .ZN(n15929) );
  NAND2_X1 U19051 ( .A1(n15930), .A2(n15929), .ZN(P1_U3004) );
  NOR2_X1 U19052 ( .A1(n15996), .A2(n15931), .ZN(n15932) );
  AOI211_X1 U19053 ( .C1(n20087), .C2(n15934), .A(n15933), .B(n15932), .ZN(
        n15941) );
  INV_X1 U19054 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15935) );
  OR2_X1 U19055 ( .A1(n15936), .A2(n15935), .ZN(n15939) );
  NAND2_X1 U19056 ( .A1(n15937), .A2(n16062), .ZN(n15938) );
  AND2_X1 U19057 ( .A1(n15939), .A2(n15938), .ZN(n15940) );
  NAND2_X1 U19058 ( .A1(n15941), .A2(n15940), .ZN(P1_U3006) );
  INV_X1 U19059 ( .A(n15942), .ZN(n15943) );
  AOI22_X1 U19060 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n13376), .B1(n15943), 
        .B2(n15835), .ZN(n15949) );
  INV_X1 U19061 ( .A(n15944), .ZN(n15947) );
  INV_X1 U19062 ( .A(n15945), .ZN(n15946) );
  AOI22_X1 U19063 ( .A1(n15947), .A2(n20087), .B1(n16062), .B2(n15946), .ZN(
        n15948) );
  OAI211_X1 U19064 ( .C1(n15950), .C2(n15835), .A(n15949), .B(n15948), .ZN(
        P1_U3008) );
  AOI22_X1 U19065 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n15951), .B1(
        n13376), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15960) );
  INV_X1 U19066 ( .A(n15952), .ZN(n15955) );
  INV_X1 U19067 ( .A(n15953), .ZN(n15954) );
  AOI22_X1 U19068 ( .A1(n15955), .A2(n20087), .B1(n16018), .B2(n15954), .ZN(
        n15959) );
  OAI211_X1 U19069 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15957), .B(n15956), .ZN(
        n15958) );
  NAND3_X1 U19070 ( .A1(n15960), .A2(n15959), .A3(n15958), .ZN(P1_U3009) );
  INV_X1 U19071 ( .A(n15961), .ZN(n15962) );
  AOI22_X1 U19072 ( .A1(n15963), .A2(n20087), .B1(n16018), .B2(n15962), .ZN(
        n15968) );
  NAND2_X1 U19073 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15964), .ZN(
        n15965) );
  OAI21_X1 U19074 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15966), .A(
        n15965), .ZN(n15967) );
  OAI211_X1 U19075 ( .C1(n20847), .C2(n15996), .A(n15968), .B(n15967), .ZN(
        P1_U3012) );
  NAND3_X1 U19076 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15970) );
  OAI21_X1 U19077 ( .B1(n15971), .B2(n15970), .A(n15969), .ZN(n15975) );
  INV_X1 U19078 ( .A(n15972), .ZN(n15973) );
  AOI22_X1 U19079 ( .A1(n15975), .A2(n15974), .B1(n16018), .B2(n15973), .ZN(
        n15977) );
  NAND2_X1 U19080 ( .A1(n13376), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15976) );
  OAI211_X1 U19081 ( .C1(n15978), .C2(n16008), .A(n15977), .B(n15976), .ZN(
        P1_U3014) );
  AOI22_X1 U19082 ( .A1(n15979), .A2(n16062), .B1(n13376), .B2(
        P1_REIP_REG_15__SCAN_IN), .ZN(n15983) );
  AOI21_X1 U19083 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15981), .A(
        n15980), .ZN(n15982) );
  OAI211_X1 U19084 ( .C1(n15984), .C2(n16008), .A(n15983), .B(n15982), .ZN(
        P1_U3016) );
  NOR3_X1 U19085 ( .A1(n20090), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        n15985), .ZN(n15988) );
  OAI22_X1 U19086 ( .A1(n20084), .A2(n15986), .B1(n14498), .B2(n15996), .ZN(
        n15987) );
  NOR2_X1 U19087 ( .A1(n15988), .A2(n15987), .ZN(n15992) );
  AOI22_X1 U19088 ( .A1(n15990), .A2(n20087), .B1(n15989), .B2(n15993), .ZN(
        n15991) );
  OAI211_X1 U19089 ( .C1(n15994), .C2(n15993), .A(n15992), .B(n15991), .ZN(
        P1_U3018) );
  INV_X1 U19090 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16004) );
  NAND3_X1 U19091 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16021), .ZN(n16015) );
  NOR3_X1 U19092 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16004), .A3(
        n16015), .ZN(n15998) );
  NAND2_X1 U19093 ( .A1(n16062), .A2(n9783), .ZN(n15995) );
  OAI21_X1 U19094 ( .B1(n20839), .B2(n15996), .A(n15995), .ZN(n15997) );
  NOR2_X1 U19095 ( .A1(n15998), .A2(n15997), .ZN(n16007) );
  OAI21_X1 U19096 ( .B1(n16004), .B2(n16000), .A(n15999), .ZN(n16001) );
  OAI211_X1 U19097 ( .C1(n16003), .C2(n16002), .A(n16026), .B(n16001), .ZN(
        n16012) );
  OAI221_X1 U19098 ( .B1(n16012), .B2(n16005), .C1(n16012), .C2(n16004), .A(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16006) );
  OAI211_X1 U19099 ( .C1(n16009), .C2(n16008), .A(n16007), .B(n16006), .ZN(
        P1_U3019) );
  AOI22_X1 U19100 ( .A1(n16062), .A2(n16010), .B1(n13376), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n16014) );
  AOI22_X1 U19101 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16012), .B1(
        n20087), .B2(n16011), .ZN(n16013) );
  OAI211_X1 U19102 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n16015), .A(
        n16014), .B(n16013), .ZN(P1_U3020) );
  AOI21_X1 U19103 ( .B1(n16018), .B2(n16017), .A(n16016), .ZN(n16025) );
  AOI22_X1 U19104 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16020), .B1(
        n20087), .B2(n16019), .ZN(n16024) );
  OAI221_X1 U19105 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n14508), .C2(n16022), .A(
        n16021), .ZN(n16023) );
  NAND3_X1 U19106 ( .A1(n16025), .A2(n16024), .A3(n16023), .ZN(P1_U3021) );
  OR2_X1 U19107 ( .A1(n16028), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16064) );
  NAND2_X1 U19108 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16030) );
  INV_X1 U19109 ( .A(n16026), .ZN(n16027) );
  AOI221_X1 U19110 ( .B1(n16030), .B2(n16029), .C1(n16028), .C2(n16029), .A(
        n16027), .ZN(n16069) );
  OAI21_X1 U19111 ( .B1(n16031), .B2(n16064), .A(n16069), .ZN(n16053) );
  AOI21_X1 U19112 ( .B1(n16036), .B2(n16032), .A(n16053), .ZN(n16050) );
  INV_X1 U19113 ( .A(n16033), .ZN(n16034) );
  AOI222_X1 U19114 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n13376), .B1(n16062), 
        .B2(n16035), .C1(n20087), .C2(n16034), .ZN(n16038) );
  INV_X1 U19115 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16049) );
  NOR2_X1 U19116 ( .A1(n16036), .A2(n16056), .ZN(n16045) );
  OAI221_X1 U19117 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16039), .C2(n16049), .A(
        n16045), .ZN(n16037) );
  OAI211_X1 U19118 ( .C1(n16050), .C2(n16039), .A(n16038), .B(n16037), .ZN(
        P1_U3023) );
  INV_X1 U19119 ( .A(n16051), .ZN(n16042) );
  INV_X1 U19120 ( .A(n16040), .ZN(n16041) );
  OAI21_X1 U19121 ( .B1(n16060), .B2(n16042), .A(n16041), .ZN(n16044) );
  AND2_X1 U19122 ( .A1(n16044), .A2(n16043), .ZN(n19996) );
  AOI22_X1 U19123 ( .A1(n16062), .A2(n19996), .B1(n13376), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16048) );
  AOI22_X1 U19124 ( .A1(n16046), .A2(n20087), .B1(n16049), .B2(n16045), .ZN(
        n16047) );
  OAI211_X1 U19125 ( .C1(n16050), .C2(n16049), .A(n16048), .B(n16047), .ZN(
        P1_U3024) );
  XNOR2_X1 U19126 ( .A(n16060), .B(n16051), .ZN(n20000) );
  AOI22_X1 U19127 ( .A1(n16062), .A2(n20000), .B1(n13376), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16055) );
  AOI22_X1 U19128 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16053), .B1(
        n16052), .B2(n20087), .ZN(n16054) );
  OAI211_X1 U19129 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16056), .A(
        n16055), .B(n16054), .ZN(P1_U3025) );
  OR2_X1 U19130 ( .A1(n16058), .A2(n16057), .ZN(n16059) );
  NAND2_X1 U19131 ( .A1(n16060), .A2(n16059), .ZN(n20004) );
  INV_X1 U19132 ( .A(n20004), .ZN(n19941) );
  AOI21_X1 U19133 ( .B1(n16062), .B2(n19941), .A(n16061), .ZN(n16063) );
  OAI21_X1 U19134 ( .B1(n16065), .B2(n16064), .A(n16063), .ZN(n16066) );
  AOI21_X1 U19135 ( .B1(n16067), .B2(n20087), .A(n16066), .ZN(n16068) );
  OAI21_X1 U19136 ( .B1(n16069), .B2(n13679), .A(n16068), .ZN(P1_U3026) );
  NAND4_X1 U19137 ( .A1(n16072), .A2(n16071), .A3(n16070), .A4(n19947), .ZN(
        n16073) );
  OAI21_X1 U19138 ( .B1(n16075), .B2(n16074), .A(n16073), .ZN(P1_U3468) );
  NAND2_X1 U19139 ( .A1(n20589), .A2(n20896), .ZN(n16082) );
  NAND4_X1 U19140 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20383), .A4(n20896), .ZN(n16076) );
  AND2_X1 U19141 ( .A1(n16077), .A2(n16076), .ZN(n20805) );
  AOI21_X1 U19142 ( .B1(n20805), .B2(n16079), .A(n16078), .ZN(n16081) );
  AOI21_X1 U19143 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n16084), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16080) );
  AOI211_X1 U19144 ( .C1(n20899), .C2(n16082), .A(n16081), .B(n16080), .ZN(
        P1_U3162) );
  OAI221_X1 U19145 ( .B1(n20589), .B2(P1_STATE2_REG_0__SCAN_IN), .C1(n20589), 
        .C2(n16084), .A(n16083), .ZN(P1_U3466) );
  AOI22_X1 U19146 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19045), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19028), .ZN(n16095) );
  AOI22_X1 U19147 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n19059), .B1(n16085), 
        .B2(n19057), .ZN(n16094) );
  INV_X1 U19148 ( .A(n16086), .ZN(n16088) );
  AOI22_X1 U19149 ( .A1(n16088), .A2(n19061), .B1(n16087), .B2(n19064), .ZN(
        n16093) );
  OAI211_X1 U19150 ( .C1(n16091), .C2(n16090), .A(n19036), .B(n16089), .ZN(
        n16092) );
  NAND4_X1 U19151 ( .A1(n16095), .A2(n16094), .A3(n16093), .A4(n16092), .ZN(
        P2_U2826) );
  AOI22_X1 U19152 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19045), .ZN(n16107) );
  AOI22_X1 U19153 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n19059), .B1(n16096), 
        .B2(n19057), .ZN(n16106) );
  INV_X1 U19154 ( .A(n16097), .ZN(n16100) );
  INV_X1 U19155 ( .A(n16098), .ZN(n16099) );
  AOI22_X1 U19156 ( .A1(n16100), .A2(n19061), .B1(n16099), .B2(n19064), .ZN(
        n16105) );
  OAI211_X1 U19157 ( .C1(n16103), .C2(n16102), .A(n19036), .B(n16101), .ZN(
        n16104) );
  NAND4_X1 U19158 ( .A1(n16107), .A2(n16106), .A3(n16105), .A4(n16104), .ZN(
        P2_U2827) );
  AOI22_X1 U19159 ( .A1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19045), .ZN(n16117) );
  AOI22_X1 U19160 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n19059), .B1(n16108), 
        .B2(n19057), .ZN(n16116) );
  AOI22_X1 U19161 ( .A1(n16110), .A2(n19061), .B1(n16109), .B2(n19064), .ZN(
        n16115) );
  OAI211_X1 U19162 ( .C1(n16113), .C2(n16112), .A(n19036), .B(n16111), .ZN(
        n16114) );
  NAND4_X1 U19163 ( .A1(n16117), .A2(n16116), .A3(n16115), .A4(n16114), .ZN(
        P2_U2828) );
  AOI22_X1 U19164 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19045), .ZN(n16128) );
  AOI22_X1 U19165 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n19059), .B1(n16118), 
        .B2(n19057), .ZN(n16127) );
  INV_X1 U19166 ( .A(n16119), .ZN(n16121) );
  AOI22_X1 U19167 ( .A1(n16121), .A2(n19061), .B1(n16120), .B2(n19064), .ZN(
        n16126) );
  OAI211_X1 U19168 ( .C1(n16124), .C2(n16123), .A(n19036), .B(n16122), .ZN(
        n16125) );
  NAND4_X1 U19169 ( .A1(n16128), .A2(n16127), .A3(n16126), .A4(n16125), .ZN(
        P2_U2829) );
  AOI22_X1 U19170 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19045), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19028), .ZN(n16140) );
  INV_X1 U19171 ( .A(n16129), .ZN(n16130) );
  AOI22_X1 U19172 ( .A1(n16130), .A2(n19057), .B1(P2_EBX_REG_25__SCAN_IN), 
        .B2(n19059), .ZN(n16139) );
  OAI22_X1 U19173 ( .A1(n16132), .A2(n19049), .B1(n16131), .B2(n19011), .ZN(
        n16133) );
  INV_X1 U19174 ( .A(n16133), .ZN(n16138) );
  OAI211_X1 U19175 ( .C1(n16136), .C2(n16135), .A(n19036), .B(n16134), .ZN(
        n16137) );
  NAND4_X1 U19176 ( .A1(n16140), .A2(n16139), .A3(n16138), .A4(n16137), .ZN(
        P2_U2830) );
  AOI22_X1 U19177 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n19045), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19028), .ZN(n16151) );
  AOI22_X1 U19178 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19059), .B1(n16141), 
        .B2(n19057), .ZN(n16150) );
  OAI22_X1 U19179 ( .A1(n16143), .A2(n19049), .B1(n16142), .B2(n19011), .ZN(
        n16144) );
  INV_X1 U19180 ( .A(n16144), .ZN(n16149) );
  OAI211_X1 U19181 ( .C1(n16147), .C2(n16146), .A(n19036), .B(n16145), .ZN(
        n16148) );
  NAND4_X1 U19182 ( .A1(n16151), .A2(n16150), .A3(n16149), .A4(n16148), .ZN(
        P2_U2831) );
  AOI22_X1 U19183 ( .A1(P2_REIP_REG_23__SCAN_IN), .A2(n19045), .B1(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19028), .ZN(n16161) );
  AOI22_X1 U19184 ( .A1(P2_EBX_REG_23__SCAN_IN), .A2(n19059), .B1(n16152), 
        .B2(n19057), .ZN(n16160) );
  OAI22_X1 U19185 ( .A1(n16153), .A2(n19049), .B1(n16166), .B2(n19011), .ZN(
        n16154) );
  INV_X1 U19186 ( .A(n16154), .ZN(n16159) );
  OAI211_X1 U19187 ( .C1(n16157), .C2(n16156), .A(n19036), .B(n16155), .ZN(
        n16158) );
  NAND4_X1 U19188 ( .A1(n16161), .A2(n16160), .A3(n16159), .A4(n16158), .ZN(
        P2_U2832) );
  INV_X1 U19189 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16162) );
  AOI22_X1 U19190 ( .A1(n19103), .A2(n16163), .B1(n16162), .B2(n19089), .ZN(
        P2_U2856) );
  AOI22_X1 U19191 ( .A1(n16164), .A2(n19100), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n19089), .ZN(n16165) );
  OAI21_X1 U19192 ( .B1(n19089), .B2(n16166), .A(n16165), .ZN(P2_U2864) );
  INV_X1 U19193 ( .A(n16167), .ZN(n16169) );
  AOI22_X1 U19194 ( .A1(n16169), .A2(n19100), .B1(n19103), .B2(n16168), .ZN(
        n16170) );
  OAI21_X1 U19195 ( .B1(n19103), .B2(n10899), .A(n16170), .ZN(P2_U2865) );
  INV_X1 U19196 ( .A(n14983), .ZN(n16173) );
  NAND2_X1 U19197 ( .A1(n14704), .A2(n16171), .ZN(n16172) );
  NAND2_X1 U19198 ( .A1(n16173), .A2(n16172), .ZN(n16185) );
  OAI22_X1 U19199 ( .A1(n16185), .A2(n19095), .B1(n19089), .B2(n16174), .ZN(
        n16175) );
  INV_X1 U19200 ( .A(n16175), .ZN(n16176) );
  OAI21_X1 U19201 ( .B1(n19103), .B2(n16177), .A(n16176), .ZN(P2_U2867) );
  OR2_X1 U19202 ( .A1(n16179), .A2(n16178), .ZN(n16180) );
  NAND2_X1 U19203 ( .A1(n14046), .A2(n16180), .ZN(n16192) );
  OAI22_X1 U19204 ( .A1(n16192), .A2(n19095), .B1(n19103), .B2(n16181), .ZN(
        n16182) );
  INV_X1 U19205 ( .A(n16182), .ZN(n16183) );
  OAI21_X1 U19206 ( .B1(n19089), .B2(n18903), .A(n16183), .ZN(P2_U2869) );
  AOI22_X1 U19207 ( .A1(n19109), .A2(n16184), .B1(n19170), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16190) );
  AOI22_X1 U19208 ( .A1(n19111), .A2(BUF2_REG_20__SCAN_IN), .B1(n19110), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n16189) );
  OAI22_X1 U19209 ( .A1(n16186), .A2(n19153), .B1(n19145), .B2(n16185), .ZN(
        n16187) );
  INV_X1 U19210 ( .A(n16187), .ZN(n16188) );
  NAND3_X1 U19211 ( .A1(n16190), .A2(n16189), .A3(n16188), .ZN(P2_U2899) );
  INV_X1 U19212 ( .A(n16191), .ZN(n19162) );
  AOI22_X1 U19213 ( .A1(n19109), .A2(n19162), .B1(n19170), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16196) );
  AOI22_X1 U19214 ( .A1(n19111), .A2(BUF2_REG_18__SCAN_IN), .B1(n19110), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n16195) );
  OAI22_X1 U19215 ( .A1(n18904), .A2(n19153), .B1(n19145), .B2(n16192), .ZN(
        n16193) );
  INV_X1 U19216 ( .A(n16193), .ZN(n16194) );
  NAND3_X1 U19217 ( .A1(n16196), .A2(n16195), .A3(n16194), .ZN(P2_U2901) );
  AOI22_X1 U19218 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19217), .B1(n16268), 
        .B2(n18930), .ZN(n16201) );
  OAI211_X1 U19219 ( .C1(n10820), .C2(n16278), .A(n16201), .B(n16200), .ZN(
        P2_U2999) );
  AOI22_X1 U19220 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19218), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19217), .ZN(n16210) );
  OAI21_X1 U19221 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16203), .A(
        n16202), .ZN(n16293) );
  NAND2_X1 U19222 ( .A1(n16205), .A2(n16204), .ZN(n16207) );
  XOR2_X1 U19223 ( .A(n16207), .B(n16206), .Z(n16289) );
  OAI22_X1 U19224 ( .A1(n16293), .A2(n19219), .B1(n19221), .B2(n16289), .ZN(
        n16208) );
  AOI21_X1 U19225 ( .B1(n19225), .B2(n18937), .A(n16208), .ZN(n16209) );
  OAI211_X1 U19226 ( .C1(n19229), .C2(n18933), .A(n16210), .B(n16209), .ZN(
        P2_U3000) );
  AOI22_X1 U19227 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19217), .B1(n16268), 
        .B2(n18941), .ZN(n16215) );
  INV_X1 U19228 ( .A(n16211), .ZN(n16212) );
  AOI222_X1 U19229 ( .A1(n16213), .A2(n16269), .B1(n11389), .B2(n16212), .C1(
        n19225), .C2(n18945), .ZN(n16214) );
  OAI211_X1 U19230 ( .C1(n16216), .C2(n16278), .A(n16215), .B(n16214), .ZN(
        P2_U3001) );
  AOI22_X1 U19231 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19217), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19218), .ZN(n16222) );
  INV_X1 U19232 ( .A(n16217), .ZN(n18962) );
  OAI22_X1 U19233 ( .A1(n16219), .A2(n19219), .B1(n16218), .B2(n19221), .ZN(
        n16220) );
  AOI21_X1 U19234 ( .B1(n19225), .B2(n18962), .A(n16220), .ZN(n16221) );
  OAI211_X1 U19235 ( .C1(n19229), .C2(n18960), .A(n16222), .B(n16221), .ZN(
        P2_U3002) );
  AOI22_X1 U19236 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19217), .B1(n16268), 
        .B2(n18971), .ZN(n16235) );
  INV_X1 U19237 ( .A(n16223), .ZN(n16224) );
  NAND2_X1 U19238 ( .A1(n16225), .A2(n16224), .ZN(n16229) );
  OR2_X1 U19239 ( .A1(n16227), .A2(n16226), .ZN(n16228) );
  XNOR2_X1 U19240 ( .A(n16229), .B(n16228), .ZN(n16305) );
  INV_X1 U19241 ( .A(n16303), .ZN(n18972) );
  NAND2_X1 U19242 ( .A1(n16230), .A2(n16300), .ZN(n16232) );
  NAND2_X1 U19243 ( .A1(n16232), .A2(n16231), .ZN(n16308) );
  INV_X1 U19244 ( .A(n16308), .ZN(n16233) );
  AOI222_X1 U19245 ( .A1(n16305), .A2(n11389), .B1(n19225), .B2(n18972), .C1(
        n16269), .C2(n16233), .ZN(n16234) );
  OAI211_X1 U19246 ( .C1(n10861), .C2(n16278), .A(n16235), .B(n16234), .ZN(
        P2_U3003) );
  AOI22_X1 U19247 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19217), .B1(n16268), 
        .B2(n18987), .ZN(n16240) );
  AOI222_X1 U19248 ( .A1(n16238), .A2(n16269), .B1(n11389), .B2(n16237), .C1(
        n19225), .C2(n16236), .ZN(n16239) );
  OAI211_X1 U19249 ( .C1(n10825), .C2(n16278), .A(n16240), .B(n16239), .ZN(
        P2_U3005) );
  AOI22_X1 U19250 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19218), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19217), .ZN(n16257) );
  NAND2_X1 U19251 ( .A1(n16241), .A2(n13303), .ZN(n16244) );
  INV_X1 U19252 ( .A(n16242), .ZN(n16243) );
  AND2_X1 U19253 ( .A1(n16244), .A2(n16243), .ZN(n19098) );
  XOR2_X1 U19254 ( .A(n16245), .B(n16246), .Z(n16315) );
  AOI21_X1 U19255 ( .B1(n13896), .B2(n16248), .A(n16247), .ZN(n16253) );
  INV_X1 U19256 ( .A(n16249), .ZN(n16251) );
  NOR2_X1 U19257 ( .A1(n16251), .A2(n16250), .ZN(n16252) );
  XNOR2_X1 U19258 ( .A(n16253), .B(n16252), .ZN(n16318) );
  AOI22_X1 U19259 ( .A1(n16315), .A2(n16269), .B1(n11389), .B2(n16318), .ZN(
        n16254) );
  INV_X1 U19260 ( .A(n16254), .ZN(n16255) );
  AOI21_X1 U19261 ( .B1(n19225), .B2(n19098), .A(n16255), .ZN(n16256) );
  OAI211_X1 U19262 ( .C1(n19229), .C2(n18997), .A(n16257), .B(n16256), .ZN(
        P2_U3006) );
  AOI22_X1 U19263 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n19218), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n19217), .ZN(n16262) );
  OAI22_X1 U19264 ( .A1(n16259), .A2(n19219), .B1(n19221), .B2(n16258), .ZN(
        n16260) );
  AOI21_X1 U19265 ( .B1(n19225), .B2(n19024), .A(n16260), .ZN(n16261) );
  OAI211_X1 U19266 ( .C1(n19229), .C2(n19022), .A(n16262), .B(n16261), .ZN(
        P2_U3008) );
  AOI22_X1 U19267 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19217), .B1(n16268), 
        .B2(n19034), .ZN(n16266) );
  AOI222_X1 U19268 ( .A1(n16264), .A2(n11389), .B1(n16269), .B2(n16263), .C1(
        n19225), .C2(n19035), .ZN(n16265) );
  OAI211_X1 U19269 ( .C1(n10838), .C2(n16278), .A(n16266), .B(n16265), .ZN(
        P2_U3009) );
  AOI22_X1 U19270 ( .A1(P2_REIP_REG_3__SCAN_IN), .A2(n19217), .B1(n16268), 
        .B2(n16267), .ZN(n16277) );
  NAND3_X1 U19271 ( .A1(n16270), .A2(n13591), .A3(n16269), .ZN(n16271) );
  OAI21_X1 U19272 ( .B1(n16273), .B2(n16272), .A(n16271), .ZN(n16274) );
  AOI21_X1 U19273 ( .B1(n16275), .B2(n11389), .A(n16274), .ZN(n16276) );
  OAI211_X1 U19274 ( .C1(n10343), .C2(n16278), .A(n16277), .B(n16276), .ZN(
        P2_U3011) );
  AOI21_X1 U19275 ( .B1(n16281), .B2(n16280), .A(n16279), .ZN(n19120) );
  NOR2_X1 U19276 ( .A1(n16283), .A2(n16282), .ZN(n16286) );
  INV_X1 U19277 ( .A(n16284), .ZN(n16285) );
  MUX2_X1 U19278 ( .A(n16286), .B(n16285), .S(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n16288) );
  INV_X1 U19279 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19778) );
  NOR2_X1 U19280 ( .A1(n19046), .A2(n19778), .ZN(n16287) );
  AOI211_X1 U19281 ( .C1(n19120), .C2(n16312), .A(n16288), .B(n16287), .ZN(
        n16292) );
  INV_X1 U19282 ( .A(n16289), .ZN(n16290) );
  AOI22_X1 U19283 ( .A1(n16290), .A2(n16317), .B1(n16316), .B2(n18937), .ZN(
        n16291) );
  OAI211_X1 U19284 ( .C1(n16339), .C2(n16293), .A(n16292), .B(n16291), .ZN(
        P2_U3032) );
  AOI211_X1 U19285 ( .C1(n10651), .C2(n16300), .A(n16295), .B(n16294), .ZN(
        n16302) );
  OAI21_X1 U19286 ( .B1(n16298), .B2(n16297), .A(n16296), .ZN(n19130) );
  OAI22_X1 U19287 ( .A1(n19130), .A2(n16330), .B1(n16300), .B2(n16299), .ZN(
        n16301) );
  AOI211_X1 U19288 ( .C1(n19217), .C2(P2_REIP_REG_11__SCAN_IN), .A(n16302), 
        .B(n16301), .ZN(n16307) );
  NOR2_X1 U19289 ( .A1(n16327), .A2(n16303), .ZN(n16304) );
  AOI21_X1 U19290 ( .B1(n16305), .B2(n16317), .A(n16304), .ZN(n16306) );
  OAI211_X1 U19291 ( .C1(n16339), .C2(n16308), .A(n16307), .B(n16306), .ZN(
        P2_U3035) );
  AOI21_X1 U19292 ( .B1(n16311), .B2(n16310), .A(n16309), .ZN(n19137) );
  AOI22_X1 U19293 ( .A1(n16313), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16312), .B2(n19137), .ZN(n16324) );
  AOI222_X1 U19294 ( .A1(n16318), .A2(n16317), .B1(n16316), .B2(n19098), .C1(
        n16315), .C2(n16314), .ZN(n16323) );
  NAND2_X1 U19295 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19217), .ZN(n16322) );
  OAI221_X1 U19296 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C1(n9956), .C2(n16320), .A(n16319), .ZN(n16321) );
  NAND4_X1 U19297 ( .A1(n16324), .A2(n16323), .A3(n16322), .A4(n16321), .ZN(
        P2_U3038) );
  OAI22_X1 U19298 ( .A1(n16328), .A2(n16327), .B1(n16326), .B2(n16325), .ZN(
        n16333) );
  OAI22_X1 U19299 ( .A1(n16331), .A2(n16335), .B1(n16330), .B2(n16329), .ZN(
        n16332) );
  AOI211_X1 U19300 ( .C1(n16335), .C2(n16334), .A(n16333), .B(n16332), .ZN(
        n16337) );
  OAI211_X1 U19301 ( .C1(n16339), .C2(n16338), .A(n16337), .B(n16336), .ZN(
        P2_U3046) );
  INV_X1 U19302 ( .A(n16340), .ZN(n16354) );
  AOI21_X1 U19303 ( .B1(n16343), .B2(n16342), .A(n16341), .ZN(n16344) );
  NOR2_X1 U19304 ( .A1(n16345), .A2(n16344), .ZN(n16349) );
  NAND2_X1 U19305 ( .A1(n16346), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19848) );
  AOI21_X1 U19306 ( .B1(n16347), .B2(n19848), .A(n16342), .ZN(n16348) );
  AOI211_X1 U19307 ( .C1(n16351), .C2(n16350), .A(n16349), .B(n16348), .ZN(
        n16353) );
  OAI211_X1 U19308 ( .C1(n16355), .C2(n16354), .A(n16353), .B(n16352), .ZN(
        P2_U3176) );
  NOR2_X1 U19309 ( .A1(n17767), .A2(n16357), .ZN(n16365) );
  NAND2_X1 U19310 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17767), .ZN(
        n16360) );
  OAI211_X1 U19311 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n17767), .A(
        n16358), .B(n16360), .ZN(n16364) );
  OAI21_X1 U19312 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16416), .A(
        n16359), .ZN(n16362) );
  OAI22_X1 U19313 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17767), .B1(
        n16360), .B2(n16416), .ZN(n16361) );
  OAI21_X1 U19314 ( .B1(n16365), .B2(n16362), .A(n16361), .ZN(n16363) );
  OAI21_X1 U19315 ( .B1(n16365), .B2(n16364), .A(n16363), .ZN(n16421) );
  INV_X1 U19316 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16546) );
  INV_X1 U19317 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16580) );
  NAND2_X1 U19318 ( .A1(n17806), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n16738) );
  NOR2_X1 U19319 ( .A1(n21064), .A2(n17761), .ZN(n16774) );
  NAND2_X1 U19320 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17692) );
  NAND2_X1 U19321 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17651) );
  NAND2_X1 U19322 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17613) );
  NAND2_X1 U19323 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17583) );
  NAND2_X1 U19324 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17562), .ZN(
        n17535) );
  NAND2_X1 U19325 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17536) );
  NAND2_X1 U19326 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16392), .ZN(
        n16382) );
  XOR2_X2 U19327 ( .A(n16546), .B(n16382), .Z(n16872) );
  INV_X1 U19328 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18777) );
  NOR2_X1 U19329 ( .A1(n18777), .A2(n18077), .ZN(n16412) );
  INV_X1 U19330 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16564) );
  NAND3_X1 U19331 ( .A1(n17493), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16395) );
  NOR2_X1 U19332 ( .A1(n16580), .A2(n16395), .ZN(n16367) );
  NAND2_X1 U19333 ( .A1(n18843), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18702) );
  INV_X1 U19334 ( .A(n17691), .ZN(n17492) );
  NAND2_X1 U19335 ( .A1(n16367), .A2(n17492), .ZN(n16381) );
  NOR2_X1 U19336 ( .A1(n16564), .A2(n16381), .ZN(n16372) );
  NOR2_X1 U19337 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17600), .ZN(
        n16397) );
  NOR2_X1 U19338 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16381), .ZN(
        n16370) );
  INV_X1 U19339 ( .A(n18702), .ZN(n17687) );
  INV_X1 U19340 ( .A(n16367), .ZN(n16368) );
  AOI22_X1 U19341 ( .A1(n17687), .A2(n16552), .B1(n18566), .B2(n16368), .ZN(
        n16369) );
  NAND2_X1 U19342 ( .A1(n16369), .A2(n17858), .ZN(n16393) );
  NOR3_X1 U19343 ( .A1(n16397), .A2(n16370), .A3(n16393), .ZN(n16380) );
  INV_X1 U19344 ( .A(n16380), .ZN(n16371) );
  MUX2_X1 U19345 ( .A(n16372), .B(n16371), .S(
        P3_PHYADDRPOINTER_REG_31__SCAN_IN), .Z(n16373) );
  INV_X1 U19346 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18802) );
  NAND2_X1 U19347 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16388), .ZN(
        n16374) );
  XOR2_X1 U19348 ( .A(n18802), .B(n16374), .Z(n16413) );
  NAND2_X1 U19349 ( .A1(n17341), .A2(n16375), .ZN(n17546) );
  NAND2_X1 U19350 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16387), .ZN(
        n16376) );
  XOR2_X1 U19351 ( .A(n18802), .B(n16376), .Z(n16417) );
  AOI22_X1 U19352 ( .A1(n17850), .A2(n16413), .B1(n17770), .B2(n16417), .ZN(
        n16377) );
  OAI211_X1 U19353 ( .C1(n17742), .C2(n16421), .A(n16378), .B(n16377), .ZN(
        P3_U2799) );
  NOR2_X2 U19354 ( .A1(n17647), .A2(n17755), .ZN(n17641) );
  INV_X1 U19355 ( .A(n17641), .ZN(n17658) );
  NOR2_X1 U19356 ( .A1(n16379), .A2(n17658), .ZN(n17519) );
  AOI21_X1 U19357 ( .B1(n16564), .B2(n16381), .A(n16380), .ZN(n16385) );
  OAI21_X1 U19358 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16392), .A(
        n16382), .ZN(n16563) );
  OAI21_X1 U19359 ( .B1(n17696), .B2(n16563), .A(n16383), .ZN(n16384) );
  AOI211_X1 U19360 ( .C1(n17519), .C2(n16386), .A(n16385), .B(n16384), .ZN(
        n16390) );
  NOR2_X1 U19361 ( .A1(n16387), .A2(n17546), .ZN(n16401) );
  NOR2_X1 U19362 ( .A1(n16388), .A2(n17862), .ZN(n16404) );
  OAI21_X1 U19363 ( .B1(n16401), .B2(n16404), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16389) );
  OAI211_X1 U19364 ( .C1(n16391), .C2(n17742), .A(n16390), .B(n16389), .ZN(
        P3_U2800) );
  AOI21_X1 U19365 ( .B1(n16580), .B2(n16552), .A(n16392), .ZN(n16574) );
  INV_X1 U19366 ( .A(n16393), .ZN(n16394) );
  AOI221_X1 U19367 ( .B1(n17816), .B2(n16580), .C1(n16395), .C2(n16580), .A(
        n16394), .ZN(n16396) );
  AOI221_X1 U19368 ( .B1(n16397), .B2(n16574), .C1(n17706), .C2(n16574), .A(
        n16396), .ZN(n16409) );
  NAND2_X1 U19369 ( .A1(n16399), .A2(n16398), .ZN(n16400) );
  AOI22_X1 U19370 ( .A1(n17768), .A2(n16402), .B1(n16401), .B2(n16400), .ZN(
        n16408) );
  NOR2_X1 U19371 ( .A1(n17498), .A2(n16403), .ZN(n16405) );
  OAI21_X1 U19372 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n16405), .A(
        n16404), .ZN(n16406) );
  NAND4_X1 U19373 ( .A1(n16409), .A2(n16408), .A3(n16407), .A4(n16406), .ZN(
        P3_U2801) );
  INV_X1 U19374 ( .A(n18140), .ZN(n18170) );
  AOI221_X1 U19375 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16410), 
        .C1(n18160), .C2(n16410), .A(n18802), .ZN(n16411) );
  AOI211_X1 U19376 ( .C1(n16413), .C2(n18170), .A(n16412), .B(n16411), .ZN(
        n16420) );
  NOR4_X1 U19377 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16416), .A3(
        n16415), .A4(n16414), .ZN(n16418) );
  OAI221_X1 U19378 ( .B1(n16418), .B2(n16417), .C1(n16418), .C2(n18031), .A(
        n18158), .ZN(n16419) );
  OAI211_X1 U19379 ( .C1(n16421), .C2(n18070), .A(n16420), .B(n16419), .ZN(
        P3_U2831) );
  NOR3_X1 U19380 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16423) );
  NOR4_X1 U19381 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16422) );
  NAND4_X1 U19382 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16423), .A3(n16422), .A4(
        U215), .ZN(U213) );
  INV_X1 U19383 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19180) );
  NOR2_X2 U19384 ( .A1(n16464), .A2(n16424), .ZN(n16473) );
  OAI222_X1 U19385 ( .A1(U212), .A2(n19180), .B1(n16477), .B2(n16425), .C1(
        U214), .C2(n16513), .ZN(U216) );
  INV_X1 U19386 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16427) );
  AOI22_X1 U19387 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16475), .ZN(n16426) );
  OAI21_X1 U19388 ( .B1(n16427), .B2(n16477), .A(n16426), .ZN(U217) );
  INV_X1 U19389 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16429) );
  AOI22_X1 U19390 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16475), .ZN(n16428) );
  OAI21_X1 U19391 ( .B1(n16429), .B2(n16477), .A(n16428), .ZN(U218) );
  INV_X1 U19392 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16431) );
  AOI22_X1 U19393 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16475), .ZN(n16430) );
  OAI21_X1 U19394 ( .B1(n16431), .B2(n16477), .A(n16430), .ZN(U219) );
  INV_X1 U19395 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16433) );
  AOI22_X1 U19396 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16475), .ZN(n16432) );
  OAI21_X1 U19397 ( .B1(n16433), .B2(n16477), .A(n16432), .ZN(U220) );
  INV_X1 U19398 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20945) );
  AOI22_X1 U19399 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16475), .ZN(n16434) );
  OAI21_X1 U19400 ( .B1(n20945), .B2(n16477), .A(n16434), .ZN(U221) );
  INV_X1 U19401 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16436) );
  AOI22_X1 U19402 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16475), .ZN(n16435) );
  OAI21_X1 U19403 ( .B1(n16436), .B2(n16477), .A(n16435), .ZN(U222) );
  INV_X1 U19404 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16438) );
  AOI22_X1 U19405 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16475), .ZN(n16437) );
  OAI21_X1 U19406 ( .B1(n16438), .B2(n16477), .A(n16437), .ZN(U223) );
  INV_X1 U19407 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16440) );
  AOI22_X1 U19408 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16475), .ZN(n16439) );
  OAI21_X1 U19409 ( .B1(n16440), .B2(n16477), .A(n16439), .ZN(U224) );
  INV_X1 U19410 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n16442) );
  AOI22_X1 U19411 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16475), .ZN(n16441) );
  OAI21_X1 U19412 ( .B1(n16442), .B2(n16477), .A(n16441), .ZN(U225) );
  AOI22_X1 U19413 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16475), .ZN(n16443) );
  OAI21_X1 U19414 ( .B1(n16444), .B2(n16477), .A(n16443), .ZN(U226) );
  INV_X1 U19415 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n20956) );
  AOI22_X1 U19416 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16464), .ZN(n16445) );
  OAI21_X1 U19417 ( .B1(n20956), .B2(U212), .A(n16445), .ZN(U227) );
  INV_X1 U19418 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16447) );
  AOI22_X1 U19419 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16475), .ZN(n16446) );
  OAI21_X1 U19420 ( .B1(n16447), .B2(n16477), .A(n16446), .ZN(U228) );
  AOI22_X1 U19421 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16475), .ZN(n16448) );
  OAI21_X1 U19422 ( .B1(n14393), .B2(n16477), .A(n16448), .ZN(U229) );
  INV_X1 U19423 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n21074) );
  AOI22_X1 U19424 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16475), .ZN(n16449) );
  OAI21_X1 U19425 ( .B1(n21074), .B2(n16477), .A(n16449), .ZN(U230) );
  AOI222_X1 U19426 ( .A1(n16475), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n16473), 
        .B2(BUF1_REG_16__SCAN_IN), .C1(n16464), .C2(P1_DATAO_REG_16__SCAN_IN), 
        .ZN(n16450) );
  INV_X1 U19427 ( .A(n16450), .ZN(U231) );
  INV_X1 U19428 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n16452) );
  AOI22_X1 U19429 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16464), .ZN(n16451) );
  OAI21_X1 U19430 ( .B1(n16452), .B2(U212), .A(n16451), .ZN(U232) );
  INV_X1 U19431 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16454) );
  AOI22_X1 U19432 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16464), .ZN(n16453) );
  OAI21_X1 U19433 ( .B1(n16454), .B2(U212), .A(n16453), .ZN(U233) );
  INV_X1 U19434 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16456) );
  AOI22_X1 U19435 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16464), .ZN(n16455) );
  OAI21_X1 U19436 ( .B1(n16456), .B2(U212), .A(n16455), .ZN(U234) );
  INV_X1 U19437 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n16458) );
  AOI22_X1 U19438 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16475), .ZN(n16457) );
  OAI21_X1 U19439 ( .B1(n16458), .B2(n16477), .A(n16457), .ZN(U235) );
  INV_X1 U19440 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16490) );
  AOI22_X1 U19441 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16464), .ZN(n16459) );
  OAI21_X1 U19442 ( .B1(n16490), .B2(U212), .A(n16459), .ZN(U236) );
  INV_X1 U19443 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16461) );
  AOI22_X1 U19444 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n16475), .ZN(n16460) );
  OAI21_X1 U19445 ( .B1(n16461), .B2(n16477), .A(n16460), .ZN(U237) );
  INV_X1 U19446 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16488) );
  AOI22_X1 U19447 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16464), .ZN(n16462) );
  OAI21_X1 U19448 ( .B1(n16488), .B2(U212), .A(n16462), .ZN(U238) );
  INV_X1 U19449 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16487) );
  INV_X1 U19450 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n21043) );
  OAI222_X1 U19451 ( .A1(U212), .A2(n16487), .B1(n16477), .B2(n16463), .C1(
        U214), .C2(n21043), .ZN(U239) );
  INV_X1 U19452 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16486) );
  AOI22_X1 U19453 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16464), .ZN(n16465) );
  OAI21_X1 U19454 ( .B1(n16486), .B2(U212), .A(n16465), .ZN(U240) );
  INV_X1 U19455 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16485) );
  AOI22_X1 U19456 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16464), .ZN(n16466) );
  OAI21_X1 U19457 ( .B1(n16485), .B2(U212), .A(n16466), .ZN(U241) );
  INV_X1 U19458 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16484) );
  AOI22_X1 U19459 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16464), .ZN(n16467) );
  OAI21_X1 U19460 ( .B1(n16484), .B2(U212), .A(n16467), .ZN(U242) );
  INV_X1 U19461 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16469) );
  AOI22_X1 U19462 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16475), .ZN(n16468) );
  OAI21_X1 U19463 ( .B1(n16469), .B2(n16477), .A(n16468), .ZN(U243) );
  INV_X1 U19464 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16482) );
  AOI22_X1 U19465 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16464), .ZN(n16470) );
  OAI21_X1 U19466 ( .B1(n16482), .B2(U212), .A(n16470), .ZN(U244) );
  INV_X1 U19467 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16472) );
  AOI22_X1 U19468 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16475), .ZN(n16471) );
  OAI21_X1 U19469 ( .B1(n16472), .B2(n16477), .A(n16471), .ZN(U245) );
  INV_X1 U19470 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16480) );
  AOI22_X1 U19471 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16473), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16464), .ZN(n16474) );
  OAI21_X1 U19472 ( .B1(n16480), .B2(U212), .A(n16474), .ZN(U246) );
  INV_X1 U19473 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16478) );
  AOI22_X1 U19474 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16464), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16475), .ZN(n16476) );
  OAI21_X1 U19475 ( .B1(n16478), .B2(n16477), .A(n16476), .ZN(U247) );
  OAI22_X1 U19476 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16511), .ZN(n16479) );
  INV_X1 U19477 ( .A(n16479), .ZN(U251) );
  INV_X1 U19478 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18191) );
  AOI22_X1 U19479 ( .A1(n16511), .A2(n16480), .B1(n18191), .B2(U215), .ZN(U252) );
  OAI22_X1 U19480 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16499), .ZN(n16481) );
  INV_X1 U19481 ( .A(n16481), .ZN(U253) );
  INV_X1 U19482 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18199) );
  AOI22_X1 U19483 ( .A1(n16511), .A2(n16482), .B1(n18199), .B2(U215), .ZN(U254) );
  OAI22_X1 U19484 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16499), .ZN(n16483) );
  INV_X1 U19485 ( .A(n16483), .ZN(U255) );
  INV_X1 U19486 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18207) );
  AOI22_X1 U19487 ( .A1(n16511), .A2(n16484), .B1(n18207), .B2(U215), .ZN(U256) );
  INV_X1 U19488 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18211) );
  AOI22_X1 U19489 ( .A1(n16511), .A2(n16485), .B1(n18211), .B2(U215), .ZN(U257) );
  INV_X1 U19490 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18216) );
  AOI22_X1 U19491 ( .A1(n16511), .A2(n16486), .B1(n18216), .B2(U215), .ZN(U258) );
  INV_X1 U19492 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17471) );
  AOI22_X1 U19493 ( .A1(n16511), .A2(n16487), .B1(n17471), .B2(U215), .ZN(U259) );
  INV_X1 U19494 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17473) );
  AOI22_X1 U19495 ( .A1(n16511), .A2(n16488), .B1(n17473), .B2(U215), .ZN(U260) );
  OAI22_X1 U19496 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16499), .ZN(n16489) );
  INV_X1 U19497 ( .A(n16489), .ZN(U261) );
  INV_X1 U19498 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n21082) );
  AOI22_X1 U19499 ( .A1(n16511), .A2(n16490), .B1(n21082), .B2(U215), .ZN(U262) );
  OAI22_X1 U19500 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16499), .ZN(n16491) );
  INV_X1 U19501 ( .A(n16491), .ZN(U263) );
  OAI22_X1 U19502 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16499), .ZN(n16492) );
  INV_X1 U19503 ( .A(n16492), .ZN(U264) );
  OAI22_X1 U19504 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16499), .ZN(n16493) );
  INV_X1 U19505 ( .A(n16493), .ZN(U265) );
  OAI22_X1 U19506 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16499), .ZN(n16494) );
  INV_X1 U19507 ( .A(n16494), .ZN(U266) );
  OAI22_X1 U19508 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16511), .ZN(n16495) );
  INV_X1 U19509 ( .A(n16495), .ZN(U267) );
  OAI22_X1 U19510 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16499), .ZN(n16496) );
  INV_X1 U19511 ( .A(n16496), .ZN(U268) );
  OAI22_X1 U19512 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16511), .ZN(n16497) );
  INV_X1 U19513 ( .A(n16497), .ZN(U269) );
  OAI22_X1 U19514 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16499), .ZN(n16498) );
  INV_X1 U19515 ( .A(n16498), .ZN(U270) );
  OAI22_X1 U19516 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16499), .ZN(n16500) );
  INV_X1 U19517 ( .A(n16500), .ZN(U271) );
  OAI22_X1 U19518 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16511), .ZN(n16501) );
  INV_X1 U19519 ( .A(n16501), .ZN(U272) );
  OAI22_X1 U19520 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16511), .ZN(n16502) );
  INV_X1 U19521 ( .A(n16502), .ZN(U273) );
  OAI22_X1 U19522 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16511), .ZN(n16503) );
  INV_X1 U19523 ( .A(n16503), .ZN(U274) );
  OAI22_X1 U19524 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16511), .ZN(n16504) );
  INV_X1 U19525 ( .A(n16504), .ZN(U275) );
  OAI22_X1 U19526 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16511), .ZN(n16505) );
  INV_X1 U19527 ( .A(n16505), .ZN(U276) );
  OAI22_X1 U19528 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16511), .ZN(n16506) );
  INV_X1 U19529 ( .A(n16506), .ZN(U277) );
  OAI22_X1 U19530 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16511), .ZN(n16507) );
  INV_X1 U19531 ( .A(n16507), .ZN(U278) );
  OAI22_X1 U19532 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16511), .ZN(n16508) );
  INV_X1 U19533 ( .A(n16508), .ZN(U279) );
  OAI22_X1 U19534 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16511), .ZN(n16509) );
  INV_X1 U19535 ( .A(n16509), .ZN(U280) );
  OAI22_X1 U19536 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16511), .ZN(n16510) );
  INV_X1 U19537 ( .A(n16510), .ZN(U281) );
  OAI22_X1 U19538 ( .A1(U215), .A2(P2_DATAO_REG_31__SCAN_IN), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n16511), .ZN(n16512) );
  INV_X1 U19539 ( .A(n16512), .ZN(U282) );
  INV_X1 U19540 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17379) );
  AOI222_X1 U19541 ( .A1(n16513), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n17379), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16514) );
  INV_X2 U19542 ( .A(n16516), .ZN(n16515) );
  INV_X1 U19543 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18737) );
  INV_X1 U19544 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19771) );
  AOI22_X1 U19545 ( .A1(n16515), .A2(n18737), .B1(n19771), .B2(n16516), .ZN(
        U347) );
  INV_X1 U19546 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18735) );
  INV_X1 U19547 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19769) );
  AOI22_X1 U19548 ( .A1(n16515), .A2(n18735), .B1(n19769), .B2(n16516), .ZN(
        U348) );
  INV_X1 U19549 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18733) );
  INV_X1 U19550 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19767) );
  AOI22_X1 U19551 ( .A1(n16515), .A2(n18733), .B1(n19767), .B2(n16516), .ZN(
        U349) );
  INV_X1 U19552 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18731) );
  INV_X1 U19553 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19765) );
  AOI22_X1 U19554 ( .A1(n16515), .A2(n18731), .B1(n19765), .B2(n16516), .ZN(
        U350) );
  INV_X1 U19555 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18729) );
  INV_X1 U19556 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19763) );
  AOI22_X1 U19557 ( .A1(n16515), .A2(n18729), .B1(n19763), .B2(n16516), .ZN(
        U351) );
  INV_X1 U19558 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18726) );
  INV_X1 U19559 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19761) );
  AOI22_X1 U19560 ( .A1(n16515), .A2(n18726), .B1(n19761), .B2(n16516), .ZN(
        U352) );
  INV_X1 U19561 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18725) );
  INV_X1 U19562 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19759) );
  AOI22_X1 U19563 ( .A1(n16515), .A2(n18725), .B1(n19759), .B2(n16516), .ZN(
        U353) );
  INV_X1 U19564 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18723) );
  AOI22_X1 U19565 ( .A1(n16515), .A2(n18723), .B1(n19757), .B2(n16516), .ZN(
        U354) );
  INV_X1 U19566 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18779) );
  INV_X1 U19567 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19807) );
  AOI22_X1 U19568 ( .A1(n16515), .A2(n18779), .B1(n19807), .B2(n16516), .ZN(
        U355) );
  INV_X1 U19569 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18776) );
  INV_X1 U19570 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19804) );
  AOI22_X1 U19571 ( .A1(n16515), .A2(n18776), .B1(n19804), .B2(n16516), .ZN(
        U356) );
  INV_X1 U19572 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18773) );
  INV_X1 U19573 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19802) );
  AOI22_X1 U19574 ( .A1(n16515), .A2(n18773), .B1(n19802), .B2(n16516), .ZN(
        U357) );
  INV_X1 U19575 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18772) );
  INV_X1 U19576 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19800) );
  AOI22_X1 U19577 ( .A1(n16515), .A2(n18772), .B1(n19800), .B2(n16516), .ZN(
        U358) );
  INV_X1 U19578 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18769) );
  INV_X1 U19579 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19799) );
  AOI22_X1 U19580 ( .A1(n16515), .A2(n18769), .B1(n19799), .B2(n16516), .ZN(
        U359) );
  INV_X1 U19581 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18767) );
  INV_X1 U19582 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19798) );
  AOI22_X1 U19583 ( .A1(n16515), .A2(n18767), .B1(n19798), .B2(n16516), .ZN(
        U360) );
  INV_X1 U19584 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18765) );
  INV_X1 U19585 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19796) );
  AOI22_X1 U19586 ( .A1(n16515), .A2(n18765), .B1(n19796), .B2(n16516), .ZN(
        U361) );
  INV_X1 U19587 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18762) );
  INV_X1 U19588 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19795) );
  AOI22_X1 U19589 ( .A1(n16515), .A2(n18762), .B1(n19795), .B2(n16516), .ZN(
        U362) );
  INV_X1 U19590 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18761) );
  INV_X1 U19591 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19793) );
  AOI22_X1 U19592 ( .A1(n16515), .A2(n18761), .B1(n19793), .B2(n16516), .ZN(
        U363) );
  INV_X1 U19593 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18758) );
  INV_X1 U19594 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19791) );
  AOI22_X1 U19595 ( .A1(n16515), .A2(n18758), .B1(n19791), .B2(n16516), .ZN(
        U364) );
  INV_X1 U19596 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18722) );
  INV_X1 U19597 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19755) );
  AOI22_X1 U19598 ( .A1(n16515), .A2(n18722), .B1(n19755), .B2(n16516), .ZN(
        U365) );
  INV_X1 U19599 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18757) );
  INV_X1 U19600 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n21075) );
  AOI22_X1 U19601 ( .A1(n16515), .A2(n18757), .B1(n21075), .B2(n16516), .ZN(
        U366) );
  INV_X1 U19602 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18755) );
  INV_X1 U19603 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19788) );
  AOI22_X1 U19604 ( .A1(n16515), .A2(n18755), .B1(n19788), .B2(n16516), .ZN(
        U367) );
  INV_X1 U19605 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18753) );
  INV_X1 U19606 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19786) );
  AOI22_X1 U19607 ( .A1(n16515), .A2(n18753), .B1(n19786), .B2(n16516), .ZN(
        U368) );
  INV_X1 U19608 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18751) );
  INV_X1 U19609 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19785) );
  AOI22_X1 U19610 ( .A1(n16515), .A2(n18751), .B1(n19785), .B2(n16516), .ZN(
        U369) );
  INV_X1 U19611 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18749) );
  INV_X1 U19612 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19783) );
  AOI22_X1 U19613 ( .A1(n16515), .A2(n18749), .B1(n19783), .B2(n16516), .ZN(
        U370) );
  INV_X1 U19614 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18747) );
  INV_X1 U19615 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19781) );
  AOI22_X1 U19616 ( .A1(n16515), .A2(n18747), .B1(n19781), .B2(n16516), .ZN(
        U371) );
  INV_X1 U19617 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18744) );
  INV_X1 U19618 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19779) );
  AOI22_X1 U19619 ( .A1(n16515), .A2(n18744), .B1(n19779), .B2(n16516), .ZN(
        U372) );
  INV_X1 U19620 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18743) );
  INV_X1 U19621 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19777) );
  AOI22_X1 U19622 ( .A1(n16515), .A2(n18743), .B1(n19777), .B2(n16516), .ZN(
        U373) );
  INV_X1 U19623 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18741) );
  INV_X1 U19624 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19775) );
  AOI22_X1 U19625 ( .A1(n16515), .A2(n18741), .B1(n19775), .B2(n16516), .ZN(
        U374) );
  INV_X1 U19626 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18739) );
  INV_X1 U19627 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19773) );
  AOI22_X1 U19628 ( .A1(n16515), .A2(n18739), .B1(n19773), .B2(n16516), .ZN(
        U375) );
  INV_X1 U19629 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18719) );
  INV_X1 U19630 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19754) );
  AOI22_X1 U19631 ( .A1(n16515), .A2(n18719), .B1(n19754), .B2(n16516), .ZN(
        U376) );
  NAND2_X1 U19632 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18718), .ZN(n18707) );
  AOI22_X1 U19633 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18707), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18710), .ZN(n18787) );
  AOI21_X1 U19634 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18787), .ZN(n16517) );
  INV_X1 U19635 ( .A(n16517), .ZN(P3_U2633) );
  OAI21_X1 U19636 ( .B1(n16523), .B2(n17378), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16518) );
  OAI21_X1 U19637 ( .B1(n16519), .B2(n18693), .A(n16518), .ZN(P3_U2634) );
  INV_X2 U19638 ( .A(n18849), .ZN(n18778) );
  AOI21_X1 U19639 ( .B1(n18710), .B2(n18718), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16520) );
  AOI22_X1 U19640 ( .A1(n18778), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16520), 
        .B2(n18849), .ZN(P3_U2635) );
  OAI21_X1 U19641 ( .B1(n18704), .B2(BS16), .A(n18787), .ZN(n18785) );
  OAI21_X1 U19642 ( .B1(n18787), .B2(n16542), .A(n18785), .ZN(P3_U2636) );
  INV_X1 U19643 ( .A(n16521), .ZN(n16522) );
  NOR3_X1 U19644 ( .A1(n16523), .A2(n18623), .A3(n16522), .ZN(n18629) );
  NOR2_X1 U19645 ( .A1(n18629), .A2(n18690), .ZN(n18832) );
  OAI21_X1 U19646 ( .B1(n18832), .B2(n18178), .A(n16524), .ZN(P3_U2637) );
  NOR4_X1 U19647 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16528) );
  NOR4_X1 U19648 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16527) );
  NOR4_X1 U19649 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16526) );
  NOR4_X1 U19650 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16525) );
  NAND4_X1 U19651 ( .A1(n16528), .A2(n16527), .A3(n16526), .A4(n16525), .ZN(
        n16534) );
  NOR4_X1 U19652 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16532) );
  AOI211_X1 U19653 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_25__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16531) );
  NOR4_X1 U19654 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16530) );
  NOR4_X1 U19655 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16529) );
  NAND4_X1 U19656 ( .A1(n16532), .A2(n16531), .A3(n16530), .A4(n16529), .ZN(
        n16533) );
  NOR2_X1 U19657 ( .A1(n16534), .A2(n16533), .ZN(n18822) );
  INV_X1 U19658 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16536) );
  INV_X1 U19659 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18786) );
  NAND2_X1 U19660 ( .A1(n18822), .A2(n18786), .ZN(n18823) );
  NOR3_X1 U19661 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A3(n18823), .ZN(n16537) );
  INV_X1 U19662 ( .A(n16537), .ZN(n16535) );
  NAND2_X1 U19663 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18822), .ZN(n18826) );
  OAI211_X1 U19664 ( .C1(n18822), .C2(n16536), .A(n16535), .B(n18826), .ZN(
        P3_U2638) );
  NOR2_X1 U19665 ( .A1(n16537), .A2(n18826), .ZN(n16539) );
  NOR2_X1 U19666 ( .A1(P3_BYTEENABLE_REG_3__SCAN_IN), .A2(n18822), .ZN(n16538)
         );
  AOI211_X1 U19667 ( .C1(n18822), .C2(P3_DATAWIDTH_REG_1__SCAN_IN), .A(n16539), 
        .B(n16538), .ZN(P3_U2639) );
  NAND2_X1 U19668 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18840), .ZN(n16541) );
  AOI211_X4 U19669 ( .C1(n16542), .C2(n18834), .A(n16543), .B(n16541), .ZN(
        n16883) );
  NOR3_X1 U19670 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16892) );
  INV_X1 U19671 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17200) );
  NAND2_X1 U19672 ( .A1(n16892), .A2(n17200), .ZN(n16882) );
  NOR2_X1 U19673 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16882), .ZN(n16858) );
  NAND2_X1 U19674 ( .A1(n16858), .A2(n16853), .ZN(n16852) );
  NAND2_X1 U19675 ( .A1(n16841), .A2(n17191), .ZN(n16829) );
  NAND2_X1 U19676 ( .A1(n16811), .A2(n16808), .ZN(n16807) );
  INV_X1 U19677 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16785) );
  NAND2_X1 U19678 ( .A1(n16788), .A2(n16785), .ZN(n16777) );
  NAND2_X1 U19679 ( .A1(n16761), .A2(n16756), .ZN(n16755) );
  INV_X1 U19680 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16731) );
  NAND2_X1 U19681 ( .A1(n16735), .A2(n16731), .ZN(n16730) );
  INV_X1 U19682 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17062) );
  NAND2_X1 U19683 ( .A1(n16712), .A2(n17062), .ZN(n16708) );
  INV_X1 U19684 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16681) );
  NAND2_X1 U19685 ( .A1(n16688), .A2(n16681), .ZN(n16679) );
  NAND2_X1 U19686 ( .A1(n16667), .A2(n16661), .ZN(n16663) );
  NAND2_X1 U19687 ( .A1(n16643), .A2(n16639), .ZN(n16638) );
  NAND2_X1 U19688 ( .A1(n16626), .A2(n16620), .ZN(n16619) );
  NOR2_X1 U19689 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16619), .ZN(n16604) );
  NAND2_X1 U19690 ( .A1(n16604), .A2(n16598), .ZN(n16597) );
  INV_X1 U19691 ( .A(n16597), .ZN(n16586) );
  NAND2_X1 U19692 ( .A1(n16585), .A2(n16586), .ZN(n16584) );
  NOR2_X1 U19693 ( .A1(n16913), .A2(n16562), .ZN(n16568) );
  INV_X1 U19694 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n21042) );
  INV_X1 U19695 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18780) );
  OAI211_X1 U19696 ( .C1(n18840), .C2(n18839), .A(n18834), .B(n16542), .ZN(
        n18682) );
  INV_X1 U19697 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18766) );
  INV_X1 U19698 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18763) );
  INV_X1 U19699 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18742) );
  INV_X1 U19700 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18738) );
  INV_X1 U19701 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18734) );
  NAND3_X1 U19702 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16857) );
  NAND2_X1 U19703 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(P3_REIP_REG_4__SCAN_IN), 
        .ZN(n16794) );
  NOR2_X1 U19704 ( .A1(n16857), .A2(n16794), .ZN(n16813) );
  NAND4_X1 U19705 ( .A1(n16813), .A2(P3_REIP_REG_8__SCAN_IN), .A3(
        P3_REIP_REG_7__SCAN_IN), .A4(P3_REIP_REG_6__SCAN_IN), .ZN(n16793) );
  NOR2_X1 U19706 ( .A1(n18734), .A2(n16793), .ZN(n16787) );
  NAND2_X1 U19707 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n16787), .ZN(n16771) );
  NOR2_X1 U19708 ( .A1(n18738), .A2(n16771), .ZN(n16764) );
  NAND2_X1 U19709 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16764), .ZN(n16748) );
  NOR2_X1 U19710 ( .A1(n18742), .A2(n16748), .ZN(n16736) );
  NAND2_X1 U19711 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16736), .ZN(n16647) );
  INV_X1 U19712 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18750) );
  NAND2_X1 U19713 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16715) );
  NOR2_X1 U19714 ( .A1(n18750), .A2(n16715), .ZN(n16684) );
  NAND4_X1 U19715 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(P3_REIP_REG_19__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .A4(n16684), .ZN(n16646) );
  NAND2_X1 U19716 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .ZN(n16649) );
  NOR4_X1 U19717 ( .A1(n18763), .A2(n16647), .A3(n16646), .A4(n16649), .ZN(
        n16625) );
  NAND2_X1 U19718 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16625), .ZN(n16616) );
  NOR2_X1 U19719 ( .A1(n18766), .A2(n16616), .ZN(n16603) );
  NAND2_X1 U19720 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16603), .ZN(n16550) );
  NOR2_X1 U19721 ( .A1(n16904), .A2(n16550), .ZN(n16587) );
  NAND4_X1 U19722 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16587), .ZN(n16549) );
  NOR3_X1 U19723 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18780), .A3(n16549), 
        .ZN(n16548) );
  NAND4_X1 U19724 ( .A1(n18851), .A2(n18843), .A3(n16542), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n18698) );
  NAND2_X1 U19725 ( .A1(n18851), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18560) );
  NOR2_X1 U19726 ( .A1(n18693), .A2(n18560), .ZN(n18687) );
  NOR4_X4 U19727 ( .A1(n9654), .A2(n18854), .A3(n16881), .A4(n18687), .ZN(
        n16912) );
  INV_X1 U19728 ( .A(P3_EBX_REG_31__SCAN_IN), .ZN(n16545) );
  INV_X1 U19729 ( .A(n16543), .ZN(n16544) );
  OAI211_X2 U19730 ( .C1(n16545), .C2(n18192), .A(n18682), .B(n16544), .ZN(
        n16914) );
  OAI22_X1 U19731 ( .A1(n16546), .A2(n16894), .B1(n16545), .B2(n16914), .ZN(
        n16547) );
  AOI211_X1 U19732 ( .C1(n16568), .C2(n21042), .A(n16548), .B(n16547), .ZN(
        n16561) );
  NOR2_X1 U19733 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16549), .ZN(n16567) );
  NAND3_X1 U19734 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16551) );
  AND2_X1 U19735 ( .A1(n16873), .A2(n16550), .ZN(n16602) );
  NOR2_X1 U19736 ( .A1(n16912), .A2(n16602), .ZN(n16601) );
  INV_X1 U19737 ( .A(n16601), .ZN(n16609) );
  AOI21_X1 U19738 ( .B1(n16873), .B2(n16551), .A(n16609), .ZN(n16565) );
  INV_X1 U19739 ( .A(n16565), .ZN(n16577) );
  OAI21_X1 U19740 ( .B1(n16567), .B2(n16577), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n16560) );
  INV_X1 U19741 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17495) );
  NOR2_X1 U19742 ( .A1(n16554), .A2(n17495), .ZN(n16553) );
  OAI21_X1 U19743 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n16553), .A(
        n16552), .ZN(n17510) );
  INV_X1 U19744 ( .A(n17510), .ZN(n16582) );
  AOI21_X1 U19745 ( .B1(n16554), .B2(n17495), .A(n16553), .ZN(n17511) );
  INV_X1 U19746 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16612) );
  NAND2_X1 U19747 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17524), .ZN(
        n17491) );
  AOI21_X1 U19748 ( .B1(n16612), .B2(n17491), .A(n9900), .ZN(n17528) );
  INV_X1 U19749 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17549) );
  INV_X1 U19750 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16652) );
  INV_X1 U19751 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17851) );
  NOR2_X1 U19752 ( .A1(n17851), .A2(n17612), .ZN(n17611) );
  INV_X1 U19753 ( .A(n17611), .ZN(n16699) );
  NOR2_X1 U19754 ( .A1(n17613), .A2(n16699), .ZN(n17573) );
  INV_X1 U19755 ( .A(n17573), .ZN(n16676) );
  NOR2_X1 U19756 ( .A1(n9895), .A2(n16676), .ZN(n16558) );
  NAND2_X1 U19757 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16558), .ZN(
        n16557) );
  NOR2_X1 U19758 ( .A1(n16652), .A2(n16557), .ZN(n17533) );
  NAND2_X1 U19759 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17533), .ZN(
        n16556) );
  NOR2_X1 U19760 ( .A1(n17549), .A2(n16556), .ZN(n16555) );
  OAI21_X1 U19761 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16555), .A(
        n17491), .ZN(n17538) );
  INV_X1 U19762 ( .A(n17538), .ZN(n16614) );
  AOI21_X1 U19763 ( .B1(n17549), .B2(n16556), .A(n16555), .ZN(n17547) );
  OAI21_X1 U19764 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17533), .A(
        n16556), .ZN(n17558) );
  INV_X1 U19765 ( .A(n17558), .ZN(n16634) );
  AOI21_X1 U19766 ( .B1(n16652), .B2(n16557), .A(n17533), .ZN(n17575) );
  OAI21_X1 U19767 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n16558), .A(
        n16557), .ZN(n17587) );
  INV_X1 U19768 ( .A(n17587), .ZN(n16658) );
  AOI21_X1 U19769 ( .B1(n9895), .B2(n16676), .A(n16558), .ZN(n17604) );
  NOR2_X1 U19770 ( .A1(n17851), .A2(n17650), .ZN(n17649) );
  NAND2_X1 U19771 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17649), .ZN(
        n16724) );
  NOR2_X1 U19772 ( .A1(n16724), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16691) );
  INV_X1 U19773 ( .A(n16691), .ZN(n16729) );
  NAND2_X1 U19774 ( .A1(n16872), .A2(n16729), .ZN(n16717) );
  OAI21_X1 U19775 ( .B1(n17573), .B2(n16835), .A(n16717), .ZN(n16670) );
  NOR2_X1 U19776 ( .A1(n17604), .A2(n16670), .ZN(n16669) );
  NOR2_X1 U19777 ( .A1(n16669), .A2(n16835), .ZN(n16657) );
  NOR2_X1 U19778 ( .A1(n16634), .A2(n9700), .ZN(n16633) );
  NOR2_X1 U19779 ( .A1(n16633), .A2(n16835), .ZN(n16628) );
  NOR2_X1 U19780 ( .A1(n17528), .A2(n16606), .ZN(n16605) );
  NOR2_X1 U19781 ( .A1(n16581), .A2(n16835), .ZN(n16573) );
  NOR2_X1 U19782 ( .A1(n16574), .A2(n16573), .ZN(n16572) );
  NAND4_X1 U19783 ( .A1(n16872), .A2(n16881), .A3(n16572), .A4(n16563), .ZN(
        n16559) );
  NAND3_X1 U19784 ( .A1(n16561), .A2(n16560), .A3(n16559), .ZN(P3_U2640) );
  NAND2_X1 U19785 ( .A1(n16883), .A2(n16562), .ZN(n16571) );
  OAI22_X1 U19786 ( .A1(n16565), .A2(n18780), .B1(n16564), .B2(n16894), .ZN(
        n16566) );
  OAI21_X1 U19787 ( .B1(n16875), .B2(n16568), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16569) );
  INV_X1 U19788 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18771) );
  NOR3_X1 U19789 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n18774), .A3(n18771), 
        .ZN(n16570) );
  AOI22_X1 U19790 ( .A1(n16875), .A2(P3_EBX_REG_29__SCAN_IN), .B1(n16587), 
        .B2(n16570), .ZN(n16579) );
  AOI21_X1 U19791 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16584), .A(n16571), .ZN(
        n16576) );
  AOI211_X1 U19792 ( .C1(n16574), .C2(n16573), .A(n16572), .B(n18698), .ZN(
        n16575) );
  AOI211_X1 U19793 ( .C1(P3_REIP_REG_29__SCAN_IN), .C2(n16577), .A(n16576), 
        .B(n16575), .ZN(n16578) );
  OAI211_X1 U19794 ( .C1(n16580), .C2(n16894), .A(n16579), .B(n16578), .ZN(
        P3_U2642) );
  AOI22_X1 U19795 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16902), .B1(
        n16875), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16591) );
  AND2_X1 U19796 ( .A1(n18771), .A2(n16587), .ZN(n16596) );
  AOI211_X1 U19797 ( .C1(n16582), .C2(n9885), .A(n16581), .B(n18698), .ZN(
        n16583) );
  AOI221_X1 U19798 ( .B1(n16596), .B2(P3_REIP_REG_28__SCAN_IN), .C1(n16609), 
        .C2(P3_REIP_REG_28__SCAN_IN), .A(n16583), .ZN(n16590) );
  OAI211_X1 U19799 ( .C1(n16586), .C2(n16585), .A(n16883), .B(n16584), .ZN(
        n16589) );
  NAND3_X1 U19800 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16587), .A3(n18774), 
        .ZN(n16588) );
  NAND4_X1 U19801 ( .A1(n16591), .A2(n16590), .A3(n16589), .A4(n16588), .ZN(
        P3_U2643) );
  AOI211_X1 U19802 ( .C1(n17511), .C2(n16593), .A(n16592), .B(n18698), .ZN(
        n16595) );
  OAI22_X1 U19803 ( .A1(n17495), .A2(n16894), .B1(n16914), .B2(n16598), .ZN(
        n16594) );
  NOR3_X1 U19804 ( .A1(n16596), .A2(n16595), .A3(n16594), .ZN(n16600) );
  OAI211_X1 U19805 ( .C1(n16604), .C2(n16598), .A(n16883), .B(n16597), .ZN(
        n16599) );
  OAI211_X1 U19806 ( .C1(n16601), .C2(n18771), .A(n16600), .B(n16599), .ZN(
        P3_U2644) );
  AOI22_X1 U19807 ( .A1(n16875), .A2(P3_EBX_REG_26__SCAN_IN), .B1(n16603), 
        .B2(n16602), .ZN(n16611) );
  AOI211_X1 U19808 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16619), .A(n16604), .B(
        n16913), .ZN(n16608) );
  AOI211_X1 U19809 ( .C1(n17528), .C2(n16606), .A(n16605), .B(n18698), .ZN(
        n16607) );
  AOI211_X1 U19810 ( .C1(P3_REIP_REG_26__SCAN_IN), .C2(n16609), .A(n16608), 
        .B(n16607), .ZN(n16610) );
  OAI211_X1 U19811 ( .C1(n16612), .C2(n16894), .A(n16611), .B(n16610), .ZN(
        P3_U2645) );
  INV_X1 U19812 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18764) );
  INV_X1 U19813 ( .A(n16912), .ZN(n16753) );
  OAI21_X1 U19814 ( .B1(n16625), .B2(n16904), .A(n16753), .ZN(n16637) );
  AOI21_X1 U19815 ( .B1(n16873), .B2(n18764), .A(n16637), .ZN(n16623) );
  AOI211_X1 U19816 ( .C1(n16614), .C2(n16613), .A(n9770), .B(n18698), .ZN(
        n16618) );
  NAND2_X1 U19817 ( .A1(n16873), .A2(n18766), .ZN(n16615) );
  OAI22_X1 U19818 ( .A1(n16914), .A2(n16620), .B1(n16616), .B2(n16615), .ZN(
        n16617) );
  AOI211_X1 U19819 ( .C1(n16902), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16618), .B(n16617), .ZN(n16622) );
  OAI211_X1 U19820 ( .C1(n16626), .C2(n16620), .A(n16883), .B(n16619), .ZN(
        n16621) );
  OAI211_X1 U19821 ( .C1(n16623), .C2(n18766), .A(n16622), .B(n16621), .ZN(
        P3_U2646) );
  NOR2_X1 U19822 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16904), .ZN(n16624) );
  AOI22_X1 U19823 ( .A1(n16875), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16625), 
        .B2(n16624), .ZN(n16632) );
  AOI211_X1 U19824 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16638), .A(n16626), .B(
        n16913), .ZN(n16630) );
  AOI211_X1 U19825 ( .C1(n17547), .C2(n16628), .A(n16627), .B(n18698), .ZN(
        n16629) );
  AOI211_X1 U19826 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16637), .A(n16630), 
        .B(n16629), .ZN(n16631) );
  OAI211_X1 U19827 ( .C1(n17549), .C2(n16894), .A(n16632), .B(n16631), .ZN(
        P3_U2647) );
  NAND3_X1 U19828 ( .A1(n16873), .A2(P3_REIP_REG_14__SCAN_IN), .A3(n16736), 
        .ZN(n16698) );
  NOR2_X1 U19829 ( .A1(n16646), .A2(n16698), .ZN(n16660) );
  NAND2_X1 U19830 ( .A1(n16660), .A2(n18763), .ZN(n16642) );
  AOI211_X1 U19831 ( .C1(n16634), .C2(n9700), .A(n16633), .B(n18698), .ZN(
        n16636) );
  INV_X1 U19832 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17559) );
  OAI22_X1 U19833 ( .A1(n17559), .A2(n16894), .B1(n16914), .B2(n16639), .ZN(
        n16635) );
  AOI211_X1 U19834 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n16637), .A(n16636), 
        .B(n16635), .ZN(n16641) );
  OAI211_X1 U19835 ( .C1(n16643), .C2(n16639), .A(n16883), .B(n16638), .ZN(
        n16640) );
  OAI211_X1 U19836 ( .C1(n16649), .C2(n16642), .A(n16641), .B(n16640), .ZN(
        P3_U2648) );
  AOI211_X1 U19837 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16663), .A(n16643), .B(
        n16913), .ZN(n16655) );
  AOI211_X1 U19838 ( .C1(n17575), .C2(n16645), .A(n16644), .B(n18698), .ZN(
        n16654) );
  INV_X1 U19839 ( .A(n16646), .ZN(n16648) );
  NOR2_X1 U19840 ( .A1(n16912), .A2(n16647), .ZN(n16714) );
  NAND2_X1 U19841 ( .A1(n16753), .A2(n16904), .ZN(n16917) );
  AOI21_X1 U19842 ( .B1(n16648), .B2(n16714), .A(n16823), .ZN(n16673) );
  AOI22_X1 U19843 ( .A1(n16875), .A2(P3_EBX_REG_22__SCAN_IN), .B1(
        P3_REIP_REG_22__SCAN_IN), .B2(n16673), .ZN(n16651) );
  OAI211_X1 U19844 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(P3_REIP_REG_22__SCAN_IN), .A(n16660), .B(n16649), .ZN(n16650) );
  OAI211_X1 U19845 ( .C1(n16894), .C2(n16652), .A(n16651), .B(n16650), .ZN(
        n16653) );
  OR3_X1 U19846 ( .A1(n16655), .A2(n16654), .A3(n16653), .ZN(P3_U2649) );
  INV_X1 U19847 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17590) );
  INV_X1 U19848 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18759) );
  AOI211_X1 U19849 ( .C1(n16658), .C2(n16657), .A(n16656), .B(n18698), .ZN(
        n16659) );
  AOI221_X1 U19850 ( .B1(n16673), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n16660), 
        .C2(n18759), .A(n16659), .ZN(n16666) );
  OAI21_X1 U19851 ( .B1(n16661), .B2(n16667), .A(n16883), .ZN(n16662) );
  INV_X1 U19852 ( .A(n16662), .ZN(n16664) );
  OAI221_X1 U19853 ( .B1(n16664), .B2(P3_EBX_REG_21__SCAN_IN), .C1(n16664), 
        .C2(n16875), .A(n16663), .ZN(n16665) );
  OAI211_X1 U19854 ( .C1(n16894), .C2(n17590), .A(n16666), .B(n16665), .ZN(
        P3_U2650) );
  AOI211_X1 U19855 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16679), .A(n16667), .B(
        n16913), .ZN(n16668) );
  AOI21_X1 U19856 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16875), .A(n16668), .ZN(
        n16675) );
  INV_X1 U19857 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18754) );
  INV_X1 U19858 ( .A(n16698), .ZN(n16728) );
  NAND3_X1 U19859 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16684), .A3(n16728), 
        .ZN(n16687) );
  NOR2_X1 U19860 ( .A1(n18754), .A2(n16687), .ZN(n16672) );
  INV_X1 U19861 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18756) );
  AOI211_X1 U19862 ( .C1(n17604), .C2(n16670), .A(n16669), .B(n18698), .ZN(
        n16671) );
  AOI221_X1 U19863 ( .B1(n16673), .B2(P3_REIP_REG_20__SCAN_IN), .C1(n16672), 
        .C2(n18756), .A(n16671), .ZN(n16674) );
  OAI211_X1 U19864 ( .C1(n9895), .C2(n16894), .A(n16675), .B(n16674), .ZN(
        P3_U2651) );
  NAND2_X1 U19865 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17611), .ZN(
        n16690) );
  OAI21_X1 U19866 ( .B1(n16690), .B2(n16729), .A(n16872), .ZN(n16693) );
  INV_X1 U19867 ( .A(n16690), .ZN(n16677) );
  OAI21_X1 U19868 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16677), .A(
        n16676), .ZN(n17615) );
  OAI21_X1 U19869 ( .B1(n16693), .B2(n17615), .A(n16881), .ZN(n16678) );
  AOI21_X1 U19870 ( .B1(n16693), .B2(n17615), .A(n16678), .ZN(n16683) );
  OAI211_X1 U19871 ( .C1(n16688), .C2(n16681), .A(n16883), .B(n16679), .ZN(
        n16680) );
  OAI211_X1 U19872 ( .C1(n16914), .C2(n16681), .A(n18077), .B(n16680), .ZN(
        n16682) );
  AOI211_X1 U19873 ( .C1(n16902), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16683), .B(n16682), .ZN(n16686) );
  AOI21_X1 U19874 ( .B1(n16684), .B2(n16714), .A(n16823), .ZN(n16707) );
  INV_X1 U19875 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18752) );
  AND3_X1 U19876 ( .A1(n18752), .A2(n16684), .A3(n16728), .ZN(n16695) );
  OAI21_X1 U19877 ( .B1(n16707), .B2(n16695), .A(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n16685) );
  OAI211_X1 U19878 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(n16687), .A(n16686), 
        .B(n16685), .ZN(P3_U2652) );
  INV_X1 U19879 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17627) );
  AOI211_X1 U19880 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16708), .A(n16688), .B(
        n16913), .ZN(n16689) );
  AOI211_X1 U19881 ( .C1(n16875), .C2(P3_EBX_REG_18__SCAN_IN), .A(n9654), .B(
        n16689), .ZN(n16697) );
  OAI21_X1 U19882 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17611), .A(
        n16690), .ZN(n17624) );
  NAND2_X1 U19883 ( .A1(n16881), .A2(n16835), .ZN(n16901) );
  OAI221_X1 U19884 ( .B1(n17624), .B2(n16691), .C1(n17624), .C2(n17627), .A(
        n16881), .ZN(n16692) );
  AOI22_X1 U19885 ( .A1(n16693), .A2(n17624), .B1(n16901), .B2(n16692), .ZN(
        n16694) );
  AOI211_X1 U19886 ( .C1(n16707), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16695), 
        .B(n16694), .ZN(n16696) );
  OAI211_X1 U19887 ( .C1(n17627), .C2(n16894), .A(n16697), .B(n16696), .ZN(
        P3_U2653) );
  AOI22_X1 U19888 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16902), .B1(
        n16875), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16711) );
  NOR2_X1 U19889 ( .A1(n16715), .A2(n16698), .ZN(n16706) );
  INV_X1 U19890 ( .A(n17649), .ZN(n16740) );
  NOR2_X1 U19891 ( .A1(n17651), .A2(n16740), .ZN(n16700) );
  OAI21_X1 U19892 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16700), .A(
        n16699), .ZN(n17644) );
  INV_X1 U19893 ( .A(n16724), .ZN(n16702) );
  INV_X1 U19894 ( .A(n16700), .ZN(n16701) );
  OAI21_X1 U19895 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16702), .A(
        n16701), .ZN(n17654) );
  NAND2_X1 U19896 ( .A1(n16717), .A2(n17654), .ZN(n16716) );
  NAND2_X1 U19897 ( .A1(n16872), .A2(n16716), .ZN(n16704) );
  OAI21_X1 U19898 ( .B1(n17644), .B2(n16704), .A(n16881), .ZN(n16703) );
  AOI21_X1 U19899 ( .B1(n17644), .B2(n16704), .A(n16703), .ZN(n16705) );
  AOI221_X1 U19900 ( .B1(n16707), .B2(P3_REIP_REG_17__SCAN_IN), .C1(n16706), 
        .C2(n18750), .A(n16705), .ZN(n16710) );
  OAI211_X1 U19901 ( .C1(n16712), .C2(n17062), .A(n16883), .B(n16708), .ZN(
        n16709) );
  NAND4_X1 U19902 ( .A1(n16711), .A2(n16710), .A3(n18077), .A4(n16709), .ZN(
        P3_U2654) );
  AOI211_X1 U19903 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16730), .A(n16712), .B(
        n16913), .ZN(n16713) );
  AOI211_X1 U19904 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n16902), .A(
        n9654), .B(n16713), .ZN(n16722) );
  NOR2_X1 U19905 ( .A1(n16823), .A2(n16714), .ZN(n16737) );
  OAI211_X1 U19906 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16728), .B(n16715), .ZN(n16719) );
  OAI211_X1 U19907 ( .C1(n16717), .C2(n17654), .A(n16881), .B(n16716), .ZN(
        n16718) );
  NAND2_X1 U19908 ( .A1(n16719), .A2(n16718), .ZN(n16720) );
  AOI21_X1 U19909 ( .B1(P3_REIP_REG_16__SCAN_IN), .B2(n16737), .A(n16720), 
        .ZN(n16721) );
  OAI211_X1 U19910 ( .C1(n16914), .C2(n16723), .A(n16722), .B(n16721), .ZN(
        P3_U2655) );
  INV_X1 U19911 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18746) );
  OAI21_X1 U19912 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17649), .A(
        n16724), .ZN(n17659) );
  INV_X1 U19913 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16911) );
  OAI21_X1 U19914 ( .B1(n16835), .B2(n16911), .A(n16881), .ZN(n16910) );
  AOI211_X1 U19915 ( .C1(n16872), .C2(n16740), .A(n17659), .B(n16910), .ZN(
        n16725) );
  AOI21_X1 U19916 ( .B1(n16902), .B2(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16725), .ZN(n16726) );
  OAI21_X1 U19917 ( .B1(n16914), .B2(n16731), .A(n16726), .ZN(n16727) );
  AOI221_X1 U19918 ( .B1(n16737), .B2(P3_REIP_REG_15__SCAN_IN), .C1(n16728), 
        .C2(n18746), .A(n16727), .ZN(n16734) );
  NOR2_X1 U19919 ( .A1(n16835), .A2(n18698), .ZN(n16903) );
  NAND3_X1 U19920 ( .A1(n16903), .A2(n16729), .A3(n17659), .ZN(n16733) );
  OAI211_X1 U19921 ( .C1(n16735), .C2(n16731), .A(n16883), .B(n16730), .ZN(
        n16732) );
  NAND4_X1 U19922 ( .A1(n16734), .A2(n18077), .A3(n16733), .A4(n16732), .ZN(
        P3_U2656) );
  AOI211_X1 U19923 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16755), .A(n16735), .B(
        n16913), .ZN(n16746) );
  AOI21_X1 U19924 ( .B1(n16873), .B2(n16736), .A(P3_REIP_REG_14__SCAN_IN), 
        .ZN(n16744) );
  INV_X1 U19925 ( .A(n16737), .ZN(n16743) );
  NOR2_X1 U19926 ( .A1(n17851), .A2(n16738), .ZN(n16847) );
  NAND2_X1 U19927 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16847), .ZN(
        n16833) );
  INV_X1 U19928 ( .A(n16833), .ZN(n16825) );
  NAND2_X1 U19929 ( .A1(n17690), .A2(n16825), .ZN(n17686) );
  OAI21_X1 U19930 ( .B1(n17686), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n16872), .ZN(n16766) );
  INV_X1 U19931 ( .A(n16766), .ZN(n16739) );
  AOI21_X1 U19932 ( .B1(n16872), .B2(n17692), .A(n16739), .ZN(n16750) );
  NAND2_X1 U19933 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17674), .ZN(
        n16751) );
  INV_X1 U19934 ( .A(n16751), .ZN(n16741) );
  OAI21_X1 U19935 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16741), .A(
        n16740), .ZN(n17675) );
  XNOR2_X1 U19936 ( .A(n16750), .B(n17675), .ZN(n16742) );
  OAI22_X1 U19937 ( .A1(n16744), .A2(n16743), .B1(n18698), .B2(n16742), .ZN(
        n16745) );
  AOI211_X1 U19938 ( .C1(n16902), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16746), .B(n16745), .ZN(n16747) );
  OAI211_X1 U19939 ( .C1(n16914), .C2(n17106), .A(n16747), .B(n18077), .ZN(
        P3_U2657) );
  NOR3_X1 U19940 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16904), .A3(n16748), 
        .ZN(n16749) );
  AOI211_X1 U19941 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n16902), .A(
        n9654), .B(n16749), .ZN(n16760) );
  NOR2_X1 U19942 ( .A1(n16750), .A2(n18698), .ZN(n16752) );
  INV_X1 U19943 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17714) );
  NOR2_X1 U19944 ( .A1(n17714), .A2(n17686), .ZN(n16765) );
  OAI21_X1 U19945 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16765), .A(
        n16751), .ZN(n17695) );
  AOI22_X1 U19946 ( .A1(n16875), .A2(P3_EBX_REG_13__SCAN_IN), .B1(n16752), 
        .B2(n17695), .ZN(n16759) );
  OAI21_X1 U19947 ( .B1(n16764), .B2(n16904), .A(n16753), .ZN(n16783) );
  NOR2_X1 U19948 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16904), .ZN(n16763) );
  AOI211_X1 U19949 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n16872), .A(
        n17695), .B(n16910), .ZN(n16754) );
  AOI221_X1 U19950 ( .B1(n16783), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n16763), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n16754), .ZN(n16758) );
  OAI211_X1 U19951 ( .C1(n16761), .C2(n16756), .A(n16883), .B(n16755), .ZN(
        n16757) );
  NAND4_X1 U19952 ( .A1(n16760), .A2(n16759), .A3(n16758), .A4(n16757), .ZN(
        P3_U2658) );
  AOI22_X1 U19953 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16902), .B1(
        n16875), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n16770) );
  AOI211_X1 U19954 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16777), .A(n16761), .B(
        n16913), .ZN(n16762) );
  AOI211_X1 U19955 ( .C1(n16764), .C2(n16763), .A(n9654), .B(n16762), .ZN(
        n16769) );
  AOI21_X1 U19956 ( .B1(n17714), .B2(n17686), .A(n16765), .ZN(n17705) );
  XNOR2_X1 U19957 ( .A(n17705), .B(n16766), .ZN(n16767) );
  AOI22_X1 U19958 ( .A1(n16881), .A2(n16767), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n16783), .ZN(n16768) );
  NAND3_X1 U19959 ( .A1(n16770), .A2(n16769), .A3(n16768), .ZN(P3_U2659) );
  OAI21_X1 U19960 ( .B1(n16904), .B2(n16771), .A(n18738), .ZN(n16782) );
  INV_X1 U19961 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16780) );
  INV_X1 U19962 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17733) );
  NAND2_X1 U19963 ( .A1(n17775), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16772) );
  NOR2_X1 U19964 ( .A1(n17851), .A2(n16772), .ZN(n16773) );
  INV_X1 U19965 ( .A(n16773), .ZN(n16824) );
  NOR2_X1 U19966 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16824), .ZN(
        n16815) );
  AOI21_X1 U19967 ( .B1(n16774), .B2(n16815), .A(n16835), .ZN(n16792) );
  AOI21_X1 U19968 ( .B1(n16872), .B2(n17733), .A(n16792), .ZN(n16776) );
  NAND2_X1 U19969 ( .A1(n16774), .A2(n16773), .ZN(n16800) );
  NOR2_X1 U19970 ( .A1(n17733), .A2(n16800), .ZN(n16790) );
  OAI21_X1 U19971 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16790), .A(
        n17686), .ZN(n17722) );
  AOI21_X1 U19972 ( .B1(n16776), .B2(n17722), .A(n18698), .ZN(n16775) );
  OAI21_X1 U19973 ( .B1(n16776), .B2(n17722), .A(n16775), .ZN(n16779) );
  OAI211_X1 U19974 ( .C1(n16788), .C2(n16785), .A(n16883), .B(n16777), .ZN(
        n16778) );
  OAI211_X1 U19975 ( .C1(n16894), .C2(n16780), .A(n16779), .B(n16778), .ZN(
        n16781) );
  AOI21_X1 U19976 ( .B1(n16783), .B2(n16782), .A(n16781), .ZN(n16784) );
  OAI211_X1 U19977 ( .C1(n16914), .C2(n16785), .A(n16784), .B(n18077), .ZN(
        P3_U2660) );
  NOR2_X1 U19978 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(n16904), .ZN(n16786) );
  AOI22_X1 U19979 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n16902), .B1(
        n16787), .B2(n16786), .ZN(n16799) );
  AOI211_X1 U19980 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16807), .A(n16788), .B(
        n16913), .ZN(n16789) );
  AOI211_X1 U19981 ( .C1(n16875), .C2(P3_EBX_REG_10__SCAN_IN), .A(n9654), .B(
        n16789), .ZN(n16798) );
  AOI21_X1 U19982 ( .B1(n17733), .B2(n16800), .A(n16790), .ZN(n17736) );
  INV_X1 U19983 ( .A(n17736), .ZN(n16791) );
  INV_X1 U19984 ( .A(n16792), .ZN(n16802) );
  OAI221_X1 U19985 ( .B1(n17736), .B2(n16792), .C1(n16791), .C2(n16802), .A(
        n16881), .ZN(n16797) );
  NOR3_X1 U19986 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16904), .A3(n16793), .ZN(
        n16803) );
  INV_X1 U19987 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18732) );
  INV_X1 U19988 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18730) );
  INV_X1 U19989 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18728) );
  NOR3_X1 U19990 ( .A1(n18732), .A2(n18730), .A3(n18728), .ZN(n16795) );
  AOI221_X1 U19991 ( .B1(n16857), .B2(n16873), .C1(n16794), .C2(n16873), .A(
        n16912), .ZN(n16849) );
  OAI21_X1 U19992 ( .B1(n16795), .B2(n16823), .A(n16849), .ZN(n16812) );
  OAI21_X1 U19993 ( .B1(n16803), .B2(n16812), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n16796) );
  NAND4_X1 U19994 ( .A1(n16799), .A2(n16798), .A3(n16797), .A4(n16796), .ZN(
        P3_U2661) );
  NOR2_X1 U19995 ( .A1(n17761), .A2(n16824), .ZN(n16814) );
  OAI21_X1 U19996 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16814), .A(
        n16800), .ZN(n17748) );
  OAI221_X1 U19997 ( .B1(n17748), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C1(
        n17748), .C2(n16815), .A(n16881), .ZN(n16801) );
  AOI22_X1 U19998 ( .A1(n17748), .A2(n16802), .B1(n16901), .B2(n16801), .ZN(
        n16806) );
  AOI211_X1 U19999 ( .C1(n16875), .C2(P3_EBX_REG_9__SCAN_IN), .A(n9654), .B(
        n16803), .ZN(n16804) );
  INV_X1 U20000 ( .A(n16804), .ZN(n16805) );
  AOI211_X1 U20001 ( .C1(P3_REIP_REG_9__SCAN_IN), .C2(n16812), .A(n16806), .B(
        n16805), .ZN(n16810) );
  OAI211_X1 U20002 ( .C1(n16811), .C2(n16808), .A(n16883), .B(n16807), .ZN(
        n16809) );
  OAI211_X1 U20003 ( .C1(n16894), .C2(n21064), .A(n16810), .B(n16809), .ZN(
        P3_U2662) );
  AOI211_X1 U20004 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16829), .A(n16811), .B(
        n16913), .ZN(n16821) );
  INV_X1 U20005 ( .A(n16812), .ZN(n16819) );
  NAND2_X1 U20006 ( .A1(n16873), .A2(n16813), .ZN(n16840) );
  NOR2_X1 U20007 ( .A1(n18728), .A2(n16840), .ZN(n16828) );
  AOI21_X1 U20008 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(n16828), .A(
        P3_REIP_REG_8__SCAN_IN), .ZN(n16818) );
  AOI21_X1 U20009 ( .B1(n17761), .B2(n16824), .A(n16814), .ZN(n17764) );
  NOR2_X1 U20010 ( .A1(n16815), .A2(n16835), .ZN(n16816) );
  XNOR2_X1 U20011 ( .A(n17764), .B(n16816), .ZN(n16817) );
  OAI22_X1 U20012 ( .A1(n16819), .A2(n16818), .B1(n18698), .B2(n16817), .ZN(
        n16820) );
  AOI211_X1 U20013 ( .C1(n16902), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16821), .B(n16820), .ZN(n16822) );
  OAI211_X1 U20014 ( .C1(n16914), .C2(n17184), .A(n16822), .B(n18077), .ZN(
        P3_U2663) );
  AOI22_X1 U20015 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16902), .B1(
        n16875), .B2(P3_EBX_REG_7__SCAN_IN), .ZN(n16832) );
  OAI21_X1 U20016 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16823), .A(n16849), .ZN(
        n16838) );
  OAI21_X1 U20017 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16825), .A(
        n16824), .ZN(n17782) );
  OAI21_X1 U20018 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16833), .A(
        n16872), .ZN(n16836) );
  OAI21_X1 U20019 ( .B1(n17782), .B2(n16836), .A(n16881), .ZN(n16826) );
  AOI21_X1 U20020 ( .B1(n17782), .B2(n16836), .A(n16826), .ZN(n16827) );
  AOI221_X1 U20021 ( .B1(n16828), .B2(n18730), .C1(n16838), .C2(
        P3_REIP_REG_7__SCAN_IN), .A(n16827), .ZN(n16831) );
  OAI211_X1 U20022 ( .C1(n16841), .C2(n17191), .A(n16883), .B(n16829), .ZN(
        n16830) );
  NAND4_X1 U20023 ( .A1(n16832), .A2(n16831), .A3(n18077), .A4(n16830), .ZN(
        P3_U2664) );
  OAI21_X1 U20024 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16847), .A(
        n16833), .ZN(n16834) );
  INV_X1 U20025 ( .A(n16834), .ZN(n17795) );
  OAI21_X1 U20026 ( .B1(n16847), .B2(n16835), .A(n17795), .ZN(n16846) );
  NOR3_X1 U20027 ( .A1(n17795), .A2(n18698), .A3(n16836), .ZN(n16837) );
  AOI211_X1 U20028 ( .C1(n16875), .C2(P3_EBX_REG_6__SCAN_IN), .A(n9654), .B(
        n16837), .ZN(n16845) );
  INV_X1 U20029 ( .A(n16838), .ZN(n16839) );
  AOI21_X1 U20030 ( .B1(n18728), .B2(n16840), .A(n16839), .ZN(n16843) );
  AOI211_X1 U20031 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16852), .A(n16841), .B(
        n16913), .ZN(n16842) );
  AOI211_X1 U20032 ( .C1(n16902), .C2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n16843), .B(n16842), .ZN(n16844) );
  OAI211_X1 U20033 ( .C1(n16910), .C2(n16846), .A(n16845), .B(n16844), .ZN(
        P3_U2665) );
  INV_X1 U20034 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16856) );
  NOR2_X1 U20035 ( .A1(n16904), .A2(n16857), .ZN(n16865) );
  AOI21_X1 U20036 ( .B1(P3_REIP_REG_4__SCAN_IN), .B2(n16865), .A(
        P3_REIP_REG_5__SCAN_IN), .ZN(n16850) );
  NAND2_X1 U20037 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17806), .ZN(
        n16862) );
  AOI21_X1 U20038 ( .B1(n16856), .B2(n16862), .A(n16847), .ZN(n17804) );
  OAI21_X1 U20039 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16862), .A(
        n16872), .ZN(n16863) );
  XOR2_X1 U20040 ( .A(n17804), .B(n16863), .Z(n16848) );
  OAI22_X1 U20041 ( .A1(n16850), .A2(n16849), .B1(n18698), .B2(n16848), .ZN(
        n16851) );
  AOI211_X1 U20042 ( .C1(n16875), .C2(P3_EBX_REG_5__SCAN_IN), .A(n9654), .B(
        n16851), .ZN(n16855) );
  OAI211_X1 U20043 ( .C1(n16858), .C2(n16853), .A(n16883), .B(n16852), .ZN(
        n16854) );
  OAI211_X1 U20044 ( .C1(n16894), .C2(n16856), .A(n16855), .B(n16854), .ZN(
        P3_U2666) );
  INV_X1 U20045 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18724) );
  AOI21_X1 U20046 ( .B1(n16873), .B2(n16857), .A(n16912), .ZN(n16877) );
  AOI211_X1 U20047 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16882), .A(n16858), .B(
        n16913), .ZN(n16861) );
  NAND2_X1 U20048 ( .A1(n18188), .A2(n18854), .ZN(n16919) );
  INV_X1 U20049 ( .A(n16919), .ZN(n18856) );
  OAI21_X1 U20050 ( .B1(n17171), .B2(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n18856), .ZN(n16859) );
  OAI211_X1 U20051 ( .C1(n17824), .C2(n16894), .A(n18077), .B(n16859), .ZN(
        n16860) );
  AOI211_X1 U20052 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16875), .A(n16861), .B(
        n16860), .ZN(n16870) );
  NOR2_X1 U20053 ( .A1(n17851), .A2(n17809), .ZN(n16871) );
  OAI21_X1 U20054 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16871), .A(
        n16862), .ZN(n17820) );
  INV_X1 U20055 ( .A(n17820), .ZN(n16864) );
  NAND2_X1 U20056 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16911), .ZN(
        n16890) );
  OR2_X1 U20057 ( .A1(n17809), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17815) );
  OAI22_X1 U20058 ( .A1(n16864), .A2(n16863), .B1(n16890), .B2(n17815), .ZN(
        n16868) );
  INV_X1 U20059 ( .A(n16865), .ZN(n16866) );
  OAI22_X1 U20060 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16866), .B1(n16901), 
        .B2(n17820), .ZN(n16867) );
  AOI21_X1 U20061 ( .B1(n16881), .B2(n16868), .A(n16867), .ZN(n16869) );
  OAI211_X1 U20062 ( .C1(n18724), .C2(n16877), .A(n16870), .B(n16869), .ZN(
        P3_U2667) );
  INV_X1 U20063 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16886) );
  NAND2_X1 U20064 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16887) );
  AOI21_X1 U20065 ( .B1(n16886), .B2(n16887), .A(n16871), .ZN(n17833) );
  INV_X1 U20066 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17844) );
  OAI21_X1 U20067 ( .B1(n17844), .B2(n16890), .A(n16872), .ZN(n16889) );
  XNOR2_X1 U20068 ( .A(n17833), .B(n16889), .ZN(n16880) );
  NAND3_X1 U20069 ( .A1(n16873), .A2(P3_REIP_REG_1__SCAN_IN), .A3(
        P3_REIP_REG_2__SCAN_IN), .ZN(n16878) );
  INV_X1 U20070 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n21058) );
  NOR2_X1 U20071 ( .A1(n18820), .A2(n18659), .ZN(n16888) );
  INV_X1 U20072 ( .A(n16888), .ZN(n18643) );
  AOI21_X1 U20073 ( .B1(n18643), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n17159), .ZN(n16874) );
  INV_X1 U20074 ( .A(n16874), .ZN(n18791) );
  AOI22_X1 U20075 ( .A1(n16875), .A2(P3_EBX_REG_3__SCAN_IN), .B1(n18856), .B2(
        n18791), .ZN(n16876) );
  OAI221_X1 U20076 ( .B1(P3_REIP_REG_3__SCAN_IN), .B2(n16878), .C1(n21058), 
        .C2(n16877), .A(n16876), .ZN(n16879) );
  AOI21_X1 U20077 ( .B1(n16881), .B2(n16880), .A(n16879), .ZN(n16885) );
  OAI211_X1 U20078 ( .C1(n16892), .C2(n17200), .A(n16883), .B(n16882), .ZN(
        n16884) );
  OAI211_X1 U20079 ( .C1(n16894), .C2(n16886), .A(n16885), .B(n16884), .ZN(
        P3_U2668) );
  OAI21_X1 U20080 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16887), .ZN(n17841) );
  AOI21_X1 U20081 ( .B1(n18807), .B2(n18665), .A(n16888), .ZN(n18803) );
  AOI22_X1 U20082 ( .A1(n16912), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n18803), 
        .B2(n18856), .ZN(n16900) );
  INV_X1 U20083 ( .A(n17841), .ZN(n16891) );
  AOI211_X1 U20084 ( .C1(n16891), .C2(n16890), .A(n18698), .B(n16889), .ZN(
        n16898) );
  INV_X1 U20085 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18720) );
  INV_X1 U20086 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18721) );
  AOI221_X1 U20087 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_2__SCAN_IN), 
        .C1(n18720), .C2(n18721), .A(n16904), .ZN(n16897) );
  INV_X1 U20088 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17223) );
  INV_X1 U20089 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17217) );
  NAND2_X1 U20090 ( .A1(n17223), .A2(n17217), .ZN(n16893) );
  AOI211_X1 U20091 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16893), .A(n16892), .B(
        n16913), .ZN(n16896) );
  OAI22_X1 U20092 ( .A1(n17844), .A2(n16894), .B1(n16914), .B2(n17212), .ZN(
        n16895) );
  NOR4_X1 U20093 ( .A1(n16898), .A2(n16897), .A3(n16896), .A4(n16895), .ZN(
        n16899) );
  OAI211_X1 U20094 ( .C1(n17841), .C2(n16901), .A(n16900), .B(n16899), .ZN(
        P3_U2669) );
  AOI21_X1 U20095 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16903), .A(
        n16902), .ZN(n16909) );
  OAI22_X1 U20096 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16904), .B1(n16914), 
        .B2(n17217), .ZN(n16907) );
  OAI21_X1 U20097 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17210), .ZN(n17219) );
  NAND2_X1 U20098 ( .A1(n16905), .A2(n18665), .ZN(n18808) );
  OAI22_X1 U20099 ( .A1(n16913), .A2(n17219), .B1(n18808), .B2(n16919), .ZN(
        n16906) );
  AOI211_X1 U20100 ( .C1(n16912), .C2(P3_REIP_REG_1__SCAN_IN), .A(n16907), .B(
        n16906), .ZN(n16908) );
  OAI221_X1 U20101 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16910), .C1(
        n17851), .C2(n16909), .A(n16908), .ZN(P3_U2670) );
  INV_X1 U20102 ( .A(n18794), .ZN(n18852) );
  NOR3_X1 U20103 ( .A1(n18852), .A2(n16912), .A3(n16911), .ZN(n16916) );
  AOI21_X1 U20104 ( .B1(n16914), .B2(n16913), .A(n17223), .ZN(n16915) );
  AOI211_X1 U20105 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(n16917), .A(n16916), .B(
        n16915), .ZN(n16918) );
  OAI21_X1 U20106 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n16919), .A(
        n16918), .ZN(P3_U2671) );
  INV_X1 U20107 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16920) );
  NOR2_X1 U20108 ( .A1(n16920), .A2(n17035), .ZN(n16997) );
  INV_X1 U20109 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16958) );
  NAND4_X1 U20110 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n16921)
         );
  NOR3_X1 U20111 ( .A1(n16958), .A2(n16955), .A3(n16921), .ZN(n16922) );
  NAND4_X1 U20112 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n16997), .A4(n16922), .ZN(n16925) );
  NOR2_X1 U20113 ( .A1(n21042), .A2(n16925), .ZN(n16950) );
  NAND2_X1 U20114 ( .A1(n17214), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16924) );
  NAND2_X1 U20115 ( .A1(n16950), .A2(n18219), .ZN(n16923) );
  OAI22_X1 U20116 ( .A1(n16950), .A2(n16924), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16923), .ZN(P3_U2672) );
  NAND2_X1 U20117 ( .A1(n21042), .A2(n16925), .ZN(n16926) );
  NAND2_X1 U20118 ( .A1(n16926), .A2(n17214), .ZN(n16949) );
  AOI22_X1 U20119 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16930) );
  AOI22_X1 U20120 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16929) );
  AOI22_X1 U20121 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16928) );
  AOI22_X1 U20122 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16927) );
  NAND4_X1 U20123 ( .A1(n16930), .A2(n16929), .A3(n16928), .A4(n16927), .ZN(
        n16936) );
  AOI22_X1 U20124 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16934) );
  AOI22_X1 U20125 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16933) );
  AOI22_X1 U20126 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16932) );
  AOI22_X1 U20127 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16931) );
  NAND4_X1 U20128 ( .A1(n16934), .A2(n16933), .A3(n16932), .A4(n16931), .ZN(
        n16935) );
  NOR2_X1 U20129 ( .A1(n16936), .A2(n16935), .ZN(n16948) );
  AOI22_X1 U20130 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16947) );
  AOI22_X1 U20131 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16946) );
  AOI22_X1 U20132 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16937) );
  OAI21_X1 U20133 ( .B1(n16938), .B2(n21092), .A(n16937), .ZN(n16944) );
  AOI22_X1 U20134 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16942) );
  AOI22_X1 U20135 ( .A1(n15559), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16941) );
  AOI22_X1 U20136 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16940) );
  AOI22_X1 U20137 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16939) );
  NAND4_X1 U20138 ( .A1(n16942), .A2(n16941), .A3(n16940), .A4(n16939), .ZN(
        n16943) );
  AOI211_X1 U20139 ( .C1(n17050), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n16944), .B(n16943), .ZN(n16945) );
  NAND3_X1 U20140 ( .A1(n16947), .A2(n16946), .A3(n16945), .ZN(n16952) );
  NAND2_X1 U20141 ( .A1(n16953), .A2(n16952), .ZN(n16951) );
  XNOR2_X1 U20142 ( .A(n16948), .B(n16951), .ZN(n17234) );
  OAI22_X1 U20143 ( .A1(n16950), .A2(n16949), .B1(n17234), .B2(n17214), .ZN(
        P3_U2673) );
  OAI21_X1 U20144 ( .B1(n16953), .B2(n16952), .A(n16951), .ZN(n17238) );
  INV_X1 U20145 ( .A(n16954), .ZN(n16957) );
  OAI21_X1 U20146 ( .B1(n16964), .B2(n16955), .A(n16958), .ZN(n16956) );
  OAI21_X1 U20147 ( .B1(n16958), .B2(n16957), .A(n16956), .ZN(n16959) );
  OAI21_X1 U20148 ( .B1(n17238), .B2(n17214), .A(n16959), .ZN(P3_U2674) );
  OAI21_X1 U20149 ( .B1(n16962), .B2(n16961), .A(n16960), .ZN(n17248) );
  NAND3_X1 U20150 ( .A1(n16964), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17214), 
        .ZN(n16963) );
  OAI221_X1 U20151 ( .B1(n16964), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17214), 
        .C2(n17248), .A(n16963), .ZN(P3_U2676) );
  INV_X1 U20152 ( .A(n16964), .ZN(n16967) );
  AOI21_X1 U20153 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17214), .A(n16973), .ZN(
        n16966) );
  XNOR2_X1 U20154 ( .A(n16965), .B(n16969), .ZN(n17253) );
  OAI22_X1 U20155 ( .A1(n16967), .A2(n16966), .B1(n17214), .B2(n17253), .ZN(
        P3_U2677) );
  INV_X1 U20156 ( .A(n16968), .ZN(n16976) );
  AOI21_X1 U20157 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17214), .A(n16976), .ZN(
        n16972) );
  OAI21_X1 U20158 ( .B1(n16971), .B2(n16970), .A(n16969), .ZN(n17258) );
  OAI22_X1 U20159 ( .A1(n16973), .A2(n16972), .B1(n17214), .B2(n17258), .ZN(
        P3_U2678) );
  AOI21_X1 U20160 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17214), .A(n16982), .ZN(
        n16975) );
  XNOR2_X1 U20161 ( .A(n16974), .B(n16978), .ZN(n17263) );
  OAI22_X1 U20162 ( .A1(n16976), .A2(n16975), .B1(n17214), .B2(n17263), .ZN(
        P3_U2679) );
  INV_X1 U20163 ( .A(n16977), .ZN(n16996) );
  AOI21_X1 U20164 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17214), .A(n16996), .ZN(
        n16981) );
  OAI21_X1 U20165 ( .B1(n16980), .B2(n16979), .A(n16978), .ZN(n17268) );
  OAI22_X1 U20166 ( .A1(n16982), .A2(n16981), .B1(n17214), .B2(n17268), .ZN(
        P3_U2680) );
  AOI21_X1 U20167 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17214), .A(n16983), .ZN(
        n16995) );
  AOI22_X1 U20168 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16993) );
  AOI22_X1 U20169 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16992) );
  AOI22_X1 U20170 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16984) );
  OAI21_X1 U20171 ( .B1(n10156), .B2(n21092), .A(n16984), .ZN(n16990) );
  AOI22_X1 U20172 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11485), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16988) );
  AOI22_X1 U20173 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16987) );
  AOI22_X1 U20174 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16986) );
  AOI22_X1 U20175 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n9652), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16985) );
  NAND4_X1 U20176 ( .A1(n16988), .A2(n16987), .A3(n16986), .A4(n16985), .ZN(
        n16989) );
  AOI211_X1 U20177 ( .C1(n17055), .C2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n16990), .B(n16989), .ZN(n16991) );
  NAND3_X1 U20178 ( .A1(n16993), .A2(n16992), .A3(n16991), .ZN(n17269) );
  INV_X1 U20179 ( .A(n17269), .ZN(n16994) );
  OAI22_X1 U20180 ( .A1(n16996), .A2(n16995), .B1(n16994), .B2(n17214), .ZN(
        P3_U2681) );
  NOR2_X1 U20181 ( .A1(n17221), .A2(n16997), .ZN(n17021) );
  AOI22_X1 U20182 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15557), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17001) );
  AOI22_X1 U20183 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17000) );
  AOI22_X1 U20184 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16999) );
  AOI22_X1 U20185 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n9652), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16998) );
  NAND4_X1 U20186 ( .A1(n17001), .A2(n17000), .A3(n16999), .A4(n16998), .ZN(
        n17007) );
  AOI22_X1 U20187 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17005) );
  AOI22_X1 U20188 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17004) );
  AOI22_X1 U20189 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20190 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17002) );
  NAND4_X1 U20191 ( .A1(n17005), .A2(n17004), .A3(n17003), .A4(n17002), .ZN(
        n17006) );
  OR2_X1 U20192 ( .A1(n17007), .A2(n17006), .ZN(n17276) );
  AOI22_X1 U20193 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17021), .B1(n17221), 
        .B2(n17276), .ZN(n17008) );
  OAI21_X1 U20194 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17009), .A(n17008), .ZN(
        P3_U2682) );
  AOI22_X1 U20195 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17020) );
  AOI22_X1 U20196 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17019) );
  AOI22_X1 U20197 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17010) );
  OAI21_X1 U20198 ( .B1(n10155), .B2(n21097), .A(n17010), .ZN(n17016) );
  AOI22_X1 U20199 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17014) );
  AOI22_X1 U20200 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17013) );
  AOI22_X1 U20201 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17012) );
  AOI22_X1 U20202 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17011) );
  NAND4_X1 U20203 ( .A1(n17014), .A2(n17013), .A3(n17012), .A4(n17011), .ZN(
        n17015) );
  AOI211_X1 U20204 ( .C1(n17017), .C2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n17016), .B(n17015), .ZN(n17018) );
  NAND3_X1 U20205 ( .A1(n17020), .A2(n17019), .A3(n17018), .ZN(n17280) );
  INV_X1 U20206 ( .A(n17280), .ZN(n17024) );
  OAI21_X1 U20207 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17022), .A(n17021), .ZN(
        n17023) );
  OAI21_X1 U20208 ( .B1(n17024), .B2(n17214), .A(n17023), .ZN(P3_U2683) );
  AOI22_X1 U20209 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20210 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11485), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17027) );
  AOI22_X1 U20211 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17026) );
  AOI22_X1 U20212 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17025) );
  NAND4_X1 U20213 ( .A1(n17028), .A2(n17027), .A3(n17026), .A4(n17025), .ZN(
        n17034) );
  AOI22_X1 U20214 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17032) );
  AOI22_X1 U20215 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9667), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17031) );
  AOI22_X1 U20216 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17030) );
  AOI22_X1 U20217 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17029) );
  NAND4_X1 U20218 ( .A1(n17032), .A2(n17031), .A3(n17030), .A4(n17029), .ZN(
        n17033) );
  NOR2_X1 U20219 ( .A1(n17034), .A2(n17033), .ZN(n17289) );
  OAI21_X1 U20220 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17049), .A(n17035), .ZN(
        n17036) );
  AOI22_X1 U20221 ( .A1(n17221), .A2(n17289), .B1(n17036), .B2(n17214), .ZN(
        P3_U2684) );
  OAI21_X1 U20222 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17037), .A(n17214), .ZN(
        n17048) );
  AOI22_X1 U20223 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20224 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17040) );
  AOI22_X1 U20225 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20226 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17038) );
  NAND4_X1 U20227 ( .A1(n17041), .A2(n17040), .A3(n17039), .A4(n17038), .ZN(
        n17047) );
  AOI22_X1 U20228 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11485), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17045) );
  AOI22_X1 U20229 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U20230 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U20231 ( .A1(n17151), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17042) );
  NAND4_X1 U20232 ( .A1(n17045), .A2(n17044), .A3(n17043), .A4(n17042), .ZN(
        n17046) );
  NOR2_X1 U20233 ( .A1(n17047), .A2(n17046), .ZN(n17294) );
  OAI22_X1 U20234 ( .A1(n17049), .A2(n17048), .B1(n17294), .B2(n17214), .ZN(
        P3_U2685) );
  AOI22_X1 U20235 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n9653), .ZN(n17054) );
  AOI22_X1 U20236 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17160), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17151), .ZN(n17053) );
  AOI22_X1 U20237 ( .A1(n17050), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17052) );
  AOI22_X1 U20238 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n9655), .ZN(n17051) );
  NAND4_X1 U20239 ( .A1(n17054), .A2(n17053), .A3(n17052), .A4(n17051), .ZN(
        n17061) );
  AOI22_X1 U20240 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17149), .ZN(n17059) );
  AOI22_X1 U20241 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17058) );
  AOI22_X1 U20242 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17055), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17057) );
  AOI22_X1 U20243 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17159), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17056) );
  NAND4_X1 U20244 ( .A1(n17059), .A2(n17058), .A3(n17057), .A4(n17056), .ZN(
        n17060) );
  NOR2_X1 U20245 ( .A1(n17061), .A2(n17060), .ZN(n17299) );
  NOR2_X1 U20246 ( .A1(n17221), .A2(n17063), .ZN(n17076) );
  OAI21_X1 U20247 ( .B1(n17299), .B2(n17214), .A(n17064), .ZN(P3_U2686) );
  AOI22_X1 U20248 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U20249 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17067) );
  AOI22_X1 U20250 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11485), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17066) );
  AOI22_X1 U20251 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17065) );
  NAND4_X1 U20252 ( .A1(n17068), .A2(n17067), .A3(n17066), .A4(n17065), .ZN(
        n17075) );
  AOI22_X1 U20253 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U20254 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17072) );
  AOI22_X1 U20255 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U20256 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17070) );
  NAND4_X1 U20257 ( .A1(n17073), .A2(n17072), .A3(n17071), .A4(n17070), .ZN(
        n17074) );
  NOR2_X1 U20258 ( .A1(n17075), .A2(n17074), .ZN(n17305) );
  INV_X1 U20259 ( .A(n17089), .ZN(n17077) );
  OAI21_X1 U20260 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17077), .A(n17076), .ZN(
        n17078) );
  OAI21_X1 U20261 ( .B1(n17305), .B2(n17214), .A(n17078), .ZN(P3_U2687) );
  AOI22_X1 U20262 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n17082) );
  AOI22_X1 U20263 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17081) );
  AOI22_X1 U20264 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17080) );
  AOI22_X1 U20265 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17079) );
  NAND4_X1 U20266 ( .A1(n17082), .A2(n17081), .A3(n17080), .A4(n17079), .ZN(
        n17088) );
  AOI22_X1 U20267 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17086) );
  AOI22_X1 U20268 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11446), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17085) );
  AOI22_X1 U20269 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20270 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17083) );
  NAND4_X1 U20271 ( .A1(n17086), .A2(n17085), .A3(n17084), .A4(n17083), .ZN(
        n17087) );
  NOR2_X1 U20272 ( .A1(n17088), .A2(n17087), .ZN(n17309) );
  OAI21_X1 U20273 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17090), .A(n17089), .ZN(
        n17091) );
  AOI22_X1 U20274 ( .A1(n17221), .A2(n17309), .B1(n17091), .B2(n17214), .ZN(
        P3_U2688) );
  AOI22_X1 U20275 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(n9667), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17101) );
  AOI22_X1 U20276 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U20277 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17092) );
  OAI21_X1 U20278 ( .B1(n10155), .B2(n21092), .A(n17092), .ZN(n17098) );
  AOI22_X1 U20279 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20280 ( .A1(n17149), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17095) );
  AOI22_X1 U20281 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17094) );
  AOI22_X1 U20282 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17093) );
  NAND4_X1 U20283 ( .A1(n17096), .A2(n17095), .A3(n17094), .A4(n17093), .ZN(
        n17097) );
  AOI211_X1 U20284 ( .C1(n11524), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n17098), .B(n17097), .ZN(n17099) );
  NAND3_X1 U20285 ( .A1(n17101), .A2(n17100), .A3(n17099), .ZN(n17313) );
  NOR2_X1 U20286 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17102), .ZN(n17103) );
  AOI22_X1 U20287 ( .A1(n17221), .A2(n17313), .B1(n17220), .B2(n17103), .ZN(
        n17104) );
  OAI221_X1 U20288 ( .B1(n17106), .B2(n17118), .C1(n17106), .C2(n17105), .A(
        n17104), .ZN(P3_U2689) );
  AOI22_X1 U20289 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U20290 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17109) );
  AOI22_X1 U20291 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17108) );
  AOI22_X1 U20292 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17107) );
  NAND4_X1 U20293 ( .A1(n17110), .A2(n17109), .A3(n17108), .A4(n17107), .ZN(
        n17116) );
  AOI22_X1 U20294 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17114) );
  AOI22_X1 U20295 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17113) );
  AOI22_X1 U20296 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17176), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17112) );
  AOI22_X1 U20297 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17111) );
  NAND4_X1 U20298 ( .A1(n17114), .A2(n17113), .A3(n17112), .A4(n17111), .ZN(
        n17115) );
  NOR2_X1 U20299 ( .A1(n17116), .A2(n17115), .ZN(n17322) );
  AND2_X1 U20300 ( .A1(n17117), .A2(n17131), .ZN(n17119) );
  OAI22_X1 U20301 ( .A1(n17322), .A2(n17214), .B1(n17119), .B2(n17118), .ZN(
        P3_U2691) );
  AOI22_X1 U20302 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17123) );
  AOI22_X1 U20303 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17122) );
  AOI22_X1 U20304 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17121) );
  AOI22_X1 U20305 ( .A1(n17171), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17120) );
  NAND4_X1 U20306 ( .A1(n17123), .A2(n17122), .A3(n17121), .A4(n17120), .ZN(
        n17130) );
  AOI22_X1 U20307 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17128) );
  AOI22_X1 U20308 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20309 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n15558), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U20310 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17125) );
  NAND4_X1 U20311 ( .A1(n17128), .A2(n17127), .A3(n17126), .A4(n17125), .ZN(
        n17129) );
  NOR2_X1 U20312 ( .A1(n17130), .A2(n17129), .ZN(n17326) );
  OAI21_X1 U20313 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17132), .A(n17131), .ZN(
        n17133) );
  AOI22_X1 U20314 ( .A1(n17221), .A2(n17326), .B1(n17133), .B2(n17214), .ZN(
        P3_U2692) );
  AOI22_X1 U20315 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9651), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17137) );
  AOI22_X1 U20316 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17149), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17136) );
  AOI22_X1 U20317 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17135) );
  AOI22_X1 U20318 ( .A1(n15559), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17134) );
  NAND4_X1 U20319 ( .A1(n17137), .A2(n17136), .A3(n17135), .A4(n17134), .ZN(
        n17144) );
  AOI22_X1 U20320 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17142) );
  AOI22_X1 U20321 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U20322 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U20323 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17151), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17139) );
  NAND4_X1 U20324 ( .A1(n17142), .A2(n17141), .A3(n17140), .A4(n17139), .ZN(
        n17143) );
  NOR2_X1 U20325 ( .A1(n17144), .A2(n17143), .ZN(n17332) );
  OAI33_X1 U20326 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17311), .A3(n17168), 
        .B1(n17146), .B2(n17221), .B3(n17145), .ZN(n17147) );
  INV_X1 U20327 ( .A(n17147), .ZN(n17148) );
  OAI21_X1 U20328 ( .B1(n17332), .B2(n17214), .A(n17148), .ZN(P3_U2693) );
  AOI22_X1 U20329 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17149), .ZN(n17158) );
  AOI22_X1 U20330 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17151), .ZN(n17157) );
  AOI22_X1 U20331 ( .A1(n17153), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17176), .ZN(n17156) );
  AOI22_X1 U20332 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17154), .B1(
        n9655), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17155) );
  NAND4_X1 U20333 ( .A1(n17158), .A2(n17157), .A3(n17156), .A4(n17155), .ZN(
        n17167) );
  AOI22_X1 U20334 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17171), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17165) );
  AOI22_X1 U20335 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17164) );
  AOI22_X1 U20336 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17124), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17163) );
  AOI22_X1 U20337 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n9653), .ZN(n17162) );
  NAND4_X1 U20338 ( .A1(n17165), .A2(n17164), .A3(n17163), .A4(n17162), .ZN(
        n17166) );
  NOR2_X1 U20339 ( .A1(n17167), .A2(n17166), .ZN(n17333) );
  AOI21_X1 U20340 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17183), .A(
        P3_EBX_REG_9__SCAN_IN), .ZN(n17170) );
  NAND2_X1 U20341 ( .A1(n17214), .A2(n17168), .ZN(n17169) );
  OAI22_X1 U20342 ( .A1(n17333), .A2(n17214), .B1(n17170), .B2(n17169), .ZN(
        P3_U2694) );
  AOI22_X1 U20343 ( .A1(n17017), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9652), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17175) );
  AOI22_X1 U20344 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17174) );
  AOI22_X1 U20345 ( .A1(n17138), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17171), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17173) );
  AOI22_X1 U20346 ( .A1(n9655), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11446), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17172) );
  NAND4_X1 U20347 ( .A1(n17175), .A2(n17174), .A3(n17173), .A4(n17172), .ZN(
        n17182) );
  AOI22_X1 U20348 ( .A1(n9667), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17055), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17180) );
  AOI22_X1 U20349 ( .A1(n9651), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17050), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U20350 ( .A1(n15559), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11485), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17178) );
  AOI22_X1 U20351 ( .A1(n17176), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9653), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17177) );
  NAND4_X1 U20352 ( .A1(n17180), .A2(n17179), .A3(n17178), .A4(n17177), .ZN(
        n17181) );
  NOR2_X1 U20353 ( .A1(n17182), .A2(n17181), .ZN(n17339) );
  OAI33_X1 U20354 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17311), .A3(n17185), .B1(
        n17184), .B2(n17221), .B3(n17183), .ZN(n17186) );
  INV_X1 U20355 ( .A(n17186), .ZN(n17187) );
  OAI21_X1 U20356 ( .B1(n17339), .B2(n17214), .A(n17187), .ZN(P3_U2695) );
  NAND2_X1 U20357 ( .A1(n17214), .A2(n17188), .ZN(n17193) );
  NOR3_X1 U20358 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17311), .A3(n17188), .ZN(
        n17189) );
  AOI21_X1 U20359 ( .B1(n17221), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n17189), .ZN(n17190) );
  OAI21_X1 U20360 ( .B1(n17191), .B2(n17193), .A(n17190), .ZN(P3_U2696) );
  NOR2_X1 U20361 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n17198), .ZN(n17194) );
  INV_X1 U20362 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17192) );
  OAI22_X1 U20363 ( .A1(n17194), .A2(n17193), .B1(n17192), .B2(n17214), .ZN(
        P3_U2697) );
  NOR2_X1 U20364 ( .A1(n17211), .A2(n17201), .ZN(n17195) );
  OAI21_X1 U20365 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17195), .A(n17214), .ZN(
        n17197) );
  INV_X1 U20366 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17196) );
  OAI22_X1 U20367 ( .A1(n17198), .A2(n17197), .B1(n17196), .B2(n17214), .ZN(
        P3_U2698) );
  NAND2_X1 U20368 ( .A1(n17199), .A2(n17220), .ZN(n17205) );
  NOR2_X1 U20369 ( .A1(n17200), .A2(n17205), .ZN(n17208) );
  AOI21_X1 U20370 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17214), .A(n17208), .ZN(
        n17204) );
  NOR2_X1 U20371 ( .A1(n17201), .A2(n17218), .ZN(n17203) );
  INV_X1 U20372 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17202) );
  OAI22_X1 U20373 ( .A1(n17204), .A2(n17203), .B1(n17202), .B2(n17214), .ZN(
        P3_U2699) );
  INV_X1 U20374 ( .A(n17205), .ZN(n17209) );
  AOI21_X1 U20375 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17214), .A(n17209), .ZN(
        n17207) );
  INV_X1 U20376 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17206) );
  OAI22_X1 U20377 ( .A1(n17208), .A2(n17207), .B1(n17206), .B2(n17214), .ZN(
        P3_U2700) );
  AOI221_X1 U20378 ( .B1(n17212), .B2(n17211), .C1(n17212), .C2(n17210), .A(
        n17209), .ZN(n17213) );
  OAI22_X1 U20379 ( .A1(n17214), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17213), .B2(n17221), .ZN(n17215) );
  INV_X1 U20380 ( .A(n17215), .ZN(P3_U2701) );
  OAI222_X1 U20381 ( .A1(n17219), .A2(n17218), .B1(n17217), .B2(n17224), .C1(
        n17216), .C2(n17214), .ZN(P3_U2702) );
  AOI22_X1 U20382 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17221), .B1(
        n17220), .B2(n17223), .ZN(n17222) );
  OAI21_X1 U20383 ( .B1(n17224), .B2(n17223), .A(n17222), .ZN(P3_U2703) );
  INV_X1 U20384 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17384) );
  INV_X1 U20385 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17388) );
  INV_X1 U20386 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17449) );
  INV_X1 U20387 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17489) );
  NAND2_X1 U20388 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n17371) );
  NAND2_X1 U20389 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .ZN(n17340) );
  NAND4_X1 U20390 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17225) );
  INV_X1 U20391 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17421) );
  INV_X1 U20392 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17482) );
  NAND4_X1 U20393 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(P3_EAX_REG_9__SCAN_IN), 
        .A3(P3_EAX_REG_12__SCAN_IN), .A4(P3_EAX_REG_11__SCAN_IN), .ZN(n17226)
         );
  NOR3_X1 U20394 ( .A1(n17421), .A2(n17482), .A3(n17226), .ZN(n17312) );
  NAND3_X1 U20395 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17310), .A3(n17312), 
        .ZN(n17314) );
  INV_X1 U20396 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17403) );
  INV_X1 U20397 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17443) );
  NOR2_X1 U20398 ( .A1(n17403), .A2(n17443), .ZN(n17270) );
  NAND4_X1 U20399 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17270), .A3(
        P3_EAX_REG_20__SCAN_IN), .A4(P3_EAX_REG_19__SCAN_IN), .ZN(n17275) );
  NAND2_X1 U20400 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17265), .ZN(n17264) );
  NAND2_X1 U20401 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17260), .ZN(n17259) );
  NAND2_X1 U20402 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17249), .ZN(n17245) );
  NAND2_X1 U20403 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17241), .ZN(n17235) );
  NAND2_X1 U20404 ( .A1(n17231), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17230) );
  NOR2_X2 U20405 ( .A1(n18212), .A2(n17363), .ZN(n17300) );
  OAI22_X1 U20406 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17361), .B1(n17347), 
        .B2(n17231), .ZN(n17227) );
  AOI22_X1 U20407 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17300), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17227), .ZN(n17228) );
  OAI21_X1 U20408 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17230), .A(n17228), .ZN(
        P3_U2704) );
  NOR2_X2 U20409 ( .A1(n17229), .A2(n17363), .ZN(n17301) );
  AOI22_X1 U20410 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17301), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17300), .ZN(n17233) );
  OAI211_X1 U20411 ( .C1(n17231), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17363), .B(
        n17230), .ZN(n17232) );
  OAI211_X1 U20412 ( .C1(n17234), .C2(n17375), .A(n17233), .B(n17232), .ZN(
        P3_U2705) );
  AOI22_X1 U20413 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17301), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17300), .ZN(n17237) );
  OAI211_X1 U20414 ( .C1(n17241), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17363), .B(
        n17235), .ZN(n17236) );
  OAI211_X1 U20415 ( .C1(n17238), .C2(n17375), .A(n17237), .B(n17236), .ZN(
        P3_U2706) );
  AOI22_X1 U20416 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17301), .B1(n17345), .B2(
        n17239), .ZN(n17240) );
  INV_X1 U20417 ( .A(n17240), .ZN(n17243) );
  AOI211_X1 U20418 ( .C1(n17384), .C2(n17245), .A(n17241), .B(n17347), .ZN(
        n17242) );
  AOI211_X1 U20419 ( .C1(n17300), .C2(BUF2_REG_28__SCAN_IN), .A(n17243), .B(
        n17242), .ZN(n17244) );
  INV_X1 U20420 ( .A(n17244), .ZN(P3_U2707) );
  AOI22_X1 U20421 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17301), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17300), .ZN(n17247) );
  OAI211_X1 U20422 ( .C1(n17249), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17363), .B(
        n17245), .ZN(n17246) );
  OAI211_X1 U20423 ( .C1(n17248), .C2(n17375), .A(n17247), .B(n17246), .ZN(
        P3_U2708) );
  AOI22_X1 U20424 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17301), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17300), .ZN(n17252) );
  AOI211_X1 U20425 ( .C1(n17388), .C2(n17254), .A(n17249), .B(n17347), .ZN(
        n17250) );
  INV_X1 U20426 ( .A(n17250), .ZN(n17251) );
  OAI211_X1 U20427 ( .C1(n17253), .C2(n17375), .A(n17252), .B(n17251), .ZN(
        P3_U2709) );
  AOI22_X1 U20428 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17301), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17300), .ZN(n17257) );
  OAI211_X1 U20429 ( .C1(n17255), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17363), .B(
        n17254), .ZN(n17256) );
  OAI211_X1 U20430 ( .C1(n17258), .C2(n17375), .A(n17257), .B(n17256), .ZN(
        P3_U2710) );
  AOI22_X1 U20431 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17301), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17300), .ZN(n17262) );
  OAI211_X1 U20432 ( .C1(n17260), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17363), .B(
        n17259), .ZN(n17261) );
  OAI211_X1 U20433 ( .C1(n17263), .C2(n17375), .A(n17262), .B(n17261), .ZN(
        P3_U2711) );
  AOI22_X1 U20434 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17301), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17300), .ZN(n17267) );
  OAI211_X1 U20435 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17265), .A(n17363), .B(
        n17264), .ZN(n17266) );
  OAI211_X1 U20436 ( .C1(n17268), .C2(n17375), .A(n17267), .B(n17266), .ZN(
        P3_U2712) );
  NAND2_X1 U20437 ( .A1(n17296), .A2(n17449), .ZN(n17274) );
  AOI22_X1 U20438 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17300), .B1(n17345), .B2(
        n17269), .ZN(n17273) );
  NAND3_X1 U20439 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(n17290), .ZN(n17281) );
  NAND2_X1 U20440 ( .A1(n17363), .A2(n17281), .ZN(n17285) );
  OAI21_X1 U20441 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17361), .A(n17285), .ZN(
        n17271) );
  AOI22_X1 U20442 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17301), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17271), .ZN(n17272) );
  OAI211_X1 U20443 ( .C1(n17275), .C2(n17274), .A(n17273), .B(n17272), .ZN(
        P3_U2713) );
  INV_X1 U20444 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17397) );
  AOI22_X1 U20445 ( .A1(n17276), .A2(n17345), .B1(BUF2_REG_21__SCAN_IN), .B2(
        n17300), .ZN(n17277) );
  INV_X1 U20446 ( .A(n17277), .ZN(n17278) );
  AOI21_X1 U20447 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17301), .A(n17278), .ZN(
        n17279) );
  OAI221_X1 U20448 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17281), .C1(n17397), 
        .C2(n17285), .A(n17279), .ZN(P3_U2714) );
  INV_X1 U20449 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17399) );
  AOI22_X1 U20450 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17300), .B1(n17345), .B2(
        n17280), .ZN(n17284) );
  NAND2_X1 U20451 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17290), .ZN(n17286) );
  INV_X1 U20452 ( .A(n17286), .ZN(n17282) );
  AOI22_X1 U20453 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17301), .B1(n17282), .B2(
        n17281), .ZN(n17283) );
  OAI211_X1 U20454 ( .C1(n17399), .C2(n17285), .A(n17284), .B(n17283), .ZN(
        P3_U2715) );
  AOI22_X1 U20455 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17301), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17300), .ZN(n17288) );
  OAI211_X1 U20456 ( .C1(n17290), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17363), .B(
        n17286), .ZN(n17287) );
  OAI211_X1 U20457 ( .C1(n17289), .C2(n17375), .A(n17288), .B(n17287), .ZN(
        P3_U2716) );
  AOI22_X1 U20458 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17301), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17300), .ZN(n17293) );
  NAND2_X1 U20459 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17296), .ZN(n17295) );
  AOI211_X1 U20460 ( .C1(n17403), .C2(n17295), .A(n17290), .B(n17347), .ZN(
        n17291) );
  INV_X1 U20461 ( .A(n17291), .ZN(n17292) );
  OAI211_X1 U20462 ( .C1(n17294), .C2(n17375), .A(n17293), .B(n17292), .ZN(
        P3_U2717) );
  AOI22_X1 U20463 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17301), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17300), .ZN(n17298) );
  OAI211_X1 U20464 ( .C1(n17296), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17363), .B(
        n17295), .ZN(n17297) );
  OAI211_X1 U20465 ( .C1(n17299), .C2(n17375), .A(n17298), .B(n17297), .ZN(
        P3_U2718) );
  AOI22_X1 U20466 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17301), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17300), .ZN(n17304) );
  OAI211_X1 U20467 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17306), .A(n17363), .B(
        n17302), .ZN(n17303) );
  OAI211_X1 U20468 ( .C1(n17305), .C2(n17375), .A(n17304), .B(n17303), .ZN(
        P3_U2719) );
  AOI211_X1 U20469 ( .C1(n17489), .C2(n17314), .A(n17347), .B(n17306), .ZN(
        n17307) );
  AOI21_X1 U20470 ( .B1(n17370), .B2(BUF2_REG_15__SCAN_IN), .A(n17307), .ZN(
        n17308) );
  OAI21_X1 U20471 ( .B1(n17309), .B2(n17375), .A(n17308), .ZN(P3_U2720) );
  INV_X1 U20472 ( .A(n17310), .ZN(n17336) );
  NAND2_X1 U20473 ( .A1(n17312), .A2(n17343), .ZN(n17317) );
  AOI22_X1 U20474 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17370), .B1(n17345), .B2(
        n17313), .ZN(n17316) );
  NAND3_X1 U20475 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17363), .A3(n17314), 
        .ZN(n17315) );
  OAI211_X1 U20476 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17317), .A(n17316), .B(
        n17315), .ZN(P3_U2721) );
  INV_X1 U20477 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17415) );
  NAND2_X1 U20478 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17335), .ZN(n17329) );
  NOR2_X1 U20479 ( .A1(n17415), .A2(n17329), .ZN(n17328) );
  NAND2_X1 U20480 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17328), .ZN(n17321) );
  NAND2_X1 U20481 ( .A1(n17321), .A2(P3_EAX_REG_13__SCAN_IN), .ZN(n17320) );
  AOI22_X1 U20482 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17370), .B1(n17345), .B2(
        n17318), .ZN(n17319) );
  OAI221_X1 U20483 ( .B1(n17321), .B2(P3_EAX_REG_13__SCAN_IN), .C1(n17320), 
        .C2(n17347), .A(n17319), .ZN(P3_U2722) );
  INV_X1 U20484 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17480) );
  INV_X1 U20485 ( .A(n17321), .ZN(n17324) );
  AOI21_X1 U20486 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17363), .A(n17328), .ZN(
        n17323) );
  OAI222_X1 U20487 ( .A1(n17368), .A2(n17480), .B1(n17324), .B2(n17323), .C1(
        n17375), .C2(n17322), .ZN(P3_U2723) );
  OAI21_X1 U20488 ( .B1(n17415), .B2(n17347), .A(n17329), .ZN(n17325) );
  INV_X1 U20489 ( .A(n17325), .ZN(n17327) );
  OAI222_X1 U20490 ( .A1(n17368), .A2(n21082), .B1(n17328), .B2(n17327), .C1(
        n17375), .C2(n17326), .ZN(P3_U2724) );
  OAI211_X1 U20491 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17335), .A(n17363), .B(
        n17329), .ZN(n17331) );
  NAND2_X1 U20492 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17370), .ZN(n17330) );
  OAI211_X1 U20493 ( .C1(n17332), .C2(n17375), .A(n17331), .B(n17330), .ZN(
        P3_U2725) );
  AOI22_X1 U20494 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17343), .B1(
        P3_EAX_REG_9__SCAN_IN), .B2(n17363), .ZN(n17334) );
  OAI222_X1 U20495 ( .A1(n17368), .A2(n17473), .B1(n17335), .B2(n17334), .C1(
        n17375), .C2(n17333), .ZN(P3_U2726) );
  AOI22_X1 U20496 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17370), .B1(n17343), .B2(
        n17421), .ZN(n17338) );
  NAND3_X1 U20497 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17363), .A3(n17336), .ZN(
        n17337) );
  OAI211_X1 U20498 ( .C1(n17339), .C2(n17375), .A(n17338), .B(n17337), .ZN(
        P3_U2727) );
  INV_X1 U20499 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17431) );
  NAND2_X1 U20500 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17367), .ZN(n17353) );
  NOR2_X1 U20501 ( .A1(n17340), .A2(n17353), .ZN(n17352) );
  AOI22_X1 U20502 ( .A1(n17352), .A2(P3_EAX_REG_6__SCAN_IN), .B1(
        P3_EAX_REG_7__SCAN_IN), .B2(n17363), .ZN(n17342) );
  OAI222_X1 U20503 ( .A1(n17368), .A2(n18216), .B1(n17343), .B2(n17342), .C1(
        n17375), .C2(n17341), .ZN(P3_U2728) );
  INV_X1 U20504 ( .A(n17352), .ZN(n17349) );
  NAND2_X1 U20505 ( .A1(n17349), .A2(P3_EAX_REG_6__SCAN_IN), .ZN(n17348) );
  AOI22_X1 U20506 ( .A1(n17370), .A2(BUF2_REG_6__SCAN_IN), .B1(n17345), .B2(
        n17344), .ZN(n17346) );
  OAI221_X1 U20507 ( .B1(n17349), .B2(P3_EAX_REG_6__SCAN_IN), .C1(n17348), 
        .C2(n17347), .A(n17346), .ZN(P3_U2729) );
  INV_X1 U20508 ( .A(n17353), .ZN(n17360) );
  AOI22_X1 U20509 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17363), .B1(
        P3_EAX_REG_4__SCAN_IN), .B2(n17360), .ZN(n17351) );
  OAI222_X1 U20510 ( .A1(n18207), .A2(n17368), .B1(n17352), .B2(n17351), .C1(
        n17375), .C2(n17350), .ZN(P3_U2730) );
  INV_X1 U20511 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18203) );
  INV_X1 U20512 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17427) );
  NOR2_X1 U20513 ( .A1(n17427), .A2(n17353), .ZN(n17357) );
  AOI21_X1 U20514 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17363), .A(n17360), .ZN(
        n17356) );
  INV_X1 U20515 ( .A(n17354), .ZN(n17355) );
  OAI222_X1 U20516 ( .A1(n18203), .A2(n17368), .B1(n17357), .B2(n17356), .C1(
        n17375), .C2(n17355), .ZN(P3_U2731) );
  AOI21_X1 U20517 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17363), .A(n17367), .ZN(
        n17359) );
  OAI222_X1 U20518 ( .A1(n18199), .A2(n17368), .B1(n17360), .B2(n17359), .C1(
        n17375), .C2(n17358), .ZN(P3_U2732) );
  INV_X1 U20519 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18195) );
  NOR2_X1 U20520 ( .A1(n17371), .A2(n17361), .ZN(n17362) );
  AOI21_X1 U20521 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17363), .A(n17362), .ZN(
        n17366) );
  INV_X1 U20522 ( .A(n17364), .ZN(n17365) );
  OAI222_X1 U20523 ( .A1(n18195), .A2(n17368), .B1(n17367), .B2(n17366), .C1(
        n17375), .C2(n17365), .ZN(P3_U2733) );
  AOI22_X1 U20524 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17370), .B1(n17369), .B2(
        P3_EAX_REG_1__SCAN_IN), .ZN(n17374) );
  OAI211_X1 U20525 ( .C1(P3_EAX_REG_1__SCAN_IN), .C2(P3_EAX_REG_0__SCAN_IN), 
        .A(n17372), .B(n17371), .ZN(n17373) );
  OAI211_X1 U20526 ( .C1(n17376), .C2(n17375), .A(n17374), .B(n17373), .ZN(
        P3_U2734) );
  NOR2_X1 U20527 ( .A1(n18800), .A2(n18702), .ZN(n18835) );
  NOR2_X1 U20528 ( .A1(n17404), .A2(n17379), .ZN(P3_U2736) );
  INV_X1 U20529 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17459) );
  NOR2_X1 U20530 ( .A1(n17436), .A2(n18188), .ZN(n17393) );
  INV_X2 U20531 ( .A(n17404), .ZN(n17433) );
  AOI22_X1 U20532 ( .A1(n18835), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17381) );
  OAI21_X1 U20533 ( .B1(n17459), .B2(n17407), .A(n17381), .ZN(P3_U2737) );
  INV_X1 U20534 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17457) );
  AOI22_X1 U20535 ( .A1(n18835), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17382) );
  OAI21_X1 U20536 ( .B1(n17457), .B2(n17407), .A(n17382), .ZN(P3_U2738) );
  AOI22_X1 U20537 ( .A1(n18835), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17383) );
  OAI21_X1 U20538 ( .B1(n17384), .B2(n17407), .A(n17383), .ZN(P3_U2739) );
  INV_X1 U20539 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17386) );
  AOI22_X1 U20540 ( .A1(n18835), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17385) );
  OAI21_X1 U20541 ( .B1(n17386), .B2(n17407), .A(n17385), .ZN(P3_U2740) );
  AOI22_X1 U20542 ( .A1(n18835), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17387) );
  OAI21_X1 U20543 ( .B1(n17388), .B2(n17407), .A(n17387), .ZN(P3_U2741) );
  INV_X1 U20544 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17390) );
  AOI22_X1 U20545 ( .A1(n18835), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17389) );
  OAI21_X1 U20546 ( .B1(n17390), .B2(n17407), .A(n17389), .ZN(P3_U2742) );
  INV_X1 U20547 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17392) );
  CLKBUF_X1 U20548 ( .A(n18835), .Z(n17434) );
  AOI22_X1 U20549 ( .A1(n17434), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17391) );
  OAI21_X1 U20550 ( .B1(n17392), .B2(n17407), .A(n17391), .ZN(P3_U2743) );
  INV_X1 U20551 ( .A(P3_DATAO_REG_23__SCAN_IN), .ZN(n20936) );
  AOI22_X1 U20552 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17393), .B1(n18835), 
        .B2(P3_UWORD_REG_7__SCAN_IN), .ZN(n17394) );
  OAI21_X1 U20553 ( .B1(n20936), .B2(n17404), .A(n17394), .ZN(P3_U2744) );
  AOI22_X1 U20554 ( .A1(n17434), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17395) );
  OAI21_X1 U20555 ( .B1(n17449), .B2(n17407), .A(n17395), .ZN(P3_U2745) );
  AOI22_X1 U20556 ( .A1(n17434), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17396) );
  OAI21_X1 U20557 ( .B1(n17397), .B2(n17407), .A(n17396), .ZN(P3_U2746) );
  AOI22_X1 U20558 ( .A1(n17434), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17398) );
  OAI21_X1 U20559 ( .B1(n17399), .B2(n17407), .A(n17398), .ZN(P3_U2747) );
  INV_X1 U20560 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17401) );
  AOI22_X1 U20561 ( .A1(n17434), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17400) );
  OAI21_X1 U20562 ( .B1(n17401), .B2(n17407), .A(n17400), .ZN(P3_U2748) );
  AOI22_X1 U20563 ( .A1(n17434), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17402) );
  OAI21_X1 U20564 ( .B1(n17403), .B2(n17407), .A(n17402), .ZN(P3_U2749) );
  AOI22_X1 U20565 ( .A1(n17434), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17405) );
  OAI21_X1 U20566 ( .B1(n17443), .B2(n17407), .A(n17405), .ZN(P3_U2750) );
  INV_X1 U20567 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17408) );
  AOI22_X1 U20568 ( .A1(n17434), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17406) );
  OAI21_X1 U20569 ( .B1(n17408), .B2(n17407), .A(n17406), .ZN(P3_U2751) );
  AOI22_X1 U20570 ( .A1(n17434), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17409) );
  OAI21_X1 U20571 ( .B1(n17489), .B2(n17436), .A(n17409), .ZN(P3_U2752) );
  INV_X1 U20572 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17484) );
  AOI22_X1 U20573 ( .A1(n17434), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17410) );
  OAI21_X1 U20574 ( .B1(n17484), .B2(n17436), .A(n17410), .ZN(P3_U2753) );
  AOI22_X1 U20575 ( .A1(n17434), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17411) );
  OAI21_X1 U20576 ( .B1(n17482), .B2(n17436), .A(n17411), .ZN(P3_U2754) );
  INV_X1 U20577 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17413) );
  AOI22_X1 U20578 ( .A1(n17434), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17412) );
  OAI21_X1 U20579 ( .B1(n17413), .B2(n17436), .A(n17412), .ZN(P3_U2755) );
  AOI22_X1 U20580 ( .A1(n17434), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17414) );
  OAI21_X1 U20581 ( .B1(n17415), .B2(n17436), .A(n17414), .ZN(P3_U2756) );
  INV_X1 U20582 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17417) );
  AOI22_X1 U20583 ( .A1(n17434), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17416) );
  OAI21_X1 U20584 ( .B1(n17417), .B2(n17436), .A(n17416), .ZN(P3_U2757) );
  INV_X1 U20585 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17419) );
  AOI22_X1 U20586 ( .A1(n17434), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17418) );
  OAI21_X1 U20587 ( .B1(n17419), .B2(n17436), .A(n17418), .ZN(P3_U2758) );
  AOI22_X1 U20588 ( .A1(n17434), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17420) );
  OAI21_X1 U20589 ( .B1(n17421), .B2(n17436), .A(n17420), .ZN(P3_U2759) );
  INV_X1 U20590 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17423) );
  AOI22_X1 U20591 ( .A1(n17434), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17422) );
  OAI21_X1 U20592 ( .B1(n17423), .B2(n17436), .A(n17422), .ZN(P3_U2760) );
  INV_X1 U20593 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17468) );
  AOI22_X1 U20594 ( .A1(n17434), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17424) );
  OAI21_X1 U20595 ( .B1(n17468), .B2(n17436), .A(n17424), .ZN(P3_U2761) );
  INV_X1 U20596 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n21094) );
  AOI22_X1 U20597 ( .A1(n17434), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17425) );
  OAI21_X1 U20598 ( .B1(n21094), .B2(n17436), .A(n17425), .ZN(P3_U2762) );
  AOI22_X1 U20599 ( .A1(n17434), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17426) );
  OAI21_X1 U20600 ( .B1(n17427), .B2(n17436), .A(n17426), .ZN(P3_U2763) );
  INV_X1 U20601 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17429) );
  AOI22_X1 U20602 ( .A1(n17434), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17428) );
  OAI21_X1 U20603 ( .B1(n17429), .B2(n17436), .A(n17428), .ZN(P3_U2764) );
  AOI22_X1 U20604 ( .A1(n17434), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17430) );
  OAI21_X1 U20605 ( .B1(n17431), .B2(n17436), .A(n17430), .ZN(P3_U2765) );
  INV_X1 U20606 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17462) );
  AOI22_X1 U20607 ( .A1(n17434), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17432) );
  OAI21_X1 U20608 ( .B1(n17462), .B2(n17436), .A(n17432), .ZN(P3_U2766) );
  AOI22_X1 U20609 ( .A1(n17434), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17433), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17435) );
  OAI21_X1 U20610 ( .B1(n17437), .B2(n17436), .A(n17435), .ZN(P3_U2767) );
  INV_X1 U20611 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18184) );
  NAND2_X1 U20612 ( .A1(n17440), .A2(n17439), .ZN(n17488) );
  AOI22_X1 U20613 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17477), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17476), .ZN(n17441) );
  OAI21_X1 U20614 ( .B1(n18184), .B2(n17479), .A(n17441), .ZN(P3_U2768) );
  AOI22_X1 U20615 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17486), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17476), .ZN(n17442) );
  OAI21_X1 U20616 ( .B1(n17443), .B2(n17488), .A(n17442), .ZN(P3_U2769) );
  AOI22_X1 U20617 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17477), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17476), .ZN(n17444) );
  OAI21_X1 U20618 ( .B1(n18195), .B2(n17479), .A(n17444), .ZN(P3_U2770) );
  AOI22_X1 U20619 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17477), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17476), .ZN(n17445) );
  OAI21_X1 U20620 ( .B1(n18199), .B2(n17479), .A(n17445), .ZN(P3_U2771) );
  AOI22_X1 U20621 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17477), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17476), .ZN(n17446) );
  OAI21_X1 U20622 ( .B1(n18203), .B2(n17479), .A(n17446), .ZN(P3_U2772) );
  AOI22_X1 U20623 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17477), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17476), .ZN(n17447) );
  OAI21_X1 U20624 ( .B1(n18207), .B2(n17479), .A(n17447), .ZN(P3_U2773) );
  AOI22_X1 U20625 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17486), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17476), .ZN(n17448) );
  OAI21_X1 U20626 ( .B1(n17449), .B2(n17488), .A(n17448), .ZN(P3_U2774) );
  AOI22_X1 U20627 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17477), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17476), .ZN(n17450) );
  OAI21_X1 U20628 ( .B1(n18216), .B2(n17479), .A(n17450), .ZN(P3_U2775) );
  AOI22_X1 U20629 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17477), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17476), .ZN(n17451) );
  OAI21_X1 U20630 ( .B1(n17471), .B2(n17479), .A(n17451), .ZN(P3_U2776) );
  AOI22_X1 U20631 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17477), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17476), .ZN(n17452) );
  OAI21_X1 U20632 ( .B1(n17473), .B2(n17479), .A(n17452), .ZN(P3_U2777) );
  INV_X1 U20633 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n20958) );
  AOI22_X1 U20634 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17477), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17476), .ZN(n17453) );
  OAI21_X1 U20635 ( .B1(n20958), .B2(n17479), .A(n17453), .ZN(P3_U2778) );
  AOI22_X1 U20636 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17477), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17476), .ZN(n17454) );
  OAI21_X1 U20637 ( .B1(n21082), .B2(n17479), .A(n17454), .ZN(P3_U2779) );
  AOI22_X1 U20638 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17477), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17476), .ZN(n17455) );
  OAI21_X1 U20639 ( .B1(n17480), .B2(n17479), .A(n17455), .ZN(P3_U2780) );
  AOI22_X1 U20640 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17486), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17476), .ZN(n17456) );
  OAI21_X1 U20641 ( .B1(n17457), .B2(n17488), .A(n17456), .ZN(P3_U2781) );
  AOI22_X1 U20642 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17486), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17476), .ZN(n17458) );
  OAI21_X1 U20643 ( .B1(n17459), .B2(n17488), .A(n17458), .ZN(P3_U2782) );
  AOI22_X1 U20644 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17477), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17476), .ZN(n17460) );
  OAI21_X1 U20645 ( .B1(n18184), .B2(n17479), .A(n17460), .ZN(P3_U2783) );
  AOI22_X1 U20646 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17486), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17476), .ZN(n17461) );
  OAI21_X1 U20647 ( .B1(n17462), .B2(n17488), .A(n17461), .ZN(P3_U2784) );
  AOI22_X1 U20648 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17477), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17476), .ZN(n17463) );
  OAI21_X1 U20649 ( .B1(n18195), .B2(n17479), .A(n17463), .ZN(P3_U2785) );
  AOI22_X1 U20650 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17477), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17476), .ZN(n17464) );
  OAI21_X1 U20651 ( .B1(n18199), .B2(n17479), .A(n17464), .ZN(P3_U2786) );
  AOI22_X1 U20652 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17477), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17485), .ZN(n17465) );
  OAI21_X1 U20653 ( .B1(n18203), .B2(n17479), .A(n17465), .ZN(P3_U2787) );
  AOI22_X1 U20654 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17477), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17485), .ZN(n17466) );
  OAI21_X1 U20655 ( .B1(n18207), .B2(n17479), .A(n17466), .ZN(P3_U2788) );
  AOI22_X1 U20656 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17486), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17485), .ZN(n17467) );
  OAI21_X1 U20657 ( .B1(n17468), .B2(n17488), .A(n17467), .ZN(P3_U2789) );
  AOI22_X1 U20658 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17477), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17485), .ZN(n17469) );
  OAI21_X1 U20659 ( .B1(n18216), .B2(n17479), .A(n17469), .ZN(P3_U2790) );
  AOI22_X1 U20660 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17477), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17485), .ZN(n17470) );
  OAI21_X1 U20661 ( .B1(n17471), .B2(n17479), .A(n17470), .ZN(P3_U2791) );
  AOI22_X1 U20662 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17477), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17485), .ZN(n17472) );
  OAI21_X1 U20663 ( .B1(n17473), .B2(n17479), .A(n17472), .ZN(P3_U2792) );
  AOI22_X1 U20664 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17477), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17485), .ZN(n17474) );
  OAI21_X1 U20665 ( .B1(n20958), .B2(n17479), .A(n17474), .ZN(P3_U2793) );
  AOI22_X1 U20666 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17477), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17476), .ZN(n17475) );
  OAI21_X1 U20667 ( .B1(n21082), .B2(n17479), .A(n17475), .ZN(P3_U2794) );
  AOI22_X1 U20668 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17477), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17476), .ZN(n17478) );
  OAI21_X1 U20669 ( .B1(n17480), .B2(n17479), .A(n17478), .ZN(P3_U2795) );
  AOI22_X1 U20670 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17486), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17485), .ZN(n17481) );
  OAI21_X1 U20671 ( .B1(n17482), .B2(n17488), .A(n17481), .ZN(P3_U2796) );
  AOI22_X1 U20672 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17486), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17485), .ZN(n17483) );
  OAI21_X1 U20673 ( .B1(n17484), .B2(n17488), .A(n17483), .ZN(P3_U2797) );
  AOI22_X1 U20674 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17486), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17485), .ZN(n17487) );
  OAI21_X1 U20675 ( .B1(n17489), .B2(n17488), .A(n17487), .ZN(P3_U2798) );
  INV_X1 U20676 ( .A(n17810), .ZN(n17689) );
  OAI21_X1 U20677 ( .B1(n17493), .B2(n17689), .A(n17858), .ZN(n17490) );
  AOI21_X1 U20678 ( .B1(n17687), .B2(n17491), .A(n17490), .ZN(n17526) );
  OAI21_X1 U20679 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17600), .A(
        n17526), .ZN(n17512) );
  INV_X1 U20680 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17494) );
  NAND2_X1 U20681 ( .A1(n17493), .A2(n17492), .ZN(n17517) );
  AOI221_X1 U20682 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C1(n17495), .C2(n17494), .A(
        n17517), .ZN(n17497) );
  AOI211_X1 U20683 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17512), .A(
        n17497), .B(n17496), .ZN(n17509) );
  NOR2_X1 U20684 ( .A1(n17850), .A2(n17770), .ZN(n17605) );
  INV_X1 U20685 ( .A(n17498), .ZN(n17868) );
  INV_X1 U20686 ( .A(n17499), .ZN(n17867) );
  OAI22_X1 U20687 ( .A1(n17868), .A2(n17862), .B1(n17867), .B2(n17546), .ZN(
        n17529) );
  NOR2_X1 U20688 ( .A1(n9931), .A2(n17529), .ZN(n17501) );
  NOR3_X1 U20689 ( .A1(n17605), .A2(n17501), .A3(n17500), .ZN(n17506) );
  AOI211_X1 U20690 ( .C1(n17504), .C2(n17503), .A(n17502), .B(n17742), .ZN(
        n17505) );
  AOI211_X1 U20691 ( .C1(n17507), .C2(n17641), .A(n17506), .B(n17505), .ZN(
        n17508) );
  OAI211_X1 U20692 ( .C1(n17696), .C2(n17510), .A(n17509), .B(n17508), .ZN(
        P3_U2802) );
  AOI22_X1 U20693 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17512), .B1(
        n17706), .B2(n17511), .ZN(n17521) );
  INV_X1 U20694 ( .A(n17513), .ZN(n17515) );
  OAI22_X1 U20695 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17517), .B1(
        n17876), .B2(n17742), .ZN(n17518) );
  AOI221_X1 U20696 ( .B1(n17519), .B2(n9931), .C1(n17529), .C2(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n17518), .ZN(n17520) );
  OAI211_X1 U20697 ( .C1(n18077), .C2(n18771), .A(n17521), .B(n17520), .ZN(
        P3_U2803) );
  AOI21_X1 U20698 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17523), .A(
        n17522), .ZN(n17882) );
  AOI21_X1 U20699 ( .B1(n17524), .B2(n18215), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17525) );
  INV_X1 U20700 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18768) );
  OAI22_X1 U20701 ( .A1(n17526), .A2(n17525), .B1(n18077), .B2(n18768), .ZN(
        n17527) );
  AOI221_X1 U20702 ( .B1(n17706), .B2(n17528), .C1(n16366), .C2(n17528), .A(
        n17527), .ZN(n17531) );
  NOR3_X1 U20703 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17892), .A3(
        n17884), .ZN(n17878) );
  AOI22_X1 U20704 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17529), .B1(
        n17641), .B2(n17878), .ZN(n17530) );
  OAI211_X1 U20705 ( .C1(n17882), .C2(n17742), .A(n17531), .B(n17530), .ZN(
        P3_U2804) );
  XOR2_X1 U20706 ( .A(n17892), .B(n17532), .Z(n17886) );
  INV_X1 U20707 ( .A(n17533), .ZN(n17534) );
  AND2_X1 U20708 ( .A1(n17535), .A2(n18566), .ZN(n17563) );
  AOI211_X1 U20709 ( .C1(n17687), .C2(n17534), .A(n17845), .B(n17563), .ZN(
        n17560) );
  OAI21_X1 U20710 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17600), .A(
        n17560), .ZN(n17548) );
  NOR2_X1 U20711 ( .A1(n17691), .A2(n17535), .ZN(n17550) );
  OAI211_X1 U20712 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17550), .B(n17536), .ZN(n17537) );
  NAND2_X1 U20713 ( .A1(n9654), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17894) );
  OAI211_X1 U20714 ( .C1(n17696), .C2(n17538), .A(n17537), .B(n17894), .ZN(
        n17544) );
  XOR2_X1 U20715 ( .A(n17539), .B(n17892), .Z(n17887) );
  OAI21_X1 U20716 ( .B1(n17645), .B2(n17541), .A(n17540), .ZN(n17542) );
  XOR2_X1 U20717 ( .A(n17542), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17891) );
  OAI22_X1 U20718 ( .A1(n17862), .A2(n17887), .B1(n17742), .B2(n17891), .ZN(
        n17543) );
  AOI211_X1 U20719 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17548), .A(
        n17544), .B(n17543), .ZN(n17545) );
  OAI21_X1 U20720 ( .B1(n17546), .B2(n17886), .A(n17545), .ZN(P3_U2805) );
  INV_X1 U20721 ( .A(n17547), .ZN(n17557) );
  NOR2_X1 U20722 ( .A1(n18077), .A2(n18764), .ZN(n17909) );
  AOI221_X1 U20723 ( .B1(n17550), .B2(n17549), .C1(n17548), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17909), .ZN(n17556) );
  NOR2_X1 U20724 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17551), .ZN(
        n17910) );
  OAI21_X1 U20725 ( .B1(n17551), .B2(n17920), .A(n17770), .ZN(n17564) );
  OAI21_X1 U20726 ( .B1(n18008), .B2(n17551), .A(n17850), .ZN(n17565) );
  AND2_X1 U20727 ( .A1(n17564), .A2(n17565), .ZN(n17572) );
  AOI21_X1 U20728 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17553), .A(
        n17552), .ZN(n17912) );
  OAI22_X1 U20729 ( .A1(n17572), .A2(n17906), .B1(n17912), .B2(n17742), .ZN(
        n17554) );
  AOI21_X1 U20730 ( .B1(n17641), .B2(n17910), .A(n17554), .ZN(n17555) );
  OAI211_X1 U20731 ( .C1(n17696), .C2(n17557), .A(n17556), .B(n17555), .ZN(
        P3_U2806) );
  NOR2_X1 U20732 ( .A1(n18077), .A2(n18763), .ZN(n17914) );
  OAI22_X1 U20733 ( .A1(n17560), .A2(n17559), .B1(n17842), .B2(n17558), .ZN(
        n17561) );
  AOI211_X1 U20734 ( .C1(n17563), .C2(n17562), .A(n17914), .B(n17561), .ZN(
        n17571) );
  OAI22_X1 U20735 ( .A1(n18008), .A2(n17565), .B1(n17920), .B2(n17564), .ZN(
        n17569) );
  AOI22_X1 U20736 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17645), .B1(
        n17566), .B2(n17576), .ZN(n17567) );
  NAND2_X1 U20737 ( .A1(n17606), .A2(n17567), .ZN(n17568) );
  XOR2_X1 U20738 ( .A(n17568), .B(n17918), .Z(n17915) );
  AOI22_X1 U20739 ( .A1(n17913), .A2(n17569), .B1(n17768), .B2(n17915), .ZN(
        n17570) );
  OAI211_X1 U20740 ( .C1(n17572), .C2(n17918), .A(n17571), .B(n17570), .ZN(
        P3_U2807) );
  OAI21_X1 U20741 ( .B1(n17573), .B2(n18702), .A(n17858), .ZN(n17574) );
  AOI21_X1 U20742 ( .B1(n17810), .B2(n17582), .A(n17574), .ZN(n17602) );
  OAI21_X1 U20743 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17600), .A(
        n17602), .ZN(n17589) );
  AOI22_X1 U20744 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17589), .B1(
        n17706), .B2(n17575), .ZN(n17586) );
  AOI22_X1 U20745 ( .A1(n17850), .A2(n18008), .B1(n17770), .B2(n17920), .ZN(
        n17657) );
  OAI21_X1 U20746 ( .B1(n17932), .B2(n17605), .A(n17657), .ZN(n17597) );
  NAND2_X1 U20747 ( .A1(n17932), .A2(n17641), .ZN(n17580) );
  INV_X1 U20748 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17928) );
  INV_X1 U20749 ( .A(n17576), .ZN(n17578) );
  OAI221_X1 U20750 ( .B1(n17578), .B2(n17932), .C1(n17578), .C2(n17577), .A(
        n17606), .ZN(n17579) );
  XNOR2_X1 U20751 ( .A(n17928), .B(n17579), .ZN(n17935) );
  OAI22_X1 U20752 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17580), .B1(
        n17935), .B2(n17742), .ZN(n17581) );
  AOI21_X1 U20753 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17597), .A(
        n17581), .ZN(n17585) );
  NAND2_X1 U20754 ( .A1(n9654), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17934) );
  NOR2_X1 U20755 ( .A1(n17691), .A2(n17582), .ZN(n17591) );
  OAI211_X1 U20756 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17591), .B(n17583), .ZN(n17584) );
  NAND4_X1 U20757 ( .A1(n17586), .A2(n17585), .A3(n17934), .A4(n17584), .ZN(
        P3_U2808) );
  NAND2_X1 U20758 ( .A1(n17942), .A2(n17596), .ZN(n17946) );
  NAND2_X1 U20759 ( .A1(n17971), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17921) );
  INV_X1 U20760 ( .A(n17921), .ZN(n17938) );
  NAND2_X1 U20761 ( .A1(n17641), .A2(n17938), .ZN(n17622) );
  OAI22_X1 U20762 ( .A1(n18077), .A2(n18759), .B1(n17696), .B2(n17587), .ZN(
        n17588) );
  AOI221_X1 U20763 ( .B1(n17591), .B2(n17590), .C1(n17589), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17588), .ZN(n17599) );
  INV_X1 U20764 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17623) );
  NOR3_X1 U20765 ( .A1(n17623), .A2(n17645), .A3(n17592), .ZN(n17617) );
  INV_X1 U20766 ( .A(n17593), .ZN(n17630) );
  AOI22_X1 U20767 ( .A1(n17942), .A2(n17617), .B1(n17630), .B2(n17594), .ZN(
        n17595) );
  XOR2_X1 U20768 ( .A(n17596), .B(n17595), .Z(n17937) );
  AOI22_X1 U20769 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17597), .B1(
        n17768), .B2(n17937), .ZN(n17598) );
  OAI211_X1 U20770 ( .C1(n17946), .C2(n17622), .A(n17599), .B(n17598), .ZN(
        P3_U2809) );
  NAND2_X1 U20771 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17608), .ZN(
        n17957) );
  AOI21_X1 U20772 ( .B1(n9798), .B2(n18215), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17601) );
  OAI22_X1 U20773 ( .A1(n17602), .A2(n17601), .B1(n18077), .B2(n18756), .ZN(
        n17603) );
  AOI221_X1 U20774 ( .B1(n17706), .B2(n17604), .C1(n16366), .C2(n17604), .A(
        n17603), .ZN(n17610) );
  NOR2_X1 U20775 ( .A1(n17964), .A2(n17921), .ZN(n17948) );
  OAI21_X1 U20776 ( .B1(n17605), .B2(n17948), .A(n17657), .ZN(n17619) );
  OAI221_X1 U20777 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17629), 
        .C1(n17964), .C2(n17617), .A(n17606), .ZN(n17607) );
  XOR2_X1 U20778 ( .A(n17608), .B(n17607), .Z(n17953) );
  AOI22_X1 U20779 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17619), .B1(
        n17768), .B2(n17953), .ZN(n17609) );
  OAI211_X1 U20780 ( .C1(n17622), .C2(n17957), .A(n17610), .B(n17609), .ZN(
        P3_U2810) );
  AOI21_X1 U20781 ( .B1(n17810), .B2(n17612), .A(n17845), .ZN(n17637) );
  OAI21_X1 U20782 ( .B1(n17611), .B2(n18702), .A(n17637), .ZN(n17626) );
  NOR2_X1 U20783 ( .A1(n17691), .A2(n17612), .ZN(n17628) );
  OAI211_X1 U20784 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17628), .B(n17613), .ZN(n17614) );
  NAND2_X1 U20785 ( .A1(n9654), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17961) );
  OAI211_X1 U20786 ( .C1(n17696), .C2(n17615), .A(n17614), .B(n17961), .ZN(
        n17616) );
  AOI21_X1 U20787 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17626), .A(
        n17616), .ZN(n17621) );
  AOI21_X1 U20788 ( .B1(n17629), .B2(n17630), .A(n17617), .ZN(n17618) );
  XOR2_X1 U20789 ( .A(n17964), .B(n17618), .Z(n17960) );
  AOI22_X1 U20790 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17619), .B1(
        n17768), .B2(n17960), .ZN(n17620) );
  OAI211_X1 U20791 ( .C1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n17622), .A(
        n17621), .B(n17620), .ZN(P3_U2811) );
  NAND2_X1 U20792 ( .A1(n17971), .A2(n17623), .ZN(n17978) );
  OAI22_X1 U20793 ( .A1(n18077), .A2(n18752), .B1(n17696), .B2(n17624), .ZN(
        n17625) );
  AOI221_X1 U20794 ( .B1(n17628), .B2(n17627), .C1(n17626), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17625), .ZN(n17633) );
  OAI21_X1 U20795 ( .B1(n17971), .B2(n17658), .A(n17657), .ZN(n17640) );
  AOI21_X1 U20796 ( .B1(n17767), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17629), .ZN(n17631) );
  XOR2_X1 U20797 ( .A(n17631), .B(n17630), .Z(n17974) );
  AOI22_X1 U20798 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17640), .B1(
        n17768), .B2(n17974), .ZN(n17632) );
  OAI211_X1 U20799 ( .C1(n17658), .C2(n17978), .A(n17633), .B(n17632), .ZN(
        P3_U2812) );
  OAI21_X1 U20800 ( .B1(n17635), .B2(n17979), .A(n17634), .ZN(n17983) );
  AOI21_X1 U20801 ( .B1(n17636), .B2(n18566), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17638) );
  OAI22_X1 U20802 ( .A1(n17638), .A2(n17637), .B1(n18077), .B2(n18750), .ZN(
        n17639) );
  AOI21_X1 U20803 ( .B1(n17768), .B2(n17983), .A(n17639), .ZN(n17643) );
  OAI221_X1 U20804 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17641), .A(n17640), .ZN(
        n17642) );
  OAI211_X1 U20805 ( .C1(n17842), .C2(n17644), .A(n17643), .B(n17642), .ZN(
        P3_U2813) );
  INV_X1 U20806 ( .A(n17744), .ZN(n17718) );
  OAI21_X1 U20807 ( .B1(n17647), .B2(n17718), .A(n17646), .ZN(n17648) );
  XOR2_X1 U20808 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17648), .Z(
        n17992) );
  AOI21_X1 U20809 ( .B1(n17810), .B2(n17650), .A(n17845), .ZN(n17677) );
  OAI21_X1 U20810 ( .B1(n17649), .B2(n18702), .A(n17677), .ZN(n17661) );
  AOI22_X1 U20811 ( .A1(n9654), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17661), .ZN(n17653) );
  NOR2_X1 U20812 ( .A1(n17691), .A2(n17650), .ZN(n17663) );
  OAI211_X1 U20813 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17663), .B(n17651), .ZN(n17652) );
  OAI211_X1 U20814 ( .C1(n17696), .C2(n17654), .A(n17653), .B(n17652), .ZN(
        n17655) );
  AOI21_X1 U20815 ( .B1(n17768), .B2(n17992), .A(n17655), .ZN(n17656) );
  OAI221_X1 U20816 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17658), 
        .C1(n17995), .C2(n17657), .A(n17656), .ZN(P3_U2814) );
  NOR2_X1 U20817 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17679), .ZN(
        n17997) );
  NAND2_X1 U20818 ( .A1(n17770), .A2(n17920), .ZN(n17672) );
  INV_X1 U20819 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17662) );
  OAI22_X1 U20820 ( .A1(n18077), .A2(n18746), .B1(n17696), .B2(n17659), .ZN(
        n17660) );
  AOI221_X1 U20821 ( .B1(n17663), .B2(n17662), .C1(n17661), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17660), .ZN(n17671) );
  INV_X1 U20822 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18039) );
  AND2_X1 U20823 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17664) );
  NAND3_X1 U20824 ( .A1(n18027), .A2(n17664), .A3(n18050), .ZN(n17665) );
  NAND2_X1 U20825 ( .A1(n17666), .A2(n17665), .ZN(n17667) );
  OAI221_X1 U20826 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18026), 
        .C1(n18039), .C2(n17767), .A(n17667), .ZN(n17668) );
  XOR2_X1 U20827 ( .A(n18004), .B(n17668), .Z(n18006) );
  NOR2_X1 U20828 ( .A1(n17897), .A2(n17862), .ZN(n17669) );
  NOR2_X1 U20829 ( .A1(n17728), .A2(n18013), .ZN(n18028) );
  NAND3_X1 U20830 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n18028), .ZN(n17673) );
  NAND2_X1 U20831 ( .A1(n18004), .A2(n17673), .ZN(n18007) );
  AOI22_X1 U20832 ( .A1(n17768), .A2(n18006), .B1(n17669), .B2(n18007), .ZN(
        n17670) );
  OAI211_X1 U20833 ( .C1(n17997), .C2(n17672), .A(n17671), .B(n17670), .ZN(
        P3_U2815) );
  OAI221_X1 U20834 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18028), .A(n17673), .ZN(
        n18020) );
  AOI21_X1 U20835 ( .B1(n17674), .B2(n18566), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17676) );
  OAI22_X1 U20836 ( .A1(n17677), .A2(n17676), .B1(n17842), .B2(n17675), .ZN(
        n17678) );
  AOI21_X1 U20837 ( .B1(n9654), .B2(P3_REIP_REG_14__SCAN_IN), .A(n17678), .ZN(
        n17684) );
  NOR2_X1 U20838 ( .A1(n18013), .A2(n18015), .ZN(n17998) );
  INV_X1 U20839 ( .A(n17998), .ZN(n17680) );
  AOI221_X1 U20840 ( .B1(n17766), .B2(n18026), .C1(n17680), .C2(n18026), .A(
        n17679), .ZN(n18019) );
  AOI21_X1 U20841 ( .B1(n17744), .B2(n17998), .A(n17681), .ZN(n17682) );
  XOR2_X1 U20842 ( .A(n18026), .B(n17682), .Z(n18023) );
  AOI22_X1 U20843 ( .A1(n17770), .A2(n18019), .B1(n17768), .B2(n18023), .ZN(
        n17683) );
  OAI211_X1 U20844 ( .C1(n17862), .C2(n18020), .A(n17684), .B(n17683), .ZN(
        P3_U2816) );
  INV_X1 U20845 ( .A(n18028), .ZN(n17685) );
  NOR2_X1 U20846 ( .A1(n18013), .A2(n17766), .ZN(n17700) );
  INV_X1 U20847 ( .A(n17700), .ZN(n18030) );
  AOI22_X1 U20848 ( .A1(n17850), .A2(n17685), .B1(n17770), .B2(n18030), .ZN(
        n17709) );
  OAI21_X1 U20849 ( .B1(n17775), .B2(n17689), .A(n17858), .ZN(n17773) );
  AOI21_X1 U20850 ( .B1(n17687), .B2(n17686), .A(n17773), .ZN(n17688) );
  OAI21_X1 U20851 ( .B1(n17690), .B2(n17689), .A(n17688), .ZN(n17707) );
  NOR2_X1 U20852 ( .A1(n17691), .A2(n17721), .ZN(n17715) );
  OAI211_X1 U20853 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17715), .B(n17692), .ZN(n17694) );
  NAND2_X1 U20854 ( .A1(n9654), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17693) );
  OAI211_X1 U20855 ( .C1(n17696), .C2(n17695), .A(n17694), .B(n17693), .ZN(
        n17697) );
  AOI21_X1 U20856 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17707), .A(
        n17697), .ZN(n17703) );
  NOR2_X1 U20857 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17767), .ZN(
        n17699) );
  OAI22_X1 U20858 ( .A1(n17700), .A2(n17699), .B1(n17767), .B2(n17698), .ZN(
        n17701) );
  XOR2_X1 U20859 ( .A(n18015), .B(n17701), .Z(n18035) );
  NOR2_X1 U20860 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18013), .ZN(
        n18034) );
  INV_X1 U20861 ( .A(n17755), .ZN(n17727) );
  AOI22_X1 U20862 ( .A1(n17768), .A2(n18035), .B1(n18034), .B2(n17727), .ZN(
        n17702) );
  OAI211_X1 U20863 ( .C1(n17709), .C2(n18015), .A(n17703), .B(n17702), .ZN(
        P3_U2817) );
  AOI21_X1 U20864 ( .B1(n17744), .B2(n18027), .A(n17698), .ZN(n17704) );
  XOR2_X1 U20865 ( .A(n17704), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18047) );
  AOI22_X1 U20866 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17707), .B1(
        n17706), .B2(n17705), .ZN(n17708) );
  NAND2_X1 U20867 ( .A1(n9654), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n18045) );
  NAND2_X1 U20868 ( .A1(n17708), .A2(n18045), .ZN(n17713) );
  NOR2_X1 U20869 ( .A1(n17755), .A2(n18038), .ZN(n17711) );
  INV_X1 U20870 ( .A(n17709), .ZN(n17710) );
  MUX2_X1 U20871 ( .A(n17711), .B(n17710), .S(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n17712) );
  AOI211_X1 U20872 ( .C1(n17715), .C2(n17714), .A(n17713), .B(n17712), .ZN(
        n17716) );
  OAI21_X1 U20873 ( .B1(n18047), .B2(n17742), .A(n17716), .ZN(P3_U2818) );
  OAI21_X1 U20874 ( .B1(n17720), .B2(n17718), .A(n17717), .ZN(n17719) );
  XNOR2_X1 U20875 ( .A(n17719), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18063) );
  NOR2_X1 U20876 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17720), .ZN(
        n18048) );
  NOR2_X1 U20877 ( .A1(n18077), .A2(n18738), .ZN(n17726) );
  INV_X1 U20878 ( .A(n17793), .ZN(n17853) );
  NAND3_X1 U20879 ( .A1(n17775), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A3(
        n18566), .ZN(n17762) );
  NOR2_X1 U20880 ( .A1(n17761), .A2(n17762), .ZN(n17747) );
  NAND2_X1 U20881 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17747), .ZN(
        n17746) );
  NOR2_X1 U20882 ( .A1(n17733), .A2(n17746), .ZN(n17732) );
  AOI21_X1 U20883 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n17853), .A(
        n17732), .ZN(n17724) );
  NOR2_X1 U20884 ( .A1(n17721), .A2(n17816), .ZN(n17723) );
  OAI22_X1 U20885 ( .A1(n17724), .A2(n17723), .B1(n17842), .B2(n17722), .ZN(
        n17725) );
  AOI211_X1 U20886 ( .C1(n18048), .C2(n17727), .A(n17726), .B(n17725), .ZN(
        n17730) );
  NOR2_X1 U20887 ( .A1(n18056), .A2(n17755), .ZN(n17738) );
  AOI22_X1 U20888 ( .A1(n17766), .A2(n17770), .B1(n17850), .B2(n17728), .ZN(
        n17754) );
  INV_X1 U20889 ( .A(n17754), .ZN(n17739) );
  OAI21_X1 U20890 ( .B1(n17738), .B2(n17739), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17729) );
  OAI211_X1 U20891 ( .C1(n18063), .C2(n17742), .A(n17730), .B(n17729), .ZN(
        P3_U2819) );
  AOI22_X1 U20892 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17744), .B1(
        n17743), .B2(n18073), .ZN(n17731) );
  XOR2_X1 U20893 ( .A(n17731), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .Z(
        n18071) );
  AOI211_X1 U20894 ( .C1(n17746), .C2(n17733), .A(n17793), .B(n17732), .ZN(
        n17735) );
  INV_X1 U20895 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18736) );
  NOR2_X1 U20896 ( .A1(n18077), .A2(n18736), .ZN(n17734) );
  AOI211_X1 U20897 ( .C1(n17736), .C2(n17852), .A(n17735), .B(n17734), .ZN(
        n17741) );
  NAND2_X1 U20898 ( .A1(n18073), .A2(n18067), .ZN(n17737) );
  AOI22_X1 U20899 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17739), .B1(
        n17738), .B2(n17737), .ZN(n17740) );
  OAI211_X1 U20900 ( .C1(n18071), .C2(n17742), .A(n17741), .B(n17740), .ZN(
        P3_U2820) );
  NOR2_X1 U20901 ( .A1(n17744), .A2(n17743), .ZN(n17745) );
  XOR2_X1 U20902 ( .A(n17745), .B(n18073), .Z(n18075) );
  NOR2_X1 U20903 ( .A1(n18077), .A2(n18734), .ZN(n17752) );
  INV_X1 U20904 ( .A(n17746), .ZN(n17750) );
  AOI21_X1 U20905 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17853), .A(
        n17747), .ZN(n17749) );
  OAI22_X1 U20906 ( .A1(n17750), .A2(n17749), .B1(n17842), .B2(n17748), .ZN(
        n17751) );
  AOI211_X1 U20907 ( .C1(n17768), .C2(n18075), .A(n17752), .B(n17751), .ZN(
        n17753) );
  OAI221_X1 U20908 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17755), .C1(
        n18073), .C2(n17754), .A(n17753), .ZN(P3_U2821) );
  OAI21_X1 U20909 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17757), .A(
        n17756), .ZN(n18097) );
  INV_X1 U20910 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17758) );
  AOI21_X1 U20911 ( .B1(n18215), .B2(n17758), .A(n17773), .ZN(n17760) );
  NAND2_X1 U20912 ( .A1(n9654), .A2(P3_REIP_REG_8__SCAN_IN), .ZN(n17759) );
  OAI221_X1 U20913 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17762), .C1(
        n17761), .C2(n17760), .A(n17759), .ZN(n17763) );
  AOI21_X1 U20914 ( .B1(n17764), .B2(n17852), .A(n17763), .ZN(n17772) );
  NAND2_X1 U20915 ( .A1(n17766), .A2(n17765), .ZN(n18090) );
  INV_X1 U20916 ( .A(n18090), .ZN(n17769) );
  XOR2_X1 U20917 ( .A(n17767), .B(n18090), .Z(n18092) );
  AOI22_X1 U20918 ( .A1(n17770), .A2(n17769), .B1(n17768), .B2(n18092), .ZN(
        n17771) );
  OAI211_X1 U20919 ( .C1(n17862), .C2(n18097), .A(n17772), .B(n17771), .ZN(
        P3_U2822) );
  NOR2_X1 U20920 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17816), .ZN(
        n17774) );
  AOI22_X1 U20921 ( .A1(n17775), .A2(n17774), .B1(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n17773), .ZN(n17785) );
  AOI21_X1 U20922 ( .B1(n17778), .B2(n17777), .A(n17776), .ZN(n17779) );
  XOR2_X1 U20923 ( .A(n17779), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18103) );
  OAI21_X1 U20924 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17781), .A(
        n17780), .ZN(n18099) );
  OAI22_X1 U20925 ( .A1(n17842), .A2(n17782), .B1(n17861), .B2(n18099), .ZN(
        n17783) );
  AOI21_X1 U20926 ( .B1(n17850), .B2(n18103), .A(n17783), .ZN(n17784) );
  OAI211_X1 U20927 ( .C1(n18077), .C2(n18730), .A(n17785), .B(n17784), .ZN(
        P3_U2823) );
  OAI21_X1 U20928 ( .B1(n17787), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n17786), .ZN(n18114) );
  NAND2_X1 U20929 ( .A1(n17794), .A2(n18566), .ZN(n17791) );
  OAI21_X1 U20930 ( .B1(n17790), .B2(n17789), .A(n17788), .ZN(n18109) );
  OAI22_X1 U20931 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17791), .B1(
        n17861), .B2(n18109), .ZN(n17792) );
  AOI21_X1 U20932 ( .B1(n9654), .B2(P3_REIP_REG_6__SCAN_IN), .A(n17792), .ZN(
        n17797) );
  AOI21_X1 U20933 ( .B1(n18566), .B2(n17794), .A(n17793), .ZN(n17805) );
  AOI22_X1 U20934 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17805), .B1(
        n17795), .B2(n17852), .ZN(n17796) );
  OAI211_X1 U20935 ( .C1(n17862), .C2(n18114), .A(n17797), .B(n17796), .ZN(
        P3_U2824) );
  OAI21_X1 U20936 ( .B1(n17800), .B2(n17799), .A(n17798), .ZN(n18123) );
  OAI21_X1 U20937 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n17802), .A(
        n17801), .ZN(n18116) );
  INV_X1 U20938 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18727) );
  OAI22_X1 U20939 ( .A1(n17861), .A2(n18116), .B1(n18077), .B2(n18727), .ZN(
        n17803) );
  AOI21_X1 U20940 ( .B1(n17804), .B2(n17852), .A(n17803), .ZN(n17808) );
  OAI221_X1 U20941 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17806), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n17858), .A(n17805), .ZN(n17807) );
  OAI211_X1 U20942 ( .C1(n17862), .C2(n18123), .A(n17808), .B(n17807), .ZN(
        P3_U2825) );
  AOI21_X1 U20943 ( .B1(n17810), .B2(n17809), .A(n17845), .ZN(n17831) );
  OAI21_X1 U20944 ( .B1(n17813), .B2(n17812), .A(n17811), .ZN(n17814) );
  XOR2_X1 U20945 ( .A(n17814), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18124) );
  OAI22_X1 U20946 ( .A1(n17862), .A2(n18124), .B1(n17816), .B2(n17815), .ZN(
        n17822) );
  OAI21_X1 U20947 ( .B1(n17819), .B2(n17818), .A(n17817), .ZN(n18130) );
  OAI22_X1 U20948 ( .A1(n17842), .A2(n17820), .B1(n17861), .B2(n18130), .ZN(
        n17821) );
  AOI211_X1 U20949 ( .C1(n9654), .C2(P3_REIP_REG_4__SCAN_IN), .A(n17822), .B(
        n17821), .ZN(n17823) );
  OAI21_X1 U20950 ( .B1(n17831), .B2(n17824), .A(n17823), .ZN(P3_U2826) );
  OAI21_X1 U20951 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17826), .A(
        n17825), .ZN(n18135) );
  AOI21_X1 U20952 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17858), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17830) );
  OAI21_X1 U20953 ( .B1(n17829), .B2(n17828), .A(n17827), .ZN(n18139) );
  OAI22_X1 U20954 ( .A1(n17831), .A2(n17830), .B1(n17862), .B2(n18139), .ZN(
        n17832) );
  AOI21_X1 U20955 ( .B1(n17833), .B2(n17852), .A(n17832), .ZN(n17834) );
  NAND2_X1 U20956 ( .A1(n9654), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18134) );
  OAI211_X1 U20957 ( .C1(n17861), .C2(n18135), .A(n17834), .B(n18134), .ZN(
        P3_U2827) );
  OAI21_X1 U20958 ( .B1(n17837), .B2(n17836), .A(n17835), .ZN(n18156) );
  OAI21_X1 U20959 ( .B1(n17840), .B2(n17839), .A(n17838), .ZN(n18151) );
  OAI22_X1 U20960 ( .A1(n17842), .A2(n17841), .B1(n17862), .B2(n18151), .ZN(
        n17843) );
  AOI221_X1 U20961 ( .B1(n17845), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18566), .C2(n17844), .A(n17843), .ZN(n17846) );
  NAND2_X1 U20962 ( .A1(n9654), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18154) );
  OAI211_X1 U20963 ( .C1(n17861), .C2(n18156), .A(n17846), .B(n18154), .ZN(
        P3_U2828) );
  OAI21_X1 U20964 ( .B1(n17848), .B2(n17856), .A(n17847), .ZN(n18167) );
  NAND2_X1 U20965 ( .A1(n18817), .A2(n17857), .ZN(n17849) );
  XNOR2_X1 U20966 ( .A(n17849), .B(n17848), .ZN(n18163) );
  AOI22_X1 U20967 ( .A1(n17850), .A2(n18163), .B1(n9654), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17855) );
  AOI22_X1 U20968 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17853), .B1(
        n17852), .B2(n17851), .ZN(n17854) );
  OAI211_X1 U20969 ( .C1(n17861), .C2(n18167), .A(n17855), .B(n17854), .ZN(
        P3_U2829) );
  AOI21_X1 U20970 ( .B1(n17857), .B2(n18817), .A(n17856), .ZN(n18171) );
  INV_X1 U20971 ( .A(n18171), .ZN(n18169) );
  NAND3_X1 U20972 ( .A1(n18800), .A2(n18702), .A3(n17858), .ZN(n17859) );
  AOI22_X1 U20973 ( .A1(n9654), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17859), .ZN(n17860) );
  OAI221_X1 U20974 ( .B1(n18171), .B2(n17862), .C1(n18169), .C2(n17861), .A(
        n17860), .ZN(P3_U2830) );
  AOI21_X1 U20975 ( .B1(n17863), .B2(n9931), .A(n18173), .ZN(n17873) );
  INV_X1 U20976 ( .A(n17968), .ZN(n17865) );
  OAI211_X1 U20977 ( .C1(n18059), .C2(n17987), .A(n17932), .B(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17864) );
  INV_X1 U20978 ( .A(n18143), .ZN(n18082) );
  OAI21_X1 U20979 ( .B1(n17865), .B2(n17864), .A(n18082), .ZN(n17901) );
  OAI221_X1 U20980 ( .B1(n18143), .B2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), 
        .C1(n18143), .C2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A(n17901), .ZN(
        n17883) );
  OAI22_X1 U20981 ( .A1(n18646), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n18059), .B2(n17866), .ZN(n17870) );
  OAI22_X1 U20982 ( .A1(n17868), .A2(n18627), .B1(n17867), .B2(n18091), .ZN(
        n17869) );
  NOR4_X1 U20983 ( .A1(n17871), .A2(n17883), .A3(n17870), .A4(n17869), .ZN(
        n17877) );
  OAI211_X1 U20984 ( .C1(n18646), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17877), .ZN(n17872) );
  AOI22_X1 U20985 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18153), .B1(
        n17873), .B2(n17872), .ZN(n17875) );
  NAND2_X1 U20986 ( .A1(n9654), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17874) );
  OAI211_X1 U20987 ( .C1(n17876), .C2(n18070), .A(n17875), .B(n17874), .ZN(
        P3_U2835) );
  AOI22_X1 U20988 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18153), .B1(
        n9654), .B2(P3_REIP_REG_26__SCAN_IN), .ZN(n17881) );
  NOR2_X1 U20989 ( .A1(n17877), .A2(n18173), .ZN(n17879) );
  AOI22_X1 U20990 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17879), .B1(
        n17936), .B2(n17878), .ZN(n17880) );
  OAI211_X1 U20991 ( .C1(n17882), .C2(n18070), .A(n17881), .B(n17880), .ZN(
        P3_U2836) );
  INV_X1 U20992 ( .A(n17903), .ZN(n17969) );
  AOI221_X1 U20993 ( .B1(n18635), .B2(n17884), .C1(n18635), .C2(n17969), .A(
        n17883), .ZN(n17885) );
  INV_X1 U20994 ( .A(n17885), .ZN(n17889) );
  OAI22_X1 U20995 ( .A1(n18627), .A2(n17887), .B1(n18091), .B2(n17886), .ZN(
        n17888) );
  AOI221_X1 U20996 ( .B1(n17890), .B2(n17892), .C1(n17889), .C2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(n17888), .ZN(n17896) );
  OAI22_X1 U20997 ( .A1(n17892), .A2(n18159), .B1(n18070), .B2(n17891), .ZN(
        n17893) );
  INV_X1 U20998 ( .A(n17893), .ZN(n17895) );
  OAI211_X1 U20999 ( .C1(n17896), .C2(n18173), .A(n17895), .B(n17894), .ZN(
        P3_U2837) );
  INV_X1 U21000 ( .A(n17990), .ZN(n18085) );
  NAND2_X1 U21001 ( .A1(n17897), .A2(n17898), .ZN(n17900) );
  NAND2_X1 U21002 ( .A1(n17898), .A2(n17577), .ZN(n17899) );
  AOI22_X1 U21003 ( .A1(n17923), .A2(n17900), .B1(n18031), .B2(n17899), .ZN(
        n17902) );
  NAND3_X1 U21004 ( .A1(n17902), .A2(n18159), .A3(n17901), .ZN(n17905) );
  INV_X1 U21005 ( .A(n17905), .ZN(n17907) );
  OAI221_X1 U21006 ( .B1(n18662), .B2(n17913), .C1(n18662), .C2(n17903), .A(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17904) );
  OAI21_X1 U21007 ( .B1(n17905), .B2(n17904), .A(n18077), .ZN(n17919) );
  AOI211_X1 U21008 ( .C1(n18085), .C2(n17907), .A(n17906), .B(n17919), .ZN(
        n17908) );
  AOI211_X1 U21009 ( .C1(n17910), .C2(n17936), .A(n17909), .B(n17908), .ZN(
        n17911) );
  OAI21_X1 U21010 ( .B1(n17912), .B2(n18070), .A(n17911), .ZN(P3_U2838) );
  NAND3_X1 U21011 ( .A1(n17913), .A2(n18159), .A3(n17931), .ZN(n17917) );
  AOI21_X1 U21012 ( .B1(n17915), .B2(n18093), .A(n17914), .ZN(n17916) );
  OAI221_X1 U21013 ( .B1(n17919), .B2(n17918), .C1(n17919), .C2(n17917), .A(
        n17916), .ZN(P3_U2839) );
  OAI221_X1 U21014 ( .B1(n18059), .B2(n17932), .C1(n18059), .C2(n17987), .A(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17927) );
  OAI22_X1 U21015 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18064), .B1(
        n17942), .B2(n18662), .ZN(n17926) );
  AOI22_X1 U21016 ( .A1(n17923), .A2(n18008), .B1(n18031), .B2(n17920), .ZN(
        n17939) );
  OAI21_X1 U21017 ( .B1(n17969), .B2(n17921), .A(n18635), .ZN(n17922) );
  OAI221_X1 U21018 ( .B1(n18646), .B2(n17968), .C1(n18646), .C2(n17948), .A(
        n17922), .ZN(n17950) );
  NOR2_X1 U21019 ( .A1(n17923), .A2(n18031), .ZN(n18055) );
  OAI22_X1 U21020 ( .A1(n18646), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17932), .B2(n18055), .ZN(n17924) );
  NOR2_X1 U21021 ( .A1(n17950), .A2(n17924), .ZN(n17941) );
  NAND2_X1 U21022 ( .A1(n17939), .A2(n17941), .ZN(n17925) );
  NOR3_X1 U21023 ( .A1(n17927), .A2(n17926), .A3(n17925), .ZN(n17929) );
  OAI22_X1 U21024 ( .A1(n17929), .A2(n18173), .B1(n17928), .B2(n18159), .ZN(
        n17930) );
  OAI221_X1 U21025 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17932), 
        .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17931), .A(n17930), .ZN(
        n17933) );
  OAI211_X1 U21026 ( .C1(n17935), .C2(n18070), .A(n17934), .B(n17933), .ZN(
        P3_U2840) );
  NAND2_X1 U21027 ( .A1(n17936), .A2(n17938), .ZN(n17958) );
  AOI22_X1 U21028 ( .A1(n9654), .A2(P3_REIP_REG_21__SCAN_IN), .B1(n18093), 
        .B2(n17937), .ZN(n17945) );
  NAND2_X1 U21029 ( .A1(n18662), .A2(n18059), .ZN(n18157) );
  INV_X1 U21030 ( .A(n18157), .ZN(n17952) );
  AOI21_X1 U21031 ( .B1(n17987), .B2(n17938), .A(n18059), .ZN(n17940) );
  NAND2_X1 U21032 ( .A1(n18158), .A2(n17939), .ZN(n17991) );
  NOR2_X1 U21033 ( .A1(n17940), .A2(n17991), .ZN(n17947) );
  OAI211_X1 U21034 ( .C1(n17942), .C2(n17952), .A(n17941), .B(n17947), .ZN(
        n17943) );
  NAND3_X1 U21035 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n18077), .A3(
        n17943), .ZN(n17944) );
  OAI211_X1 U21036 ( .C1(n17958), .C2(n17946), .A(n17945), .B(n17944), .ZN(
        P3_U2841) );
  NAND2_X1 U21037 ( .A1(n17964), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17951) );
  OAI21_X1 U21038 ( .B1(n17948), .B2(n18055), .A(n17947), .ZN(n17949) );
  OAI21_X1 U21039 ( .B1(n17950), .B2(n17949), .A(n18077), .ZN(n17963) );
  OAI21_X1 U21040 ( .B1(n17952), .B2(n17951), .A(n17963), .ZN(n17954) );
  AOI22_X1 U21041 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17954), .B1(
        n18093), .B2(n17953), .ZN(n17956) );
  NAND2_X1 U21042 ( .A1(n9654), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17955) );
  OAI211_X1 U21043 ( .C1(n17957), .C2(n17958), .A(n17956), .B(n17955), .ZN(
        P3_U2842) );
  INV_X1 U21044 ( .A(n17958), .ZN(n17959) );
  AOI22_X1 U21045 ( .A1(n18093), .A2(n17960), .B1(n17959), .B2(n17964), .ZN(
        n17962) );
  OAI211_X1 U21046 ( .C1(n17964), .C2(n17963), .A(n17962), .B(n17961), .ZN(
        P3_U2843) );
  AOI22_X1 U21047 ( .A1(n18635), .A2(n18144), .B1(n18148), .B2(n18079), .ZN(
        n18133) );
  NOR2_X1 U21048 ( .A1(n18133), .A2(n17965), .ZN(n17999) );
  NOR2_X1 U21049 ( .A1(n17999), .A2(n17966), .ZN(n18040) );
  NAND2_X1 U21050 ( .A1(n17967), .A2(n18074), .ZN(n17996) );
  NAND2_X1 U21051 ( .A1(n18656), .A2(n18817), .ZN(n18141) );
  NAND3_X1 U21052 ( .A1(n17968), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18141), .ZN(n17973) );
  NAND2_X1 U21053 ( .A1(n18635), .A2(n17969), .ZN(n17970) );
  AOI22_X1 U21054 ( .A1(n17971), .A2(n17970), .B1(n18055), .B2(n18662), .ZN(
        n17972) );
  AOI211_X1 U21055 ( .C1(n18082), .C2(n17973), .A(n17972), .B(n17991), .ZN(
        n17980) );
  AOI221_X1 U21056 ( .B1(n18143), .B2(n17980), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17980), .A(n9654), .ZN(
        n17975) );
  AOI22_X1 U21057 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17975), .B1(
        n18093), .B2(n17974), .ZN(n17977) );
  NAND2_X1 U21058 ( .A1(n9654), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17976) );
  OAI211_X1 U21059 ( .C1(n17978), .C2(n17996), .A(n17977), .B(n17976), .ZN(
        P3_U2844) );
  NOR3_X1 U21060 ( .A1(n9654), .A2(n17980), .A3(n17979), .ZN(n17982) );
  NOR3_X1 U21061 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17995), .A3(
        n17996), .ZN(n17981) );
  AOI211_X1 U21062 ( .C1(n18093), .C2(n17983), .A(n17982), .B(n17981), .ZN(
        n17984) );
  OAI21_X1 U21063 ( .B1(n18077), .B2(n18750), .A(n17984), .ZN(P3_U2845) );
  AOI22_X1 U21064 ( .A1(n18635), .A2(n17986), .B1(n18633), .B2(n17985), .ZN(
        n18054) );
  AOI21_X1 U21065 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18059), .A(
        n17987), .ZN(n17988) );
  INV_X1 U21066 ( .A(n17988), .ZN(n17989) );
  OAI211_X1 U21067 ( .C1(n18012), .C2(n18064), .A(n18054), .B(n17989), .ZN(
        n18001) );
  OAI221_X1 U21068 ( .B1(n17991), .B2(n17990), .C1(n17991), .C2(n18001), .A(
        n18077), .ZN(n17994) );
  AOI22_X1 U21069 ( .A1(n9654), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18093), 
        .B2(n17992), .ZN(n17993) );
  OAI221_X1 U21070 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17996), 
        .C1(n17995), .C2(n17994), .A(n17993), .ZN(P3_U2846) );
  NOR2_X1 U21071 ( .A1(n17577), .A2(n18091), .ZN(n18003) );
  INV_X1 U21072 ( .A(n17997), .ZN(n18002) );
  NAND2_X1 U21073 ( .A1(n17999), .A2(n17998), .ZN(n18016) );
  OAI21_X1 U21074 ( .B1(n18026), .B2(n18016), .A(n18004), .ZN(n18000) );
  AOI22_X1 U21075 ( .A1(n18003), .A2(n18002), .B1(n18001), .B2(n18000), .ZN(
        n18011) );
  OAI22_X1 U21076 ( .A1(n18004), .A2(n18159), .B1(n18077), .B2(n18746), .ZN(
        n18005) );
  AOI21_X1 U21077 ( .B1(n18093), .B2(n18006), .A(n18005), .ZN(n18010) );
  NAND3_X1 U21078 ( .A1(n18170), .A2(n18008), .A3(n18007), .ZN(n18009) );
  OAI211_X1 U21079 ( .C1(n18011), .C2(n18173), .A(n18010), .B(n18009), .ZN(
        P3_U2847) );
  AOI21_X1 U21080 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18064), .A(
        n18012), .ZN(n18014) );
  NOR2_X1 U21081 ( .A1(n18013), .A2(n18052), .ZN(n18042) );
  NOR2_X1 U21082 ( .A1(n18059), .A2(n18042), .ZN(n18033) );
  AOI211_X1 U21083 ( .C1(n18015), .C2(n18157), .A(n18014), .B(n18033), .ZN(
        n18017) );
  AOI22_X1 U21084 ( .A1(n18017), .A2(n18054), .B1(n18026), .B2(n18016), .ZN(
        n18018) );
  AOI21_X1 U21085 ( .B1(n18019), .B2(n18031), .A(n18018), .ZN(n18021) );
  OAI22_X1 U21086 ( .A1(n18021), .A2(n18173), .B1(n18140), .B2(n18020), .ZN(
        n18022) );
  AOI21_X1 U21087 ( .B1(n18093), .B2(n18023), .A(n18022), .ZN(n18025) );
  NAND2_X1 U21088 ( .A1(n9654), .A2(P3_REIP_REG_14__SCAN_IN), .ZN(n18024) );
  OAI211_X1 U21089 ( .C1(n18159), .C2(n18026), .A(n18025), .B(n18024), .ZN(
        P3_U2848) );
  OR2_X1 U21090 ( .A1(n18027), .A2(n18064), .ZN(n18058) );
  OAI211_X1 U21091 ( .C1(n18028), .C2(n18627), .A(n18054), .B(n18058), .ZN(
        n18029) );
  AOI21_X1 U21092 ( .B1(n18031), .B2(n18030), .A(n18029), .ZN(n18041) );
  OAI211_X1 U21093 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18064), .A(
        n18158), .B(n18041), .ZN(n18032) );
  OAI21_X1 U21094 ( .B1(n18033), .B2(n18032), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n18037) );
  AOI22_X1 U21095 ( .A1(n18093), .A2(n18035), .B1(n18074), .B2(n18034), .ZN(
        n18036) );
  OAI221_X1 U21096 ( .B1(n9654), .B2(n18037), .C1(n18077), .C2(n18742), .A(
        n18036), .ZN(P3_U2849) );
  AOI221_X1 U21097 ( .B1(n18040), .B2(n18039), .C1(n18038), .C2(n18039), .A(
        n18173), .ZN(n18044) );
  OAI211_X1 U21098 ( .C1(n18042), .C2(n18059), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n18041), .ZN(n18043) );
  AOI22_X1 U21099 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18153), .B1(
        n18044), .B2(n18043), .ZN(n18046) );
  OAI211_X1 U21100 ( .C1(n18047), .C2(n18070), .A(n18046), .B(n18045), .ZN(
        P3_U2850) );
  AOI22_X1 U21101 ( .A1(n9654), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18074), 
        .B2(n18048), .ZN(n18062) );
  OAI22_X1 U21102 ( .A1(n18050), .A2(n18091), .B1(n18627), .B2(n18049), .ZN(
        n18051) );
  AOI211_X1 U21103 ( .C1(n18656), .C2(n18052), .A(n18173), .B(n18051), .ZN(
        n18053) );
  NAND2_X1 U21104 ( .A1(n18054), .A2(n18053), .ZN(n18072) );
  OAI22_X1 U21105 ( .A1(n18059), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n18056), .B2(n18055), .ZN(n18057) );
  NOR2_X1 U21106 ( .A1(n18072), .A2(n18057), .ZN(n18065) );
  OAI211_X1 U21107 ( .C1(n18059), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18065), .B(n18058), .ZN(n18060) );
  NAND3_X1 U21108 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18077), .A3(
        n18060), .ZN(n18061) );
  OAI211_X1 U21109 ( .C1(n18063), .C2(n18070), .A(n18062), .B(n18061), .ZN(
        P3_U2851) );
  AOI221_X1 U21110 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18065), .C1(
        n18064), .C2(n18065), .A(n18067), .ZN(n18066) );
  AOI22_X1 U21111 ( .A1(n9654), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18066), 
        .B2(n18077), .ZN(n18069) );
  NAND3_X1 U21112 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18074), .A3(
        n18067), .ZN(n18068) );
  OAI211_X1 U21113 ( .C1(n18071), .C2(n18070), .A(n18069), .B(n18068), .ZN(
        P3_U2852) );
  NAND2_X1 U21114 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18072), .ZN(
        n18078) );
  AOI22_X1 U21115 ( .A1(n18093), .A2(n18075), .B1(n18074), .B2(n18073), .ZN(
        n18076) );
  OAI221_X1 U21116 ( .B1(n9654), .B2(n18078), .C1(n18077), .C2(n18734), .A(
        n18076), .ZN(P3_U2853) );
  INV_X1 U21117 ( .A(n18079), .ZN(n18081) );
  OAI211_X1 U21118 ( .C1(n18662), .C2(n18144), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18141), .ZN(n18080) );
  AOI21_X1 U21119 ( .B1(n18082), .B2(n18081), .A(n18080), .ZN(n18131) );
  NOR2_X1 U21120 ( .A1(n18131), .A2(n18160), .ZN(n18127) );
  NOR2_X1 U21121 ( .A1(n18117), .A2(n20931), .ZN(n18083) );
  AOI21_X1 U21122 ( .B1(n18083), .B2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n18160), .ZN(n18084) );
  AOI211_X1 U21123 ( .C1(n18158), .C2(n18106), .A(n18127), .B(n18084), .ZN(
        n18101) );
  OAI21_X1 U21124 ( .B1(n18085), .B2(n18101), .A(n18159), .ZN(n18086) );
  AOI22_X1 U21125 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18086), .B1(
        n9654), .B2(P3_REIP_REG_8__SCAN_IN), .ZN(n18096) );
  INV_X1 U21126 ( .A(n18133), .ZN(n18115) );
  NAND2_X1 U21127 ( .A1(n18087), .A2(n18115), .ZN(n18107) );
  NAND3_X1 U21128 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n18088), .ZN(n18089) );
  OAI22_X1 U21129 ( .A1(n18091), .A2(n18090), .B1(n18107), .B2(n18089), .ZN(
        n18094) );
  AOI22_X1 U21130 ( .A1(n18158), .A2(n18094), .B1(n18093), .B2(n18092), .ZN(
        n18095) );
  OAI211_X1 U21131 ( .C1(n18140), .C2(n18097), .A(n18096), .B(n18095), .ZN(
        P3_U2854) );
  INV_X1 U21132 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18110) );
  OAI21_X1 U21133 ( .B1(n18110), .B2(n18107), .A(n18106), .ZN(n18098) );
  INV_X1 U21134 ( .A(n18098), .ZN(n18100) );
  OAI22_X1 U21135 ( .A1(n18101), .A2(n18100), .B1(n18166), .B2(n18099), .ZN(
        n18102) );
  AOI21_X1 U21136 ( .B1(n18170), .B2(n18103), .A(n18102), .ZN(n18105) );
  NAND2_X1 U21137 ( .A1(n9654), .A2(P3_REIP_REG_7__SCAN_IN), .ZN(n18104) );
  OAI211_X1 U21138 ( .C1(n18159), .C2(n18106), .A(n18105), .B(n18104), .ZN(
        P3_U2855) );
  NOR3_X1 U21139 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18173), .A3(
        n18107), .ZN(n18112) );
  AOI21_X1 U21140 ( .B1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n18160), .ZN(n18108) );
  NOR3_X1 U21141 ( .A1(n18153), .A2(n18127), .A3(n18108), .ZN(n18118) );
  OAI22_X1 U21142 ( .A1(n18118), .A2(n18110), .B1(n18166), .B2(n18109), .ZN(
        n18111) );
  AOI211_X1 U21143 ( .C1(P3_REIP_REG_6__SCAN_IN), .C2(n9654), .A(n18112), .B(
        n18111), .ZN(n18113) );
  OAI21_X1 U21144 ( .B1(n18140), .B2(n18114), .A(n18113), .ZN(P3_U2856) );
  NAND3_X1 U21145 ( .A1(n18158), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18115), .ZN(n18125) );
  NOR2_X1 U21146 ( .A1(n18125), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n18120) );
  OAI22_X1 U21147 ( .A1(n18118), .A2(n18117), .B1(n18166), .B2(n18116), .ZN(
        n18119) );
  AOI21_X1 U21148 ( .B1(n18120), .B2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n18119), .ZN(n18122) );
  NAND2_X1 U21149 ( .A1(n9654), .A2(P3_REIP_REG_5__SCAN_IN), .ZN(n18121) );
  OAI211_X1 U21150 ( .C1(n18123), .C2(n18140), .A(n18122), .B(n18121), .ZN(
        P3_U2857) );
  OAI22_X1 U21151 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18125), .B1(
        n18124), .B2(n18140), .ZN(n18126) );
  AOI221_X1 U21152 ( .B1(n18153), .B2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(
        n18127), .C2(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n18126), .ZN(
        n18129) );
  NAND2_X1 U21153 ( .A1(n9654), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n18128) );
  OAI211_X1 U21154 ( .C1(n18130), .C2(n18166), .A(n18129), .B(n18128), .ZN(
        P3_U2858) );
  AOI211_X1 U21155 ( .C1(n18133), .C2(n18132), .A(n18131), .B(n18173), .ZN(
        n18137) );
  OAI21_X1 U21156 ( .B1(n18166), .B2(n18135), .A(n18134), .ZN(n18136) );
  AOI211_X1 U21157 ( .C1(n18153), .C2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n18137), .B(n18136), .ZN(n18138) );
  OAI21_X1 U21158 ( .B1(n18140), .B2(n18139), .A(n18138), .ZN(P3_U2859) );
  NAND3_X1 U21159 ( .A1(n18635), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18142) );
  OAI211_X1 U21160 ( .C1(n18143), .C2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n18142), .B(n18141), .ZN(n18146) );
  NOR2_X1 U21161 ( .A1(n18662), .A2(n18144), .ZN(n18145) );
  AOI21_X1 U21162 ( .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18146), .A(
        n18145), .ZN(n18150) );
  NAND3_X1 U21163 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18148), .A3(
        n18147), .ZN(n18149) );
  OAI211_X1 U21164 ( .C1(n18151), .C2(n18627), .A(n18150), .B(n18149), .ZN(
        n18152) );
  AOI22_X1 U21165 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18153), .B1(
        n18158), .B2(n18152), .ZN(n18155) );
  OAI211_X1 U21166 ( .C1(n18166), .C2(n18156), .A(n18155), .B(n18154), .ZN(
        P3_U2860) );
  NAND3_X1 U21167 ( .A1(n18158), .A2(n18817), .A3(n18157), .ZN(n18175) );
  AOI21_X1 U21168 ( .B1(n18159), .B2(n18175), .A(n18801), .ZN(n18162) );
  AOI211_X1 U21169 ( .C1(n18646), .C2(n18817), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18160), .ZN(n18161) );
  AOI211_X1 U21170 ( .C1(n18170), .C2(n18163), .A(n18162), .B(n18161), .ZN(
        n18165) );
  NAND2_X1 U21171 ( .A1(n9654), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18164) );
  OAI211_X1 U21172 ( .C1(n18167), .C2(n18166), .A(n18165), .B(n18164), .ZN(
        P3_U2861) );
  INV_X1 U21173 ( .A(P3_REIP_REG_0__SCAN_IN), .ZN(n18828) );
  NOR2_X1 U21174 ( .A1(n18077), .A2(n18828), .ZN(n18168) );
  AOI221_X1 U21175 ( .B1(n18172), .B2(n18171), .C1(n18170), .C2(n18169), .A(
        n18168), .ZN(n18176) );
  OAI211_X1 U21176 ( .C1(n18633), .C2(n18173), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18077), .ZN(n18174) );
  NAND3_X1 U21177 ( .A1(n18176), .A2(n18175), .A3(n18174), .ZN(P3_U2862) );
  INV_X1 U21178 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18469) );
  AOI211_X1 U21179 ( .C1(n18178), .C2(n18177), .A(n18851), .B(n18800), .ZN(
        n18684) );
  OAI21_X1 U21180 ( .B1(n18684), .B2(n18223), .A(n18183), .ZN(n18179) );
  OAI221_X1 U21181 ( .B1(n18469), .B2(n18837), .C1(n18469), .C2(n18183), .A(
        n18179), .ZN(P3_U2863) );
  INV_X1 U21182 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18673) );
  NAND2_X1 U21183 ( .A1(n18673), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18359) );
  NOR2_X1 U21184 ( .A1(n18673), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18447) );
  NAND2_X1 U21185 ( .A1(n18524), .A2(n18447), .ZN(n18471) );
  AND2_X1 U21186 ( .A1(n18359), .A2(n18471), .ZN(n18181) );
  OAI22_X1 U21187 ( .A1(n18182), .A2(n18673), .B1(n18181), .B2(n18180), .ZN(
        P3_U2866) );
  NOR2_X1 U21188 ( .A1(n18674), .A2(n18183), .ZN(P3_U2867) );
  NOR2_X1 U21189 ( .A1(n18670), .A2(n18673), .ZN(n18497) );
  NAND2_X1 U21190 ( .A1(n18649), .A2(n18497), .ZN(n18495) );
  NOR2_X2 U21191 ( .A1(n18469), .A2(n18495), .ZN(n18603) );
  INV_X1 U21192 ( .A(n18603), .ZN(n18619) );
  NAND2_X1 U21193 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18566), .ZN(n18528) );
  NOR2_X2 U21194 ( .A1(n18288), .A2(n18184), .ZN(n18561) );
  NAND2_X1 U21195 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18653) );
  INV_X1 U21196 ( .A(n18497), .ZN(n18185) );
  NOR2_X2 U21197 ( .A1(n18653), .A2(n18185), .ZN(n18614) );
  NOR2_X1 U21198 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18652) );
  NOR2_X1 U21199 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18265) );
  NAND2_X1 U21200 ( .A1(n18652), .A2(n18265), .ZN(n18285) );
  NAND2_X1 U21201 ( .A1(n18263), .A2(n18285), .ZN(n18243) );
  AND2_X1 U21202 ( .A1(n18560), .A2(n18243), .ZN(n18217) );
  NAND2_X1 U21203 ( .A1(n18215), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18570) );
  INV_X1 U21204 ( .A(n18570), .ZN(n18521) );
  NOR2_X1 U21205 ( .A1(n18649), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18332) );
  NAND2_X1 U21206 ( .A1(n18497), .A2(n18332), .ZN(n18242) );
  INV_X1 U21207 ( .A(n18242), .ZN(n18556) );
  AOI22_X1 U21208 ( .A1(n18561), .A2(n18217), .B1(n18521), .B2(n18556), .ZN(
        n18190) );
  INV_X1 U21209 ( .A(n18332), .ZN(n18424) );
  NAND2_X1 U21210 ( .A1(n18649), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18403) );
  AND2_X1 U21211 ( .A1(n18424), .A2(n18403), .ZN(n18472) );
  NOR2_X1 U21212 ( .A1(n18472), .A2(n18185), .ZN(n18525) );
  AOI21_X1 U21213 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18288), .ZN(n18522) );
  AOI22_X1 U21214 ( .A1(n18566), .A2(n18525), .B1(n18522), .B2(n18243), .ZN(
        n18220) );
  INV_X1 U21215 ( .A(n18285), .ZN(n18278) );
  NAND2_X1 U21216 ( .A1(n18187), .A2(n18186), .ZN(n18218) );
  NOR2_X2 U21217 ( .A1(n18188), .A2(n18218), .ZN(n18567) );
  AOI22_X1 U21218 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18220), .B1(
        n18278), .B2(n18567), .ZN(n18189) );
  OAI211_X1 U21219 ( .C1(n18619), .C2(n18528), .A(n18190), .B(n18189), .ZN(
        P3_U2868) );
  NAND2_X1 U21220 ( .A1(n18215), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18532) );
  NAND2_X1 U21221 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18566), .ZN(n18576) );
  INV_X1 U21222 ( .A(n18576), .ZN(n18529) );
  NOR2_X2 U21223 ( .A1(n18288), .A2(n18191), .ZN(n18571) );
  AOI22_X1 U21224 ( .A1(n18603), .A2(n18529), .B1(n18217), .B2(n18571), .ZN(
        n18194) );
  NOR2_X2 U21225 ( .A1(n18192), .A2(n18218), .ZN(n18573) );
  AOI22_X1 U21226 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18220), .B1(
        n18278), .B2(n18573), .ZN(n18193) );
  OAI211_X1 U21227 ( .C1(n18242), .C2(n18532), .A(n18194), .B(n18193), .ZN(
        P3_U2869) );
  NAND2_X1 U21228 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18566), .ZN(n18536) );
  NOR2_X2 U21229 ( .A1(n18288), .A2(n18195), .ZN(n18577) );
  NAND2_X1 U21230 ( .A1(n18215), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18582) );
  INV_X1 U21231 ( .A(n18582), .ZN(n18533) );
  AOI22_X1 U21232 ( .A1(n18217), .A2(n18577), .B1(n18556), .B2(n18533), .ZN(
        n18198) );
  NOR2_X2 U21233 ( .A1(n18196), .A2(n18218), .ZN(n18579) );
  AOI22_X1 U21234 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18220), .B1(
        n18278), .B2(n18579), .ZN(n18197) );
  OAI211_X1 U21235 ( .C1(n18619), .C2(n18536), .A(n18198), .B(n18197), .ZN(
        P3_U2870) );
  NAND2_X1 U21236 ( .A1(n18215), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18588) );
  NAND2_X1 U21237 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18566), .ZN(n18541) );
  INV_X1 U21238 ( .A(n18541), .ZN(n18583) );
  NOR2_X2 U21239 ( .A1(n18288), .A2(n18199), .ZN(n18584) );
  AOI22_X1 U21240 ( .A1(n18603), .A2(n18583), .B1(n18217), .B2(n18584), .ZN(
        n18202) );
  NOR2_X2 U21241 ( .A1(n18200), .A2(n18218), .ZN(n18585) );
  AOI22_X1 U21242 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18220), .B1(
        n18278), .B2(n18585), .ZN(n18201) );
  OAI211_X1 U21243 ( .C1(n18242), .C2(n18588), .A(n18202), .B(n18201), .ZN(
        P3_U2871) );
  NAND2_X1 U21244 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n18566), .ZN(n18594) );
  NOR2_X2 U21245 ( .A1(n18288), .A2(n18203), .ZN(n18589) );
  NAND2_X1 U21246 ( .A1(n18215), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18545) );
  INV_X1 U21247 ( .A(n18545), .ZN(n18590) );
  AOI22_X1 U21248 ( .A1(n18217), .A2(n18589), .B1(n18556), .B2(n18590), .ZN(
        n18206) );
  NOR2_X2 U21249 ( .A1(n18204), .A2(n18218), .ZN(n18591) );
  AOI22_X1 U21250 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18220), .B1(
        n18278), .B2(n18591), .ZN(n18205) );
  OAI211_X1 U21251 ( .C1(n18619), .C2(n18594), .A(n18206), .B(n18205), .ZN(
        P3_U2872) );
  NAND2_X1 U21252 ( .A1(n18566), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18549) );
  NAND2_X1 U21253 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18566), .ZN(n18600) );
  INV_X1 U21254 ( .A(n18600), .ZN(n18546) );
  NOR2_X2 U21255 ( .A1(n18288), .A2(n18207), .ZN(n18595) );
  AOI22_X1 U21256 ( .A1(n18603), .A2(n18546), .B1(n18217), .B2(n18595), .ZN(
        n18210) );
  NOR2_X2 U21257 ( .A1(n18208), .A2(n18218), .ZN(n18597) );
  AOI22_X1 U21258 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18220), .B1(
        n18278), .B2(n18597), .ZN(n18209) );
  OAI211_X1 U21259 ( .C1(n18242), .C2(n18549), .A(n18210), .B(n18209), .ZN(
        P3_U2873) );
  NAND2_X1 U21260 ( .A1(n18566), .A2(BUF2_REG_22__SCAN_IN), .ZN(n18553) );
  NAND2_X1 U21261 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18566), .ZN(n18608) );
  NOR2_X2 U21262 ( .A1(n18288), .A2(n18211), .ZN(n18601) );
  AOI22_X1 U21263 ( .A1(n18603), .A2(n18550), .B1(n18217), .B2(n18601), .ZN(
        n18214) );
  NOR2_X2 U21264 ( .A1(n18212), .A2(n18218), .ZN(n18604) );
  AOI22_X1 U21265 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18220), .B1(
        n18278), .B2(n18604), .ZN(n18213) );
  OAI211_X1 U21266 ( .C1(n18242), .C2(n18553), .A(n18214), .B(n18213), .ZN(
        P3_U2874) );
  NAND2_X1 U21267 ( .A1(n18215), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18520) );
  NOR2_X2 U21268 ( .A1(n18216), .A2(n18288), .ZN(n18610) );
  NAND2_X1 U21269 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18566), .ZN(n18618) );
  INV_X1 U21270 ( .A(n18618), .ZN(n18515) );
  AOI22_X1 U21271 ( .A1(n18217), .A2(n18610), .B1(n18556), .B2(n18515), .ZN(
        n18222) );
  NOR2_X2 U21272 ( .A1(n18219), .A2(n18218), .ZN(n18613) );
  AOI22_X1 U21273 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18220), .B1(
        n18278), .B2(n18613), .ZN(n18221) );
  OAI211_X1 U21274 ( .C1(n18619), .C2(n18520), .A(n18222), .B(n18221), .ZN(
        P3_U2875) );
  INV_X1 U21275 ( .A(n18560), .ZN(n18694) );
  INV_X1 U21276 ( .A(n18265), .ZN(n18310) );
  AOI22_X1 U21277 ( .A1(n18614), .A2(n18521), .B1(n18561), .B2(n18238), .ZN(
        n18225) );
  NOR2_X1 U21278 ( .A1(n18673), .A2(n18401), .ZN(n18563) );
  NOR2_X1 U21279 ( .A1(n18288), .A2(n18223), .ZN(n18564) );
  AND2_X1 U21280 ( .A1(n18649), .A2(n18564), .ZN(n18496) );
  AOI22_X1 U21281 ( .A1(n18566), .A2(n18563), .B1(n18265), .B2(n18496), .ZN(
        n18239) );
  NOR2_X2 U21282 ( .A1(n18310), .A2(n18403), .ZN(n18306) );
  AOI22_X1 U21283 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18239), .B1(
        n18567), .B2(n18306), .ZN(n18224) );
  OAI211_X1 U21284 ( .C1(n18528), .C2(n18242), .A(n18225), .B(n18224), .ZN(
        P3_U2876) );
  INV_X1 U21285 ( .A(n18532), .ZN(n18572) );
  AOI22_X1 U21286 ( .A1(n18614), .A2(n18572), .B1(n18571), .B2(n18238), .ZN(
        n18227) );
  AOI22_X1 U21287 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18239), .B1(
        n18573), .B2(n18306), .ZN(n18226) );
  OAI211_X1 U21288 ( .C1(n18242), .C2(n18576), .A(n18227), .B(n18226), .ZN(
        P3_U2877) );
  INV_X1 U21289 ( .A(n18536), .ZN(n18578) );
  AOI22_X1 U21290 ( .A1(n18556), .A2(n18578), .B1(n18577), .B2(n18238), .ZN(
        n18229) );
  AOI22_X1 U21291 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18239), .B1(
        n18579), .B2(n18306), .ZN(n18228) );
  OAI211_X1 U21292 ( .C1(n18263), .C2(n18582), .A(n18229), .B(n18228), .ZN(
        P3_U2878) );
  AOI22_X1 U21293 ( .A1(n18556), .A2(n18583), .B1(n18584), .B2(n18238), .ZN(
        n18231) );
  AOI22_X1 U21294 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18239), .B1(
        n18585), .B2(n18306), .ZN(n18230) );
  OAI211_X1 U21295 ( .C1(n18263), .C2(n18588), .A(n18231), .B(n18230), .ZN(
        P3_U2879) );
  INV_X1 U21296 ( .A(n18594), .ZN(n18542) );
  AOI22_X1 U21297 ( .A1(n18556), .A2(n18542), .B1(n18589), .B2(n18238), .ZN(
        n18233) );
  AOI22_X1 U21298 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18239), .B1(
        n18591), .B2(n18306), .ZN(n18232) );
  OAI211_X1 U21299 ( .C1(n18263), .C2(n18545), .A(n18233), .B(n18232), .ZN(
        P3_U2880) );
  AOI22_X1 U21300 ( .A1(n18556), .A2(n18546), .B1(n18595), .B2(n18238), .ZN(
        n18235) );
  AOI22_X1 U21301 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18239), .B1(
        n18597), .B2(n18306), .ZN(n18234) );
  OAI211_X1 U21302 ( .C1(n18263), .C2(n18549), .A(n18235), .B(n18234), .ZN(
        P3_U2881) );
  INV_X1 U21303 ( .A(n18553), .ZN(n18602) );
  AOI22_X1 U21304 ( .A1(n18614), .A2(n18602), .B1(n18601), .B2(n18238), .ZN(
        n18237) );
  AOI22_X1 U21305 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18239), .B1(
        n18604), .B2(n18306), .ZN(n18236) );
  OAI211_X1 U21306 ( .C1(n18242), .C2(n18608), .A(n18237), .B(n18236), .ZN(
        P3_U2882) );
  AOI22_X1 U21307 ( .A1(n18614), .A2(n18515), .B1(n18610), .B2(n18238), .ZN(
        n18241) );
  AOI22_X1 U21308 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18239), .B1(
        n18613), .B2(n18306), .ZN(n18240) );
  OAI211_X1 U21309 ( .C1(n18242), .C2(n18520), .A(n18241), .B(n18240), .ZN(
        P3_U2883) );
  NOR2_X2 U21310 ( .A1(n18310), .A2(n18424), .ZN(n18324) );
  NOR2_X1 U21311 ( .A1(n18306), .A2(n18324), .ZN(n18287) );
  INV_X1 U21312 ( .A(n18287), .ZN(n18244) );
  OAI221_X1 U21313 ( .B1(n18244), .B2(n18524), .C1(n18244), .C2(n18243), .A(
        n18522), .ZN(n18260) );
  NOR2_X1 U21314 ( .A1(n18694), .A2(n18287), .ZN(n18259) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18260), .B1(
        n18561), .B2(n18259), .ZN(n18246) );
  AOI22_X1 U21316 ( .A1(n18278), .A2(n18521), .B1(n18567), .B2(n18324), .ZN(
        n18245) );
  OAI211_X1 U21317 ( .C1(n18528), .C2(n18263), .A(n18246), .B(n18245), .ZN(
        P3_U2884) );
  AOI22_X1 U21318 ( .A1(n18614), .A2(n18529), .B1(n18571), .B2(n18259), .ZN(
        n18248) );
  AOI22_X1 U21319 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18260), .B1(
        n18573), .B2(n18324), .ZN(n18247) );
  OAI211_X1 U21320 ( .C1(n18285), .C2(n18532), .A(n18248), .B(n18247), .ZN(
        P3_U2885) );
  AOI22_X1 U21321 ( .A1(n18278), .A2(n18533), .B1(n18577), .B2(n18259), .ZN(
        n18250) );
  AOI22_X1 U21322 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18260), .B1(
        n18579), .B2(n18324), .ZN(n18249) );
  OAI211_X1 U21323 ( .C1(n18263), .C2(n18536), .A(n18250), .B(n18249), .ZN(
        P3_U2886) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18260), .B1(
        n18584), .B2(n18259), .ZN(n18252) );
  AOI22_X1 U21325 ( .A1(n18614), .A2(n18583), .B1(n18585), .B2(n18324), .ZN(
        n18251) );
  OAI211_X1 U21326 ( .C1(n18285), .C2(n18588), .A(n18252), .B(n18251), .ZN(
        P3_U2887) );
  AOI22_X1 U21327 ( .A1(n18278), .A2(n18590), .B1(n18589), .B2(n18259), .ZN(
        n18254) );
  AOI22_X1 U21328 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18260), .B1(
        n18591), .B2(n18324), .ZN(n18253) );
  OAI211_X1 U21329 ( .C1(n18263), .C2(n18594), .A(n18254), .B(n18253), .ZN(
        P3_U2888) );
  INV_X1 U21330 ( .A(n18549), .ZN(n18596) );
  AOI22_X1 U21331 ( .A1(n18278), .A2(n18596), .B1(n18595), .B2(n18259), .ZN(
        n18256) );
  AOI22_X1 U21332 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18260), .B1(
        n18597), .B2(n18324), .ZN(n18255) );
  OAI211_X1 U21333 ( .C1(n18263), .C2(n18600), .A(n18256), .B(n18255), .ZN(
        P3_U2889) );
  AOI22_X1 U21334 ( .A1(n18278), .A2(n18602), .B1(n18601), .B2(n18259), .ZN(
        n18258) );
  AOI22_X1 U21335 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18260), .B1(
        n18604), .B2(n18324), .ZN(n18257) );
  OAI211_X1 U21336 ( .C1(n18263), .C2(n18608), .A(n18258), .B(n18257), .ZN(
        P3_U2890) );
  AOI22_X1 U21337 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18260), .B1(
        n18610), .B2(n18259), .ZN(n18262) );
  AOI22_X1 U21338 ( .A1(n18278), .A2(n18515), .B1(n18613), .B2(n18324), .ZN(
        n18261) );
  OAI211_X1 U21339 ( .C1(n18263), .C2(n18520), .A(n18262), .B(n18261), .ZN(
        P3_U2891) );
  INV_X1 U21340 ( .A(n18306), .ZN(n18300) );
  INV_X1 U21341 ( .A(n18528), .ZN(n18562) );
  AOI22_X1 U21342 ( .A1(n18562), .A2(n18278), .B1(n18561), .B2(n18281), .ZN(
        n18267) );
  NOR2_X1 U21343 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18524), .ZN(
        n18264) );
  AOI211_X1 U21344 ( .C1(P3_STATE2_REG_3__SCAN_IN), .C2(n18653), .A(n18264), 
        .B(n18288), .ZN(n18358) );
  NAND2_X1 U21345 ( .A1(n18265), .A2(n18358), .ZN(n18282) );
  NOR2_X2 U21346 ( .A1(n18653), .A2(n18310), .ZN(n18353) );
  AOI22_X1 U21347 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18282), .B1(
        n18567), .B2(n18353), .ZN(n18266) );
  OAI211_X1 U21348 ( .C1(n18570), .C2(n18300), .A(n18267), .B(n18266), .ZN(
        P3_U2892) );
  AOI22_X1 U21349 ( .A1(n18572), .A2(n18306), .B1(n18571), .B2(n18281), .ZN(
        n18269) );
  AOI22_X1 U21350 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18282), .B1(
        n18573), .B2(n18353), .ZN(n18268) );
  OAI211_X1 U21351 ( .C1(n18285), .C2(n18576), .A(n18269), .B(n18268), .ZN(
        P3_U2893) );
  AOI22_X1 U21352 ( .A1(n18577), .A2(n18281), .B1(n18533), .B2(n18306), .ZN(
        n18271) );
  AOI22_X1 U21353 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18282), .B1(
        n18579), .B2(n18353), .ZN(n18270) );
  OAI211_X1 U21354 ( .C1(n18285), .C2(n18536), .A(n18271), .B(n18270), .ZN(
        P3_U2894) );
  INV_X1 U21355 ( .A(n18588), .ZN(n18537) );
  AOI22_X1 U21356 ( .A1(n18537), .A2(n18306), .B1(n18584), .B2(n18281), .ZN(
        n18273) );
  AOI22_X1 U21357 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18282), .B1(
        n18585), .B2(n18353), .ZN(n18272) );
  OAI211_X1 U21358 ( .C1(n18285), .C2(n18541), .A(n18273), .B(n18272), .ZN(
        P3_U2895) );
  AOI22_X1 U21359 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18282), .B1(
        n18589), .B2(n18281), .ZN(n18275) );
  AOI22_X1 U21360 ( .A1(n18591), .A2(n18353), .B1(n18590), .B2(n18306), .ZN(
        n18274) );
  OAI211_X1 U21361 ( .C1(n18285), .C2(n18594), .A(n18275), .B(n18274), .ZN(
        P3_U2896) );
  AOI22_X1 U21362 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18282), .B1(
        n18595), .B2(n18281), .ZN(n18277) );
  AOI22_X1 U21363 ( .A1(n18278), .A2(n18546), .B1(n18597), .B2(n18353), .ZN(
        n18276) );
  OAI211_X1 U21364 ( .C1(n18549), .C2(n18300), .A(n18277), .B(n18276), .ZN(
        P3_U2897) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18282), .B1(
        n18601), .B2(n18281), .ZN(n18280) );
  AOI22_X1 U21366 ( .A1(n18278), .A2(n18550), .B1(n18604), .B2(n18353), .ZN(
        n18279) );
  OAI211_X1 U21367 ( .C1(n18553), .C2(n18300), .A(n18280), .B(n18279), .ZN(
        P3_U2898) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18282), .B1(
        n18610), .B2(n18281), .ZN(n18284) );
  AOI22_X1 U21369 ( .A1(n18613), .A2(n18353), .B1(n18515), .B2(n18306), .ZN(
        n18283) );
  OAI211_X1 U21370 ( .C1(n18285), .C2(n18520), .A(n18284), .B(n18283), .ZN(
        P3_U2899) );
  INV_X1 U21371 ( .A(n18652), .ZN(n18286) );
  NOR2_X2 U21372 ( .A1(n18286), .A2(n18359), .ZN(n18376) );
  INV_X1 U21373 ( .A(n18376), .ZN(n18372) );
  AOI21_X1 U21374 ( .B1(n18351), .B2(n18372), .A(n18694), .ZN(n18305) );
  AOI22_X1 U21375 ( .A1(n18561), .A2(n18305), .B1(n18521), .B2(n18324), .ZN(
        n18291) );
  AOI221_X1 U21376 ( .B1(n18287), .B2(n18351), .C1(n18334), .C2(n18351), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18289) );
  INV_X1 U21377 ( .A(n18288), .ZN(n18474) );
  OAI21_X1 U21378 ( .B1(n18376), .B2(n18289), .A(n18474), .ZN(n18307) );
  AOI22_X1 U21379 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18307), .B1(
        n18567), .B2(n18376), .ZN(n18290) );
  OAI211_X1 U21380 ( .C1(n18528), .C2(n18300), .A(n18291), .B(n18290), .ZN(
        P3_U2900) );
  AOI22_X1 U21381 ( .A1(n18572), .A2(n18324), .B1(n18571), .B2(n18305), .ZN(
        n18293) );
  AOI22_X1 U21382 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18307), .B1(
        n18573), .B2(n18376), .ZN(n18292) );
  OAI211_X1 U21383 ( .C1(n18576), .C2(n18300), .A(n18293), .B(n18292), .ZN(
        P3_U2901) );
  AOI22_X1 U21384 ( .A1(n18577), .A2(n18305), .B1(n18533), .B2(n18324), .ZN(
        n18295) );
  AOI22_X1 U21385 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18307), .B1(
        n18579), .B2(n18376), .ZN(n18294) );
  OAI211_X1 U21386 ( .C1(n18536), .C2(n18300), .A(n18295), .B(n18294), .ZN(
        P3_U2902) );
  AOI22_X1 U21387 ( .A1(n18537), .A2(n18324), .B1(n18584), .B2(n18305), .ZN(
        n18297) );
  AOI22_X1 U21388 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18307), .B1(
        n18585), .B2(n18376), .ZN(n18296) );
  OAI211_X1 U21389 ( .C1(n18541), .C2(n18300), .A(n18297), .B(n18296), .ZN(
        P3_U2903) );
  AOI22_X1 U21390 ( .A1(n18590), .A2(n18324), .B1(n18589), .B2(n18305), .ZN(
        n18299) );
  AOI22_X1 U21391 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18307), .B1(
        n18591), .B2(n18376), .ZN(n18298) );
  OAI211_X1 U21392 ( .C1(n18594), .C2(n18300), .A(n18299), .B(n18298), .ZN(
        P3_U2904) );
  INV_X1 U21393 ( .A(n18324), .ZN(n18331) );
  AOI22_X1 U21394 ( .A1(n18546), .A2(n18306), .B1(n18595), .B2(n18305), .ZN(
        n18302) );
  AOI22_X1 U21395 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18307), .B1(
        n18597), .B2(n18376), .ZN(n18301) );
  OAI211_X1 U21396 ( .C1(n18549), .C2(n18331), .A(n18302), .B(n18301), .ZN(
        P3_U2905) );
  AOI22_X1 U21397 ( .A1(n18550), .A2(n18306), .B1(n18601), .B2(n18305), .ZN(
        n18304) );
  AOI22_X1 U21398 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18307), .B1(
        n18604), .B2(n18376), .ZN(n18303) );
  OAI211_X1 U21399 ( .C1(n18553), .C2(n18331), .A(n18304), .B(n18303), .ZN(
        P3_U2906) );
  INV_X1 U21400 ( .A(n18520), .ZN(n18612) );
  AOI22_X1 U21401 ( .A1(n18612), .A2(n18306), .B1(n18610), .B2(n18305), .ZN(
        n18309) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18307), .B1(
        n18613), .B2(n18376), .ZN(n18308) );
  OAI211_X1 U21403 ( .C1(n18618), .C2(n18331), .A(n18309), .B(n18308), .ZN(
        P3_U2907) );
  AOI22_X1 U21404 ( .A1(n18561), .A2(n18327), .B1(n18521), .B2(n18353), .ZN(
        n18313) );
  NOR2_X1 U21405 ( .A1(n18649), .A2(n18310), .ZN(n18311) );
  INV_X1 U21406 ( .A(n18359), .ZN(n18357) );
  AOI22_X1 U21407 ( .A1(n18566), .A2(n18311), .B1(n18496), .B2(n18357), .ZN(
        n18328) );
  NOR2_X2 U21408 ( .A1(n18403), .A2(n18359), .ZN(n18398) );
  AOI22_X1 U21409 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18328), .B1(
        n18567), .B2(n18398), .ZN(n18312) );
  OAI211_X1 U21410 ( .C1(n18528), .C2(n18331), .A(n18313), .B(n18312), .ZN(
        P3_U2908) );
  AOI22_X1 U21411 ( .A1(n18529), .A2(n18324), .B1(n18571), .B2(n18327), .ZN(
        n18315) );
  AOI22_X1 U21412 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18328), .B1(
        n18573), .B2(n18398), .ZN(n18314) );
  OAI211_X1 U21413 ( .C1(n18532), .C2(n18351), .A(n18315), .B(n18314), .ZN(
        P3_U2909) );
  AOI22_X1 U21414 ( .A1(n18577), .A2(n18327), .B1(n18533), .B2(n18353), .ZN(
        n18317) );
  AOI22_X1 U21415 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18328), .B1(
        n18579), .B2(n18398), .ZN(n18316) );
  OAI211_X1 U21416 ( .C1(n18536), .C2(n18331), .A(n18317), .B(n18316), .ZN(
        P3_U2910) );
  AOI22_X1 U21417 ( .A1(n18537), .A2(n18353), .B1(n18584), .B2(n18327), .ZN(
        n18319) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18328), .B1(
        n18585), .B2(n18398), .ZN(n18318) );
  OAI211_X1 U21419 ( .C1(n18541), .C2(n18331), .A(n18319), .B(n18318), .ZN(
        P3_U2911) );
  AOI22_X1 U21420 ( .A1(n18542), .A2(n18324), .B1(n18589), .B2(n18327), .ZN(
        n18321) );
  AOI22_X1 U21421 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18328), .B1(
        n18591), .B2(n18398), .ZN(n18320) );
  OAI211_X1 U21422 ( .C1(n18545), .C2(n18351), .A(n18321), .B(n18320), .ZN(
        P3_U2912) );
  AOI22_X1 U21423 ( .A1(n18546), .A2(n18324), .B1(n18595), .B2(n18327), .ZN(
        n18323) );
  AOI22_X1 U21424 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18328), .B1(
        n18597), .B2(n18398), .ZN(n18322) );
  OAI211_X1 U21425 ( .C1(n18549), .C2(n18351), .A(n18323), .B(n18322), .ZN(
        P3_U2913) );
  AOI22_X1 U21426 ( .A1(n18550), .A2(n18324), .B1(n18601), .B2(n18327), .ZN(
        n18326) );
  AOI22_X1 U21427 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18328), .B1(
        n18604), .B2(n18398), .ZN(n18325) );
  OAI211_X1 U21428 ( .C1(n18553), .C2(n18351), .A(n18326), .B(n18325), .ZN(
        P3_U2914) );
  AOI22_X1 U21429 ( .A1(n18515), .A2(n18353), .B1(n18610), .B2(n18327), .ZN(
        n18330) );
  AOI22_X1 U21430 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18328), .B1(
        n18613), .B2(n18398), .ZN(n18329) );
  OAI211_X1 U21431 ( .C1(n18520), .C2(n18331), .A(n18330), .B(n18329), .ZN(
        P3_U2915) );
  NAND2_X1 U21432 ( .A1(n18332), .A2(n18357), .ZN(n18418) );
  NAND2_X1 U21433 ( .A1(n18393), .A2(n18418), .ZN(n18380) );
  INV_X1 U21434 ( .A(n18380), .ZN(n18333) );
  NOR2_X1 U21435 ( .A1(n18694), .A2(n18333), .ZN(n18352) );
  AOI22_X1 U21436 ( .A1(n18561), .A2(n18352), .B1(n18521), .B2(n18376), .ZN(
        n18338) );
  NOR2_X1 U21437 ( .A1(n18353), .A2(n18376), .ZN(n18335) );
  OAI21_X1 U21438 ( .B1(n18335), .B2(n18334), .A(n18333), .ZN(n18336) );
  OAI211_X1 U21439 ( .C1(n18420), .C2(n18790), .A(n18474), .B(n18336), .ZN(
        n18354) );
  AOI22_X1 U21440 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18354), .B1(
        n18567), .B2(n18420), .ZN(n18337) );
  OAI211_X1 U21441 ( .C1(n18528), .C2(n18351), .A(n18338), .B(n18337), .ZN(
        P3_U2916) );
  AOI22_X1 U21442 ( .A1(n18572), .A2(n18376), .B1(n18571), .B2(n18352), .ZN(
        n18340) );
  AOI22_X1 U21443 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18354), .B1(
        n18573), .B2(n18420), .ZN(n18339) );
  OAI211_X1 U21444 ( .C1(n18576), .C2(n18351), .A(n18340), .B(n18339), .ZN(
        P3_U2917) );
  AOI22_X1 U21445 ( .A1(n18578), .A2(n18353), .B1(n18577), .B2(n18352), .ZN(
        n18342) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18354), .B1(
        n18579), .B2(n18420), .ZN(n18341) );
  OAI211_X1 U21447 ( .C1(n18582), .C2(n18372), .A(n18342), .B(n18341), .ZN(
        P3_U2918) );
  AOI22_X1 U21448 ( .A1(n18537), .A2(n18376), .B1(n18584), .B2(n18352), .ZN(
        n18344) );
  AOI22_X1 U21449 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18354), .B1(
        n18585), .B2(n18420), .ZN(n18343) );
  OAI211_X1 U21450 ( .C1(n18541), .C2(n18351), .A(n18344), .B(n18343), .ZN(
        P3_U2919) );
  AOI22_X1 U21451 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18354), .B1(
        n18589), .B2(n18352), .ZN(n18346) );
  AOI22_X1 U21452 ( .A1(n18542), .A2(n18353), .B1(n18591), .B2(n18420), .ZN(
        n18345) );
  OAI211_X1 U21453 ( .C1(n18545), .C2(n18372), .A(n18346), .B(n18345), .ZN(
        P3_U2920) );
  AOI22_X1 U21454 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18354), .B1(
        n18595), .B2(n18352), .ZN(n18348) );
  AOI22_X1 U21455 ( .A1(n18596), .A2(n18376), .B1(n18597), .B2(n18420), .ZN(
        n18347) );
  OAI211_X1 U21456 ( .C1(n18600), .C2(n18351), .A(n18348), .B(n18347), .ZN(
        P3_U2921) );
  AOI22_X1 U21457 ( .A1(n18602), .A2(n18376), .B1(n18601), .B2(n18352), .ZN(
        n18350) );
  AOI22_X1 U21458 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18354), .B1(
        n18604), .B2(n18420), .ZN(n18349) );
  OAI211_X1 U21459 ( .C1(n18608), .C2(n18351), .A(n18350), .B(n18349), .ZN(
        P3_U2922) );
  AOI22_X1 U21460 ( .A1(n18612), .A2(n18353), .B1(n18610), .B2(n18352), .ZN(
        n18356) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18354), .B1(
        n18613), .B2(n18420), .ZN(n18355) );
  OAI211_X1 U21462 ( .C1(n18618), .C2(n18372), .A(n18356), .B(n18355), .ZN(
        P3_U2923) );
  AOI22_X1 U21463 ( .A1(n18562), .A2(n18376), .B1(n18561), .B2(n18375), .ZN(
        n18361) );
  NAND2_X1 U21464 ( .A1(n18358), .A2(n18357), .ZN(n18377) );
  NOR2_X2 U21465 ( .A1(n18653), .A2(n18359), .ZN(n18435) );
  AOI22_X1 U21466 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18377), .B1(
        n18567), .B2(n18435), .ZN(n18360) );
  OAI211_X1 U21467 ( .C1(n18570), .C2(n18393), .A(n18361), .B(n18360), .ZN(
        P3_U2924) );
  AOI22_X1 U21468 ( .A1(n18529), .A2(n18376), .B1(n18571), .B2(n18375), .ZN(
        n18363) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18377), .B1(
        n18573), .B2(n18435), .ZN(n18362) );
  OAI211_X1 U21470 ( .C1(n18532), .C2(n18393), .A(n18363), .B(n18362), .ZN(
        P3_U2925) );
  AOI22_X1 U21471 ( .A1(n18577), .A2(n18375), .B1(n18533), .B2(n18398), .ZN(
        n18365) );
  AOI22_X1 U21472 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18377), .B1(
        n18579), .B2(n18435), .ZN(n18364) );
  OAI211_X1 U21473 ( .C1(n18536), .C2(n18372), .A(n18365), .B(n18364), .ZN(
        P3_U2926) );
  AOI22_X1 U21474 ( .A1(n18584), .A2(n18375), .B1(n18583), .B2(n18376), .ZN(
        n18367) );
  AOI22_X1 U21475 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18377), .B1(
        n18585), .B2(n18435), .ZN(n18366) );
  OAI211_X1 U21476 ( .C1(n18588), .C2(n18393), .A(n18367), .B(n18366), .ZN(
        P3_U2927) );
  AOI22_X1 U21477 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18377), .B1(
        n18589), .B2(n18375), .ZN(n18369) );
  AOI22_X1 U21478 ( .A1(n18591), .A2(n18435), .B1(n18590), .B2(n18398), .ZN(
        n18368) );
  OAI211_X1 U21479 ( .C1(n18594), .C2(n18372), .A(n18369), .B(n18368), .ZN(
        P3_U2928) );
  AOI22_X1 U21480 ( .A1(n18596), .A2(n18398), .B1(n18595), .B2(n18375), .ZN(
        n18371) );
  AOI22_X1 U21481 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18377), .B1(
        n18597), .B2(n18435), .ZN(n18370) );
  OAI211_X1 U21482 ( .C1(n18600), .C2(n18372), .A(n18371), .B(n18370), .ZN(
        P3_U2929) );
  AOI22_X1 U21483 ( .A1(n18550), .A2(n18376), .B1(n18601), .B2(n18375), .ZN(
        n18374) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18377), .B1(
        n18604), .B2(n18435), .ZN(n18373) );
  OAI211_X1 U21485 ( .C1(n18553), .C2(n18393), .A(n18374), .B(n18373), .ZN(
        P3_U2930) );
  AOI22_X1 U21486 ( .A1(n18612), .A2(n18376), .B1(n18610), .B2(n18375), .ZN(
        n18379) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18377), .B1(
        n18613), .B2(n18435), .ZN(n18378) );
  OAI211_X1 U21488 ( .C1(n18618), .C2(n18393), .A(n18379), .B(n18378), .ZN(
        P3_U2931) );
  NAND2_X1 U21489 ( .A1(n18652), .A2(n18447), .ZN(n18461) );
  NAND2_X1 U21490 ( .A1(n18446), .A2(n18461), .ZN(n18425) );
  AND2_X1 U21491 ( .A1(n18560), .A2(n18425), .ZN(n18396) );
  AOI22_X1 U21492 ( .A1(n18561), .A2(n18396), .B1(n18521), .B2(n18420), .ZN(
        n18382) );
  OAI221_X1 U21493 ( .B1(n18425), .B2(n18524), .C1(n18425), .C2(n18380), .A(
        n18522), .ZN(n18397) );
  INV_X1 U21494 ( .A(n18461), .ZN(n18465) );
  AOI22_X1 U21495 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18397), .B1(
        n18567), .B2(n18465), .ZN(n18381) );
  OAI211_X1 U21496 ( .C1(n18528), .C2(n18393), .A(n18382), .B(n18381), .ZN(
        P3_U2932) );
  AOI22_X1 U21497 ( .A1(n18572), .A2(n18420), .B1(n18571), .B2(n18396), .ZN(
        n18384) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18397), .B1(
        n18573), .B2(n18465), .ZN(n18383) );
  OAI211_X1 U21499 ( .C1(n18576), .C2(n18393), .A(n18384), .B(n18383), .ZN(
        P3_U2933) );
  AOI22_X1 U21500 ( .A1(n18578), .A2(n18398), .B1(n18577), .B2(n18396), .ZN(
        n18386) );
  AOI22_X1 U21501 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18397), .B1(
        n18579), .B2(n18465), .ZN(n18385) );
  OAI211_X1 U21502 ( .C1(n18582), .C2(n18418), .A(n18386), .B(n18385), .ZN(
        P3_U2934) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18397), .B1(
        n18584), .B2(n18396), .ZN(n18388) );
  AOI22_X1 U21504 ( .A1(n18537), .A2(n18420), .B1(n18585), .B2(n18465), .ZN(
        n18387) );
  OAI211_X1 U21505 ( .C1(n18541), .C2(n18393), .A(n18388), .B(n18387), .ZN(
        P3_U2935) );
  AOI22_X1 U21506 ( .A1(n18542), .A2(n18398), .B1(n18589), .B2(n18396), .ZN(
        n18390) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18397), .B1(
        n18591), .B2(n18465), .ZN(n18389) );
  OAI211_X1 U21508 ( .C1(n18545), .C2(n18418), .A(n18390), .B(n18389), .ZN(
        P3_U2936) );
  AOI22_X1 U21509 ( .A1(n18596), .A2(n18420), .B1(n18595), .B2(n18396), .ZN(
        n18392) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18397), .B1(
        n18597), .B2(n18465), .ZN(n18391) );
  OAI211_X1 U21511 ( .C1(n18600), .C2(n18393), .A(n18392), .B(n18391), .ZN(
        P3_U2937) );
  AOI22_X1 U21512 ( .A1(n18550), .A2(n18398), .B1(n18601), .B2(n18396), .ZN(
        n18395) );
  AOI22_X1 U21513 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18397), .B1(
        n18604), .B2(n18465), .ZN(n18394) );
  OAI211_X1 U21514 ( .C1(n18553), .C2(n18418), .A(n18395), .B(n18394), .ZN(
        P3_U2938) );
  AOI22_X1 U21515 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18397), .B1(
        n18610), .B2(n18396), .ZN(n18400) );
  AOI22_X1 U21516 ( .A1(n18612), .A2(n18398), .B1(n18613), .B2(n18465), .ZN(
        n18399) );
  OAI211_X1 U21517 ( .C1(n18618), .C2(n18418), .A(n18400), .B(n18399), .ZN(
        P3_U2939) );
  INV_X1 U21518 ( .A(n18447), .ZN(n18448) );
  AOI22_X1 U21519 ( .A1(n18562), .A2(n18420), .B1(n18561), .B2(n18419), .ZN(
        n18405) );
  NOR2_X1 U21520 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18401), .ZN(
        n18402) );
  AOI22_X1 U21521 ( .A1(n18566), .A2(n18402), .B1(n18496), .B2(n18447), .ZN(
        n18421) );
  NOR2_X2 U21522 ( .A1(n18403), .A2(n18448), .ZN(n18491) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18421), .B1(
        n18567), .B2(n18491), .ZN(n18404) );
  OAI211_X1 U21524 ( .C1(n18570), .C2(n18446), .A(n18405), .B(n18404), .ZN(
        P3_U2940) );
  AOI22_X1 U21525 ( .A1(n18529), .A2(n18420), .B1(n18571), .B2(n18419), .ZN(
        n18407) );
  AOI22_X1 U21526 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18421), .B1(
        n18573), .B2(n18491), .ZN(n18406) );
  OAI211_X1 U21527 ( .C1(n18532), .C2(n18446), .A(n18407), .B(n18406), .ZN(
        P3_U2941) );
  AOI22_X1 U21528 ( .A1(n18578), .A2(n18420), .B1(n18577), .B2(n18419), .ZN(
        n18409) );
  AOI22_X1 U21529 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18421), .B1(
        n18579), .B2(n18491), .ZN(n18408) );
  OAI211_X1 U21530 ( .C1(n18582), .C2(n18446), .A(n18409), .B(n18408), .ZN(
        P3_U2942) );
  AOI22_X1 U21531 ( .A1(n18537), .A2(n18435), .B1(n18584), .B2(n18419), .ZN(
        n18411) );
  AOI22_X1 U21532 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18421), .B1(
        n18585), .B2(n18491), .ZN(n18410) );
  OAI211_X1 U21533 ( .C1(n18541), .C2(n18418), .A(n18411), .B(n18410), .ZN(
        P3_U2943) );
  AOI22_X1 U21534 ( .A1(n18542), .A2(n18420), .B1(n18589), .B2(n18419), .ZN(
        n18413) );
  AOI22_X1 U21535 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18421), .B1(
        n18591), .B2(n18491), .ZN(n18412) );
  OAI211_X1 U21536 ( .C1(n18545), .C2(n18446), .A(n18413), .B(n18412), .ZN(
        P3_U2944) );
  AOI22_X1 U21537 ( .A1(n18546), .A2(n18420), .B1(n18595), .B2(n18419), .ZN(
        n18415) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18421), .B1(
        n18597), .B2(n18491), .ZN(n18414) );
  OAI211_X1 U21539 ( .C1(n18549), .C2(n18446), .A(n18415), .B(n18414), .ZN(
        P3_U2945) );
  AOI22_X1 U21540 ( .A1(n18602), .A2(n18435), .B1(n18601), .B2(n18419), .ZN(
        n18417) );
  AOI22_X1 U21541 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18421), .B1(
        n18604), .B2(n18491), .ZN(n18416) );
  OAI211_X1 U21542 ( .C1(n18608), .C2(n18418), .A(n18417), .B(n18416), .ZN(
        P3_U2946) );
  AOI22_X1 U21543 ( .A1(n18612), .A2(n18420), .B1(n18610), .B2(n18419), .ZN(
        n18423) );
  AOI22_X1 U21544 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18421), .B1(
        n18613), .B2(n18491), .ZN(n18422) );
  OAI211_X1 U21545 ( .C1(n18618), .C2(n18446), .A(n18423), .B(n18422), .ZN(
        P3_U2947) );
  INV_X1 U21546 ( .A(n18491), .ZN(n18481) );
  NOR2_X2 U21547 ( .A1(n18424), .A2(n18448), .ZN(n18511) );
  AOI21_X1 U21548 ( .B1(n18481), .B2(n18519), .A(n18694), .ZN(n18442) );
  AOI22_X1 U21549 ( .A1(n18562), .A2(n18435), .B1(n18561), .B2(n18442), .ZN(
        n18428) );
  NAND2_X1 U21550 ( .A1(n18481), .A2(n18519), .ZN(n18426) );
  OAI221_X1 U21551 ( .B1(n18426), .B2(n18524), .C1(n18426), .C2(n18425), .A(
        n18522), .ZN(n18443) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18443), .B1(
        n18567), .B2(n18511), .ZN(n18427) );
  OAI211_X1 U21553 ( .C1(n18570), .C2(n18461), .A(n18428), .B(n18427), .ZN(
        P3_U2948) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18443), .B1(
        n18571), .B2(n18442), .ZN(n18430) );
  AOI22_X1 U21555 ( .A1(n18572), .A2(n18465), .B1(n18573), .B2(n18511), .ZN(
        n18429) );
  OAI211_X1 U21556 ( .C1(n18576), .C2(n18446), .A(n18430), .B(n18429), .ZN(
        P3_U2949) );
  AOI22_X1 U21557 ( .A1(n18578), .A2(n18435), .B1(n18577), .B2(n18442), .ZN(
        n18432) );
  AOI22_X1 U21558 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18443), .B1(
        n18579), .B2(n18511), .ZN(n18431) );
  OAI211_X1 U21559 ( .C1(n18582), .C2(n18461), .A(n18432), .B(n18431), .ZN(
        P3_U2950) );
  AOI22_X1 U21560 ( .A1(n18584), .A2(n18442), .B1(n18583), .B2(n18435), .ZN(
        n18434) );
  AOI22_X1 U21561 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18443), .B1(
        n18585), .B2(n18511), .ZN(n18433) );
  OAI211_X1 U21562 ( .C1(n18588), .C2(n18461), .A(n18434), .B(n18433), .ZN(
        P3_U2951) );
  AOI22_X1 U21563 ( .A1(n18542), .A2(n18435), .B1(n18589), .B2(n18442), .ZN(
        n18437) );
  AOI22_X1 U21564 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18443), .B1(
        n18591), .B2(n18511), .ZN(n18436) );
  OAI211_X1 U21565 ( .C1(n18545), .C2(n18461), .A(n18437), .B(n18436), .ZN(
        P3_U2952) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18443), .B1(
        n18595), .B2(n18442), .ZN(n18439) );
  AOI22_X1 U21567 ( .A1(n18596), .A2(n18465), .B1(n18597), .B2(n18511), .ZN(
        n18438) );
  OAI211_X1 U21568 ( .C1(n18600), .C2(n18446), .A(n18439), .B(n18438), .ZN(
        P3_U2953) );
  AOI22_X1 U21569 ( .A1(n18602), .A2(n18465), .B1(n18601), .B2(n18442), .ZN(
        n18441) );
  AOI22_X1 U21570 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18443), .B1(
        n18604), .B2(n18511), .ZN(n18440) );
  OAI211_X1 U21571 ( .C1(n18608), .C2(n18446), .A(n18441), .B(n18440), .ZN(
        P3_U2954) );
  AOI22_X1 U21572 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18443), .B1(
        n18610), .B2(n18442), .ZN(n18445) );
  AOI22_X1 U21573 ( .A1(n18613), .A2(n18511), .B1(n18515), .B2(n18465), .ZN(
        n18444) );
  OAI211_X1 U21574 ( .C1(n18520), .C2(n18446), .A(n18445), .B(n18444), .ZN(
        P3_U2955) );
  NOR2_X1 U21575 ( .A1(n18649), .A2(n18448), .ZN(n18498) );
  AND2_X1 U21576 ( .A1(n18560), .A2(n18498), .ZN(n18464) );
  AOI22_X1 U21577 ( .A1(n18561), .A2(n18464), .B1(n18521), .B2(n18491), .ZN(
        n18450) );
  OAI211_X1 U21578 ( .C1(n18566), .C2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n18564), .B(n18447), .ZN(n18466) );
  NOR2_X2 U21579 ( .A1(n18653), .A2(n18448), .ZN(n18555) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18466), .B1(
        n18567), .B2(n18555), .ZN(n18449) );
  OAI211_X1 U21581 ( .C1(n18528), .C2(n18461), .A(n18450), .B(n18449), .ZN(
        P3_U2956) );
  AOI22_X1 U21582 ( .A1(n18529), .A2(n18465), .B1(n18571), .B2(n18464), .ZN(
        n18452) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18466), .B1(
        n18573), .B2(n18555), .ZN(n18451) );
  OAI211_X1 U21584 ( .C1(n18532), .C2(n18481), .A(n18452), .B(n18451), .ZN(
        P3_U2957) );
  AOI22_X1 U21585 ( .A1(n18578), .A2(n18465), .B1(n18577), .B2(n18464), .ZN(
        n18454) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18466), .B1(
        n18579), .B2(n18555), .ZN(n18453) );
  OAI211_X1 U21587 ( .C1(n18582), .C2(n18481), .A(n18454), .B(n18453), .ZN(
        P3_U2958) );
  AOI22_X1 U21588 ( .A1(n18537), .A2(n18491), .B1(n18584), .B2(n18464), .ZN(
        n18456) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18466), .B1(
        n18585), .B2(n18555), .ZN(n18455) );
  OAI211_X1 U21590 ( .C1(n18541), .C2(n18461), .A(n18456), .B(n18455), .ZN(
        P3_U2959) );
  AOI22_X1 U21591 ( .A1(n18542), .A2(n18465), .B1(n18589), .B2(n18464), .ZN(
        n18458) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18466), .B1(
        n18591), .B2(n18555), .ZN(n18457) );
  OAI211_X1 U21593 ( .C1(n18545), .C2(n18481), .A(n18458), .B(n18457), .ZN(
        P3_U2960) );
  AOI22_X1 U21594 ( .A1(n18596), .A2(n18491), .B1(n18595), .B2(n18464), .ZN(
        n18460) );
  AOI22_X1 U21595 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18466), .B1(
        n18597), .B2(n18555), .ZN(n18459) );
  OAI211_X1 U21596 ( .C1(n18600), .C2(n18461), .A(n18460), .B(n18459), .ZN(
        P3_U2961) );
  AOI22_X1 U21597 ( .A1(n18550), .A2(n18465), .B1(n18601), .B2(n18464), .ZN(
        n18463) );
  AOI22_X1 U21598 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18466), .B1(
        n18604), .B2(n18555), .ZN(n18462) );
  OAI211_X1 U21599 ( .C1(n18553), .C2(n18481), .A(n18463), .B(n18462), .ZN(
        P3_U2962) );
  AOI22_X1 U21600 ( .A1(n18612), .A2(n18465), .B1(n18610), .B2(n18464), .ZN(
        n18468) );
  AOI22_X1 U21601 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18466), .B1(
        n18613), .B2(n18555), .ZN(n18467) );
  OAI211_X1 U21602 ( .C1(n18618), .C2(n18481), .A(n18468), .B(n18467), .ZN(
        P3_U2963) );
  INV_X1 U21603 ( .A(n18555), .ZN(n18540) );
  INV_X1 U21604 ( .A(n18495), .ZN(n18565) );
  NAND2_X1 U21605 ( .A1(n18469), .A2(n18565), .ZN(n18607) );
  NAND2_X1 U21606 ( .A1(n18540), .A2(n18607), .ZN(n18523) );
  INV_X1 U21607 ( .A(n18523), .ZN(n18470) );
  NOR2_X1 U21608 ( .A1(n18694), .A2(n18470), .ZN(n18490) );
  AOI22_X1 U21609 ( .A1(n18562), .A2(n18491), .B1(n18561), .B2(n18490), .ZN(
        n18476) );
  INV_X1 U21610 ( .A(n18607), .ZN(n18611) );
  OAI21_X1 U21611 ( .B1(n18472), .B2(n18471), .A(n18470), .ZN(n18473) );
  OAI211_X1 U21612 ( .C1(n18611), .C2(n18790), .A(n18474), .B(n18473), .ZN(
        n18492) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18492), .B1(
        n18567), .B2(n18611), .ZN(n18475) );
  OAI211_X1 U21614 ( .C1(n18570), .C2(n18519), .A(n18476), .B(n18475), .ZN(
        P3_U2964) );
  AOI22_X1 U21615 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18492), .B1(
        n18571), .B2(n18490), .ZN(n18478) );
  AOI22_X1 U21616 ( .A1(n18572), .A2(n18511), .B1(n18573), .B2(n18611), .ZN(
        n18477) );
  OAI211_X1 U21617 ( .C1(n18576), .C2(n18481), .A(n18478), .B(n18477), .ZN(
        P3_U2965) );
  AOI22_X1 U21618 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18492), .B1(
        n18577), .B2(n18490), .ZN(n18480) );
  AOI22_X1 U21619 ( .A1(n18579), .A2(n18611), .B1(n18533), .B2(n18511), .ZN(
        n18479) );
  OAI211_X1 U21620 ( .C1(n18536), .C2(n18481), .A(n18480), .B(n18479), .ZN(
        P3_U2966) );
  AOI22_X1 U21621 ( .A1(n18584), .A2(n18490), .B1(n18583), .B2(n18491), .ZN(
        n18483) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18492), .B1(
        n18585), .B2(n18611), .ZN(n18482) );
  OAI211_X1 U21623 ( .C1(n18588), .C2(n18519), .A(n18483), .B(n18482), .ZN(
        P3_U2967) );
  AOI22_X1 U21624 ( .A1(n18542), .A2(n18491), .B1(n18589), .B2(n18490), .ZN(
        n18485) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18492), .B1(
        n18591), .B2(n18611), .ZN(n18484) );
  OAI211_X1 U21626 ( .C1(n18545), .C2(n18519), .A(n18485), .B(n18484), .ZN(
        P3_U2968) );
  AOI22_X1 U21627 ( .A1(n18546), .A2(n18491), .B1(n18595), .B2(n18490), .ZN(
        n18487) );
  AOI22_X1 U21628 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18492), .B1(
        n18597), .B2(n18611), .ZN(n18486) );
  OAI211_X1 U21629 ( .C1(n18549), .C2(n18519), .A(n18487), .B(n18486), .ZN(
        P3_U2969) );
  AOI22_X1 U21630 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18492), .B1(
        n18601), .B2(n18490), .ZN(n18489) );
  AOI22_X1 U21631 ( .A1(n18604), .A2(n18611), .B1(n18550), .B2(n18491), .ZN(
        n18488) );
  OAI211_X1 U21632 ( .C1(n18553), .C2(n18519), .A(n18489), .B(n18488), .ZN(
        P3_U2970) );
  AOI22_X1 U21633 ( .A1(n18612), .A2(n18491), .B1(n18610), .B2(n18490), .ZN(
        n18494) );
  AOI22_X1 U21634 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18492), .B1(
        n18613), .B2(n18611), .ZN(n18493) );
  OAI211_X1 U21635 ( .C1(n18618), .C2(n18519), .A(n18494), .B(n18493), .ZN(
        P3_U2971) );
  NOR2_X1 U21636 ( .A1(n18694), .A2(n18495), .ZN(n18514) );
  AOI22_X1 U21637 ( .A1(n18562), .A2(n18511), .B1(n18561), .B2(n18514), .ZN(
        n18500) );
  AOI22_X1 U21638 ( .A1(n18566), .A2(n18498), .B1(n18497), .B2(n18496), .ZN(
        n18516) );
  AOI22_X1 U21639 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18516), .B1(
        n18603), .B2(n18567), .ZN(n18499) );
  OAI211_X1 U21640 ( .C1(n18570), .C2(n18540), .A(n18500), .B(n18499), .ZN(
        P3_U2972) );
  AOI22_X1 U21641 ( .A1(n18572), .A2(n18555), .B1(n18571), .B2(n18514), .ZN(
        n18502) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18516), .B1(
        n18603), .B2(n18573), .ZN(n18501) );
  OAI211_X1 U21643 ( .C1(n18576), .C2(n18519), .A(n18502), .B(n18501), .ZN(
        P3_U2973) );
  AOI22_X1 U21644 ( .A1(n18577), .A2(n18514), .B1(n18533), .B2(n18555), .ZN(
        n18504) );
  AOI22_X1 U21645 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18516), .B1(
        n18603), .B2(n18579), .ZN(n18503) );
  OAI211_X1 U21646 ( .C1(n18536), .C2(n18519), .A(n18504), .B(n18503), .ZN(
        P3_U2974) );
  AOI22_X1 U21647 ( .A1(n18537), .A2(n18555), .B1(n18584), .B2(n18514), .ZN(
        n18506) );
  AOI22_X1 U21648 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18516), .B1(
        n18603), .B2(n18585), .ZN(n18505) );
  OAI211_X1 U21649 ( .C1(n18541), .C2(n18519), .A(n18506), .B(n18505), .ZN(
        P3_U2975) );
  AOI22_X1 U21650 ( .A1(n18590), .A2(n18555), .B1(n18589), .B2(n18514), .ZN(
        n18508) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18516), .B1(
        n18603), .B2(n18591), .ZN(n18507) );
  OAI211_X1 U21652 ( .C1(n18594), .C2(n18519), .A(n18508), .B(n18507), .ZN(
        P3_U2976) );
  AOI22_X1 U21653 ( .A1(n18596), .A2(n18555), .B1(n18595), .B2(n18514), .ZN(
        n18510) );
  AOI22_X1 U21654 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18516), .B1(
        n18603), .B2(n18597), .ZN(n18509) );
  OAI211_X1 U21655 ( .C1(n18600), .C2(n18519), .A(n18510), .B(n18509), .ZN(
        P3_U2977) );
  AOI22_X1 U21656 ( .A1(n18550), .A2(n18511), .B1(n18601), .B2(n18514), .ZN(
        n18513) );
  AOI22_X1 U21657 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18516), .B1(
        n18603), .B2(n18604), .ZN(n18512) );
  OAI211_X1 U21658 ( .C1(n18553), .C2(n18540), .A(n18513), .B(n18512), .ZN(
        P3_U2978) );
  AOI22_X1 U21659 ( .A1(n18515), .A2(n18555), .B1(n18610), .B2(n18514), .ZN(
        n18518) );
  AOI22_X1 U21660 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18516), .B1(
        n18603), .B2(n18613), .ZN(n18517) );
  OAI211_X1 U21661 ( .C1(n18520), .C2(n18519), .A(n18518), .B(n18517), .ZN(
        P3_U2979) );
  AND2_X1 U21662 ( .A1(n18560), .A2(n18525), .ZN(n18554) );
  AOI22_X1 U21663 ( .A1(n18561), .A2(n18554), .B1(n18521), .B2(n18611), .ZN(
        n18527) );
  OAI221_X1 U21664 ( .B1(n18525), .B2(n18524), .C1(n18525), .C2(n18523), .A(
        n18522), .ZN(n18557) );
  AOI22_X1 U21665 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18557), .B1(
        n18567), .B2(n18556), .ZN(n18526) );
  OAI211_X1 U21666 ( .C1(n18528), .C2(n18540), .A(n18527), .B(n18526), .ZN(
        P3_U2980) );
  AOI22_X1 U21667 ( .A1(n18529), .A2(n18555), .B1(n18571), .B2(n18554), .ZN(
        n18531) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18557), .B1(
        n18556), .B2(n18573), .ZN(n18530) );
  OAI211_X1 U21669 ( .C1(n18532), .C2(n18607), .A(n18531), .B(n18530), .ZN(
        P3_U2981) );
  AOI22_X1 U21670 ( .A1(n18577), .A2(n18554), .B1(n18533), .B2(n18611), .ZN(
        n18535) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18557), .B1(
        n18556), .B2(n18579), .ZN(n18534) );
  OAI211_X1 U21672 ( .C1(n18536), .C2(n18540), .A(n18535), .B(n18534), .ZN(
        P3_U2982) );
  AOI22_X1 U21673 ( .A1(n18537), .A2(n18611), .B1(n18584), .B2(n18554), .ZN(
        n18539) );
  AOI22_X1 U21674 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18557), .B1(
        n18556), .B2(n18585), .ZN(n18538) );
  OAI211_X1 U21675 ( .C1(n18541), .C2(n18540), .A(n18539), .B(n18538), .ZN(
        P3_U2983) );
  AOI22_X1 U21676 ( .A1(n18542), .A2(n18555), .B1(n18589), .B2(n18554), .ZN(
        n18544) );
  AOI22_X1 U21677 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18557), .B1(
        n18556), .B2(n18591), .ZN(n18543) );
  OAI211_X1 U21678 ( .C1(n18545), .C2(n18607), .A(n18544), .B(n18543), .ZN(
        P3_U2984) );
  AOI22_X1 U21679 ( .A1(n18546), .A2(n18555), .B1(n18595), .B2(n18554), .ZN(
        n18548) );
  AOI22_X1 U21680 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18557), .B1(
        n18556), .B2(n18597), .ZN(n18547) );
  OAI211_X1 U21681 ( .C1(n18549), .C2(n18607), .A(n18548), .B(n18547), .ZN(
        P3_U2985) );
  AOI22_X1 U21682 ( .A1(n18550), .A2(n18555), .B1(n18601), .B2(n18554), .ZN(
        n18552) );
  AOI22_X1 U21683 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18557), .B1(
        n18556), .B2(n18604), .ZN(n18551) );
  OAI211_X1 U21684 ( .C1(n18553), .C2(n18607), .A(n18552), .B(n18551), .ZN(
        P3_U2986) );
  AOI22_X1 U21685 ( .A1(n18612), .A2(n18555), .B1(n18610), .B2(n18554), .ZN(
        n18559) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18557), .B1(
        n18556), .B2(n18613), .ZN(n18558) );
  OAI211_X1 U21687 ( .C1(n18618), .C2(n18607), .A(n18559), .B(n18558), .ZN(
        P3_U2987) );
  AND2_X1 U21688 ( .A1(n18560), .A2(n18563), .ZN(n18609) );
  AOI22_X1 U21689 ( .A1(n18562), .A2(n18611), .B1(n18561), .B2(n18609), .ZN(
        n18569) );
  AOI22_X1 U21690 ( .A1(n18566), .A2(n18565), .B1(n18564), .B2(n18563), .ZN(
        n18615) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18615), .B1(
        n18614), .B2(n18567), .ZN(n18568) );
  OAI211_X1 U21692 ( .C1(n18619), .C2(n18570), .A(n18569), .B(n18568), .ZN(
        P3_U2988) );
  AOI22_X1 U21693 ( .A1(n18603), .A2(n18572), .B1(n18571), .B2(n18609), .ZN(
        n18575) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18615), .B1(
        n18614), .B2(n18573), .ZN(n18574) );
  OAI211_X1 U21695 ( .C1(n18576), .C2(n18607), .A(n18575), .B(n18574), .ZN(
        P3_U2989) );
  AOI22_X1 U21696 ( .A1(n18578), .A2(n18611), .B1(n18577), .B2(n18609), .ZN(
        n18581) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18615), .B1(
        n18614), .B2(n18579), .ZN(n18580) );
  OAI211_X1 U21698 ( .C1(n18619), .C2(n18582), .A(n18581), .B(n18580), .ZN(
        P3_U2990) );
  AOI22_X1 U21699 ( .A1(n18584), .A2(n18609), .B1(n18583), .B2(n18611), .ZN(
        n18587) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18615), .B1(
        n18614), .B2(n18585), .ZN(n18586) );
  OAI211_X1 U21701 ( .C1(n18619), .C2(n18588), .A(n18587), .B(n18586), .ZN(
        P3_U2991) );
  AOI22_X1 U21702 ( .A1(n18603), .A2(n18590), .B1(n18589), .B2(n18609), .ZN(
        n18593) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18615), .B1(
        n18614), .B2(n18591), .ZN(n18592) );
  OAI211_X1 U21704 ( .C1(n18594), .C2(n18607), .A(n18593), .B(n18592), .ZN(
        P3_U2992) );
  AOI22_X1 U21705 ( .A1(n18603), .A2(n18596), .B1(n18595), .B2(n18609), .ZN(
        n18599) );
  AOI22_X1 U21706 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18615), .B1(
        n18614), .B2(n18597), .ZN(n18598) );
  OAI211_X1 U21707 ( .C1(n18600), .C2(n18607), .A(n18599), .B(n18598), .ZN(
        P3_U2993) );
  AOI22_X1 U21708 ( .A1(n18603), .A2(n18602), .B1(n18601), .B2(n18609), .ZN(
        n18606) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18615), .B1(
        n18614), .B2(n18604), .ZN(n18605) );
  OAI211_X1 U21710 ( .C1(n18608), .C2(n18607), .A(n18606), .B(n18605), .ZN(
        P3_U2994) );
  AOI22_X1 U21711 ( .A1(n18612), .A2(n18611), .B1(n18610), .B2(n18609), .ZN(
        n18617) );
  AOI22_X1 U21712 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18615), .B1(
        n18614), .B2(n18613), .ZN(n18616) );
  OAI211_X1 U21713 ( .C1(n18619), .C2(n18618), .A(n18617), .B(n18616), .ZN(
        P3_U2995) );
  INV_X1 U21714 ( .A(n18620), .ZN(n18628) );
  NAND2_X1 U21715 ( .A1(n18621), .A2(n18661), .ZN(n18622) );
  AOI22_X1 U21716 ( .A1(n18625), .A2(n18624), .B1(n18623), .B2(n18622), .ZN(
        n18626) );
  OAI221_X1 U21717 ( .B1(n18628), .B2(n18662), .C1(n18628), .C2(n18627), .A(
        n18626), .ZN(n18833) );
  INV_X1 U21718 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18632) );
  OAI21_X1 U21719 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18629), .ZN(n18631) );
  OAI211_X1 U21720 ( .C1(n18667), .C2(n18632), .A(n18631), .B(n18630), .ZN(
        n18679) );
  NOR2_X1 U21721 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18633), .ZN(
        n18647) );
  INV_X1 U21722 ( .A(n18647), .ZN(n18636) );
  NAND2_X1 U21723 ( .A1(n18807), .A2(n18665), .ZN(n18634) );
  AOI22_X1 U21724 ( .A1(n18641), .A2(n18636), .B1(n18635), .B2(n18634), .ZN(
        n18637) );
  NOR2_X1 U21725 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18637), .ZN(
        n18792) );
  AOI21_X1 U21726 ( .B1(n18640), .B2(n18639), .A(n18638), .ZN(n18655) );
  OAI21_X1 U21727 ( .B1(n18641), .B2(n18646), .A(n18655), .ZN(n18642) );
  AOI22_X1 U21728 ( .A1(n18807), .A2(n18665), .B1(n18643), .B2(n18642), .ZN(
        n18793) );
  NAND2_X1 U21729 ( .A1(n18667), .A2(n18793), .ZN(n18644) );
  AOI22_X1 U21730 ( .A1(n18667), .A2(n18792), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18644), .ZN(n18677) );
  NOR2_X1 U21731 ( .A1(n18656), .A2(n18645), .ZN(n18648) );
  OAI22_X1 U21732 ( .A1(n18820), .A2(n18646), .B1(n18648), .B2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18816) );
  OAI22_X1 U21733 ( .A1(n18648), .A2(n18808), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18647), .ZN(n18812) );
  OAI221_X1 U21734 ( .B1(n18812), .B2(n18816), .C1(n18812), .C2(n18649), .A(
        n18667), .ZN(n18650) );
  INV_X1 U21735 ( .A(n18650), .ZN(n18651) );
  OAI22_X1 U21736 ( .A1(n18653), .A2(n18816), .B1(n18652), .B2(n18651), .ZN(
        n18654) );
  INV_X1 U21737 ( .A(n18654), .ZN(n18671) );
  INV_X1 U21738 ( .A(n18667), .ZN(n18668) );
  AOI221_X1 U21739 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18655), 
        .C1(n18658), .C2(n18655), .A(n18807), .ZN(n18666) );
  NAND2_X1 U21740 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18656), .ZN(
        n18657) );
  AOI211_X1 U21741 ( .C1(n18658), .C2(n18657), .A(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n18814), .ZN(n18664) );
  OAI21_X1 U21742 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n18659), .ZN(n18660) );
  OAI22_X1 U21743 ( .A1(n18803), .A2(n18662), .B1(n18661), .B2(n18660), .ZN(
        n18663) );
  AOI211_X1 U21744 ( .C1(n18666), .C2(n18665), .A(n18664), .B(n18663), .ZN(
        n18799) );
  AOI22_X1 U21745 ( .A1(n18668), .A2(n18807), .B1(n18799), .B2(n18667), .ZN(
        n18672) );
  AND2_X1 U21746 ( .A1(n18671), .A2(n18672), .ZN(n18669) );
  OAI221_X1 U21747 ( .B1(n18671), .B2(n18672), .C1(n18670), .C2(n18669), .A(
        n18674), .ZN(n18676) );
  AOI21_X1 U21748 ( .B1(n18674), .B2(n18673), .A(n18672), .ZN(n18675) );
  AOI222_X1 U21749 ( .A1(n18677), .A2(n18676), .B1(n18677), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18676), .C2(n18675), .ZN(
        n18678) );
  NOR4_X1 U21750 ( .A1(n18680), .A2(n18833), .A3(n18679), .A4(n18678), .ZN(
        n18691) );
  AOI22_X1 U21751 ( .A1(n18815), .A2(n18846), .B1(n18841), .B2(n18835), .ZN(
        n18681) );
  INV_X1 U21752 ( .A(n18681), .ZN(n18686) );
  OAI211_X1 U21753 ( .C1(n18683), .C2(n18682), .A(n18838), .B(n18691), .ZN(
        n18789) );
  OAI21_X1 U21754 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18834), .A(n18789), 
        .ZN(n18692) );
  NOR2_X1 U21755 ( .A1(n18684), .A2(n18692), .ZN(n18685) );
  MUX2_X1 U21756 ( .A(n18686), .B(n18685), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18689) );
  INV_X1 U21757 ( .A(n18687), .ZN(n18688) );
  OAI211_X1 U21758 ( .C1(n18691), .C2(n18690), .A(n18689), .B(n18688), .ZN(
        P3_U2996) );
  NAND2_X1 U21759 ( .A1(n18841), .A2(n18835), .ZN(n18697) );
  NOR4_X1 U21760 ( .A1(n18843), .A2(n18800), .A3(n18834), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18700) );
  INV_X1 U21761 ( .A(n18700), .ZN(n18696) );
  OR3_X1 U21762 ( .A1(n18694), .A2(n18693), .A3(n18692), .ZN(n18695) );
  NAND4_X1 U21763 ( .A1(n18698), .A2(n18697), .A3(n18696), .A4(n18695), .ZN(
        P3_U2997) );
  OAI21_X1 U21764 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18699), .ZN(n18701) );
  AOI21_X1 U21765 ( .B1(n18702), .B2(n18701), .A(n18700), .ZN(P3_U2998) );
  AND2_X1 U21766 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18703), .ZN(
        P3_U2999) );
  AND2_X1 U21767 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18703), .ZN(
        P3_U3000) );
  AND2_X1 U21768 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18703), .ZN(
        P3_U3001) );
  AND2_X1 U21769 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18703), .ZN(
        P3_U3002) );
  AND2_X1 U21770 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18703), .ZN(
        P3_U3003) );
  AND2_X1 U21771 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18703), .ZN(
        P3_U3004) );
  INV_X1 U21772 ( .A(P3_DATAWIDTH_REG_25__SCAN_IN), .ZN(n21065) );
  NOR2_X1 U21773 ( .A1(n21065), .A2(n18787), .ZN(P3_U3005) );
  AND2_X1 U21774 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18703), .ZN(
        P3_U3006) );
  AND2_X1 U21775 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18703), .ZN(
        P3_U3007) );
  AND2_X1 U21776 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18703), .ZN(
        P3_U3008) );
  AND2_X1 U21777 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18703), .ZN(
        P3_U3009) );
  AND2_X1 U21778 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18703), .ZN(
        P3_U3010) );
  AND2_X1 U21779 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18703), .ZN(
        P3_U3011) );
  AND2_X1 U21780 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18703), .ZN(
        P3_U3012) );
  AND2_X1 U21781 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18703), .ZN(
        P3_U3013) );
  AND2_X1 U21782 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18703), .ZN(
        P3_U3014) );
  AND2_X1 U21783 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18703), .ZN(
        P3_U3015) );
  AND2_X1 U21784 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18703), .ZN(
        P3_U3016) );
  AND2_X1 U21785 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18703), .ZN(
        P3_U3017) );
  AND2_X1 U21786 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18703), .ZN(
        P3_U3018) );
  AND2_X1 U21787 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18703), .ZN(
        P3_U3019) );
  AND2_X1 U21788 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18703), .ZN(
        P3_U3020) );
  AND2_X1 U21789 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18703), .ZN(P3_U3021) );
  AND2_X1 U21790 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18703), .ZN(P3_U3022) );
  AND2_X1 U21791 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18703), .ZN(P3_U3023) );
  AND2_X1 U21792 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18703), .ZN(P3_U3024) );
  AND2_X1 U21793 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18703), .ZN(P3_U3025) );
  AND2_X1 U21794 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18703), .ZN(P3_U3026) );
  AND2_X1 U21795 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18703), .ZN(P3_U3027) );
  AND2_X1 U21796 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18703), .ZN(P3_U3028) );
  OAI21_X1 U21797 ( .B1(n18704), .B2(n20809), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18705) );
  AOI22_X1 U21798 ( .A1(n18710), .A2(n18718), .B1(n18849), .B2(n18705), .ZN(
        n18706) );
  INV_X1 U21799 ( .A(NA), .ZN(n20818) );
  OR3_X1 U21800 ( .A1(n20818), .A2(P3_STATE_REG_0__SCAN_IN), .A3(
        P3_STATE_REG_1__SCAN_IN), .ZN(n18709) );
  OAI211_X1 U21801 ( .C1(n18834), .C2(n18707), .A(n18706), .B(n18709), .ZN(
        P3_U3029) );
  OAI22_X1 U21802 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(n20809), .B2(n18718), .ZN(n18712)
         );
  OAI21_X1 U21803 ( .B1(P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18714) );
  INV_X1 U21804 ( .A(n18839), .ZN(n18708) );
  NAND2_X1 U21805 ( .A1(n18841), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18711) );
  OAI211_X1 U21806 ( .C1(n18712), .C2(n18714), .A(n18708), .B(n18711), .ZN(
        P3_U3030) );
  AOI22_X1 U21807 ( .A1(n18841), .A2(P3_STATE_REG_1__SCAN_IN), .B1(n18710), 
        .B2(n18709), .ZN(n18716) );
  INV_X1 U21808 ( .A(n18711), .ZN(n18713) );
  AOI21_X1 U21809 ( .B1(n18713), .B2(n20818), .A(n18712), .ZN(n18715) );
  OAI22_X1 U21810 ( .A1(n18716), .A2(n18718), .B1(n18715), .B2(n18714), .ZN(
        P3_U3031) );
  OAI222_X1 U21811 ( .A1(n18720), .A2(n18781), .B1(n18719), .B2(n18778), .C1(
        n18721), .C2(n18770), .ZN(P3_U3032) );
  OAI222_X1 U21812 ( .A1(n18770), .A2(n21058), .B1(n18722), .B2(n18778), .C1(
        n18721), .C2(n18781), .ZN(P3_U3033) );
  OAI222_X1 U21813 ( .A1(n21058), .A2(n18781), .B1(n18723), .B2(n18778), .C1(
        n18724), .C2(n18770), .ZN(P3_U3034) );
  OAI222_X1 U21814 ( .A1(n18770), .A2(n18727), .B1(n18725), .B2(n18778), .C1(
        n18724), .C2(n18781), .ZN(P3_U3035) );
  OAI222_X1 U21815 ( .A1(n18727), .A2(n18781), .B1(n18726), .B2(n18778), .C1(
        n18728), .C2(n18770), .ZN(P3_U3036) );
  OAI222_X1 U21816 ( .A1(n18770), .A2(n18730), .B1(n18729), .B2(n18778), .C1(
        n18728), .C2(n18781), .ZN(P3_U3037) );
  OAI222_X1 U21817 ( .A1(n18770), .A2(n18732), .B1(n18731), .B2(n18778), .C1(
        n18730), .C2(n18781), .ZN(P3_U3038) );
  OAI222_X1 U21818 ( .A1(n18770), .A2(n18734), .B1(n18733), .B2(n18778), .C1(
        n18732), .C2(n18781), .ZN(P3_U3039) );
  OAI222_X1 U21819 ( .A1(n18770), .A2(n18736), .B1(n18735), .B2(n18778), .C1(
        n18734), .C2(n18781), .ZN(P3_U3040) );
  OAI222_X1 U21820 ( .A1(n18770), .A2(n18738), .B1(n18737), .B2(n18778), .C1(
        n18736), .C2(n18781), .ZN(P3_U3041) );
  INV_X1 U21821 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18740) );
  OAI222_X1 U21822 ( .A1(n18770), .A2(n18740), .B1(n18739), .B2(n18778), .C1(
        n18738), .C2(n18781), .ZN(P3_U3042) );
  OAI222_X1 U21823 ( .A1(n18770), .A2(n18742), .B1(n18741), .B2(n18778), .C1(
        n18740), .C2(n18781), .ZN(P3_U3043) );
  INV_X1 U21824 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18745) );
  OAI222_X1 U21825 ( .A1(n18770), .A2(n18745), .B1(n18743), .B2(n18778), .C1(
        n18742), .C2(n18781), .ZN(P3_U3044) );
  OAI222_X1 U21826 ( .A1(n18745), .A2(n18781), .B1(n18744), .B2(n18778), .C1(
        n18746), .C2(n18770), .ZN(P3_U3045) );
  INV_X1 U21827 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18748) );
  OAI222_X1 U21828 ( .A1(n18770), .A2(n18748), .B1(n18747), .B2(n18778), .C1(
        n18746), .C2(n18781), .ZN(P3_U3046) );
  OAI222_X1 U21829 ( .A1(n18770), .A2(n18750), .B1(n18749), .B2(n18778), .C1(
        n18748), .C2(n18781), .ZN(P3_U3047) );
  OAI222_X1 U21830 ( .A1(n18770), .A2(n18752), .B1(n18751), .B2(n18778), .C1(
        n18750), .C2(n18781), .ZN(P3_U3048) );
  OAI222_X1 U21831 ( .A1(n18770), .A2(n18754), .B1(n18753), .B2(n18778), .C1(
        n18752), .C2(n18781), .ZN(P3_U3049) );
  OAI222_X1 U21832 ( .A1(n18770), .A2(n18756), .B1(n18755), .B2(n18778), .C1(
        n18754), .C2(n18781), .ZN(P3_U3050) );
  OAI222_X1 U21833 ( .A1(n18770), .A2(n18759), .B1(n18757), .B2(n18778), .C1(
        n18756), .C2(n18781), .ZN(P3_U3051) );
  INV_X1 U21834 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18760) );
  OAI222_X1 U21835 ( .A1(n18759), .A2(n18781), .B1(n18758), .B2(n18778), .C1(
        n18760), .C2(n18770), .ZN(P3_U3052) );
  OAI222_X1 U21836 ( .A1(n18770), .A2(n18763), .B1(n18761), .B2(n18778), .C1(
        n18760), .C2(n18781), .ZN(P3_U3053) );
  OAI222_X1 U21837 ( .A1(n18763), .A2(n18781), .B1(n18762), .B2(n18778), .C1(
        n18764), .C2(n18770), .ZN(P3_U3054) );
  OAI222_X1 U21838 ( .A1(n18770), .A2(n18766), .B1(n18765), .B2(n18778), .C1(
        n18764), .C2(n18781), .ZN(P3_U3055) );
  OAI222_X1 U21839 ( .A1(n18770), .A2(n18768), .B1(n18767), .B2(n18778), .C1(
        n18766), .C2(n18781), .ZN(P3_U3056) );
  OAI222_X1 U21840 ( .A1(n18770), .A2(n18771), .B1(n18769), .B2(n18778), .C1(
        n18768), .C2(n18781), .ZN(P3_U3057) );
  OAI222_X1 U21841 ( .A1(n18770), .A2(n18774), .B1(n18772), .B2(n18778), .C1(
        n18771), .C2(n18781), .ZN(P3_U3058) );
  INV_X1 U21842 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18775) );
  OAI222_X1 U21843 ( .A1(n18774), .A2(n18781), .B1(n18773), .B2(n18778), .C1(
        n18775), .C2(n18770), .ZN(P3_U3059) );
  OAI222_X1 U21844 ( .A1(n18770), .A2(n18780), .B1(n18776), .B2(n18778), .C1(
        n18775), .C2(n18781), .ZN(P3_U3060) );
  OAI222_X1 U21845 ( .A1(n18781), .A2(n18780), .B1(n18779), .B2(n18778), .C1(
        n18777), .C2(n18770), .ZN(P3_U3061) );
  MUX2_X1 U21846 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .B(P3_BE_N_REG_3__SCAN_IN), .S(n18849), .Z(P3_U3274) );
  MUX2_X1 U21847 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .B(P3_BE_N_REG_2__SCAN_IN), .S(n18849), .Z(P3_U3275) );
  OAI22_X1 U21848 ( .A1(n18849), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18778), .ZN(n18782) );
  INV_X1 U21849 ( .A(n18782), .ZN(P3_U3276) );
  OAI22_X1 U21850 ( .A1(n18849), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18778), .ZN(n18783) );
  INV_X1 U21851 ( .A(n18783), .ZN(P3_U3277) );
  OAI21_X1 U21852 ( .B1(n18787), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18785), 
        .ZN(n18784) );
  INV_X1 U21853 ( .A(n18784), .ZN(P3_U3280) );
  OAI21_X1 U21854 ( .B1(n18787), .B2(n18786), .A(n18785), .ZN(P3_U3281) );
  OAI221_X1 U21855 ( .B1(n18790), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18790), 
        .C2(n18789), .A(n18788), .ZN(P3_U3282) );
  AOI22_X1 U21856 ( .A1(n18852), .A2(n18792), .B1(n18815), .B2(n18791), .ZN(
        n18798) );
  INV_X1 U21857 ( .A(n18821), .ZN(n18818) );
  OAI21_X1 U21858 ( .B1(n18794), .B2(n18793), .A(n18818), .ZN(n18795) );
  INV_X1 U21859 ( .A(n18795), .ZN(n18797) );
  OAI22_X1 U21860 ( .A1(n18821), .A2(n18798), .B1(n18797), .B2(n18796), .ZN(
        P3_U3285) );
  INV_X1 U21861 ( .A(n18799), .ZN(n18805) );
  NOR2_X1 U21862 ( .A1(n18800), .A2(n18817), .ZN(n18809) );
  OAI22_X1 U21863 ( .A1(n18802), .A2(n18801), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18810) );
  INV_X1 U21864 ( .A(n18810), .ZN(n18804) );
  AOI222_X1 U21865 ( .A1(n18805), .A2(n18852), .B1(n18809), .B2(n18804), .C1(
        n18815), .C2(n18803), .ZN(n18806) );
  AOI22_X1 U21866 ( .A1(n18821), .A2(n18807), .B1(n18806), .B2(n18818), .ZN(
        P3_U3288) );
  INV_X1 U21867 ( .A(n18808), .ZN(n18811) );
  AOI222_X1 U21868 ( .A1(n18812), .A2(n18852), .B1(n18815), .B2(n18811), .C1(
        n18810), .C2(n18809), .ZN(n18813) );
  AOI22_X1 U21869 ( .A1(n18821), .A2(n18814), .B1(n18813), .B2(n18818), .ZN(
        P3_U3289) );
  AOI222_X1 U21870 ( .A1(n18817), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18852), 
        .B2(n18816), .C1(n18820), .C2(n18815), .ZN(n18819) );
  AOI22_X1 U21871 ( .A1(n18821), .A2(n18820), .B1(n18819), .B2(n18818), .ZN(
        P3_U3290) );
  INV_X1 U21872 ( .A(n18822), .ZN(n18829) );
  AOI211_X1 U21873 ( .C1(P3_REIP_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_REIP_REG_1__SCAN_IN), .B(n18823), 
        .ZN(n18824) );
  AOI21_X1 U21874 ( .B1(P3_BYTEENABLE_REG_2__SCAN_IN), .B2(n18829), .A(n18824), 
        .ZN(n18825) );
  OAI21_X1 U21875 ( .B1(n18828), .B2(n18826), .A(n18825), .ZN(P3_U3292) );
  INV_X1 U21876 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18830) );
  NOR2_X1 U21877 ( .A1(n18829), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18827) );
  AOI22_X1 U21878 ( .A1(n18830), .A2(n18829), .B1(n18828), .B2(n18827), .ZN(
        P3_U3293) );
  INV_X1 U21879 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18855) );
  OAI22_X1 U21880 ( .A1(n18849), .A2(n18855), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n18778), .ZN(n18831) );
  INV_X1 U21881 ( .A(n18831), .ZN(P3_U3294) );
  MUX2_X1 U21882 ( .A(P3_MORE_REG_SCAN_IN), .B(n18833), .S(n18832), .Z(
        P3_U3295) );
  AOI21_X1 U21883 ( .B1(n18835), .B2(n18834), .A(n18854), .ZN(n18836) );
  OAI21_X1 U21884 ( .B1(n18838), .B2(n18837), .A(n18836), .ZN(n18848) );
  INV_X1 U21885 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n20937) );
  OAI21_X1 U21886 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n18840), .A(n18839), 
        .ZN(n18842) );
  AOI211_X1 U21887 ( .C1(n18853), .C2(n18842), .A(n18841), .B(n18851), .ZN(
        n18844) );
  NOR2_X1 U21888 ( .A1(n18844), .A2(n18843), .ZN(n18845) );
  OAI21_X1 U21889 ( .B1(n18846), .B2(n18845), .A(n18848), .ZN(n18847) );
  OAI21_X1 U21890 ( .B1(n18848), .B2(n20937), .A(n18847), .ZN(P3_U3296) );
  OAI22_X1 U21891 ( .A1(n18849), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18778), .ZN(n18850) );
  INV_X1 U21892 ( .A(n18850), .ZN(P3_U3297) );
  AOI21_X1 U21893 ( .B1(n18852), .B2(n18851), .A(n18854), .ZN(n18858) );
  AOI22_X1 U21894 ( .A1(n18858), .A2(n18855), .B1(n18854), .B2(n18853), .ZN(
        P3_U3298) );
  INV_X1 U21895 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18857) );
  AOI21_X1 U21896 ( .B1(n18858), .B2(n18857), .A(n18856), .ZN(P3_U3299) );
  INV_X1 U21897 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19732) );
  NAND2_X1 U21898 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19752), .ZN(n19741) );
  NAND2_X1 U21899 ( .A1(n19732), .A2(n18859), .ZN(n19738) );
  OAI21_X1 U21900 ( .B1(n19732), .B2(n19741), .A(n19738), .ZN(n19816) );
  AOI21_X1 U21901 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19816), .ZN(n18860) );
  INV_X1 U21902 ( .A(n18860), .ZN(P2_U2815) );
  INV_X1 U21903 ( .A(n18861), .ZN(n18863) );
  INV_X1 U21904 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n20921) );
  OAI22_X1 U21905 ( .A1(n18863), .A2(n20921), .B1(n16342), .B2(n18862), .ZN(
        P2_U2816) );
  NAND2_X1 U21906 ( .A1(n19732), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19867) );
  INV_X2 U21907 ( .A(n19867), .ZN(n19866) );
  AOI21_X1 U21908 ( .B1(n19732), .B2(n19752), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18864) );
  AOI22_X1 U21909 ( .A1(n19866), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18864), 
        .B2(n19867), .ZN(P2_U2817) );
  OAI21_X1 U21910 ( .B1(n19745), .B2(BS16), .A(n19816), .ZN(n19814) );
  OAI21_X1 U21911 ( .B1(n19816), .B2(n19818), .A(n19814), .ZN(P2_U2818) );
  NOR4_X1 U21912 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18868) );
  NOR4_X1 U21913 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18867) );
  NOR4_X1 U21914 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18866) );
  NOR4_X1 U21915 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18865) );
  NAND4_X1 U21916 ( .A1(n18868), .A2(n18867), .A3(n18866), .A4(n18865), .ZN(
        n18874) );
  NOR4_X1 U21917 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18872) );
  AOI211_X1 U21918 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_16__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18871) );
  NOR4_X1 U21919 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18870) );
  NOR4_X1 U21920 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18869) );
  NAND4_X1 U21921 ( .A1(n18872), .A2(n18871), .A3(n18870), .A4(n18869), .ZN(
        n18873) );
  NOR2_X1 U21922 ( .A1(n18874), .A2(n18873), .ZN(n18884) );
  INV_X1 U21923 ( .A(n18884), .ZN(n18882) );
  NOR2_X1 U21924 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18882), .ZN(n18877) );
  INV_X1 U21925 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18875) );
  AOI22_X1 U21926 ( .A1(n18877), .A2(n12852), .B1(n18882), .B2(n18875), .ZN(
        P2_U2820) );
  OR3_X1 U21927 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18881) );
  INV_X1 U21928 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18876) );
  AOI22_X1 U21929 ( .A1(n18877), .A2(n18881), .B1(n18882), .B2(n18876), .ZN(
        P2_U2821) );
  INV_X1 U21930 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19815) );
  NAND2_X1 U21931 ( .A1(n18877), .A2(n19815), .ZN(n18880) );
  OAI21_X1 U21932 ( .B1(n12852), .B2(n19753), .A(n18884), .ZN(n18878) );
  OAI21_X1 U21933 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18884), .A(n18878), 
        .ZN(n18879) );
  OAI221_X1 U21934 ( .B1(n18880), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18880), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18879), .ZN(P2_U2822) );
  INV_X1 U21935 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18883) );
  OAI221_X1 U21936 ( .B1(n18884), .B2(n18883), .C1(n18882), .C2(n18881), .A(
        n18880), .ZN(P2_U2823) );
  AOI22_X1 U21937 ( .A1(P2_REIP_REG_21__SCAN_IN), .A2(n19045), .B1(
        P2_EBX_REG_21__SCAN_IN), .B2(n19059), .ZN(n18889) );
  OAI211_X1 U21938 ( .C1(n18887), .C2(n18886), .A(n19036), .B(n18885), .ZN(
        n18888) );
  OAI211_X1 U21939 ( .C1(n19071), .C2(n18890), .A(n18889), .B(n18888), .ZN(
        n18894) );
  OAI22_X1 U21940 ( .A1(n18892), .A2(n19043), .B1(n18891), .B2(n19011), .ZN(
        n18893) );
  AOI211_X1 U21941 ( .C1(n18895), .C2(n19061), .A(n18894), .B(n18893), .ZN(
        n18896) );
  INV_X1 U21942 ( .A(n18896), .ZN(P2_U2834) );
  NOR2_X1 U21943 ( .A1(n19041), .A2(n18897), .ZN(n18899) );
  XOR2_X1 U21944 ( .A(n18899), .B(n18898), .Z(n18908) );
  AOI22_X1 U21945 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(n19059), .B1(n18900), 
        .B2(n19057), .ZN(n18901) );
  OAI211_X1 U21946 ( .C1(n15192), .C2(n19068), .A(n18901), .B(n19046), .ZN(
        n18902) );
  AOI21_X1 U21947 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n19028), .A(
        n18902), .ZN(n18907) );
  OAI22_X1 U21948 ( .A1(n18904), .A2(n19049), .B1(n18903), .B2(n19011), .ZN(
        n18905) );
  INV_X1 U21949 ( .A(n18905), .ZN(n18906) );
  OAI211_X1 U21950 ( .C1(n19077), .C2(n18908), .A(n18907), .B(n18906), .ZN(
        P2_U2837) );
  INV_X1 U21951 ( .A(n18909), .ZN(n18912) );
  NAND2_X1 U21952 ( .A1(n18910), .A2(n18912), .ZN(n18931) );
  AOI211_X1 U21953 ( .C1(n11360), .C2(n18912), .A(n18911), .B(n19077), .ZN(
        n18916) );
  AOI22_X1 U21954 ( .A1(P2_REIP_REG_16__SCAN_IN), .A2(n19045), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n19028), .ZN(n18913) );
  OAI211_X1 U21955 ( .C1(n18914), .C2(n19043), .A(n18913), .B(n19046), .ZN(
        n18915) );
  AOI211_X1 U21956 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n19059), .A(n18916), .B(
        n18915), .ZN(n18919) );
  OAI22_X1 U21957 ( .A1(n19113), .A2(n19049), .B1(n19082), .B2(n19011), .ZN(
        n18917) );
  INV_X1 U21958 ( .A(n18917), .ZN(n18918) );
  OAI211_X1 U21959 ( .C1(n18920), .C2(n18931), .A(n18919), .B(n18918), .ZN(
        P2_U2839) );
  INV_X1 U21960 ( .A(n18930), .ZN(n18922) );
  AOI22_X1 U21961 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_15__SCAN_IN), .B2(n19045), .ZN(n18921) );
  OAI211_X1 U21962 ( .C1(n18922), .C2(n18943), .A(n18921), .B(n19046), .ZN(
        n18927) );
  OAI22_X1 U21963 ( .A1(n19001), .A2(n10821), .B1(n18923), .B2(n19043), .ZN(
        n18926) );
  OAI22_X1 U21964 ( .A1(n19119), .A2(n19049), .B1(n18924), .B2(n19011), .ZN(
        n18925) );
  NOR3_X1 U21965 ( .A1(n18927), .A2(n18926), .A3(n18925), .ZN(n18928) );
  OAI221_X1 U21966 ( .B1(n18931), .B2(n18930), .C1(n18931), .C2(n18929), .A(
        n18928), .ZN(P2_U2840) );
  NOR2_X1 U21967 ( .A1(n19041), .A2(n18932), .ZN(n18951) );
  XOR2_X1 U21968 ( .A(n18951), .B(n18933), .Z(n18940) );
  AOI22_X1 U21969 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n19028), .B1(
        P2_EBX_REG_14__SCAN_IN), .B2(n19059), .ZN(n18934) );
  OAI21_X1 U21970 ( .B1(n18935), .B2(n19043), .A(n18934), .ZN(n18936) );
  AOI211_X1 U21971 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n19045), .A(n19217), 
        .B(n18936), .ZN(n18939) );
  AOI22_X1 U21972 ( .A1(n19120), .A2(n19061), .B1(n18937), .B2(n19064), .ZN(
        n18938) );
  OAI211_X1 U21973 ( .C1(n19077), .C2(n18940), .A(n18939), .B(n18938), .ZN(
        P2_U2841) );
  AOI22_X1 U21974 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19045), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19028), .ZN(n18947) );
  INV_X1 U21975 ( .A(n18941), .ZN(n18952) );
  AOI21_X1 U21976 ( .B1(n19059), .B2(P2_EBX_REG_13__SCAN_IN), .A(n19217), .ZN(
        n18942) );
  OAI21_X1 U21977 ( .B1(n18952), .B2(n18943), .A(n18942), .ZN(n18944) );
  AOI21_X1 U21978 ( .B1(n18945), .B2(n19064), .A(n18944), .ZN(n18946) );
  OAI211_X1 U21979 ( .C1(n18948), .C2(n19043), .A(n18947), .B(n18946), .ZN(
        n18949) );
  INV_X1 U21980 ( .A(n18949), .ZN(n18955) );
  INV_X1 U21981 ( .A(n18950), .ZN(n18953) );
  OAI211_X1 U21982 ( .C1(n18953), .C2(n18952), .A(n19036), .B(n18951), .ZN(
        n18954) );
  OAI211_X1 U21983 ( .C1(n19049), .C2(n19125), .A(n18955), .B(n18954), .ZN(
        P2_U2842) );
  AOI22_X1 U21984 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19028), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n19059), .ZN(n18956) );
  OAI21_X1 U21985 ( .B1(n18957), .B2(n19043), .A(n18956), .ZN(n18958) );
  AOI211_X1 U21986 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19045), .A(n19217), 
        .B(n18958), .ZN(n18965) );
  NOR2_X1 U21987 ( .A1(n19041), .A2(n18959), .ZN(n18961) );
  XNOR2_X1 U21988 ( .A(n18961), .B(n18960), .ZN(n18963) );
  AOI22_X1 U21989 ( .A1(n18963), .A2(n19036), .B1(n18962), .B2(n19064), .ZN(
        n18964) );
  OAI211_X1 U21990 ( .C1(n19128), .C2(n19049), .A(n18965), .B(n18964), .ZN(
        P2_U2843) );
  AOI22_X1 U21991 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n19059), .B1(n18966), 
        .B2(n19057), .ZN(n18967) );
  OAI21_X1 U21992 ( .B1(n10861), .B2(n19071), .A(n18967), .ZN(n18968) );
  AOI211_X1 U21993 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n19045), .A(n19217), 
        .B(n18968), .ZN(n18975) );
  NAND2_X1 U21994 ( .A1(n11360), .A2(n18969), .ZN(n18970) );
  XNOR2_X1 U21995 ( .A(n18971), .B(n18970), .ZN(n18973) );
  AOI22_X1 U21996 ( .A1(n18973), .A2(n19036), .B1(n18972), .B2(n19064), .ZN(
        n18974) );
  OAI211_X1 U21997 ( .C1(n19130), .C2(n19049), .A(n18975), .B(n18974), .ZN(
        P2_U2844) );
  NOR2_X1 U21998 ( .A1(n19041), .A2(n18976), .ZN(n18978) );
  XOR2_X1 U21999 ( .A(n18978), .B(n18977), .Z(n18985) );
  OAI21_X1 U22000 ( .B1(n19770), .B2(n19068), .A(n19046), .ZN(n18981) );
  OAI22_X1 U22001 ( .A1(n19001), .A2(n10857), .B1(n18979), .B2(n19043), .ZN(
        n18980) );
  AOI211_X1 U22002 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n19028), .A(
        n18981), .B(n18980), .ZN(n18984) );
  INV_X1 U22003 ( .A(n19090), .ZN(n18982) );
  AOI22_X1 U22004 ( .A1(n19131), .A2(n19061), .B1(n18982), .B2(n19064), .ZN(
        n18983) );
  OAI211_X1 U22005 ( .C1(n19077), .C2(n18985), .A(n18984), .B(n18983), .ZN(
        P2_U2845) );
  NAND2_X1 U22006 ( .A1(n9690), .A2(n18986), .ZN(n18988) );
  XOR2_X1 U22007 ( .A(n18988), .B(n18987), .Z(n18995) );
  AOI22_X1 U22008 ( .A1(P2_EBX_REG_9__SCAN_IN), .A2(n19059), .B1(n19057), .B2(
        n18989), .ZN(n18990) );
  OAI211_X1 U22009 ( .C1(n19768), .C2(n19068), .A(n18990), .B(n19046), .ZN(
        n18993) );
  OAI22_X1 U22010 ( .A1(n19136), .A2(n19049), .B1(n18991), .B2(n19011), .ZN(
        n18992) );
  AOI211_X1 U22011 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19028), .A(
        n18993), .B(n18992), .ZN(n18994) );
  OAI21_X1 U22012 ( .B1(n18995), .B2(n19077), .A(n18994), .ZN(P2_U2846) );
  NOR2_X1 U22013 ( .A1(n19041), .A2(n18996), .ZN(n18998) );
  XOR2_X1 U22014 ( .A(n18998), .B(n18997), .Z(n19005) );
  AOI22_X1 U22015 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19028), .B1(
        n18999), .B2(n19057), .ZN(n19000) );
  OAI21_X1 U22016 ( .B1(n19001), .B2(n10853), .A(n19000), .ZN(n19002) );
  AOI211_X1 U22017 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19045), .A(n19217), .B(
        n19002), .ZN(n19004) );
  AOI22_X1 U22018 ( .A1(n19098), .A2(n19064), .B1(n19061), .B2(n19137), .ZN(
        n19003) );
  OAI211_X1 U22019 ( .C1(n19077), .C2(n19005), .A(n19004), .B(n19003), .ZN(
        P2_U2847) );
  NAND2_X1 U22020 ( .A1(n9690), .A2(n19006), .ZN(n19008) );
  XOR2_X1 U22021 ( .A(n19008), .B(n19007), .Z(n19016) );
  AOI22_X1 U22022 ( .A1(P2_EBX_REG_7__SCAN_IN), .A2(n19059), .B1(n19009), .B2(
        n19057), .ZN(n19010) );
  OAI211_X1 U22023 ( .C1(n19764), .C2(n19068), .A(n19010), .B(n19046), .ZN(
        n19014) );
  OAI22_X1 U22024 ( .A1(n19141), .A2(n19049), .B1(n19012), .B2(n19011), .ZN(
        n19013) );
  AOI211_X1 U22025 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19028), .A(
        n19014), .B(n19013), .ZN(n19015) );
  OAI21_X1 U22026 ( .B1(n19016), .B2(n19077), .A(n19015), .ZN(P2_U2848) );
  OAI21_X1 U22027 ( .B1(n19762), .B2(n19068), .A(n19046), .ZN(n19020) );
  AOI22_X1 U22028 ( .A1(n19059), .A2(P2_EBX_REG_6__SCAN_IN), .B1(n19017), .B2(
        n19057), .ZN(n19018) );
  INV_X1 U22029 ( .A(n19018), .ZN(n19019) );
  AOI211_X1 U22030 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19028), .A(
        n19020), .B(n19019), .ZN(n19027) );
  NOR2_X1 U22031 ( .A1(n19041), .A2(n19021), .ZN(n19023) );
  XNOR2_X1 U22032 ( .A(n19023), .B(n19022), .ZN(n19025) );
  AOI22_X1 U22033 ( .A1(n19025), .A2(n19036), .B1(n19064), .B2(n19024), .ZN(
        n19026) );
  OAI211_X1 U22034 ( .C1(n19049), .C2(n19142), .A(n19027), .B(n19026), .ZN(
        P2_U2849) );
  AOI22_X1 U22035 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19028), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(n19059), .ZN(n19029) );
  OAI21_X1 U22036 ( .B1(n19030), .B2(n19043), .A(n19029), .ZN(n19031) );
  AOI211_X1 U22037 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19045), .A(n19217), .B(
        n19031), .ZN(n19039) );
  NAND2_X1 U22038 ( .A1(n11360), .A2(n19032), .ZN(n19033) );
  XNOR2_X1 U22039 ( .A(n19034), .B(n19033), .ZN(n19037) );
  AOI22_X1 U22040 ( .A1(n19037), .A2(n19036), .B1(n19064), .B2(n19035), .ZN(
        n19038) );
  OAI211_X1 U22041 ( .C1(n19049), .C2(n19150), .A(n19039), .B(n19038), .ZN(
        P2_U2850) );
  NOR2_X1 U22042 ( .A1(n19041), .A2(n19040), .ZN(n19042) );
  XOR2_X1 U22043 ( .A(n19042), .B(n19228), .Z(n19054) );
  NOR2_X1 U22044 ( .A1(n19044), .A2(n19043), .ZN(n19051) );
  AOI22_X1 U22045 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19028), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19045), .ZN(n19047) );
  OAI211_X1 U22046 ( .C1(n19049), .C2(n19048), .A(n19047), .B(n19046), .ZN(
        n19050) );
  AOI211_X1 U22047 ( .C1(P2_EBX_REG_4__SCAN_IN), .C2(n19059), .A(n19051), .B(
        n19050), .ZN(n19053) );
  INV_X1 U22048 ( .A(n19146), .ZN(n19101) );
  AOI22_X1 U22049 ( .A1(n19101), .A2(n19074), .B1(n19064), .B2(n19224), .ZN(
        n19052) );
  OAI211_X1 U22050 ( .C1(n19077), .C2(n19054), .A(n19053), .B(n19052), .ZN(
        P2_U2851) );
  NAND2_X1 U22051 ( .A1(n19057), .A2(n19056), .ZN(n19063) );
  AOI22_X1 U22052 ( .A1(n19061), .A2(n19060), .B1(P2_EBX_REG_0__SCAN_IN), .B2(
        n19059), .ZN(n19062) );
  AND2_X1 U22053 ( .A1(n19063), .A2(n19062), .ZN(n19067) );
  NAND2_X1 U22054 ( .A1(n9647), .A2(n19064), .ZN(n19066) );
  OAI211_X1 U22055 ( .C1(n19068), .C2(n12852), .A(n19067), .B(n19066), .ZN(
        n19069) );
  INV_X1 U22056 ( .A(n19069), .ZN(n19076) );
  INV_X1 U22057 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19070) );
  NOR2_X1 U22058 ( .A1(n19071), .A2(n19070), .ZN(n19072) );
  AOI21_X1 U22059 ( .B1(n19074), .B2(n19073), .A(n19072), .ZN(n19075) );
  OAI211_X1 U22060 ( .C1(n19077), .C2(n15450), .A(n19076), .B(n19075), .ZN(
        P2_U2855) );
  OR2_X1 U22061 ( .A1(n13837), .A2(n19078), .ZN(n19080) );
  NAND2_X1 U22062 ( .A1(n19080), .A2(n19079), .ZN(n19081) );
  NAND2_X1 U22063 ( .A1(n13860), .A2(n19081), .ZN(n19112) );
  OAI22_X1 U22064 ( .A1(n19112), .A2(n19095), .B1(n19089), .B2(n19082), .ZN(
        n19083) );
  INV_X1 U22065 ( .A(n19083), .ZN(n19084) );
  OAI21_X1 U22066 ( .B1(n19103), .B2(n10877), .A(n19084), .ZN(P2_U2871) );
  AOI21_X1 U22067 ( .B1(n9751), .B2(n19086), .A(n19085), .ZN(n19087) );
  OR3_X1 U22068 ( .A1(n19087), .A2(n9752), .A3(n19095), .ZN(n19088) );
  OAI21_X1 U22069 ( .B1(n19090), .B2(n19089), .A(n19088), .ZN(n19091) );
  INV_X1 U22070 ( .A(n19091), .ZN(n19092) );
  OAI21_X1 U22071 ( .B1(n19103), .B2(n10857), .A(n19092), .ZN(P2_U2877) );
  AOI21_X1 U22072 ( .B1(n19094), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A(
        n19093), .ZN(n19096) );
  NOR3_X1 U22073 ( .A1(n19096), .A2(n9751), .A3(n19095), .ZN(n19097) );
  AOI21_X1 U22074 ( .B1(n19098), .B2(n19103), .A(n19097), .ZN(n19099) );
  OAI21_X1 U22075 ( .B1(n19103), .B2(n10853), .A(n19099), .ZN(P2_U2879) );
  AOI22_X1 U22076 ( .A1(n19101), .A2(n19100), .B1(n19103), .B2(n19224), .ZN(
        n19102) );
  OAI21_X1 U22077 ( .B1(n19103), .B2(n10549), .A(n19102), .ZN(P2_U2883) );
  AOI22_X1 U22078 ( .A1(n19104), .A2(n19171), .B1(n19110), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n19106) );
  AOI22_X1 U22079 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19170), .B1(n19111), 
        .B2(BUF2_REG_31__SCAN_IN), .ZN(n19105) );
  NAND2_X1 U22080 ( .A1(n19106), .A2(n19105), .ZN(P2_U2888) );
  INV_X1 U22081 ( .A(n19107), .ZN(n19108) );
  AOI22_X1 U22082 ( .A1(n19109), .A2(n19108), .B1(n19170), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19117) );
  AOI22_X1 U22083 ( .A1(n19111), .A2(BUF2_REG_16__SCAN_IN), .B1(n19110), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19116) );
  OAI22_X1 U22084 ( .A1(n19113), .A2(n19153), .B1(n19145), .B2(n19112), .ZN(
        n19114) );
  INV_X1 U22085 ( .A(n19114), .ZN(n19115) );
  NAND3_X1 U22086 ( .A1(n19117), .A2(n19116), .A3(n19115), .ZN(P2_U2903) );
  OAI222_X1 U22087 ( .A1(n19119), .A2(n19151), .B1(n19185), .B2(n19169), .C1(
        n19118), .C2(n19179), .ZN(P2_U2904) );
  INV_X1 U22088 ( .A(n19120), .ZN(n19123) );
  AOI22_X1 U22089 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19170), .B1(n19121), 
        .B2(n19161), .ZN(n19122) );
  OAI21_X1 U22090 ( .B1(n19151), .B2(n19123), .A(n19122), .ZN(P2_U2905) );
  INV_X1 U22091 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n21088) );
  OAI222_X1 U22092 ( .A1(n19125), .A2(n19151), .B1(n21088), .B2(n19169), .C1(
        n19179), .C2(n19124), .ZN(P2_U2906) );
  AOI22_X1 U22093 ( .A1(P2_EAX_REG_12__SCAN_IN), .A2(n19170), .B1(n19126), 
        .B2(n19161), .ZN(n19127) );
  OAI21_X1 U22094 ( .B1(n19151), .B2(n19128), .A(n19127), .ZN(P2_U2907) );
  INV_X1 U22095 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19193) );
  OAI222_X1 U22096 ( .A1(n19130), .A2(n19151), .B1(n19193), .B2(n19169), .C1(
        n19179), .C2(n19129), .ZN(P2_U2908) );
  INV_X1 U22097 ( .A(n19131), .ZN(n19134) );
  AOI22_X1 U22098 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19170), .B1(n19132), 
        .B2(n19161), .ZN(n19133) );
  OAI21_X1 U22099 ( .B1(n19151), .B2(n19134), .A(n19133), .ZN(P2_U2909) );
  INV_X1 U22100 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19197) );
  OAI222_X1 U22101 ( .A1(n19136), .A2(n19151), .B1(n19197), .B2(n19169), .C1(
        n19179), .C2(n19135), .ZN(P2_U2910) );
  INV_X1 U22102 ( .A(n19137), .ZN(n19140) );
  AOI22_X1 U22103 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19170), .B1(n19138), .B2(
        n19161), .ZN(n19139) );
  OAI21_X1 U22104 ( .B1(n19151), .B2(n19140), .A(n19139), .ZN(P2_U2911) );
  OAI222_X1 U22105 ( .A1(n19141), .A2(n19151), .B1(n19201), .B2(n19169), .C1(
        n19179), .C2(n19259), .ZN(P2_U2912) );
  OAI222_X1 U22106 ( .A1(n19142), .A2(n19151), .B1(n19203), .B2(n19169), .C1(
        n19179), .C2(n19252), .ZN(P2_U2913) );
  INV_X1 U22107 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19205) );
  OAI22_X1 U22108 ( .A1(n19205), .A2(n19169), .B1(n19143), .B2(n19179), .ZN(
        n19144) );
  INV_X1 U22109 ( .A(n19144), .ZN(n19149) );
  OR3_X1 U22110 ( .A1(n19147), .A2(n19146), .A3(n19145), .ZN(n19148) );
  OAI211_X1 U22111 ( .C1(n19151), .C2(n19150), .A(n19149), .B(n19148), .ZN(
        P2_U2914) );
  INV_X1 U22112 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19152) );
  OAI22_X1 U22113 ( .A1(n19826), .A2(n19153), .B1(n19169), .B2(n19152), .ZN(
        n19154) );
  INV_X1 U22114 ( .A(n19154), .ZN(n19160) );
  OAI21_X1 U22115 ( .B1(n19157), .B2(n19156), .A(n19155), .ZN(n19158) );
  NAND2_X1 U22116 ( .A1(n19158), .A2(n19175), .ZN(n19159) );
  OAI211_X1 U22117 ( .C1(n19240), .C2(n19179), .A(n19160), .B(n19159), .ZN(
        P2_U2916) );
  AOI22_X1 U22118 ( .A1(n19835), .A2(n19171), .B1(n19162), .B2(n19161), .ZN(
        n19168) );
  OAI21_X1 U22119 ( .B1(n19165), .B2(n19164), .A(n19163), .ZN(n19166) );
  NAND2_X1 U22120 ( .A1(n19166), .A2(n19175), .ZN(n19167) );
  OAI211_X1 U22121 ( .C1(n19169), .C2(n19209), .A(n19168), .B(n19167), .ZN(
        P2_U2917) );
  AOI22_X1 U22122 ( .A1(n19171), .A2(n19844), .B1(n19170), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19178) );
  OAI21_X1 U22123 ( .B1(n19174), .B2(n19173), .A(n19172), .ZN(n19176) );
  NAND2_X1 U22124 ( .A1(n19176), .A2(n19175), .ZN(n19177) );
  OAI211_X1 U22125 ( .C1(n19232), .C2(n19179), .A(n19178), .B(n19177), .ZN(
        P2_U2918) );
  NOR2_X1 U22126 ( .A1(n19183), .A2(n19180), .ZN(P2_U2920) );
  AOI22_X1 U22127 ( .A1(n19181), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n19214), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n19182) );
  OAI21_X1 U22128 ( .B1(n20956), .B2(n19183), .A(n19182), .ZN(P2_U2931) );
  AOI22_X1 U22129 ( .A1(n19214), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19184) );
  OAI21_X1 U22130 ( .B1(n19185), .B2(n19216), .A(n19184), .ZN(P2_U2936) );
  AOI22_X1 U22131 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19186), .B1(n19213), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19187) );
  OAI21_X1 U22132 ( .B1(n20924), .B2(n19188), .A(n19187), .ZN(P2_U2937) );
  AOI22_X1 U22133 ( .A1(n19214), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19189) );
  OAI21_X1 U22134 ( .B1(n21088), .B2(n19216), .A(n19189), .ZN(P2_U2938) );
  AOI22_X1 U22135 ( .A1(n19214), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19190) );
  OAI21_X1 U22136 ( .B1(n19191), .B2(n19216), .A(n19190), .ZN(P2_U2939) );
  AOI22_X1 U22137 ( .A1(n19214), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19192) );
  OAI21_X1 U22138 ( .B1(n19193), .B2(n19216), .A(n19192), .ZN(P2_U2940) );
  AOI22_X1 U22139 ( .A1(n19214), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19194) );
  OAI21_X1 U22140 ( .B1(n19195), .B2(n19216), .A(n19194), .ZN(P2_U2941) );
  AOI22_X1 U22141 ( .A1(n19214), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19196) );
  OAI21_X1 U22142 ( .B1(n19197), .B2(n19216), .A(n19196), .ZN(P2_U2942) );
  AOI22_X1 U22143 ( .A1(n19214), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19198) );
  OAI21_X1 U22144 ( .B1(n19199), .B2(n19216), .A(n19198), .ZN(P2_U2943) );
  AOI22_X1 U22145 ( .A1(n19214), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19200) );
  OAI21_X1 U22146 ( .B1(n19201), .B2(n19216), .A(n19200), .ZN(P2_U2944) );
  AOI22_X1 U22147 ( .A1(n19214), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19202) );
  OAI21_X1 U22148 ( .B1(n19203), .B2(n19216), .A(n19202), .ZN(P2_U2945) );
  AOI22_X1 U22149 ( .A1(n19214), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19204) );
  OAI21_X1 U22150 ( .B1(n19205), .B2(n19216), .A(n19204), .ZN(P2_U2946) );
  AOI22_X1 U22151 ( .A1(n19214), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19206) );
  OAI21_X1 U22152 ( .B1(n12897), .B2(n19216), .A(n19206), .ZN(P2_U2947) );
  AOI22_X1 U22153 ( .A1(n19214), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19207) );
  OAI21_X1 U22154 ( .B1(n19152), .B2(n19216), .A(n19207), .ZN(P2_U2948) );
  AOI22_X1 U22155 ( .A1(n19214), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19208) );
  OAI21_X1 U22156 ( .B1(n19209), .B2(n19216), .A(n19208), .ZN(P2_U2949) );
  AOI22_X1 U22157 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(n19213), .B1(n19210), 
        .B2(P2_LWORD_REG_1__SCAN_IN), .ZN(n19211) );
  OAI21_X1 U22158 ( .B1(n19212), .B2(n19216), .A(n19211), .ZN(P2_U2950) );
  AOI22_X1 U22159 ( .A1(n19214), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19213), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19215) );
  OAI21_X1 U22160 ( .B1(n12845), .B2(n19216), .A(n19215), .ZN(P2_U2951) );
  AOI22_X1 U22161 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19218), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19217), .ZN(n19227) );
  OAI22_X1 U22162 ( .A1(n19222), .A2(n19221), .B1(n19220), .B2(n19219), .ZN(
        n19223) );
  AOI21_X1 U22163 ( .B1(n19225), .B2(n19224), .A(n19223), .ZN(n19226) );
  OAI211_X1 U22164 ( .C1(n19229), .C2(n19228), .A(n19227), .B(n19226), .ZN(
        P2_U3010) );
  AOI22_X2 U22165 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19261), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19260), .ZN(n19690) );
  INV_X1 U22166 ( .A(n19690), .ZN(n19576) );
  NOR2_X2 U22167 ( .A1(n19231), .A2(n19230), .ZN(n19685) );
  AOI22_X1 U22168 ( .A1(n19576), .A2(n19725), .B1(n19258), .B2(n19685), .ZN(
        n19235) );
  NOR2_X2 U22169 ( .A1(n19232), .A2(n19442), .ZN(n19686) );
  AOI22_X1 U22170 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19260), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19261), .ZN(n19233) );
  AOI22_X1 U22171 ( .A1(n19686), .A2(n19262), .B1(n19286), .B2(n19687), .ZN(
        n19234) );
  OAI211_X1 U22172 ( .C1(n19266), .C2(n19236), .A(n19235), .B(n19234), .ZN(
        P2_U3049) );
  INV_X1 U22173 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19239) );
  AOI22_X1 U22174 ( .A1(n19725), .A2(n19539), .B1(n19691), .B2(n19258), .ZN(
        n19238) );
  AOI22_X1 U22175 ( .A1(n13433), .A2(n19262), .B1(n19286), .B2(n19692), .ZN(
        n19237) );
  OAI211_X1 U22176 ( .C1(n19266), .C2(n19239), .A(n19238), .B(n19237), .ZN(
        P2_U3050) );
  AOI22_X1 U22177 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19261), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19260), .ZN(n19701) );
  AOI22_X1 U22178 ( .A1(n19725), .A2(n19579), .B1(n19258), .B2(n19696), .ZN(
        n19242) );
  NOR2_X2 U22179 ( .A1(n19240), .A2(n19442), .ZN(n19697) );
  AOI22_X1 U22180 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19260), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19261), .ZN(n19545) );
  AOI22_X1 U22181 ( .A1(n19697), .A2(n19262), .B1(n19286), .B2(n19698), .ZN(
        n19241) );
  OAI211_X1 U22182 ( .C1(n19266), .C2(n19243), .A(n19242), .B(n19241), .ZN(
        P2_U3051) );
  AOI22_X1 U22183 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n19260), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19261), .ZN(n19707) );
  AOI22_X1 U22184 ( .A1(n19725), .A2(n19647), .B1(n19258), .B2(n19702), .ZN(
        n19247) );
  NOR2_X2 U22185 ( .A1(n19245), .A2(n19442), .ZN(n19703) );
  AOI22_X1 U22186 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19260), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19261), .ZN(n19650) );
  INV_X1 U22187 ( .A(n19650), .ZN(n19704) );
  AOI22_X1 U22188 ( .A1(n19703), .A2(n19262), .B1(n19286), .B2(n19704), .ZN(
        n19246) );
  OAI211_X1 U22189 ( .C1(n19266), .C2(n19248), .A(n19247), .B(n19246), .ZN(
        P2_U3052) );
  AOI22_X1 U22190 ( .A1(n19725), .A2(n19651), .B1(n19708), .B2(n19258), .ZN(
        n19250) );
  AOI22_X1 U22191 ( .A1(n19709), .A2(n19262), .B1(n19286), .B2(n19710), .ZN(
        n19249) );
  OAI211_X1 U22192 ( .C1(n19266), .C2(n21045), .A(n19250), .B(n19249), .ZN(
        P2_U3053) );
  AOI22_X1 U22193 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19261), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19260), .ZN(n19719) );
  INV_X1 U22194 ( .A(n19719), .ZN(n19655) );
  AND2_X1 U22195 ( .A1(n19251), .A2(n19256), .ZN(n19714) );
  AOI22_X1 U22196 ( .A1(n19725), .A2(n19655), .B1(n19258), .B2(n19714), .ZN(
        n19254) );
  NOR2_X2 U22197 ( .A1(n19252), .A2(n19442), .ZN(n19715) );
  AOI22_X1 U22198 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19260), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19261), .ZN(n19658) );
  AOI22_X1 U22199 ( .A1(n19715), .A2(n19262), .B1(n19286), .B2(n19716), .ZN(
        n19253) );
  OAI211_X1 U22200 ( .C1(n19266), .C2(n19255), .A(n19254), .B(n19253), .ZN(
        P2_U3054) );
  AOI22_X1 U22201 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19260), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19261), .ZN(n19730) );
  INV_X1 U22202 ( .A(n19730), .ZN(n19660) );
  AOI22_X1 U22203 ( .A1(n19725), .A2(n19660), .B1(n19258), .B2(n19720), .ZN(
        n19264) );
  NOR2_X2 U22204 ( .A1(n19259), .A2(n19442), .ZN(n19722) );
  AOI22_X1 U22205 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19261), .B1(
        BUF1_REG_23__SCAN_IN), .B2(n19260), .ZN(n19666) );
  AOI22_X1 U22206 ( .A1(n19722), .A2(n19262), .B1(n19286), .B2(n19724), .ZN(
        n19263) );
  OAI211_X1 U22207 ( .C1(n19266), .C2(n19265), .A(n19264), .B(n19263), .ZN(
        P2_U3055) );
  NOR2_X1 U22208 ( .A1(n19496), .A2(n19330), .ZN(n19289) );
  AOI21_X1 U22209 ( .B1(n19593), .B2(n19270), .A(n19437), .ZN(n19268) );
  AOI22_X1 U22210 ( .A1(n19290), .A2(n19672), .B1(n19671), .B2(n19289), .ZN(
        n19275) );
  AND2_X1 U22211 ( .A1(n19269), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19440) );
  OAI21_X1 U22212 ( .B1(n19378), .B2(n19497), .A(n19270), .ZN(n19272) );
  AND2_X1 U22213 ( .A1(n19272), .A2(n19271), .ZN(n19273) );
  OAI211_X1 U22214 ( .C1(n19289), .C2(n19825), .A(n19273), .B(n19679), .ZN(
        n19291) );
  AOI22_X1 U22215 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19291), .B1(
        n19286), .B2(n19604), .ZN(n19274) );
  OAI211_X1 U22216 ( .C1(n19607), .C2(n19321), .A(n19275), .B(n19274), .ZN(
        P2_U3056) );
  AOI22_X1 U22217 ( .A1(n19290), .A2(n19686), .B1(n19685), .B2(n19289), .ZN(
        n19277) );
  AOI22_X1 U22218 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19291), .B1(
        n19324), .B2(n19687), .ZN(n19276) );
  OAI211_X1 U22219 ( .C1(n19690), .C2(n19294), .A(n19277), .B(n19276), .ZN(
        P2_U3057) );
  AOI22_X1 U22220 ( .A1(n19290), .A2(n13433), .B1(n19691), .B2(n19289), .ZN(
        n19279) );
  AOI22_X1 U22221 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19291), .B1(
        n19286), .B2(n19539), .ZN(n19278) );
  OAI211_X1 U22222 ( .C1(n19542), .C2(n19321), .A(n19279), .B(n19278), .ZN(
        P2_U3058) );
  AOI22_X1 U22223 ( .A1(n19290), .A2(n19697), .B1(n19696), .B2(n19289), .ZN(
        n19281) );
  AOI22_X1 U22224 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19291), .B1(
        n19324), .B2(n19698), .ZN(n19280) );
  OAI211_X1 U22225 ( .C1(n19701), .C2(n19294), .A(n19281), .B(n19280), .ZN(
        P2_U3059) );
  AOI22_X1 U22226 ( .A1(n19290), .A2(n19703), .B1(n19702), .B2(n19289), .ZN(
        n19283) );
  AOI22_X1 U22227 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19291), .B1(
        n19324), .B2(n19704), .ZN(n19282) );
  OAI211_X1 U22228 ( .C1(n19707), .C2(n19294), .A(n19283), .B(n19282), .ZN(
        P2_U3060) );
  AOI22_X1 U22229 ( .A1(n19290), .A2(n19709), .B1(n19708), .B2(n19289), .ZN(
        n19285) );
  AOI22_X1 U22230 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19291), .B1(
        n19324), .B2(n19710), .ZN(n19284) );
  OAI211_X1 U22231 ( .C1(n19713), .C2(n19294), .A(n19285), .B(n19284), .ZN(
        P2_U3061) );
  AOI22_X1 U22232 ( .A1(n19290), .A2(n19715), .B1(n19714), .B2(n19289), .ZN(
        n19288) );
  AOI22_X1 U22233 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19291), .B1(
        n19286), .B2(n19655), .ZN(n19287) );
  OAI211_X1 U22234 ( .C1(n19658), .C2(n19321), .A(n19288), .B(n19287), .ZN(
        P2_U3062) );
  AOI22_X1 U22235 ( .A1(n19290), .A2(n19722), .B1(n19720), .B2(n19289), .ZN(
        n19293) );
  AOI22_X1 U22236 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19291), .B1(
        n19324), .B2(n19724), .ZN(n19292) );
  OAI211_X1 U22237 ( .C1(n19730), .C2(n19294), .A(n19293), .B(n19292), .ZN(
        P2_U3063) );
  NOR2_X1 U22238 ( .A1(n19526), .A2(n19330), .ZN(n19322) );
  OAI21_X1 U22239 ( .B1(n19295), .B2(n19322), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19297) );
  INV_X1 U22240 ( .A(n19330), .ZN(n19296) );
  NAND2_X1 U22241 ( .A1(n19525), .A2(n19296), .ZN(n19302) );
  NAND2_X1 U22242 ( .A1(n19297), .A2(n19302), .ZN(n19323) );
  AOI22_X1 U22243 ( .A1(n19323), .A2(n19672), .B1(n19671), .B2(n19322), .ZN(
        n19308) );
  INV_X1 U22244 ( .A(n19322), .ZN(n19298) );
  OAI21_X1 U22245 ( .B1(n19299), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19298), 
        .ZN(n19305) );
  INV_X1 U22246 ( .A(n19407), .ZN(n19301) );
  OAI21_X1 U22247 ( .B1(n19350), .B2(n19324), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19303) );
  NAND2_X1 U22248 ( .A1(n19303), .A2(n19302), .ZN(n19304) );
  MUX2_X1 U22249 ( .A(n19305), .B(n19304), .S(n19830), .Z(n19306) );
  NAND2_X1 U22250 ( .A1(n19306), .A2(n19679), .ZN(n19325) );
  AOI22_X1 U22251 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19325), .B1(
        n19350), .B2(n19681), .ZN(n19307) );
  OAI211_X1 U22252 ( .C1(n19684), .C2(n19321), .A(n19308), .B(n19307), .ZN(
        P2_U3064) );
  AOI22_X1 U22253 ( .A1(n19323), .A2(n19686), .B1(n19685), .B2(n19322), .ZN(
        n19310) );
  AOI22_X1 U22254 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19325), .B1(
        n19350), .B2(n19687), .ZN(n19309) );
  OAI211_X1 U22255 ( .C1(n19690), .C2(n19321), .A(n19310), .B(n19309), .ZN(
        P2_U3065) );
  AOI22_X1 U22256 ( .A1(n19323), .A2(n13433), .B1(n19691), .B2(n19322), .ZN(
        n19312) );
  AOI22_X1 U22257 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19325), .B1(
        n19350), .B2(n19692), .ZN(n19311) );
  OAI211_X1 U22258 ( .C1(n19695), .C2(n19321), .A(n19312), .B(n19311), .ZN(
        P2_U3066) );
  AOI22_X1 U22259 ( .A1(n19323), .A2(n19697), .B1(n19696), .B2(n19322), .ZN(
        n19314) );
  AOI22_X1 U22260 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19325), .B1(
        n19350), .B2(n19698), .ZN(n19313) );
  OAI211_X1 U22261 ( .C1(n19701), .C2(n19321), .A(n19314), .B(n19313), .ZN(
        P2_U3067) );
  AOI22_X1 U22262 ( .A1(n19323), .A2(n19703), .B1(n19702), .B2(n19322), .ZN(
        n19316) );
  AOI22_X1 U22263 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19325), .B1(
        n19324), .B2(n19647), .ZN(n19315) );
  OAI211_X1 U22264 ( .C1(n19650), .C2(n19358), .A(n19316), .B(n19315), .ZN(
        P2_U3068) );
  AOI22_X1 U22265 ( .A1(n19323), .A2(n19709), .B1(n19708), .B2(n19322), .ZN(
        n19318) );
  AOI22_X1 U22266 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19325), .B1(
        n19324), .B2(n19651), .ZN(n19317) );
  OAI211_X1 U22267 ( .C1(n19654), .C2(n19358), .A(n19318), .B(n19317), .ZN(
        P2_U3069) );
  AOI22_X1 U22268 ( .A1(n19323), .A2(n19715), .B1(n19714), .B2(n19322), .ZN(
        n19320) );
  AOI22_X1 U22269 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19325), .B1(
        n19350), .B2(n19716), .ZN(n19319) );
  OAI211_X1 U22270 ( .C1(n19719), .C2(n19321), .A(n19320), .B(n19319), .ZN(
        P2_U3070) );
  AOI22_X1 U22271 ( .A1(n19323), .A2(n19722), .B1(n19720), .B2(n19322), .ZN(
        n19327) );
  AOI22_X1 U22272 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19325), .B1(
        n19324), .B2(n19660), .ZN(n19326) );
  OAI211_X1 U22273 ( .C1(n19666), .C2(n19358), .A(n19327), .B(n19326), .ZN(
        P2_U3071) );
  NOR2_X1 U22274 ( .A1(n19328), .A2(n19330), .ZN(n19353) );
  AOI22_X1 U22275 ( .A1(n19350), .A2(n19604), .B1(n19671), .B2(n19353), .ZN(
        n19339) );
  OAI21_X1 U22276 ( .B1(n19378), .B2(n19329), .A(n19830), .ZN(n19337) );
  NOR2_X1 U22277 ( .A1(n19846), .A2(n19330), .ZN(n19334) );
  OAI21_X1 U22278 ( .B1(n10579), .B2(n19593), .A(n19825), .ZN(n19332) );
  INV_X1 U22279 ( .A(n19353), .ZN(n19331) );
  AOI21_X1 U22280 ( .B1(n19332), .B2(n19331), .A(n19442), .ZN(n19333) );
  OAI21_X1 U22281 ( .B1(n19337), .B2(n19334), .A(n19333), .ZN(n19355) );
  INV_X1 U22282 ( .A(n19334), .ZN(n19336) );
  OAI21_X1 U22283 ( .B1(n10579), .B2(n19353), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19335) );
  OAI21_X1 U22284 ( .B1(n19337), .B2(n19336), .A(n19335), .ZN(n19354) );
  AOI22_X1 U22285 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19355), .B1(
        n19672), .B2(n19354), .ZN(n19338) );
  OAI211_X1 U22286 ( .C1(n19607), .C2(n19365), .A(n19339), .B(n19338), .ZN(
        P2_U3072) );
  AOI22_X1 U22287 ( .A1(n19374), .A2(n19687), .B1(n19353), .B2(n19685), .ZN(
        n19341) );
  AOI22_X1 U22288 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19355), .B1(
        n19686), .B2(n19354), .ZN(n19340) );
  OAI211_X1 U22289 ( .C1(n19690), .C2(n19358), .A(n19341), .B(n19340), .ZN(
        P2_U3073) );
  AOI22_X1 U22290 ( .A1(n19350), .A2(n19539), .B1(n19691), .B2(n19353), .ZN(
        n19343) );
  AOI22_X1 U22291 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19355), .B1(
        n13433), .B2(n19354), .ZN(n19342) );
  OAI211_X1 U22292 ( .C1(n19542), .C2(n19365), .A(n19343), .B(n19342), .ZN(
        P2_U3074) );
  AOI22_X1 U22293 ( .A1(n19350), .A2(n19579), .B1(n19353), .B2(n19696), .ZN(
        n19345) );
  AOI22_X1 U22294 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19355), .B1(
        n19697), .B2(n19354), .ZN(n19344) );
  OAI211_X1 U22295 ( .C1(n19545), .C2(n19365), .A(n19345), .B(n19344), .ZN(
        P2_U3075) );
  AOI22_X1 U22296 ( .A1(n19350), .A2(n19647), .B1(n19353), .B2(n19702), .ZN(
        n19347) );
  AOI22_X1 U22297 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19355), .B1(
        n19703), .B2(n19354), .ZN(n19346) );
  OAI211_X1 U22298 ( .C1(n19650), .C2(n19365), .A(n19347), .B(n19346), .ZN(
        P2_U3076) );
  AOI22_X1 U22299 ( .A1(n19350), .A2(n19651), .B1(n19708), .B2(n19353), .ZN(
        n19349) );
  AOI22_X1 U22300 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19355), .B1(
        n19709), .B2(n19354), .ZN(n19348) );
  OAI211_X1 U22301 ( .C1(n19654), .C2(n19365), .A(n19349), .B(n19348), .ZN(
        P2_U3077) );
  AOI22_X1 U22302 ( .A1(n19350), .A2(n19655), .B1(n19353), .B2(n19714), .ZN(
        n19352) );
  AOI22_X1 U22303 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19355), .B1(
        n19715), .B2(n19354), .ZN(n19351) );
  OAI211_X1 U22304 ( .C1(n19658), .C2(n19365), .A(n19352), .B(n19351), .ZN(
        P2_U3078) );
  AOI22_X1 U22305 ( .A1(n19724), .A2(n19374), .B1(n19353), .B2(n19720), .ZN(
        n19357) );
  AOI22_X1 U22306 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19355), .B1(
        n19722), .B2(n19354), .ZN(n19356) );
  OAI211_X1 U22307 ( .C1(n19730), .C2(n19358), .A(n19357), .B(n19356), .ZN(
        P2_U3079) );
  AOI22_X1 U22308 ( .A1(n19373), .A2(n19686), .B1(n19685), .B2(n19372), .ZN(
        n19360) );
  AOI22_X1 U22309 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19375), .B1(
        n19395), .B2(n19687), .ZN(n19359) );
  OAI211_X1 U22310 ( .C1(n19690), .C2(n19365), .A(n19360), .B(n19359), .ZN(
        P2_U3081) );
  AOI22_X1 U22311 ( .A1(n19373), .A2(n13433), .B1(n19691), .B2(n19372), .ZN(
        n19362) );
  AOI22_X1 U22312 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19375), .B1(
        n19395), .B2(n19692), .ZN(n19361) );
  OAI211_X1 U22313 ( .C1(n19695), .C2(n19365), .A(n19362), .B(n19361), .ZN(
        P2_U3082) );
  AOI22_X1 U22314 ( .A1(n19373), .A2(n19697), .B1(n19696), .B2(n19372), .ZN(
        n19364) );
  AOI22_X1 U22315 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19375), .B1(
        n19395), .B2(n19698), .ZN(n19363) );
  OAI211_X1 U22316 ( .C1(n19701), .C2(n19365), .A(n19364), .B(n19363), .ZN(
        P2_U3083) );
  AOI22_X1 U22317 ( .A1(n19373), .A2(n19703), .B1(n19702), .B2(n19372), .ZN(
        n19367) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19375), .B1(
        n19374), .B2(n19647), .ZN(n19366) );
  OAI211_X1 U22319 ( .C1(n19650), .C2(n19406), .A(n19367), .B(n19366), .ZN(
        P2_U3084) );
  AOI22_X1 U22320 ( .A1(n19373), .A2(n19709), .B1(n19708), .B2(n19372), .ZN(
        n19369) );
  AOI22_X1 U22321 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19375), .B1(
        n19374), .B2(n19651), .ZN(n19368) );
  OAI211_X1 U22322 ( .C1(n19654), .C2(n19406), .A(n19369), .B(n19368), .ZN(
        P2_U3085) );
  AOI22_X1 U22323 ( .A1(n19373), .A2(n19715), .B1(n19714), .B2(n19372), .ZN(
        n19371) );
  AOI22_X1 U22324 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19375), .B1(
        n19374), .B2(n19655), .ZN(n19370) );
  OAI211_X1 U22325 ( .C1(n19658), .C2(n19406), .A(n19371), .B(n19370), .ZN(
        P2_U3086) );
  AOI22_X1 U22326 ( .A1(n19373), .A2(n19722), .B1(n19720), .B2(n19372), .ZN(
        n19377) );
  AOI22_X1 U22327 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19375), .B1(
        n19374), .B2(n19660), .ZN(n19376) );
  OAI211_X1 U22328 ( .C1(n19666), .C2(n19406), .A(n19377), .B(n19376), .ZN(
        P2_U3087) );
  NOR2_X1 U22329 ( .A1(n19855), .A2(n19385), .ZN(n19411) );
  AOI22_X1 U22330 ( .A1(n19604), .A2(n19395), .B1(n19671), .B2(n19411), .ZN(
        n19388) );
  OAI21_X1 U22331 ( .B1(n19378), .B2(n19597), .A(n19830), .ZN(n19386) );
  INV_X1 U22332 ( .A(n19383), .ZN(n19380) );
  INV_X1 U22333 ( .A(n19411), .ZN(n19379) );
  OAI211_X1 U22334 ( .C1(n19380), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19676), 
        .B(n19379), .ZN(n19381) );
  OAI211_X1 U22335 ( .C1(n19386), .C2(n19382), .A(n19679), .B(n19381), .ZN(
        n19403) );
  OAI21_X1 U22336 ( .B1(n19383), .B2(n19411), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19384) );
  OAI21_X1 U22337 ( .B1(n19386), .B2(n19385), .A(n19384), .ZN(n19402) );
  AOI22_X1 U22338 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19403), .B1(
        n19672), .B2(n19402), .ZN(n19387) );
  OAI211_X1 U22339 ( .C1(n19607), .C2(n19434), .A(n19388), .B(n19387), .ZN(
        P2_U3088) );
  AOI22_X1 U22340 ( .A1(n19422), .A2(n19687), .B1(n19685), .B2(n19411), .ZN(
        n19390) );
  AOI22_X1 U22341 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19403), .B1(
        n19686), .B2(n19402), .ZN(n19389) );
  OAI211_X1 U22342 ( .C1(n19690), .C2(n19406), .A(n19390), .B(n19389), .ZN(
        P2_U3089) );
  AOI22_X1 U22343 ( .A1(n19539), .A2(n19395), .B1(n19691), .B2(n19411), .ZN(
        n19392) );
  AOI22_X1 U22344 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19403), .B1(
        n13433), .B2(n19402), .ZN(n19391) );
  OAI211_X1 U22345 ( .C1(n19542), .C2(n19434), .A(n19392), .B(n19391), .ZN(
        P2_U3090) );
  AOI22_X1 U22346 ( .A1(n19579), .A2(n19395), .B1(n19411), .B2(n19696), .ZN(
        n19394) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19403), .B1(
        n19697), .B2(n19402), .ZN(n19393) );
  OAI211_X1 U22348 ( .C1(n19545), .C2(n19434), .A(n19394), .B(n19393), .ZN(
        P2_U3091) );
  AOI22_X1 U22349 ( .A1(n19647), .A2(n19395), .B1(n19411), .B2(n19702), .ZN(
        n19397) );
  AOI22_X1 U22350 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19403), .B1(
        n19703), .B2(n19402), .ZN(n19396) );
  OAI211_X1 U22351 ( .C1(n19650), .C2(n19434), .A(n19397), .B(n19396), .ZN(
        P2_U3092) );
  AOI22_X1 U22352 ( .A1(n19710), .A2(n19422), .B1(n19708), .B2(n19411), .ZN(
        n19399) );
  AOI22_X1 U22353 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19403), .B1(
        n19709), .B2(n19402), .ZN(n19398) );
  OAI211_X1 U22354 ( .C1(n19713), .C2(n19406), .A(n19399), .B(n19398), .ZN(
        P2_U3093) );
  AOI22_X1 U22355 ( .A1(n19716), .A2(n19422), .B1(n19411), .B2(n19714), .ZN(
        n19401) );
  AOI22_X1 U22356 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19403), .B1(
        n19715), .B2(n19402), .ZN(n19400) );
  OAI211_X1 U22357 ( .C1(n19719), .C2(n19406), .A(n19401), .B(n19400), .ZN(
        P2_U3094) );
  AOI22_X1 U22358 ( .A1(n19724), .A2(n19422), .B1(n19720), .B2(n19411), .ZN(
        n19405) );
  AOI22_X1 U22359 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19403), .B1(
        n19722), .B2(n19402), .ZN(n19404) );
  OAI211_X1 U22360 ( .C1(n19730), .C2(n19406), .A(n19405), .B(n19404), .ZN(
        P2_U3095) );
  NAND2_X1 U22361 ( .A1(n19829), .A2(n19667), .ZN(n19438) );
  NOR2_X1 U22362 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19438), .ZN(
        n19429) );
  NOR2_X1 U22363 ( .A1(n19411), .A2(n19429), .ZN(n19408) );
  OR2_X1 U22364 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19408), .ZN(n19409) );
  NOR3_X1 U22365 ( .A1(n10580), .A2(n19429), .A3(n19593), .ZN(n19412) );
  AOI21_X1 U22366 ( .B1(n19593), .B2(n19409), .A(n19412), .ZN(n19430) );
  AOI22_X1 U22367 ( .A1(n19430), .A2(n19672), .B1(n19671), .B2(n19429), .ZN(
        n19415) );
  AOI21_X1 U22368 ( .B1(n19434), .B2(n19464), .A(n19818), .ZN(n19410) );
  AOI221_X1 U22369 ( .B1(n19825), .B2(n19411), .C1(n19825), .C2(n19410), .A(
        n19429), .ZN(n19413) );
  AOI22_X1 U22370 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19431), .B1(
        n19422), .B2(n19604), .ZN(n19414) );
  OAI211_X1 U22371 ( .C1(n19607), .C2(n19464), .A(n19415), .B(n19414), .ZN(
        P2_U3096) );
  AOI22_X1 U22372 ( .A1(n19430), .A2(n19686), .B1(n19685), .B2(n19429), .ZN(
        n19417) );
  AOI22_X1 U22373 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19431), .B1(
        n19457), .B2(n19687), .ZN(n19416) );
  OAI211_X1 U22374 ( .C1(n19690), .C2(n19434), .A(n19417), .B(n19416), .ZN(
        P2_U3097) );
  AOI22_X1 U22375 ( .A1(n19430), .A2(n13433), .B1(n19691), .B2(n19429), .ZN(
        n19419) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19431), .B1(
        n19457), .B2(n19692), .ZN(n19418) );
  OAI211_X1 U22377 ( .C1(n19695), .C2(n19434), .A(n19419), .B(n19418), .ZN(
        P2_U3098) );
  AOI22_X1 U22378 ( .A1(n19430), .A2(n19697), .B1(n19696), .B2(n19429), .ZN(
        n19421) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19431), .B1(
        n19422), .B2(n19579), .ZN(n19420) );
  OAI211_X1 U22380 ( .C1(n19545), .C2(n19464), .A(n19421), .B(n19420), .ZN(
        P2_U3099) );
  AOI22_X1 U22381 ( .A1(n19430), .A2(n19703), .B1(n19702), .B2(n19429), .ZN(
        n19424) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19431), .B1(
        n19422), .B2(n19647), .ZN(n19423) );
  OAI211_X1 U22383 ( .C1(n19650), .C2(n19464), .A(n19424), .B(n19423), .ZN(
        P2_U3100) );
  AOI22_X1 U22384 ( .A1(n19430), .A2(n19709), .B1(n19708), .B2(n19429), .ZN(
        n19426) );
  AOI22_X1 U22385 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19431), .B1(
        n19457), .B2(n19710), .ZN(n19425) );
  OAI211_X1 U22386 ( .C1(n19713), .C2(n19434), .A(n19426), .B(n19425), .ZN(
        P2_U3101) );
  AOI22_X1 U22387 ( .A1(n19430), .A2(n19715), .B1(n19714), .B2(n19429), .ZN(
        n19428) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19431), .B1(
        n19457), .B2(n19716), .ZN(n19427) );
  OAI211_X1 U22389 ( .C1(n19719), .C2(n19434), .A(n19428), .B(n19427), .ZN(
        P2_U3102) );
  AOI22_X1 U22390 ( .A1(n19430), .A2(n19722), .B1(n19720), .B2(n19429), .ZN(
        n19433) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19431), .B1(
        n19457), .B2(n19724), .ZN(n19432) );
  OAI211_X1 U22392 ( .C1(n19730), .C2(n19434), .A(n19433), .B(n19432), .ZN(
        P2_U3103) );
  INV_X1 U22393 ( .A(n19435), .ZN(n19436) );
  INV_X1 U22394 ( .A(n19819), .ZN(n19439) );
  NOR2_X1 U22395 ( .A1(n19855), .A2(n19438), .ZN(n19471) );
  NOR3_X1 U22396 ( .A1(n10416), .A2(n19471), .A3(n19593), .ZN(n19441) );
  AOI211_X2 U22397 ( .C1(n19438), .C2(n19593), .A(n19437), .B(n19441), .ZN(
        n19460) );
  AOI22_X1 U22398 ( .A1(n19460), .A2(n19672), .B1(n19671), .B2(n19471), .ZN(
        n19446) );
  INV_X1 U22399 ( .A(n19438), .ZN(n19444) );
  AND2_X1 U22400 ( .A1(n19440), .A2(n19439), .ZN(n19817) );
  INV_X1 U22401 ( .A(n19471), .ZN(n19468) );
  AOI211_X1 U22402 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19468), .A(n19442), 
        .B(n19441), .ZN(n19443) );
  OAI21_X1 U22403 ( .B1(n19444), .B2(n19817), .A(n19443), .ZN(n19461) );
  AOI22_X1 U22404 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19461), .B1(
        n19457), .B2(n19604), .ZN(n19445) );
  OAI211_X1 U22405 ( .C1(n19607), .C2(n19489), .A(n19446), .B(n19445), .ZN(
        P2_U3104) );
  AOI22_X1 U22406 ( .A1(n19460), .A2(n19686), .B1(n19685), .B2(n19471), .ZN(
        n19448) );
  AOI22_X1 U22407 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19461), .B1(
        n19491), .B2(n19687), .ZN(n19447) );
  OAI211_X1 U22408 ( .C1(n19690), .C2(n19464), .A(n19448), .B(n19447), .ZN(
        P2_U3105) );
  AOI22_X1 U22409 ( .A1(n19460), .A2(n13433), .B1(n19691), .B2(n19471), .ZN(
        n19450) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19461), .B1(
        n19457), .B2(n19539), .ZN(n19449) );
  OAI211_X1 U22411 ( .C1(n19542), .C2(n19489), .A(n19450), .B(n19449), .ZN(
        P2_U3106) );
  AOI22_X1 U22412 ( .A1(n19460), .A2(n19697), .B1(n19696), .B2(n19471), .ZN(
        n19452) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19461), .B1(
        n19457), .B2(n19579), .ZN(n19451) );
  OAI211_X1 U22414 ( .C1(n19545), .C2(n19489), .A(n19452), .B(n19451), .ZN(
        P2_U3107) );
  AOI22_X1 U22415 ( .A1(n19460), .A2(n19703), .B1(n19702), .B2(n19471), .ZN(
        n19454) );
  AOI22_X1 U22416 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19461), .B1(
        n19457), .B2(n19647), .ZN(n19453) );
  OAI211_X1 U22417 ( .C1(n19650), .C2(n19489), .A(n19454), .B(n19453), .ZN(
        P2_U3108) );
  AOI22_X1 U22418 ( .A1(n19460), .A2(n19709), .B1(n19708), .B2(n19471), .ZN(
        n19456) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19461), .B1(
        n19457), .B2(n19651), .ZN(n19455) );
  OAI211_X1 U22420 ( .C1(n19654), .C2(n19489), .A(n19456), .B(n19455), .ZN(
        P2_U3109) );
  AOI22_X1 U22421 ( .A1(n19460), .A2(n19715), .B1(n19714), .B2(n19471), .ZN(
        n19459) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19461), .B1(
        n19457), .B2(n19655), .ZN(n19458) );
  OAI211_X1 U22423 ( .C1(n19658), .C2(n19489), .A(n19459), .B(n19458), .ZN(
        P2_U3110) );
  AOI22_X1 U22424 ( .A1(n19460), .A2(n19722), .B1(n19720), .B2(n19471), .ZN(
        n19463) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19461), .B1(
        n19491), .B2(n19724), .ZN(n19462) );
  OAI211_X1 U22426 ( .C1(n19730), .C2(n19464), .A(n19463), .B(n19462), .ZN(
        P2_U3111) );
  NOR2_X1 U22427 ( .A1(n19529), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19500) );
  INV_X1 U22428 ( .A(n19500), .ZN(n19503) );
  NOR2_X1 U22429 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19503), .ZN(
        n19490) );
  AOI22_X1 U22430 ( .A1(n19520), .A2(n19681), .B1(n19671), .B2(n19490), .ZN(
        n19476) );
  AOI21_X1 U22431 ( .B1(n19515), .B2(n19489), .A(n19818), .ZN(n19465) );
  NOR2_X1 U22432 ( .A1(n19465), .A2(n19676), .ZN(n19470) );
  INV_X1 U22433 ( .A(n19466), .ZN(n19472) );
  OAI21_X1 U22434 ( .B1(n19472), .B2(n19593), .A(n19825), .ZN(n19467) );
  AOI21_X1 U22435 ( .B1(n19470), .B2(n19468), .A(n19467), .ZN(n19469) );
  OAI21_X1 U22436 ( .B1(n19490), .B2(n19469), .A(n19679), .ZN(n19493) );
  OAI21_X1 U22437 ( .B1(n19490), .B2(n19471), .A(n19470), .ZN(n19474) );
  OAI21_X1 U22438 ( .B1(n19472), .B2(n19490), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19473) );
  AOI22_X1 U22439 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19493), .B1(
        n19672), .B2(n19492), .ZN(n19475) );
  OAI211_X1 U22440 ( .C1(n19684), .C2(n19489), .A(n19476), .B(n19475), .ZN(
        P2_U3112) );
  AOI22_X1 U22441 ( .A1(n19520), .A2(n19687), .B1(n19685), .B2(n19490), .ZN(
        n19478) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19493), .B1(
        n19492), .B2(n19686), .ZN(n19477) );
  OAI211_X1 U22443 ( .C1(n19690), .C2(n19489), .A(n19478), .B(n19477), .ZN(
        P2_U3113) );
  AOI22_X1 U22444 ( .A1(n19491), .A2(n19539), .B1(n19691), .B2(n19490), .ZN(
        n19480) );
  AOI22_X1 U22445 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19493), .B1(
        n19492), .B2(n13433), .ZN(n19479) );
  OAI211_X1 U22446 ( .C1(n19542), .C2(n19515), .A(n19480), .B(n19479), .ZN(
        P2_U3114) );
  AOI22_X1 U22447 ( .A1(n19491), .A2(n19579), .B1(n19696), .B2(n19490), .ZN(
        n19482) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19493), .B1(
        n19492), .B2(n19697), .ZN(n19481) );
  OAI211_X1 U22449 ( .C1(n19545), .C2(n19515), .A(n19482), .B(n19481), .ZN(
        P2_U3115) );
  AOI22_X1 U22450 ( .A1(n19491), .A2(n19647), .B1(n19702), .B2(n19490), .ZN(
        n19484) );
  AOI22_X1 U22451 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19493), .B1(
        n19492), .B2(n19703), .ZN(n19483) );
  OAI211_X1 U22452 ( .C1(n19650), .C2(n19515), .A(n19484), .B(n19483), .ZN(
        P2_U3116) );
  AOI22_X1 U22453 ( .A1(n19520), .A2(n19710), .B1(n19708), .B2(n19490), .ZN(
        n19486) );
  AOI22_X1 U22454 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19493), .B1(
        n19492), .B2(n19709), .ZN(n19485) );
  OAI211_X1 U22455 ( .C1(n19713), .C2(n19489), .A(n19486), .B(n19485), .ZN(
        P2_U3117) );
  AOI22_X1 U22456 ( .A1(n19520), .A2(n19716), .B1(n19714), .B2(n19490), .ZN(
        n19488) );
  AOI22_X1 U22457 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19493), .B1(
        n19492), .B2(n19715), .ZN(n19487) );
  OAI211_X1 U22458 ( .C1(n19719), .C2(n19489), .A(n19488), .B(n19487), .ZN(
        P2_U3118) );
  AOI22_X1 U22459 ( .A1(n19491), .A2(n19660), .B1(n19720), .B2(n19490), .ZN(
        n19495) );
  AOI22_X1 U22460 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19493), .B1(
        n19492), .B2(n19722), .ZN(n19494) );
  OAI211_X1 U22461 ( .C1(n19666), .C2(n19515), .A(n19495), .B(n19494), .ZN(
        P2_U3119) );
  NOR2_X1 U22462 ( .A1(n19496), .A2(n19529), .ZN(n19531) );
  AOI22_X1 U22463 ( .A1(n19555), .A2(n19681), .B1(n19671), .B2(n19531), .ZN(
        n19506) );
  INV_X1 U22464 ( .A(n19599), .ZN(n19674) );
  OAI21_X1 U22465 ( .B1(n19674), .B2(n19497), .A(n19830), .ZN(n19504) );
  INV_X1 U22466 ( .A(n19531), .ZN(n19498) );
  OAI211_X1 U22467 ( .C1(n10571), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19676), 
        .B(n19498), .ZN(n19499) );
  OAI211_X1 U22468 ( .C1(n19504), .C2(n19500), .A(n19679), .B(n19499), .ZN(
        n19522) );
  OAI21_X1 U22469 ( .B1(n19501), .B2(n19531), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19502) );
  OAI21_X1 U22470 ( .B1(n19504), .B2(n19503), .A(n19502), .ZN(n19521) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19522), .B1(
        n19672), .B2(n19521), .ZN(n19505) );
  OAI211_X1 U22472 ( .C1(n19684), .C2(n19515), .A(n19506), .B(n19505), .ZN(
        P2_U3120) );
  AOI22_X1 U22473 ( .A1(n19555), .A2(n19687), .B1(n19685), .B2(n19531), .ZN(
        n19508) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19522), .B1(
        n19686), .B2(n19521), .ZN(n19507) );
  OAI211_X1 U22475 ( .C1(n19690), .C2(n19515), .A(n19508), .B(n19507), .ZN(
        P2_U3121) );
  AOI22_X1 U22476 ( .A1(n19555), .A2(n19692), .B1(n19691), .B2(n19531), .ZN(
        n19510) );
  AOI22_X1 U22477 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19522), .B1(
        n13433), .B2(n19521), .ZN(n19509) );
  OAI211_X1 U22478 ( .C1(n19695), .C2(n19515), .A(n19510), .B(n19509), .ZN(
        P2_U3122) );
  AOI22_X1 U22479 ( .A1(n19520), .A2(n19579), .B1(n19696), .B2(n19531), .ZN(
        n19512) );
  AOI22_X1 U22480 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19522), .B1(
        n19697), .B2(n19521), .ZN(n19511) );
  OAI211_X1 U22481 ( .C1(n19545), .C2(n19552), .A(n19512), .B(n19511), .ZN(
        P2_U3123) );
  AOI22_X1 U22482 ( .A1(n19704), .A2(n19555), .B1(n19702), .B2(n19531), .ZN(
        n19514) );
  AOI22_X1 U22483 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19522), .B1(
        n19703), .B2(n19521), .ZN(n19513) );
  OAI211_X1 U22484 ( .C1(n19707), .C2(n19515), .A(n19514), .B(n19513), .ZN(
        P2_U3124) );
  AOI22_X1 U22485 ( .A1(n19520), .A2(n19651), .B1(n19708), .B2(n19531), .ZN(
        n19517) );
  AOI22_X1 U22486 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19522), .B1(
        n19709), .B2(n19521), .ZN(n19516) );
  OAI211_X1 U22487 ( .C1(n19654), .C2(n19552), .A(n19517), .B(n19516), .ZN(
        P2_U3125) );
  AOI22_X1 U22488 ( .A1(n19520), .A2(n19655), .B1(n19714), .B2(n19531), .ZN(
        n19519) );
  AOI22_X1 U22489 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19522), .B1(
        n19715), .B2(n19521), .ZN(n19518) );
  OAI211_X1 U22490 ( .C1(n19658), .C2(n19552), .A(n19519), .B(n19518), .ZN(
        P2_U3126) );
  AOI22_X1 U22491 ( .A1(n19520), .A2(n19660), .B1(n19720), .B2(n19531), .ZN(
        n19524) );
  AOI22_X1 U22492 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19522), .B1(
        n19722), .B2(n19521), .ZN(n19523) );
  OAI211_X1 U22493 ( .C1(n19666), .C2(n19552), .A(n19524), .B(n19523), .ZN(
        P2_U3127) );
  INV_X1 U22494 ( .A(n19525), .ZN(n19528) );
  NOR2_X1 U22495 ( .A1(n19526), .A2(n19529), .ZN(n19553) );
  OAI21_X1 U22496 ( .B1(n19530), .B2(n19553), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19527) );
  OAI21_X1 U22497 ( .B1(n19529), .B2(n19528), .A(n19527), .ZN(n19554) );
  AOI22_X1 U22498 ( .A1(n19554), .A2(n19672), .B1(n19671), .B2(n19553), .ZN(
        n19536) );
  INV_X1 U22499 ( .A(n19530), .ZN(n19533) );
  AOI221_X1 U22500 ( .B1(n19555), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19559), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19531), .ZN(n19532) );
  AOI211_X1 U22501 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19533), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19532), .ZN(n19534) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19556), .B1(
        n19559), .B2(n19681), .ZN(n19535) );
  OAI211_X1 U22503 ( .C1(n19684), .C2(n19552), .A(n19536), .B(n19535), .ZN(
        P2_U3128) );
  AOI22_X1 U22504 ( .A1(n19554), .A2(n19686), .B1(n19685), .B2(n19553), .ZN(
        n19538) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19556), .B1(
        n19559), .B2(n19687), .ZN(n19537) );
  OAI211_X1 U22506 ( .C1(n19690), .C2(n19552), .A(n19538), .B(n19537), .ZN(
        P2_U3129) );
  AOI22_X1 U22507 ( .A1(n19554), .A2(n13433), .B1(n19691), .B2(n19553), .ZN(
        n19541) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19556), .B1(
        n19555), .B2(n19539), .ZN(n19540) );
  OAI211_X1 U22509 ( .C1(n19542), .C2(n19575), .A(n19541), .B(n19540), .ZN(
        P2_U3130) );
  AOI22_X1 U22510 ( .A1(n19554), .A2(n19697), .B1(n19696), .B2(n19553), .ZN(
        n19544) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19556), .B1(
        n19555), .B2(n19579), .ZN(n19543) );
  OAI211_X1 U22512 ( .C1(n19545), .C2(n19575), .A(n19544), .B(n19543), .ZN(
        P2_U3131) );
  AOI22_X1 U22513 ( .A1(n19554), .A2(n19703), .B1(n19702), .B2(n19553), .ZN(
        n19547) );
  AOI22_X1 U22514 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19556), .B1(
        n19555), .B2(n19647), .ZN(n19546) );
  OAI211_X1 U22515 ( .C1(n19650), .C2(n19575), .A(n19547), .B(n19546), .ZN(
        P2_U3132) );
  AOI22_X1 U22516 ( .A1(n19554), .A2(n19709), .B1(n19708), .B2(n19553), .ZN(
        n19549) );
  AOI22_X1 U22517 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19556), .B1(
        n19559), .B2(n19710), .ZN(n19548) );
  OAI211_X1 U22518 ( .C1(n19713), .C2(n19552), .A(n19549), .B(n19548), .ZN(
        P2_U3133) );
  AOI22_X1 U22519 ( .A1(n19554), .A2(n19715), .B1(n19714), .B2(n19553), .ZN(
        n19551) );
  AOI22_X1 U22520 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19556), .B1(
        n19559), .B2(n19716), .ZN(n19550) );
  OAI211_X1 U22521 ( .C1(n19719), .C2(n19552), .A(n19551), .B(n19550), .ZN(
        P2_U3134) );
  AOI22_X1 U22522 ( .A1(n19554), .A2(n19722), .B1(n19720), .B2(n19553), .ZN(
        n19558) );
  AOI22_X1 U22523 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19556), .B1(
        n19555), .B2(n19660), .ZN(n19557) );
  OAI211_X1 U22524 ( .C1(n19666), .C2(n19575), .A(n19558), .B(n19557), .ZN(
        P2_U3135) );
  AOI22_X1 U22525 ( .A1(n19571), .A2(n19686), .B1(n19570), .B2(n19685), .ZN(
        n19561) );
  AOI22_X1 U22526 ( .A1(n19588), .A2(n19687), .B1(n19559), .B2(n19576), .ZN(
        n19560) );
  OAI211_X1 U22527 ( .C1(n19563), .C2(n19562), .A(n19561), .B(n19560), .ZN(
        P2_U3137) );
  AOI22_X1 U22528 ( .A1(n19571), .A2(n19697), .B1(n19570), .B2(n19696), .ZN(
        n19565) );
  INV_X1 U22529 ( .A(n19563), .ZN(n19572) );
  AOI22_X1 U22530 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19572), .B1(
        n19588), .B2(n19698), .ZN(n19564) );
  OAI211_X1 U22531 ( .C1(n19701), .C2(n19575), .A(n19565), .B(n19564), .ZN(
        P2_U3139) );
  AOI22_X1 U22532 ( .A1(n19571), .A2(n19703), .B1(n19570), .B2(n19702), .ZN(
        n19567) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19572), .B1(
        n19588), .B2(n19704), .ZN(n19566) );
  OAI211_X1 U22534 ( .C1(n19707), .C2(n19575), .A(n19567), .B(n19566), .ZN(
        P2_U3140) );
  AOI22_X1 U22535 ( .A1(n19571), .A2(n19715), .B1(n19570), .B2(n19714), .ZN(
        n19569) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19572), .B1(
        n19588), .B2(n19716), .ZN(n19568) );
  OAI211_X1 U22537 ( .C1(n19719), .C2(n19575), .A(n19569), .B(n19568), .ZN(
        P2_U3142) );
  AOI22_X1 U22538 ( .A1(n19571), .A2(n19722), .B1(n19570), .B2(n19720), .ZN(
        n19574) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19572), .B1(
        n19588), .B2(n19724), .ZN(n19573) );
  OAI211_X1 U22540 ( .C1(n19730), .C2(n19575), .A(n19574), .B(n19573), .ZN(
        P2_U3143) );
  AOI22_X1 U22541 ( .A1(n19587), .A2(n19686), .B1(n19586), .B2(n19685), .ZN(
        n19578) );
  AOI22_X1 U22542 ( .A1(n19614), .A2(n19687), .B1(n19588), .B2(n19576), .ZN(
        n19577) );
  OAI211_X1 U22543 ( .C1(n19591), .C2(n13828), .A(n19578), .B(n19577), .ZN(
        P2_U3145) );
  AOI22_X1 U22544 ( .A1(n19587), .A2(n19697), .B1(n19586), .B2(n19696), .ZN(
        n19581) );
  AOI22_X1 U22545 ( .A1(n19588), .A2(n19579), .B1(n19614), .B2(n19698), .ZN(
        n19580) );
  OAI211_X1 U22546 ( .C1(n19591), .C2(n14037), .A(n19581), .B(n19580), .ZN(
        P2_U3147) );
  AOI22_X1 U22547 ( .A1(n19587), .A2(n19703), .B1(n19586), .B2(n19702), .ZN(
        n19583) );
  AOI22_X1 U22548 ( .A1(n19588), .A2(n19647), .B1(n19614), .B2(n19704), .ZN(
        n19582) );
  OAI211_X1 U22549 ( .C1(n19591), .C2(n14695), .A(n19583), .B(n19582), .ZN(
        P2_U3148) );
  AOI22_X1 U22550 ( .A1(n19587), .A2(n19715), .B1(n19586), .B2(n19714), .ZN(
        n19585) );
  AOI22_X1 U22551 ( .A1(n19614), .A2(n19716), .B1(n19588), .B2(n19655), .ZN(
        n19584) );
  OAI211_X1 U22552 ( .C1(n19591), .C2(n14737), .A(n19585), .B(n19584), .ZN(
        P2_U3150) );
  AOI22_X1 U22553 ( .A1(n19587), .A2(n19722), .B1(n19586), .B2(n19720), .ZN(
        n19590) );
  AOI22_X1 U22554 ( .A1(n19588), .A2(n19660), .B1(n19614), .B2(n19724), .ZN(
        n19589) );
  OAI211_X1 U22555 ( .C1(n19591), .C2(n11257), .A(n19590), .B(n19589), .ZN(
        P2_U3151) );
  INV_X1 U22556 ( .A(n10417), .ZN(n19594) );
  NOR2_X1 U22557 ( .A1(n19855), .A2(n19601), .ZN(n19628) );
  NOR3_X1 U22558 ( .A1(n19594), .A2(n19628), .A3(n19593), .ZN(n19600) );
  INV_X1 U22559 ( .A(n19601), .ZN(n19595) );
  AOI21_X1 U22560 ( .B1(n19825), .B2(n19595), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19596) );
  NOR2_X1 U22561 ( .A1(n19600), .A2(n19596), .ZN(n19621) );
  AOI22_X1 U22562 ( .A1(n19621), .A2(n19672), .B1(n19671), .B2(n19628), .ZN(
        n19606) );
  INV_X1 U22563 ( .A(n19597), .ZN(n19598) );
  NAND2_X1 U22564 ( .A1(n19599), .A2(n19598), .ZN(n19602) );
  AOI21_X1 U22565 ( .B1(n19602), .B2(n19601), .A(n19600), .ZN(n19603) );
  OAI211_X1 U22566 ( .C1(n19628), .C2(n19825), .A(n19603), .B(n19679), .ZN(
        n19622) );
  AOI22_X1 U22567 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19622), .B1(
        n19614), .B2(n19604), .ZN(n19605) );
  OAI211_X1 U22568 ( .C1(n19607), .C2(n19646), .A(n19606), .B(n19605), .ZN(
        P2_U3152) );
  AOI22_X1 U22569 ( .A1(n19621), .A2(n19686), .B1(n19685), .B2(n19628), .ZN(
        n19609) );
  AOI22_X1 U22570 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19622), .B1(
        n19661), .B2(n19687), .ZN(n19608) );
  OAI211_X1 U22571 ( .C1(n19690), .C2(n19625), .A(n19609), .B(n19608), .ZN(
        P2_U3153) );
  AOI22_X1 U22572 ( .A1(n19621), .A2(n13433), .B1(n19691), .B2(n19628), .ZN(
        n19611) );
  AOI22_X1 U22573 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19622), .B1(
        n19661), .B2(n19692), .ZN(n19610) );
  OAI211_X1 U22574 ( .C1(n19695), .C2(n19625), .A(n19611), .B(n19610), .ZN(
        P2_U3154) );
  AOI22_X1 U22575 ( .A1(n19621), .A2(n19697), .B1(n19696), .B2(n19628), .ZN(
        n19613) );
  AOI22_X1 U22576 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19622), .B1(
        n19661), .B2(n19698), .ZN(n19612) );
  OAI211_X1 U22577 ( .C1(n19701), .C2(n19625), .A(n19613), .B(n19612), .ZN(
        P2_U3155) );
  AOI22_X1 U22578 ( .A1(n19621), .A2(n19703), .B1(n19702), .B2(n19628), .ZN(
        n19616) );
  AOI22_X1 U22579 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19622), .B1(
        n19614), .B2(n19647), .ZN(n19615) );
  OAI211_X1 U22580 ( .C1(n19650), .C2(n19646), .A(n19616), .B(n19615), .ZN(
        P2_U3156) );
  AOI22_X1 U22581 ( .A1(n19621), .A2(n19709), .B1(n19708), .B2(n19628), .ZN(
        n19618) );
  AOI22_X1 U22582 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19622), .B1(
        n19661), .B2(n19710), .ZN(n19617) );
  OAI211_X1 U22583 ( .C1(n19713), .C2(n19625), .A(n19618), .B(n19617), .ZN(
        P2_U3157) );
  AOI22_X1 U22584 ( .A1(n19621), .A2(n19715), .B1(n19714), .B2(n19628), .ZN(
        n19620) );
  AOI22_X1 U22585 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19622), .B1(
        n19661), .B2(n19716), .ZN(n19619) );
  OAI211_X1 U22586 ( .C1(n19719), .C2(n19625), .A(n19620), .B(n19619), .ZN(
        P2_U3158) );
  AOI22_X1 U22587 ( .A1(n19621), .A2(n19722), .B1(n19720), .B2(n19628), .ZN(
        n19624) );
  AOI22_X1 U22588 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19622), .B1(
        n19661), .B2(n19724), .ZN(n19623) );
  OAI211_X1 U22589 ( .C1(n19730), .C2(n19625), .A(n19624), .B(n19623), .ZN(
        P2_U3159) );
  INV_X1 U22590 ( .A(n19667), .ZN(n19673) );
  NOR3_X2 U22591 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19829), .A3(
        n19673), .ZN(n19659) );
  AOI22_X1 U22592 ( .A1(n19643), .A2(n19681), .B1(n19671), .B2(n19659), .ZN(
        n19638) );
  OAI21_X1 U22593 ( .B1(n19661), .B2(n19643), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19627) );
  NAND2_X1 U22594 ( .A1(n19627), .A2(n19830), .ZN(n19636) );
  NOR2_X1 U22595 ( .A1(n19659), .A2(n19628), .ZN(n19635) );
  INV_X1 U22596 ( .A(n19635), .ZN(n19632) );
  INV_X1 U22597 ( .A(n19633), .ZN(n19630) );
  INV_X1 U22598 ( .A(n19659), .ZN(n19629) );
  OAI211_X1 U22599 ( .C1(n19630), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19676), 
        .B(n19629), .ZN(n19631) );
  OAI211_X1 U22600 ( .C1(n19636), .C2(n19632), .A(n19679), .B(n19631), .ZN(
        n19663) );
  OAI21_X1 U22601 ( .B1(n19633), .B2(n19659), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19634) );
  AOI22_X1 U22602 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19663), .B1(
        n19672), .B2(n19662), .ZN(n19637) );
  OAI211_X1 U22603 ( .C1(n19684), .C2(n19646), .A(n19638), .B(n19637), .ZN(
        P2_U3160) );
  AOI22_X1 U22604 ( .A1(n19643), .A2(n19687), .B1(n19685), .B2(n19659), .ZN(
        n19640) );
  AOI22_X1 U22605 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19663), .B1(
        n19686), .B2(n19662), .ZN(n19639) );
  OAI211_X1 U22606 ( .C1(n19690), .C2(n19646), .A(n19640), .B(n19639), .ZN(
        P2_U3161) );
  AOI22_X1 U22607 ( .A1(n19643), .A2(n19692), .B1(n19691), .B2(n19659), .ZN(
        n19642) );
  AOI22_X1 U22608 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19663), .B1(
        n13433), .B2(n19662), .ZN(n19641) );
  OAI211_X1 U22609 ( .C1(n19695), .C2(n19646), .A(n19642), .B(n19641), .ZN(
        P2_U3162) );
  AOI22_X1 U22610 ( .A1(n19643), .A2(n19698), .B1(n19696), .B2(n19659), .ZN(
        n19645) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19663), .B1(
        n19697), .B2(n19662), .ZN(n19644) );
  OAI211_X1 U22612 ( .C1(n19701), .C2(n19646), .A(n19645), .B(n19644), .ZN(
        P2_U3163) );
  AOI22_X1 U22613 ( .A1(n19661), .A2(n19647), .B1(n19702), .B2(n19659), .ZN(
        n19649) );
  AOI22_X1 U22614 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19663), .B1(
        n19703), .B2(n19662), .ZN(n19648) );
  OAI211_X1 U22615 ( .C1(n19650), .C2(n19729), .A(n19649), .B(n19648), .ZN(
        P2_U3164) );
  AOI22_X1 U22616 ( .A1(n19661), .A2(n19651), .B1(n19708), .B2(n19659), .ZN(
        n19653) );
  AOI22_X1 U22617 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19663), .B1(
        n19709), .B2(n19662), .ZN(n19652) );
  OAI211_X1 U22618 ( .C1(n19654), .C2(n19729), .A(n19653), .B(n19652), .ZN(
        P2_U3165) );
  AOI22_X1 U22619 ( .A1(n19661), .A2(n19655), .B1(n19714), .B2(n19659), .ZN(
        n19657) );
  AOI22_X1 U22620 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19663), .B1(
        n19715), .B2(n19662), .ZN(n19656) );
  OAI211_X1 U22621 ( .C1(n19658), .C2(n19729), .A(n19657), .B(n19656), .ZN(
        P2_U3166) );
  AOI22_X1 U22622 ( .A1(n19661), .A2(n19660), .B1(n19720), .B2(n19659), .ZN(
        n19665) );
  AOI22_X1 U22623 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19663), .B1(
        n19722), .B2(n19662), .ZN(n19664) );
  OAI211_X1 U22624 ( .C1(n19666), .C2(n19729), .A(n19665), .B(n19664), .ZN(
        P2_U3167) );
  NAND2_X1 U22625 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19667), .ZN(
        n19670) );
  INV_X1 U22626 ( .A(n19677), .ZN(n19668) );
  INV_X1 U22627 ( .A(n19675), .ZN(n19721) );
  OAI21_X1 U22628 ( .B1(n19668), .B2(n19721), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19669) );
  OAI21_X1 U22629 ( .B1(n19670), .B2(n19676), .A(n19669), .ZN(n19723) );
  AOI22_X1 U22630 ( .A1(n19723), .A2(n19672), .B1(n19721), .B2(n19671), .ZN(
        n19683) );
  OAI22_X1 U22631 ( .A1(n19674), .A2(n19819), .B1(n19829), .B2(n19673), .ZN(
        n19680) );
  OAI211_X1 U22632 ( .C1(n19677), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19676), 
        .B(n19675), .ZN(n19678) );
  NAND3_X1 U22633 ( .A1(n19680), .A2(n19679), .A3(n19678), .ZN(n19726) );
  AOI22_X1 U22634 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19726), .B1(
        n19725), .B2(n19681), .ZN(n19682) );
  OAI211_X1 U22635 ( .C1(n19684), .C2(n19729), .A(n19683), .B(n19682), .ZN(
        P2_U3168) );
  AOI22_X1 U22636 ( .A1(n19723), .A2(n19686), .B1(n19721), .B2(n19685), .ZN(
        n19689) );
  AOI22_X1 U22637 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19726), .B1(
        n19725), .B2(n19687), .ZN(n19688) );
  OAI211_X1 U22638 ( .C1(n19690), .C2(n19729), .A(n19689), .B(n19688), .ZN(
        P2_U3169) );
  AOI22_X1 U22639 ( .A1(n19723), .A2(n13433), .B1(n19721), .B2(n19691), .ZN(
        n19694) );
  AOI22_X1 U22640 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19726), .B1(
        n19725), .B2(n19692), .ZN(n19693) );
  OAI211_X1 U22641 ( .C1(n19695), .C2(n19729), .A(n19694), .B(n19693), .ZN(
        P2_U3170) );
  AOI22_X1 U22642 ( .A1(n19723), .A2(n19697), .B1(n19721), .B2(n19696), .ZN(
        n19700) );
  AOI22_X1 U22643 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19726), .B1(
        n19725), .B2(n19698), .ZN(n19699) );
  OAI211_X1 U22644 ( .C1(n19701), .C2(n19729), .A(n19700), .B(n19699), .ZN(
        P2_U3171) );
  AOI22_X1 U22645 ( .A1(n19723), .A2(n19703), .B1(n19721), .B2(n19702), .ZN(
        n19706) );
  AOI22_X1 U22646 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19726), .B1(
        n19725), .B2(n19704), .ZN(n19705) );
  OAI211_X1 U22647 ( .C1(n19707), .C2(n19729), .A(n19706), .B(n19705), .ZN(
        P2_U3172) );
  AOI22_X1 U22648 ( .A1(n19723), .A2(n19709), .B1(n19721), .B2(n19708), .ZN(
        n19712) );
  AOI22_X1 U22649 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19726), .B1(
        n19725), .B2(n19710), .ZN(n19711) );
  OAI211_X1 U22650 ( .C1(n19713), .C2(n19729), .A(n19712), .B(n19711), .ZN(
        P2_U3173) );
  AOI22_X1 U22651 ( .A1(n19723), .A2(n19715), .B1(n19721), .B2(n19714), .ZN(
        n19718) );
  AOI22_X1 U22652 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19726), .B1(
        n19725), .B2(n19716), .ZN(n19717) );
  OAI211_X1 U22653 ( .C1(n19719), .C2(n19729), .A(n19718), .B(n19717), .ZN(
        P2_U3174) );
  AOI22_X1 U22654 ( .A1(n19723), .A2(n19722), .B1(n19721), .B2(n19720), .ZN(
        n19728) );
  AOI22_X1 U22655 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19726), .B1(
        n19725), .B2(n19724), .ZN(n19727) );
  OAI211_X1 U22656 ( .C1(n19730), .C2(n19729), .A(n19728), .B(n19727), .ZN(
        P2_U3175) );
  AND2_X1 U22657 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19731), .ZN(
        P2_U3179) );
  AND2_X1 U22658 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19731), .ZN(
        P2_U3180) );
  AND2_X1 U22659 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19731), .ZN(
        P2_U3181) );
  AND2_X1 U22660 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19731), .ZN(
        P2_U3182) );
  AND2_X1 U22661 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19731), .ZN(
        P2_U3183) );
  AND2_X1 U22662 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19731), .ZN(
        P2_U3184) );
  AND2_X1 U22663 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19731), .ZN(
        P2_U3185) );
  AND2_X1 U22664 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19731), .ZN(
        P2_U3186) );
  AND2_X1 U22665 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19731), .ZN(
        P2_U3187) );
  AND2_X1 U22666 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19731), .ZN(
        P2_U3188) );
  AND2_X1 U22667 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19731), .ZN(
        P2_U3189) );
  AND2_X1 U22668 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19731), .ZN(
        P2_U3190) );
  AND2_X1 U22669 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19731), .ZN(
        P2_U3191) );
  AND2_X1 U22670 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19731), .ZN(
        P2_U3192) );
  AND2_X1 U22671 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19731), .ZN(
        P2_U3193) );
  INV_X1 U22672 ( .A(P2_DATAWIDTH_REG_16__SCAN_IN), .ZN(n21062) );
  NOR2_X1 U22673 ( .A1(n21062), .A2(n19816), .ZN(P2_U3194) );
  AND2_X1 U22674 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19731), .ZN(
        P2_U3195) );
  AND2_X1 U22675 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19731), .ZN(
        P2_U3196) );
  AND2_X1 U22676 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19731), .ZN(
        P2_U3197) );
  AND2_X1 U22677 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19731), .ZN(
        P2_U3198) );
  AND2_X1 U22678 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19731), .ZN(
        P2_U3199) );
  AND2_X1 U22679 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19731), .ZN(
        P2_U3200) );
  AND2_X1 U22680 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19731), .ZN(P2_U3201) );
  AND2_X1 U22681 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19731), .ZN(P2_U3202) );
  AND2_X1 U22682 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19731), .ZN(P2_U3203) );
  AND2_X1 U22683 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19731), .ZN(P2_U3204) );
  AND2_X1 U22684 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19731), .ZN(P2_U3205) );
  AND2_X1 U22685 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19731), .ZN(P2_U3206) );
  AND2_X1 U22686 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19731), .ZN(P2_U3207) );
  AND2_X1 U22687 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19731), .ZN(P2_U3208) );
  NOR2_X1 U22688 ( .A1(n20818), .A2(n19738), .ZN(n19751) );
  NOR2_X1 U22689 ( .A1(n19732), .A2(n19736), .ZN(n19733) );
  NAND2_X1 U22690 ( .A1(n19743), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19746) );
  AOI21_X1 U22691 ( .B1(n19733), .B2(n19746), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19735) );
  AOI211_X1 U22692 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20809), .A(
        n19745), .B(n19866), .ZN(n19734) );
  OR3_X1 U22693 ( .A1(n19751), .A2(n19735), .A3(n19734), .ZN(P2_U3209) );
  AOI21_X1 U22694 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20809), .A(n19752), 
        .ZN(n19742) );
  NOR2_X1 U22695 ( .A1(n19736), .A2(n19742), .ZN(n19739) );
  AOI21_X1 U22696 ( .B1(n19739), .B2(n19738), .A(n19737), .ZN(n19740) );
  OAI211_X1 U22697 ( .C1(n20809), .C2(n19741), .A(n19740), .B(n19746), .ZN(
        P2_U3210) );
  AOI21_X1 U22698 ( .B1(n19744), .B2(n19743), .A(n19742), .ZN(n19750) );
  INV_X1 U22699 ( .A(n19745), .ZN(n19747) );
  OAI22_X1 U22700 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19747), .B1(NA), 
        .B2(n19746), .ZN(n19748) );
  OAI211_X1 U22701 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19748), .ZN(n19749) );
  OAI21_X1 U22702 ( .B1(n19751), .B2(n19750), .A(n19749), .ZN(P2_U3211) );
  INV_X1 U22703 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19756) );
  OAI222_X1 U22704 ( .A1(n19809), .A2(n19756), .B1(n19754), .B2(n19866), .C1(
        n19753), .C2(n19805), .ZN(P2_U3212) );
  OAI222_X1 U22705 ( .A1(n19805), .A2(n19756), .B1(n19755), .B2(n19866), .C1(
        n19758), .C2(n19809), .ZN(P2_U3213) );
  OAI222_X1 U22706 ( .A1(n19805), .A2(n19758), .B1(n19757), .B2(n19866), .C1(
        n10835), .C2(n19809), .ZN(P2_U3214) );
  INV_X1 U22707 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19760) );
  OAI222_X1 U22708 ( .A1(n19809), .A2(n19760), .B1(n19759), .B2(n19866), .C1(
        n10835), .C2(n19805), .ZN(P2_U3215) );
  OAI222_X1 U22709 ( .A1(n19809), .A2(n19762), .B1(n19761), .B2(n19866), .C1(
        n19760), .C2(n19805), .ZN(P2_U3216) );
  OAI222_X1 U22710 ( .A1(n19809), .A2(n19764), .B1(n19763), .B2(n19866), .C1(
        n19762), .C2(n19805), .ZN(P2_U3217) );
  INV_X1 U22711 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19766) );
  OAI222_X1 U22712 ( .A1(n19809), .A2(n19766), .B1(n19765), .B2(n19866), .C1(
        n19764), .C2(n19805), .ZN(P2_U3218) );
  OAI222_X1 U22713 ( .A1(n19809), .A2(n19768), .B1(n19767), .B2(n19866), .C1(
        n19766), .C2(n19805), .ZN(P2_U3219) );
  OAI222_X1 U22714 ( .A1(n19809), .A2(n19770), .B1(n19769), .B2(n19866), .C1(
        n19768), .C2(n19805), .ZN(P2_U3220) );
  INV_X1 U22715 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19772) );
  OAI222_X1 U22716 ( .A1(n19809), .A2(n19772), .B1(n19771), .B2(n19866), .C1(
        n19770), .C2(n19805), .ZN(P2_U3221) );
  OAI222_X1 U22717 ( .A1(n19809), .A2(n19774), .B1(n19773), .B2(n19866), .C1(
        n19772), .C2(n19805), .ZN(P2_U3222) );
  INV_X1 U22718 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19776) );
  OAI222_X1 U22719 ( .A1(n19809), .A2(n19776), .B1(n19775), .B2(n19866), .C1(
        n19774), .C2(n19805), .ZN(P2_U3223) );
  OAI222_X1 U22720 ( .A1(n19809), .A2(n19778), .B1(n19777), .B2(n19866), .C1(
        n19776), .C2(n19805), .ZN(P2_U3224) );
  INV_X1 U22721 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19780) );
  OAI222_X1 U22722 ( .A1(n19809), .A2(n19780), .B1(n19779), .B2(n19866), .C1(
        n19778), .C2(n19805), .ZN(P2_U3225) );
  INV_X1 U22723 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19782) );
  OAI222_X1 U22724 ( .A1(n19809), .A2(n19782), .B1(n19781), .B2(n19866), .C1(
        n19780), .C2(n19805), .ZN(P2_U3226) );
  OAI222_X1 U22725 ( .A1(n19809), .A2(n19784), .B1(n19783), .B2(n19866), .C1(
        n19782), .C2(n19805), .ZN(P2_U3227) );
  OAI222_X1 U22726 ( .A1(n19809), .A2(n15192), .B1(n19785), .B2(n19866), .C1(
        n19784), .C2(n19805), .ZN(P2_U3228) );
  OAI222_X1 U22727 ( .A1(n19809), .A2(n19787), .B1(n19786), .B2(n19866), .C1(
        n15192), .C2(n19805), .ZN(P2_U3229) );
  OAI222_X1 U22728 ( .A1(n19809), .A2(n19789), .B1(n19788), .B2(n19866), .C1(
        n19787), .C2(n19805), .ZN(P2_U3230) );
  OAI222_X1 U22729 ( .A1(n19809), .A2(n19790), .B1(n21075), .B2(n19866), .C1(
        n19789), .C2(n19805), .ZN(P2_U3231) );
  OAI222_X1 U22730 ( .A1(n19809), .A2(n19792), .B1(n19791), .B2(n19866), .C1(
        n19790), .C2(n19805), .ZN(P2_U3232) );
  OAI222_X1 U22731 ( .A1(n19809), .A2(n19794), .B1(n19793), .B2(n19866), .C1(
        n19792), .C2(n19805), .ZN(P2_U3233) );
  OAI222_X1 U22732 ( .A1(n19809), .A2(n15117), .B1(n19795), .B2(n19866), .C1(
        n19794), .C2(n19805), .ZN(P2_U3234) );
  OAI222_X1 U22733 ( .A1(n19809), .A2(n19797), .B1(n19796), .B2(n19866), .C1(
        n15117), .C2(n19805), .ZN(P2_U3235) );
  OAI222_X1 U22734 ( .A1(n19809), .A2(n11404), .B1(n19798), .B2(n19866), .C1(
        n19797), .C2(n19805), .ZN(P2_U3236) );
  OAI222_X1 U22735 ( .A1(n19809), .A2(n19801), .B1(n19799), .B2(n19866), .C1(
        n11404), .C2(n19805), .ZN(P2_U3237) );
  OAI222_X1 U22736 ( .A1(n19805), .A2(n19801), .B1(n19800), .B2(n19866), .C1(
        n11294), .C2(n19809), .ZN(P2_U3238) );
  OAI222_X1 U22737 ( .A1(n19809), .A2(n19803), .B1(n19802), .B2(n19866), .C1(
        n11294), .C2(n19805), .ZN(P2_U3239) );
  INV_X1 U22738 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19806) );
  OAI222_X1 U22739 ( .A1(n19809), .A2(n19806), .B1(n19804), .B2(n19866), .C1(
        n19803), .C2(n19805), .ZN(P2_U3240) );
  OAI222_X1 U22740 ( .A1(n19809), .A2(n19808), .B1(n19807), .B2(n19866), .C1(
        n19806), .C2(n19805), .ZN(P2_U3241) );
  OAI22_X1 U22741 ( .A1(n19867), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19866), .ZN(n19810) );
  INV_X1 U22742 ( .A(n19810), .ZN(P2_U3585) );
  MUX2_X1 U22743 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19867), .Z(P2_U3586) );
  OAI22_X1 U22744 ( .A1(n19867), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19866), .ZN(n19811) );
  INV_X1 U22745 ( .A(n19811), .ZN(P2_U3587) );
  OAI22_X1 U22746 ( .A1(n19867), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19866), .ZN(n19812) );
  INV_X1 U22747 ( .A(n19812), .ZN(P2_U3588) );
  OAI21_X1 U22748 ( .B1(n19816), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19814), 
        .ZN(n19813) );
  INV_X1 U22749 ( .A(n19813), .ZN(P2_U3591) );
  OAI21_X1 U22750 ( .B1(n19816), .B2(n19815), .A(n19814), .ZN(P2_U3592) );
  NAND2_X1 U22751 ( .A1(n19817), .A2(n19830), .ZN(n19824) );
  OAI21_X1 U22752 ( .B1(n19819), .B2(n19818), .A(n19830), .ZN(n19821) );
  NAND2_X1 U22753 ( .A1(n19821), .A2(n19820), .ZN(n19834) );
  NAND2_X1 U22754 ( .A1(n19834), .A2(n19822), .ZN(n19823) );
  OAI211_X1 U22755 ( .C1(n19826), .C2(n19825), .A(n19824), .B(n19823), .ZN(
        n19827) );
  INV_X1 U22756 ( .A(n19827), .ZN(n19828) );
  AOI22_X1 U22757 ( .A1(n19853), .A2(n19829), .B1(n19828), .B2(n19854), .ZN(
        P2_U3602) );
  NAND2_X1 U22758 ( .A1(n19830), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19841) );
  OAI21_X1 U22759 ( .B1(n19832), .B2(n19841), .A(n19831), .ZN(n19833) );
  AOI22_X1 U22760 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19835), .B1(n19834), 
        .B2(n19833), .ZN(n19836) );
  AOI22_X1 U22761 ( .A1(n19853), .A2(n19837), .B1(n19836), .B2(n19854), .ZN(
        P2_U3603) );
  INV_X1 U22762 ( .A(n19838), .ZN(n19839) );
  NAND3_X1 U22763 ( .A1(n19842), .A2(n19847), .A3(n19839), .ZN(n19840) );
  OAI21_X1 U22764 ( .B1(n19842), .B2(n19841), .A(n19840), .ZN(n19843) );
  AOI21_X1 U22765 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19844), .A(n19843), 
        .ZN(n19845) );
  AOI22_X1 U22766 ( .A1(n19853), .A2(n19846), .B1(n19845), .B2(n19854), .ZN(
        P2_U3604) );
  INV_X1 U22767 ( .A(n19847), .ZN(n19849) );
  OAI21_X1 U22768 ( .B1(n19850), .B2(n19849), .A(n19848), .ZN(n19851) );
  AOI21_X1 U22769 ( .B1(n19855), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19851), 
        .ZN(n19852) );
  OAI22_X1 U22770 ( .A1(n19855), .A2(n19854), .B1(n19853), .B2(n19852), .ZN(
        P2_U3605) );
  INV_X1 U22771 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19856) );
  AOI22_X1 U22772 ( .A1(n19866), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19856), 
        .B2(n19867), .ZN(P2_U3608) );
  INV_X1 U22773 ( .A(n19857), .ZN(n19858) );
  NAND2_X1 U22774 ( .A1(n19859), .A2(n19858), .ZN(n19860) );
  OAI211_X1 U22775 ( .C1(n19863), .C2(n19862), .A(n19861), .B(n19860), .ZN(
        n19865) );
  MUX2_X1 U22776 ( .A(P2_MORE_REG_SCAN_IN), .B(n19865), .S(n19864), .Z(
        P2_U3609) );
  OAI22_X1 U22777 ( .A1(n19867), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19866), .ZN(n19868) );
  INV_X1 U22778 ( .A(n19868), .ZN(P2_U3611) );
  AND2_X1 U22779 ( .A1(n20813), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n19870) );
  INV_X1 U22780 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19869) );
  AOI21_X1 U22781 ( .B1(n19870), .B2(n19869), .A(n20904), .ZN(P1_U2802) );
  OAI21_X1 U22782 ( .B1(n19872), .B2(n19871), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19873) );
  OAI21_X1 U22783 ( .B1(n19874), .B2(n20804), .A(n19873), .ZN(P1_U2803) );
  INV_X1 U22784 ( .A(n20904), .ZN(n20905) );
  NOR2_X1 U22785 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19876) );
  OAI21_X1 U22786 ( .B1(n19876), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20905), .ZN(
        n19875) );
  OAI21_X1 U22787 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20905), .A(n19875), 
        .ZN(P1_U2804) );
  AOI21_X1 U22788 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20813), .A(n20904), 
        .ZN(n20807) );
  OAI21_X1 U22789 ( .B1(BS16), .B2(n19876), .A(n20807), .ZN(n20872) );
  OAI21_X1 U22790 ( .B1(n20807), .B2(n20466), .A(n20872), .ZN(P1_U2805) );
  OAI21_X1 U22791 ( .B1(n19879), .B2(n19878), .A(n19877), .ZN(P1_U2806) );
  NOR4_X1 U22792 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19883) );
  NOR4_X1 U22793 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19882) );
  NOR4_X1 U22794 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_29__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19881) );
  NOR4_X1 U22795 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19880) );
  NAND4_X1 U22796 ( .A1(n19883), .A2(n19882), .A3(n19881), .A4(n19880), .ZN(
        n19889) );
  NOR4_X1 U22797 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19887) );
  AOI211_X1 U22798 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19886) );
  NOR4_X1 U22799 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19885) );
  NOR4_X1 U22800 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19884) );
  NAND4_X1 U22801 ( .A1(n19887), .A2(n19886), .A3(n19885), .A4(n19884), .ZN(
        n19888) );
  NOR2_X1 U22802 ( .A1(n19889), .A2(n19888), .ZN(n20892) );
  INV_X1 U22803 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19891) );
  NOR3_X1 U22804 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19892) );
  OAI21_X1 U22805 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19892), .A(n20892), .ZN(
        n19890) );
  OAI21_X1 U22806 ( .B1(n20892), .B2(n19891), .A(n19890), .ZN(P1_U2807) );
  INV_X1 U22807 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19894) );
  NOR2_X1 U22808 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20886) );
  OAI21_X1 U22809 ( .B1(n19892), .B2(n20886), .A(n20892), .ZN(n19893) );
  OAI21_X1 U22810 ( .B1(n20892), .B2(n19894), .A(n19893), .ZN(P1_U2808) );
  NOR2_X1 U22811 ( .A1(n19965), .A2(n19895), .ZN(n19896) );
  NOR2_X1 U22812 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19896), .ZN(n19906) );
  NAND2_X1 U22813 ( .A1(n19932), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n19897) );
  OAI211_X1 U22814 ( .C1(n19899), .C2(n19898), .A(n19897), .B(n19921), .ZN(
        n19900) );
  AOI21_X1 U22815 ( .B1(n19940), .B2(n19901), .A(n19900), .ZN(n19905) );
  AOI22_X1 U22816 ( .A1(n19903), .A2(n19916), .B1(n19979), .B2(n19902), .ZN(
        n19904) );
  OAI211_X1 U22817 ( .C1(n19907), .C2(n19906), .A(n19905), .B(n19904), .ZN(
        P1_U2831) );
  AOI221_X1 U22818 ( .B1(n19931), .B2(n19961), .C1(n19913), .C2(n19961), .A(
        n19960), .ZN(n19929) );
  NOR2_X1 U22819 ( .A1(n19965), .A2(n19931), .ZN(n19933) );
  NAND2_X1 U22820 ( .A1(n19933), .A2(n19918), .ZN(n19914) );
  AOI21_X1 U22821 ( .B1(n19978), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19946), .ZN(n19908) );
  OAI21_X1 U22822 ( .B1(n19909), .B2(n19935), .A(n19908), .ZN(n19911) );
  NOR2_X1 U22823 ( .A1(n19987), .A2(n19999), .ZN(n19910) );
  AOI211_X1 U22824 ( .C1(n19996), .C2(n19940), .A(n19911), .B(n19910), .ZN(
        n19912) );
  OAI21_X1 U22825 ( .B1(n19914), .B2(n19913), .A(n19912), .ZN(n19915) );
  AOI21_X1 U22826 ( .B1(n19916), .B2(n19997), .A(n19915), .ZN(n19917) );
  OAI21_X1 U22827 ( .B1(n19918), .B2(n19929), .A(n19917), .ZN(P1_U2833) );
  INV_X1 U22828 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n19930) );
  NOR2_X1 U22829 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n19944), .ZN(n19919) );
  AOI22_X1 U22830 ( .A1(n19933), .A2(n19919), .B1(n19940), .B2(n20000), .ZN(
        n19928) );
  NAND2_X1 U22831 ( .A1(n19978), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n19920) );
  OAI211_X1 U22832 ( .C1(n19935), .C2(n19922), .A(n19921), .B(n19920), .ZN(
        n19926) );
  NOR2_X1 U22833 ( .A1(n19924), .A2(n19923), .ZN(n19925) );
  AOI211_X1 U22834 ( .C1(n19932), .C2(P1_EBX_REG_6__SCAN_IN), .A(n19926), .B(
        n19925), .ZN(n19927) );
  OAI211_X1 U22835 ( .C1(n19930), .C2(n19929), .A(n19928), .B(n19927), .ZN(
        P1_U2834) );
  AOI21_X1 U22836 ( .B1(n19961), .B2(n19931), .A(n19960), .ZN(n19958) );
  AOI22_X1 U22837 ( .A1(n19933), .A2(n19944), .B1(n19932), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n19943) );
  AOI21_X1 U22838 ( .B1(n19978), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n19946), .ZN(n19934) );
  OAI21_X1 U22839 ( .B1(n19936), .B2(n19935), .A(n19934), .ZN(n19939) );
  NOR2_X1 U22840 ( .A1(n20006), .A2(n19937), .ZN(n19938) );
  AOI211_X1 U22841 ( .C1(n19941), .C2(n19940), .A(n19939), .B(n19938), .ZN(
        n19942) );
  OAI211_X1 U22842 ( .C1(n19944), .C2(n19958), .A(n19943), .B(n19942), .ZN(
        P1_U2835) );
  INV_X1 U22843 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n19975) );
  NAND2_X1 U22844 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n19962) );
  NOR2_X1 U22845 ( .A1(n19975), .A2(n19962), .ZN(n19945) );
  AOI21_X1 U22846 ( .B1(n19961), .B2(n19945), .A(P1_REIP_REG_4__SCAN_IN), .ZN(
        n19959) );
  AOI21_X1 U22847 ( .B1(n19978), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n19946), .ZN(n19949) );
  INV_X1 U22848 ( .A(n19981), .ZN(n19966) );
  NAND2_X1 U22849 ( .A1(n19966), .A2(n19947), .ZN(n19948) );
  OAI211_X1 U22850 ( .C1(n19985), .C2(n19950), .A(n19949), .B(n19948), .ZN(
        n19953) );
  NOR2_X1 U22851 ( .A1(n19987), .A2(n19951), .ZN(n19952) );
  NOR2_X1 U22852 ( .A1(n19953), .A2(n19952), .ZN(n19957) );
  AOI22_X1 U22853 ( .A1(n19955), .A2(n19991), .B1(n19954), .B2(n19979), .ZN(
        n19956) );
  OAI211_X1 U22854 ( .C1(n19959), .C2(n19958), .A(n19957), .B(n19956), .ZN(
        P1_U2836) );
  AOI21_X1 U22855 ( .B1(n19961), .B2(n19962), .A(n19960), .ZN(n19995) );
  INV_X1 U22856 ( .A(n19962), .ZN(n19963) );
  NAND2_X1 U22857 ( .A1(n19963), .A2(n19975), .ZN(n19964) );
  OAI22_X1 U22858 ( .A1(n19965), .A2(n19964), .B1(n19985), .B2(n20010), .ZN(
        n19970) );
  INV_X1 U22859 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n20015) );
  NAND2_X1 U22860 ( .A1(n19966), .A2(n13145), .ZN(n19968) );
  NAND2_X1 U22861 ( .A1(n19978), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n19967) );
  OAI211_X1 U22862 ( .C1(n19987), .C2(n20015), .A(n19968), .B(n19967), .ZN(
        n19969) );
  NOR2_X1 U22863 ( .A1(n19970), .A2(n19969), .ZN(n19974) );
  INV_X1 U22864 ( .A(n19971), .ZN(n20013) );
  AOI22_X1 U22865 ( .A1(n20013), .A2(n19991), .B1(n19972), .B2(n19979), .ZN(
        n19973) );
  OAI211_X1 U22866 ( .C1(n19995), .C2(n19975), .A(n19974), .B(n19973), .ZN(
        P1_U2837) );
  AOI21_X1 U22867 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19976), .A(
        P1_REIP_REG_2__SCAN_IN), .ZN(n19994) );
  INV_X1 U22868 ( .A(n19977), .ZN(n19980) );
  AOI22_X1 U22869 ( .A1(n19980), .A2(n19979), .B1(n19978), .B2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n19983) );
  OR2_X1 U22870 ( .A1(n19981), .A2(n13122), .ZN(n19982) );
  OAI211_X1 U22871 ( .C1(n19985), .C2(n19984), .A(n19983), .B(n19982), .ZN(
        n19989) );
  NOR2_X1 U22872 ( .A1(n19987), .A2(n19986), .ZN(n19988) );
  NOR2_X1 U22873 ( .A1(n19989), .A2(n19988), .ZN(n19993) );
  NAND2_X1 U22874 ( .A1(n19991), .A2(n19990), .ZN(n19992) );
  OAI211_X1 U22875 ( .C1(n19995), .C2(n19994), .A(n19993), .B(n19992), .ZN(
        P1_U2838) );
  AOI22_X1 U22876 ( .A1(n19997), .A2(n12640), .B1(n20012), .B2(n19996), .ZN(
        n19998) );
  OAI21_X1 U22877 ( .B1(n20016), .B2(n19999), .A(n19998), .ZN(P1_U2865) );
  AOI22_X1 U22878 ( .A1(n20001), .A2(n12640), .B1(n20012), .B2(n20000), .ZN(
        n20002) );
  OAI21_X1 U22879 ( .B1(n20016), .B2(n20003), .A(n20002), .ZN(P1_U2866) );
  OAI22_X1 U22880 ( .A1(n20006), .A2(n14350), .B1(n20005), .B2(n20004), .ZN(
        n20007) );
  INV_X1 U22881 ( .A(n20007), .ZN(n20008) );
  OAI21_X1 U22882 ( .B1(n20016), .B2(n20009), .A(n20008), .ZN(P1_U2867) );
  INV_X1 U22883 ( .A(n20010), .ZN(n20011) );
  AOI22_X1 U22884 ( .A1(n20013), .A2(n12640), .B1(n20012), .B2(n20011), .ZN(
        n20014) );
  OAI21_X1 U22885 ( .B1(n20016), .B2(n20015), .A(n20014), .ZN(P1_U2869) );
  AOI22_X1 U22886 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20017) );
  OAI21_X1 U22887 ( .B1(n12265), .B2(n20041), .A(n20017), .ZN(P1_U2921) );
  INV_X1 U22888 ( .A(P1_LWORD_REG_14__SCAN_IN), .ZN(n21098) );
  AOI22_X1 U22889 ( .A1(P1_EAX_REG_14__SCAN_IN), .A2(n20026), .B1(n20038), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20018) );
  OAI21_X1 U22890 ( .B1(n21098), .B2(n20019), .A(n20018), .ZN(P1_U2922) );
  AOI22_X1 U22891 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20020) );
  OAI21_X1 U22892 ( .B1(n14065), .B2(n20041), .A(n20020), .ZN(P1_U2923) );
  AOI22_X1 U22893 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20021) );
  OAI21_X1 U22894 ( .B1(n13967), .B2(n20041), .A(n20021), .ZN(P1_U2924) );
  AOI22_X1 U22895 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20022) );
  OAI21_X1 U22896 ( .B1(n13892), .B2(n20041), .A(n20022), .ZN(P1_U2925) );
  AOI22_X1 U22897 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20023) );
  OAI21_X1 U22898 ( .B1(n13804), .B2(n20041), .A(n20023), .ZN(P1_U2926) );
  INV_X1 U22899 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20025) );
  AOI22_X1 U22900 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20024) );
  OAI21_X1 U22901 ( .B1(n20025), .B2(n20041), .A(n20024), .ZN(P1_U2927) );
  AOI22_X1 U22902 ( .A1(P1_EAX_REG_8__SCAN_IN), .A2(n20026), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20039), .ZN(n20027) );
  OAI21_X1 U22903 ( .B1(n21043), .B2(n20028), .A(n20027), .ZN(P1_U2928) );
  AOI22_X1 U22904 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20029) );
  OAI21_X1 U22905 ( .B1(n13514), .B2(n20041), .A(n20029), .ZN(P1_U2929) );
  AOI22_X1 U22906 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20030) );
  OAI21_X1 U22907 ( .B1(n20031), .B2(n20041), .A(n20030), .ZN(P1_U2930) );
  AOI22_X1 U22908 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20032) );
  OAI21_X1 U22909 ( .B1(n12105), .B2(n20041), .A(n20032), .ZN(P1_U2931) );
  AOI22_X1 U22910 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20033) );
  OAI21_X1 U22911 ( .B1(n20034), .B2(n20041), .A(n20033), .ZN(P1_U2932) );
  AOI22_X1 U22912 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20035) );
  OAI21_X1 U22913 ( .B1(n13104), .B2(n20041), .A(n20035), .ZN(P1_U2933) );
  AOI22_X1 U22914 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20036) );
  OAI21_X1 U22915 ( .B1(n12071), .B2(n20041), .A(n20036), .ZN(P1_U2934) );
  AOI22_X1 U22916 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20037) );
  OAI21_X1 U22917 ( .B1(n12064), .B2(n20041), .A(n20037), .ZN(P1_U2935) );
  AOI22_X1 U22918 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20039), .B1(n20038), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20040) );
  OAI21_X1 U22919 ( .B1(n20042), .B2(n20041), .A(n20040), .ZN(P1_U2936) );
  AOI22_X1 U22920 ( .A1(n20069), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20066), .ZN(n20044) );
  NAND2_X1 U22921 ( .A1(n20054), .A2(n20043), .ZN(n20056) );
  NAND2_X1 U22922 ( .A1(n20044), .A2(n20056), .ZN(P1_U2945) );
  AOI22_X1 U22923 ( .A1(n20069), .A2(P1_EAX_REG_25__SCAN_IN), .B1(n20066), 
        .B2(P1_UWORD_REG_9__SCAN_IN), .ZN(n20046) );
  NAND2_X1 U22924 ( .A1(n20054), .A2(n20045), .ZN(n20058) );
  NAND2_X1 U22925 ( .A1(n20046), .A2(n20058), .ZN(P1_U2946) );
  AOI22_X1 U22926 ( .A1(n20069), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20066), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20048) );
  NAND2_X1 U22927 ( .A1(n20054), .A2(n20047), .ZN(n20060) );
  NAND2_X1 U22928 ( .A1(n20048), .A2(n20060), .ZN(P1_U2947) );
  AOI22_X1 U22929 ( .A1(n20069), .A2(P1_EAX_REG_28__SCAN_IN), .B1(n20066), 
        .B2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20050) );
  NAND2_X1 U22930 ( .A1(n20054), .A2(n20049), .ZN(n20064) );
  NAND2_X1 U22931 ( .A1(n20050), .A2(n20064), .ZN(P1_U2949) );
  AOI22_X1 U22932 ( .A1(n20069), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20066), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20052) );
  NAND2_X1 U22933 ( .A1(n20054), .A2(n20051), .ZN(n20067) );
  NAND2_X1 U22934 ( .A1(n20052), .A2(n20067), .ZN(P1_U2950) );
  AOI22_X1 U22935 ( .A1(n20069), .A2(P1_EAX_REG_30__SCAN_IN), .B1(n20066), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20055) );
  NAND2_X1 U22936 ( .A1(n20054), .A2(n20053), .ZN(n20070) );
  NAND2_X1 U22937 ( .A1(n20055), .A2(n20070), .ZN(P1_U2951) );
  AOI22_X1 U22938 ( .A1(n20069), .A2(P1_EAX_REG_8__SCAN_IN), .B1(n20066), .B2(
        P1_LWORD_REG_8__SCAN_IN), .ZN(n20057) );
  NAND2_X1 U22939 ( .A1(n20057), .A2(n20056), .ZN(P1_U2960) );
  AOI22_X1 U22940 ( .A1(n20069), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20066), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20059) );
  NAND2_X1 U22941 ( .A1(n20059), .A2(n20058), .ZN(P1_U2961) );
  AOI22_X1 U22942 ( .A1(n20069), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20066), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20061) );
  NAND2_X1 U22943 ( .A1(n20061), .A2(n20060), .ZN(P1_U2962) );
  AOI22_X1 U22944 ( .A1(n20069), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20066), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20063) );
  NAND2_X1 U22945 ( .A1(n20063), .A2(n20062), .ZN(P1_U2963) );
  AOI22_X1 U22946 ( .A1(n20069), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20066), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20065) );
  NAND2_X1 U22947 ( .A1(n20065), .A2(n20064), .ZN(P1_U2964) );
  AOI22_X1 U22948 ( .A1(n20069), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20066), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20068) );
  NAND2_X1 U22949 ( .A1(n20068), .A2(n20067), .ZN(P1_U2965) );
  AOI22_X1 U22950 ( .A1(n20069), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20066), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20071) );
  NAND2_X1 U22951 ( .A1(n20071), .A2(n20070), .ZN(P1_U2966) );
  AOI21_X1 U22952 ( .B1(n20073), .B2(n20091), .A(n20072), .ZN(n20086) );
  AOI22_X1 U22953 ( .A1(n20074), .A2(n20086), .B1(n13376), .B2(
        P1_REIP_REG_0__SCAN_IN), .ZN(n20078) );
  OAI21_X1 U22954 ( .B1(n20076), .B2(n20075), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20077) );
  OAI211_X1 U22955 ( .C1(n20079), .C2(n20101), .A(n20078), .B(n20077), .ZN(
        P1_U2999) );
  AOI21_X1 U22956 ( .B1(n13376), .B2(P1_REIP_REG_0__SCAN_IN), .A(n20080), .ZN(
        n20082) );
  OAI211_X1 U22957 ( .C1(n20084), .C2(n20083), .A(n20082), .B(n20081), .ZN(
        n20085) );
  AOI21_X1 U22958 ( .B1(n20087), .B2(n20086), .A(n20085), .ZN(n20088) );
  OAI221_X1 U22959 ( .B1(n20091), .B2(n20090), .C1(n20091), .C2(n20089), .A(
        n20088), .ZN(P1_U3031) );
  INV_X1 U22960 ( .A(n20883), .ZN(n20092) );
  AND2_X1 U22961 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n20092), .ZN(
        P1_U3032) );
  NAND2_X1 U22962 ( .A1(n13020), .A2(n13227), .ZN(n20551) );
  NAND3_X1 U22963 ( .A1(n20911), .A2(n20741), .A3(n20909), .ZN(n20093) );
  NAND2_X1 U22964 ( .A1(n20741), .A2(n20466), .ZN(n20585) );
  NAND2_X1 U22965 ( .A1(n20093), .A2(n20585), .ZN(n20109) );
  OR2_X1 U22966 ( .A1(n13145), .A2(n20094), .ZN(n20224) );
  NOR2_X1 U22967 ( .A1(n20224), .A2(n9946), .ZN(n20107) );
  NAND2_X1 U22968 ( .A1(n20109), .A2(n20107), .ZN(n20098) );
  INV_X1 U22969 ( .A(n20420), .ZN(n20095) );
  AND2_X1 U22970 ( .A1(n20095), .A2(n20501), .ZN(n20265) );
  NAND2_X1 U22971 ( .A1(n20106), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20507) );
  INV_X1 U22972 ( .A(n20507), .ZN(n20096) );
  NAND2_X1 U22973 ( .A1(n20265), .A2(n20096), .ZN(n20097) );
  AOI22_X2 U22974 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n9636), .B1(DATAI_24_), 
        .B2(n9632), .ZN(n20692) );
  NAND2_X1 U22975 ( .A1(n20173), .A2(n20104), .ZN(n20738) );
  NAND2_X1 U22976 ( .A1(n20882), .A2(n20419), .ZN(n20186) );
  OR2_X1 U22977 ( .A1(n20583), .A2(n20186), .ZN(n20907) );
  OAI22_X1 U22978 ( .A1(n20692), .A2(n20909), .B1(n20738), .B2(n20907), .ZN(
        n20105) );
  INV_X1 U22979 ( .A(n20105), .ZN(n20112) );
  OR2_X1 U22980 ( .A1(n20106), .A2(n20383), .ZN(n20592) );
  INV_X1 U22981 ( .A(n20107), .ZN(n20108) );
  AOI22_X1 U22982 ( .A1(n20109), .A2(n20108), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20907), .ZN(n20110) );
  OAI211_X1 U22983 ( .C1(n20265), .C2(n20383), .A(n20504), .B(n20110), .ZN(
        n20917) );
  AOI22_X1 U22984 ( .A1(DATAI_16_), .A2(n9632), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n9636), .ZN(n20753) );
  INV_X1 U22985 ( .A(n20753), .ZN(n20689) );
  AOI22_X1 U22986 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20917), .B1(
        n20181), .B2(n20689), .ZN(n20111) );
  OAI211_X1 U22987 ( .C1(n20914), .C2(n20739), .A(n20112), .B(n20111), .ZN(
        P1_U3033) );
  NAND2_X1 U22988 ( .A1(n20173), .A2(n20114), .ZN(n20754) );
  OAI22_X1 U22989 ( .A1(n20697), .A2(n20909), .B1(n20754), .B2(n20907), .ZN(
        n20115) );
  INV_X1 U22990 ( .A(n20115), .ZN(n20117) );
  AOI22_X1 U22991 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n9636), .B1(DATAI_17_), 
        .B2(n9632), .ZN(n20760) );
  INV_X1 U22992 ( .A(n20760), .ZN(n20694) );
  AOI22_X1 U22993 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20917), .B1(
        n20181), .B2(n20694), .ZN(n20116) );
  OAI211_X1 U22994 ( .C1(n20914), .C2(n20755), .A(n20117), .B(n20116), .ZN(
        P1_U3034) );
  AOI22_X1 U22995 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n9636), .B1(DATAI_26_), 
        .B2(n9632), .ZN(n20702) );
  NAND2_X1 U22996 ( .A1(n20173), .A2(n20119), .ZN(n20761) );
  OAI22_X1 U22997 ( .A1(n20702), .A2(n20909), .B1(n20761), .B2(n20907), .ZN(
        n20120) );
  INV_X1 U22998 ( .A(n20120), .ZN(n20122) );
  INV_X1 U22999 ( .A(n20767), .ZN(n20699) );
  AOI22_X1 U23000 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20917), .B1(
        n20181), .B2(n20699), .ZN(n20121) );
  OAI211_X1 U23001 ( .C1(n20914), .C2(n20762), .A(n20122), .B(n20121), .ZN(
        P1_U3035) );
  AOI22_X2 U23002 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n9636), .B1(DATAI_27_), 
        .B2(n9632), .ZN(n20707) );
  NAND2_X1 U23003 ( .A1(n20173), .A2(n20124), .ZN(n20768) );
  OAI22_X1 U23004 ( .A1(n20707), .A2(n20909), .B1(n20768), .B2(n20907), .ZN(
        n20125) );
  INV_X1 U23005 ( .A(n20125), .ZN(n20127) );
  AOI22_X1 U23006 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n9636), .B1(DATAI_19_), 
        .B2(n9632), .ZN(n20774) );
  INV_X1 U23007 ( .A(n20774), .ZN(n20704) );
  AOI22_X1 U23008 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20917), .B1(
        n20181), .B2(n20704), .ZN(n20126) );
  OAI211_X1 U23009 ( .C1(n20914), .C2(n20769), .A(n20127), .B(n20126), .ZN(
        P1_U3036) );
  AOI22_X2 U23010 ( .A1(DATAI_20_), .A2(n9632), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n9636), .ZN(n20781) );
  AOI22_X1 U23011 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n9636), .B1(DATAI_28_), 
        .B2(n9632), .ZN(n20712) );
  NAND2_X1 U23012 ( .A1(n20173), .A2(n11878), .ZN(n20775) );
  OAI22_X1 U23013 ( .A1(n20712), .A2(n20909), .B1(n20775), .B2(n20907), .ZN(
        n20128) );
  INV_X1 U23014 ( .A(n20128), .ZN(n20131) );
  INV_X1 U23015 ( .A(n20914), .ZN(n20139) );
  AOI22_X1 U23016 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20917), .B1(
        n20612), .B2(n20139), .ZN(n20130) );
  OAI211_X1 U23017 ( .C1(n20781), .C2(n20911), .A(n20131), .B(n20130), .ZN(
        P1_U3037) );
  AOI22_X1 U23018 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n9636), .B1(DATAI_21_), 
        .B2(n9632), .ZN(n20788) );
  NAND2_X1 U23019 ( .A1(n20173), .A2(n11877), .ZN(n20782) );
  OAI22_X1 U23020 ( .A1(n20717), .A2(n20909), .B1(n20782), .B2(n20907), .ZN(
        n20132) );
  INV_X1 U23021 ( .A(n20132), .ZN(n20135) );
  INV_X1 U23022 ( .A(n20783), .ZN(n20616) );
  AOI22_X1 U23023 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20917), .B1(
        n20616), .B2(n20139), .ZN(n20134) );
  OAI211_X1 U23024 ( .C1(n20788), .C2(n20911), .A(n20135), .B(n20134), .ZN(
        P1_U3038) );
  NAND2_X1 U23025 ( .A1(n20173), .A2(n20136), .ZN(n20789) );
  OAI22_X1 U23026 ( .A1(n20722), .A2(n20909), .B1(n20789), .B2(n20907), .ZN(
        n20137) );
  INV_X1 U23027 ( .A(n20137), .ZN(n20141) );
  AOI22_X1 U23028 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20917), .B1(
        n20620), .B2(n20139), .ZN(n20140) );
  OAI211_X1 U23029 ( .C1(n20795), .C2(n20911), .A(n20141), .B(n20140), .ZN(
        P1_U3039) );
  OR2_X1 U23030 ( .A1(n20224), .A2(n20634), .ZN(n20143) );
  NOR2_X1 U23031 ( .A1(n20186), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20150) );
  INV_X1 U23032 ( .A(n20150), .ZN(n20142) );
  OR2_X1 U23033 ( .A1(n20635), .A2(n20142), .ZN(n20177) );
  NAND2_X1 U23034 ( .A1(n20143), .A2(n20177), .ZN(n20147) );
  NAND2_X1 U23035 ( .A1(n20147), .A2(n20741), .ZN(n20145) );
  NAND2_X1 U23036 ( .A1(n20150), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20144) );
  OAI22_X1 U23037 ( .A1(n20739), .A2(n20176), .B1(n20738), .B2(n20177), .ZN(
        n20146) );
  INV_X1 U23038 ( .A(n20146), .ZN(n20152) );
  INV_X1 U23039 ( .A(n20147), .ZN(n20148) );
  OAI211_X1 U23040 ( .C1(n20229), .C2(n20466), .A(n20741), .B(n20148), .ZN(
        n20149) );
  OAI211_X1 U23041 ( .C1(n20741), .C2(n20150), .A(n20748), .B(n20149), .ZN(
        n20182) );
  INV_X1 U23042 ( .A(n20221), .ZN(n20169) );
  AOI22_X1 U23043 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20182), .B1(
        n20169), .B2(n20689), .ZN(n20151) );
  OAI211_X1 U23044 ( .C1(n20692), .C2(n20911), .A(n20152), .B(n20151), .ZN(
        P1_U3041) );
  OAI22_X1 U23045 ( .A1(n20755), .A2(n20176), .B1(n20754), .B2(n20177), .ZN(
        n20153) );
  INV_X1 U23046 ( .A(n20153), .ZN(n20155) );
  INV_X1 U23047 ( .A(n20697), .ZN(n20757) );
  AOI22_X1 U23048 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20182), .B1(
        n20181), .B2(n20757), .ZN(n20154) );
  OAI211_X1 U23049 ( .C1(n20760), .C2(n20221), .A(n20155), .B(n20154), .ZN(
        P1_U3042) );
  OAI22_X1 U23050 ( .A1(n20762), .A2(n20176), .B1(n20761), .B2(n20177), .ZN(
        n20156) );
  INV_X1 U23051 ( .A(n20156), .ZN(n20158) );
  INV_X1 U23052 ( .A(n20702), .ZN(n20764) );
  AOI22_X1 U23053 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20182), .B1(
        n20181), .B2(n20764), .ZN(n20157) );
  OAI211_X1 U23054 ( .C1(n20767), .C2(n20221), .A(n20158), .B(n20157), .ZN(
        P1_U3043) );
  OAI22_X1 U23055 ( .A1(n20769), .A2(n20176), .B1(n20768), .B2(n20177), .ZN(
        n20159) );
  INV_X1 U23056 ( .A(n20159), .ZN(n20161) );
  AOI22_X1 U23057 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20182), .B1(
        n20169), .B2(n20704), .ZN(n20160) );
  OAI211_X1 U23058 ( .C1(n20707), .C2(n20911), .A(n20161), .B(n20160), .ZN(
        P1_U3044) );
  OAI22_X1 U23059 ( .A1(n20776), .A2(n20176), .B1(n20775), .B2(n20177), .ZN(
        n20162) );
  INV_X1 U23060 ( .A(n20162), .ZN(n20164) );
  INV_X1 U23061 ( .A(n20712), .ZN(n20778) );
  AOI22_X1 U23062 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20182), .B1(
        n20181), .B2(n20778), .ZN(n20163) );
  OAI211_X1 U23063 ( .C1(n20781), .C2(n20221), .A(n20164), .B(n20163), .ZN(
        P1_U3045) );
  OAI22_X1 U23064 ( .A1(n20783), .A2(n20176), .B1(n20782), .B2(n20177), .ZN(
        n20165) );
  INV_X1 U23065 ( .A(n20165), .ZN(n20167) );
  INV_X1 U23066 ( .A(n20717), .ZN(n20785) );
  AOI22_X1 U23067 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20182), .B1(
        n20181), .B2(n20785), .ZN(n20166) );
  OAI211_X1 U23068 ( .C1(n20788), .C2(n20221), .A(n20167), .B(n20166), .ZN(
        P1_U3046) );
  OAI22_X1 U23069 ( .A1(n20790), .A2(n20176), .B1(n20789), .B2(n20177), .ZN(
        n20168) );
  INV_X1 U23070 ( .A(n20168), .ZN(n20171) );
  AOI22_X1 U23072 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20182), .B1(
        n20169), .B2(n9633), .ZN(n20170) );
  OAI211_X1 U23073 ( .C1(n20722), .C2(n20911), .A(n20171), .B(n20170), .ZN(
        P1_U3047) );
  AOI22_X1 U23074 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n9636), .B1(DATAI_23_), 
        .B2(n9632), .ZN(n20912) );
  NAND2_X1 U23075 ( .A1(n20173), .A2(n20172), .ZN(n20908) );
  NOR2_X1 U23076 ( .A1(n20175), .A2(n20174), .ZN(n20626) );
  OAI22_X1 U23077 ( .A1(n20908), .A2(n20177), .B1(n20176), .B2(n20913), .ZN(
        n20178) );
  INV_X1 U23078 ( .A(n20178), .ZN(n20184) );
  INV_X1 U23079 ( .A(n20910), .ZN(n20799) );
  AOI22_X1 U23080 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20182), .B1(
        n20181), .B2(n20799), .ZN(n20183) );
  OAI211_X1 U23081 ( .C1(n20912), .C2(n20221), .A(n20184), .B(n20183), .ZN(
        P1_U3048) );
  INV_X1 U23082 ( .A(n20186), .ZN(n20222) );
  NAND2_X1 U23083 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20222), .ZN(
        n20233) );
  NOR2_X1 U23084 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20233), .ZN(
        n20189) );
  INV_X1 U23085 ( .A(n20189), .ZN(n20215) );
  OAI22_X1 U23086 ( .A1(n20257), .A2(n20753), .B1(n20738), .B2(n20215), .ZN(
        n20187) );
  INV_X1 U23087 ( .A(n20187), .ZN(n20196) );
  NAND2_X1 U23088 ( .A1(n20257), .A2(n20221), .ZN(n20188) );
  AOI21_X1 U23089 ( .B1(n20188), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20744), 
        .ZN(n20192) );
  OR2_X1 U23090 ( .A1(n20224), .A2(n20673), .ZN(n20193) );
  NOR2_X1 U23091 ( .A1(n20189), .A2(n20589), .ZN(n20190) );
  AOI21_X1 U23092 ( .B1(n20192), .B2(n20193), .A(n20190), .ZN(n20191) );
  OR2_X1 U23093 ( .A1(n20501), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20342) );
  NAND2_X1 U23094 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20342), .ZN(n20349) );
  NAND3_X1 U23095 ( .A1(n20504), .A2(n20191), .A3(n20349), .ZN(n20218) );
  INV_X1 U23096 ( .A(n20739), .ZN(n20596) );
  INV_X1 U23097 ( .A(n20192), .ZN(n20194) );
  OAI22_X1 U23098 ( .A1(n20194), .A2(n20193), .B1(n20507), .B2(n20342), .ZN(
        n20217) );
  AOI22_X1 U23099 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20218), .B1(
        n20596), .B2(n20217), .ZN(n20195) );
  OAI211_X1 U23100 ( .C1(n20692), .C2(n20221), .A(n20196), .B(n20195), .ZN(
        P1_U3049) );
  OAI22_X1 U23101 ( .A1(n20257), .A2(n20760), .B1(n20215), .B2(n20754), .ZN(
        n20197) );
  INV_X1 U23102 ( .A(n20197), .ZN(n20199) );
  INV_X1 U23103 ( .A(n20755), .ZN(n20600) );
  AOI22_X1 U23104 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20218), .B1(
        n20600), .B2(n20217), .ZN(n20198) );
  OAI211_X1 U23105 ( .C1(n20697), .C2(n20221), .A(n20199), .B(n20198), .ZN(
        P1_U3050) );
  OAI22_X1 U23106 ( .A1(n20221), .A2(n20702), .B1(n20215), .B2(n20761), .ZN(
        n20200) );
  INV_X1 U23107 ( .A(n20200), .ZN(n20202) );
  INV_X1 U23108 ( .A(n20762), .ZN(n20604) );
  AOI22_X1 U23109 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20218), .B1(
        n20604), .B2(n20217), .ZN(n20201) );
  OAI211_X1 U23110 ( .C1(n20767), .C2(n20257), .A(n20202), .B(n20201), .ZN(
        P1_U3051) );
  OAI22_X1 U23111 ( .A1(n20257), .A2(n20774), .B1(n20215), .B2(n20768), .ZN(
        n20203) );
  INV_X1 U23112 ( .A(n20203), .ZN(n20205) );
  INV_X1 U23113 ( .A(n20769), .ZN(n20608) );
  AOI22_X1 U23114 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20218), .B1(
        n20608), .B2(n20217), .ZN(n20204) );
  OAI211_X1 U23115 ( .C1(n20707), .C2(n20221), .A(n20205), .B(n20204), .ZN(
        P1_U3052) );
  OAI22_X1 U23116 ( .A1(n20221), .A2(n20712), .B1(n20215), .B2(n20775), .ZN(
        n20206) );
  INV_X1 U23117 ( .A(n20206), .ZN(n20208) );
  AOI22_X1 U23118 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20218), .B1(
        n20612), .B2(n20217), .ZN(n20207) );
  OAI211_X1 U23119 ( .C1(n20781), .C2(n20257), .A(n20208), .B(n20207), .ZN(
        P1_U3053) );
  OAI22_X1 U23120 ( .A1(n20257), .A2(n20788), .B1(n20215), .B2(n20782), .ZN(
        n20209) );
  INV_X1 U23121 ( .A(n20209), .ZN(n20211) );
  AOI22_X1 U23122 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20218), .B1(
        n20616), .B2(n20217), .ZN(n20210) );
  OAI211_X1 U23123 ( .C1(n20717), .C2(n20221), .A(n20211), .B(n20210), .ZN(
        P1_U3054) );
  OAI22_X1 U23124 ( .A1(n20257), .A2(n20795), .B1(n20215), .B2(n20789), .ZN(
        n20212) );
  INV_X1 U23125 ( .A(n20212), .ZN(n20214) );
  AOI22_X1 U23126 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20218), .B1(
        n20620), .B2(n20217), .ZN(n20213) );
  OAI211_X1 U23127 ( .C1(n20722), .C2(n20221), .A(n20214), .B(n20213), .ZN(
        P1_U3055) );
  OAI22_X1 U23128 ( .A1(n20257), .A2(n20912), .B1(n20215), .B2(n20908), .ZN(
        n20216) );
  INV_X1 U23129 ( .A(n20216), .ZN(n20220) );
  AOI22_X1 U23130 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20218), .B1(
        n20626), .B2(n20217), .ZN(n20219) );
  OAI211_X1 U23131 ( .C1(n20910), .C2(n20221), .A(n20220), .B(n20219), .ZN(
        P1_U3056) );
  NAND2_X1 U23132 ( .A1(n20734), .A2(n20222), .ZN(n20256) );
  OAI22_X1 U23133 ( .A1(n20304), .A2(n20753), .B1(n20738), .B2(n20256), .ZN(
        n20223) );
  INV_X1 U23134 ( .A(n20223), .ZN(n20237) );
  INV_X1 U23135 ( .A(n20224), .ZN(n20228) );
  AND2_X1 U23136 ( .A1(n20226), .A2(n20225), .ZN(n20539) );
  INV_X1 U23137 ( .A(n20256), .ZN(n20227) );
  AOI21_X1 U23138 ( .B1(n20228), .B2(n20539), .A(n20227), .ZN(n20235) );
  OR2_X1 U23139 ( .A1(n20229), .A2(n20742), .ZN(n20230) );
  AOI22_X1 U23140 ( .A1(n20235), .A2(n20232), .B1(n20744), .B2(n20233), .ZN(
        n20231) );
  NAND2_X1 U23141 ( .A1(n20748), .A2(n20231), .ZN(n20260) );
  INV_X1 U23142 ( .A(n20232), .ZN(n20234) );
  OAI22_X1 U23143 ( .A1(n20235), .A2(n20234), .B1(n20383), .B2(n20233), .ZN(
        n20259) );
  AOI22_X1 U23144 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20260), .B1(
        n20596), .B2(n20259), .ZN(n20236) );
  OAI211_X1 U23145 ( .C1(n20692), .C2(n20257), .A(n20237), .B(n20236), .ZN(
        P1_U3057) );
  OAI22_X1 U23146 ( .A1(n20257), .A2(n20697), .B1(n20754), .B2(n20256), .ZN(
        n20238) );
  INV_X1 U23147 ( .A(n20238), .ZN(n20240) );
  AOI22_X1 U23148 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20260), .B1(
        n20600), .B2(n20259), .ZN(n20239) );
  OAI211_X1 U23149 ( .C1(n20760), .C2(n20304), .A(n20240), .B(n20239), .ZN(
        P1_U3058) );
  OAI22_X1 U23150 ( .A1(n20257), .A2(n20702), .B1(n20256), .B2(n20761), .ZN(
        n20241) );
  INV_X1 U23151 ( .A(n20241), .ZN(n20243) );
  AOI22_X1 U23152 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20260), .B1(
        n20604), .B2(n20259), .ZN(n20242) );
  OAI211_X1 U23153 ( .C1(n20767), .C2(n20304), .A(n20243), .B(n20242), .ZN(
        P1_U3059) );
  OAI22_X1 U23154 ( .A1(n20257), .A2(n20707), .B1(n20768), .B2(n20256), .ZN(
        n20244) );
  INV_X1 U23155 ( .A(n20244), .ZN(n20246) );
  AOI22_X1 U23156 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20260), .B1(
        n20608), .B2(n20259), .ZN(n20245) );
  OAI211_X1 U23157 ( .C1(n20774), .C2(n20304), .A(n20246), .B(n20245), .ZN(
        P1_U3060) );
  OAI22_X1 U23158 ( .A1(n20304), .A2(n20781), .B1(n20256), .B2(n20775), .ZN(
        n20247) );
  INV_X1 U23159 ( .A(n20247), .ZN(n20249) );
  AOI22_X1 U23160 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20260), .B1(
        n20612), .B2(n20259), .ZN(n20248) );
  OAI211_X1 U23161 ( .C1(n20712), .C2(n20257), .A(n20249), .B(n20248), .ZN(
        P1_U3061) );
  OAI22_X1 U23162 ( .A1(n20304), .A2(n20788), .B1(n20782), .B2(n20256), .ZN(
        n20250) );
  INV_X1 U23163 ( .A(n20250), .ZN(n20252) );
  AOI22_X1 U23164 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20260), .B1(
        n20616), .B2(n20259), .ZN(n20251) );
  OAI211_X1 U23165 ( .C1(n20717), .C2(n20257), .A(n20252), .B(n20251), .ZN(
        P1_U3062) );
  OAI22_X1 U23166 ( .A1(n20304), .A2(n20795), .B1(n20789), .B2(n20256), .ZN(
        n20253) );
  INV_X1 U23167 ( .A(n20253), .ZN(n20255) );
  AOI22_X1 U23168 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20260), .B1(
        n20620), .B2(n20259), .ZN(n20254) );
  OAI211_X1 U23169 ( .C1(n20722), .C2(n20257), .A(n20255), .B(n20254), .ZN(
        P1_U3063) );
  OAI22_X1 U23170 ( .A1(n20257), .A2(n20910), .B1(n20908), .B2(n20256), .ZN(
        n20258) );
  INV_X1 U23171 ( .A(n20258), .ZN(n20262) );
  AOI22_X1 U23172 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20260), .B1(
        n20626), .B2(n20259), .ZN(n20261) );
  OAI211_X1 U23173 ( .C1(n20912), .C2(n20304), .A(n20262), .B(n20261), .ZN(
        P1_U3064) );
  OR2_X1 U23174 ( .A1(n13122), .A2(n20263), .ZN(n20382) );
  NAND2_X1 U23175 ( .A1(n20673), .A2(n20741), .ZN(n20264) );
  OR2_X1 U23176 ( .A1(n20382), .A2(n20264), .ZN(n20267) );
  INV_X1 U23177 ( .A(n20592), .ZN(n20677) );
  NAND2_X1 U23178 ( .A1(n20265), .A2(n20677), .ZN(n20266) );
  OR2_X1 U23179 ( .A1(n20583), .A2(n20344), .ZN(n20298) );
  OAI22_X1 U23180 ( .A1(n20739), .A2(n20297), .B1(n20738), .B2(n20298), .ZN(
        n20268) );
  INV_X1 U23181 ( .A(n20268), .ZN(n20277) );
  INV_X1 U23182 ( .A(n20298), .ZN(n20275) );
  INV_X1 U23183 ( .A(n20382), .ZN(n20271) );
  AOI21_X1 U23184 ( .B1(n20304), .B2(n20340), .A(n20466), .ZN(n20270) );
  AOI21_X1 U23185 ( .B1(n20271), .B2(n20673), .A(n20270), .ZN(n20272) );
  NOR2_X1 U23186 ( .A1(n20272), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20274) );
  AOI22_X1 U23187 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20301), .B1(
        n20300), .B2(n20689), .ZN(n20276) );
  OAI211_X1 U23188 ( .C1(n20692), .C2(n20304), .A(n20277), .B(n20276), .ZN(
        P1_U3065) );
  OAI22_X1 U23189 ( .A1(n20755), .A2(n20297), .B1(n20754), .B2(n20298), .ZN(
        n20278) );
  INV_X1 U23190 ( .A(n20278), .ZN(n20280) );
  AOI22_X1 U23191 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20301), .B1(
        n20300), .B2(n20694), .ZN(n20279) );
  OAI211_X1 U23192 ( .C1(n20697), .C2(n20304), .A(n20280), .B(n20279), .ZN(
        P1_U3066) );
  OAI22_X1 U23193 ( .A1(n20762), .A2(n20297), .B1(n20761), .B2(n20298), .ZN(
        n20281) );
  INV_X1 U23194 ( .A(n20281), .ZN(n20283) );
  INV_X1 U23195 ( .A(n20304), .ZN(n20288) );
  AOI22_X1 U23196 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20301), .B1(
        n20288), .B2(n20764), .ZN(n20282) );
  OAI211_X1 U23197 ( .C1(n20767), .C2(n20340), .A(n20283), .B(n20282), .ZN(
        P1_U3067) );
  OAI22_X1 U23198 ( .A1(n20769), .A2(n20297), .B1(n20768), .B2(n20298), .ZN(
        n20284) );
  INV_X1 U23199 ( .A(n20284), .ZN(n20286) );
  AOI22_X1 U23200 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20301), .B1(
        n20300), .B2(n20704), .ZN(n20285) );
  OAI211_X1 U23201 ( .C1(n20707), .C2(n20304), .A(n20286), .B(n20285), .ZN(
        P1_U3068) );
  OAI22_X1 U23202 ( .A1(n20776), .A2(n20297), .B1(n20775), .B2(n20298), .ZN(
        n20287) );
  INV_X1 U23203 ( .A(n20287), .ZN(n20290) );
  AOI22_X1 U23204 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20301), .B1(
        n20288), .B2(n20778), .ZN(n20289) );
  OAI211_X1 U23205 ( .C1(n20781), .C2(n20340), .A(n20290), .B(n20289), .ZN(
        P1_U3069) );
  OAI22_X1 U23206 ( .A1(n20783), .A2(n20297), .B1(n20782), .B2(n20298), .ZN(
        n20291) );
  INV_X1 U23207 ( .A(n20291), .ZN(n20293) );
  INV_X1 U23208 ( .A(n20788), .ZN(n20714) );
  AOI22_X1 U23209 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20301), .B1(
        n20300), .B2(n20714), .ZN(n20292) );
  OAI211_X1 U23210 ( .C1(n20717), .C2(n20304), .A(n20293), .B(n20292), .ZN(
        P1_U3070) );
  OAI22_X1 U23211 ( .A1(n20790), .A2(n20297), .B1(n20789), .B2(n20298), .ZN(
        n20294) );
  INV_X1 U23212 ( .A(n20294), .ZN(n20296) );
  AOI22_X1 U23213 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20301), .B1(
        n20300), .B2(n9633), .ZN(n20295) );
  OAI211_X1 U23214 ( .C1(n20722), .C2(n20304), .A(n20296), .B(n20295), .ZN(
        P1_U3071) );
  OAI22_X1 U23215 ( .A1(n20908), .A2(n20298), .B1(n20297), .B2(n20913), .ZN(
        n20299) );
  INV_X1 U23216 ( .A(n20299), .ZN(n20303) );
  INV_X1 U23217 ( .A(n20912), .ZN(n20726) );
  AOI22_X1 U23218 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20301), .B1(
        n20300), .B2(n20726), .ZN(n20302) );
  OAI211_X1 U23219 ( .C1(n20910), .C2(n20304), .A(n20303), .B(n20302), .ZN(
        P1_U3072) );
  OR2_X1 U23220 ( .A1(n20382), .A2(n20634), .ZN(n20306) );
  NOR2_X1 U23221 ( .A1(n20344), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20313) );
  INV_X1 U23222 ( .A(n20313), .ZN(n20305) );
  OR2_X1 U23223 ( .A1(n20635), .A2(n20305), .ZN(n20335) );
  NAND2_X1 U23224 ( .A1(n20306), .A2(n20335), .ZN(n20310) );
  NAND2_X1 U23225 ( .A1(n20310), .A2(n20741), .ZN(n20308) );
  NAND2_X1 U23226 ( .A1(n20313), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20307) );
  AND2_X1 U23227 ( .A1(n20308), .A2(n20307), .ZN(n20334) );
  OAI22_X1 U23228 ( .A1(n20739), .A2(n20334), .B1(n20738), .B2(n20335), .ZN(
        n20309) );
  INV_X1 U23229 ( .A(n20309), .ZN(n20315) );
  INV_X1 U23230 ( .A(n20585), .ZN(n20642) );
  INV_X1 U23231 ( .A(n20310), .ZN(n20311) );
  OAI21_X1 U23232 ( .B1(n20390), .B2(n20642), .A(n20311), .ZN(n20312) );
  OAI211_X1 U23233 ( .C1(n20741), .C2(n20313), .A(n20748), .B(n20312), .ZN(
        n20337) );
  AOI22_X1 U23234 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20337), .B1(
        n20370), .B2(n20689), .ZN(n20314) );
  OAI211_X1 U23235 ( .C1(n20692), .C2(n20340), .A(n20315), .B(n20314), .ZN(
        P1_U3073) );
  OAI22_X1 U23236 ( .A1(n20755), .A2(n20334), .B1(n20754), .B2(n20335), .ZN(
        n20316) );
  INV_X1 U23237 ( .A(n20316), .ZN(n20318) );
  AOI22_X1 U23238 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20337), .B1(
        n20370), .B2(n20694), .ZN(n20317) );
  OAI211_X1 U23239 ( .C1(n20697), .C2(n20340), .A(n20318), .B(n20317), .ZN(
        P1_U3074) );
  OAI22_X1 U23240 ( .A1(n20762), .A2(n20334), .B1(n20761), .B2(n20335), .ZN(
        n20319) );
  INV_X1 U23241 ( .A(n20319), .ZN(n20321) );
  AOI22_X1 U23242 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20337), .B1(
        n20370), .B2(n20699), .ZN(n20320) );
  OAI211_X1 U23243 ( .C1(n20702), .C2(n20340), .A(n20321), .B(n20320), .ZN(
        P1_U3075) );
  OAI22_X1 U23244 ( .A1(n20769), .A2(n20334), .B1(n20768), .B2(n20335), .ZN(
        n20322) );
  INV_X1 U23245 ( .A(n20322), .ZN(n20324) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20337), .B1(
        n20370), .B2(n20704), .ZN(n20323) );
  OAI211_X1 U23247 ( .C1(n20707), .C2(n20340), .A(n20324), .B(n20323), .ZN(
        P1_U3076) );
  OAI22_X1 U23248 ( .A1(n20776), .A2(n20334), .B1(n20775), .B2(n20335), .ZN(
        n20325) );
  INV_X1 U23249 ( .A(n20325), .ZN(n20327) );
  INV_X1 U23250 ( .A(n20781), .ZN(n20709) );
  AOI22_X1 U23251 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20337), .B1(
        n20370), .B2(n20709), .ZN(n20326) );
  OAI211_X1 U23252 ( .C1(n20712), .C2(n20340), .A(n20327), .B(n20326), .ZN(
        P1_U3077) );
  OAI22_X1 U23253 ( .A1(n20783), .A2(n20334), .B1(n20782), .B2(n20335), .ZN(
        n20328) );
  INV_X1 U23254 ( .A(n20328), .ZN(n20330) );
  AOI22_X1 U23255 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20337), .B1(
        n20370), .B2(n20714), .ZN(n20329) );
  OAI211_X1 U23256 ( .C1(n20717), .C2(n20340), .A(n20330), .B(n20329), .ZN(
        P1_U3078) );
  OAI22_X1 U23257 ( .A1(n20790), .A2(n20334), .B1(n20789), .B2(n20335), .ZN(
        n20331) );
  INV_X1 U23258 ( .A(n20331), .ZN(n20333) );
  AOI22_X1 U23259 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20337), .B1(
        n20370), .B2(n9633), .ZN(n20332) );
  OAI211_X1 U23260 ( .C1(n20722), .C2(n20340), .A(n20333), .B(n20332), .ZN(
        P1_U3079) );
  OAI22_X1 U23261 ( .A1(n20908), .A2(n20335), .B1(n20334), .B2(n20913), .ZN(
        n20336) );
  INV_X1 U23262 ( .A(n20336), .ZN(n20339) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20337), .B1(
        n20370), .B2(n20726), .ZN(n20338) );
  OAI211_X1 U23264 ( .C1(n20910), .C2(n20340), .A(n20339), .B(n20338), .ZN(
        P1_U3080) );
  NAND3_X1 U23265 ( .A1(n20368), .A2(n20374), .A3(n20741), .ZN(n20341) );
  NAND2_X1 U23266 ( .A1(n20341), .A2(n20585), .ZN(n20348) );
  NOR2_X1 U23267 ( .A1(n20382), .A2(n20673), .ZN(n20346) );
  INV_X1 U23268 ( .A(n20342), .ZN(n20343) );
  AOI22_X1 U23269 ( .A1(n20348), .A2(n20346), .B1(n20343), .B2(n20677), .ZN(
        n20379) );
  NOR2_X1 U23270 ( .A1(n20746), .A2(n20344), .ZN(n20391) );
  NAND2_X1 U23271 ( .A1(n20635), .A2(n20391), .ZN(n20373) );
  OAI22_X1 U23272 ( .A1(n20692), .A2(n20374), .B1(n20738), .B2(n20373), .ZN(
        n20345) );
  INV_X1 U23273 ( .A(n20345), .ZN(n20352) );
  INV_X1 U23274 ( .A(n20346), .ZN(n20347) );
  AOI22_X1 U23275 ( .A1(n20348), .A2(n20347), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20373), .ZN(n20350) );
  NAND3_X1 U23276 ( .A1(n20686), .A2(n20350), .A3(n20349), .ZN(n20376) );
  AOI22_X1 U23277 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20376), .B1(
        n20415), .B2(n20689), .ZN(n20351) );
  OAI211_X1 U23278 ( .C1(n20379), .C2(n20739), .A(n20352), .B(n20351), .ZN(
        P1_U3081) );
  OAI22_X1 U23279 ( .A1(n20697), .A2(n20374), .B1(n20754), .B2(n20373), .ZN(
        n20353) );
  INV_X1 U23280 ( .A(n20353), .ZN(n20355) );
  AOI22_X1 U23281 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20376), .B1(
        n20415), .B2(n20694), .ZN(n20354) );
  OAI211_X1 U23282 ( .C1(n20379), .C2(n20755), .A(n20355), .B(n20354), .ZN(
        P1_U3082) );
  OAI22_X1 U23283 ( .A1(n20702), .A2(n20374), .B1(n20761), .B2(n20373), .ZN(
        n20356) );
  INV_X1 U23284 ( .A(n20356), .ZN(n20358) );
  AOI22_X1 U23285 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20376), .B1(
        n20415), .B2(n20699), .ZN(n20357) );
  OAI211_X1 U23286 ( .C1(n20379), .C2(n20762), .A(n20358), .B(n20357), .ZN(
        P1_U3083) );
  OAI22_X1 U23287 ( .A1(n20707), .A2(n20374), .B1(n20768), .B2(n20373), .ZN(
        n20359) );
  INV_X1 U23288 ( .A(n20359), .ZN(n20361) );
  AOI22_X1 U23289 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20376), .B1(
        n20415), .B2(n20704), .ZN(n20360) );
  OAI211_X1 U23290 ( .C1(n20379), .C2(n20769), .A(n20361), .B(n20360), .ZN(
        P1_U3084) );
  OAI22_X1 U23291 ( .A1(n20781), .A2(n20368), .B1(n20775), .B2(n20373), .ZN(
        n20362) );
  INV_X1 U23292 ( .A(n20362), .ZN(n20364) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20376), .B1(
        n20370), .B2(n20778), .ZN(n20363) );
  OAI211_X1 U23294 ( .C1(n20379), .C2(n20776), .A(n20364), .B(n20363), .ZN(
        P1_U3085) );
  OAI22_X1 U23295 ( .A1(n20717), .A2(n20374), .B1(n20782), .B2(n20373), .ZN(
        n20365) );
  INV_X1 U23296 ( .A(n20365), .ZN(n20367) );
  AOI22_X1 U23297 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20376), .B1(
        n20415), .B2(n20714), .ZN(n20366) );
  OAI211_X1 U23298 ( .C1(n20379), .C2(n20783), .A(n20367), .B(n20366), .ZN(
        P1_U3086) );
  OAI22_X1 U23299 ( .A1(n20795), .A2(n20368), .B1(n20789), .B2(n20373), .ZN(
        n20369) );
  INV_X1 U23300 ( .A(n20369), .ZN(n20372) );
  INV_X1 U23301 ( .A(n20722), .ZN(n20792) );
  AOI22_X1 U23302 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20376), .B1(
        n20370), .B2(n20792), .ZN(n20371) );
  OAI211_X1 U23303 ( .C1(n20379), .C2(n20790), .A(n20372), .B(n20371), .ZN(
        P1_U3087) );
  OAI22_X1 U23304 ( .A1(n20910), .A2(n20374), .B1(n20908), .B2(n20373), .ZN(
        n20375) );
  INV_X1 U23305 ( .A(n20375), .ZN(n20378) );
  AOI22_X1 U23306 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20376), .B1(
        n20415), .B2(n20726), .ZN(n20377) );
  OAI211_X1 U23307 ( .C1(n20379), .C2(n20913), .A(n20378), .B(n20377), .ZN(
        P1_U3088) );
  INV_X1 U23308 ( .A(n20390), .ZN(n20381) );
  INV_X1 U23309 ( .A(n20551), .ZN(n20380) );
  INV_X1 U23310 ( .A(n20539), .ZN(n20731) );
  OAI21_X1 U23311 ( .B1(n20382), .B2(n20731), .A(n20413), .ZN(n20386) );
  INV_X1 U23312 ( .A(n20391), .ZN(n20384) );
  NOR2_X1 U23313 ( .A1(n20384), .A2(n20383), .ZN(n20385) );
  AOI21_X1 U23314 ( .B1(n20386), .B2(n20741), .A(n20385), .ZN(n20412) );
  OAI22_X1 U23315 ( .A1(n20739), .A2(n20412), .B1(n20738), .B2(n20413), .ZN(
        n20387) );
  INV_X1 U23316 ( .A(n20387), .ZN(n20393) );
  INV_X1 U23317 ( .A(n20388), .ZN(n20389) );
  NOR2_X1 U23318 ( .A1(n20390), .A2(n20389), .ZN(n20876) );
  OAI21_X1 U23319 ( .B1(n20391), .B2(n20876), .A(n20748), .ZN(n20416) );
  INV_X1 U23320 ( .A(n20692), .ZN(n20750) );
  AOI22_X1 U23321 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20750), .ZN(n20392) );
  OAI211_X1 U23322 ( .C1(n20753), .C2(n20457), .A(n20393), .B(n20392), .ZN(
        P1_U3089) );
  OAI22_X1 U23323 ( .A1(n20755), .A2(n20412), .B1(n20754), .B2(n20413), .ZN(
        n20394) );
  INV_X1 U23324 ( .A(n20394), .ZN(n20396) );
  AOI22_X1 U23325 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20757), .ZN(n20395) );
  OAI211_X1 U23326 ( .C1(n20760), .C2(n20457), .A(n20396), .B(n20395), .ZN(
        P1_U3090) );
  OAI22_X1 U23327 ( .A1(n20762), .A2(n20412), .B1(n20761), .B2(n20413), .ZN(
        n20397) );
  INV_X1 U23328 ( .A(n20397), .ZN(n20399) );
  AOI22_X1 U23329 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20764), .ZN(n20398) );
  OAI211_X1 U23330 ( .C1(n20767), .C2(n20457), .A(n20399), .B(n20398), .ZN(
        P1_U3091) );
  OAI22_X1 U23331 ( .A1(n20769), .A2(n20412), .B1(n20768), .B2(n20413), .ZN(
        n20400) );
  INV_X1 U23332 ( .A(n20400), .ZN(n20402) );
  INV_X1 U23333 ( .A(n20707), .ZN(n20771) );
  AOI22_X1 U23334 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20771), .ZN(n20401) );
  OAI211_X1 U23335 ( .C1(n20774), .C2(n20457), .A(n20402), .B(n20401), .ZN(
        P1_U3092) );
  OAI22_X1 U23336 ( .A1(n20776), .A2(n20412), .B1(n20775), .B2(n20413), .ZN(
        n20403) );
  INV_X1 U23337 ( .A(n20403), .ZN(n20405) );
  AOI22_X1 U23338 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20778), .ZN(n20404) );
  OAI211_X1 U23339 ( .C1(n20781), .C2(n20457), .A(n20405), .B(n20404), .ZN(
        P1_U3093) );
  OAI22_X1 U23340 ( .A1(n20783), .A2(n20412), .B1(n20782), .B2(n20413), .ZN(
        n20406) );
  INV_X1 U23341 ( .A(n20406), .ZN(n20408) );
  AOI22_X1 U23342 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20785), .ZN(n20407) );
  OAI211_X1 U23343 ( .C1(n20788), .C2(n20457), .A(n20408), .B(n20407), .ZN(
        P1_U3094) );
  OAI22_X1 U23344 ( .A1(n20790), .A2(n20412), .B1(n20789), .B2(n20413), .ZN(
        n20409) );
  INV_X1 U23345 ( .A(n20409), .ZN(n20411) );
  AOI22_X1 U23346 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20792), .ZN(n20410) );
  OAI211_X1 U23347 ( .C1(n20795), .C2(n20457), .A(n20411), .B(n20410), .ZN(
        P1_U3095) );
  OAI22_X1 U23348 ( .A1(n20908), .A2(n20413), .B1(n20412), .B2(n20913), .ZN(
        n20414) );
  INV_X1 U23349 ( .A(n20414), .ZN(n20418) );
  AOI22_X1 U23350 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20416), .B1(
        n20415), .B2(n20799), .ZN(n20417) );
  OAI211_X1 U23351 ( .C1(n20912), .C2(n20457), .A(n20418), .B(n20417), .ZN(
        P1_U3096) );
  AND2_X1 U23352 ( .A1(n13145), .A2(n13122), .ZN(n20540) );
  NAND2_X1 U23353 ( .A1(n20419), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20537) );
  OR2_X1 U23354 ( .A1(n20583), .A2(n20537), .ZN(n20452) );
  INV_X1 U23355 ( .A(n20452), .ZN(n20430) );
  AOI21_X1 U23356 ( .B1(n20540), .B2(n20673), .A(n20430), .ZN(n20427) );
  OR2_X1 U23357 ( .A1(n20427), .A2(n20744), .ZN(n20422) );
  NAND2_X1 U23358 ( .A1(n20420), .A2(n20501), .ZN(n20593) );
  OR2_X1 U23359 ( .A1(n20593), .A2(n20507), .ZN(n20421) );
  OAI22_X1 U23360 ( .A1(n20739), .A2(n20451), .B1(n20738), .B2(n20452), .ZN(
        n20423) );
  INV_X1 U23361 ( .A(n20423), .ZN(n20432) );
  INV_X1 U23362 ( .A(n20424), .ZN(n20425) );
  INV_X1 U23363 ( .A(n20457), .ZN(n20426) );
  OAI21_X1 U23364 ( .B1(n20493), .B2(n20426), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20428) );
  NAND2_X1 U23365 ( .A1(n20428), .A2(n20427), .ZN(n20429) );
  AOI22_X1 U23366 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20454), .B1(
        n20493), .B2(n20689), .ZN(n20431) );
  OAI211_X1 U23367 ( .C1(n20692), .C2(n20457), .A(n20432), .B(n20431), .ZN(
        P1_U3097) );
  OAI22_X1 U23368 ( .A1(n20755), .A2(n20451), .B1(n20754), .B2(n20452), .ZN(
        n20433) );
  INV_X1 U23369 ( .A(n20433), .ZN(n20435) );
  AOI22_X1 U23370 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20454), .B1(
        n20493), .B2(n20694), .ZN(n20434) );
  OAI211_X1 U23371 ( .C1(n20697), .C2(n20457), .A(n20435), .B(n20434), .ZN(
        P1_U3098) );
  OAI22_X1 U23372 ( .A1(n20762), .A2(n20451), .B1(n20761), .B2(n20452), .ZN(
        n20436) );
  INV_X1 U23373 ( .A(n20436), .ZN(n20438) );
  AOI22_X1 U23374 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20454), .B1(
        n20493), .B2(n20699), .ZN(n20437) );
  OAI211_X1 U23375 ( .C1(n20702), .C2(n20457), .A(n20438), .B(n20437), .ZN(
        P1_U3099) );
  OAI22_X1 U23376 ( .A1(n20769), .A2(n20451), .B1(n20768), .B2(n20452), .ZN(
        n20439) );
  INV_X1 U23377 ( .A(n20439), .ZN(n20441) );
  AOI22_X1 U23378 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20454), .B1(
        n20493), .B2(n20704), .ZN(n20440) );
  OAI211_X1 U23379 ( .C1(n20707), .C2(n20457), .A(n20441), .B(n20440), .ZN(
        P1_U3100) );
  OAI22_X1 U23380 ( .A1(n20776), .A2(n20451), .B1(n20775), .B2(n20452), .ZN(
        n20442) );
  INV_X1 U23381 ( .A(n20442), .ZN(n20444) );
  AOI22_X1 U23382 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20454), .B1(
        n20493), .B2(n20709), .ZN(n20443) );
  OAI211_X1 U23383 ( .C1(n20712), .C2(n20457), .A(n20444), .B(n20443), .ZN(
        P1_U3101) );
  OAI22_X1 U23384 ( .A1(n20783), .A2(n20451), .B1(n20782), .B2(n20452), .ZN(
        n20445) );
  INV_X1 U23385 ( .A(n20445), .ZN(n20447) );
  AOI22_X1 U23386 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20454), .B1(
        n20493), .B2(n20714), .ZN(n20446) );
  OAI211_X1 U23387 ( .C1(n20717), .C2(n20457), .A(n20447), .B(n20446), .ZN(
        P1_U3102) );
  OAI22_X1 U23388 ( .A1(n20790), .A2(n20451), .B1(n20789), .B2(n20452), .ZN(
        n20448) );
  INV_X1 U23389 ( .A(n20448), .ZN(n20450) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20454), .B1(
        n20493), .B2(n9633), .ZN(n20449) );
  OAI211_X1 U23391 ( .C1(n20722), .C2(n20457), .A(n20450), .B(n20449), .ZN(
        P1_U3103) );
  OAI22_X1 U23392 ( .A1(n20908), .A2(n20452), .B1(n20451), .B2(n20913), .ZN(
        n20453) );
  INV_X1 U23393 ( .A(n20453), .ZN(n20456) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20454), .B1(
        n20493), .B2(n20726), .ZN(n20455) );
  OAI211_X1 U23395 ( .C1(n20910), .C2(n20457), .A(n20456), .B(n20455), .ZN(
        P1_U3104) );
  INV_X1 U23396 ( .A(n20634), .ZN(n20458) );
  NAND2_X1 U23397 ( .A1(n20540), .A2(n20458), .ZN(n20460) );
  NOR2_X1 U23398 ( .A1(n20537), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20468) );
  INV_X1 U23399 ( .A(n20468), .ZN(n20459) );
  OR2_X1 U23400 ( .A1(n20635), .A2(n20459), .ZN(n20491) );
  NAND2_X1 U23401 ( .A1(n20460), .A2(n20491), .ZN(n20464) );
  NAND2_X1 U23402 ( .A1(n20464), .A2(n20741), .ZN(n20462) );
  NAND2_X1 U23403 ( .A1(n20468), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20461) );
  AND2_X1 U23404 ( .A1(n20462), .A2(n20461), .ZN(n20490) );
  OAI22_X1 U23405 ( .A1(n20739), .A2(n20490), .B1(n20738), .B2(n20491), .ZN(
        n20463) );
  INV_X1 U23406 ( .A(n20463), .ZN(n20470) );
  INV_X1 U23407 ( .A(n20464), .ZN(n20465) );
  OAI211_X1 U23408 ( .C1(n20552), .C2(n20466), .A(n20741), .B(n20465), .ZN(
        n20467) );
  OAI211_X1 U23409 ( .C1(n20741), .C2(n20468), .A(n20748), .B(n20467), .ZN(
        n20494) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20494), .B1(
        n20499), .B2(n20689), .ZN(n20469) );
  OAI211_X1 U23411 ( .C1(n20692), .C2(n20480), .A(n20470), .B(n20469), .ZN(
        P1_U3105) );
  OAI22_X1 U23412 ( .A1(n20755), .A2(n20490), .B1(n20754), .B2(n20491), .ZN(
        n20471) );
  INV_X1 U23413 ( .A(n20471), .ZN(n20473) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20494), .B1(
        n20499), .B2(n20694), .ZN(n20472) );
  OAI211_X1 U23415 ( .C1(n20697), .C2(n20480), .A(n20473), .B(n20472), .ZN(
        P1_U3106) );
  OAI22_X1 U23416 ( .A1(n20762), .A2(n20490), .B1(n20761), .B2(n20491), .ZN(
        n20474) );
  INV_X1 U23417 ( .A(n20474), .ZN(n20476) );
  AOI22_X1 U23418 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20764), .ZN(n20475) );
  OAI211_X1 U23419 ( .C1(n20767), .C2(n20536), .A(n20476), .B(n20475), .ZN(
        P1_U3107) );
  OAI22_X1 U23420 ( .A1(n20769), .A2(n20490), .B1(n20768), .B2(n20491), .ZN(
        n20477) );
  INV_X1 U23421 ( .A(n20477), .ZN(n20479) );
  AOI22_X1 U23422 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20494), .B1(
        n20499), .B2(n20704), .ZN(n20478) );
  OAI211_X1 U23423 ( .C1(n20707), .C2(n20480), .A(n20479), .B(n20478), .ZN(
        P1_U3108) );
  OAI22_X1 U23424 ( .A1(n20776), .A2(n20490), .B1(n20775), .B2(n20491), .ZN(
        n20481) );
  INV_X1 U23425 ( .A(n20481), .ZN(n20483) );
  AOI22_X1 U23426 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20778), .ZN(n20482) );
  OAI211_X1 U23427 ( .C1(n20781), .C2(n20536), .A(n20483), .B(n20482), .ZN(
        P1_U3109) );
  OAI22_X1 U23428 ( .A1(n20783), .A2(n20490), .B1(n20782), .B2(n20491), .ZN(
        n20484) );
  INV_X1 U23429 ( .A(n20484), .ZN(n20486) );
  AOI22_X1 U23430 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20785), .ZN(n20485) );
  OAI211_X1 U23431 ( .C1(n20788), .C2(n20536), .A(n20486), .B(n20485), .ZN(
        P1_U3110) );
  OAI22_X1 U23432 ( .A1(n20790), .A2(n20490), .B1(n20789), .B2(n20491), .ZN(
        n20487) );
  INV_X1 U23433 ( .A(n20487), .ZN(n20489) );
  AOI22_X1 U23434 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20792), .ZN(n20488) );
  OAI211_X1 U23435 ( .C1(n20795), .C2(n20536), .A(n20489), .B(n20488), .ZN(
        P1_U3111) );
  OAI22_X1 U23436 ( .A1(n20908), .A2(n20491), .B1(n20490), .B2(n20913), .ZN(
        n20492) );
  INV_X1 U23437 ( .A(n20492), .ZN(n20496) );
  AOI22_X1 U23438 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20494), .B1(
        n20493), .B2(n20799), .ZN(n20495) );
  OAI211_X1 U23439 ( .C1(n20912), .C2(n20536), .A(n20496), .B(n20495), .ZN(
        P1_U3112) );
  NOR2_X1 U23440 ( .A1(n20746), .A2(n20537), .ZN(n20550) );
  INV_X1 U23441 ( .A(n20550), .ZN(n20497) );
  NOR2_X1 U23442 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20497), .ZN(
        n20502) );
  INV_X1 U23443 ( .A(n20502), .ZN(n20530) );
  OAI22_X1 U23444 ( .A1(n20581), .A2(n20753), .B1(n20738), .B2(n20530), .ZN(
        n20498) );
  INV_X1 U23445 ( .A(n20498), .ZN(n20511) );
  OAI21_X1 U23446 ( .B1(n20565), .B2(n20499), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20500) );
  NAND2_X1 U23447 ( .A1(n20500), .A2(n20741), .ZN(n20509) );
  AND2_X1 U23448 ( .A1(n20540), .A2(n9946), .ZN(n20506) );
  OR2_X1 U23449 ( .A1(n20501), .A2(n20882), .ZN(n20675) );
  NAND2_X1 U23450 ( .A1(n20675), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20685) );
  OAI21_X1 U23451 ( .B1(n20589), .B2(n20502), .A(n20685), .ZN(n20503) );
  INV_X1 U23452 ( .A(n20503), .ZN(n20505) );
  INV_X1 U23453 ( .A(n20506), .ZN(n20508) );
  AOI22_X1 U23454 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20533), .B1(
        n20596), .B2(n20532), .ZN(n20510) );
  OAI211_X1 U23455 ( .C1(n20692), .C2(n20536), .A(n20511), .B(n20510), .ZN(
        P1_U3113) );
  OAI22_X1 U23456 ( .A1(n20536), .A2(n20697), .B1(n20754), .B2(n20530), .ZN(
        n20512) );
  INV_X1 U23457 ( .A(n20512), .ZN(n20514) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20533), .B1(
        n20600), .B2(n20532), .ZN(n20513) );
  OAI211_X1 U23459 ( .C1(n20760), .C2(n20581), .A(n20514), .B(n20513), .ZN(
        P1_U3114) );
  OAI22_X1 U23460 ( .A1(n20581), .A2(n20767), .B1(n20761), .B2(n20530), .ZN(
        n20515) );
  INV_X1 U23461 ( .A(n20515), .ZN(n20517) );
  AOI22_X1 U23462 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20533), .B1(
        n20604), .B2(n20532), .ZN(n20516) );
  OAI211_X1 U23463 ( .C1(n20702), .C2(n20536), .A(n20517), .B(n20516), .ZN(
        P1_U3115) );
  OAI22_X1 U23464 ( .A1(n20581), .A2(n20774), .B1(n20768), .B2(n20530), .ZN(
        n20518) );
  INV_X1 U23465 ( .A(n20518), .ZN(n20520) );
  AOI22_X1 U23466 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20533), .B1(
        n20608), .B2(n20532), .ZN(n20519) );
  OAI211_X1 U23467 ( .C1(n20707), .C2(n20536), .A(n20520), .B(n20519), .ZN(
        P1_U3116) );
  OAI22_X1 U23468 ( .A1(n20536), .A2(n20712), .B1(n20775), .B2(n20530), .ZN(
        n20521) );
  INV_X1 U23469 ( .A(n20521), .ZN(n20523) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20533), .B1(
        n20612), .B2(n20532), .ZN(n20522) );
  OAI211_X1 U23471 ( .C1(n20781), .C2(n20581), .A(n20523), .B(n20522), .ZN(
        P1_U3117) );
  OAI22_X1 U23472 ( .A1(n20536), .A2(n20717), .B1(n20782), .B2(n20530), .ZN(
        n20524) );
  INV_X1 U23473 ( .A(n20524), .ZN(n20526) );
  AOI22_X1 U23474 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20533), .B1(
        n20616), .B2(n20532), .ZN(n20525) );
  OAI211_X1 U23475 ( .C1(n20788), .C2(n20581), .A(n20526), .B(n20525), .ZN(
        P1_U3118) );
  OAI22_X1 U23476 ( .A1(n20536), .A2(n20722), .B1(n20789), .B2(n20530), .ZN(
        n20527) );
  INV_X1 U23477 ( .A(n20527), .ZN(n20529) );
  AOI22_X1 U23478 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20533), .B1(
        n20620), .B2(n20532), .ZN(n20528) );
  OAI211_X1 U23479 ( .C1(n20795), .C2(n20581), .A(n20529), .B(n20528), .ZN(
        P1_U3119) );
  OAI22_X1 U23480 ( .A1(n20581), .A2(n20912), .B1(n20908), .B2(n20530), .ZN(
        n20531) );
  INV_X1 U23481 ( .A(n20531), .ZN(n20535) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20533), .B1(
        n20626), .B2(n20532), .ZN(n20534) );
  OAI211_X1 U23483 ( .C1(n20910), .C2(n20536), .A(n20535), .B(n20534), .ZN(
        P1_U3120) );
  NOR2_X1 U23484 ( .A1(n20538), .A2(n20537), .ZN(n20543) );
  AOI21_X1 U23485 ( .B1(n20540), .B2(n20539), .A(n20543), .ZN(n20546) );
  OR2_X1 U23486 ( .A1(n20546), .A2(n20744), .ZN(n20542) );
  NAND2_X1 U23487 ( .A1(n20550), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20541) );
  INV_X1 U23488 ( .A(n20543), .ZN(n20575) );
  OAI22_X1 U23489 ( .A1(n20739), .A2(n20574), .B1(n20738), .B2(n20575), .ZN(
        n20544) );
  INV_X1 U23490 ( .A(n20544), .ZN(n20554) );
  INV_X1 U23491 ( .A(n20552), .ZN(n20545) );
  NOR2_X1 U23492 ( .A1(n20545), .A2(n20744), .ZN(n20547) );
  OAI21_X1 U23493 ( .B1(n20548), .B2(n20547), .A(n20546), .ZN(n20549) );
  OAI211_X1 U23494 ( .C1(n20741), .C2(n20550), .A(n20748), .B(n20549), .ZN(
        n20578) );
  INV_X1 U23495 ( .A(n20630), .ZN(n20577) );
  AOI22_X1 U23496 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20689), .ZN(n20553) );
  OAI211_X1 U23497 ( .C1(n20692), .C2(n20581), .A(n20554), .B(n20553), .ZN(
        P1_U3121) );
  OAI22_X1 U23498 ( .A1(n20755), .A2(n20574), .B1(n20754), .B2(n20575), .ZN(
        n20555) );
  INV_X1 U23499 ( .A(n20555), .ZN(n20557) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20578), .B1(
        n20565), .B2(n20757), .ZN(n20556) );
  OAI211_X1 U23501 ( .C1(n20760), .C2(n20630), .A(n20557), .B(n20556), .ZN(
        P1_U3122) );
  OAI22_X1 U23502 ( .A1(n20762), .A2(n20574), .B1(n20761), .B2(n20575), .ZN(
        n20558) );
  INV_X1 U23503 ( .A(n20558), .ZN(n20560) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20578), .B1(
        n20565), .B2(n20764), .ZN(n20559) );
  OAI211_X1 U23505 ( .C1(n20767), .C2(n20630), .A(n20560), .B(n20559), .ZN(
        P1_U3123) );
  OAI22_X1 U23506 ( .A1(n20769), .A2(n20574), .B1(n20768), .B2(n20575), .ZN(
        n20561) );
  INV_X1 U23507 ( .A(n20561), .ZN(n20563) );
  AOI22_X1 U23508 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20704), .ZN(n20562) );
  OAI211_X1 U23509 ( .C1(n20707), .C2(n20581), .A(n20563), .B(n20562), .ZN(
        P1_U3124) );
  OAI22_X1 U23510 ( .A1(n20776), .A2(n20574), .B1(n20775), .B2(n20575), .ZN(
        n20564) );
  INV_X1 U23511 ( .A(n20564), .ZN(n20567) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20578), .B1(
        n20565), .B2(n20778), .ZN(n20566) );
  OAI211_X1 U23513 ( .C1(n20781), .C2(n20630), .A(n20567), .B(n20566), .ZN(
        P1_U3125) );
  OAI22_X1 U23514 ( .A1(n20783), .A2(n20574), .B1(n20782), .B2(n20575), .ZN(
        n20568) );
  INV_X1 U23515 ( .A(n20568), .ZN(n20570) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20714), .ZN(n20569) );
  OAI211_X1 U23517 ( .C1(n20717), .C2(n20581), .A(n20570), .B(n20569), .ZN(
        P1_U3126) );
  OAI22_X1 U23518 ( .A1(n20790), .A2(n20574), .B1(n20789), .B2(n20575), .ZN(
        n20571) );
  INV_X1 U23519 ( .A(n20571), .ZN(n20573) );
  AOI22_X1 U23520 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n9633), .ZN(n20572) );
  OAI211_X1 U23521 ( .C1(n20722), .C2(n20581), .A(n20573), .B(n20572), .ZN(
        P1_U3127) );
  OAI22_X1 U23522 ( .A1(n20908), .A2(n20575), .B1(n20574), .B2(n20913), .ZN(
        n20576) );
  INV_X1 U23523 ( .A(n20576), .ZN(n20580) );
  AOI22_X1 U23524 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20578), .B1(
        n20577), .B2(n20726), .ZN(n20579) );
  OAI211_X1 U23525 ( .C1(n20910), .C2(n20581), .A(n20580), .B(n20579), .ZN(
        P1_U3128) );
  NAND2_X1 U23526 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20745) );
  OR2_X1 U23527 ( .A1(n20583), .A2(n20745), .ZN(n20623) );
  OAI22_X1 U23528 ( .A1(n20753), .A2(n20645), .B1(n20738), .B2(n20623), .ZN(
        n20584) );
  INV_X1 U23529 ( .A(n20584), .ZN(n20598) );
  INV_X1 U23530 ( .A(n20623), .ZN(n20590) );
  NAND3_X1 U23531 ( .A1(n20630), .A2(n20741), .A3(n20645), .ZN(n20586) );
  NAND2_X1 U23532 ( .A1(n20586), .A2(n20585), .ZN(n20591) );
  OR2_X1 U23533 ( .A1(n13122), .A2(n20587), .ZN(n20732) );
  OR2_X1 U23534 ( .A1(n20732), .A2(n9946), .ZN(n20594) );
  AOI22_X1 U23535 ( .A1(n20591), .A2(n20594), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20593), .ZN(n20588) );
  OAI211_X1 U23536 ( .C1(n20590), .C2(n20589), .A(n20686), .B(n20588), .ZN(
        n20627) );
  INV_X1 U23537 ( .A(n20591), .ZN(n20595) );
  AOI22_X1 U23538 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20627), .B1(
        n20596), .B2(n20625), .ZN(n20597) );
  OAI211_X1 U23539 ( .C1(n20692), .C2(n20630), .A(n20598), .B(n20597), .ZN(
        P1_U3129) );
  OAI22_X1 U23540 ( .A1(n20760), .A2(n20645), .B1(n20754), .B2(n20623), .ZN(
        n20599) );
  INV_X1 U23541 ( .A(n20599), .ZN(n20602) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20627), .B1(
        n20600), .B2(n20625), .ZN(n20601) );
  OAI211_X1 U23543 ( .C1(n20697), .C2(n20630), .A(n20602), .B(n20601), .ZN(
        P1_U3130) );
  OAI22_X1 U23544 ( .A1(n20767), .A2(n20645), .B1(n20761), .B2(n20623), .ZN(
        n20603) );
  INV_X1 U23545 ( .A(n20603), .ZN(n20606) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20627), .B1(
        n20604), .B2(n20625), .ZN(n20605) );
  OAI211_X1 U23547 ( .C1(n20702), .C2(n20630), .A(n20606), .B(n20605), .ZN(
        P1_U3131) );
  OAI22_X1 U23548 ( .A1(n20774), .A2(n20645), .B1(n20768), .B2(n20623), .ZN(
        n20607) );
  INV_X1 U23549 ( .A(n20607), .ZN(n20610) );
  AOI22_X1 U23550 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20627), .B1(
        n20608), .B2(n20625), .ZN(n20609) );
  OAI211_X1 U23551 ( .C1(n20707), .C2(n20630), .A(n20610), .B(n20609), .ZN(
        P1_U3132) );
  OAI22_X1 U23552 ( .A1(n20781), .A2(n20645), .B1(n20775), .B2(n20623), .ZN(
        n20611) );
  INV_X1 U23553 ( .A(n20611), .ZN(n20614) );
  AOI22_X1 U23554 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20627), .B1(
        n20612), .B2(n20625), .ZN(n20613) );
  OAI211_X1 U23555 ( .C1(n20712), .C2(n20630), .A(n20614), .B(n20613), .ZN(
        P1_U3133) );
  OAI22_X1 U23556 ( .A1(n20788), .A2(n20645), .B1(n20782), .B2(n20623), .ZN(
        n20615) );
  INV_X1 U23557 ( .A(n20615), .ZN(n20618) );
  AOI22_X1 U23558 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20627), .B1(
        n20616), .B2(n20625), .ZN(n20617) );
  OAI211_X1 U23559 ( .C1(n20717), .C2(n20630), .A(n20618), .B(n20617), .ZN(
        P1_U3134) );
  OAI22_X1 U23560 ( .A1(n20795), .A2(n20645), .B1(n20789), .B2(n20623), .ZN(
        n20619) );
  INV_X1 U23561 ( .A(n20619), .ZN(n20622) );
  AOI22_X1 U23562 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20627), .B1(
        n20620), .B2(n20625), .ZN(n20621) );
  OAI211_X1 U23563 ( .C1(n20722), .C2(n20630), .A(n20622), .B(n20621), .ZN(
        P1_U3135) );
  OAI22_X1 U23564 ( .A1(n20912), .A2(n20645), .B1(n20908), .B2(n20623), .ZN(
        n20624) );
  INV_X1 U23565 ( .A(n20624), .ZN(n20629) );
  AOI22_X1 U23566 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20627), .B1(
        n20626), .B2(n20625), .ZN(n20628) );
  OAI211_X1 U23567 ( .C1(n20910), .C2(n20630), .A(n20629), .B(n20628), .ZN(
        P1_U3136) );
  INV_X1 U23568 ( .A(n20743), .ZN(n20633) );
  INV_X1 U23569 ( .A(n20631), .ZN(n20632) );
  OR2_X1 U23570 ( .A1(n20732), .A2(n20634), .ZN(n20636) );
  OR3_X1 U23571 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20635), .A3(
        n20745), .ZN(n20667) );
  NAND2_X1 U23572 ( .A1(n20636), .A2(n20667), .ZN(n20640) );
  NAND2_X1 U23573 ( .A1(n20640), .A2(n20741), .ZN(n20638) );
  NOR2_X1 U23574 ( .A1(n20745), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n20644) );
  NAND2_X1 U23575 ( .A1(n20644), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20637) );
  AND2_X1 U23576 ( .A1(n20638), .A2(n20637), .ZN(n20666) );
  OAI22_X1 U23577 ( .A1(n20739), .A2(n20666), .B1(n20738), .B2(n20667), .ZN(
        n20639) );
  INV_X1 U23578 ( .A(n20639), .ZN(n20647) );
  INV_X1 U23579 ( .A(n20640), .ZN(n20641) );
  OAI21_X1 U23580 ( .B1(n20743), .B2(n20642), .A(n20641), .ZN(n20643) );
  OAI211_X1 U23581 ( .C1(n20741), .C2(n20644), .A(n20748), .B(n20643), .ZN(
        n20670) );
  AOI22_X1 U23582 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20750), .ZN(n20646) );
  OAI211_X1 U23583 ( .C1(n20753), .C2(n20730), .A(n20647), .B(n20646), .ZN(
        P1_U3137) );
  OAI22_X1 U23584 ( .A1(n20755), .A2(n20666), .B1(n20754), .B2(n20667), .ZN(
        n20648) );
  INV_X1 U23585 ( .A(n20648), .ZN(n20650) );
  AOI22_X1 U23586 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20757), .ZN(n20649) );
  OAI211_X1 U23587 ( .C1(n20760), .C2(n20730), .A(n20650), .B(n20649), .ZN(
        P1_U3138) );
  OAI22_X1 U23588 ( .A1(n20762), .A2(n20666), .B1(n20761), .B2(n20667), .ZN(
        n20651) );
  INV_X1 U23589 ( .A(n20651), .ZN(n20653) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20764), .ZN(n20652) );
  OAI211_X1 U23591 ( .C1(n20767), .C2(n20730), .A(n20653), .B(n20652), .ZN(
        P1_U3139) );
  OAI22_X1 U23592 ( .A1(n20769), .A2(n20666), .B1(n20768), .B2(n20667), .ZN(
        n20654) );
  INV_X1 U23593 ( .A(n20654), .ZN(n20656) );
  AOI22_X1 U23594 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20771), .ZN(n20655) );
  OAI211_X1 U23595 ( .C1(n20774), .C2(n20730), .A(n20656), .B(n20655), .ZN(
        P1_U3140) );
  OAI22_X1 U23596 ( .A1(n20776), .A2(n20666), .B1(n20775), .B2(n20667), .ZN(
        n20657) );
  INV_X1 U23597 ( .A(n20657), .ZN(n20659) );
  AOI22_X1 U23598 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20778), .ZN(n20658) );
  OAI211_X1 U23599 ( .C1(n20781), .C2(n20730), .A(n20659), .B(n20658), .ZN(
        P1_U3141) );
  OAI22_X1 U23600 ( .A1(n20783), .A2(n20666), .B1(n20782), .B2(n20667), .ZN(
        n20660) );
  INV_X1 U23601 ( .A(n20660), .ZN(n20662) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20785), .ZN(n20661) );
  OAI211_X1 U23603 ( .C1(n20788), .C2(n20730), .A(n20662), .B(n20661), .ZN(
        P1_U3142) );
  OAI22_X1 U23604 ( .A1(n20790), .A2(n20666), .B1(n20789), .B2(n20667), .ZN(
        n20663) );
  INV_X1 U23605 ( .A(n20663), .ZN(n20665) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20792), .ZN(n20664) );
  OAI211_X1 U23607 ( .C1(n20795), .C2(n20730), .A(n20665), .B(n20664), .ZN(
        P1_U3143) );
  OAI22_X1 U23608 ( .A1(n20908), .A2(n20667), .B1(n20666), .B2(n20913), .ZN(
        n20668) );
  INV_X1 U23609 ( .A(n20668), .ZN(n20672) );
  AOI22_X1 U23610 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20670), .B1(
        n20669), .B2(n20799), .ZN(n20671) );
  OAI211_X1 U23611 ( .C1(n20912), .C2(n20730), .A(n20672), .B(n20671), .ZN(
        P1_U3144) );
  OR2_X1 U23612 ( .A1(n20732), .A2(n20673), .ZN(n20683) );
  INV_X1 U23613 ( .A(n20683), .ZN(n20674) );
  NAND2_X1 U23614 ( .A1(n20674), .A2(n20741), .ZN(n20679) );
  INV_X1 U23615 ( .A(n20675), .ZN(n20676) );
  NAND2_X1 U23616 ( .A1(n20677), .A2(n20676), .ZN(n20678) );
  AND2_X1 U23617 ( .A1(n20679), .A2(n20678), .ZN(n20723) );
  NOR3_X1 U23618 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20746), .A3(
        n20745), .ZN(n20688) );
  INV_X1 U23619 ( .A(n20688), .ZN(n20724) );
  OAI22_X1 U23620 ( .A1(n20739), .A2(n20723), .B1(n20738), .B2(n20724), .ZN(
        n20680) );
  INV_X1 U23621 ( .A(n20680), .ZN(n20691) );
  INV_X1 U23622 ( .A(n20730), .ZN(n20682) );
  NOR2_X2 U23623 ( .A1(n20743), .A2(n20681), .ZN(n20800) );
  OAI21_X1 U23624 ( .B1(n20682), .B2(n20800), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20684) );
  AOI21_X1 U23625 ( .B1(n20684), .B2(n20683), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n20687) );
  AOI22_X1 U23626 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20727), .B1(
        n20800), .B2(n20689), .ZN(n20690) );
  OAI211_X1 U23627 ( .C1(n20692), .C2(n20730), .A(n20691), .B(n20690), .ZN(
        P1_U3145) );
  OAI22_X1 U23628 ( .A1(n20755), .A2(n20723), .B1(n20754), .B2(n20724), .ZN(
        n20693) );
  INV_X1 U23629 ( .A(n20693), .ZN(n20696) );
  AOI22_X1 U23630 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20727), .B1(
        n20800), .B2(n20694), .ZN(n20695) );
  OAI211_X1 U23631 ( .C1(n20697), .C2(n20730), .A(n20696), .B(n20695), .ZN(
        P1_U3146) );
  OAI22_X1 U23632 ( .A1(n20762), .A2(n20723), .B1(n20761), .B2(n20724), .ZN(
        n20698) );
  INV_X1 U23633 ( .A(n20698), .ZN(n20701) );
  AOI22_X1 U23634 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20727), .B1(
        n20800), .B2(n20699), .ZN(n20700) );
  OAI211_X1 U23635 ( .C1(n20702), .C2(n20730), .A(n20701), .B(n20700), .ZN(
        P1_U3147) );
  OAI22_X1 U23636 ( .A1(n20769), .A2(n20723), .B1(n20768), .B2(n20724), .ZN(
        n20703) );
  INV_X1 U23637 ( .A(n20703), .ZN(n20706) );
  AOI22_X1 U23638 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20727), .B1(
        n20800), .B2(n20704), .ZN(n20705) );
  OAI211_X1 U23639 ( .C1(n20707), .C2(n20730), .A(n20706), .B(n20705), .ZN(
        P1_U3148) );
  OAI22_X1 U23640 ( .A1(n20776), .A2(n20723), .B1(n20775), .B2(n20724), .ZN(
        n20708) );
  INV_X1 U23641 ( .A(n20708), .ZN(n20711) );
  AOI22_X1 U23642 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20727), .B1(
        n20800), .B2(n20709), .ZN(n20710) );
  OAI211_X1 U23643 ( .C1(n20712), .C2(n20730), .A(n20711), .B(n20710), .ZN(
        P1_U3149) );
  OAI22_X1 U23644 ( .A1(n20783), .A2(n20723), .B1(n20782), .B2(n20724), .ZN(
        n20713) );
  INV_X1 U23645 ( .A(n20713), .ZN(n20716) );
  AOI22_X1 U23646 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20727), .B1(
        n20800), .B2(n20714), .ZN(n20715) );
  OAI211_X1 U23647 ( .C1(n20717), .C2(n20730), .A(n20716), .B(n20715), .ZN(
        P1_U3150) );
  OAI22_X1 U23648 ( .A1(n20790), .A2(n20723), .B1(n20789), .B2(n20724), .ZN(
        n20718) );
  INV_X1 U23649 ( .A(n20718), .ZN(n20721) );
  AOI22_X1 U23650 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20727), .B1(
        n20800), .B2(n9633), .ZN(n20720) );
  OAI211_X1 U23651 ( .C1(n20722), .C2(n20730), .A(n20721), .B(n20720), .ZN(
        P1_U3151) );
  OAI22_X1 U23652 ( .A1(n20908), .A2(n20724), .B1(n20723), .B2(n20913), .ZN(
        n20725) );
  INV_X1 U23653 ( .A(n20725), .ZN(n20729) );
  AOI22_X1 U23654 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20727), .B1(
        n20800), .B2(n20726), .ZN(n20728) );
  OAI211_X1 U23655 ( .C1(n20910), .C2(n20730), .A(n20729), .B(n20728), .ZN(
        P1_U3152) );
  OR2_X1 U23656 ( .A1(n20732), .A2(n20731), .ZN(n20735) );
  INV_X1 U23657 ( .A(n20745), .ZN(n20733) );
  NAND2_X1 U23658 ( .A1(n20734), .A2(n20733), .ZN(n20797) );
  NAND2_X1 U23659 ( .A1(n20735), .A2(n20797), .ZN(n20749) );
  NAND2_X1 U23660 ( .A1(n20749), .A2(n20741), .ZN(n20737) );
  NAND2_X1 U23661 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n10162), .ZN(n20736) );
  AND2_X1 U23662 ( .A1(n20737), .A2(n20736), .ZN(n20796) );
  OAI22_X1 U23663 ( .A1(n20739), .A2(n20796), .B1(n20738), .B2(n20797), .ZN(
        n20740) );
  INV_X1 U23664 ( .A(n20740), .ZN(n20752) );
  OAI21_X1 U23665 ( .B1(n20743), .B2(n20742), .A(n20741), .ZN(n20879) );
  OAI21_X1 U23666 ( .B1(n20746), .B2(n20745), .A(n20744), .ZN(n20747) );
  OAI211_X1 U23667 ( .C1(n20879), .C2(n20749), .A(n20748), .B(n20747), .ZN(
        n20801) );
  AOI22_X1 U23668 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20801), .B1(
        n20800), .B2(n20750), .ZN(n20751) );
  OAI211_X1 U23669 ( .C1(n20753), .C2(n20909), .A(n20752), .B(n20751), .ZN(
        P1_U3153) );
  OAI22_X1 U23670 ( .A1(n20755), .A2(n20796), .B1(n20754), .B2(n20797), .ZN(
        n20756) );
  INV_X1 U23671 ( .A(n20756), .ZN(n20759) );
  AOI22_X1 U23672 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20801), .B1(
        n20800), .B2(n20757), .ZN(n20758) );
  OAI211_X1 U23673 ( .C1(n20760), .C2(n20909), .A(n20759), .B(n20758), .ZN(
        P1_U3154) );
  OAI22_X1 U23674 ( .A1(n20762), .A2(n20796), .B1(n20761), .B2(n20797), .ZN(
        n20763) );
  INV_X1 U23675 ( .A(n20763), .ZN(n20766) );
  AOI22_X1 U23676 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20801), .B1(
        n20800), .B2(n20764), .ZN(n20765) );
  OAI211_X1 U23677 ( .C1(n20767), .C2(n20909), .A(n20766), .B(n20765), .ZN(
        P1_U3155) );
  OAI22_X1 U23678 ( .A1(n20769), .A2(n20796), .B1(n20768), .B2(n20797), .ZN(
        n20770) );
  INV_X1 U23679 ( .A(n20770), .ZN(n20773) );
  AOI22_X1 U23680 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20801), .B1(
        n20800), .B2(n20771), .ZN(n20772) );
  OAI211_X1 U23681 ( .C1(n20774), .C2(n20909), .A(n20773), .B(n20772), .ZN(
        P1_U3156) );
  OAI22_X1 U23682 ( .A1(n20776), .A2(n20796), .B1(n20775), .B2(n20797), .ZN(
        n20777) );
  INV_X1 U23683 ( .A(n20777), .ZN(n20780) );
  AOI22_X1 U23684 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20801), .B1(
        n20800), .B2(n20778), .ZN(n20779) );
  OAI211_X1 U23685 ( .C1(n20781), .C2(n20909), .A(n20780), .B(n20779), .ZN(
        P1_U3157) );
  OAI22_X1 U23686 ( .A1(n20783), .A2(n20796), .B1(n20782), .B2(n20797), .ZN(
        n20784) );
  INV_X1 U23687 ( .A(n20784), .ZN(n20787) );
  AOI22_X1 U23688 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20801), .B1(
        n20800), .B2(n20785), .ZN(n20786) );
  OAI211_X1 U23689 ( .C1(n20788), .C2(n20909), .A(n20787), .B(n20786), .ZN(
        P1_U3158) );
  OAI22_X1 U23690 ( .A1(n20790), .A2(n20796), .B1(n20789), .B2(n20797), .ZN(
        n20791) );
  INV_X1 U23691 ( .A(n20791), .ZN(n20794) );
  AOI22_X1 U23692 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20801), .B1(
        n20800), .B2(n20792), .ZN(n20793) );
  OAI211_X1 U23693 ( .C1(n20795), .C2(n20909), .A(n20794), .B(n20793), .ZN(
        P1_U3159) );
  OAI22_X1 U23694 ( .A1(n20908), .A2(n20797), .B1(n20796), .B2(n20913), .ZN(
        n20798) );
  INV_X1 U23695 ( .A(n20798), .ZN(n20803) );
  AOI22_X1 U23696 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20801), .B1(
        n20800), .B2(n20799), .ZN(n20802) );
  OAI211_X1 U23697 ( .C1(n20912), .C2(n20909), .A(n20803), .B(n20802), .ZN(
        P1_U3160) );
  NOR2_X1 U23698 ( .A1(n20804), .A2(n21068), .ZN(n20806) );
  OAI21_X1 U23699 ( .B1(n20806), .B2(n20383), .A(n20805), .ZN(P1_U3163) );
  INV_X1 U23700 ( .A(P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n21049) );
  NOR2_X1 U23701 ( .A1(n20807), .A2(n21049), .ZN(P1_U3164) );
  AND2_X1 U23702 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20874), .ZN(
        P1_U3165) );
  AND2_X1 U23703 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20874), .ZN(
        P1_U3166) );
  AND2_X1 U23704 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20874), .ZN(
        P1_U3167) );
  AND2_X1 U23705 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20874), .ZN(
        P1_U3168) );
  AND2_X1 U23706 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20874), .ZN(
        P1_U3169) );
  AND2_X1 U23707 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20874), .ZN(
        P1_U3170) );
  AND2_X1 U23708 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20874), .ZN(
        P1_U3171) );
  AND2_X1 U23709 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20874), .ZN(
        P1_U3172) );
  AND2_X1 U23710 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20874), .ZN(
        P1_U3173) );
  AND2_X1 U23711 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20874), .ZN(
        P1_U3174) );
  AND2_X1 U23712 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20874), .ZN(
        P1_U3175) );
  AND2_X1 U23713 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20874), .ZN(
        P1_U3176) );
  AND2_X1 U23714 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20874), .ZN(
        P1_U3177) );
  AND2_X1 U23715 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20874), .ZN(
        P1_U3178) );
  AND2_X1 U23716 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20874), .ZN(
        P1_U3179) );
  AND2_X1 U23717 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20874), .ZN(
        P1_U3180) );
  AND2_X1 U23718 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20874), .ZN(
        P1_U3181) );
  AND2_X1 U23719 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20874), .ZN(
        P1_U3182) );
  AND2_X1 U23720 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20874), .ZN(
        P1_U3183) );
  AND2_X1 U23721 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20874), .ZN(
        P1_U3184) );
  AND2_X1 U23722 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20874), .ZN(
        P1_U3185) );
  AND2_X1 U23723 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20874), .ZN(P1_U3186) );
  AND2_X1 U23724 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20874), .ZN(P1_U3187) );
  AND2_X1 U23725 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20874), .ZN(P1_U3188) );
  AND2_X1 U23726 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20874), .ZN(P1_U3189) );
  AND2_X1 U23727 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20874), .ZN(P1_U3190) );
  AND2_X1 U23728 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20874), .ZN(P1_U3191) );
  AND2_X1 U23729 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20874), .ZN(P1_U3192) );
  AND2_X1 U23730 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20874), .ZN(P1_U3193) );
  NOR2_X1 U23731 ( .A1(n20808), .A2(n20819), .ZN(n20816) );
  NOR2_X1 U23732 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20810) );
  OAI22_X1 U23733 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20818), .B1(n20810), 
        .B2(n20809), .ZN(n20811) );
  NOR2_X1 U23734 ( .A1(n20815), .A2(n20811), .ZN(n20812) );
  OAI22_X1 U23735 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20816), .B1(n20904), 
        .B2(n20812), .ZN(P1_U3194) );
  AOI21_X1 U23736 ( .B1(n20814), .B2(n20818), .A(n20813), .ZN(n20823) );
  OAI211_X1 U23737 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20815), .A(
        P1_STATE_REG_0__SCAN_IN), .B(HOLD), .ZN(n20822) );
  INV_X1 U23738 ( .A(n20816), .ZN(n20817) );
  OAI211_X1 U23739 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20818), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20817), .ZN(n20821) );
  NAND4_X1 U23740 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(
        P1_STATE_REG_0__SCAN_IN), .A3(n20819), .A4(n20818), .ZN(n20820) );
  OAI211_X1 U23741 ( .C1(n20823), .C2(n20822), .A(n20821), .B(n20820), .ZN(
        P1_U3196) );
  INV_X1 U23742 ( .A(n20864), .ZN(n20861) );
  OAI222_X1 U23743 ( .A1(n20866), .A2(n20827), .B1(n20826), .B2(n20904), .C1(
        n20825), .C2(n20861), .ZN(P1_U3197) );
  AOI222_X1 U23744 ( .A1(n20864), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20859), .ZN(n20828) );
  INV_X1 U23745 ( .A(n20828), .ZN(P1_U3198) );
  AOI222_X1 U23746 ( .A1(n20864), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20859), .ZN(n20829) );
  INV_X1 U23747 ( .A(n20829), .ZN(P1_U3199) );
  AOI222_X1 U23748 ( .A1(n20859), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20864), .ZN(n20830) );
  INV_X1 U23749 ( .A(n20830), .ZN(P1_U3200) );
  AOI222_X1 U23750 ( .A1(n20864), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20859), .ZN(n20831) );
  INV_X1 U23751 ( .A(n20831), .ZN(P1_U3201) );
  AOI222_X1 U23752 ( .A1(n20864), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20859), .ZN(n20832) );
  INV_X1 U23753 ( .A(n20832), .ZN(P1_U3202) );
  AOI222_X1 U23754 ( .A1(n20864), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20859), .ZN(n20833) );
  INV_X1 U23755 ( .A(n20833), .ZN(P1_U3203) );
  INV_X1 U23756 ( .A(P1_ADDRESS_REG_7__SCAN_IN), .ZN(n21091) );
  INV_X1 U23757 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20834) );
  OAI222_X1 U23758 ( .A1(n20866), .A2(n20836), .B1(n21091), .B2(n20904), .C1(
        n20834), .C2(n20861), .ZN(P1_U3204) );
  AOI22_X1 U23759 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n20905), .B1(
        P1_REIP_REG_10__SCAN_IN), .B2(n20859), .ZN(n20835) );
  OAI21_X1 U23760 ( .B1(n20836), .B2(n20861), .A(n20835), .ZN(P1_U3205) );
  AOI22_X1 U23761 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(n20905), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n20859), .ZN(n20837) );
  OAI21_X1 U23762 ( .B1(n14511), .B2(n20861), .A(n20837), .ZN(P1_U3206) );
  AOI22_X1 U23763 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(n20905), .B1(
        P1_REIP_REG_11__SCAN_IN), .B2(n20864), .ZN(n20838) );
  OAI21_X1 U23764 ( .B1(n20839), .B2(n20866), .A(n20838), .ZN(P1_U3207) );
  INV_X1 U23765 ( .A(P1_ADDRESS_REG_11__SCAN_IN), .ZN(n21032) );
  OAI222_X1 U23766 ( .A1(n20861), .A2(n20839), .B1(n21032), .B2(n20904), .C1(
        n14498), .C2(n20866), .ZN(P1_U3208) );
  AOI222_X1 U23767 ( .A1(n20864), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20859), .ZN(n20840) );
  INV_X1 U23768 ( .A(n20840), .ZN(P1_U3209) );
  AOI222_X1 U23769 ( .A1(n20859), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20864), .ZN(n20841) );
  INV_X1 U23770 ( .A(n20841), .ZN(P1_U3210) );
  AOI222_X1 U23771 ( .A1(n20864), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20859), .ZN(n20842) );
  INV_X1 U23772 ( .A(n20842), .ZN(P1_U3211) );
  AOI222_X1 U23773 ( .A1(n20864), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20859), .ZN(n20843) );
  INV_X1 U23774 ( .A(n20843), .ZN(P1_U3212) );
  AOI222_X1 U23775 ( .A1(n20864), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20859), .ZN(n20844) );
  INV_X1 U23776 ( .A(n20844), .ZN(P1_U3213) );
  AOI222_X1 U23777 ( .A1(n20864), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20859), .ZN(n20845) );
  INV_X1 U23778 ( .A(n20845), .ZN(P1_U3214) );
  AOI22_X1 U23779 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20905), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20859), .ZN(n20846) );
  OAI21_X1 U23780 ( .B1(n20847), .B2(n20861), .A(n20846), .ZN(P1_U3215) );
  AOI22_X1 U23781 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20905), .B1(
        P1_REIP_REG_20__SCAN_IN), .B2(n20864), .ZN(n20848) );
  OAI21_X1 U23782 ( .B1(n20849), .B2(n20866), .A(n20848), .ZN(P1_U3216) );
  AOI222_X1 U23783 ( .A1(n20864), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20859), .ZN(n20850) );
  INV_X1 U23784 ( .A(n20850), .ZN(P1_U3217) );
  AOI22_X1 U23785 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20905), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20859), .ZN(n20851) );
  OAI21_X1 U23786 ( .B1(n14463), .B2(n20861), .A(n20851), .ZN(P1_U3218) );
  AOI22_X1 U23787 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20905), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20864), .ZN(n20852) );
  OAI21_X1 U23788 ( .B1(n20853), .B2(n20866), .A(n20852), .ZN(P1_U3219) );
  AOI222_X1 U23789 ( .A1(n20864), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20859), .ZN(n20854) );
  INV_X1 U23790 ( .A(n20854), .ZN(P1_U3220) );
  AOI222_X1 U23791 ( .A1(n20864), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20859), .ZN(n20855) );
  INV_X1 U23792 ( .A(n20855), .ZN(P1_U3221) );
  AOI222_X1 U23793 ( .A1(n20864), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20859), .ZN(n20856) );
  INV_X1 U23794 ( .A(n20856), .ZN(P1_U3222) );
  AOI222_X1 U23795 ( .A1(n20864), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20859), .ZN(n20857) );
  INV_X1 U23796 ( .A(n20857), .ZN(P1_U3223) );
  AOI222_X1 U23797 ( .A1(n20864), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20863), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20859), .ZN(n20858) );
  INV_X1 U23798 ( .A(n20858), .ZN(P1_U3224) );
  AOI22_X1 U23799 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20859), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20863), .ZN(n20860) );
  OAI21_X1 U23800 ( .B1(n20862), .B2(n20861), .A(n20860), .ZN(P1_U3225) );
  INV_X1 U23801 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20867) );
  AOI22_X1 U23802 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(n20864), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20863), .ZN(n20865) );
  OAI21_X1 U23803 ( .B1(n20867), .B2(n20866), .A(n20865), .ZN(P1_U3226) );
  OAI22_X1 U23804 ( .A1(n20905), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20904), .ZN(n20868) );
  INV_X1 U23805 ( .A(n20868), .ZN(P1_U3458) );
  OAI22_X1 U23806 ( .A1(n20905), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20904), .ZN(n20869) );
  INV_X1 U23807 ( .A(n20869), .ZN(P1_U3459) );
  OAI22_X1 U23808 ( .A1(n20905), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20904), .ZN(n20870) );
  INV_X1 U23809 ( .A(n20870), .ZN(P1_U3460) );
  OAI22_X1 U23810 ( .A1(n20905), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20904), .ZN(n20871) );
  INV_X1 U23811 ( .A(n20871), .ZN(P1_U3461) );
  INV_X1 U23812 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n20885) );
  INV_X1 U23813 ( .A(n20872), .ZN(n20873) );
  AOI21_X1 U23814 ( .B1(n20885), .B2(n20874), .A(n20873), .ZN(P1_U3464) );
  AOI21_X1 U23815 ( .B1(n20874), .B2(P1_DATAWIDTH_REG_1__SCAN_IN), .A(n20873), 
        .ZN(n20875) );
  INV_X1 U23816 ( .A(n20875), .ZN(P1_U3465) );
  AOI21_X1 U23817 ( .B1(n13145), .B2(n20877), .A(n20876), .ZN(n20878) );
  OAI21_X1 U23818 ( .B1(n13353), .B2(n20879), .A(n20878), .ZN(n20880) );
  NAND2_X1 U23819 ( .A1(n20883), .A2(n20880), .ZN(n20881) );
  OAI21_X1 U23820 ( .B1(n20883), .B2(n20882), .A(n20881), .ZN(P1_U3475) );
  NOR3_X1 U23821 ( .A1(n20885), .A2(P1_REIP_REG_0__SCAN_IN), .A3(
        P1_REIP_REG_1__SCAN_IN), .ZN(n20884) );
  AOI221_X1 U23822 ( .B1(n20886), .B2(n20885), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n20884), .ZN(n20888) );
  INV_X1 U23823 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20887) );
  INV_X1 U23824 ( .A(n20892), .ZN(n20889) );
  AOI22_X1 U23825 ( .A1(n20892), .A2(n20888), .B1(n20887), .B2(n20889), .ZN(
        P1_U3481) );
  NOR2_X1 U23826 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .ZN(n20891) );
  INV_X1 U23827 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20890) );
  AOI22_X1 U23828 ( .A1(n20892), .A2(n20891), .B1(n20890), .B2(n20889), .ZN(
        P1_U3482) );
  AOI22_X1 U23829 ( .A1(n20904), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20893), 
        .B2(n20905), .ZN(P1_U3483) );
  AOI211_X1 U23830 ( .C1(n20039), .C2(n20896), .A(n20895), .B(n20894), .ZN(
        n20903) );
  OAI211_X1 U23831 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20898), .A(n20897), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20900) );
  AOI21_X1 U23832 ( .B1(n20900), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20899), 
        .ZN(n20902) );
  NAND2_X1 U23833 ( .A1(n20903), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20901) );
  OAI21_X1 U23834 ( .B1(n20903), .B2(n20902), .A(n20901), .ZN(P1_U3485) );
  OAI22_X1 U23835 ( .A1(n20905), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n20904), .ZN(n20906) );
  INV_X1 U23836 ( .A(n20906), .ZN(P1_U3486) );
  OAI22_X1 U23837 ( .A1(n20910), .A2(n20909), .B1(n20908), .B2(n20907), .ZN(
        n20916) );
  OAI22_X1 U23838 ( .A1(n20914), .A2(n20913), .B1(n20912), .B2(n20911), .ZN(
        n20915) );
  AOI211_X1 U23839 ( .C1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .C2(n20917), .A(
        n20916), .B(n20915), .ZN(n21112) );
  INV_X1 U23840 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n20919) );
  AOI22_X1 U23841 ( .A1(n21042), .A2(keyinput87), .B1(n20919), .B2(keyinput118), .ZN(n20918) );
  OAI221_X1 U23842 ( .B1(n21042), .B2(keyinput87), .C1(n20919), .C2(
        keyinput118), .A(n20918), .ZN(n20929) );
  AOI22_X1 U23843 ( .A1(n12874), .A2(keyinput91), .B1(keyinput89), .B2(n20921), 
        .ZN(n20920) );
  OAI221_X1 U23844 ( .B1(n12874), .B2(keyinput91), .C1(n20921), .C2(keyinput89), .A(n20920), .ZN(n20928) );
  AOI22_X1 U23845 ( .A1(n20924), .A2(keyinput107), .B1(n20923), .B2(keyinput85), .ZN(n20922) );
  OAI221_X1 U23846 ( .B1(n20924), .B2(keyinput107), .C1(n20923), .C2(
        keyinput85), .A(n20922), .ZN(n20927) );
  INV_X1 U23847 ( .A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n21046) );
  AOI22_X1 U23848 ( .A1(n21079), .A2(keyinput108), .B1(keyinput71), .B2(n21046), .ZN(n20925) );
  OAI221_X1 U23849 ( .B1(n21079), .B2(keyinput108), .C1(n21046), .C2(
        keyinput71), .A(n20925), .ZN(n20926) );
  NOR4_X1 U23850 ( .A1(n20929), .A2(n20928), .A3(n20927), .A4(n20926), .ZN(
        n20967) );
  AOI22_X1 U23851 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(keyinput78), .B1(n20931), .B2(keyinput115), .ZN(n20930) );
  OAI221_X1 U23852 ( .B1(P1_LWORD_REG_14__SCAN_IN), .B2(keyinput78), .C1(
        n20931), .C2(keyinput115), .A(n20930), .ZN(n20941) );
  AOI22_X1 U23853 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(keyinput84), .B1(
        P2_ADDRESS_REG_19__SCAN_IN), .B2(keyinput121), .ZN(n20932) );
  OAI221_X1 U23854 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(keyinput84), .C1(
        P2_ADDRESS_REG_19__SCAN_IN), .C2(keyinput121), .A(n20932), .ZN(n20940)
         );
  AOI22_X1 U23855 ( .A1(n21064), .A2(keyinput67), .B1(n20934), .B2(keyinput112), .ZN(n20933) );
  OAI221_X1 U23856 ( .B1(n21064), .B2(keyinput67), .C1(n20934), .C2(
        keyinput112), .A(n20933), .ZN(n20939) );
  AOI22_X1 U23857 ( .A1(n20937), .A2(keyinput116), .B1(keyinput72), .B2(n20936), .ZN(n20935) );
  OAI221_X1 U23858 ( .B1(n20937), .B2(keyinput116), .C1(n20936), .C2(
        keyinput72), .A(n20935), .ZN(n20938) );
  NOR4_X1 U23859 ( .A1(n20941), .A2(n20940), .A3(n20939), .A4(n20938), .ZN(
        n20966) );
  INV_X1 U23860 ( .A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n21059) );
  AOI22_X1 U23861 ( .A1(n21059), .A2(keyinput102), .B1(n21082), .B2(keyinput68), .ZN(n20942) );
  OAI221_X1 U23862 ( .B1(n21059), .B2(keyinput102), .C1(n21082), .C2(
        keyinput68), .A(n20942), .ZN(n20951) );
  AOI22_X1 U23863 ( .A1(n21074), .A2(keyinput109), .B1(keyinput99), .B2(n21049), .ZN(n20943) );
  OAI221_X1 U23864 ( .B1(n21074), .B2(keyinput109), .C1(n21049), .C2(
        keyinput99), .A(n20943), .ZN(n20950) );
  AOI22_X1 U23865 ( .A1(n21094), .A2(keyinput93), .B1(n20945), .B2(keyinput110), .ZN(n20944) );
  OAI221_X1 U23866 ( .B1(n21094), .B2(keyinput93), .C1(n20945), .C2(
        keyinput110), .A(n20944), .ZN(n20949) );
  INV_X1 U23867 ( .A(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n20947) );
  INV_X1 U23868 ( .A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n21048) );
  AOI22_X1 U23869 ( .A1(n20947), .A2(keyinput79), .B1(keyinput96), .B2(n21048), 
        .ZN(n20946) );
  OAI221_X1 U23870 ( .B1(n20947), .B2(keyinput79), .C1(n21048), .C2(keyinput96), .A(n20946), .ZN(n20948) );
  NOR4_X1 U23871 ( .A1(n20951), .A2(n20950), .A3(n20949), .A4(n20948), .ZN(
        n20965) );
  AOI22_X1 U23872 ( .A1(n21067), .A2(keyinput64), .B1(n20953), .B2(keyinput95), 
        .ZN(n20952) );
  OAI221_X1 U23873 ( .B1(n21067), .B2(keyinput64), .C1(n20953), .C2(keyinput95), .A(n20952), .ZN(n20963) );
  INV_X1 U23874 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n20955) );
  AOI22_X1 U23875 ( .A1(n20956), .A2(keyinput103), .B1(n20955), .B2(keyinput73), .ZN(n20954) );
  OAI221_X1 U23876 ( .B1(n20956), .B2(keyinput103), .C1(n20955), .C2(
        keyinput73), .A(n20954), .ZN(n20962) );
  AOI22_X1 U23877 ( .A1(n21058), .A2(keyinput80), .B1(n20958), .B2(keyinput98), 
        .ZN(n20957) );
  OAI221_X1 U23878 ( .B1(n21058), .B2(keyinput80), .C1(n20958), .C2(keyinput98), .A(n20957), .ZN(n20961) );
  AOI22_X1 U23879 ( .A1(n10820), .A2(keyinput77), .B1(keyinput94), .B2(n21065), 
        .ZN(n20959) );
  OAI221_X1 U23880 ( .B1(n10820), .B2(keyinput77), .C1(n21065), .C2(keyinput94), .A(n20959), .ZN(n20960) );
  NOR4_X1 U23881 ( .A1(n20963), .A2(n20962), .A3(n20961), .A4(n20960), .ZN(
        n20964) );
  AND4_X1 U23882 ( .A1(n20967), .A2(n20966), .A3(n20965), .A4(n20964), .ZN(
        n21110) );
  OAI22_X1 U23883 ( .A1(P2_EAX_REG_26__SCAN_IN), .A2(keyinput126), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(keyinput74), .ZN(n20968) );
  AOI221_X1 U23884 ( .B1(P2_EAX_REG_26__SCAN_IN), .B2(keyinput126), .C1(
        keyinput74), .C2(P2_M_IO_N_REG_SCAN_IN), .A(n20968), .ZN(n20975) );
  OAI22_X1 U23885 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(keyinput114), 
        .B1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput83), .ZN(n20969) );
  AOI221_X1 U23886 ( .B1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B2(keyinput114), 
        .C1(keyinput83), .C2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A(n20969), 
        .ZN(n20974) );
  OAI22_X1 U23887 ( .A1(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(keyinput86), 
        .B1(keyinput82), .B2(P3_EAX_REG_18__SCAN_IN), .ZN(n20970) );
  AOI221_X1 U23888 ( .B1(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput86), 
        .C1(P3_EAX_REG_18__SCAN_IN), .C2(keyinput82), .A(n20970), .ZN(n20973)
         );
  OAI22_X1 U23889 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(keyinput122), 
        .B1(keyinput117), .B2(P3_REIP_REG_20__SCAN_IN), .ZN(n20971) );
  AOI221_X1 U23890 ( .B1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B2(keyinput122), 
        .C1(P3_REIP_REG_20__SCAN_IN), .C2(keyinput117), .A(n20971), .ZN(n20972) );
  NAND4_X1 U23891 ( .A1(n20975), .A2(n20974), .A3(n20973), .A4(n20972), .ZN(
        n21003) );
  OAI22_X1 U23892 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput65), .B1(
        P2_DATAWIDTH_REG_16__SCAN_IN), .B2(keyinput105), .ZN(n20976) );
  AOI221_X1 U23893 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput65), .C1(
        keyinput105), .C2(P2_DATAWIDTH_REG_16__SCAN_IN), .A(n20976), .ZN(
        n20983) );
  OAI22_X1 U23894 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(keyinput100), 
        .B1(P3_EBX_REG_14__SCAN_IN), .B2(keyinput101), .ZN(n20977) );
  AOI221_X1 U23895 ( .B1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B2(keyinput100), 
        .C1(keyinput101), .C2(P3_EBX_REG_14__SCAN_IN), .A(n20977), .ZN(n20982)
         );
  OAI22_X1 U23896 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(keyinput127), 
        .B1(keyinput75), .B2(P2_EBX_REG_26__SCAN_IN), .ZN(n20978) );
  AOI221_X1 U23897 ( .B1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B2(keyinput127), 
        .C1(P2_EBX_REG_26__SCAN_IN), .C2(keyinput75), .A(n20978), .ZN(n20981)
         );
  OAI22_X1 U23898 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(keyinput106), 
        .B1(keyinput111), .B2(P3_EAX_REG_31__SCAN_IN), .ZN(n20979) );
  AOI221_X1 U23899 ( .B1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B2(keyinput106), 
        .C1(P3_EAX_REG_31__SCAN_IN), .C2(keyinput111), .A(n20979), .ZN(n20980)
         );
  NAND4_X1 U23900 ( .A1(n20983), .A2(n20982), .A3(n20981), .A4(n20980), .ZN(
        n21002) );
  OAI22_X1 U23901 ( .A1(P2_EAX_REG_13__SCAN_IN), .A2(keyinput124), .B1(
        keyinput92), .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n20984) );
  AOI221_X1 U23902 ( .B1(P2_EAX_REG_13__SCAN_IN), .B2(keyinput124), .C1(
        P1_DATAO_REG_16__SCAN_IN), .C2(keyinput92), .A(n20984), .ZN(n20991) );
  OAI22_X1 U23903 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(keyinput123), .B1(
        P3_INSTQUEUE_REG_10__2__SCAN_IN), .B2(keyinput120), .ZN(n20985) );
  AOI221_X1 U23904 ( .B1(P1_ADDRESS_REG_7__SCAN_IN), .B2(keyinput123), .C1(
        keyinput120), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(n20985), .ZN(
        n20990) );
  OAI22_X1 U23905 ( .A1(P2_EBX_REG_8__SCAN_IN), .A2(keyinput119), .B1(
        P1_EAX_REG_2__SCAN_IN), .B2(keyinput81), .ZN(n20986) );
  AOI221_X1 U23906 ( .B1(P2_EBX_REG_8__SCAN_IN), .B2(keyinput119), .C1(
        keyinput81), .C2(P1_EAX_REG_2__SCAN_IN), .A(n20986), .ZN(n20989) );
  OAI22_X1 U23907 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(keyinput66), 
        .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput76), .ZN(n20987)
         );
  AOI221_X1 U23908 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(keyinput66), 
        .C1(keyinput76), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(n20987), 
        .ZN(n20988) );
  NAND4_X1 U23909 ( .A1(n20991), .A2(n20990), .A3(n20989), .A4(n20988), .ZN(
        n21001) );
  OAI22_X1 U23910 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(keyinput104), 
        .B1(P1_ADDRESS_REG_11__SCAN_IN), .B2(keyinput97), .ZN(n20992) );
  AOI221_X1 U23911 ( .B1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B2(keyinput104), 
        .C1(keyinput97), .C2(P1_ADDRESS_REG_11__SCAN_IN), .A(n20992), .ZN(
        n20999) );
  OAI22_X1 U23912 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(keyinput69), .B1(
        P1_DATAO_REG_8__SCAN_IN), .B2(keyinput90), .ZN(n20993) );
  AOI221_X1 U23913 ( .B1(P2_DATAO_REG_1__SCAN_IN), .B2(keyinput69), .C1(
        keyinput90), .C2(P1_DATAO_REG_8__SCAN_IN), .A(n20993), .ZN(n20998) );
  OAI22_X1 U23914 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(keyinput88), .B1(
        keyinput70), .B2(P3_REIP_REG_17__SCAN_IN), .ZN(n20994) );
  AOI221_X1 U23915 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(keyinput88), .C1(
        P3_REIP_REG_17__SCAN_IN), .C2(keyinput70), .A(n20994), .ZN(n20997) );
  OAI22_X1 U23916 ( .A1(P2_UWORD_REG_0__SCAN_IN), .A2(keyinput113), .B1(
        P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput125), .ZN(n20995) );
  AOI221_X1 U23917 ( .B1(P2_UWORD_REG_0__SCAN_IN), .B2(keyinput113), .C1(
        keyinput125), .C2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n20995), .ZN(n20996)
         );
  NAND4_X1 U23918 ( .A1(n20999), .A2(n20998), .A3(n20997), .A4(n20996), .ZN(
        n21000) );
  NOR4_X1 U23919 ( .A1(n21003), .A2(n21002), .A3(n21001), .A4(n21000), .ZN(
        n21109) );
  AOI22_X1 U23920 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(keyinput18), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(keyinput55), .ZN(n21004) );
  OAI221_X1 U23921 ( .B1(P3_EAX_REG_18__SCAN_IN), .B2(keyinput18), .C1(
        P2_EBX_REG_8__SCAN_IN), .C2(keyinput55), .A(n21004), .ZN(n21011) );
  AOI22_X1 U23922 ( .A1(P2_CODEFETCH_REG_SCAN_IN), .A2(keyinput25), .B1(
        P3_INSTQUEUE_REG_13__4__SCAN_IN), .B2(keyinput36), .ZN(n21005) );
  OAI221_X1 U23923 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(keyinput25), .C1(
        P3_INSTQUEUE_REG_13__4__SCAN_IN), .C2(keyinput36), .A(n21005), .ZN(
        n21010) );
  AOI22_X1 U23924 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(keyinput47), .B1(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(keyinput51), .ZN(n21006) );
  OAI221_X1 U23925 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(keyinput47), .C1(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(keyinput51), .A(n21006), .ZN(
        n21009) );
  AOI22_X1 U23926 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput61), .B1(
        P1_INSTQUEUE_REG_14__7__SCAN_IN), .B2(keyinput50), .ZN(n21007) );
  OAI221_X1 U23927 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput61), .C1(
        P1_INSTQUEUE_REG_14__7__SCAN_IN), .C2(keyinput50), .A(n21007), .ZN(
        n21008) );
  NOR4_X1 U23928 ( .A1(n21011), .A2(n21010), .A3(n21009), .A4(n21008), .ZN(
        n21040) );
  AOI22_X1 U23929 ( .A1(P3_DATAO_REG_23__SCAN_IN), .A2(keyinput8), .B1(
        P3_EAX_REG_8__SCAN_IN), .B2(keyinput20), .ZN(n21012) );
  OAI221_X1 U23930 ( .B1(P3_DATAO_REG_23__SCAN_IN), .B2(keyinput8), .C1(
        P3_EAX_REG_8__SCAN_IN), .C2(keyinput20), .A(n21012), .ZN(n21019) );
  AOI22_X1 U23931 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(keyinput6), .B1(
        P2_INSTQUEUE_REG_15__6__SCAN_IN), .B2(keyinput54), .ZN(n21013) );
  OAI221_X1 U23932 ( .B1(P3_REIP_REG_17__SCAN_IN), .B2(keyinput6), .C1(
        P2_INSTQUEUE_REG_15__6__SCAN_IN), .C2(keyinput54), .A(n21013), .ZN(
        n21018) );
  AOI22_X1 U23933 ( .A1(P2_LWORD_REG_14__SCAN_IN), .A2(keyinput43), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(keyinput5), .ZN(n21014) );
  OAI221_X1 U23934 ( .B1(P2_LWORD_REG_14__SCAN_IN), .B2(keyinput43), .C1(
        P2_DATAO_REG_1__SCAN_IN), .C2(keyinput5), .A(n21014), .ZN(n21017) );
  AOI22_X1 U23935 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(keyinput37), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(keyinput13), .ZN(n21015) );
  OAI221_X1 U23936 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(keyinput37), .C1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(keyinput13), .A(n21015), .ZN(
        n21016) );
  NOR4_X1 U23937 ( .A1(n21019), .A2(n21018), .A3(n21017), .A4(n21016), .ZN(
        n21039) );
  AOI22_X1 U23938 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(keyinput52), .B1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .B2(keyinput31), .ZN(n21020) );
  OAI221_X1 U23939 ( .B1(P3_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput52), .C1(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .C2(keyinput31), .A(n21020), .ZN(
        n21027) );
  AOI22_X1 U23940 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(keyinput27), .B1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(keyinput48), .ZN(n21021) );
  OAI221_X1 U23941 ( .B1(P2_DATAO_REG_16__SCAN_IN), .B2(keyinput27), .C1(
        P1_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(keyinput48), .A(n21021), .ZN(
        n21026) );
  AOI22_X1 U23942 ( .A1(BUF2_REG_10__SCAN_IN), .A2(keyinput34), .B1(
        P1_INSTQUEUE_REG_11__4__SCAN_IN), .B2(keyinput9), .ZN(n21022) );
  OAI221_X1 U23943 ( .B1(BUF2_REG_10__SCAN_IN), .B2(keyinput34), .C1(
        P1_INSTQUEUE_REG_11__4__SCAN_IN), .C2(keyinput9), .A(n21022), .ZN(
        n21025) );
  AOI22_X1 U23944 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(keyinput28), .B1(
        P2_INSTQUEUE_REG_10__7__SCAN_IN), .B2(keyinput40), .ZN(n21023) );
  OAI221_X1 U23945 ( .B1(P1_DATAO_REG_16__SCAN_IN), .B2(keyinput28), .C1(
        P2_INSTQUEUE_REG_10__7__SCAN_IN), .C2(keyinput40), .A(n21023), .ZN(
        n21024) );
  NOR4_X1 U23946 ( .A1(n21027), .A2(n21026), .A3(n21025), .A4(n21024), .ZN(
        n21038) );
  AOI22_X1 U23947 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(keyinput10), .B1(
        P3_INSTQUEUE_REG_10__2__SCAN_IN), .B2(keyinput56), .ZN(n21028) );
  OAI221_X1 U23948 ( .B1(P2_M_IO_N_REG_SCAN_IN), .B2(keyinput10), .C1(
        P3_INSTQUEUE_REG_10__2__SCAN_IN), .C2(keyinput56), .A(n21028), .ZN(
        n21036) );
  AOI22_X1 U23949 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(keyinput15), 
        .B1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(keyinput21), .ZN(n21029)
         );
  OAI221_X1 U23950 ( .B1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B2(keyinput15), 
        .C1(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(keyinput21), .A(n21029), 
        .ZN(n21035) );
  AOI22_X1 U23951 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(keyinput39), .B1(
        P3_REIP_REG_20__SCAN_IN), .B2(keyinput53), .ZN(n21030) );
  OAI221_X1 U23952 ( .B1(P2_DATAO_REG_20__SCAN_IN), .B2(keyinput39), .C1(
        P3_REIP_REG_20__SCAN_IN), .C2(keyinput53), .A(n21030), .ZN(n21034) );
  AOI22_X1 U23953 ( .A1(BUF1_REG_26__SCAN_IN), .A2(keyinput46), .B1(n21032), 
        .B2(keyinput33), .ZN(n21031) );
  OAI221_X1 U23954 ( .B1(BUF1_REG_26__SCAN_IN), .B2(keyinput46), .C1(n21032), 
        .C2(keyinput33), .A(n21031), .ZN(n21033) );
  NOR4_X1 U23955 ( .A1(n21036), .A2(n21035), .A3(n21034), .A4(n21033), .ZN(
        n21037) );
  NAND4_X1 U23956 ( .A1(n21040), .A2(n21039), .A3(n21038), .A4(n21037), .ZN(
        n21108) );
  AOI22_X1 U23957 ( .A1(n21043), .A2(keyinput26), .B1(n21042), .B2(keyinput23), 
        .ZN(n21041) );
  OAI221_X1 U23958 ( .B1(n21043), .B2(keyinput26), .C1(n21042), .C2(keyinput23), .A(n21041), .ZN(n21056) );
  AOI22_X1 U23959 ( .A1(n21046), .A2(keyinput7), .B1(n21045), .B2(keyinput63), 
        .ZN(n21044) );
  OAI221_X1 U23960 ( .B1(n21046), .B2(keyinput7), .C1(n21045), .C2(keyinput63), 
        .A(n21044), .ZN(n21055) );
  AOI22_X1 U23961 ( .A1(n21049), .A2(keyinput35), .B1(n21048), .B2(keyinput32), 
        .ZN(n21047) );
  OAI221_X1 U23962 ( .B1(n21049), .B2(keyinput35), .C1(n21048), .C2(keyinput32), .A(n21047), .ZN(n21054) );
  INV_X1 U23963 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21051) );
  AOI22_X1 U23964 ( .A1(n21052), .A2(keyinput49), .B1(n21051), .B2(keyinput1), 
        .ZN(n21050) );
  OAI221_X1 U23965 ( .B1(n21052), .B2(keyinput49), .C1(n21051), .C2(keyinput1), 
        .A(n21050), .ZN(n21053) );
  NOR4_X1 U23966 ( .A1(n21056), .A2(n21055), .A3(n21054), .A4(n21053), .ZN(
        n21106) );
  AOI22_X1 U23967 ( .A1(n21059), .A2(keyinput38), .B1(keyinput16), .B2(n21058), 
        .ZN(n21057) );
  OAI221_X1 U23968 ( .B1(n21059), .B2(keyinput38), .C1(n21058), .C2(keyinput16), .A(n21057), .ZN(n21072) );
  AOI22_X1 U23969 ( .A1(n21062), .A2(keyinput41), .B1(n21061), .B2(keyinput2), 
        .ZN(n21060) );
  OAI221_X1 U23970 ( .B1(n21062), .B2(keyinput41), .C1(n21061), .C2(keyinput2), 
        .A(n21060), .ZN(n21071) );
  AOI22_X1 U23971 ( .A1(n21065), .A2(keyinput30), .B1(n21064), .B2(keyinput3), 
        .ZN(n21063) );
  OAI221_X1 U23972 ( .B1(n21065), .B2(keyinput30), .C1(n21064), .C2(keyinput3), 
        .A(n21063), .ZN(n21070) );
  AOI22_X1 U23973 ( .A1(n21068), .A2(keyinput24), .B1(keyinput0), .B2(n21067), 
        .ZN(n21066) );
  OAI221_X1 U23974 ( .B1(n21068), .B2(keyinput24), .C1(n21067), .C2(keyinput0), 
        .A(n21066), .ZN(n21069) );
  NOR4_X1 U23975 ( .A1(n21072), .A2(n21071), .A3(n21070), .A4(n21069), .ZN(
        n21105) );
  AOI22_X1 U23976 ( .A1(n21075), .A2(keyinput57), .B1(keyinput45), .B2(n21074), 
        .ZN(n21073) );
  OAI221_X1 U23977 ( .B1(n21075), .B2(keyinput57), .C1(n21074), .C2(keyinput45), .A(n21073), .ZN(n21086) );
  AOI22_X1 U23978 ( .A1(n14740), .A2(keyinput58), .B1(keyinput11), .B2(n21077), 
        .ZN(n21076) );
  OAI221_X1 U23979 ( .B1(n14740), .B2(keyinput58), .C1(n21077), .C2(keyinput11), .A(n21076), .ZN(n21085) );
  AOI22_X1 U23980 ( .A1(n21079), .A2(keyinput44), .B1(keyinput17), .B2(n12071), 
        .ZN(n21078) );
  OAI221_X1 U23981 ( .B1(n21079), .B2(keyinput44), .C1(n12071), .C2(keyinput17), .A(n21078), .ZN(n21084) );
  AOI22_X1 U23982 ( .A1(n21082), .A2(keyinput4), .B1(n21081), .B2(keyinput62), 
        .ZN(n21080) );
  OAI221_X1 U23983 ( .B1(n21082), .B2(keyinput4), .C1(n21081), .C2(keyinput62), 
        .A(n21080), .ZN(n21083) );
  NOR4_X1 U23984 ( .A1(n21086), .A2(n21085), .A3(n21084), .A4(n21083), .ZN(
        n21104) );
  AOI22_X1 U23985 ( .A1(n21089), .A2(keyinput22), .B1(n21088), .B2(keyinput60), 
        .ZN(n21087) );
  OAI221_X1 U23986 ( .B1(n21089), .B2(keyinput22), .C1(n21088), .C2(keyinput60), .A(n21087), .ZN(n21102) );
  AOI22_X1 U23987 ( .A1(n21092), .A2(keyinput42), .B1(n21091), .B2(keyinput59), 
        .ZN(n21090) );
  OAI221_X1 U23988 ( .B1(n21092), .B2(keyinput42), .C1(n21091), .C2(keyinput59), .A(n21090), .ZN(n21101) );
  INV_X1 U23989 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n21095) );
  AOI22_X1 U23990 ( .A1(n21095), .A2(keyinput12), .B1(keyinput29), .B2(n21094), 
        .ZN(n21093) );
  OAI221_X1 U23991 ( .B1(n21095), .B2(keyinput12), .C1(n21094), .C2(keyinput29), .A(n21093), .ZN(n21100) );
  AOI22_X1 U23992 ( .A1(n21098), .A2(keyinput14), .B1(n21097), .B2(keyinput19), 
        .ZN(n21096) );
  OAI221_X1 U23993 ( .B1(n21098), .B2(keyinput14), .C1(n21097), .C2(keyinput19), .A(n21096), .ZN(n21099) );
  NOR4_X1 U23994 ( .A1(n21102), .A2(n21101), .A3(n21100), .A4(n21099), .ZN(
        n21103) );
  NAND4_X1 U23995 ( .A1(n21106), .A2(n21105), .A3(n21104), .A4(n21103), .ZN(
        n21107) );
  AOI211_X1 U23996 ( .C1(n21110), .C2(n21109), .A(n21108), .B(n21107), .ZN(
        n21111) );
  XNOR2_X1 U23997 ( .A(n21112), .B(n21111), .ZN(P1_U3040) );
  INV_X4 U11235 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9846) );
  CLKBUF_X2 U11440 ( .A(n13472), .Z(n9678) );
  AOI211_X1 U11170 ( .C1(n18188), .C2(n11655), .A(n11654), .B(n11653), .ZN(
        n11677) );
  XNOR2_X1 U11202 ( .A(n12107), .B(n12108), .ZN(n13673) );
  CLKBUF_X1 U11403 ( .A(n14152), .Z(n15832) );
  CLKBUF_X1 U11420 ( .A(n10582), .Z(n19530) );
  CLKBUF_X1 U12317 ( .A(n10581), .Z(n19633) );
  CLKBUF_X1 U12723 ( .A(n11880), .Z(n14096) );
  CLKBUF_X1 U12837 ( .A(n14793), .Z(n15064) );
  AOI211_X1 U12849 ( .C1(n15889), .C2(n14434), .A(n14433), .B(n14432), .ZN(
        n14435) );
  CLKBUF_X1 U14846 ( .A(n16499), .Z(n16511) );
endmodule

