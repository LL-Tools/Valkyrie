

module b21_C_2inp_gates_syn ( P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63 );
  input P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
         P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
         P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
         P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
         P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
         P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
         P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
         P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
         P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
         P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
         P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
         P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
         P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
         P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
         P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
         P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
         P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
         P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
         P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
         P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
         P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
         P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4243, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224;

  INV_X4 U4747 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NAND2_X1 U4748 ( .A1(n9262), .A2(n5643), .ZN(n9340) );
  NAND2_X1 U4749 ( .A1(n6219), .A2(n6218), .ZN(n7761) );
  AND4_X1 U4750 ( .A1(n5217), .A2(n5216), .A3(n5215), .A4(n5214), .ZN(n7519)
         );
  CLKBUF_X2 U4751 ( .A(n6166), .Z(n6443) );
  INV_X2 U4753 ( .A(n5173), .ZN(n5586) );
  INV_X2 U4754 ( .A(n6322), .ZN(n6410) );
  CLKBUF_X2 U4755 ( .A(n6148), .Z(n6421) );
  NAND2_X1 U4756 ( .A1(n6463), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6464) );
  CLKBUF_X2 U4758 ( .A(n4251), .Z(n4440) );
  INV_X1 U4759 ( .A(n9066), .ZN(n4243) );
  INV_X2 U4760 ( .A(n4243), .ZN(P1_U3084) );
  INV_X1 U4761 ( .A(P1_STATE_REG_SCAN_IN), .ZN(n9066) );
  AND2_X1 U4762 ( .A1(n4631), .A2(n4974), .ZN(n4636) );
  INV_X1 U4763 ( .A(n6003), .ZN(n6040) );
  NAND2_X1 U4764 ( .A1(n9438), .A2(n9439), .ZN(n9437) );
  BUF_X1 U4765 ( .A(n6149), .Z(n6444) );
  NAND2_X1 U4766 ( .A1(n6507), .A2(n7813), .ZN(n7823) );
  INV_X1 U4767 ( .A(n8637), .ZN(n7606) );
  AND3_X1 U4768 ( .A1(n5178), .A2(n5177), .A3(n5176), .ZN(n9958) );
  NAND2_X1 U4769 ( .A1(n5616), .A2(n7857), .ZN(n7890) );
  NAND2_X2 U4770 ( .A1(n7182), .A2(n5785), .ZN(n7426) );
  NAND2_X1 U4771 ( .A1(n5119), .A2(n5118), .ZN(n9514) );
  INV_X1 U4772 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n9779) );
  BUF_X1 U4773 ( .A(n6075), .Z(n4250) );
  NAND2_X1 U4774 ( .A1(n5530), .A2(n5529), .ZN(n9541) );
  AND4_X1 U4775 ( .A1(n5195), .A2(n5194), .A3(n5193), .A4(n5192), .ZN(n7532)
         );
  AND2_X1 U4776 ( .A1(n9265), .A2(n5730), .ZN(n9314) );
  OAI211_X1 U4777 ( .C1(n5173), .C2(n6743), .A(n5169), .B(n4891), .ZN(n7400)
         );
  MUX2_X1 U4778 ( .A(n8215), .B(n8214), .S(n8637), .Z(n8216) );
  NAND2_X1 U4779 ( .A1(n5571), .A2(n5570), .ZN(n9315) );
  INV_X1 U4780 ( .A(n5083), .ZN(n8219) );
  INV_X1 U4781 ( .A(n5164), .ZN(n5435) );
  XNOR2_X1 U4782 ( .A(n8189), .B(n8188), .ZN(n8187) );
  AND2_X2 U4783 ( .A1(n4522), .A2(n4521), .ZN(n8189) );
  NAND4_X2 U4784 ( .A1(n6194), .A2(n6193), .A3(n6192), .A4(n6191), .ZN(n8521)
         );
  NAND2_X2 U4785 ( .A1(n7460), .A2(n7459), .ZN(n7492) );
  NOR2_X2 U4786 ( .A1(n5657), .A2(n4889), .ZN(n5069) );
  NAND2_X1 U4787 ( .A1(n7606), .A2(n6709), .ZN(n7235) );
  XNOR2_X2 U4788 ( .A(n5283), .B(n5282), .ZN(n6779) );
  NAND2_X2 U4789 ( .A1(n4963), .A2(n4962), .ZN(n5314) );
  AOI21_X2 U4790 ( .B1(n4636), .B2(n4986), .A(n4635), .ZN(n4634) );
  NOR2_X2 U4791 ( .A1(n4894), .A2(n4897), .ZN(n4986) );
  OR2_X2 U4792 ( .A1(n8566), .A2(n8565), .ZN(n4519) );
  NOR2_X2 U4793 ( .A1(n5197), .A2(P1_IR_REG_5__SCAN_IN), .ZN(n5196) );
  NOR4_X2 U4794 ( .A1(n8807), .A2(n6484), .A3(n8231), .A4(n8037), .ZN(n6485)
         );
  OR2_X2 U4795 ( .A1(n7148), .A2(n7149), .ZN(n4515) );
  INV_X2 U4796 ( .A(n7426), .ZN(n5794) );
  OAI21_X2 U4797 ( .B1(n4824), .B2(n8729), .A(n8240), .ZN(n8721) );
  XNOR2_X2 U4798 ( .A(n6176), .B(P2_IR_REG_4__SCAN_IN), .ZN(n6916) );
  XNOR2_X2 U4799 ( .A(n7761), .B(n10061), .ZN(n7763) );
  NAND2_X2 U4800 ( .A1(n6160), .A2(n6159), .ZN(n6888) );
  NAND2_X1 U4801 ( .A1(n9333), .A2(n9239), .ZN(n9241) );
  AOI21_X1 U4802 ( .B1(n9107), .B2(n9109), .A(n9106), .ZN(n9013) );
  NAND2_X1 U4803 ( .A1(n9306), .A2(n9296), .ZN(n9297) );
  INV_X2 U4804 ( .A(n8618), .ZN(n4772) );
  CLKBUF_X1 U4805 ( .A(n9470), .Z(n4356) );
  NAND2_X1 U4806 ( .A1(n6704), .A2(n6703), .ZN(n7299) );
  NAND2_X1 U4807 ( .A1(n10015), .A2(n10039), .ZN(n7813) );
  NAND2_X1 U4808 ( .A1(n5340), .A2(n5339), .ZN(n9594) );
  INV_X1 U4809 ( .A(n7755), .ZN(n4245) );
  AND2_X1 U4810 ( .A1(n5706), .A2(n7552), .ZN(n7550) );
  NOR2_X1 U4811 ( .A1(n7547), .A2(n5705), .ZN(n7553) );
  NAND2_X2 U4812 ( .A1(n7212), .A2(n7211), .ZN(n7210) );
  NAND2_X1 U4813 ( .A1(n7519), .A2(n7537), .ZN(n5629) );
  INV_X2 U4814 ( .A(n5207), .ZN(n9964) );
  NAND2_X1 U4815 ( .A1(n9156), .A2(n9958), .ZN(n7546) );
  NAND2_X1 U4816 ( .A1(n6134), .A2(n6133), .ZN(n6513) );
  INV_X1 U4817 ( .A(n6630), .ZN(n6624) );
  INV_X1 U4818 ( .A(n7443), .ZN(n7447) );
  AND3_X1 U4819 ( .A1(n6164), .A2(n6163), .A3(n6162), .ZN(n7241) );
  BUF_X4 U4820 ( .A(n6150), .Z(n6273) );
  CLKBUF_X2 U4821 ( .A(n5224), .Z(n5596) );
  INV_X2 U4822 ( .A(n9785), .ZN(n5109) );
  AND4_X2 U4823 ( .A1(n6315), .A2(n6063), .A3(n6104), .A4(n6465), .ZN(n4284)
         );
  OR3_X1 U4824 ( .A1(n5673), .A2(n7188), .A3(n5766), .ZN(n4899) );
  AOI21_X1 U4825 ( .B1(n4569), .B2(n4567), .A(n4564), .ZN(n5673) );
  AOI21_X1 U4826 ( .B1(n4502), .B2(n10080), .A(n4500), .ZN(n8864) );
  OR2_X1 U4827 ( .A1(n5674), .A2(n5650), .ZN(n5651) );
  AND2_X1 U4828 ( .A1(n6013), .A2(n4413), .ZN(n4410) );
  AND2_X1 U4829 ( .A1(n5735), .A2(n5734), .ZN(n5762) );
  NOR2_X1 U4830 ( .A1(n9217), .A2(n9275), .ZN(n9216) );
  NAND2_X1 U4831 ( .A1(n4349), .A2(n4348), .ZN(n9275) );
  INV_X1 U4832 ( .A(n9297), .ZN(n4349) );
  NAND2_X1 U4833 ( .A1(n4519), .A2(n4518), .ZN(n4517) );
  NAND3_X1 U4834 ( .A1(n4457), .A2(n4458), .A3(n4455), .ZN(n9343) );
  AND2_X1 U4835 ( .A1(n9261), .A2(n4459), .ZN(n4458) );
  INV_X1 U4836 ( .A(n9511), .ZN(n4348) );
  NAND2_X1 U4837 ( .A1(n8337), .A2(n8291), .ZN(n8444) );
  NAND2_X1 U4838 ( .A1(n6418), .A2(n6417), .ZN(n8856) );
  NOR2_X1 U4839 ( .A1(n8552), .A2(n4520), .ZN(n8566) );
  NAND2_X1 U4840 ( .A1(n5101), .A2(n5100), .ZN(n9511) );
  OR2_X1 U4841 ( .A1(n9520), .A2(n9288), .ZN(n9265) );
  NOR2_X1 U4842 ( .A1(n4855), .A2(n4398), .ZN(n4397) );
  NAND2_X1 U4843 ( .A1(n4854), .A2(n4859), .ZN(n4853) );
  OR2_X1 U4844 ( .A1(n8861), .A2(n8608), .ZN(n6617) );
  XNOR2_X1 U4845 ( .A(n5117), .B(n5116), .ZN(n9788) );
  NAND2_X1 U4846 ( .A1(n6412), .A2(n6411), .ZN(n8861) );
  OAI21_X1 U4847 ( .B1(n9470), .B2(n4386), .A(n4664), .ZN(n9229) );
  NAND2_X1 U4848 ( .A1(n5575), .A2(n5574), .ZN(n9527) );
  OR2_X1 U4849 ( .A1(n9366), .A2(n9053), .ZN(n5725) );
  OR2_X1 U4850 ( .A1(n9533), .A2(n9140), .ZN(n9262) );
  XNOR2_X1 U4851 ( .A(n5585), .B(n5584), .ZN(n8997) );
  NAND2_X1 U4852 ( .A1(n6401), .A2(n6400), .ZN(n8867) );
  NAND2_X1 U4853 ( .A1(n6391), .A2(n6390), .ZN(n8873) );
  NAND2_X1 U4854 ( .A1(n6375), .A2(n6374), .ZN(n8883) );
  INV_X1 U4855 ( .A(n9288), .ZN(n9322) );
  NAND2_X1 U4856 ( .A1(n5518), .A2(n5517), .ZN(n9366) );
  AND2_X1 U4857 ( .A1(n5514), .A2(n5513), .ZN(n9140) );
  INV_X1 U4858 ( .A(n8692), .ZN(n8888) );
  AOI21_X1 U4859 ( .B1(n7626), .B2(n8051), .A(n7625), .ZN(n7627) );
  AND2_X1 U4860 ( .A1(n6362), .A2(n6361), .ZN(n8692) );
  OR2_X1 U4861 ( .A1(n9051), .A2(n5535), .ZN(n5514) );
  NAND2_X1 U4862 ( .A1(n8137), .A2(n4268), .ZN(n8136) );
  NAND2_X1 U4863 ( .A1(n7876), .A2(n7875), .ZN(n8022) );
  NAND2_X1 U4864 ( .A1(n7492), .A2(n7491), .ZN(n7970) );
  NAND2_X1 U4865 ( .A1(n7367), .A2(n4333), .ZN(n7370) );
  NOR2_X1 U4866 ( .A1(n4877), .A2(n4450), .ZN(n4449) );
  NAND2_X1 U4867 ( .A1(n7270), .A2(n7269), .ZN(n7367) );
  NAND2_X1 U4868 ( .A1(n5466), .A2(n5465), .ZN(n9556) );
  OAI21_X1 U4869 ( .B1(n7299), .B2(n4740), .A(n4737), .ZN(n7460) );
  AND2_X1 U4870 ( .A1(n4515), .A2(n4514), .ZN(n7270) );
  NAND2_X1 U4871 ( .A1(n5020), .A2(n5019), .ZN(n5490) );
  OR2_X2 U4872 ( .A1(n8006), .A2(n9599), .ZN(n8007) );
  NAND2_X1 U4873 ( .A1(n4607), .A2(n4331), .ZN(n5020) );
  NAND2_X1 U4874 ( .A1(n5106), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n5534) );
  AOI21_X1 U4875 ( .B1(n10083), .B2(n7663), .A(n4900), .ZN(n10063) );
  NAND2_X1 U4876 ( .A1(n6343), .A2(n6342), .ZN(n8909) );
  NAND2_X1 U4877 ( .A1(n5438), .A2(n5437), .ZN(n9568) );
  INV_X1 U4878 ( .A(n8228), .ZN(n8028) );
  NAND2_X1 U4879 ( .A1(n7658), .A2(n7657), .ZN(n10083) );
  NAND2_X1 U4880 ( .A1(n6334), .A2(n6333), .ZN(n8915) );
  AOI21_X1 U4881 ( .B1(n4741), .B2(n4739), .A(n4738), .ZN(n4737) );
  NAND2_X1 U4882 ( .A1(n5420), .A2(n5419), .ZN(n9573) );
  AND2_X1 U4883 ( .A1(n7363), .A2(n7357), .ZN(n4741) );
  NOR2_X1 U4884 ( .A1(n9590), .A2(n9594), .ZN(n4755) );
  AND2_X1 U4885 ( .A1(n7854), .A2(n5617), .ZN(n7853) );
  NAND2_X1 U4886 ( .A1(n7028), .A2(n4297), .ZN(n7045) );
  AND2_X1 U4887 ( .A1(n7573), .A2(n7571), .ZN(n7557) );
  NAND2_X1 U4888 ( .A1(n6325), .A2(n6324), .ZN(n8919) );
  OAI21_X1 U4889 ( .B1(n5412), .B2(n5002), .A(n5001), .ZN(n5432) );
  NAND2_X1 U4890 ( .A1(n6289), .A2(n6288), .ZN(n8934) );
  NAND2_X1 U4891 ( .A1(n6282), .A2(n6281), .ZN(n8929) );
  NAND2_X1 U4892 ( .A1(n4828), .A2(n6242), .ZN(n10015) );
  NAND2_X1 U4893 ( .A1(n4998), .A2(n4997), .ZN(n5412) );
  NAND2_X1 U4894 ( .A1(n5287), .A2(n5286), .ZN(n7709) );
  NAND2_X1 U4895 ( .A1(n5361), .A2(n5360), .ZN(n9590) );
  AND2_X1 U4896 ( .A1(n6549), .A2(n6548), .ZN(n10064) );
  NAND2_X2 U4897 ( .A1(n5322), .A2(n5321), .ZN(n9599) );
  NAND2_X1 U4898 ( .A1(n6230), .A2(n6229), .ZN(n8957) );
  AND2_X1 U4899 ( .A1(n5623), .A2(n5622), .ZN(n7549) );
  XNOR2_X1 U4900 ( .A(n5336), .B(n5335), .ZN(n7074) );
  NAND2_X1 U4901 ( .A1(n6252), .A2(n6251), .ZN(n10051) );
  AND2_X1 U4902 ( .A1(n7315), .A2(n7320), .ZN(n7421) );
  XNOR2_X1 U4903 ( .A(n5248), .B(n5247), .ZN(n6747) );
  NAND2_X1 U4904 ( .A1(n7614), .A2(n6538), .ZN(n7597) );
  OR2_X1 U4905 ( .A1(n6111), .A2(n8447), .ZN(n6364) );
  NAND2_X1 U4906 ( .A1(n6909), .A2(n4294), .ZN(n6963) );
  OAI21_X1 U4907 ( .B1(n5334), .B2(n5333), .A(n5332), .ZN(n5336) );
  INV_X1 U4908 ( .A(n7537), .ZN(n9971) );
  XNOR2_X1 U4909 ( .A(n5277), .B(n5276), .ZN(n6756) );
  OAI21_X1 U4910 ( .B1(n5314), .B2(n5313), .A(n5315), .ZN(n5334) );
  INV_X2 U4911 ( .A(n9463), .ZN(n4246) );
  NAND2_X1 U4912 ( .A1(n6894), .A2(n6895), .ZN(n6909) );
  NAND2_X1 U4913 ( .A1(n6198), .A2(n6197), .ZN(n10141) );
  NOR2_X2 U4914 ( .A1(n9201), .A2(n7071), .ZN(n9929) );
  INV_X1 U4915 ( .A(n7739), .ZN(n10138) );
  NAND2_X1 U4916 ( .A1(n6186), .A2(n6185), .ZN(n7739) );
  NAND2_X1 U4917 ( .A1(n6937), .A2(n6938), .ZN(n6936) );
  NAND2_X1 U4918 ( .A1(n4606), .A2(n4945), .ZN(n5234) );
  OR2_X1 U4919 ( .A1(n5348), .A2(n4983), .ZN(n4974) );
  NAND2_X1 U4920 ( .A1(n7331), .A2(n7447), .ZN(n9944) );
  AND4_X1 U4921 ( .A1(n6203), .A2(n6202), .A3(n6201), .A4(n6200), .ZN(n7350)
         );
  XNOR2_X1 U4922 ( .A(n5204), .B(n5203), .ZN(n6726) );
  NAND2_X1 U4923 ( .A1(n4942), .A2(n4941), .ZN(n5219) );
  NAND2_X1 U4924 ( .A1(n5785), .A2(n7183), .ZN(n5786) );
  OR2_X1 U4925 ( .A1(n4982), .A2(n4981), .ZN(n5349) );
  OR2_X1 U4926 ( .A1(n5313), .A2(n4982), .ZN(n5348) );
  INV_X2 U4927 ( .A(n6712), .ZN(n4247) );
  INV_X1 U4928 ( .A(n6702), .ZN(n4742) );
  INV_X2 U4929 ( .A(n7400), .ZN(n9952) );
  CLKBUF_X1 U4930 ( .A(n5694), .Z(n9160) );
  NAND2_X1 U4931 ( .A1(n4367), .A2(n4972), .ZN(n4982) );
  NAND2_X1 U4932 ( .A1(n6948), .A2(n4505), .ZN(n6923) );
  NAND4_X2 U4933 ( .A1(n5141), .A2(n5140), .A3(n5139), .A4(n5138), .ZN(n9161)
         );
  NAND4_X2 U4934 ( .A1(n5149), .A2(n5148), .A3(n5147), .A4(n5146), .ZN(n9158)
         );
  NAND2_X1 U4935 ( .A1(n6949), .A2(n6950), .ZN(n6948) );
  NOR2_X1 U4936 ( .A1(n4863), .A2(n4605), .ZN(n4604) );
  AOI21_X1 U4937 ( .B1(n4864), .B2(n5233), .A(n4862), .ZN(n4861) );
  INV_X1 U4938 ( .A(n4980), .ZN(n5335) );
  NAND2_X1 U4939 ( .A1(n6014), .A2(n5664), .ZN(n5783) );
  XNOR2_X1 U4940 ( .A(n5656), .B(P1_IR_REG_24__SCAN_IN), .ZN(n6014) );
  INV_X1 U4941 ( .A(n5173), .ZN(n4248) );
  NAND2_X1 U4942 ( .A1(n8985), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6083) );
  OAI21_X1 U4943 ( .B1(n5665), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5656) );
  NAND2_X1 U4944 ( .A1(n6466), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6468) );
  NAND2_X1 U4945 ( .A1(n5080), .A2(n9780), .ZN(n9785) );
  NAND2_X1 U4946 ( .A1(n6101), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6341) );
  INV_X2 U4947 ( .A(n8989), .ZN(n9000) );
  MUX2_X1 U4948 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5079), .S(
        P1_IR_REG_29__SCAN_IN), .Z(n5080) );
  XNOR2_X1 U4949 ( .A(n4937), .B(SI_4_), .ZN(n5172) );
  MUX2_X1 U4950 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5074), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n5076) );
  NAND2_X1 U4951 ( .A1(n6081), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6652) );
  INV_X2 U4952 ( .A(n8994), .ZN(n4249) );
  OAI21_X1 U4953 ( .B1(n5660), .B2(P1_IR_REG_26__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5074) );
  CLKBUF_X3 U4954 ( .A(n6075), .Z(n4251) );
  NAND2_X1 U4955 ( .A1(n5071), .A2(n4870), .ZN(n4869) );
  NAND3_X1 U4956 ( .A1(n9207), .A2(n4796), .A3(n4795), .ZN(n4799) );
  NAND3_X1 U4957 ( .A1(n4797), .A2(P1_ADDR_REG_19__SCAN_IN), .A3(
        P2_ADDR_REG_19__SCAN_IN), .ZN(n4798) );
  INV_X1 U4958 ( .A(P1_RD_REG_SCAN_IN), .ZN(n4795) );
  OR2_X1 U4959 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), .ZN(
        n4889) );
  NOR2_X1 U4960 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n6069) );
  AND3_X2 U4961 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n5188) );
  INV_X1 U4962 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n9207) );
  NOR2_X1 U4963 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), .ZN(
        n5066) );
  NOR2_X1 U4964 ( .A1(P2_IR_REG_23__SCAN_IN), .A2(P2_IR_REG_22__SCAN_IN), .ZN(
        n6067) );
  NOR2_X1 U4965 ( .A1(P2_IR_REG_2__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n6068) );
  NOR2_X1 U4966 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n4909) );
  INV_X1 U4967 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n5065) );
  NOR2_X1 U4968 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n4904) );
  INV_X1 U4969 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n5413) );
  INV_X1 U4970 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6239) );
  BUF_X2 U4971 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n9003) );
  INV_X1 U4972 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n5356) );
  INV_X1 U4973 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n6063) );
  INV_X1 U4974 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6096) );
  INV_X1 U4975 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6453) );
  AND2_X2 U4976 ( .A1(n4794), .A2(n4793), .ZN(n4275) );
  NAND2_X1 U4977 ( .A1(n6524), .A2(n6515), .ZN(n7234) );
  AND2_X1 U4978 ( .A1(n6087), .A2(n8993), .ZN(n6166) );
  NOR2_X2 U4979 ( .A1(n7370), .A2(n7371), .ZN(n7625) );
  INV_X1 U4980 ( .A(n6086), .ZN(n8993) );
  INV_X2 U4981 ( .A(n5135), .ZN(n5155) );
  XNOR2_X2 U4982 ( .A(n5590), .B(P1_REG3_REG_27__SCAN_IN), .ZN(n9307) );
  NAND2_X1 U4983 ( .A1(n5135), .A2(n4252), .ZN(n5173) );
  NOR2_X2 U4984 ( .A1(n4752), .A2(n8007), .ZN(n9208) );
  XNOR2_X1 U4985 ( .A(n4640), .B(n7277), .ZN(n7187) );
  BUF_X4 U4986 ( .A(n6075), .Z(n4252) );
  NAND2_X2 U4987 ( .A1(n4799), .A2(n4798), .ZN(n6075) );
  AND2_X1 U4988 ( .A1(n6504), .A2(n6507), .ZN(n6556) );
  NAND2_X1 U4989 ( .A1(n4592), .A2(n4591), .ZN(n6504) );
  NAND2_X1 U4990 ( .A1(n6505), .A2(n6624), .ZN(n4592) );
  NOR2_X1 U4991 ( .A1(n5247), .A2(n4865), .ZN(n4864) );
  INV_X1 U4992 ( .A(n4948), .ZN(n4865) );
  NAND2_X1 U4993 ( .A1(n8022), .A2(n8021), .ZN(n8027) );
  AND2_X1 U4994 ( .A1(n8037), .A2(n8035), .ZN(n8021) );
  INV_X1 U4995 ( .A(n6565), .ZN(n4504) );
  OR2_X1 U4996 ( .A1(n9514), .A2(n9318), .ZN(n9266) );
  AND2_X1 U4997 ( .A1(n7642), .A2(n9277), .ZN(n6051) );
  INV_X1 U4998 ( .A(n5568), .ZN(n5592) );
  INV_X1 U4999 ( .A(n5563), .ZN(n5535) );
  BUF_X1 U5000 ( .A(n5256), .Z(n5568) );
  NAND2_X1 U5001 ( .A1(n9785), .A2(n5083), .ZN(n5256) );
  AND2_X1 U5002 ( .A1(n6556), .A2(n6555), .ZN(n6563) );
  OAI21_X1 U5003 ( .B1(n5679), .B2(n5608), .A(n4552), .ZN(n4551) );
  NAND2_X1 U5004 ( .A1(n4553), .A2(n5608), .ZN(n4552) );
  NAND2_X1 U5005 ( .A1(n5613), .A2(n9251), .ZN(n4553) );
  NAND2_X1 U5006 ( .A1(n4600), .A2(n5003), .ZN(n4599) );
  NAND2_X1 U5007 ( .A1(n5002), .A2(n5001), .ZN(n4600) );
  AOI21_X1 U5008 ( .B1(n4603), .B2(n4861), .A(n4315), .ZN(n4602) );
  OR2_X1 U5009 ( .A1(n5284), .A2(P1_IR_REG_9__SCAN_IN), .ZN(n5358) );
  NAND2_X1 U5010 ( .A1(n4950), .A2(n4949), .ZN(n4953) );
  OR2_X1 U5011 ( .A1(n8856), .A2(n8355), .ZN(n6620) );
  NAND2_X1 U5012 ( .A1(n4772), .A2(n6615), .ZN(n4771) );
  INV_X1 U5013 ( .A(n4770), .ZN(n4769) );
  OAI21_X1 U5014 ( .B1(n4901), .B2(n4771), .A(n6617), .ZN(n4770) );
  OR2_X1 U5015 ( .A1(n8867), .A2(n8321), .ZN(n6613) );
  NAND2_X1 U5016 ( .A1(n8867), .A2(n8321), .ZN(n6615) );
  OR2_X1 U5017 ( .A1(n8681), .A2(n4857), .ZN(n4854) );
  INV_X1 U5018 ( .A(n4860), .ZN(n4857) );
  NAND2_X1 U5019 ( .A1(n8721), .A2(n4401), .ZN(n4399) );
  AND2_X1 U5020 ( .A1(n4404), .A2(n8727), .ZN(n4401) );
  OR2_X1 U5021 ( .A1(n8898), .A2(n8744), .ZN(n8710) );
  OR2_X1 U5022 ( .A1(n8915), .A2(n8477), .ZN(n6498) );
  OR2_X1 U5023 ( .A1(n8934), .A2(n8068), .ZN(n6568) );
  INV_X1 U5024 ( .A(n8049), .ZN(n4802) );
  INV_X1 U5025 ( .A(n8828), .ZN(n4812) );
  AND2_X1 U5026 ( .A1(n8247), .A2(n4473), .ZN(n8636) );
  INV_X1 U5027 ( .A(n8867), .ZN(n4473) );
  INV_X1 U5028 ( .A(n6548), .ZN(n4490) );
  AND2_X1 U5029 ( .A1(n9075), .A2(n4709), .ZN(n4707) );
  INV_X1 U5030 ( .A(n5930), .ZN(n4709) );
  NAND2_X1 U5031 ( .A1(n7788), .A2(n5880), .ZN(n5898) );
  OR2_X1 U5032 ( .A1(n9496), .A2(n9213), .ZN(n5611) );
  AND2_X1 U5033 ( .A1(n9263), .A2(n9262), .ZN(n4888) );
  OR2_X1 U5034 ( .A1(n9541), .A2(n9387), .ZN(n9234) );
  OAI21_X1 U5035 ( .B1(n4668), .B2(n4257), .A(n4290), .ZN(n4665) );
  AND2_X1 U5036 ( .A1(n9478), .A2(n4879), .ZN(n4878) );
  NAND2_X1 U5037 ( .A1(n9245), .A2(n9244), .ZN(n4879) );
  OR2_X1 U5038 ( .A1(n9580), .A2(n9483), .ZN(n9244) );
  NOR2_X1 U5039 ( .A1(n4651), .A2(n4650), .ZN(n4649) );
  INV_X1 U5040 ( .A(n7842), .ZN(n4650) );
  INV_X1 U5041 ( .A(n4652), .ZN(n4651) );
  AND2_X1 U5042 ( .A1(n7993), .A2(n4444), .ZN(n7841) );
  OR2_X1 U5043 ( .A1(n9599), .A2(n7893), .ZN(n7854) );
  NAND2_X1 U5044 ( .A1(n5170), .A2(n5700), .ZN(n7555) );
  INV_X1 U5045 ( .A(n4610), .ZN(n4609) );
  OAI21_X1 U5046 ( .B1(n4614), .B2(n4611), .A(n5055), .ZN(n4610) );
  OAI21_X1 U5047 ( .B1(n5505), .B2(n5504), .A(n5037), .ZN(n5573) );
  AND2_X1 U5048 ( .A1(n5042), .A2(n5041), .ZN(n5572) );
  NAND2_X1 U5049 ( .A1(n5011), .A2(n5010), .ZN(n5464) );
  NAND2_X1 U5050 ( .A1(n4594), .A2(n4299), .ZN(n5011) );
  INV_X1 U5051 ( .A(n5450), .ZN(n4593) );
  AND2_X1 U5052 ( .A1(n5016), .A2(n5015), .ZN(n5463) );
  NOR2_X1 U5053 ( .A1(n4638), .A2(n5377), .ZN(n4637) );
  INV_X1 U5054 ( .A(n4986), .ZN(n4638) );
  INV_X1 U5055 ( .A(n4992), .ZN(n4635) );
  INV_X1 U5056 ( .A(n5377), .ZN(n4631) );
  NAND2_X1 U5057 ( .A1(n5163), .A2(n5162), .ZN(n4831) );
  NOR2_X1 U5058 ( .A1(n6210), .A2(n6209), .ZN(n6221) );
  OAI21_X1 U5059 ( .B1(n8444), .B2(n4734), .A(n4731), .ZN(n8304) );
  INV_X1 U5060 ( .A(n4735), .ZN(n4734) );
  AND2_X1 U5061 ( .A1(n6680), .A2(n6679), .ZN(n10022) );
  NAND2_X1 U5062 ( .A1(n4718), .A2(n4717), .ZN(n8353) );
  AOI21_X1 U5063 ( .B1(n4719), .B2(n8387), .A(n4283), .ZN(n4717) );
  INV_X1 U5064 ( .A(n6421), .ZN(n6435) );
  INV_X1 U5065 ( .A(n6166), .ZN(n6388) );
  NAND2_X1 U5066 ( .A1(n8988), .A2(n6086), .ZN(n6148) );
  XNOR2_X1 U5067 ( .A(n4517), .B(n4516), .ZN(n8580) );
  NAND2_X1 U5068 ( .A1(n4836), .A2(n4843), .ZN(n4835) );
  OAI21_X1 U5069 ( .B1(n4840), .B2(n4842), .A(n8618), .ZN(n4836) );
  INV_X1 U5070 ( .A(n4843), .ZN(n4837) );
  AOI21_X1 U5071 ( .B1(n4483), .B2(n4485), .A(n8235), .ZN(n4481) );
  INV_X1 U5072 ( .A(n4486), .ZN(n4485) );
  NAND2_X1 U5073 ( .A1(n6314), .A2(n6574), .ZN(n4482) );
  NAND2_X1 U5074 ( .A1(n8027), .A2(n4260), .ZN(n4832) );
  OR2_X1 U5075 ( .A1(n8924), .A2(n8270), .ZN(n6574) );
  NAND2_X1 U5076 ( .A1(n4828), .A2(n4826), .ZN(n6507) );
  NOR2_X1 U5077 ( .A1(n10039), .A2(n4827), .ZN(n4826) );
  INV_X1 U5078 ( .A(n6242), .ZN(n4827) );
  INV_X1 U5079 ( .A(n8844), .ZN(n8259) );
  AND2_X1 U5080 ( .A1(n7508), .A2(n6710), .ZN(n8903) );
  AND2_X1 U5081 ( .A1(n5500), .A2(n5499), .ZN(n9038) );
  OR2_X1 U5082 ( .A1(n9511), .A2(n9287), .ZN(n5612) );
  NAND2_X1 U5083 ( .A1(n4673), .A2(n4678), .ZN(n9502) );
  AND2_X1 U5084 ( .A1(n9292), .A2(n9242), .ZN(n4678) );
  AND2_X1 U5085 ( .A1(n5126), .A2(n5125), .ZN(n9318) );
  OR2_X1 U5086 ( .A1(n9294), .A2(n5535), .ZN(n5126) );
  NAND2_X1 U5087 ( .A1(n5589), .A2(n5588), .ZN(n9520) );
  NAND2_X1 U5088 ( .A1(n8997), .A2(n5586), .ZN(n5589) );
  NOR2_X2 U5089 ( .A1(n9327), .A2(n9527), .ZN(n9209) );
  NAND2_X1 U5090 ( .A1(n9343), .A2(n4888), .ZN(n9311) );
  AND2_X1 U5091 ( .A1(n9343), .A2(n9262), .ZN(n9321) );
  NOR2_X1 U5092 ( .A1(n9556), .A2(n9440), .ZN(n9230) );
  NOR2_X1 U5093 ( .A1(n9252), .A2(n4873), .ZN(n4872) );
  OR2_X1 U5094 ( .A1(n9573), .A2(n9125), .ZN(n9247) );
  NAND2_X1 U5095 ( .A1(n7191), .A2(n7190), .ZN(n9454) );
  INV_X1 U5096 ( .A(n9519), .ZN(n9522) );
  AND2_X1 U5097 ( .A1(n6033), .A2(n7328), .ZN(n9607) );
  OR2_X1 U5098 ( .A1(n5081), .A2(n9779), .ZN(n5082) );
  AOI21_X1 U5099 ( .B1(n4780), .B2(n4285), .A(n4773), .ZN(n6462) );
  OAI21_X1 U5100 ( .B1(n4775), .B2(n4777), .A(n4774), .ZN(n4773) );
  NAND2_X1 U5101 ( .A1(n4584), .A2(n4585), .ZN(n4582) );
  NAND2_X1 U5102 ( .A1(n6657), .A2(n7508), .ZN(n4585) );
  AND2_X1 U5103 ( .A1(n4892), .A2(n6013), .ZN(n4701) );
  MUX2_X1 U5104 ( .A(n6512), .B(n6511), .S(n6624), .Z(n6564) );
  AND2_X1 U5105 ( .A1(n8028), .A2(n6569), .ZN(n4578) );
  NAND2_X1 U5106 ( .A1(n4580), .A2(n4579), .ZN(n6596) );
  AND2_X1 U5107 ( .A1(n6580), .A2(n6582), .ZN(n4579) );
  NAND2_X1 U5108 ( .A1(n4261), .A2(n4550), .ZN(n4549) );
  NAND2_X1 U5109 ( .A1(n5678), .A2(n7096), .ZN(n4550) );
  AND2_X1 U5110 ( .A1(n5614), .A2(n5615), .ZN(n4554) );
  NOR2_X1 U5111 ( .A1(n4551), .A2(n5548), .ZN(n4548) );
  INV_X1 U5112 ( .A(n4549), .ZN(n4545) );
  INV_X1 U5113 ( .A(n4548), .ZN(n4546) );
  OAI21_X1 U5114 ( .B1(n4252), .B2(P1_DATAO_REG_13__SCAN_IN), .A(n4385), .ZN(
        n4967) );
  NAND2_X1 U5115 ( .A1(n4251), .A2(n4965), .ZN(n4385) );
  INV_X1 U5116 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n4965) );
  NOR4_X1 U5117 ( .A1(n7825), .A2(n6482), .A3(n7823), .A4(n7668), .ZN(n6483)
         );
  NOR2_X1 U5118 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n4478) );
  NOR2_X1 U5119 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n4479) );
  NOR2_X1 U5120 ( .A1(n4696), .A2(n4694), .ZN(n4693) );
  INV_X1 U5121 ( .A(n9095), .ZN(n4694) );
  INV_X1 U5122 ( .A(n9033), .ZN(n4696) );
  OR2_X1 U5123 ( .A1(n9568), .A2(n9485), .ZN(n5615) );
  NAND2_X1 U5124 ( .A1(n5007), .A2(n5006), .ZN(n5010) );
  INV_X1 U5125 ( .A(n4637), .ZN(n4629) );
  INV_X1 U5126 ( .A(n4895), .ZN(n4633) );
  NAND2_X1 U5127 ( .A1(n4252), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n4379) );
  NAND2_X1 U5128 ( .A1(n5219), .A2(n4943), .ZN(n4606) );
  INV_X1 U5129 ( .A(n4935), .ZN(n4829) );
  OR2_X1 U5130 ( .A1(n8852), .A2(n8607), .ZN(n6625) );
  NAND2_X1 U5131 ( .A1(n8624), .A2(n8608), .ZN(n4843) );
  AND2_X1 U5132 ( .A1(n8888), .A2(n8677), .ZN(n6496) );
  AND2_X1 U5133 ( .A1(n8692), .A2(n8715), .ZN(n6588) );
  NAND2_X1 U5134 ( .A1(n4317), .A2(n4404), .ZN(n4400) );
  NOR2_X1 U5135 ( .A1(n8711), .A2(n4782), .ZN(n4781) );
  OAI21_X1 U5136 ( .B1(n8235), .B2(n4850), .A(n8239), .ZN(n4849) );
  NAND2_X1 U5137 ( .A1(n4763), .A2(n6507), .ZN(n4762) );
  INV_X1 U5138 ( .A(n6553), .ZN(n4763) );
  INV_X1 U5139 ( .A(n6557), .ZN(n4761) );
  NOR2_X1 U5140 ( .A1(n7763), .A2(n4393), .ZN(n4392) );
  INV_X1 U5141 ( .A(n7664), .ZN(n4393) );
  INV_X1 U5142 ( .A(n7762), .ZN(n4391) );
  OR2_X1 U5143 ( .A1(n10051), .A2(n10008), .ZN(n6557) );
  OAI21_X1 U5144 ( .B1(n6421), .B2(P2_REG3_REG_3__SCAN_IN), .A(n6117), .ZN(
        n4499) );
  OR2_X1 U5145 ( .A1(n10102), .A2(n7221), .ZN(n7599) );
  AND2_X1 U5146 ( .A1(n8903), .A2(n7621), .ZN(n7222) );
  OR2_X1 U5147 ( .A1(n6183), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n6204) );
  NOR2_X1 U5148 ( .A1(n4433), .A2(n4430), .ZN(n4429) );
  INV_X1 U5149 ( .A(n5854), .ZN(n4430) );
  NOR2_X1 U5150 ( .A1(n7646), .A2(n5860), .ZN(n4433) );
  NAND2_X1 U5151 ( .A1(n4425), .A2(n4424), .ZN(n5962) );
  NOR2_X1 U5152 ( .A1(n4426), .A2(n4304), .ZN(n4424) );
  NAND2_X1 U5153 ( .A1(n5825), .A2(n4266), .ZN(n7510) );
  NAND2_X1 U5154 ( .A1(n4685), .A2(n4688), .ZN(n5914) );
  AND2_X1 U5155 ( .A1(n4689), .A2(n5907), .ZN(n4688) );
  INV_X1 U5156 ( .A(n5532), .ZN(n5106) );
  INV_X1 U5157 ( .A(n4384), .ZN(n5521) );
  INV_X1 U5158 ( .A(n4645), .ZN(n4644) );
  OAI21_X1 U5159 ( .B1(n9405), .B2(n4646), .A(n9233), .ZN(n4645) );
  INV_X1 U5160 ( .A(n9232), .ZN(n4646) );
  INV_X1 U5161 ( .A(n4667), .ZN(n4386) );
  AND2_X1 U5162 ( .A1(n9580), .A2(n9483), .ZN(n9245) );
  NAND2_X1 U5163 ( .A1(n9225), .A2(n9224), .ZN(n9470) );
  AND2_X1 U5164 ( .A1(n8107), .A2(n7855), .ZN(n4883) );
  NOR2_X1 U5165 ( .A1(n8097), .A2(n4653), .ZN(n4652) );
  INV_X1 U5166 ( .A(n7844), .ZN(n4653) );
  INV_X1 U5167 ( .A(n4657), .ZN(n4656) );
  OAI21_X1 U5168 ( .B1(n7543), .B2(n4658), .A(n4661), .ZN(n4657) );
  INV_X1 U5169 ( .A(n7557), .ZN(n7543) );
  INV_X1 U5170 ( .A(n7308), .ZN(n5705) );
  AOI21_X1 U5171 ( .B1(n4616), .B2(n5116), .A(n4335), .ZN(n4615) );
  INV_X1 U5172 ( .A(n5049), .ZN(n4616) );
  INV_X1 U5173 ( .A(n5116), .ZN(n4617) );
  INV_X1 U5174 ( .A(n4869), .ZN(n4663) );
  NAND2_X1 U5175 ( .A1(n5043), .A2(n5042), .ZN(n5585) );
  AND2_X1 U5176 ( .A1(n5049), .A2(n5048), .ZN(n5584) );
  NAND2_X1 U5177 ( .A1(n4620), .A2(n4619), .ZN(n5505) );
  AOI21_X1 U5178 ( .B1(n4621), .B2(n4622), .A(n4336), .ZN(n4619) );
  AOI21_X1 U5179 ( .B1(n5527), .B2(n4626), .A(n4625), .ZN(n4624) );
  INV_X1 U5180 ( .A(n5024), .ZN(n4626) );
  INV_X1 U5181 ( .A(n5030), .ZN(n4625) );
  NAND2_X1 U5182 ( .A1(n5527), .A2(n4623), .ZN(n4622) );
  INV_X1 U5183 ( .A(n5489), .ZN(n4623) );
  NAND2_X1 U5184 ( .A1(n5464), .A2(n5463), .ZN(n4607) );
  INV_X1 U5185 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n4912) );
  AND2_X1 U5186 ( .A1(n5196), .A2(n5068), .ZN(n4914) );
  INV_X1 U5187 ( .A(n4598), .ZN(n4597) );
  OAI21_X1 U5188 ( .B1(n4599), .B2(n5001), .A(n5005), .ZN(n4598) );
  INV_X1 U5189 ( .A(n4599), .ZN(n4595) );
  NOR2_X1 U5190 ( .A1(n4983), .A2(n5349), .ZN(n4894) );
  XNOR2_X1 U5191 ( .A(n4977), .B(SI_11_), .ZN(n5301) );
  OR2_X1 U5192 ( .A1(n4961), .A2(n4960), .ZN(n4962) );
  NAND2_X1 U5193 ( .A1(n4954), .A2(n9632), .ZN(n5278) );
  NAND2_X1 U5194 ( .A1(n4952), .A2(n4953), .ZN(n5247) );
  NAND2_X1 U5195 ( .A1(n6143), .A2(SI_1_), .ZN(n4807) );
  NOR2_X1 U5196 ( .A1(n6728), .A2(n5132), .ZN(n4808) );
  NAND2_X1 U5197 ( .A1(n4808), .A2(n5133), .ZN(n4805) );
  NOR2_X1 U5198 ( .A1(n10012), .A2(n4716), .ZN(n4715) );
  INV_X1 U5199 ( .A(n7969), .ZN(n4716) );
  NAND2_X1 U5200 ( .A1(n6779), .A2(n6457), .ZN(n4828) );
  AND2_X1 U5201 ( .A1(n8305), .A2(n8308), .ZN(n8416) );
  NAND2_X1 U5202 ( .A1(n4713), .A2(n10022), .ZN(n10027) );
  INV_X1 U5203 ( .A(n7298), .ZN(n4739) );
  INV_X1 U5204 ( .A(n7457), .ZN(n4738) );
  OR2_X1 U5205 ( .A1(n6675), .A2(n10020), .ZN(n6677) );
  INV_X1 U5206 ( .A(n8276), .ZN(n4725) );
  INV_X1 U5207 ( .A(n8281), .ZN(n4724) );
  AND2_X1 U5208 ( .A1(n8411), .A2(n4729), .ZN(n4728) );
  NAND2_X1 U5209 ( .A1(n8271), .A2(n8276), .ZN(n4729) );
  NOR2_X1 U5210 ( .A1(n6456), .A2(n4338), .ZN(n4778) );
  INV_X1 U5211 ( .A(n6626), .ZN(n4776) );
  AND2_X1 U5212 ( .A1(n6427), .A2(n6426), .ZN(n8355) );
  AND3_X1 U5213 ( .A1(n6340), .A2(n6339), .A3(n6338), .ZN(n8477) );
  AND3_X1 U5214 ( .A1(n6330), .A2(n6329), .A3(n6328), .ZN(n8501) );
  AND4_X1 U5215 ( .A1(n6215), .A2(n6214), .A3(n6213), .A4(n6212), .ZN(n7464)
         );
  OR2_X1 U5216 ( .A1(n7627), .A2(n7628), .ZN(n4522) );
  NAND2_X1 U5217 ( .A1(n8204), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n4518) );
  AND2_X1 U5218 ( .A1(n6625), .A2(n6626), .ZN(n8244) );
  AND2_X1 U5219 ( .A1(n4835), .A2(n8605), .ZN(n4833) );
  INV_X1 U5220 ( .A(n8244), .ZN(n8221) );
  NAND2_X1 U5221 ( .A1(n4768), .A2(n4767), .ZN(n8610) );
  AOI21_X1 U5222 ( .B1(n4769), .B2(n4771), .A(n8605), .ZN(n4767) );
  NAND2_X1 U5223 ( .A1(n8636), .A2(n4820), .ZN(n8601) );
  INV_X1 U5224 ( .A(n4822), .ZN(n4820) );
  NAND2_X1 U5225 ( .A1(n8636), .A2(n8624), .ZN(n8619) );
  NOR2_X1 U5226 ( .A1(n8632), .A2(n8646), .ZN(n4842) );
  INV_X1 U5227 ( .A(n4845), .ZN(n4841) );
  NAND2_X1 U5228 ( .A1(n8631), .A2(n6615), .ZN(n4503) );
  OR2_X1 U5229 ( .A1(n8873), .A2(n8661), .ZN(n8630) );
  AND2_X1 U5230 ( .A1(n6613), .A2(n6615), .ZN(n8632) );
  NAND2_X1 U5231 ( .A1(n8644), .A2(n4901), .ZN(n8631) );
  NOR2_X1 U5232 ( .A1(n8873), .A2(n4846), .ZN(n4845) );
  AND2_X1 U5233 ( .A1(n6402), .A2(n6395), .ZN(n8650) );
  OR2_X1 U5234 ( .A1(n8667), .A2(n8512), .ZN(n8241) );
  INV_X1 U5235 ( .A(n8663), .ZN(n8657) );
  NAND2_X1 U5236 ( .A1(n8664), .A2(n8663), .ZN(n8662) );
  NAND2_X1 U5237 ( .A1(n8692), .A2(n8677), .ZN(n4860) );
  INV_X1 U5238 ( .A(n4854), .ZN(n4856) );
  NAND2_X1 U5239 ( .A1(n4399), .A2(n4400), .ZN(n8688) );
  OR2_X1 U5240 ( .A1(n4786), .A2(n6360), .ZN(n4784) );
  NAND2_X1 U5241 ( .A1(n8797), .A2(n4289), .ZN(n8751) );
  OR2_X1 U5242 ( .A1(n8755), .A2(n8760), .ZN(n4851) );
  AND2_X1 U5243 ( .A1(n6594), .A2(n8709), .ZN(n8738) );
  AOI21_X1 U5244 ( .B1(n4271), .B2(n6574), .A(n4487), .ZN(n4486) );
  INV_X1 U5245 ( .A(n6579), .ZN(n4487) );
  NAND2_X1 U5246 ( .A1(n4832), .A2(n4281), .ZN(n8806) );
  AND2_X1 U5247 ( .A1(n6568), .A2(n8142), .ZN(n4352) );
  NAND2_X1 U5248 ( .A1(n6574), .A2(n6573), .ZN(n8231) );
  OR2_X1 U5249 ( .A1(n8929), .A2(n8499), .ZN(n8142) );
  AND3_X1 U5250 ( .A1(n6312), .A2(n6311), .A3(n6310), .ZN(n8270) );
  NAND2_X1 U5251 ( .A1(n6268), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6308) );
  NAND2_X1 U5252 ( .A1(n6253), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6270) );
  NAND2_X1 U5253 ( .A1(n10057), .A2(n10064), .ZN(n10056) );
  OR2_X1 U5254 ( .A1(n10088), .A2(n10072), .ZN(n10069) );
  NOR2_X1 U5255 ( .A1(n4810), .A2(n8434), .ZN(n4809) );
  AND2_X1 U5256 ( .A1(n6178), .A2(n6177), .ZN(n7610) );
  NAND2_X1 U5257 ( .A1(n8826), .A2(n10128), .ZN(n8828) );
  INV_X1 U5258 ( .A(n10080), .ZN(n8820) );
  AND2_X1 U5259 ( .A1(n4890), .A2(n7241), .ZN(n8826) );
  AND2_X1 U5260 ( .A1(n6855), .A2(n6655), .ZN(n10058) );
  INV_X1 U5261 ( .A(n8823), .ZN(n10060) );
  NAND2_X1 U5262 ( .A1(n7236), .A2(n7235), .ZN(n10080) );
  AND2_X1 U5263 ( .A1(n6131), .A2(n4406), .ZN(n4896) );
  INV_X1 U5264 ( .A(n8247), .ZN(n8649) );
  NAND2_X1 U5265 ( .A1(n6077), .A2(n6076), .ZN(n8898) );
  INV_X1 U5266 ( .A(n10149), .ZN(n8950) );
  INV_X1 U5267 ( .A(n6126), .ZN(n10128) );
  INV_X1 U5268 ( .A(n6702), .ZN(n10116) );
  OAI211_X1 U5269 ( .C1(n6082), .C2(n4496), .A(n4493), .B(n4491), .ZN(n6086)
         );
  NAND2_X1 U5270 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n6085), .ZN(n4496) );
  NAND2_X1 U5271 ( .A1(n4495), .A2(n4494), .ZN(n4493) );
  NAND2_X1 U5272 ( .A1(n6082), .A2(n4492), .ZN(n4491) );
  NOR2_X1 U5273 ( .A1(n4417), .A2(n4418), .ZN(n4416) );
  NAND2_X1 U5274 ( .A1(n6012), .A2(n4259), .ZN(n4414) );
  NAND2_X1 U5275 ( .A1(n4705), .A2(n4704), .ZN(n4703) );
  NOR2_X1 U5276 ( .A1(n6044), .A2(n9132), .ZN(n4704) );
  INV_X1 U5277 ( .A(n4898), .ZN(n4705) );
  INV_X1 U5278 ( .A(n5815), .ZN(n4683) );
  AND2_X1 U5279 ( .A1(n5797), .A2(n5796), .ZN(n7067) );
  NAND2_X1 U5280 ( .A1(n7067), .A2(n7066), .ZN(n7065) );
  NAND2_X1 U5281 ( .A1(n5962), .A2(n9095), .ZN(n9098) );
  NAND2_X1 U5282 ( .A1(n5898), .A2(n5897), .ZN(n7948) );
  INV_X1 U5283 ( .A(n4416), .ZN(n4413) );
  NAND2_X1 U5284 ( .A1(n5604), .A2(n5605), .ZN(n4570) );
  MUX2_X1 U5285 ( .A(n5127), .B(n5675), .S(n7096), .Z(n5605) );
  NAND2_X1 U5286 ( .A1(n5769), .A2(n5608), .ZN(n4565) );
  NAND2_X1 U5287 ( .A1(n5607), .A2(n4568), .ZN(n4566) );
  INV_X1 U5288 ( .A(n5761), .ZN(n4568) );
  NOR2_X1 U5289 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(n9779), .ZN(n4437) );
  NAND2_X1 U5290 ( .A1(n4913), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5609) );
  AND2_X1 U5291 ( .A1(n4420), .A2(n4422), .ZN(n4419) );
  NAND2_X1 U5292 ( .A1(n5611), .A2(n5096), .ZN(n5769) );
  OR2_X1 U5293 ( .A1(n9496), .A2(n5610), .ZN(n5096) );
  OR2_X1 U5294 ( .A1(n5256), .A2(n6787), .ZN(n5158) );
  OR2_X1 U5295 ( .A1(n7133), .A2(n7134), .ZN(n7131) );
  OR2_X1 U5296 ( .A1(n7137), .A2(n7138), .ZN(n7135) );
  NAND2_X1 U5297 ( .A1(n4529), .A2(n4528), .ZN(n6845) );
  AOI21_X1 U5298 ( .B1(n4253), .B2(n7138), .A(n4302), .ZN(n4528) );
  OR2_X1 U5299 ( .A1(n7112), .A2(n7111), .ZN(n7109) );
  OAI21_X1 U5300 ( .B1(n9839), .B2(P1_REG1_REG_12__SCAN_IN), .A(n9835), .ZN(
        n9854) );
  AOI21_X1 U5301 ( .B1(n9197), .B2(n9924), .A(n9920), .ZN(n9198) );
  INV_X1 U5302 ( .A(n9242), .ZN(n4676) );
  INV_X1 U5303 ( .A(n9314), .ZN(n4679) );
  INV_X1 U5304 ( .A(n4888), .ZN(n4887) );
  AOI21_X1 U5305 ( .B1(n9337), .B2(n9238), .A(n9237), .ZN(n9333) );
  NAND2_X1 U5306 ( .A1(n9322), .A2(n9449), .ZN(n9324) );
  NAND2_X1 U5307 ( .A1(n4460), .A2(n9256), .ZN(n4457) );
  NAND2_X1 U5308 ( .A1(n4456), .A2(n9386), .ZN(n4455) );
  NAND2_X1 U5309 ( .A1(n9406), .A2(n9405), .ZN(n9404) );
  AOI21_X1 U5310 ( .B1(n4668), .B2(n9227), .A(n4257), .ZN(n4667) );
  AND2_X1 U5311 ( .A1(n5614), .A2(n9251), .ZN(n9439) );
  NAND2_X1 U5312 ( .A1(n4353), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n5455) );
  NAND2_X1 U5313 ( .A1(n4672), .A2(n4671), .ZN(n4670) );
  NOR2_X1 U5314 ( .A1(n4301), .A2(n4880), .ZN(n4874) );
  NAND2_X1 U5315 ( .A1(n4875), .A2(n4878), .ZN(n9487) );
  NAND2_X1 U5316 ( .A1(n9246), .A2(n9244), .ZN(n4875) );
  NAND2_X1 U5317 ( .A1(n4383), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n5421) );
  AND3_X1 U5318 ( .A1(n5426), .A2(n5425), .A3(n5424), .ZN(n9125) );
  AND3_X1 U5319 ( .A1(n5390), .A2(n5389), .A3(n5388), .ZN(n9067) );
  NAND2_X1 U5320 ( .A1(n5104), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n5342) );
  INV_X1 U5321 ( .A(n5324), .ZN(n5104) );
  NAND2_X1 U5322 ( .A1(n7843), .A2(n7842), .ZN(n7888) );
  AOI21_X1 U5323 ( .B1(n7853), .B2(n5370), .A(n4443), .ZN(n4442) );
  INV_X1 U5324 ( .A(n7854), .ZN(n4443) );
  OR2_X1 U5325 ( .A1(n7840), .A2(n7839), .ZN(n7993) );
  AND4_X1 U5326 ( .A1(n5347), .A2(n5346), .A3(n5345), .A4(n5344), .ZN(n8125)
         );
  NAND2_X1 U5327 ( .A1(n5289), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n5324) );
  NAND2_X1 U5328 ( .A1(n5103), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n5268) );
  INV_X1 U5329 ( .A(n5254), .ZN(n5103) );
  OR2_X1 U5330 ( .A1(n9981), .A2(n7750), .ZN(n7573) );
  NAND2_X1 U5331 ( .A1(n7572), .A2(n7571), .ZN(n7718) );
  NAND2_X1 U5332 ( .A1(n4662), .A2(n7543), .ZN(n7570) );
  INV_X1 U5333 ( .A(n7544), .ZN(n4662) );
  INV_X1 U5334 ( .A(n9451), .ZN(n9482) );
  AND2_X1 U5335 ( .A1(n7189), .A2(n7642), .ZN(n7278) );
  INV_X1 U5336 ( .A(n9484), .ZN(n9449) );
  OR2_X1 U5337 ( .A1(n7194), .A2(n7195), .ZN(n9484) );
  INV_X1 U5338 ( .A(n9272), .ZN(n9273) );
  AOI21_X1 U5339 ( .B1(n9271), .B2(n9451), .A(n9270), .ZN(n9272) );
  NAND2_X1 U5340 ( .A1(n5479), .A2(n5478), .ZN(n9552) );
  NAND2_X1 U5341 ( .A1(n5453), .A2(n5452), .ZN(n9561) );
  OR2_X1 U5342 ( .A1(n5173), .A2(n6730), .ZN(n5178) );
  INV_X1 U5343 ( .A(n9984), .ZN(n9945) );
  NAND2_X1 U5344 ( .A1(n5164), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4641) );
  NAND2_X1 U5345 ( .A1(n4248), .A2(n6130), .ZN(n4639) );
  XNOR2_X1 U5346 ( .A(n5064), .B(n5063), .ZN(n8984) );
  OAI22_X1 U5347 ( .A1(n5090), .A2(n5059), .B1(SI_30_), .B2(n5088), .ZN(n5064)
         );
  NAND2_X1 U5348 ( .A1(n4914), .A2(n4912), .ZN(n5655) );
  OR2_X1 U5349 ( .A1(n5319), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5337) );
  AND2_X1 U5350 ( .A1(n5285), .A2(n5302), .ZN(n6993) );
  NOR2_X1 U5351 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n5154) );
  NOR2_X1 U5352 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n4744) );
  OAI211_X1 U5353 ( .C1(n4251), .C2(P1_DATAO_REG_2__SCAN_IN), .A(SI_2_), .B(
        n4441), .ZN(n4930) );
  NAND2_X1 U5354 ( .A1(n4251), .A2(n6740), .ZN(n4441) );
  XNOR2_X1 U5355 ( .A(n4933), .B(SI_3_), .ZN(n5162) );
  INV_X1 U5356 ( .A(P2_RD_REG_SCAN_IN), .ZN(n4797) );
  NOR2_X1 U5357 ( .A1(n9813), .A2(n9812), .ZN(n9814) );
  NAND2_X1 U5358 ( .A1(n9824), .A2(n9825), .ZN(n9826) );
  AND2_X1 U5359 ( .A1(n6409), .A2(n6408), .ZN(n8321) );
  AOI21_X1 U5360 ( .B1(n8353), .B2(n8352), .A(n8351), .ZN(n8367) );
  INV_X1 U5361 ( .A(n8760), .ZN(n8729) );
  NAND2_X1 U5362 ( .A1(n6303), .A2(n6302), .ZN(n8924) );
  OAI21_X1 U5363 ( .B1(n8354), .B2(n6473), .A(n6637), .ZN(n6474) );
  INV_X1 U5364 ( .A(n8321), .ZN(n8615) );
  AND4_X1 U5365 ( .A1(n6248), .A2(n6247), .A3(n6246), .A4(n6245), .ZN(n10039)
         );
  NAND2_X1 U5366 ( .A1(n6923), .A2(n6924), .ZN(n6922) );
  NAND2_X1 U5367 ( .A1(n6963), .A2(n6964), .ZN(n6962) );
  NAND2_X1 U5368 ( .A1(n7045), .A2(n7044), .ZN(n7043) );
  NAND2_X1 U5369 ( .A1(n7034), .A2(n7033), .ZN(n7145) );
  NAND2_X1 U5370 ( .A1(n7267), .A2(n7266), .ZN(n4514) );
  NAND2_X1 U5371 ( .A1(n10174), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n4816) );
  NAND2_X1 U5372 ( .A1(n10165), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n4819) );
  NOR2_X1 U5373 ( .A1(n8596), .A2(n8847), .ZN(n8260) );
  OR2_X1 U5374 ( .A1(n6105), .A2(n6104), .ZN(n6106) );
  NOR2_X1 U5375 ( .A1(n4703), .A2(n4417), .ZN(n4697) );
  OR2_X1 U5376 ( .A1(n4703), .A2(n6013), .ZN(n4699) );
  AND2_X1 U5377 ( .A1(n5474), .A2(n5473), .ZN(n9036) );
  NOR2_X1 U5378 ( .A1(n5986), .A2(n5983), .ZN(n5992) );
  OR2_X1 U5379 ( .A1(n5990), .A2(n9048), .ZN(n5991) );
  AND2_X1 U5380 ( .A1(n6053), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9137) );
  AND2_X1 U5381 ( .A1(n5462), .A2(n5461), .ZN(n9124) );
  AND4_X1 U5382 ( .A1(n5369), .A2(n5368), .A3(n5367), .A4(n5366), .ZN(n7907)
         );
  AND2_X1 U5383 ( .A1(n5487), .A2(n5486), .ZN(n9113) );
  OR2_X1 U5384 ( .A1(n7166), .A2(n9982), .ZN(n9145) );
  AND2_X1 U5385 ( .A1(n6049), .A2(n6035), .ZN(n9134) );
  INV_X1 U5386 ( .A(n9134), .ZN(n9132) );
  INV_X1 U5387 ( .A(n9140), .ZN(n9358) );
  INV_X1 U5388 ( .A(n9038), .ZN(n9402) );
  INV_X1 U5389 ( .A(n9113), .ZN(n9419) );
  INV_X1 U5390 ( .A(n9036), .ZN(n9440) );
  INV_X1 U5391 ( .A(n9124), .ZN(n9450) );
  XNOR2_X1 U5392 ( .A(n9182), .B(n4526), .ZN(n9203) );
  NOR2_X1 U5393 ( .A1(n9886), .A2(n9277), .ZN(n4525) );
  OR2_X1 U5394 ( .A1(P1_U3083), .A2(n7070), .ZN(n9877) );
  NAND2_X1 U5395 ( .A1(n5612), .A2(n5734), .ZN(n9508) );
  NOR2_X1 U5396 ( .A1(n4308), .A2(n9523), .ZN(n4381) );
  XNOR2_X1 U5397 ( .A(n9826), .B(P2_ADDR_REG_9__SCAN_IN), .ZN(n10215) );
  OAI21_X1 U5398 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10182), .ZN(n10211) );
  AOI21_X1 U5399 ( .B1(n6546), .B2(n6545), .A(n6544), .ZN(n6552) );
  AOI21_X1 U5400 ( .B1(n4573), .B2(n4575), .A(n4572), .ZN(n6577) );
  NOR2_X1 U5401 ( .A1(n4578), .A2(n4577), .ZN(n4572) );
  NAND2_X1 U5402 ( .A1(n6564), .A2(n6562), .ZN(n4575) );
  INV_X1 U5403 ( .A(n5275), .ZN(n4540) );
  NOR2_X1 U5404 ( .A1(n4538), .A2(n4537), .ZN(n4536) );
  NAND2_X1 U5405 ( .A1(n7854), .A2(n7850), .ZN(n4537) );
  INV_X1 U5406 ( .A(n5331), .ZN(n4538) );
  OAI211_X1 U5407 ( .C1(n6584), .C2(n6583), .A(n8710), .B(n6602), .ZN(n6585)
         );
  INV_X1 U5408 ( .A(n4551), .ZN(n4547) );
  AND2_X1 U5409 ( .A1(n5685), .A2(n4544), .ZN(n4543) );
  NAND2_X1 U5410 ( .A1(n4548), .A2(n4545), .ZN(n4544) );
  AND2_X1 U5411 ( .A1(n6604), .A2(n6606), .ZN(n4355) );
  NAND2_X1 U5412 ( .A1(n8707), .A2(n8730), .ZN(n4404) );
  NAND2_X1 U5413 ( .A1(n8759), .A2(n6582), .ZN(n6350) );
  OR2_X1 U5414 ( .A1(n10141), .A2(n7350), .ZN(n6545) );
  AND2_X1 U5415 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n6168) );
  NOR2_X1 U5416 ( .A1(n4428), .A2(n4255), .ZN(n4426) );
  NOR2_X1 U5417 ( .A1(n4691), .A2(n4687), .ZN(n4686) );
  INV_X1 U5418 ( .A(n7905), .ZN(n4691) );
  INV_X1 U5419 ( .A(n5897), .ZN(n4687) );
  NAND2_X1 U5420 ( .A1(n7905), .A2(n4690), .ZN(n4689) );
  INV_X1 U5421 ( .A(n5899), .ZN(n4690) );
  NAND2_X1 U5422 ( .A1(n4245), .A2(n7920), .ZN(n4661) );
  INV_X1 U5423 ( .A(n7569), .ZN(n4660) );
  NAND2_X1 U5424 ( .A1(n5186), .A2(n5185), .ZN(n7308) );
  INV_X1 U5425 ( .A(n9156), .ZN(n5185) );
  NAND2_X1 U5426 ( .A1(n9157), .A2(n9952), .ZN(n5702) );
  INV_X1 U5427 ( .A(n4615), .ZN(n4614) );
  NAND2_X1 U5428 ( .A1(n4617), .A2(n4612), .ZN(n4611) );
  INV_X1 U5429 ( .A(n5056), .ZN(n4612) );
  NOR2_X1 U5430 ( .A1(n4614), .A2(n5056), .ZN(n4613) );
  INV_X1 U5431 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n4908) );
  INV_X1 U5432 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n4870) );
  AND2_X1 U5433 ( .A1(n4624), .A2(n5515), .ZN(n4621) );
  NAND2_X1 U5434 ( .A1(n4989), .A2(n4988), .ZN(n4992) );
  INV_X1 U5435 ( .A(n5351), .ZN(n4983) );
  NAND2_X1 U5436 ( .A1(n5335), .A2(n4973), .ZN(n4367) );
  INV_X1 U5437 ( .A(n5332), .ZN(n4973) );
  INV_X1 U5438 ( .A(n4604), .ZN(n4603) );
  INV_X1 U5439 ( .A(n4945), .ZN(n4605) );
  INV_X1 U5440 ( .A(n4864), .ZN(n4863) );
  INV_X1 U5441 ( .A(n4953), .ZN(n4862) );
  AOI21_X1 U5442 ( .B1(n4735), .B2(n4733), .A(n4732), .ZN(n4731) );
  INV_X1 U5443 ( .A(n8296), .ZN(n4733) );
  INV_X1 U5444 ( .A(n8300), .ZN(n4732) );
  NOR2_X1 U5445 ( .A1(n8487), .A2(n4720), .ZN(n4719) );
  NOR2_X1 U5446 ( .A1(n6345), .A2(n6344), .ZN(n4361) );
  NOR2_X1 U5447 ( .A1(n6394), .A2(n6392), .ZN(n4360) );
  NOR2_X1 U5448 ( .A1(n8883), .A2(n4464), .ZN(n4463) );
  INV_X1 U5449 ( .A(n4465), .ZN(n4464) );
  NAND2_X1 U5450 ( .A1(n8883), .A2(n8658), .ZN(n4859) );
  NAND2_X1 U5451 ( .A1(n8687), .A2(n4859), .ZN(n4855) );
  INV_X1 U5452 ( .A(n4400), .ZN(n4398) );
  NOR2_X1 U5453 ( .A1(n8888), .A2(n8893), .ZN(n4465) );
  INV_X1 U5454 ( .A(n4361), .ZN(n6347) );
  NOR2_X1 U5455 ( .A1(n8909), .A2(n8915), .ZN(n4825) );
  AOI21_X1 U5456 ( .B1(n4486), .B2(n4484), .A(n8773), .ZN(n4483) );
  INV_X1 U5457 ( .A(n6574), .ZN(n4484) );
  NOR2_X1 U5458 ( .A1(n6270), .A2(n6269), .ZN(n6268) );
  INV_X1 U5459 ( .A(n10051), .ZN(n4470) );
  OR2_X1 U5460 ( .A1(n8941), .A2(n6278), .ZN(n6565) );
  NAND2_X1 U5461 ( .A1(n10065), .A2(n4392), .ZN(n4389) );
  NAND2_X1 U5462 ( .A1(n6545), .A2(n6547), .ZN(n7660) );
  INV_X1 U5463 ( .A(n10138), .ZN(n4810) );
  AND2_X1 U5464 ( .A1(n6168), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n6199) );
  OR2_X1 U5465 ( .A1(n10019), .A2(n7610), .ZN(n6519) );
  NOR2_X1 U5466 ( .A1(n6073), .A2(P2_IR_REG_28__SCAN_IN), .ZN(n6074) );
  OR2_X1 U5467 ( .A1(n6652), .A2(P2_IR_REG_27__SCAN_IN), .ZN(n4471) );
  NAND2_X1 U5468 ( .A1(n4823), .A2(n8624), .ZN(n4822) );
  NOR2_X1 U5469 ( .A1(n8665), .A2(n8873), .ZN(n8247) );
  AND2_X1 U5470 ( .A1(n4765), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n4492) );
  OAI21_X1 U5471 ( .B1(n4765), .B2(P2_IR_REG_29__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n4495) );
  NAND2_X1 U5472 ( .A1(n6084), .A2(n6085), .ZN(n4494) );
  AND2_X1 U5473 ( .A1(n4479), .A2(n4478), .ZN(n6065) );
  AND2_X1 U5474 ( .A1(n6064), .A2(n6094), .ZN(n6066) );
  INV_X1 U5475 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n6093) );
  INV_X1 U5476 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n6095) );
  OR2_X1 U5477 ( .A1(n6159), .A2(P2_IR_REG_3__SCAN_IN), .ZN(n6179) );
  NOR2_X1 U5478 ( .A1(n5480), .A2(n9035), .ZN(n4382) );
  INV_X1 U5479 ( .A(n5783), .ZN(n5787) );
  NAND2_X1 U5480 ( .A1(n7409), .A2(n5854), .ZN(n4434) );
  NAND2_X1 U5481 ( .A1(n4692), .A2(n4695), .ZN(n5974) );
  AOI21_X1 U5482 ( .B1(n9033), .B2(n5963), .A(n4303), .ZN(n4695) );
  AND3_X1 U5483 ( .A1(n5835), .A2(n4292), .A3(n7406), .ZN(n5838) );
  AND2_X1 U5484 ( .A1(n5612), .A2(n9266), .ZN(n5675) );
  INV_X1 U5485 ( .A(n4423), .ZN(n4422) );
  OAI21_X1 U5486 ( .B1(n4912), .B2(n9779), .A(n5065), .ZN(n4423) );
  NAND2_X1 U5487 ( .A1(n5109), .A2(n4555), .ZN(n4557) );
  NOR2_X1 U5488 ( .A1(n5083), .A2(n7209), .ZN(n4555) );
  NAND2_X1 U5489 ( .A1(n4535), .A2(n4534), .ZN(n4533) );
  NAND2_X1 U5490 ( .A1(n9856), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n4534) );
  INV_X1 U5491 ( .A(n9862), .ZN(n4535) );
  INV_X1 U5492 ( .A(n9261), .ZN(n4886) );
  AND2_X1 U5493 ( .A1(n9314), .A2(n9312), .ZN(n9264) );
  AND2_X1 U5494 ( .A1(n4460), .A2(n9257), .ZN(n4456) );
  NAND2_X1 U5495 ( .A1(n4460), .A2(n5542), .ZN(n4459) );
  NOR2_X1 U5496 ( .A1(n9541), .A2(n9546), .ZN(n4758) );
  NAND2_X1 U5497 ( .A1(n4382), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n5532) );
  OR2_X1 U5498 ( .A1(n9552), .A2(n9113), .ZN(n5680) );
  NAND2_X1 U5499 ( .A1(n5105), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n5467) );
  INV_X1 U5500 ( .A(n5455), .ZN(n5105) );
  NOR2_X1 U5501 ( .A1(n5421), .A2(n9730), .ZN(n4353) );
  INV_X1 U5502 ( .A(n9244), .ZN(n4876) );
  INV_X1 U5503 ( .A(n8110), .ZN(n4450) );
  INV_X1 U5504 ( .A(n4878), .ZN(n4877) );
  NAND2_X1 U5505 ( .A1(n9249), .A2(n9247), .ZN(n4880) );
  NOR2_X1 U5506 ( .A1(n5386), .A2(n8115), .ZN(n4383) );
  INV_X1 U5507 ( .A(n8007), .ZN(n4754) );
  NOR2_X1 U5508 ( .A1(n5291), .A2(n5290), .ZN(n5289) );
  NAND2_X1 U5509 ( .A1(n7718), .A2(n7717), .ZN(n4868) );
  OR2_X1 U5510 ( .A1(n7547), .A2(n7546), .ZN(n7548) );
  NOR2_X1 U5511 ( .A1(n7589), .A2(n4446), .ZN(n4445) );
  INV_X1 U5512 ( .A(n5240), .ZN(n4446) );
  AND2_X1 U5513 ( .A1(n9155), .A2(n9964), .ZN(n5621) );
  NAND2_X1 U5514 ( .A1(n9971), .A2(n5830), .ZN(n5622) );
  NAND2_X1 U5515 ( .A1(n7436), .A2(n4563), .ZN(n4560) );
  INV_X1 U5516 ( .A(n9514), .ZN(n9296) );
  NOR2_X1 U5517 ( .A1(n4869), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n4712) );
  INV_X1 U5518 ( .A(n5197), .ZN(n5070) );
  NAND2_X1 U5519 ( .A1(n4342), .A2(n4341), .ZN(n5665) );
  NOR2_X1 U5520 ( .A1(n5654), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n4341) );
  INV_X1 U5521 ( .A(n5655), .ZN(n4342) );
  INV_X1 U5522 ( .A(n5411), .ZN(n5002) );
  XNOR2_X1 U5523 ( .A(n5004), .B(SI_18_), .ZN(n5431) );
  NAND2_X1 U5524 ( .A1(n5000), .A2(SI_17_), .ZN(n5001) );
  XNOR2_X1 U5525 ( .A(n4999), .B(SI_17_), .ZN(n5411) );
  OAI21_X1 U5526 ( .B1(n4630), .B2(n5314), .A(n4628), .ZN(n4998) );
  AOI21_X1 U5527 ( .B1(n4629), .B2(n4634), .A(n4633), .ZN(n4628) );
  OR2_X1 U5528 ( .A1(n5358), .A2(n5357), .ZN(n5379) );
  XNOR2_X1 U5529 ( .A(n4984), .B(SI_14_), .ZN(n5351) );
  NAND2_X1 U5530 ( .A1(n4957), .A2(SI_10_), .ZN(n5280) );
  NAND2_X1 U5531 ( .A1(n4861), .A2(n4571), .ZN(n5277) );
  NAND2_X1 U5532 ( .A1(n4606), .A2(n4604), .ZN(n4571) );
  AND2_X1 U5533 ( .A1(n5278), .A2(n4956), .ZN(n5276) );
  OAI211_X1 U5534 ( .C1(n4830), .C2(n4831), .A(n4311), .B(n4365), .ZN(n5201)
         );
  NAND2_X1 U5535 ( .A1(n5172), .A2(n4829), .ZN(n4365) );
  AND2_X1 U5536 ( .A1(n4252), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n4928) );
  OAI21_X1 U5537 ( .B1(n4252), .B2(n9633), .A(n5150), .ZN(n4929) );
  OAI21_X1 U5538 ( .B1(n4251), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n4932), .ZN(
        n4933) );
  NAND2_X1 U5539 ( .A1(n6199), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n6210) );
  AND2_X1 U5540 ( .A1(n8373), .A2(n4736), .ZN(n4735) );
  NAND2_X1 U5541 ( .A1(n8443), .A2(n8296), .ZN(n4736) );
  NAND2_X1 U5542 ( .A1(n4357), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6336) );
  INV_X1 U5543 ( .A(n6326), .ZN(n4357) );
  NAND2_X1 U5544 ( .A1(n6079), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6345) );
  INV_X1 U5545 ( .A(n6336), .ZN(n6079) );
  OR2_X1 U5546 ( .A1(n6376), .A2(n9666), .ZN(n6394) );
  NAND2_X1 U5547 ( .A1(n10027), .A2(n6681), .ZN(n8435) );
  NAND2_X1 U5548 ( .A1(n6479), .A2(n10117), .ZN(n7698) );
  NAND2_X1 U5549 ( .A1(n4361), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6111) );
  NAND2_X1 U5551 ( .A1(n4359), .A2(n4358), .ZN(n6326) );
  NOR2_X1 U5552 ( .A1(n7629), .A2(n8500), .ZN(n4358) );
  INV_X1 U5553 ( .A(n6308), .ZN(n4359) );
  NAND2_X1 U5554 ( .A1(n4772), .A2(n4269), .ZN(n4590) );
  NOR2_X1 U5555 ( .A1(n8259), .A2(n8510), .ZN(n6632) );
  INV_X1 U5556 ( .A(n6493), .ZN(n4775) );
  INV_X1 U5557 ( .A(n6632), .ZN(n4774) );
  NAND2_X1 U5558 ( .A1(n6623), .A2(n4338), .ZN(n4777) );
  AND2_X1 U5559 ( .A1(n6629), .A2(n6628), .ZN(n6493) );
  NAND2_X1 U5560 ( .A1(n6436), .A2(n6625), .ZN(n4780) );
  NAND2_X1 U5561 ( .A1(n6166), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U5562 ( .A1(n4511), .A2(P2_IR_REG_1__SCAN_IN), .ZN(n4510) );
  INV_X1 U5563 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n4513) );
  OAI211_X1 U5564 ( .C1(n8527), .C2(P2_REG2_REG_1__SCAN_IN), .A(n8525), .B(
        n4506), .ZN(n8524) );
  NAND2_X1 U5565 ( .A1(n8527), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n4506) );
  NAND2_X1 U5566 ( .A1(n7934), .A2(n7935), .ZN(n4521) );
  INV_X1 U5567 ( .A(n4360), .ZN(n6402) );
  NAND2_X1 U5568 ( .A1(n4792), .A2(n4789), .ZN(n8645) );
  OAI21_X1 U5569 ( .B1(n8681), .B2(n4791), .A(n6606), .ZN(n4790) );
  NAND2_X2 U5570 ( .A1(n8645), .A2(n8646), .ZN(n8644) );
  NAND3_X1 U5571 ( .A1(n8722), .A2(n8877), .A3(n4463), .ZN(n8665) );
  NAND2_X1 U5572 ( .A1(n8722), .A2(n8707), .ZN(n8702) );
  NOR2_X1 U5573 ( .A1(n8898), .A2(n8751), .ZN(n8722) );
  NAND2_X1 U5574 ( .A1(n4852), .A2(n8237), .ZN(n4847) );
  INV_X1 U5575 ( .A(n4849), .ZN(n4848) );
  NAND2_X1 U5576 ( .A1(n8797), .A2(n4825), .ZN(n8762) );
  NAND2_X1 U5577 ( .A1(n8797), .A2(n8785), .ZN(n8787) );
  AND2_X1 U5578 ( .A1(n4802), .A2(n4474), .ZN(n8797) );
  NOR2_X1 U5579 ( .A1(n4476), .A2(n8919), .ZN(n4474) );
  NAND2_X1 U5580 ( .A1(n4802), .A2(n4801), .ZN(n8147) );
  NAND2_X1 U5581 ( .A1(n4802), .A2(n4475), .ZN(n8798) );
  NAND2_X1 U5582 ( .A1(n8048), .A2(n8052), .ZN(n8049) );
  AND4_X1 U5583 ( .A1(n6286), .A2(n6285), .A3(n6284), .A4(n6283), .ZN(n8499)
         );
  AND2_X1 U5584 ( .A1(n4467), .A2(n7803), .ZN(n8048) );
  NOR2_X1 U5585 ( .A1(n4469), .A2(n8941), .ZN(n4467) );
  NAND2_X1 U5586 ( .A1(n4468), .A2(n7803), .ZN(n7881) );
  INV_X1 U5587 ( .A(n4469), .ZN(n4468) );
  AOI21_X1 U5588 ( .B1(n4279), .B2(n4764), .A(n4761), .ZN(n4760) );
  INV_X1 U5589 ( .A(n6507), .ZN(n4764) );
  OAI21_X1 U5590 ( .B1(n4388), .B2(n4390), .A(n7824), .ZN(n7826) );
  OAI21_X1 U5591 ( .B1(n4392), .B2(n4391), .A(n7817), .ZN(n4390) );
  AND2_X1 U5592 ( .A1(n6243), .A2(n6078), .ZN(n6253) );
  NAND2_X1 U5593 ( .A1(n7803), .A2(n7808), .ZN(n7827) );
  AND2_X1 U5594 ( .A1(n6221), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6243) );
  NOR2_X1 U5595 ( .A1(n10069), .A2(n7761), .ZN(n7775) );
  NOR2_X1 U5596 ( .A1(n10141), .A2(n8434), .ZN(n4811) );
  INV_X1 U5597 ( .A(n7660), .ZN(n10087) );
  AND3_X1 U5598 ( .A1(n6118), .A2(n6119), .A3(n4498), .ZN(n6127) );
  INV_X1 U5599 ( .A(n4499), .ZN(n4498) );
  AND2_X1 U5600 ( .A1(n7689), .A2(n7688), .ZN(n4890) );
  NAND2_X1 U5601 ( .A1(n8636), .A2(n4821), .ZN(n8596) );
  NOR2_X1 U5602 ( .A1(n8852), .A2(n4822), .ZN(n4821) );
  AND2_X1 U5603 ( .A1(n10157), .A2(n10158), .ZN(n8949) );
  AND2_X1 U5604 ( .A1(n10101), .A2(n10109), .ZN(n6701) );
  AND2_X1 U5605 ( .A1(n7226), .A2(n7225), .ZN(n7247) );
  NAND2_X1 U5606 ( .A1(n6856), .A2(n10111), .ZN(n10102) );
  AND2_X1 U5607 ( .A1(n6073), .A2(n4766), .ZN(n4765) );
  OR2_X1 U5608 ( .A1(n6279), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n6319) );
  AND2_X1 U5609 ( .A1(n6184), .A2(n6204), .ZN(n6928) );
  NAND2_X1 U5610 ( .A1(n5188), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n5226) );
  NAND2_X1 U5611 ( .A1(n5102), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n5254) );
  INV_X1 U5612 ( .A(n5226), .ZN(n5102) );
  NAND2_X1 U5613 ( .A1(n4350), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n5386) );
  INV_X1 U5614 ( .A(n5364), .ZN(n4350) );
  AND2_X1 U5615 ( .A1(n6006), .A2(n6005), .ZN(n6044) );
  OR2_X1 U5616 ( .A1(n5467), .A2(n9101), .ZN(n5480) );
  INV_X1 U5617 ( .A(n4382), .ZN(n5493) );
  AND2_X1 U5618 ( .A1(n5987), .A2(n9047), .ZN(n5990) );
  AND2_X1 U5619 ( .A1(n5985), .A2(n5984), .ZN(n5986) );
  NAND2_X1 U5620 ( .A1(n4316), .A2(n9075), .ZN(n4708) );
  NAND2_X1 U5621 ( .A1(n4314), .A2(n5915), .ZN(n4706) );
  NAND2_X1 U5622 ( .A1(n4434), .A2(n5859), .ZN(n7643) );
  OR2_X1 U5623 ( .A1(n4434), .A2(n5859), .ZN(n7644) );
  NAND2_X1 U5624 ( .A1(n4432), .A2(n4300), .ZN(n7788) );
  NAND2_X1 U5625 ( .A1(n7409), .A2(n4429), .ZN(n4432) );
  NAND2_X1 U5626 ( .A1(n7646), .A2(n5860), .ZN(n4431) );
  NAND2_X1 U5627 ( .A1(n7065), .A2(n5798), .ZN(n5806) );
  NAND2_X1 U5628 ( .A1(n4706), .A2(n4255), .ZN(n9023) );
  NAND2_X1 U5629 ( .A1(n8121), .A2(n8124), .ZN(n5915) );
  OR2_X1 U5630 ( .A1(n5914), .A2(n5913), .ZN(n8122) );
  OR2_X1 U5631 ( .A1(n7053), .A2(n7054), .ZN(n7051) );
  NAND2_X1 U5632 ( .A1(n7131), .A2(n6819), .ZN(n9165) );
  OAI21_X1 U5633 ( .B1(n7103), .B2(n6828), .A(n6827), .ZN(n7002) );
  NOR2_X1 U5634 ( .A1(n7105), .A2(n7104), .ZN(n7103) );
  NAND2_X1 U5635 ( .A1(n7003), .A2(n7004), .ZN(n9186) );
  NAND2_X1 U5636 ( .A1(n9186), .A2(n4372), .ZN(n9837) );
  OR2_X1 U5637 ( .A1(n9187), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n4372) );
  NAND2_X1 U5638 ( .A1(n9177), .A2(n4523), .ZN(n9846) );
  OR2_X1 U5639 ( .A1(n9187), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n4523) );
  NOR2_X1 U5640 ( .A1(n9846), .A2(n9847), .ZN(n9845) );
  XNOR2_X1 U5641 ( .A(n4533), .B(n9191), .ZN(n9879) );
  NAND2_X1 U5642 ( .A1(n9872), .A2(n9871), .ZN(n9870) );
  XNOR2_X1 U5643 ( .A(n9179), .B(n4531), .ZN(n9890) );
  INV_X1 U5644 ( .A(n9885), .ZN(n4531) );
  OAI22_X1 U5645 ( .A1(n9879), .A2(n9178), .B1(n9874), .B2(n4532), .ZN(n9179)
         );
  INV_X1 U5646 ( .A(n4533), .ZN(n4532) );
  NAND2_X1 U5647 ( .A1(n9870), .A2(n4373), .ZN(n9193) );
  OR2_X1 U5648 ( .A1(n9191), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n4373) );
  NAND2_X1 U5649 ( .A1(n5092), .A2(n5091), .ZN(n9217) );
  AND2_X1 U5650 ( .A1(n5599), .A2(n5598), .ZN(n9288) );
  AND2_X1 U5651 ( .A1(n5590), .A2(n5562), .ZN(n9329) );
  INV_X1 U5652 ( .A(n9355), .ZN(n9342) );
  OR2_X1 U5653 ( .A1(n9346), .A2(n9484), .ZN(n4369) );
  AND2_X1 U5654 ( .A1(n4258), .A2(n9408), .ZN(n9363) );
  AND2_X1 U5655 ( .A1(n4461), .A2(n9258), .ZN(n9357) );
  NAND2_X1 U5656 ( .A1(n9358), .A2(n9449), .ZN(n4377) );
  NAND2_X1 U5657 ( .A1(n4643), .A2(n4642), .ZN(n9381) );
  AOI21_X1 U5658 ( .B1(n4644), .B2(n4646), .A(n4306), .ZN(n4642) );
  NAND2_X1 U5659 ( .A1(n9408), .A2(n4758), .ZN(n9377) );
  NAND2_X1 U5660 ( .A1(n9408), .A2(n9394), .ZN(n9390) );
  INV_X1 U5661 ( .A(n4665), .ZN(n4664) );
  INV_X1 U5662 ( .A(n4353), .ZN(n5439) );
  INV_X1 U5663 ( .A(n4383), .ZN(n5404) );
  NAND2_X1 U5664 ( .A1(n8136), .A2(n8110), .ZN(n9246) );
  NAND2_X1 U5665 ( .A1(n4256), .A2(n8104), .ZN(n4752) );
  INV_X1 U5666 ( .A(n7857), .ZN(n4884) );
  AOI21_X1 U5667 ( .B1(n7855), .B2(n4652), .A(n4310), .ZN(n4647) );
  NAND2_X1 U5668 ( .A1(n4754), .A2(n4755), .ZN(n8133) );
  NAND2_X1 U5669 ( .A1(n4351), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n5364) );
  INV_X1 U5670 ( .A(n5342), .ZN(n4351) );
  NOR2_X1 U5671 ( .A1(n8007), .A2(n9594), .ZN(n7896) );
  AND4_X1 U5672 ( .A1(n5296), .A2(n5295), .A3(n5294), .A4(n5293), .ZN(n7724)
         );
  AND2_X1 U5673 ( .A1(n7851), .A2(n5373), .ZN(n7850) );
  CLKBUF_X1 U5674 ( .A(n7710), .Z(n7927) );
  INV_X1 U5675 ( .A(n4749), .ZN(n4747) );
  INV_X1 U5676 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n5267) );
  OR2_X1 U5677 ( .A1(n5268), .A2(n5267), .ZN(n5291) );
  NAND2_X1 U5678 ( .A1(n7542), .A2(n7541), .ZN(n7544) );
  NAND2_X1 U5679 ( .A1(n4750), .A2(n7482), .ZN(n7562) );
  AND4_X1 U5680 ( .A1(n5260), .A2(n5259), .A3(n5258), .A4(n5257), .ZN(n7750)
         );
  NAND2_X1 U5681 ( .A1(n5629), .A2(n5628), .ZN(n7547) );
  NAND2_X1 U5682 ( .A1(n7479), .A2(n7480), .ZN(n7542) );
  AND2_X1 U5683 ( .A1(n7474), .A2(n7546), .ZN(n4559) );
  AND2_X1 U5684 ( .A1(n5628), .A2(n5626), .ZN(n7474) );
  OR2_X1 U5685 ( .A1(n9944), .A2(n7400), .ZN(n7396) );
  NOR2_X1 U5686 ( .A1(n9944), .A2(n4745), .ZN(n7429) );
  NAND2_X1 U5687 ( .A1(n9958), .A2(n9952), .ZN(n4745) );
  INV_X1 U5688 ( .A(n7314), .ZN(n7391) );
  NAND2_X1 U5689 ( .A1(n7193), .A2(n5618), .ZN(n4562) );
  INV_X1 U5690 ( .A(n9277), .ZN(n7285) );
  NAND2_X1 U5691 ( .A1(n9520), .A2(n9607), .ZN(n9521) );
  NAND2_X1 U5692 ( .A1(n5507), .A2(n5506), .ZN(n9533) );
  NAND2_X1 U5693 ( .A1(n5305), .A2(n5304), .ZN(n9606) );
  OR2_X1 U5694 ( .A1(n7329), .A2(n7198), .ZN(n9984) );
  INV_X1 U5695 ( .A(n9979), .ZN(n9611) );
  AND4_X1 U5696 ( .A1(n5068), .A2(n5069), .A3(n5070), .A4(n4710), .ZN(n5081)
         );
  AND2_X1 U5697 ( .A1(n4712), .A2(n4711), .ZN(n4710) );
  INV_X1 U5698 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4711) );
  XNOR2_X1 U5699 ( .A(n5099), .B(n5098), .ZN(n8992) );
  NAND2_X1 U5700 ( .A1(n5585), .A2(n5584), .ZN(n5050) );
  CLKBUF_X1 U5701 ( .A(n5660), .Z(n5661) );
  XNOR2_X1 U5702 ( .A(n5516), .B(n5515), .ZN(n7914) );
  NAND2_X1 U5703 ( .A1(n4618), .A2(n4624), .ZN(n5516) );
  NAND2_X1 U5704 ( .A1(n5021), .A2(n9634), .ZN(n5024) );
  XNOR2_X1 U5705 ( .A(n5609), .B(P1_IR_REG_21__SCAN_IN), .ZN(n7189) );
  NAND2_X1 U5706 ( .A1(n4607), .A2(n5016), .ZN(n5477) );
  NAND2_X1 U5707 ( .A1(n4594), .A2(n4597), .ZN(n5451) );
  AND2_X1 U5708 ( .A1(n5433), .A2(n5418), .ZN(n9184) );
  NAND2_X1 U5709 ( .A1(n4632), .A2(n4634), .ZN(n5397) );
  NAND2_X1 U5710 ( .A1(n5314), .A2(n4637), .ZN(n4632) );
  XNOR2_X1 U5711 ( .A(n5334), .B(n5333), .ZN(n7008) );
  XNOR2_X1 U5712 ( .A(n5314), .B(n5301), .ZN(n6777) );
  NAND2_X1 U5713 ( .A1(n4866), .A2(n4948), .ZN(n5248) );
  XNOR2_X1 U5714 ( .A(n5219), .B(n5218), .ZN(n6731) );
  NAND2_X1 U5715 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n4530) );
  INV_X1 U5716 ( .A(n5134), .ZN(n4803) );
  NOR2_X1 U5717 ( .A1(n9815), .A2(n10208), .ZN(n9816) );
  NAND2_X1 U5718 ( .A1(n7358), .A2(n4741), .ZN(n7458) );
  AND2_X1 U5719 ( .A1(n7358), .A2(n7357), .ZN(n7364) );
  AND4_X1 U5720 ( .A1(n6297), .A2(n6296), .A3(n6295), .A4(n6294), .ZN(n8068)
         );
  NAND2_X1 U5721 ( .A1(n7970), .A2(n7969), .ZN(n10011) );
  AND4_X1 U5722 ( .A1(n6259), .A2(n6258), .A3(n6257), .A4(n6256), .ZN(n10008)
         );
  NAND2_X1 U5723 ( .A1(n6125), .A2(n4497), .ZN(n6126) );
  AOI21_X1 U5724 ( .B1(n6410), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n4280), .ZN(
        n4497) );
  AND2_X1 U5725 ( .A1(n6092), .A2(n6091), .ZN(n8744) );
  NAND2_X1 U5726 ( .A1(n4730), .A2(n4735), .ZN(n8376) );
  NAND2_X1 U5727 ( .A1(n8444), .A2(n8296), .ZN(n4730) );
  OR2_X1 U5728 ( .A1(n8418), .A2(n8421), .ZN(n8312) );
  NAND2_X1 U5729 ( .A1(n4722), .A2(n4728), .ZN(n8476) );
  NAND2_X1 U5730 ( .A1(n4363), .A2(n8276), .ZN(n4722) );
  NAND2_X1 U5731 ( .A1(n4727), .A2(n8276), .ZN(n8410) );
  OR2_X1 U5732 ( .A1(n4363), .A2(n8271), .ZN(n4727) );
  INV_X1 U5733 ( .A(n10038), .ZN(n10029) );
  INV_X1 U5734 ( .A(n4741), .ZN(n4740) );
  OR2_X1 U5735 ( .A1(n8444), .A2(n8443), .ZN(n8445) );
  NAND2_X1 U5736 ( .A1(n7210), .A2(n6672), .ZN(n7178) );
  OR2_X1 U5737 ( .A1(n7174), .A2(n10159), .ZN(n8486) );
  INV_X1 U5738 ( .A(n4728), .ZN(n4726) );
  AOI21_X1 U5739 ( .B1(n4728), .B2(n4725), .A(n4724), .ZN(n4723) );
  NAND2_X1 U5740 ( .A1(n7299), .A2(n7298), .ZN(n7358) );
  NAND2_X1 U5741 ( .A1(n4721), .A2(n8390), .ZN(n8488) );
  OR2_X1 U5742 ( .A1(n8391), .A2(n8387), .ZN(n4721) );
  INV_X1 U5743 ( .A(n10055), .ZN(n8505) );
  INV_X1 U5744 ( .A(n8486), .ZN(n10052) );
  AOI21_X1 U5745 ( .B1(n8621), .B2(n6435), .A(n6416), .ZN(n8608) );
  INV_X1 U5746 ( .A(n6127), .ZN(n8522) );
  NAND2_X1 U5747 ( .A1(n6166), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n6152) );
  CLKBUF_X1 U5748 ( .A(n6146), .Z(n8523) );
  NAND2_X1 U5749 ( .A1(n6922), .A2(n4296), .ZN(n6937) );
  NAND2_X1 U5750 ( .A1(n6962), .A2(n4295), .ZN(n6912) );
  NAND2_X1 U5751 ( .A1(n7043), .A2(n4293), .ZN(n7034) );
  INV_X1 U5752 ( .A(n4522), .ZN(n7933) );
  AND2_X1 U5753 ( .A1(n8190), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n4520) );
  INV_X1 U5754 ( .A(n4519), .ZN(n8563) );
  INV_X1 U5755 ( .A(n4517), .ZN(n8191) );
  NAND2_X1 U5756 ( .A1(n6459), .A2(n6458), .ZN(n8844) );
  NAND2_X1 U5757 ( .A1(n6438), .A2(n6437), .ZN(n8847) );
  NAND2_X1 U5758 ( .A1(n4394), .A2(n4395), .ZN(n8245) );
  AOI21_X1 U5759 ( .B1(n4833), .B2(n4319), .A(n4309), .ZN(n4395) );
  INV_X1 U5760 ( .A(n8225), .ZN(n8226) );
  INV_X1 U5761 ( .A(n8601), .ZN(n8249) );
  NAND2_X1 U5762 ( .A1(n4834), .A2(n4835), .ZN(n8600) );
  OR2_X1 U5763 ( .A1(n8643), .A2(n4319), .ZN(n4834) );
  NAND2_X1 U5764 ( .A1(n4838), .A2(n4839), .ZN(n8617) );
  NAND2_X1 U5765 ( .A1(n8643), .A2(n4842), .ZN(n4838) );
  INV_X1 U5766 ( .A(n8861), .ZN(n8624) );
  INV_X1 U5767 ( .A(n4501), .ZN(n4500) );
  XNOR2_X1 U5768 ( .A(n4503), .B(n4772), .ZN(n4502) );
  AOI22_X1 U5769 ( .A1(n8616), .A2(n10060), .B1(n10058), .B2(n8615), .ZN(n4501) );
  AOI21_X1 U5770 ( .B1(n8643), .B2(n8242), .A(n4845), .ZN(n8629) );
  NAND2_X1 U5771 ( .A1(n4794), .A2(n4318), .ZN(n8656) );
  NAND2_X1 U5772 ( .A1(n4858), .A2(n4860), .ZN(n8680) );
  OR2_X1 U5773 ( .A1(n8688), .A2(n8694), .ZN(n4858) );
  INV_X1 U5774 ( .A(n4794), .ZN(n8673) );
  AND2_X1 U5775 ( .A1(n8697), .A2(n8696), .ZN(n8891) );
  AND3_X1 U5776 ( .A1(n4783), .A2(n4784), .A3(n4282), .ZN(n8695) );
  AND2_X1 U5777 ( .A1(n4402), .A2(n4405), .ZN(n8701) );
  NAND2_X1 U5778 ( .A1(n8721), .A2(n8727), .ZN(n4402) );
  NAND2_X1 U5779 ( .A1(n8778), .A2(n8237), .ZN(n8768) );
  NAND2_X1 U5780 ( .A1(n4482), .A2(n4486), .ZN(n8775) );
  AND2_X1 U5781 ( .A1(n4832), .A2(n8232), .ZN(n8808) );
  OAI21_X1 U5782 ( .B1(n6314), .B2(n4271), .A(n6574), .ZN(n8793) );
  NAND2_X1 U5783 ( .A1(n7799), .A2(n6507), .ZN(n7814) );
  OR2_X1 U5784 ( .A1(n8836), .A2(n7609), .ZN(n8803) );
  NAND2_X1 U5785 ( .A1(n10065), .A2(n7664), .ZN(n7764) );
  NAND2_X1 U5786 ( .A1(n10056), .A2(n6548), .ZN(n7669) );
  NOR2_X1 U5787 ( .A1(n8828), .A2(n8434), .ZN(n7736) );
  INV_X1 U5788 ( .A(n8803), .ZN(n10095) );
  OR2_X1 U5789 ( .A1(n10102), .A2(n7603), .ZN(n10090) );
  OR2_X1 U5790 ( .A1(n8908), .A2(n8907), .ZN(n8973) );
  INV_X1 U5791 ( .A(n10112), .ZN(n10108) );
  INV_X1 U5792 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n9750) );
  INV_X1 U5793 ( .A(n6709), .ZN(n7744) );
  INV_X1 U5794 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7172) );
  INV_X1 U5795 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7119) );
  INV_X1 U5796 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n7016) );
  INV_X1 U5797 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n7050) );
  INV_X1 U5798 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6836) );
  INV_X1 U5799 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n6758) );
  INV_X1 U5800 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6748) );
  INV_X1 U5801 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6727) );
  NAND2_X1 U5802 ( .A1(n4414), .A2(n4415), .ZN(n4409) );
  NAND2_X1 U5803 ( .A1(n6012), .A2(n4416), .ZN(n4415) );
  NOR3_X1 U5804 ( .A1(n4410), .A2(n4408), .A3(n6013), .ZN(n4407) );
  INV_X1 U5805 ( .A(n4414), .ZN(n4408) );
  AND4_X1 U5806 ( .A1(n5312), .A2(n5311), .A3(n5310), .A4(n5309), .ZN(n7999)
         );
  AND2_X1 U5807 ( .A1(n5445), .A2(n5444), .ZN(n9485) );
  NAND2_X1 U5808 ( .A1(n9032), .A2(n9033), .ZN(n9031) );
  NAND2_X1 U5809 ( .A1(n9098), .A2(n5964), .ZN(n9032) );
  AND2_X1 U5810 ( .A1(n5526), .A2(n5525), .ZN(n9053) );
  OR2_X1 U5811 ( .A1(n5568), .A2(n5208), .ZN(n5217) );
  NAND2_X1 U5812 ( .A1(n5564), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n5214) );
  AND2_X1 U5813 ( .A1(n5541), .A2(n5540), .ZN(n9090) );
  AOI21_X1 U5814 ( .B1(n8161), .B2(n4683), .A(n4274), .ZN(n4681) );
  NAND2_X1 U5815 ( .A1(n4680), .A2(n7644), .ZN(n7747) );
  NAND2_X1 U5816 ( .A1(n7643), .A2(n7646), .ZN(n4680) );
  NAND2_X1 U5817 ( .A1(n7904), .A2(n7905), .ZN(n7903) );
  NAND2_X1 U5818 ( .A1(n7948), .A2(n5899), .ZN(n7904) );
  AND4_X1 U5819 ( .A1(n5329), .A2(n5328), .A3(n5327), .A4(n5326), .ZN(n7893)
         );
  AND2_X1 U5820 ( .A1(n5835), .A2(n7406), .ZN(n7584) );
  AND2_X1 U5821 ( .A1(n6049), .A2(n6046), .ZN(n9016) );
  INV_X1 U5822 ( .A(n9016), .ZN(n9139) );
  AND2_X1 U5823 ( .A1(n6049), .A2(n6048), .ZN(n9142) );
  AND3_X1 U5824 ( .A1(n5408), .A2(n5407), .A3(n5406), .ZN(n9483) );
  INV_X1 U5825 ( .A(n9142), .ZN(n9037) );
  NAND2_X1 U5826 ( .A1(n5915), .A2(n8122), .ZN(n9058) );
  INV_X1 U5827 ( .A(n9145), .ZN(n9130) );
  NOR2_X1 U5828 ( .A1(n5769), .A2(n4568), .ZN(n4567) );
  NAND2_X1 U5829 ( .A1(n4566), .A2(n4565), .ZN(n4564) );
  NAND2_X1 U5830 ( .A1(n4570), .A2(n5603), .ZN(n4569) );
  NAND2_X1 U5831 ( .A1(n4438), .A2(n4436), .ZN(n7188) );
  NAND2_X1 U5832 ( .A1(n4439), .A2(n4437), .ZN(n4436) );
  NOR2_X1 U5833 ( .A1(n9740), .A2(P1_IR_REG_21__SCAN_IN), .ZN(n4435) );
  AND2_X1 U5834 ( .A1(n5115), .A2(n5114), .ZN(n9287) );
  INV_X1 U5835 ( .A(n9318), .ZN(n9271) );
  INV_X1 U5836 ( .A(n9053), .ZN(n9374) );
  INV_X1 U5837 ( .A(n9090), .ZN(n9387) );
  INV_X1 U5838 ( .A(n7907), .ZN(n9147) );
  INV_X1 U5839 ( .A(n7999), .ZN(n9150) );
  INV_X1 U5840 ( .A(n7589), .ZN(n9154) );
  NAND2_X1 U5841 ( .A1(n6989), .A2(n7064), .ZN(n6988) );
  INV_X1 U5842 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n9808) );
  NAND2_X1 U5843 ( .A1(n7135), .A2(n4253), .ZN(n9168) );
  AND2_X1 U5844 ( .A1(n7135), .A2(n6810), .ZN(n9169) );
  NOR2_X1 U5845 ( .A1(n6992), .A2(n4334), .ZN(n6994) );
  NAND2_X1 U5846 ( .A1(n6994), .A2(n6995), .ZN(n9177) );
  AND2_X1 U5847 ( .A1(n6783), .A2(n6771), .ZN(n9911) );
  NAND2_X1 U5848 ( .A1(n5077), .A2(n6663), .ZN(n9496) );
  OAI21_X1 U5849 ( .B1(n9241), .B2(n4676), .A(n4674), .ZN(n4677) );
  INV_X1 U5850 ( .A(n4675), .ZN(n4674) );
  OAI21_X1 U5851 ( .B1(n4278), .B2(n4676), .A(n9285), .ZN(n4675) );
  INV_X1 U5852 ( .A(n4454), .ZN(n4453) );
  OAI21_X1 U5853 ( .B1(n9318), .B2(n9484), .A(n9316), .ZN(n4454) );
  INV_X1 U5854 ( .A(n9209), .ZN(n9328) );
  INV_X1 U5855 ( .A(n9263), .ZN(n9332) );
  AOI21_X1 U5856 ( .B1(n9326), .B2(n9454), .A(n9325), .ZN(n9529) );
  NAND2_X1 U5857 ( .A1(n9324), .A2(n9323), .ZN(n9325) );
  NAND2_X1 U5858 ( .A1(n4893), .A2(n9311), .ZN(n9326) );
  AOI21_X1 U5859 ( .B1(n4378), .B2(n9454), .A(n4375), .ZN(n9539) );
  NAND2_X1 U5860 ( .A1(n4377), .A2(n4376), .ZN(n4375) );
  NAND2_X1 U5861 ( .A1(n9355), .A2(n4287), .ZN(n4378) );
  NAND2_X1 U5862 ( .A1(n9387), .A2(n9451), .ZN(n4376) );
  NAND2_X1 U5863 ( .A1(n9404), .A2(n9232), .ZN(n9395) );
  INV_X1 U5864 ( .A(n9552), .ZN(n9414) );
  AND2_X1 U5865 ( .A1(n4871), .A2(n9253), .ZN(n9401) );
  NAND2_X1 U5866 ( .A1(n9437), .A2(n9251), .ZN(n9418) );
  NAND2_X1 U5867 ( .A1(n4666), .A2(n4667), .ZN(n9432) );
  OR2_X1 U5868 ( .A1(n4672), .A2(n4669), .ZN(n4666) );
  NAND2_X1 U5869 ( .A1(n4670), .A2(n9226), .ZN(n9466) );
  NAND2_X1 U5870 ( .A1(n4670), .A2(n4668), .ZN(n9567) );
  AND2_X1 U5871 ( .A1(n9487), .A2(n9247), .ZN(n9448) );
  NAND2_X1 U5872 ( .A1(n7892), .A2(n7857), .ZN(n8109) );
  NAND2_X1 U5873 ( .A1(n4654), .A2(n7844), .ZN(n8098) );
  NAND2_X1 U5874 ( .A1(n7888), .A2(n7890), .ZN(n4654) );
  NAND2_X1 U5875 ( .A1(n7570), .A2(n7569), .ZN(n7706) );
  AND2_X1 U5876 ( .A1(n9463), .A2(n7333), .ZN(n9365) );
  INV_X1 U5877 ( .A(n9365), .ZN(n9475) );
  AND2_X1 U5878 ( .A1(n9512), .A2(n9506), .ZN(n4368) );
  AND2_X2 U5879 ( .A1(n7284), .A2(n7206), .ZN(n9991) );
  AND2_X1 U5880 ( .A1(n9777), .A2(n9776), .ZN(n9942) );
  INV_X1 U5881 ( .A(n7188), .ZN(n5784) );
  INV_X1 U5882 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n9755) );
  XNOR2_X1 U5883 ( .A(n5652), .B(n5065), .ZN(n7642) );
  INV_X1 U5884 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n7171) );
  INV_X1 U5885 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7018) );
  AND2_X1 U5886 ( .A1(n5337), .A2(n5320), .ZN(n9839) );
  INV_X1 U5887 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6757) );
  INV_X1 U5888 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n6750) );
  AND2_X1 U5889 ( .A1(n5239), .A2(n5249), .ZN(n9163) );
  NAND2_X1 U5890 ( .A1(n5154), .A2(n4744), .ZN(n5174) );
  NAND2_X1 U5891 ( .A1(n4440), .A2(SI_0_), .ZN(n5143) );
  INV_X1 U5892 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10181) );
  OAI21_X1 U5893 ( .B1(n10177), .B2(n10181), .A(n10179), .ZN(n10219) );
  NAND2_X1 U5894 ( .A1(n4343), .A2(n9811), .ZN(n10223) );
  NAND2_X1 U5895 ( .A1(n10221), .A2(n10222), .ZN(n4343) );
  AND2_X1 U5896 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9814), .ZN(n10207) );
  XNOR2_X1 U5897 ( .A(n9816), .B(n4347), .ZN(n10206) );
  INV_X1 U5898 ( .A(P1_ADDR_REG_6__SCAN_IN), .ZN(n4347) );
  XOR2_X1 U5899 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n9819), .Z(n10218) );
  NOR2_X1 U5900 ( .A1(n10214), .A2(n9827), .ZN(n10205) );
  NOR2_X1 U5901 ( .A1(n10205), .A2(n10204), .ZN(n10203) );
  AOI21_X1 U5902 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n10203), .ZN(n10202) );
  AOI21_X1 U5903 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10200), .ZN(n10199) );
  OAI21_X1 U5904 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10197), .ZN(n10195) );
  OAI21_X1 U5905 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10194), .ZN(n10192) );
  NAND2_X1 U5906 ( .A1(n10191), .A2(n4344), .ZN(n10189) );
  NAND2_X1 U5907 ( .A1(n4346), .A2(n4345), .ZN(n4344) );
  NAND2_X1 U5908 ( .A1(n10189), .A2(n10190), .ZN(n10188) );
  OR2_X1 U5909 ( .A1(n6635), .A2(n4263), .ZN(n4387) );
  INV_X1 U5910 ( .A(n4515), .ZN(n7265) );
  INV_X1 U5911 ( .A(n4815), .ZN(n4814) );
  OAI21_X1 U5912 ( .B1(n4272), .B2(n10174), .A(n4816), .ZN(n4815) );
  INV_X1 U5913 ( .A(n4818), .ZN(n4817) );
  OAI21_X1 U5914 ( .B1(n4272), .B2(n10165), .A(n4819), .ZN(n4818) );
  NAND2_X1 U5915 ( .A1(n4684), .A2(n5815), .ZN(n8160) );
  AND2_X1 U5916 ( .A1(n4320), .A2(n4699), .ZN(n4698) );
  NAND2_X1 U5917 ( .A1(n9204), .A2(n9277), .ZN(n4527) );
  NAND2_X1 U5918 ( .A1(n9618), .A2(n9991), .ZN(n4452) );
  INV_X1 U5919 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n4451) );
  OAI21_X1 U5920 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(n9831), .A(n10210), .ZN(
        n9833) );
  BUF_X1 U5921 ( .A(n5135), .Z(n6663) );
  INV_X1 U5922 ( .A(n4356), .ZN(n4672) );
  AND2_X1 U5923 ( .A1(n9170), .A2(n6810), .ZN(n4253) );
  NAND2_X1 U5924 ( .A1(n5130), .A2(n4267), .ZN(n5694) );
  AND2_X1 U5925 ( .A1(n8722), .A2(n4463), .ZN(n4254) );
  AND2_X1 U5926 ( .A1(n4708), .A2(n5938), .ZN(n4255) );
  INV_X1 U5927 ( .A(n9958), .ZN(n5186) );
  AND2_X1 U5928 ( .A1(n4755), .A2(n4753), .ZN(n4256) );
  AND2_X1 U5929 ( .A1(n9258), .A2(n9356), .ZN(n4460) );
  AND2_X1 U5930 ( .A1(n9568), .A2(n9441), .ZN(n4257) );
  INV_X1 U5931 ( .A(n9251), .ZN(n4873) );
  AND2_X1 U5932 ( .A1(n4758), .A2(n4757), .ZN(n4258) );
  AND2_X1 U5933 ( .A1(n6011), .A2(n6010), .ZN(n4259) );
  AND2_X1 U5934 ( .A1(n4307), .A2(n8026), .ZN(n4260) );
  NAND2_X1 U5935 ( .A1(n4554), .A2(n5608), .ZN(n4261) );
  NOR2_X1 U5936 ( .A1(n4778), .A2(n4776), .ZN(n4262) );
  NAND2_X1 U5937 ( .A1(n4754), .A2(n4256), .ZN(n4756) );
  INV_X1 U5938 ( .A(n8924), .ZN(n4477) );
  NAND2_X1 U5939 ( .A1(n7533), .A2(n9971), .ZN(n7481) );
  NAND4_X1 U5940 ( .A1(n7508), .A2(n6637), .A3(n7235), .A4(n6702), .ZN(n4263)
         );
  NAND2_X2 U5941 ( .A1(n6491), .A2(n7744), .ZN(n6630) );
  INV_X1 U5942 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n9740) );
  INV_X1 U5943 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U5944 ( .A1(n8027), .A2(n8026), .ZN(n8233) );
  INV_X1 U5945 ( .A(n8711), .ZN(n4787) );
  INV_X1 U5946 ( .A(n9136), .ZN(n4417) );
  NAND2_X1 U5947 ( .A1(n9556), .A2(n9440), .ZN(n4264) );
  NOR2_X1 U5948 ( .A1(n9050), .A2(n4418), .ZN(n4265) );
  NAND2_X1 U5949 ( .A1(n8176), .A2(n8175), .ZN(n4266) );
  AND2_X2 U5950 ( .A1(n6132), .A2(n4896), .ZN(n7689) );
  AND3_X1 U5951 ( .A1(n4558), .A2(n4557), .A3(n4556), .ZN(n4267) );
  AND2_X1 U5952 ( .A1(n5718), .A2(n8110), .ZN(n4268) );
  OR2_X1 U5953 ( .A1(n6615), .A2(n6630), .ZN(n4269) );
  OR2_X1 U5954 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n4270) );
  NAND2_X1 U5955 ( .A1(n6313), .A2(n6573), .ZN(n4271) );
  NAND2_X1 U5956 ( .A1(n6350), .A2(n6595), .ZN(n8708) );
  AND2_X1 U5957 ( .A1(n8845), .A2(n8849), .ZN(n4272) );
  AND2_X1 U5958 ( .A1(n4885), .A2(n9264), .ZN(n4273) );
  NOR2_X1 U5959 ( .A1(n5819), .A2(n5818), .ZN(n4274) );
  INV_X1 U5960 ( .A(n6623), .ZN(n4779) );
  OR2_X1 U5961 ( .A1(n6148), .A2(n7699), .ZN(n4276) );
  OR2_X1 U5962 ( .A1(n9556), .A2(n9036), .ZN(n9253) );
  OR2_X1 U5963 ( .A1(n6579), .A2(n6630), .ZN(n4277) );
  AND2_X1 U5964 ( .A1(n4679), .A2(n9240), .ZN(n4278) );
  AND2_X1 U5965 ( .A1(n6260), .A2(n4762), .ZN(n4279) );
  NAND2_X1 U5966 ( .A1(n5492), .A2(n5491), .ZN(n9546) );
  NOR2_X1 U5967 ( .A1(n6588), .A2(n6496), .ZN(n8694) );
  NAND2_X1 U5968 ( .A1(n6352), .A2(n6351), .ZN(n8893) );
  NAND2_X1 U5969 ( .A1(n6108), .A2(n6107), .ZN(n8755) );
  INV_X1 U5970 ( .A(n8755), .ZN(n4824) );
  INV_X1 U5971 ( .A(n8390), .ZN(n4720) );
  NAND2_X1 U5972 ( .A1(n6145), .A2(n10117), .ZN(n6477) );
  NAND2_X1 U5973 ( .A1(n6617), .A2(n6618), .ZN(n8618) );
  AND2_X1 U5974 ( .A1(n6861), .A2(n6942), .ZN(n4280) );
  AND2_X1 U5975 ( .A1(n8232), .A2(n8807), .ZN(n4281) );
  NAND2_X1 U5976 ( .A1(n8893), .A2(n8730), .ZN(n4282) );
  OR2_X1 U5977 ( .A1(n9541), .A2(n9090), .ZN(n9258) );
  XNOR2_X1 U5978 ( .A(n4947), .B(SI_7_), .ZN(n5233) );
  INV_X1 U5979 ( .A(n6591), .ZN(n4793) );
  AND2_X1 U5980 ( .A1(n8319), .A2(n8318), .ZN(n4283) );
  INV_X1 U5981 ( .A(n7920), .ZN(n9152) );
  AND4_X1 U5982 ( .A1(n5273), .A2(n5272), .A3(n5271), .A4(n5270), .ZN(n7920)
         );
  AND2_X1 U5983 ( .A1(n6493), .A2(n4262), .ZN(n4285) );
  NAND2_X1 U5984 ( .A1(n8630), .A2(n6494), .ZN(n8242) );
  INV_X1 U5985 ( .A(n8242), .ZN(n8646) );
  AND2_X1 U5986 ( .A1(n8893), .A2(n8513), .ZN(n4286) );
  INV_X1 U5987 ( .A(n4840), .ZN(n4839) );
  OAI21_X1 U5988 ( .B1(n8632), .B2(n4841), .A(n4844), .ZN(n4840) );
  INV_X1 U5989 ( .A(n6130), .ZN(n8156) );
  XNOR2_X1 U5990 ( .A(n4804), .B(n4803), .ZN(n6130) );
  NAND2_X1 U5991 ( .A1(n4975), .A2(n4971), .ZN(n5332) );
  OR2_X1 U5992 ( .A1(n9357), .A2(n9356), .ZN(n4287) );
  NAND2_X1 U5993 ( .A1(n5655), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5652) );
  AND2_X1 U5994 ( .A1(n4541), .A2(n4547), .ZN(n4288) );
  AND2_X1 U5995 ( .A1(n4824), .A2(n4825), .ZN(n4289) );
  INV_X1 U5996 ( .A(n9227), .ZN(n4671) );
  OR2_X1 U5997 ( .A1(n9561), .A2(n9450), .ZN(n4290) );
  AND2_X1 U5998 ( .A1(n4783), .A2(n4784), .ZN(n4291) );
  INV_X1 U5999 ( .A(n8237), .ZN(n4850) );
  NAND2_X1 U6000 ( .A1(n6429), .A2(n6428), .ZN(n8852) );
  NAND2_X1 U6001 ( .A1(n7511), .A2(n7516), .ZN(n4292) );
  OR2_X1 U6002 ( .A1(n7040), .A2(n7032), .ZN(n4293) );
  OR2_X1 U6003 ( .A1(n6910), .A2(n10092), .ZN(n4294) );
  OR2_X1 U6004 ( .A1(n6967), .A2(n6911), .ZN(n4295) );
  OR2_X1 U6005 ( .A1(n6927), .A2(n7612), .ZN(n4296) );
  OR2_X1 U6006 ( .A1(n7030), .A2(n7029), .ZN(n4297) );
  OR2_X1 U6007 ( .A1(n7555), .A2(n7554), .ZN(n4298) );
  AND2_X1 U6008 ( .A1(n4597), .A2(n4593), .ZN(n4299) );
  AND2_X1 U6009 ( .A1(n5870), .A2(n4431), .ZN(n4300) );
  NAND2_X1 U6010 ( .A1(n6266), .A2(n6265), .ZN(n8941) );
  OR2_X1 U6011 ( .A1(n7709), .A2(n7724), .ZN(n7848) );
  AND2_X1 U6012 ( .A1(n4878), .A2(n4876), .ZN(n4301) );
  NAND2_X1 U6013 ( .A1(n5402), .A2(n5401), .ZN(n9580) );
  NOR2_X1 U6014 ( .A1(n9163), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n4302) );
  NOR2_X1 U6015 ( .A1(n5969), .A2(n5968), .ZN(n4303) );
  NAND2_X1 U6016 ( .A1(n8236), .A2(n8235), .ZN(n8778) );
  OR2_X1 U6017 ( .A1(n8919), .A2(n8501), .ZN(n6497) );
  NAND2_X1 U6018 ( .A1(n5953), .A2(n9094), .ZN(n4304) );
  AND2_X1 U6019 ( .A1(n4858), .A2(n4856), .ZN(n4305) );
  AND2_X1 U6020 ( .A1(n9546), .A2(n9402), .ZN(n4306) );
  INV_X1 U6021 ( .A(n5218), .ZN(n4943) );
  XNOR2_X1 U6022 ( .A(n4944), .B(SI_6_), .ZN(n5218) );
  INV_X1 U6023 ( .A(n8856), .ZN(n4823) );
  INV_X1 U6024 ( .A(n4476), .ZN(n4475) );
  NAND2_X1 U6025 ( .A1(n4801), .A2(n4477), .ZN(n4476) );
  AND2_X1 U6026 ( .A1(n9556), .A2(n9036), .ZN(n9252) );
  AND2_X1 U6027 ( .A1(n6498), .A2(n6500), .ZN(n8781) );
  INV_X1 U6028 ( .A(n8781), .ZN(n8235) );
  AND2_X1 U6029 ( .A1(n8231), .A2(n8228), .ZN(n4307) );
  NAND2_X1 U6030 ( .A1(n9522), .A2(n9521), .ZN(n4308) );
  INV_X1 U6031 ( .A(n4577), .ZN(n4576) );
  NAND2_X1 U6032 ( .A1(n6384), .A2(n6383), .ZN(n8667) );
  NOR2_X1 U6033 ( .A1(n8856), .A2(n8616), .ZN(n4309) );
  NOR2_X1 U6034 ( .A1(n9590), .A2(n9147), .ZN(n4310) );
  INV_X1 U6035 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n5653) );
  NAND2_X1 U6036 ( .A1(n4938), .A2(SI_4_), .ZN(n4311) );
  OR2_X1 U6037 ( .A1(n8667), .A2(n8678), .ZN(n6606) );
  NAND2_X1 U6038 ( .A1(n4706), .A2(n4708), .ZN(n4312) );
  OR2_X1 U6039 ( .A1(n5300), .A2(n5299), .ZN(n4313) );
  INV_X1 U6040 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7116) );
  AND2_X1 U6041 ( .A1(n8122), .A2(n4707), .ZN(n4314) );
  NAND2_X1 U6042 ( .A1(n5276), .A2(n5280), .ZN(n4315) );
  AND2_X1 U6043 ( .A1(n5030), .A2(n5029), .ZN(n5527) );
  NAND2_X1 U6044 ( .A1(n5929), .A2(n9074), .ZN(n4316) );
  INV_X1 U6045 ( .A(n9366), .ZN(n4757) );
  OR2_X1 U6046 ( .A1(n4403), .A2(n4286), .ZN(n4317) );
  AND2_X1 U6047 ( .A1(n8657), .A2(n4793), .ZN(n4318) );
  OR2_X1 U6048 ( .A1(n4840), .A2(n4837), .ZN(n4319) );
  AND2_X1 U6049 ( .A1(n6062), .A2(n6061), .ZN(n4320) );
  AND3_X1 U6050 ( .A1(n6627), .A2(n4779), .A3(n6628), .ZN(n4321) );
  AND2_X1 U6051 ( .A1(n4861), .A2(n4943), .ZN(n4322) );
  AND2_X1 U6052 ( .A1(n9546), .A2(n9038), .ZN(n9256) );
  INV_X1 U6053 ( .A(n9256), .ZN(n4462) );
  AND2_X1 U6054 ( .A1(n6620), .A2(n6621), .ZN(n8243) );
  INV_X1 U6055 ( .A(n8243), .ZN(n8605) );
  AND2_X1 U6056 ( .A1(n9266), .A2(n5731), .ZN(n9285) );
  AND2_X1 U6057 ( .A1(n8243), .A2(n6619), .ZN(n4323) );
  AND2_X1 U6058 ( .A1(n8042), .A2(n6567), .ZN(n4324) );
  AND2_X1 U6059 ( .A1(n9254), .A2(n9253), .ZN(n4325) );
  AND2_X1 U6060 ( .A1(n4427), .A2(n4707), .ZN(n4326) );
  AND2_X1 U6061 ( .A1(n9311), .A2(n9312), .ZN(n4327) );
  OR2_X1 U6062 ( .A1(n9546), .A2(n9038), .ZN(n9257) );
  AND2_X1 U6063 ( .A1(n4765), .A2(n6085), .ZN(n4328) );
  AND2_X1 U6064 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(n9779), .ZN(n4329) );
  INV_X1 U6065 ( .A(n4659), .ZN(n4658) );
  NOR2_X1 U6066 ( .A1(n7705), .A2(n4660), .ZN(n4659) );
  AND2_X1 U6067 ( .A1(n4369), .A2(n9345), .ZN(n4330) );
  NAND2_X1 U6068 ( .A1(n8722), .A2(n4465), .ZN(n4466) );
  INV_X1 U6069 ( .A(n6322), .ZN(n6161) );
  INV_X1 U6070 ( .A(n8661), .ZN(n4846) );
  NAND2_X1 U6071 ( .A1(n4389), .A2(n7762), .ZN(n7818) );
  NAND2_X1 U6072 ( .A1(n6236), .A2(n6553), .ZN(n7799) );
  NAND2_X1 U6073 ( .A1(n7851), .A2(n7852), .ZN(n7998) );
  NAND2_X1 U6074 ( .A1(n5784), .A2(n7285), .ZN(n7096) );
  INV_X1 U6075 ( .A(n8883), .ZN(n4800) );
  AND2_X1 U6076 ( .A1(n7775), .A2(n7778), .ZN(n7803) );
  AND2_X1 U6077 ( .A1(n9421), .A2(n9426), .ZN(n9407) );
  AND2_X1 U6078 ( .A1(n9208), .A2(n9476), .ZN(n9455) );
  OAI21_X1 U6079 ( .B1(n7852), .B2(n4444), .A(n4442), .ZN(n7889) );
  AND2_X1 U6080 ( .A1(n5476), .A2(n5016), .ZN(n4331) );
  AND2_X1 U6081 ( .A1(n7323), .A2(n7546), .ZN(n4332) );
  INV_X1 U6082 ( .A(n9520), .ZN(n4371) );
  OR2_X1 U6083 ( .A1(n7481), .A2(n4747), .ZN(n4751) );
  OR2_X1 U6084 ( .A1(n7369), .A2(n7368), .ZN(n4333) );
  AND2_X1 U6085 ( .A1(n6993), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n4334) );
  INV_X1 U6086 ( .A(n7481), .ZN(n4750) );
  AND2_X1 U6087 ( .A1(n5052), .A2(n5051), .ZN(n4335) );
  AND2_X1 U6088 ( .A1(n5032), .A2(SI_24_), .ZN(n4336) );
  OR2_X1 U6089 ( .A1(n10174), .A2(n10149), .ZN(n4337) );
  INV_X1 U6090 ( .A(n4669), .ZN(n4668) );
  NAND2_X1 U6091 ( .A1(n9248), .A2(n9226), .ZN(n4669) );
  INV_X1 U6092 ( .A(n4405), .ZN(n4403) );
  NAND2_X1 U6093 ( .A1(n8898), .A2(n8714), .ZN(n4405) );
  INV_X1 U6094 ( .A(n7610), .ZN(n8434) );
  AND2_X2 U6095 ( .A1(n7247), .A2(n7227), .ZN(n10166) );
  OR2_X1 U6096 ( .A1(n8510), .A2(n7621), .ZN(n4338) );
  NAND2_X1 U6097 ( .A1(n4812), .A2(n4809), .ZN(n7735) );
  INV_X1 U6098 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n4766) );
  NAND2_X1 U6099 ( .A1(n5382), .A2(n5381), .ZN(n9583) );
  INV_X1 U6100 ( .A(n9583), .ZN(n4753) );
  INV_X1 U6101 ( .A(n8929), .ZN(n4801) );
  NAND2_X1 U6102 ( .A1(n6082), .A2(n6073), .ZN(n6653) );
  OR2_X1 U6103 ( .A1(n10165), .A2(n10149), .ZN(n4339) );
  OR2_X1 U6104 ( .A1(n9991), .A2(n4451), .ZN(n4340) );
  INV_X1 U6105 ( .A(n8202), .ZN(n4516) );
  INV_X1 U6106 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n4346) );
  INV_X1 U6107 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n4526) );
  INV_X1 U6108 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n4380) );
  INV_X1 U6109 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n4345) );
  INV_X1 U6110 ( .A(n8958), .ZN(n10159) );
  MUX2_X1 U6111 ( .A(n6493), .B(n6492), .S(n6630), .Z(n6634) );
  MUX2_X1 U6112 ( .A(n6587), .B(n6586), .S(n6630), .Z(n6590) );
  MUX2_X1 U6113 ( .A(n6520), .B(n6539), .S(n6630), .Z(n6542) );
  OR2_X2 U6114 ( .A1(n10138), .A2(n8521), .ZN(n6529) );
  AOI21_X1 U6115 ( .B1(n6542), .B2(n6531), .A(n6530), .ZN(n6532) );
  NAND2_X1 U6116 ( .A1(n6099), .A2(n6216), .ZN(n6331) );
  NAND3_X1 U6117 ( .A1(n8313), .A2(n8314), .A3(n8312), .ZN(n8391) );
  NAND2_X1 U6118 ( .A1(n8269), .A2(n8268), .ZN(n8399) );
  OAI21_X1 U6119 ( .B1(n9049), .B2(n9050), .A(n9134), .ZN(n9056) );
  NOR2_X1 U6120 ( .A1(n5974), .A2(n5973), .ZN(n9106) );
  NAND2_X1 U6121 ( .A1(n9447), .A2(n9250), .ZN(n9438) );
  NAND2_X1 U6122 ( .A1(n4882), .A2(n4881), .ZN(n8137) );
  AOI21_X2 U6123 ( .B1(n9386), .B2(n9257), .A(n9256), .ZN(n9373) );
  NAND3_X1 U6124 ( .A1(n5070), .A2(n5069), .A3(n5068), .ZN(n5660) );
  NOR2_X2 U6125 ( .A1(n4911), .A2(n4910), .ZN(n5068) );
  NAND2_X1 U6126 ( .A1(n4370), .A2(n4330), .ZN(n9531) );
  NAND2_X1 U6127 ( .A1(n4871), .A2(n4325), .ZN(n9400) );
  NAND2_X2 U6128 ( .A1(n4461), .A2(n4460), .ZN(n9355) );
  NOR2_X1 U6129 ( .A1(n10202), .A2(n10201), .ZN(n10200) );
  NOR4_X2 U6130 ( .A1(n8605), .A2(n8618), .A3(n8628), .A4(n6488), .ZN(n6489)
         );
  NOR4_X1 U6131 ( .A1(n8687), .A2(n8711), .A3(n8727), .A4(n6486), .ZN(n6487)
         );
  OAI211_X2 U6132 ( .C1(n4275), .C2(n8657), .A(n8656), .B(n10080), .ZN(n8660)
         );
  AOI211_X2 U6133 ( .C1(n8880), .C2(n10155), .A(n8879), .B(n8878), .ZN(n8881)
         );
  OAI21_X2 U6134 ( .B1(n9355), .B2(n4887), .A(n4273), .ZN(n9313) );
  NAND2_X1 U6135 ( .A1(n4384), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n5561) );
  XNOR2_X1 U6136 ( .A(n5153), .B(n5152), .ZN(n6741) );
  AND2_X2 U6137 ( .A1(n8041), .A2(n4352), .ZN(n6314) );
  NOR2_X1 U6138 ( .A1(n10057), .A2(n4490), .ZN(n4488) );
  NAND2_X1 U6139 ( .A1(n4354), .A2(n6608), .ZN(n6609) );
  NAND2_X1 U6140 ( .A1(n6605), .A2(n4355), .ZN(n4354) );
  NAND2_X1 U6141 ( .A1(n4576), .A2(n4324), .ZN(n4574) );
  OAI21_X1 U6142 ( .B1(n4974), .B2(n5314), .A(n4986), .ZN(n5378) );
  NAND2_X1 U6143 ( .A1(n6571), .A2(n6572), .ZN(n4577) );
  NAND2_X1 U6144 ( .A1(n4360), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6419) );
  OR2_X1 U6145 ( .A1(n9524), .A2(n9611), .ZN(n9525) );
  NAND2_X1 U6146 ( .A1(n9525), .A2(n4381), .ZN(n9618) );
  OAI21_X2 U6147 ( .B1(n8132), .B2(n8099), .A(n8100), .ZN(n9222) );
  AND2_X4 U6148 ( .A1(n4362), .A2(n7604), .ZN(n8306) );
  NAND3_X1 U6149 ( .A1(n6702), .A2(n7235), .A3(n7621), .ZN(n4362) );
  INV_X1 U6150 ( .A(n7177), .ZN(n4714) );
  NAND3_X1 U6151 ( .A1(n6585), .A2(n6587), .A3(n4282), .ZN(n6586) );
  NAND2_X1 U6152 ( .A1(n4596), .A2(n4595), .ZN(n4594) );
  AOI21_X1 U6153 ( .B1(n4364), .B2(n6634), .A(n6633), .ZN(n6635) );
  NAND2_X1 U6154 ( .A1(n4588), .A2(n4321), .ZN(n4364) );
  NAND2_X1 U6155 ( .A1(n4366), .A2(n6611), .ZN(n6614) );
  NAND3_X1 U6156 ( .A1(n6609), .A2(n8646), .A3(n6610), .ZN(n4366) );
  NAND2_X1 U6157 ( .A1(n6578), .A2(n4277), .ZN(n4581) );
  NAND2_X1 U6158 ( .A1(n4627), .A2(n5024), .ZN(n5528) );
  NAND2_X1 U6159 ( .A1(n4245), .A2(n4749), .ZN(n4748) );
  NAND3_X1 U6160 ( .A1(n9513), .A2(n4368), .A3(n9505), .ZN(n9616) );
  OR2_X1 U6161 ( .A1(n5228), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n5159) );
  INV_X1 U6162 ( .A(n9502), .ZN(n9504) );
  NAND2_X1 U6163 ( .A1(n4759), .A2(n4760), .ZN(n7873) );
  AOI21_X2 U6164 ( .B1(n8227), .B2(n10080), .A(n8226), .ZN(n8854) );
  OAI21_X1 U6165 ( .B1(n10064), .B2(n4490), .A(n7763), .ZN(n4489) );
  NAND2_X1 U6166 ( .A1(n5075), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5072) );
  NAND4_X1 U6167 ( .A1(n5070), .A2(n4663), .A3(n5069), .A4(n5068), .ZN(n5075)
         );
  NAND2_X2 U6168 ( .A1(n5078), .A2(n5073), .ZN(n7071) );
  NAND3_X1 U6169 ( .A1(n7548), .A2(n7550), .A3(n7549), .ZN(n7551) );
  NAND3_X1 U6170 ( .A1(n9344), .A2(n9343), .A3(n9454), .ZN(n4370) );
  NAND2_X1 U6171 ( .A1(n4602), .A2(n4601), .ZN(n4963) );
  AOI211_X2 U6172 ( .C1(n9607), .C2(n9511), .A(n9510), .B(n9509), .ZN(n9512)
         );
  AND2_X2 U6173 ( .A1(n9209), .A2(n4371), .ZN(n9306) );
  NOR2_X2 U6174 ( .A1(n9456), .A2(n9561), .ZN(n9421) );
  XNOR2_X2 U6175 ( .A(n5166), .B(P1_IR_REG_2__SCAN_IN), .ZN(n7087) );
  OAI211_X1 U6176 ( .C1(n9203), .C2(n9201), .A(n9200), .B(n4525), .ZN(n4524)
         );
  NAND2_X1 U6177 ( .A1(n4527), .A2(n4524), .ZN(n9206) );
  XNOR2_X1 U6178 ( .A(n4374), .B(n8637), .ZN(n6490) );
  NAND4_X1 U6179 ( .A1(n6489), .A2(n6492), .A3(n8244), .A4(n6493), .ZN(n4374)
         );
  OAI21_X1 U6180 ( .B1(n4929), .B2(n4928), .A(n5151), .ZN(n4931) );
  NAND4_X1 U6181 ( .A1(n4583), .A2(n6658), .A3(n4387), .A4(n4582), .ZN(
        P2_U3244) );
  OAI21_X2 U6182 ( .B1(n8085), .B2(n8084), .A(n8083), .ZN(n8269) );
  NAND3_X2 U6183 ( .A1(n6072), .A2(n6071), .A3(n6216), .ZN(n6081) );
  XNOR2_X2 U6184 ( .A(n8309), .B(n8308), .ZN(n8329) );
  OAI21_X1 U6185 ( .B1(n4252), .B2(n4380), .A(n4379), .ZN(n4947) );
  INV_X1 U6186 ( .A(n7853), .ZN(n4444) );
  NAND2_X1 U6187 ( .A1(n9373), .A2(n9259), .ZN(n4461) );
  INV_X1 U6188 ( .A(n7889), .ZN(n7856) );
  NAND2_X1 U6189 ( .A1(n5078), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5079) );
  NOR2_X2 U6190 ( .A1(n5534), .A2(n5519), .ZN(n4384) );
  NAND2_X2 U6191 ( .A1(n9239), .A2(n9240), .ZN(n9263) );
  INV_X1 U6192 ( .A(n4634), .ZN(n4630) );
  NAND2_X1 U6193 ( .A1(n4581), .A2(n8781), .ZN(n4580) );
  INV_X2 U6194 ( .A(n6081), .ZN(n6082) );
  AOI21_X1 U6195 ( .B1(n6596), .B2(n6582), .A(n6581), .ZN(n6584) );
  AOI21_X1 U6196 ( .B1(n6563), .B2(n6562), .A(n4574), .ZN(n4573) );
  OAI21_X1 U6197 ( .B1(n6616), .B2(n4590), .A(n4323), .ZN(n4589) );
  NOR2_X1 U6198 ( .A1(n10065), .A2(n4391), .ZN(n4388) );
  NAND2_X1 U6199 ( .A1(n8643), .A2(n4833), .ZN(n4394) );
  NAND2_X1 U6200 ( .A1(n4399), .A2(n4397), .ZN(n4396) );
  NAND2_X1 U6201 ( .A1(n4396), .A2(n4853), .ZN(n8664) );
  NAND2_X1 U6202 ( .A1(n6651), .A2(n6081), .ZN(n9002) );
  NAND3_X1 U6203 ( .A1(n4472), .A2(n4471), .A3(n8527), .ZN(n4406) );
  INV_X2 U6204 ( .A(n6859), .ZN(n6861) );
  NAND2_X2 U6205 ( .A1(n4472), .A2(n4471), .ZN(n6859) );
  NAND2_X1 U6206 ( .A1(n9050), .A2(n4407), .ZN(n4411) );
  OR3_X1 U6207 ( .A1(n9050), .A2(n4410), .A3(n4409), .ZN(n4412) );
  OR2_X1 U6208 ( .A1(n9050), .A2(n4413), .ZN(n9135) );
  NAND3_X1 U6209 ( .A1(n4412), .A2(n9134), .A3(n4411), .ZN(n9011) );
  AND2_X1 U6210 ( .A1(n5994), .A2(n5995), .ZN(n4418) );
  OR2_X1 U6211 ( .A1(n5068), .A2(n9779), .ZN(n4420) );
  NAND2_X1 U6212 ( .A1(n4421), .A2(n4419), .ZN(n4913) );
  OR2_X1 U6213 ( .A1(n5196), .A2(n9779), .ZN(n4421) );
  NAND3_X1 U6214 ( .A1(n5915), .A2(n4326), .A3(n8122), .ZN(n4425) );
  INV_X1 U6215 ( .A(n4428), .ZN(n4427) );
  NAND2_X1 U6216 ( .A1(n9024), .A2(n5948), .ZN(n4428) );
  NAND3_X1 U6217 ( .A1(n4744), .A2(n5154), .A3(n4903), .ZN(n5197) );
  NAND2_X1 U6218 ( .A1(n5609), .A2(n5653), .ZN(n4439) );
  AOI21_X1 U6219 ( .B1(n5609), .B2(n4435), .A(n4329), .ZN(n4438) );
  XNOR2_X1 U6220 ( .A(n5829), .B(n7426), .ZN(n5834) );
  INV_X1 U6221 ( .A(n5834), .ZN(n5831) );
  MUX2_X1 U6222 ( .A(n7119), .B(n4987), .S(n4251), .Z(n4989) );
  MUX2_X1 U6223 ( .A(n7172), .B(n7171), .S(n4440), .Z(n4994) );
  MUX2_X1 U6224 ( .A(n7218), .B(n7220), .S(n4440), .Z(n4999) );
  MUX2_X1 U6225 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n4440), .Z(n5004) );
  MUX2_X1 U6226 ( .A(n7388), .B(n7386), .S(n4440), .Z(n5007) );
  MUX2_X1 U6227 ( .A(n9750), .B(n5025), .S(n4440), .Z(n5027) );
  MUX2_X1 U6228 ( .A(n7507), .B(n7640), .S(n4440), .Z(n5013) );
  MUX2_X1 U6229 ( .A(n9646), .B(n7990), .S(n4440), .Z(n5031) );
  MUX2_X1 U6230 ( .A(n7622), .B(n9755), .S(n4440), .Z(n5017) );
  MUX2_X1 U6231 ( .A(n7745), .B(n8159), .S(n4440), .Z(n5021) );
  MUX2_X1 U6232 ( .A(n9001), .B(n9796), .S(n4440), .Z(n5039) );
  MUX2_X1 U6233 ( .A(n9757), .B(n9724), .S(n4440), .Z(n5052) );
  MUX2_X1 U6234 ( .A(n9733), .B(n5044), .S(n4440), .Z(n5046) );
  MUX2_X1 U6235 ( .A(n9665), .B(n9786), .S(n4440), .Z(n5097) );
  NAND2_X2 U6236 ( .A1(P1_U3084), .A2(n4440), .ZN(n9798) );
  MUX2_X1 U6237 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(n8984), .S(n4440), .Z(n5077) );
  NAND2_X2 U6238 ( .A1(n4447), .A2(n5240), .ZN(n5842) );
  NAND2_X1 U6239 ( .A1(n4447), .A2(n4445), .ZN(n5706) );
  NAND2_X1 U6240 ( .A1(n6737), .A2(n5586), .ZN(n4447) );
  NAND2_X1 U6241 ( .A1(n4449), .A2(n8136), .ZN(n4448) );
  NAND2_X1 U6242 ( .A1(n4448), .A2(n4874), .ZN(n9447) );
  NAND2_X1 U6243 ( .A1(n4452), .A2(n4340), .ZN(P1_U3518) );
  NAND2_X1 U6244 ( .A1(n9317), .A2(n4453), .ZN(n9523) );
  NOR2_X2 U6245 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n6094) );
  INV_X1 U6246 ( .A(n4466), .ZN(n8246) );
  NAND2_X1 U6247 ( .A1(n7808), .A2(n4470), .ZN(n4469) );
  AOI21_X1 U6248 ( .B1(n6652), .B2(P2_IR_REG_28__SCAN_IN), .A(n6074), .ZN(
        n4472) );
  INV_X1 U6249 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6317) );
  NAND2_X1 U6250 ( .A1(n6314), .A2(n4483), .ZN(n4480) );
  NAND2_X1 U6251 ( .A1(n4480), .A2(n4481), .ZN(n8772) );
  OAI21_X1 U6252 ( .B1(n4488), .B2(n4489), .A(n6509), .ZN(n7769) );
  NAND2_X1 U6253 ( .A1(n6127), .A2(n6126), .ZN(n7614) );
  OAI21_X2 U6254 ( .B1(n7873), .B2(n4504), .A(n6566), .ZN(n8041) );
  NAND2_X1 U6255 ( .A1(n6942), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n4505) );
  INV_X1 U6256 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n4511) );
  NAND2_X2 U6257 ( .A1(n4507), .A2(n4512), .ZN(n8527) );
  INV_X1 U6258 ( .A(n4508), .ZN(n4507) );
  OAI21_X1 U6259 ( .B1(n9003), .B2(n4513), .A(n4510), .ZN(n4508) );
  NAND3_X1 U6260 ( .A1(n9003), .A2(n4513), .A3(P2_IR_REG_31__SCAN_IN), .ZN(
        n4512) );
  OAI21_X1 U6261 ( .B1(n8527), .B2(n6886), .A(n4509), .ZN(n8526) );
  NAND2_X1 U6262 ( .A1(n8527), .A2(n6886), .ZN(n4509) );
  NAND2_X1 U6263 ( .A1(n7137), .A2(n4253), .ZN(n4529) );
  MUX2_X1 U6264 ( .A(P1_REG2_REG_1__SCAN_IN), .B(n5128), .S(n6980), .Z(n6989)
         );
  XNOR2_X2 U6265 ( .A(n4530), .B(P1_IR_REG_1__SCAN_IN), .ZN(n6980) );
  OAI21_X1 U6266 ( .B1(n4539), .B2(n4313), .A(n4536), .ZN(n5396) );
  AOI21_X1 U6267 ( .B1(n5261), .B2(n7557), .A(n4540), .ZN(n4539) );
  OR2_X1 U6268 ( .A1(n5475), .A2(n4546), .ZN(n4542) );
  NAND2_X1 U6269 ( .A1(n5475), .A2(n4549), .ZN(n4541) );
  NAND2_X1 U6270 ( .A1(n4542), .A2(n4543), .ZN(n5550) );
  AND2_X2 U6271 ( .A1(n5109), .A2(n5083), .ZN(n5563) );
  NAND3_X1 U6272 ( .A1(n5109), .A2(n5083), .A3(P1_REG3_REG_1__SCAN_IN), .ZN(
        n4558) );
  NAND2_X2 U6273 ( .A1(n9785), .A2(n8219), .ZN(n5180) );
  NAND3_X1 U6274 ( .A1(n8219), .A2(n9785), .A3(P1_REG0_REG_1__SCAN_IN), .ZN(
        n4556) );
  AND2_X2 U6275 ( .A1(n5109), .A2(n8219), .ZN(n5564) );
  INV_X1 U6276 ( .A(n5563), .ZN(n5228) );
  NAND4_X1 U6277 ( .A1(n5070), .A2(n4712), .A3(n5069), .A4(n5068), .ZN(n5078)
         );
  NAND2_X1 U6278 ( .A1(n7417), .A2(n5628), .ZN(n7530) );
  NAND2_X1 U6279 ( .A1(n7323), .A2(n4559), .ZN(n7417) );
  XNOR2_X1 U6280 ( .A(n7530), .B(n7096), .ZN(n5223) );
  NAND3_X1 U6281 ( .A1(n7193), .A2(n7436), .A3(n5618), .ZN(n4561) );
  NAND3_X1 U6282 ( .A1(n4561), .A2(n5697), .A3(n4560), .ZN(n5742) );
  NAND2_X1 U6283 ( .A1(n4562), .A2(n5144), .ZN(n7437) );
  INV_X1 U6284 ( .A(n5144), .ZN(n4563) );
  NAND2_X1 U6285 ( .A1(n6635), .A2(n4584), .ZN(n4583) );
  OR2_X2 U6286 ( .A1(n4587), .A2(n4586), .ZN(n4584) );
  INV_X1 U6287 ( .A(n6657), .ZN(n4586) );
  AND2_X1 U6288 ( .A1(n6636), .A2(n6637), .ZN(n4587) );
  NAND3_X1 U6289 ( .A1(n4589), .A2(n6622), .A3(n8244), .ZN(n4588) );
  NAND3_X1 U6290 ( .A1(n7813), .A2(n6553), .A3(n6630), .ZN(n4591) );
  INV_X1 U6291 ( .A(n5412), .ZN(n4596) );
  NAND2_X1 U6292 ( .A1(n5219), .A2(n4322), .ZN(n4601) );
  NAND2_X1 U6293 ( .A1(n5050), .A2(n4613), .ZN(n4608) );
  OAI21_X1 U6294 ( .B1(n5050), .B2(n4617), .A(n4615), .ZN(n5099) );
  NAND2_X1 U6295 ( .A1(n4608), .A2(n4609), .ZN(n5090) );
  NAND2_X1 U6296 ( .A1(n5050), .A2(n5049), .ZN(n5117) );
  OR2_X1 U6297 ( .A1(n5490), .A2(n4622), .ZN(n4618) );
  NAND2_X1 U6298 ( .A1(n5490), .A2(n4621), .ZN(n4620) );
  OR2_X1 U6299 ( .A1(n5490), .A2(n5489), .ZN(n4627) );
  NAND2_X1 U6300 ( .A1(n8999), .A2(n5586), .ZN(n5575) );
  INV_X1 U6301 ( .A(n4790), .ZN(n4789) );
  NAND3_X2 U6302 ( .A1(n4639), .A2(n5136), .A3(n4641), .ZN(n7277) );
  INV_X1 U6303 ( .A(n5694), .ZN(n4640) );
  INV_X1 U6304 ( .A(n7187), .ZN(n7193) );
  NAND2_X1 U6305 ( .A1(n9406), .A2(n4644), .ZN(n4643) );
  NAND2_X1 U6306 ( .A1(n7843), .A2(n4649), .ZN(n4648) );
  NAND2_X1 U6307 ( .A1(n4648), .A2(n4647), .ZN(n8132) );
  NAND2_X1 U6308 ( .A1(n7544), .A2(n4659), .ZN(n4655) );
  NAND2_X1 U6309 ( .A1(n4655), .A2(n4656), .ZN(n7835) );
  NAND2_X1 U6310 ( .A1(n9241), .A2(n4278), .ZN(n4673) );
  NAND2_X1 U6311 ( .A1(n4677), .A2(n9502), .ZN(n9518) );
  NAND2_X1 U6312 ( .A1(n9241), .A2(n9240), .ZN(n9303) );
  NAND2_X1 U6313 ( .A1(n4682), .A2(n4681), .ZN(n8178) );
  NAND3_X1 U6314 ( .A1(n7164), .A2(n7163), .A3(n8161), .ZN(n4682) );
  NAND2_X1 U6315 ( .A1(n7164), .A2(n7163), .ZN(n4684) );
  NAND2_X1 U6316 ( .A1(n5898), .A2(n4686), .ZN(n4685) );
  NAND2_X1 U6317 ( .A1(n5962), .A2(n4693), .ZN(n4692) );
  NAND2_X1 U6318 ( .A1(n4265), .A2(n4697), .ZN(n4702) );
  NAND3_X1 U6319 ( .A1(n4702), .A2(n4700), .A3(n4698), .ZN(P1_U3218) );
  NAND2_X1 U6320 ( .A1(n9135), .A2(n4701), .ZN(n4700) );
  NAND3_X1 U6321 ( .A1(n7210), .A2(n6672), .A3(n4714), .ZN(n7176) );
  NAND2_X1 U6322 ( .A1(n7176), .A2(n6677), .ZN(n4713) );
  NAND2_X1 U6323 ( .A1(n7970), .A2(n4715), .ZN(n10009) );
  NAND2_X1 U6324 ( .A1(n8391), .A2(n4719), .ZN(n4718) );
  OAI21_X1 U6325 ( .B1(n8399), .B2(n4726), .A(n4723), .ZN(n8286) );
  INV_X2 U6326 ( .A(n8310), .ZN(n8354) );
  NAND2_X4 U6327 ( .A1(n4247), .A2(n4742), .ZN(n8310) );
  OR2_X2 U6328 ( .A1(n4743), .A2(n6709), .ZN(n6702) );
  INV_X2 U6329 ( .A(n7621), .ZN(n4743) );
  NAND2_X2 U6330 ( .A1(n7508), .A2(n8637), .ZN(n6712) );
  XNOR2_X2 U6331 ( .A(n6464), .B(n6465), .ZN(n7508) );
  NOR2_X2 U6332 ( .A1(n9944), .A2(n4746), .ZN(n7533) );
  NAND3_X1 U6333 ( .A1(n9958), .A2(n9952), .A3(n9964), .ZN(n4746) );
  NOR2_X2 U6334 ( .A1(n7481), .A2(n4748), .ZN(n7710) );
  NOR2_X2 U6335 ( .A1(n9981), .A2(n5842), .ZN(n4749) );
  INV_X1 U6336 ( .A(n4751), .ZN(n7578) );
  INV_X1 U6337 ( .A(n4756), .ZN(n8101) );
  NAND3_X2 U6338 ( .A1(n9408), .A2(n9352), .A3(n4258), .ZN(n9327) );
  NAND2_X1 U6339 ( .A1(n6236), .A2(n4279), .ZN(n4759) );
  NAND2_X1 U6340 ( .A1(n6082), .A2(n4328), .ZN(n8985) );
  NAND2_X1 U6341 ( .A1(n8644), .A2(n4769), .ZN(n4768) );
  OAI21_X1 U6342 ( .B1(n8644), .B2(n4771), .A(n4769), .ZN(n8604) );
  NAND2_X1 U6343 ( .A1(n4787), .A2(n4788), .ZN(n4786) );
  NAND2_X1 U6344 ( .A1(n6350), .A2(n4781), .ZN(n4785) );
  NAND2_X1 U6345 ( .A1(n4788), .A2(n6595), .ZN(n4782) );
  CLKBUF_X1 U6346 ( .A(n4785), .Z(n4783) );
  NAND4_X1 U6347 ( .A1(n4785), .A2(n4784), .A3(n4282), .A4(n8694), .ZN(n8693)
         );
  INV_X1 U6348 ( .A(n6359), .ZN(n4788) );
  NAND2_X1 U6349 ( .A1(n8657), .A2(n4793), .ZN(n4791) );
  NAND2_X1 U6350 ( .A1(n8674), .A2(n4318), .ZN(n4792) );
  OR2_X2 U6351 ( .A1(n8674), .A2(n8675), .ZN(n4794) );
  INV_X2 U6352 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n4796) );
  OAI211_X1 U6353 ( .C1(n4808), .C2(n4807), .A(n4806), .B(n4805), .ZN(n4804)
         );
  OR2_X1 U6354 ( .A1(n6143), .A2(SI_1_), .ZN(n4806) );
  NAND3_X1 U6355 ( .A1(n4812), .A2(n10138), .A3(n4811), .ZN(n10088) );
  OR2_X1 U6356 ( .A1(n8846), .A2(n4337), .ZN(n4813) );
  NAND2_X1 U6357 ( .A1(n4813), .A2(n4814), .ZN(P2_U3551) );
  OAI21_X1 U6358 ( .B1(n8846), .B2(n4339), .A(n4817), .ZN(P2_U3519) );
  NAND2_X1 U6359 ( .A1(n4831), .A2(n4935), .ZN(n5171) );
  INV_X1 U6360 ( .A(n5172), .ZN(n4830) );
  OR2_X1 U6361 ( .A1(n8867), .A2(n8615), .ZN(n4844) );
  OAI22_X1 U6362 ( .A1(n8236), .A2(n4847), .B1(n4848), .B2(n8238), .ZN(n8737)
         );
  NAND2_X1 U6363 ( .A1(n8737), .A2(n4851), .ZN(n8240) );
  INV_X1 U6364 ( .A(n8238), .ZN(n4852) );
  NAND2_X1 U6365 ( .A1(n5234), .A2(n4946), .ZN(n4866) );
  NAND3_X1 U6366 ( .A1(n4867), .A2(n7849), .A3(n7850), .ZN(n7852) );
  NAND3_X1 U6367 ( .A1(n7718), .A2(n7717), .A3(n7848), .ZN(n4867) );
  NAND2_X1 U6368 ( .A1(n4868), .A2(n7917), .ZN(n7918) );
  NAND2_X1 U6369 ( .A1(n4868), .A2(n7720), .ZN(n7721) );
  NAND2_X1 U6370 ( .A1(n9437), .A2(n4872), .ZN(n4871) );
  OAI21_X1 U6371 ( .B1(n9246), .B2(n9245), .A(n9244), .ZN(n9477) );
  NAND2_X1 U6372 ( .A1(n7856), .A2(n7855), .ZN(n7892) );
  OAI21_X1 U6373 ( .B1(n4884), .B2(n8108), .A(n8107), .ZN(n4881) );
  NAND2_X1 U6374 ( .A1(n7856), .A2(n4883), .ZN(n4882) );
  NAND2_X1 U6375 ( .A1(n4888), .A2(n4886), .ZN(n4885) );
  CLKBUF_X1 U6376 ( .A(n5201), .Z(n5204) );
  NAND2_X1 U6377 ( .A1(n7712), .A2(n7711), .ZN(n8006) );
  INV_X1 U6378 ( .A(n7713), .ZN(n7712) );
  OR2_X1 U6379 ( .A1(n8022), .A2(n7878), .ZN(n8036) );
  XNOR2_X1 U6380 ( .A(n5573), .B(n5572), .ZN(n8999) );
  CLKBUF_X1 U6381 ( .A(n8737), .Z(n8739) );
  XNOR2_X1 U6382 ( .A(n5505), .B(n5504), .ZN(n8091) );
  XNOR2_X1 U6383 ( .A(n5090), .B(n5089), .ZN(n8218) );
  INV_X1 U6384 ( .A(n6706), .ZN(n6704) );
  INV_X1 U6385 ( .A(n7189), .ZN(n7624) );
  OR2_X1 U6386 ( .A1(n5783), .A2(n6661), .ZN(n6760) );
  CLKBUF_X1 U6387 ( .A(n7835), .Z(n7916) );
  OR2_X1 U6388 ( .A1(n6150), .A2(n6865), .ZN(n6128) );
  OR2_X1 U6389 ( .A1(n6148), .A2(n6147), .ZN(n6154) );
  NAND2_X1 U6390 ( .A1(n6100), .A2(n6063), .ZN(n6101) );
  INV_X1 U6391 ( .A(n7689), .ZN(n6133) );
  XNOR2_X1 U6392 ( .A(n8260), .B(n8259), .ZN(n8846) );
  XNOR2_X1 U6393 ( .A(n8222), .B(n8221), .ZN(n8227) );
  OR2_X1 U6394 ( .A1(n8368), .A2(n6421), .ZN(n6427) );
  OR2_X1 U6395 ( .A1(n8639), .A2(n6421), .ZN(n6409) );
  OR2_X1 U6396 ( .A1(n6149), .A2(n6887), .ZN(n6153) );
  CLKBUF_X1 U6397 ( .A(n5742), .Z(n7392) );
  NAND4_X1 U6398 ( .A1(n4276), .A2(n4902), .A3(n6129), .A4(n6128), .ZN(n6146)
         );
  AND2_X1 U6399 ( .A1(n6712), .A2(n10116), .ZN(n8958) );
  INV_X1 U6400 ( .A(n6014), .ZN(n7992) );
  NAND2_X1 U6401 ( .A1(n8988), .A2(n8993), .ZN(n6149) );
  OR2_X1 U6402 ( .A1(n6663), .A2(n6973), .ZN(n4891) );
  AND2_X1 U6403 ( .A1(n4898), .A2(n9134), .ZN(n4892) );
  OR2_X1 U6404 ( .A1(n9321), .A2(n9263), .ZN(n4893) );
  NAND2_X1 U6405 ( .A1(n5725), .A2(n9260), .ZN(n9360) );
  AND2_X1 U6406 ( .A1(n4997), .A2(n4996), .ZN(n4895) );
  AND2_X1 U6407 ( .A1(n4985), .A2(SI_14_), .ZN(n4897) );
  XOR2_X1 U6408 ( .A(n6043), .B(n6042), .Z(n4898) );
  INV_X1 U6409 ( .A(n9285), .ZN(n9292) );
  NOR2_X1 U6410 ( .A1(n9157), .A2(n7400), .ZN(n7313) );
  NOR2_X1 U6411 ( .A1(n7662), .A2(n7661), .ZN(n4900) );
  AND2_X1 U6412 ( .A1(n8632), .A2(n8630), .ZN(n4901) );
  INV_X1 U6413 ( .A(n9606), .ZN(n7711) );
  OR2_X1 U6414 ( .A1(n6149), .A2(n6886), .ZN(n4902) );
  INV_X1 U6415 ( .A(n6479), .ZN(n6145) );
  INV_X1 U6416 ( .A(n8847), .ZN(n6456) );
  OR2_X1 U6417 ( .A1(n9022), .A2(n9119), .ZN(n5948) );
  AND2_X1 U6418 ( .A1(n9269), .A2(n9268), .ZN(n9270) );
  AND2_X1 U6419 ( .A1(n7529), .A2(n7525), .ZN(n7472) );
  INV_X1 U6420 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n5071) );
  INV_X1 U6421 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n4903) );
  INV_X1 U6422 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n6209) );
  INV_X1 U6423 ( .A(n6364), .ZN(n6366) );
  AND2_X1 U6424 ( .A1(n6519), .A2(n7614), .ZN(n6528) );
  AND2_X1 U6425 ( .A1(n7823), .A2(n7819), .ZN(n7817) );
  OR2_X1 U6426 ( .A1(n7066), .A2(n5794), .ZN(n5798) );
  INV_X1 U6427 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n5290) );
  INV_X1 U6428 ( .A(n5842), .ZN(n7482) );
  INV_X1 U6429 ( .A(n5431), .ZN(n5003) );
  INV_X1 U6430 ( .A(n5301), .ZN(n5313) );
  INV_X1 U6431 ( .A(n5233), .ZN(n4946) );
  NAND2_X1 U6432 ( .A1(n8329), .A2(n8311), .ZN(n8313) );
  NAND2_X1 U6433 ( .A1(n6366), .A2(n6365), .ZN(n6376) );
  INV_X1 U6434 ( .A(n8988), .ZN(n6087) );
  NAND2_X1 U6435 ( .A1(n8909), .A2(n8743), .ZN(n6582) );
  NOR2_X1 U6436 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n6070) );
  INV_X1 U6437 ( .A(n5564), .ZN(n5224) );
  AND2_X1 U6438 ( .A1(n6783), .A2(n9792), .ZN(n6846) );
  INV_X1 U6439 ( .A(n9405), .ZN(n9254) );
  AND2_X1 U6440 ( .A1(n9340), .A2(n9338), .ZN(n9238) );
  OR2_X1 U6441 ( .A1(n9776), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6019) );
  NAND2_X1 U6442 ( .A1(n5573), .A2(n5572), .ZN(n5043) );
  NAND2_X1 U6443 ( .A1(n4994), .A2(n4993), .ZN(n4997) );
  AND2_X1 U6444 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_10__SCAN_IN), 
        .ZN(n6078) );
  OR2_X1 U6445 ( .A1(n8362), .A2(n6708), .ZN(n8386) );
  OR3_X1 U6446 ( .A1(n6419), .A2(n8322), .A3(n8369), .ZN(n6430) );
  INV_X1 U6447 ( .A(n6273), .ZN(n6385) );
  OR2_X1 U6448 ( .A1(n7263), .A2(n7264), .ZN(n7378) );
  OR2_X1 U6449 ( .A1(n8550), .A2(n8551), .ZN(n8570) );
  AOI22_X1 U6450 ( .A1(n8616), .A2(n10058), .B1(n8261), .B2(n8511), .ZN(n8225)
         );
  AND2_X1 U6451 ( .A1(n4743), .A2(n6709), .ZN(n6855) );
  AND2_X1 U6452 ( .A1(n6595), .A2(n6582), .ZN(n8767) );
  NAND2_X1 U6453 ( .A1(n7826), .A2(n7825), .ZN(n7876) );
  NAND2_X1 U6454 ( .A1(n7596), .A2(n7595), .ZN(n8825) );
  OR3_X1 U6455 ( .A1(n7915), .A2(n8092), .A3(n9002), .ZN(n6856) );
  NOR2_X1 U6456 ( .A1(n6012), .A2(n4259), .ZN(n6013) );
  INV_X1 U6457 ( .A(n5986), .ZN(n9047) );
  INV_X2 U6458 ( .A(n5802), .ZN(n5970) );
  INV_X1 U6459 ( .A(n9137), .ZN(n9128) );
  NAND2_X2 U6460 ( .A1(n7071), .A2(n9211), .ZN(n5135) );
  OR2_X1 U6461 ( .A1(n9602), .A2(n7276), .ZN(n9460) );
  AND2_X1 U6462 ( .A1(n4462), .A2(n9257), .ZN(n9396) );
  INV_X1 U6463 ( .A(n7642), .ZN(n7198) );
  INV_X1 U6464 ( .A(n9454), .ZN(n9479) );
  NAND2_X1 U6465 ( .A1(n5010), .A2(n5009), .ZN(n5450) );
  NAND2_X1 U6466 ( .A1(n4992), .A2(n4991), .ZN(n5377) );
  NOR2_X1 U6467 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10207), .ZN(n9815) );
  INV_X1 U6468 ( .A(n8386), .ZN(n8493) );
  INV_X1 U6469 ( .A(n10010), .ZN(n10043) );
  AND2_X1 U6470 ( .A1(n6893), .A2(n6891), .ZN(n8540) );
  AND2_X1 U6471 ( .A1(n6863), .A2(n6862), .ZN(n8542) );
  INV_X1 U6472 ( .A(n8564), .ZN(n8593) );
  AND2_X1 U6473 ( .A1(n8838), .A2(n8950), .ZN(n8813) );
  INV_X1 U6474 ( .A(n8836), .ZN(n10093) );
  INV_X1 U6475 ( .A(n8790), .ZN(n10099) );
  NOR2_X1 U6476 ( .A1(n10110), .A2(n6701), .ZN(n7600) );
  INV_X1 U6477 ( .A(n8949), .ZN(n10155) );
  AND2_X1 U6478 ( .A1(n6697), .A2(n6696), .ZN(n10101) );
  INV_X1 U6479 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6639) );
  AND2_X1 U6480 ( .A1(n6241), .A2(n6249), .ZN(n7153) );
  AND2_X1 U6481 ( .A1(n6662), .A2(n6760), .ZN(n6783) );
  AND2_X1 U6482 ( .A1(n9247), .A2(n5446), .ZN(n9478) );
  AND2_X1 U6483 ( .A1(n9463), .A2(n7330), .ZN(n9491) );
  AND2_X1 U6484 ( .A1(n7196), .A2(n7195), .ZN(n9451) );
  NAND2_X2 U6485 ( .A1(n7286), .A2(n9460), .ZN(n9463) );
  INV_X1 U6486 ( .A(n9607), .ZN(n9982) );
  OR2_X1 U6487 ( .A1(n7096), .A2(n7198), .ZN(n9602) );
  AND2_X1 U6488 ( .A1(n7570), .A2(n7545), .ZN(n9988) );
  AND2_X1 U6489 ( .A1(n7098), .A2(n7097), .ZN(n7206) );
  INV_X1 U6490 ( .A(n8217), .ZN(n8587) );
  INV_X1 U6491 ( .A(n8893), .ZN(n8707) );
  INV_X1 U6492 ( .A(n8667), .ZN(n8877) );
  NAND2_X1 U6493 ( .A1(n6717), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10055) );
  OR2_X1 U6494 ( .A1(n8362), .A2(n8363), .ZN(n10010) );
  INV_X1 U6495 ( .A(n8355), .ZN(n8616) );
  INV_X1 U6496 ( .A(n8540), .ZN(n8590) );
  INV_X1 U6497 ( .A(n8542), .ZN(n8584) );
  INV_X1 U6498 ( .A(n10093), .ZN(n8717) );
  AND2_X1 U6499 ( .A1(n7607), .A2(n10090), .ZN(n8836) );
  OR2_X1 U6500 ( .A1(n8836), .A2(n7605), .ZN(n8790) );
  INV_X1 U6501 ( .A(n10176), .ZN(n10174) );
  INV_X1 U6502 ( .A(n10166), .ZN(n10165) );
  NOR2_X1 U6503 ( .A1(n10102), .A2(n10101), .ZN(n10112) );
  AND2_X1 U6504 ( .A1(n6713), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10111) );
  XNOR2_X1 U6505 ( .A(n6640), .B(n6639), .ZN(n7915) );
  INV_X1 U6506 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7218) );
  INV_X1 U6507 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6781) );
  INV_X1 U6508 ( .A(n7709), .ZN(n7959) );
  INV_X1 U6509 ( .A(n9533), .ZN(n9352) );
  INV_X1 U6510 ( .A(n9546), .ZN(n9394) );
  AOI21_X1 U6511 ( .B1(n5673), .B2(n5672), .A(n5671), .ZN(n5782) );
  INV_X1 U6512 ( .A(n9483), .ZN(n9223) );
  INV_X1 U6513 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n9807) );
  INV_X1 U6514 ( .A(n9911), .ZN(n9934) );
  AND2_X1 U6515 ( .A1(n9291), .A2(n9290), .ZN(n9517) );
  INV_X1 U6516 ( .A(n10003), .ZN(n10000) );
  OR2_X1 U6517 ( .A1(n9605), .A2(n9604), .ZN(n9774) );
  INV_X1 U6518 ( .A(n9991), .ZN(n9990) );
  INV_X1 U6519 ( .A(n9942), .ZN(n9943) );
  AND2_X1 U6520 ( .A1(n5783), .A2(n5668), .ZN(n9777) );
  INV_X1 U6521 ( .A(n6015), .ZN(n9799) );
  INV_X1 U6522 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7220) );
  INV_X1 U6523 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6780) );
  INV_X1 U6524 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6746) );
  NOR2_X1 U6525 ( .A1(n10216), .A2(n10215), .ZN(n10214) );
  INV_X1 U6526 ( .A(n8518), .ZN(P2_U3966) );
  NOR2_X1 U6527 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n4907) );
  NOR2_X1 U6528 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n4906) );
  NOR2_X1 U6529 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), .ZN(
        n4905) );
  NAND4_X1 U6530 ( .A1(n4907), .A2(n4906), .A3(n4905), .A4(n4904), .ZN(n4911)
         );
  NAND4_X1 U6531 ( .A1(n4909), .A2(n5356), .A3(n5413), .A4(n4908), .ZN(n4910)
         );
  INV_X1 U6532 ( .A(n4914), .ZN(n5658) );
  NAND2_X1 U6533 ( .A1(n5658), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n4915) );
  MUX2_X1 U6534 ( .A(P1_IR_REG_31__SCAN_IN), .B(n4915), .S(
        P1_IR_REG_19__SCAN_IN), .Z(n4916) );
  NAND2_X1 U6535 ( .A1(n4916), .A2(n5655), .ZN(n9277) );
  INV_X1 U6536 ( .A(n7096), .ZN(n5608) );
  INV_X1 U6537 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n9633) );
  INV_X1 U6538 ( .A(SI_2_), .ZN(n5150) );
  NAND2_X1 U6539 ( .A1(SI_0_), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n5132) );
  INV_X1 U6540 ( .A(SI_1_), .ZN(n5133) );
  NAND2_X1 U6541 ( .A1(n5132), .A2(n5133), .ZN(n4917) );
  NAND2_X1 U6542 ( .A1(n4917), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n4920) );
  INV_X1 U6543 ( .A(n5132), .ZN(n4918) );
  NAND2_X1 U6544 ( .A1(n4918), .A2(SI_1_), .ZN(n4919) );
  NAND2_X1 U6545 ( .A1(n4920), .A2(n4919), .ZN(n4921) );
  NAND2_X1 U6546 ( .A1(n4251), .A2(n4921), .ZN(n4927) );
  INV_X2 U6547 ( .A(n4250), .ZN(n6728) );
  NOR2_X1 U6548 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4924) );
  AND2_X1 U6549 ( .A1(SI_0_), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n5131) );
  INV_X1 U6550 ( .A(n5131), .ZN(n4923) );
  NAND2_X1 U6551 ( .A1(SI_1_), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n4922) );
  OAI21_X1 U6552 ( .B1(n4924), .B2(n4923), .A(n4922), .ZN(n4925) );
  NAND2_X1 U6553 ( .A1(n6728), .A2(n4925), .ZN(n4926) );
  NAND2_X1 U6554 ( .A1(n4927), .A2(n4926), .ZN(n5151) );
  INV_X1 U6555 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6740) );
  NAND2_X1 U6556 ( .A1(n4931), .A2(n4930), .ZN(n5163) );
  INV_X1 U6557 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n6723) );
  INV_X1 U6558 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U6559 ( .A1(n4250), .A2(n6744), .ZN(n4932) );
  INV_X1 U6560 ( .A(n4933), .ZN(n4934) );
  NAND2_X1 U6561 ( .A1(n4934), .A2(SI_3_), .ZN(n4935) );
  INV_X1 U6562 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6725) );
  INV_X1 U6563 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n4936) );
  MUX2_X1 U6564 ( .A(n6725), .B(n4936), .S(n4252), .Z(n4937) );
  INV_X1 U6565 ( .A(n4937), .ZN(n4938) );
  MUX2_X1 U6566 ( .A(n6727), .B(n6746), .S(n4252), .Z(n4939) );
  XNOR2_X1 U6567 ( .A(n4939), .B(SI_5_), .ZN(n5202) );
  NAND2_X1 U6568 ( .A1(n5201), .A2(n5202), .ZN(n4942) );
  INV_X1 U6569 ( .A(n4939), .ZN(n4940) );
  NAND2_X1 U6570 ( .A1(n4940), .A2(SI_5_), .ZN(n4941) );
  MUX2_X1 U6571 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .S(n4252), .Z(n4944) );
  NAND2_X1 U6572 ( .A1(n4944), .A2(SI_6_), .ZN(n4945) );
  NAND2_X1 U6573 ( .A1(n4947), .A2(SI_7_), .ZN(n4948) );
  MUX2_X1 U6574 ( .A(n6748), .B(n6750), .S(n4251), .Z(n4950) );
  INV_X1 U6575 ( .A(SI_8_), .ZN(n4949) );
  INV_X1 U6576 ( .A(n4950), .ZN(n4951) );
  NAND2_X1 U6577 ( .A1(n4951), .A2(SI_8_), .ZN(n4952) );
  MUX2_X1 U6578 ( .A(n6758), .B(n6757), .S(n4251), .Z(n4954) );
  INV_X1 U6579 ( .A(SI_9_), .ZN(n9632) );
  INV_X1 U6580 ( .A(n4954), .ZN(n4955) );
  NAND2_X1 U6581 ( .A1(n4955), .A2(SI_9_), .ZN(n4956) );
  MUX2_X1 U6582 ( .A(n6781), .B(n6780), .S(n4252), .Z(n4959) );
  INV_X1 U6583 ( .A(n4959), .ZN(n4957) );
  INV_X1 U6584 ( .A(n5280), .ZN(n4961) );
  INV_X1 U6585 ( .A(SI_10_), .ZN(n4958) );
  NAND2_X1 U6586 ( .A1(n4959), .A2(n4958), .ZN(n5281) );
  AND2_X1 U6587 ( .A1(n5278), .A2(n5281), .ZN(n4960) );
  INV_X1 U6588 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n4964) );
  MUX2_X1 U6589 ( .A(n6836), .B(n4964), .S(n4251), .Z(n4977) );
  INV_X1 U6590 ( .A(SI_13_), .ZN(n4966) );
  NAND2_X1 U6591 ( .A1(n4967), .A2(n4966), .ZN(n4972) );
  INV_X1 U6592 ( .A(n4967), .ZN(n4968) );
  NAND2_X1 U6593 ( .A1(n4968), .A2(SI_13_), .ZN(n4969) );
  NAND2_X1 U6594 ( .A1(n4972), .A2(n4969), .ZN(n4980) );
  INV_X1 U6595 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n4970) );
  MUX2_X1 U6596 ( .A(n7050), .B(n4970), .S(n4252), .Z(n4975) );
  INV_X1 U6597 ( .A(SI_12_), .ZN(n4971) );
  MUX2_X1 U6598 ( .A(n7016), .B(n7018), .S(n4252), .Z(n4984) );
  INV_X1 U6599 ( .A(n4975), .ZN(n4976) );
  NAND2_X1 U6600 ( .A1(n4976), .A2(SI_12_), .ZN(n5316) );
  INV_X1 U6601 ( .A(n4977), .ZN(n4978) );
  NAND2_X1 U6602 ( .A1(n4978), .A2(SI_11_), .ZN(n5315) );
  NAND2_X1 U6603 ( .A1(n5316), .A2(n5315), .ZN(n4979) );
  NOR2_X1 U6604 ( .A1(n4980), .A2(n4979), .ZN(n4981) );
  INV_X1 U6605 ( .A(n4984), .ZN(n4985) );
  INV_X1 U6606 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n4987) );
  INV_X1 U6607 ( .A(SI_15_), .ZN(n4988) );
  INV_X1 U6608 ( .A(n4989), .ZN(n4990) );
  NAND2_X1 U6609 ( .A1(n4990), .A2(SI_15_), .ZN(n4991) );
  INV_X1 U6610 ( .A(SI_16_), .ZN(n4993) );
  INV_X1 U6611 ( .A(n4994), .ZN(n4995) );
  NAND2_X1 U6612 ( .A1(n4995), .A2(SI_16_), .ZN(n4996) );
  INV_X1 U6613 ( .A(n4999), .ZN(n5000) );
  NAND2_X1 U6614 ( .A1(n5004), .A2(SI_18_), .ZN(n5005) );
  INV_X1 U6615 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7388) );
  INV_X1 U6616 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7386) );
  INV_X1 U6617 ( .A(SI_19_), .ZN(n5006) );
  INV_X1 U6618 ( .A(n5007), .ZN(n5008) );
  NAND2_X1 U6619 ( .A1(n5008), .A2(SI_19_), .ZN(n5009) );
  INV_X1 U6620 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7507) );
  INV_X1 U6621 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n7640) );
  INV_X1 U6622 ( .A(SI_20_), .ZN(n5012) );
  NAND2_X1 U6623 ( .A1(n5013), .A2(n5012), .ZN(n5016) );
  INV_X1 U6624 ( .A(n5013), .ZN(n5014) );
  NAND2_X1 U6625 ( .A1(n5014), .A2(SI_20_), .ZN(n5015) );
  INV_X1 U6626 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7622) );
  XNOR2_X1 U6627 ( .A(n5017), .B(SI_21_), .ZN(n5476) );
  INV_X1 U6628 ( .A(n5017), .ZN(n5018) );
  NAND2_X1 U6629 ( .A1(n5018), .A2(SI_21_), .ZN(n5019) );
  INV_X1 U6630 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7745) );
  INV_X1 U6631 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8159) );
  INV_X1 U6632 ( .A(SI_22_), .ZN(n9634) );
  INV_X1 U6633 ( .A(n5021), .ZN(n5022) );
  NAND2_X1 U6634 ( .A1(n5022), .A2(SI_22_), .ZN(n5023) );
  NAND2_X1 U6635 ( .A1(n5024), .A2(n5023), .ZN(n5489) );
  INV_X1 U6636 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n5025) );
  INV_X1 U6637 ( .A(SI_23_), .ZN(n5026) );
  NAND2_X1 U6638 ( .A1(n5027), .A2(n5026), .ZN(n5030) );
  INV_X1 U6639 ( .A(n5027), .ZN(n5028) );
  NAND2_X1 U6640 ( .A1(n5028), .A2(SI_23_), .ZN(n5029) );
  INV_X1 U6641 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n9646) );
  INV_X1 U6642 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n7990) );
  XNOR2_X1 U6643 ( .A(n5031), .B(SI_24_), .ZN(n5515) );
  INV_X1 U6644 ( .A(n5031), .ZN(n5032) );
  INV_X1 U6645 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8093) );
  INV_X1 U6646 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8096) );
  MUX2_X1 U6647 ( .A(n8093), .B(n8096), .S(n4251), .Z(n5034) );
  INV_X1 U6648 ( .A(SI_25_), .ZN(n5033) );
  NAND2_X1 U6649 ( .A1(n5034), .A2(n5033), .ZN(n5037) );
  INV_X1 U6650 ( .A(n5034), .ZN(n5035) );
  NAND2_X1 U6651 ( .A1(n5035), .A2(SI_25_), .ZN(n5036) );
  NAND2_X1 U6652 ( .A1(n5037), .A2(n5036), .ZN(n5504) );
  INV_X1 U6653 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n9001) );
  INV_X1 U6654 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9796) );
  INV_X1 U6655 ( .A(SI_26_), .ZN(n5038) );
  NAND2_X1 U6656 ( .A1(n5039), .A2(n5038), .ZN(n5042) );
  INV_X1 U6657 ( .A(n5039), .ZN(n5040) );
  NAND2_X1 U6658 ( .A1(n5040), .A2(SI_26_), .ZN(n5041) );
  INV_X1 U6659 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n9733) );
  INV_X1 U6660 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n5044) );
  INV_X1 U6661 ( .A(SI_27_), .ZN(n5045) );
  NAND2_X1 U6662 ( .A1(n5046), .A2(n5045), .ZN(n5049) );
  INV_X1 U6663 ( .A(n5046), .ZN(n5047) );
  NAND2_X1 U6664 ( .A1(n5047), .A2(SI_27_), .ZN(n5048) );
  INV_X1 U6665 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9757) );
  INV_X1 U6666 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n9724) );
  XNOR2_X1 U6667 ( .A(n5052), .B(SI_28_), .ZN(n5116) );
  INV_X1 U6668 ( .A(SI_28_), .ZN(n5051) );
  INV_X1 U6669 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9665) );
  INV_X1 U6670 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9786) );
  INV_X1 U6671 ( .A(SI_29_), .ZN(n5053) );
  AND2_X1 U6672 ( .A1(n5097), .A2(n5053), .ZN(n5056) );
  INV_X1 U6673 ( .A(n5097), .ZN(n5054) );
  NAND2_X1 U6674 ( .A1(n5054), .A2(SI_29_), .ZN(n5055) );
  MUX2_X1 U6675 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n6728), .Z(n5088) );
  INV_X1 U6676 ( .A(n5088), .ZN(n5058) );
  INV_X1 U6677 ( .A(SI_30_), .ZN(n5057) );
  NOR2_X1 U6678 ( .A1(n5058), .A2(n5057), .ZN(n5059) );
  INV_X1 U6679 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n5061) );
  INV_X1 U6680 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n5060) );
  MUX2_X1 U6681 ( .A(n5061), .B(n5060), .S(n6728), .Z(n5062) );
  XNOR2_X1 U6682 ( .A(n5062), .B(SI_31_), .ZN(n5063) );
  NOR2_X1 U6683 ( .A1(P1_IR_REG_19__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n5067) );
  NAND4_X1 U6684 ( .A1(n5067), .A2(n5066), .A3(n5653), .A4(n5065), .ZN(n5657)
         );
  MUX2_X2 U6685 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5072), .S(
        P1_IR_REG_28__SCAN_IN), .Z(n5073) );
  NAND2_X2 U6686 ( .A1(n5076), .A2(n5075), .ZN(n9211) );
  INV_X1 U6687 ( .A(n5081), .ZN(n9780) );
  XNOR2_X2 U6688 ( .A(n5082), .B(P1_IR_REG_30__SCAN_IN), .ZN(n5083) );
  INV_X1 U6689 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n5087) );
  NAND2_X1 U6690 ( .A1(n5564), .A2(P1_REG1_REG_31__SCAN_IN), .ZN(n5086) );
  INV_X1 U6691 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n5084) );
  OR2_X1 U6692 ( .A1(n5180), .A2(n5084), .ZN(n5085) );
  OAI211_X1 U6693 ( .C1(n5568), .C2(n5087), .A(n5086), .B(n5085), .ZN(n9213)
         );
  XNOR2_X1 U6694 ( .A(n5088), .B(SI_30_), .ZN(n5089) );
  NAND2_X1 U6695 ( .A1(n8218), .A2(n5586), .ZN(n5092) );
  AND2_X2 U6696 ( .A1(n5135), .A2(n6728), .ZN(n5164) );
  NAND2_X1 U6697 ( .A1(n5587), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n5091) );
  INV_X1 U6698 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n5095) );
  NAND2_X1 U6699 ( .A1(n5592), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n5094) );
  INV_X2 U6700 ( .A(n5180), .ZN(n5591) );
  NAND2_X1 U6701 ( .A1(n5591), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n5093) );
  OAI211_X1 U6702 ( .C1(n5596), .C2(n5095), .A(n5094), .B(n5093), .ZN(n9268)
         );
  INV_X1 U6703 ( .A(n9268), .ZN(n5647) );
  OR2_X1 U6704 ( .A1(n9217), .A2(n5647), .ZN(n5610) );
  AND2_X1 U6705 ( .A1(n5611), .A2(n7096), .ZN(n5607) );
  XNOR2_X1 U6706 ( .A(n5097), .B(SI_29_), .ZN(n5098) );
  NAND2_X1 U6707 ( .A1(n8992), .A2(n5586), .ZN(n5101) );
  NAND2_X1 U6708 ( .A1(n5164), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n5100) );
  INV_X1 U6709 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n5341) );
  INV_X1 U6710 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n8115) );
  INV_X1 U6711 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n9730) );
  INV_X1 U6712 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n9101) );
  INV_X1 U6713 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n9035) );
  INV_X1 U6714 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n5519) );
  INV_X1 U6715 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n5560) );
  OR2_X2 U6716 ( .A1(n5561), .A2(n5560), .ZN(n5590) );
  INV_X1 U6717 ( .A(n5590), .ZN(n5108) );
  AND2_X1 U6718 ( .A1(P1_REG3_REG_27__SCAN_IN), .A2(P1_REG3_REG_28__SCAN_IN), 
        .ZN(n5107) );
  NAND2_X1 U6719 ( .A1(n5108), .A2(n5107), .ZN(n9279) );
  OR2_X1 U6720 ( .A1(n9279), .A2(n5535), .ZN(n5115) );
  INV_X1 U6721 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n5112) );
  NAND2_X1 U6722 ( .A1(n5592), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n5111) );
  NAND2_X1 U6723 ( .A1(n5591), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n5110) );
  OAI211_X1 U6724 ( .C1(n5112), .C2(n5596), .A(n5111), .B(n5110), .ZN(n5113)
         );
  INV_X1 U6725 ( .A(n5113), .ZN(n5114) );
  NAND2_X1 U6726 ( .A1(n9511), .A2(n9287), .ZN(n5734) );
  NAND2_X1 U6727 ( .A1(n9788), .A2(n5586), .ZN(n5119) );
  NAND2_X1 U6728 ( .A1(n5164), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n5118) );
  INV_X1 U6729 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n9008) );
  INV_X1 U6730 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n5120) );
  OAI21_X1 U6731 ( .B1(n5590), .B2(n9008), .A(n5120), .ZN(n5121) );
  NAND2_X1 U6732 ( .A1(n5121), .A2(n9279), .ZN(n9294) );
  INV_X1 U6733 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n9293) );
  NAND2_X1 U6734 ( .A1(n5564), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n5123) );
  NAND2_X1 U6735 ( .A1(n5591), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5122) );
  OAI211_X1 U6736 ( .C1(n5568), .C2(n9293), .A(n5123), .B(n5122), .ZN(n5124)
         );
  INV_X1 U6737 ( .A(n5124), .ZN(n5125) );
  NAND2_X1 U6738 ( .A1(n9514), .A2(n9318), .ZN(n5731) );
  AND2_X1 U6739 ( .A1(n5734), .A2(n5731), .ZN(n5127) );
  INV_X1 U6740 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n5128) );
  OR2_X1 U6741 ( .A1(n5256), .A2(n5128), .ZN(n5130) );
  INV_X1 U6742 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U6743 ( .A1(n6728), .A2(n5131), .ZN(n6143) );
  MUX2_X1 U6744 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4251), .Z(n5134) );
  NAND2_X1 U6745 ( .A1(n5155), .A2(n6980), .ZN(n5136) );
  NAND2_X1 U6746 ( .A1(n5563), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n5141) );
  NAND2_X1 U6747 ( .A1(n5564), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5140) );
  INV_X1 U6748 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n5137) );
  OR2_X1 U6749 ( .A1(n5180), .A2(n5137), .ZN(n5139) );
  INV_X1 U6750 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n7344) );
  OR2_X1 U6751 ( .A1(n5256), .A2(n7344), .ZN(n5138) );
  INV_X1 U6752 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n6772) );
  INV_X1 U6753 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n5142) );
  XNOR2_X1 U6754 ( .A(n5143), .B(n5142), .ZN(n6722) );
  MUX2_X2 U6755 ( .A(n6772), .B(n6722), .S(n6663), .Z(n7345) );
  NOR2_X1 U6756 ( .A1(n9161), .A2(n7345), .ZN(n5618) );
  NAND2_X1 U6757 ( .A1(n4640), .A2(n7277), .ZN(n5144) );
  NAND2_X1 U6758 ( .A1(n5563), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n5149) );
  NAND2_X1 U6759 ( .A1(n5564), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n5148) );
  INV_X1 U6760 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6785) );
  OR2_X1 U6761 ( .A1(n5256), .A2(n6785), .ZN(n5147) );
  INV_X1 U6762 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n5145) );
  OR2_X1 U6763 ( .A1(n5180), .A2(n5145), .ZN(n5146) );
  XNOR2_X1 U6764 ( .A(n5151), .B(n5150), .ZN(n5153) );
  MUX2_X1 U6765 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .S(n4251), .Z(n5152) );
  NAND2_X1 U6766 ( .A1(n5164), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5157) );
  OR2_X1 U6767 ( .A1(n5154), .A2(n9779), .ZN(n5166) );
  NAND2_X1 U6768 ( .A1(n5155), .A2(n7087), .ZN(n5156) );
  OAI211_X2 U6769 ( .C1(n5173), .C2(n6741), .A(n5157), .B(n5156), .ZN(n7443)
         );
  XNOR2_X2 U6770 ( .A(n9158), .B(n7443), .ZN(n7436) );
  INV_X1 U6771 ( .A(n9158), .ZN(n8162) );
  NAND2_X1 U6772 ( .A1(n8162), .A2(n7443), .ZN(n5697) );
  NAND2_X1 U6773 ( .A1(n5564), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n5161) );
  OR2_X1 U6774 ( .A1(n5180), .A2(n9957), .ZN(n5160) );
  INV_X1 U6775 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6787) );
  AND4_X2 U6776 ( .A1(n5161), .A2(n5160), .A3(n5159), .A4(n5158), .ZN(n8179)
         );
  INV_X2 U6777 ( .A(n8179), .ZN(n9157) );
  XNOR2_X1 U6778 ( .A(n5163), .B(n5162), .ZN(n6743) );
  NAND2_X1 U6779 ( .A1(n5164), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5169) );
  INV_X1 U6780 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n5165) );
  NAND2_X1 U6781 ( .A1(n5166), .A2(n5165), .ZN(n5167) );
  NAND2_X1 U6782 ( .A1(n5167), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5168) );
  XNOR2_X1 U6783 ( .A(n5168), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6795) );
  NAND2_X1 U6784 ( .A1(n8179), .A2(n7400), .ZN(n5700) );
  AND2_X1 U6785 ( .A1(n5702), .A2(n5700), .ZN(n7314) );
  NAND2_X1 U6786 ( .A1(n5742), .A2(n7314), .ZN(n5170) );
  XNOR2_X1 U6787 ( .A(n5171), .B(n4830), .ZN(n6724) );
  NAND2_X1 U6788 ( .A1(n5164), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6789 ( .A1(n5174), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5175) );
  XNOR2_X1 U6790 ( .A(n5175), .B(P1_IR_REG_4__SCAN_IN), .ZN(n7063) );
  NAND2_X1 U6791 ( .A1(n5155), .A2(n7063), .ZN(n5176) );
  NAND2_X1 U6792 ( .A1(n5564), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n5184) );
  INV_X1 U6793 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n8167) );
  XNOR2_X1 U6794 ( .A(n8167), .B(P1_REG3_REG_4__SCAN_IN), .ZN(n8184) );
  NAND2_X1 U6795 ( .A1(n5563), .A2(n8184), .ZN(n5183) );
  INV_X1 U6796 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n5179) );
  OR2_X1 U6797 ( .A1(n5180), .A2(n5179), .ZN(n5182) );
  INV_X1 U6798 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n7335) );
  OR2_X1 U6799 ( .A1(n5256), .A2(n7335), .ZN(n5181) );
  NAND4_X2 U6800 ( .A1(n5184), .A2(n5183), .A3(n5182), .A4(n5181), .ZN(n9156)
         );
  OR2_X1 U6801 ( .A1(n7555), .A2(n5705), .ZN(n7323) );
  NAND2_X1 U6802 ( .A1(n5564), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n5195) );
  INV_X1 U6803 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n5187) );
  OR2_X1 U6804 ( .A1(n5180), .A2(n5187), .ZN(n5194) );
  INV_X1 U6805 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7431) );
  OR2_X1 U6806 ( .A1(n5256), .A2(n7431), .ZN(n5193) );
  INV_X1 U6807 ( .A(n5188), .ZN(n5211) );
  INV_X1 U6808 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n5190) );
  NAND2_X1 U6809 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n5189) );
  NAND2_X1 U6810 ( .A1(n5190), .A2(n5189), .ZN(n5191) );
  NAND2_X1 U6811 ( .A1(n5211), .A2(n5191), .ZN(n7520) );
  OR2_X1 U6812 ( .A1(n5228), .A2(n7520), .ZN(n5192) );
  INV_X1 U6813 ( .A(n5196), .ZN(n5200) );
  NAND2_X1 U6814 ( .A1(n5197), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5198) );
  MUX2_X1 U6815 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5198), .S(
        P1_IR_REG_5__SCAN_IN), .Z(n5199) );
  NAND2_X1 U6816 ( .A1(n5200), .A2(n5199), .ZN(n6815) );
  INV_X1 U6817 ( .A(n5202), .ZN(n5203) );
  NAND2_X1 U6818 ( .A1(n6726), .A2(n4248), .ZN(n5206) );
  INV_X2 U6819 ( .A(n5435), .ZN(n5587) );
  NAND2_X1 U6820 ( .A1(n5164), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n5205) );
  OAI211_X1 U6821 ( .C1(n6663), .C2(n6815), .A(n5206), .B(n5205), .ZN(n5207)
         );
  NAND2_X1 U6822 ( .A1(n7532), .A2(n5207), .ZN(n5628) );
  INV_X1 U6823 ( .A(n7532), .ZN(n9155) );
  INV_X1 U6824 ( .A(n5621), .ZN(n5626) );
  INV_X1 U6825 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n5208) );
  INV_X1 U6826 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n5209) );
  OR2_X1 U6827 ( .A1(n5180), .A2(n5209), .ZN(n5216) );
  INV_X1 U6828 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n5210) );
  NAND2_X1 U6829 ( .A1(n5211), .A2(n5210), .ZN(n5212) );
  NAND2_X1 U6830 ( .A1(n5226), .A2(n5212), .ZN(n7590) );
  OR2_X1 U6831 ( .A1(n5228), .A2(n7590), .ZN(n5215) );
  INV_X1 U6832 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n5213) );
  NAND2_X1 U6833 ( .A1(n6731), .A2(n5586), .ZN(n5222) );
  OR2_X1 U6834 ( .A1(n5196), .A2(n9779), .ZN(n5220) );
  XNOR2_X1 U6835 ( .A(n5220), .B(P1_IR_REG_6__SCAN_IN), .ZN(n7141) );
  AOI22_X1 U6836 ( .A1(n5164), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5155), .B2(
        n7141), .ZN(n5221) );
  NAND2_X1 U6837 ( .A1(n5222), .A2(n5221), .ZN(n7537) );
  INV_X1 U6838 ( .A(n7519), .ZN(n5830) );
  NAND2_X1 U6839 ( .A1(n5629), .A2(n5622), .ZN(n7529) );
  INV_X1 U6840 ( .A(n7529), .ZN(n7527) );
  NAND2_X1 U6841 ( .A1(n5223), .A2(n7527), .ZN(n5244) );
  NAND2_X1 U6842 ( .A1(n5591), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n5232) );
  INV_X1 U6843 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n6820) );
  OR2_X1 U6844 ( .A1(n5224), .A2(n6820), .ZN(n5231) );
  INV_X1 U6845 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n5225) );
  NAND2_X1 U6846 ( .A1(n5226), .A2(n5225), .ZN(n5227) );
  NAND2_X1 U6847 ( .A1(n5254), .A2(n5227), .ZN(n7483) );
  OR2_X1 U6848 ( .A1(n5228), .A2(n7483), .ZN(n5230) );
  INV_X1 U6849 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7484) );
  OR2_X1 U6850 ( .A1(n5256), .A2(n7484), .ZN(n5229) );
  AND4_X2 U6851 ( .A1(n5232), .A2(n5231), .A3(n5230), .A4(n5229), .ZN(n7589)
         );
  XNOR2_X1 U6852 ( .A(n5234), .B(n5233), .ZN(n6737) );
  INV_X1 U6853 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n5235) );
  AND2_X1 U6854 ( .A1(n5196), .A2(n5235), .ZN(n5263) );
  NOR2_X1 U6855 ( .A1(n5263), .A2(n9779), .ZN(n5236) );
  NAND2_X1 U6856 ( .A1(n5236), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n5239) );
  INV_X1 U6857 ( .A(n5236), .ZN(n5238) );
  INV_X1 U6858 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6859 ( .A1(n5238), .A2(n5237), .ZN(n5249) );
  AOI22_X1 U6860 ( .A1(n5587), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5155), .B2(
        n9163), .ZN(n5240) );
  AND2_X1 U6861 ( .A1(n5706), .A2(n5622), .ZN(n5741) );
  NAND2_X1 U6862 ( .A1(n5842), .A2(n7589), .ZN(n7552) );
  INV_X1 U6863 ( .A(n7552), .ZN(n5241) );
  AOI21_X1 U6864 ( .B1(n5244), .B2(n5741), .A(n5241), .ZN(n5246) );
  AND2_X1 U6865 ( .A1(n7552), .A2(n5629), .ZN(n5243) );
  INV_X1 U6866 ( .A(n5706), .ZN(n5242) );
  AOI21_X1 U6867 ( .B1(n5244), .B2(n5243), .A(n5242), .ZN(n5245) );
  MUX2_X1 U6868 ( .A(n5246), .B(n5245), .S(n7096), .Z(n5261) );
  NAND2_X1 U6869 ( .A1(n6747), .A2(n5586), .ZN(n5252) );
  NAND2_X1 U6870 ( .A1(n5249), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5250) );
  XNOR2_X1 U6871 ( .A(n5250), .B(P1_IR_REG_8__SCAN_IN), .ZN(n6822) );
  AOI22_X1 U6872 ( .A1(n5587), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5155), .B2(
        n6822), .ZN(n5251) );
  NAND2_X2 U6873 ( .A1(n5252), .A2(n5251), .ZN(n9981) );
  NAND2_X1 U6874 ( .A1(n5564), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n5260) );
  INV_X1 U6875 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n5253) );
  OR2_X1 U6876 ( .A1(n5180), .A2(n5253), .ZN(n5259) );
  INV_X1 U6877 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6844) );
  NAND2_X1 U6878 ( .A1(n5254), .A2(n6844), .ZN(n5255) );
  NAND2_X1 U6879 ( .A1(n5268), .A2(n5255), .ZN(n7647) );
  OR2_X1 U6880 ( .A1(n5535), .A2(n7647), .ZN(n5258) );
  INV_X1 U6881 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7561) );
  OR2_X1 U6882 ( .A1(n5256), .A2(n7561), .ZN(n5257) );
  NAND2_X1 U6883 ( .A1(n9981), .A2(n7750), .ZN(n7571) );
  NAND2_X1 U6884 ( .A1(n6756), .A2(n5586), .ZN(n5266) );
  NOR2_X1 U6885 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n5262) );
  NAND2_X1 U6886 ( .A1(n5263), .A2(n5262), .ZN(n5284) );
  NAND2_X1 U6887 ( .A1(n5284), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5264) );
  XNOR2_X1 U6888 ( .A(n5264), .B(P1_IR_REG_9__SCAN_IN), .ZN(n6824) );
  AOI22_X1 U6889 ( .A1(n5587), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5155), .B2(
        n6824), .ZN(n5265) );
  NAND2_X2 U6890 ( .A1(n5266), .A2(n5265), .ZN(n7755) );
  NAND2_X1 U6891 ( .A1(n5591), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n5273) );
  INV_X1 U6892 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7577) );
  OR2_X1 U6893 ( .A1(n5568), .A2(n7577), .ZN(n5272) );
  NAND2_X1 U6894 ( .A1(n5268), .A2(n5267), .ZN(n5269) );
  NAND2_X1 U6895 ( .A1(n5291), .A2(n5269), .ZN(n7753) );
  OR2_X1 U6896 ( .A1(n5535), .A2(n7753), .ZN(n5271) );
  INV_X1 U6897 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n6823) );
  OR2_X1 U6898 ( .A1(n5596), .A2(n6823), .ZN(n5270) );
  OR2_X1 U6899 ( .A1(n7755), .A2(n7920), .ZN(n5297) );
  AND2_X1 U6900 ( .A1(n5297), .A2(n7573), .ZN(n7717) );
  NAND2_X1 U6901 ( .A1(n7755), .A2(n7920), .ZN(n7917) );
  AND2_X1 U6902 ( .A1(n7917), .A2(n7571), .ZN(n5274) );
  MUX2_X1 U6903 ( .A(n7717), .B(n5274), .S(n7096), .Z(n5275) );
  NAND2_X1 U6904 ( .A1(n5277), .A2(n5276), .ZN(n5279) );
  NAND2_X1 U6905 ( .A1(n5279), .A2(n5278), .ZN(n5283) );
  AND2_X1 U6906 ( .A1(n5281), .A2(n5280), .ZN(n5282) );
  NAND2_X1 U6907 ( .A1(n6779), .A2(n5586), .ZN(n5287) );
  NAND2_X1 U6908 ( .A1(n5358), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5318) );
  OR2_X1 U6909 ( .A1(n5318), .A2(n5356), .ZN(n5285) );
  NAND2_X1 U6910 ( .A1(n5318), .A2(n5356), .ZN(n5302) );
  AOI22_X1 U6911 ( .A1(n5587), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5155), .B2(
        n6993), .ZN(n5286) );
  NAND2_X1 U6912 ( .A1(n5564), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n5296) );
  INV_X1 U6913 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n7926) );
  OR2_X1 U6914 ( .A1(n5568), .A2(n7926), .ZN(n5295) );
  INV_X1 U6915 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n5288) );
  OR2_X1 U6916 ( .A1(n5180), .A2(n5288), .ZN(n5294) );
  INV_X1 U6917 ( .A(n5289), .ZN(n5307) );
  NAND2_X1 U6918 ( .A1(n5291), .A2(n5290), .ZN(n5292) );
  NAND2_X1 U6919 ( .A1(n5307), .A2(n5292), .ZN(n7928) );
  OR2_X1 U6920 ( .A1(n5535), .A2(n7928), .ZN(n5293) );
  NAND2_X1 U6921 ( .A1(n7848), .A2(n5297), .ZN(n5712) );
  INV_X1 U6922 ( .A(n7917), .ZN(n5298) );
  MUX2_X1 U6923 ( .A(n5712), .B(n5298), .S(n5608), .Z(n5300) );
  NAND2_X1 U6924 ( .A1(n7709), .A2(n7724), .ZN(n5687) );
  INV_X1 U6925 ( .A(n5687), .ZN(n5299) );
  NAND2_X1 U6926 ( .A1(n6777), .A2(n5586), .ZN(n5305) );
  NAND2_X1 U6927 ( .A1(n5302), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5303) );
  XNOR2_X1 U6928 ( .A(n5303), .B(P1_IR_REG_11__SCAN_IN), .ZN(n9187) );
  AOI22_X1 U6929 ( .A1(n5587), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n9187), .B2(
        n5155), .ZN(n5304) );
  NAND2_X1 U6930 ( .A1(n5591), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n5312) );
  INV_X1 U6931 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7727) );
  OR2_X1 U6932 ( .A1(n5568), .A2(n7727), .ZN(n5311) );
  INV_X1 U6933 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n5306) );
  NAND2_X1 U6934 ( .A1(n5307), .A2(n5306), .ZN(n5308) );
  NAND2_X1 U6935 ( .A1(n5324), .A2(n5308), .ZN(n7868) );
  OR2_X1 U6936 ( .A1(n5535), .A2(n7868), .ZN(n5310) );
  INV_X1 U6937 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7000) );
  OR2_X1 U6938 ( .A1(n5596), .A2(n7000), .ZN(n5309) );
  OR2_X1 U6939 ( .A1(n9606), .A2(n7999), .ZN(n7851) );
  NAND2_X1 U6940 ( .A1(n9606), .A2(n7999), .ZN(n5373) );
  NAND2_X1 U6941 ( .A1(n5332), .A2(n5316), .ZN(n5333) );
  NAND2_X1 U6942 ( .A1(n7008), .A2(n5586), .ZN(n5322) );
  OAI21_X1 U6943 ( .B1(P1_IR_REG_10__SCAN_IN), .B2(P1_IR_REG_11__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n5317) );
  NAND2_X1 U6944 ( .A1(n5318), .A2(n5317), .ZN(n5319) );
  NAND2_X1 U6945 ( .A1(n5319), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n5320) );
  AOI22_X1 U6946 ( .A1(n5587), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n9839), .B2(
        n5155), .ZN(n5321) );
  NAND2_X1 U6947 ( .A1(n5591), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n5329) );
  INV_X1 U6948 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n9188) );
  OR2_X1 U6949 ( .A1(n5596), .A2(n9188), .ZN(n5328) );
  INV_X1 U6950 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n5323) );
  NAND2_X1 U6951 ( .A1(n5324), .A2(n5323), .ZN(n5325) );
  NAND2_X1 U6952 ( .A1(n5342), .A2(n5325), .ZN(n8009) );
  OR2_X1 U6953 ( .A1(n5535), .A2(n8009), .ZN(n5327) );
  INV_X1 U6954 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n8004) );
  OR2_X1 U6955 ( .A1(n5568), .A2(n8004), .ZN(n5326) );
  NAND2_X1 U6956 ( .A1(n9599), .A2(n7893), .ZN(n5617) );
  AND2_X1 U6957 ( .A1(n5617), .A2(n5687), .ZN(n5330) );
  MUX2_X1 U6958 ( .A(n7848), .B(n5330), .S(n7096), .Z(n5331) );
  NAND2_X1 U6959 ( .A1(n7074), .A2(n5586), .ZN(n5340) );
  NAND2_X1 U6960 ( .A1(n5337), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5338) );
  XNOR2_X1 U6961 ( .A(n5338), .B(P1_IR_REG_13__SCAN_IN), .ZN(n9856) );
  AOI22_X1 U6962 ( .A1(n9856), .A2(n5155), .B1(n5587), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n5339) );
  NAND2_X1 U6963 ( .A1(n5592), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5347) );
  INV_X1 U6964 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n9682) );
  OR2_X1 U6965 ( .A1(n5180), .A2(n9682), .ZN(n5346) );
  NAND2_X1 U6966 ( .A1(n5342), .A2(n5341), .ZN(n5343) );
  NAND2_X1 U6967 ( .A1(n5364), .A2(n5343), .ZN(n7908) );
  OR2_X1 U6968 ( .A1(n5535), .A2(n7908), .ZN(n5345) );
  INV_X1 U6969 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n9189) );
  OR2_X1 U6970 ( .A1(n5596), .A2(n9189), .ZN(n5344) );
  OR2_X1 U6971 ( .A1(n9594), .A2(n8125), .ZN(n5616) );
  OR2_X1 U6972 ( .A1(n5314), .A2(n5348), .ZN(n5350) );
  AND2_X1 U6973 ( .A1(n5350), .A2(n5349), .ZN(n5352) );
  XNOR2_X1 U6974 ( .A(n5352), .B(n5351), .ZN(n7015) );
  NAND2_X1 U6975 ( .A1(n7015), .A2(n5586), .ZN(n5361) );
  INV_X1 U6976 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n5355) );
  INV_X1 U6977 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n5354) );
  INV_X1 U6978 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n5353) );
  NAND4_X1 U6979 ( .A1(n5356), .A2(n5355), .A3(n5354), .A4(n5353), .ZN(n5357)
         );
  NAND2_X1 U6980 ( .A1(n5379), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5359) );
  XNOR2_X1 U6981 ( .A(n5359), .B(P1_IR_REG_14__SCAN_IN), .ZN(n9191) );
  AOI22_X1 U6982 ( .A1(n5587), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5155), .B2(
        n9191), .ZN(n5360) );
  NAND2_X1 U6983 ( .A1(n5592), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5369) );
  INV_X1 U6984 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n5362) );
  OR2_X1 U6985 ( .A1(n5180), .A2(n5362), .ZN(n5368) );
  INV_X1 U6986 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n5363) );
  NAND2_X1 U6987 ( .A1(n5364), .A2(n5363), .ZN(n5365) );
  NAND2_X1 U6988 ( .A1(n5386), .A2(n5365), .ZN(n8128) );
  OR2_X1 U6989 ( .A1(n5535), .A2(n8128), .ZN(n5367) );
  INV_X1 U6990 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n9190) );
  OR2_X1 U6991 ( .A1(n5596), .A2(n9190), .ZN(n5366) );
  OR2_X1 U6992 ( .A1(n9590), .A2(n7907), .ZN(n8107) );
  NAND2_X1 U6993 ( .A1(n5616), .A2(n8107), .ZN(n5392) );
  INV_X1 U6994 ( .A(n7851), .ZN(n5370) );
  NAND2_X1 U6995 ( .A1(n5617), .A2(n5370), .ZN(n5371) );
  NAND2_X1 U6996 ( .A1(n5371), .A2(n7854), .ZN(n5372) );
  OR2_X1 U6997 ( .A1(n5392), .A2(n5372), .ZN(n5717) );
  NAND2_X1 U6998 ( .A1(n9590), .A2(n7907), .ZN(n5690) );
  AND2_X1 U6999 ( .A1(n5690), .A2(n5608), .ZN(n5391) );
  NAND2_X1 U7000 ( .A1(n5617), .A2(n5373), .ZN(n5689) );
  NAND2_X1 U7001 ( .A1(n5689), .A2(n7854), .ZN(n5374) );
  NAND2_X1 U7002 ( .A1(n9594), .A2(n8125), .ZN(n7857) );
  NAND3_X1 U7003 ( .A1(n5391), .A2(n5374), .A3(n7857), .ZN(n5375) );
  OAI21_X1 U7004 ( .B1(n5717), .B2(n5608), .A(n5375), .ZN(n5395) );
  NAND2_X1 U7005 ( .A1(n7857), .A2(n5690), .ZN(n5376) );
  NAND2_X1 U7006 ( .A1(n5376), .A2(n8107), .ZN(n5715) );
  XNOR2_X1 U7007 ( .A(n5378), .B(n5377), .ZN(n7090) );
  NAND2_X1 U7008 ( .A1(n7090), .A2(n5586), .ZN(n5382) );
  NOR2_X1 U7009 ( .A1(n5379), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n5399) );
  OR2_X1 U7010 ( .A1(n5399), .A2(n9779), .ZN(n5380) );
  XNOR2_X1 U7011 ( .A(n5380), .B(P1_IR_REG_15__SCAN_IN), .ZN(n9885) );
  AOI22_X1 U7012 ( .A1(n9885), .A2(n5155), .B1(n5587), .B2(
        P2_DATAO_REG_15__SCAN_IN), .ZN(n5381) );
  INV_X1 U7013 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n9717) );
  OR2_X1 U7014 ( .A1(n5568), .A2(n9717), .ZN(n5385) );
  INV_X1 U7015 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n5383) );
  OR2_X1 U7016 ( .A1(n5180), .A2(n5383), .ZN(n5384) );
  AND2_X1 U7017 ( .A1(n5385), .A2(n5384), .ZN(n5390) );
  NAND2_X1 U7018 ( .A1(n5386), .A2(n8115), .ZN(n5387) );
  AND2_X1 U7019 ( .A1(n5404), .A2(n5387), .ZN(n8134) );
  NAND2_X1 U7020 ( .A1(n8134), .A2(n5563), .ZN(n5389) );
  NAND2_X1 U7021 ( .A1(n5564), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n5388) );
  OR2_X1 U7022 ( .A1(n9583), .A2(n9067), .ZN(n5718) );
  NAND2_X1 U7023 ( .A1(n9583), .A2(n9067), .ZN(n8110) );
  NAND2_X1 U7024 ( .A1(n5392), .A2(n5391), .ZN(n5393) );
  OAI211_X1 U7025 ( .C1(n5608), .C2(n5715), .A(n4268), .B(n5393), .ZN(n5394)
         );
  AOI21_X1 U7026 ( .B1(n5396), .B2(n5395), .A(n5394), .ZN(n5430) );
  XNOR2_X1 U7027 ( .A(n5397), .B(n4895), .ZN(n7170) );
  NAND2_X1 U7028 ( .A1(n7170), .A2(n5586), .ZN(n5402) );
  INV_X1 U7029 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n5398) );
  NAND2_X1 U7030 ( .A1(n5399), .A2(n5398), .ZN(n5400) );
  NAND2_X1 U7031 ( .A1(n5400), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5414) );
  XNOR2_X1 U7032 ( .A(n5414), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9185) );
  AOI22_X1 U7033 ( .A1(n9185), .A2(n5155), .B1(n5587), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n5401) );
  INV_X1 U7034 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U7035 ( .A1(n5404), .A2(n5403), .ZN(n5405) );
  NAND2_X1 U7036 ( .A1(n5421), .A2(n5405), .ZN(n9070) );
  OR2_X1 U7037 ( .A1(n9070), .A2(n5535), .ZN(n5408) );
  AOI22_X1 U7038 ( .A1(n5592), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n5591), .B2(
        P1_REG0_REG_16__SCAN_IN), .ZN(n5407) );
  NAND2_X1 U7039 ( .A1(n5564), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5406) );
  INV_X1 U7040 ( .A(n9245), .ZN(n5427) );
  NAND2_X1 U7041 ( .A1(n9244), .A2(n5427), .ZN(n9221) );
  INV_X1 U7042 ( .A(n9221), .ZN(n5410) );
  MUX2_X1 U7043 ( .A(n8110), .B(n5718), .S(n7096), .Z(n5409) );
  NAND2_X1 U7044 ( .A1(n5410), .A2(n5409), .ZN(n5429) );
  XNOR2_X1 U7045 ( .A(n5412), .B(n5411), .ZN(n7217) );
  NAND2_X1 U7046 ( .A1(n7217), .A2(n5586), .ZN(n5420) );
  NAND2_X1 U7047 ( .A1(n5414), .A2(n5413), .ZN(n5415) );
  NAND2_X1 U7048 ( .A1(n5415), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5417) );
  INV_X1 U7049 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n5416) );
  NAND2_X1 U7050 ( .A1(n5417), .A2(n5416), .ZN(n5433) );
  OR2_X1 U7051 ( .A1(n5417), .A2(n5416), .ZN(n5418) );
  AOI22_X1 U7052 ( .A1(n9184), .A2(n5155), .B1(n5587), .B2(
        P2_DATAO_REG_17__SCAN_IN), .ZN(n5419) );
  NAND2_X1 U7053 ( .A1(n5421), .A2(n9730), .ZN(n5422) );
  AND2_X1 U7054 ( .A1(n5439), .A2(n5422), .ZN(n9473) );
  NAND2_X1 U7055 ( .A1(n9473), .A2(n5563), .ZN(n5426) );
  AOI22_X1 U7056 ( .A1(n5564), .A2(P1_REG1_REG_17__SCAN_IN), .B1(n5591), .B2(
        P1_REG0_REG_17__SCAN_IN), .ZN(n5425) );
  INV_X1 U7057 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n5423) );
  OR2_X1 U7058 ( .A1(n5568), .A2(n5423), .ZN(n5424) );
  NAND2_X1 U7059 ( .A1(n9573), .A2(n9125), .ZN(n5446) );
  MUX2_X1 U7060 ( .A(n9244), .B(n5427), .S(n7096), .Z(n5428) );
  OAI211_X1 U7061 ( .C1(n5430), .C2(n5429), .A(n9478), .B(n5428), .ZN(n5449)
         );
  XNOR2_X1 U7062 ( .A(n5432), .B(n5431), .ZN(n7340) );
  NAND2_X1 U7063 ( .A1(n7340), .A2(n5586), .ZN(n5438) );
  NAND2_X1 U7064 ( .A1(n5433), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5434) );
  XNOR2_X1 U7065 ( .A(n5434), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9183) );
  INV_X1 U7066 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9732) );
  NOR2_X1 U7067 ( .A1(n5435), .A2(n9732), .ZN(n5436) );
  AOI21_X1 U7068 ( .B1(n9183), .B2(n5155), .A(n5436), .ZN(n5437) );
  INV_X1 U7069 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n9712) );
  NAND2_X1 U7070 ( .A1(n5439), .A2(n9712), .ZN(n5440) );
  NAND2_X1 U7071 ( .A1(n5455), .A2(n5440), .ZN(n9461) );
  OR2_X1 U7072 ( .A1(n9461), .A2(n5535), .ZN(n5445) );
  INV_X1 U7073 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9462) );
  NAND2_X1 U7074 ( .A1(n5564), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n5442) );
  NAND2_X1 U7075 ( .A1(n5591), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n5441) );
  OAI211_X1 U7076 ( .C1(n5568), .C2(n9462), .A(n5442), .B(n5441), .ZN(n5443)
         );
  INV_X1 U7077 ( .A(n5443), .ZN(n5444) );
  NAND2_X1 U7078 ( .A1(n9568), .A2(n9485), .ZN(n9250) );
  NAND2_X1 U7079 ( .A1(n9250), .A2(n5446), .ZN(n5721) );
  NAND2_X1 U7080 ( .A1(n5615), .A2(n9247), .ZN(n5677) );
  MUX2_X1 U7081 ( .A(n5721), .B(n5677), .S(n7096), .Z(n5447) );
  INV_X1 U7082 ( .A(n5447), .ZN(n5448) );
  NAND2_X1 U7083 ( .A1(n5449), .A2(n5448), .ZN(n5475) );
  XNOR2_X1 U7084 ( .A(n5451), .B(n5450), .ZN(n7385) );
  NAND2_X1 U7085 ( .A1(n7385), .A2(n5586), .ZN(n5453) );
  AOI22_X1 U7086 ( .A1(n5587), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n7285), .B2(
        n5155), .ZN(n5452) );
  INV_X1 U7087 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n5454) );
  NAND2_X1 U7088 ( .A1(n5455), .A2(n5454), .ZN(n5456) );
  NAND2_X1 U7089 ( .A1(n5467), .A2(n5456), .ZN(n9443) );
  OR2_X1 U7090 ( .A1(n9443), .A2(n5535), .ZN(n5462) );
  INV_X1 U7091 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n5459) );
  NAND2_X1 U7092 ( .A1(n5591), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n5458) );
  NAND2_X1 U7093 ( .A1(n5592), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n5457) );
  OAI211_X1 U7094 ( .C1(n5459), .C2(n5596), .A(n5458), .B(n5457), .ZN(n5460)
         );
  INV_X1 U7095 ( .A(n5460), .ZN(n5461) );
  OR2_X1 U7096 ( .A1(n9561), .A2(n9124), .ZN(n5614) );
  NAND2_X1 U7097 ( .A1(n9561), .A2(n9124), .ZN(n9251) );
  XNOR2_X1 U7098 ( .A(n5464), .B(n5463), .ZN(n7506) );
  NAND2_X1 U7099 ( .A1(n7506), .A2(n5586), .ZN(n5466) );
  NAND2_X1 U7100 ( .A1(n5587), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n5465) );
  NAND2_X1 U7101 ( .A1(n5467), .A2(n9101), .ZN(n5468) );
  NAND2_X1 U7102 ( .A1(n5480), .A2(n5468), .ZN(n9423) );
  OR2_X1 U7103 ( .A1(n9423), .A2(n5535), .ZN(n5474) );
  INV_X1 U7104 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n5471) );
  NAND2_X1 U7105 ( .A1(n5592), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U7106 ( .A1(n5591), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n5469) );
  OAI211_X1 U7107 ( .C1(n5471), .C2(n5596), .A(n5470), .B(n5469), .ZN(n5472)
         );
  INV_X1 U7108 ( .A(n5472), .ZN(n5473) );
  INV_X1 U7109 ( .A(n9252), .ZN(n5613) );
  AND2_X1 U7110 ( .A1(n9251), .A2(n9250), .ZN(n5678) );
  AND2_X1 U7111 ( .A1(n9253), .A2(n5614), .ZN(n5679) );
  XNOR2_X1 U7112 ( .A(n5477), .B(n5476), .ZN(n7620) );
  NAND2_X1 U7113 ( .A1(n7620), .A2(n5586), .ZN(n5479) );
  NAND2_X1 U7114 ( .A1(n5587), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n5478) );
  NAND2_X1 U7115 ( .A1(n5480), .A2(n9035), .ZN(n5481) );
  AND2_X1 U7116 ( .A1(n5493), .A2(n5481), .ZN(n9411) );
  NAND2_X1 U7117 ( .A1(n9411), .A2(n5563), .ZN(n5487) );
  INV_X1 U7118 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n5484) );
  NAND2_X1 U7119 ( .A1(n5592), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n5483) );
  NAND2_X1 U7120 ( .A1(n5591), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n5482) );
  OAI211_X1 U7121 ( .C1(n5484), .C2(n5596), .A(n5483), .B(n5482), .ZN(n5485)
         );
  INV_X1 U7122 ( .A(n5485), .ZN(n5486) );
  NAND2_X1 U7123 ( .A1(n5680), .A2(n9253), .ZN(n5488) );
  NAND2_X1 U7124 ( .A1(n9552), .A2(n9113), .ZN(n9255) );
  OAI21_X1 U7125 ( .B1(n4288), .B2(n5488), .A(n9255), .ZN(n5501) );
  XNOR2_X1 U7126 ( .A(n5490), .B(n5489), .ZN(n7743) );
  NAND2_X1 U7127 ( .A1(n7743), .A2(n5586), .ZN(n5492) );
  NAND2_X1 U7128 ( .A1(n5587), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n5491) );
  INV_X1 U7129 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n9112) );
  NAND2_X1 U7130 ( .A1(n5493), .A2(n9112), .ZN(n5494) );
  NAND2_X1 U7131 ( .A1(n5532), .A2(n5494), .ZN(n9391) );
  OR2_X1 U7132 ( .A1(n9391), .A2(n5535), .ZN(n5500) );
  INV_X1 U7133 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n5497) );
  NAND2_X1 U7134 ( .A1(n5592), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n5496) );
  NAND2_X1 U7135 ( .A1(n5591), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n5495) );
  OAI211_X1 U7136 ( .C1(n5497), .C2(n5596), .A(n5496), .B(n5495), .ZN(n5498)
         );
  INV_X1 U7137 ( .A(n5498), .ZN(n5499) );
  NAND2_X1 U7138 ( .A1(n5501), .A2(n9257), .ZN(n5503) );
  NOR2_X1 U7139 ( .A1(n9256), .A2(n7096), .ZN(n5502) );
  NAND2_X1 U7140 ( .A1(n5503), .A2(n5502), .ZN(n5559) );
  NAND2_X1 U7141 ( .A1(n8091), .A2(n5586), .ZN(n5507) );
  NAND2_X1 U7142 ( .A1(n5587), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n5506) );
  INV_X1 U7143 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n5508) );
  NAND2_X1 U7144 ( .A1(n5521), .A2(n5508), .ZN(n5509) );
  NAND2_X1 U7145 ( .A1(n5561), .A2(n5509), .ZN(n9051) );
  INV_X1 U7146 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n9721) );
  NAND2_X1 U7147 ( .A1(n5592), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n5511) );
  NAND2_X1 U7148 ( .A1(n5564), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n5510) );
  OAI211_X1 U7149 ( .C1(n5180), .C2(n9721), .A(n5511), .B(n5510), .ZN(n5512)
         );
  INV_X1 U7150 ( .A(n5512), .ZN(n5513) );
  NAND2_X1 U7151 ( .A1(n9533), .A2(n9140), .ZN(n5643) );
  NAND2_X1 U7152 ( .A1(n7914), .A2(n5586), .ZN(n5518) );
  NAND2_X1 U7153 ( .A1(n5164), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n5517) );
  NAND2_X1 U7154 ( .A1(n5534), .A2(n5519), .ZN(n5520) );
  AND2_X1 U7155 ( .A1(n5521), .A2(n5520), .ZN(n9364) );
  NAND2_X1 U7156 ( .A1(n9364), .A2(n5563), .ZN(n5526) );
  INV_X1 U7157 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n9680) );
  NAND2_X1 U7158 ( .A1(n5592), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n5523) );
  NAND2_X1 U7159 ( .A1(n5564), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n5522) );
  OAI211_X1 U7160 ( .C1(n5180), .C2(n9680), .A(n5523), .B(n5522), .ZN(n5524)
         );
  INV_X1 U7161 ( .A(n5524), .ZN(n5525) );
  NAND2_X1 U7162 ( .A1(n9366), .A2(n9053), .ZN(n9260) );
  NAND2_X1 U7163 ( .A1(n5643), .A2(n9260), .ZN(n5756) );
  XNOR2_X1 U7164 ( .A(n5528), .B(n5527), .ZN(n7782) );
  NAND2_X1 U7165 ( .A1(n7782), .A2(n5586), .ZN(n5530) );
  NAND2_X1 U7166 ( .A1(n5587), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n5529) );
  INV_X1 U7167 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U7168 ( .A1(n5532), .A2(n5531), .ZN(n5533) );
  NAND2_X1 U7169 ( .A1(n5534), .A2(n5533), .ZN(n9015) );
  OR2_X1 U7170 ( .A1(n9015), .A2(n5535), .ZN(n5541) );
  INV_X1 U7171 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U7172 ( .A1(n5591), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U7173 ( .A1(n5592), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n5536) );
  OAI211_X1 U7174 ( .C1(n5538), .C2(n5596), .A(n5537), .B(n5536), .ZN(n5539)
         );
  INV_X1 U7175 ( .A(n5539), .ZN(n5540) );
  NAND2_X1 U7176 ( .A1(n9541), .A2(n9090), .ZN(n9259) );
  INV_X1 U7177 ( .A(n9259), .ZN(n5542) );
  AND2_X1 U7178 ( .A1(n5725), .A2(n5542), .ZN(n5543) );
  NOR2_X1 U7179 ( .A1(n5756), .A2(n5543), .ZN(n5545) );
  INV_X1 U7180 ( .A(n5545), .ZN(n5558) );
  XNOR2_X1 U7181 ( .A(n9541), .B(n9387), .ZN(n9382) );
  AOI21_X1 U7182 ( .B1(n5725), .B2(n9382), .A(n7096), .ZN(n5544) );
  NAND2_X1 U7183 ( .A1(n5545), .A2(n5544), .ZN(n5557) );
  INV_X1 U7184 ( .A(n5680), .ZN(n5548) );
  NAND2_X1 U7185 ( .A1(n5680), .A2(n9252), .ZN(n5546) );
  NAND2_X1 U7186 ( .A1(n5546), .A2(n9255), .ZN(n5547) );
  OR2_X1 U7187 ( .A1(n9256), .A2(n5547), .ZN(n5686) );
  INV_X1 U7188 ( .A(n5686), .ZN(n5685) );
  AND2_X1 U7189 ( .A1(n9257), .A2(n7096), .ZN(n5549) );
  AND4_X1 U7190 ( .A1(n5725), .A2(n5550), .A3(n5549), .A4(n9258), .ZN(n5555)
         );
  NAND3_X1 U7191 ( .A1(n9541), .A2(n9090), .A3(n9053), .ZN(n5553) );
  AOI21_X1 U7192 ( .B1(n9374), .B2(n9387), .A(n5608), .ZN(n5551) );
  OAI21_X1 U7193 ( .B1(n9541), .B2(n9053), .A(n5551), .ZN(n5552) );
  AOI21_X1 U7194 ( .B1(n4757), .B2(n5553), .A(n5552), .ZN(n5554) );
  OAI21_X1 U7195 ( .B1(n5555), .B2(n5554), .A(n9262), .ZN(n5556) );
  OAI211_X1 U7196 ( .C1(n5559), .C2(n5558), .A(n5557), .B(n5556), .ZN(n5580)
         );
  INV_X1 U7197 ( .A(n5580), .ZN(n5583) );
  NAND2_X1 U7198 ( .A1(n5561), .A2(n5560), .ZN(n5562) );
  NAND2_X1 U7199 ( .A1(n9329), .A2(n5563), .ZN(n5571) );
  INV_X1 U7200 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U7201 ( .A1(n5564), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n5566) );
  NAND2_X1 U7202 ( .A1(n5591), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n5565) );
  OAI211_X1 U7203 ( .C1(n5568), .C2(n5567), .A(n5566), .B(n5565), .ZN(n5569)
         );
  INV_X1 U7204 ( .A(n5569), .ZN(n5570) );
  NAND2_X1 U7205 ( .A1(n5587), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n5574) );
  MUX2_X1 U7206 ( .A(n9315), .B(n9527), .S(n5608), .Z(n5582) );
  MUX2_X1 U7207 ( .A(n9262), .B(n5643), .S(n7096), .Z(n5576) );
  NAND2_X1 U7208 ( .A1(n5582), .A2(n5576), .ZN(n5579) );
  OR2_X2 U7209 ( .A1(n9527), .A2(n9315), .ZN(n9239) );
  NOR2_X1 U7210 ( .A1(n5576), .A2(n9239), .ZN(n5578) );
  MUX2_X1 U7211 ( .A(n9315), .B(n9527), .S(n7096), .Z(n5577) );
  OAI22_X1 U7212 ( .A1(n5580), .A2(n5579), .B1(n5578), .B2(n5577), .ZN(n5581)
         );
  OAI21_X1 U7213 ( .B1(n5583), .B2(n5582), .A(n5581), .ZN(n5600) );
  NAND2_X1 U7214 ( .A1(n5587), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n5588) );
  NAND2_X1 U7215 ( .A1(n9307), .A2(n5563), .ZN(n5599) );
  INV_X1 U7216 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U7217 ( .A1(n5591), .A2(P1_REG0_REG_27__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U7218 ( .A1(n5592), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n5593) );
  OAI211_X1 U7219 ( .C1(n5596), .C2(n5595), .A(n5594), .B(n5593), .ZN(n5597)
         );
  INV_X1 U7220 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U7221 ( .A1(n9520), .A2(n9288), .ZN(n5730) );
  NAND2_X1 U7222 ( .A1(n5600), .A2(n9314), .ZN(n5602) );
  MUX2_X1 U7223 ( .A(n9265), .B(n5730), .S(n7096), .Z(n5601) );
  NAND3_X1 U7224 ( .A1(n5602), .A2(n9285), .A3(n5601), .ZN(n5604) );
  MUX2_X1 U7225 ( .A(n5734), .B(n5612), .S(n5608), .Z(n5603) );
  NAND2_X1 U7226 ( .A1(n9268), .A2(n9213), .ZN(n5606) );
  NAND2_X1 U7227 ( .A1(n9217), .A2(n5606), .ZN(n5761) );
  NAND2_X1 U7228 ( .A1(n9496), .A2(n9213), .ZN(n5649) );
  NAND2_X1 U7229 ( .A1(n5649), .A2(n7189), .ZN(n5766) );
  INV_X1 U7230 ( .A(n5649), .ZN(n5738) );
  NAND2_X1 U7231 ( .A1(n7188), .A2(n7189), .ZN(n7194) );
  NOR2_X1 U7232 ( .A1(n5738), .A2(n7194), .ZN(n5672) );
  NAND2_X1 U7233 ( .A1(n5611), .A2(n5610), .ZN(n5674) );
  INV_X1 U7234 ( .A(n9360), .ZN(n9356) );
  NAND2_X1 U7235 ( .A1(n5613), .A2(n9253), .ZN(n9427) );
  NAND2_X1 U7236 ( .A1(n5615), .A2(n9250), .ZN(n9248) );
  NAND2_X1 U7237 ( .A1(n7848), .A2(n5687), .ZN(n7919) );
  XNOR2_X1 U7238 ( .A(n7755), .B(n7920), .ZN(n7574) );
  INV_X1 U7239 ( .A(n5618), .ZN(n5619) );
  INV_X1 U7240 ( .A(n5619), .ZN(n7192) );
  AND2_X1 U7241 ( .A1(n9161), .A2(n7345), .ZN(n5693) );
  NOR2_X1 U7242 ( .A1(n7192), .A2(n5693), .ZN(n7100) );
  NAND4_X1 U7243 ( .A1(n7193), .A2(n7546), .A3(n7100), .A4(n5702), .ZN(n5620)
         );
  INV_X1 U7244 ( .A(n7436), .ZN(n7442) );
  OR2_X1 U7245 ( .A1(n5620), .A2(n7442), .ZN(n5625) );
  NAND2_X1 U7246 ( .A1(n5629), .A2(n5621), .ZN(n5623) );
  INV_X1 U7247 ( .A(n7549), .ZN(n5624) );
  NOR2_X1 U7248 ( .A1(n5625), .A2(n5624), .ZN(n5632) );
  INV_X1 U7249 ( .A(n5700), .ZN(n5627) );
  OAI211_X1 U7250 ( .C1(n5627), .C2(n5705), .A(n5626), .B(n7546), .ZN(n5631)
         );
  INV_X1 U7251 ( .A(n7547), .ZN(n5630) );
  AND2_X1 U7252 ( .A1(n5631), .A2(n5630), .ZN(n5746) );
  NAND4_X1 U7253 ( .A1(n7550), .A2(n7557), .A3(n5632), .A4(n5746), .ZN(n5633)
         );
  NOR3_X1 U7254 ( .A1(n7919), .A2(n7574), .A3(n5633), .ZN(n5634) );
  NAND3_X1 U7255 ( .A1(n7853), .A2(n7850), .A3(n5634), .ZN(n5635) );
  NOR2_X1 U7256 ( .A1(n7890), .A2(n5635), .ZN(n5637) );
  XNOR2_X1 U7257 ( .A(n9590), .B(n7907), .ZN(n8108) );
  INV_X1 U7258 ( .A(n8108), .ZN(n5636) );
  NAND3_X1 U7259 ( .A1(n4268), .A2(n5637), .A3(n5636), .ZN(n5638) );
  NOR2_X1 U7260 ( .A1(n9221), .A2(n5638), .ZN(n5639) );
  NAND4_X1 U7261 ( .A1(n9439), .A2(n9478), .A3(n9249), .A4(n5639), .ZN(n5640)
         );
  OR2_X1 U7262 ( .A1(n9427), .A2(n5640), .ZN(n5641) );
  NAND2_X1 U7263 ( .A1(n5680), .A2(n9255), .ZN(n9405) );
  NOR2_X1 U7264 ( .A1(n5641), .A2(n9405), .ZN(n5642) );
  NAND4_X1 U7265 ( .A1(n9356), .A2(n9396), .A3(n5642), .A4(n9382), .ZN(n5644)
         );
  NOR2_X1 U7266 ( .A1(n5644), .A2(n9340), .ZN(n5645) );
  NAND2_X1 U7267 ( .A1(n9527), .A2(n9315), .ZN(n9240) );
  NAND4_X1 U7268 ( .A1(n9285), .A2(n9314), .A3(n5645), .A4(n9263), .ZN(n5646)
         );
  NOR2_X1 U7269 ( .A1(n9508), .A2(n5646), .ZN(n5648) );
  NAND2_X1 U7270 ( .A1(n9217), .A2(n5647), .ZN(n5736) );
  NAND3_X1 U7271 ( .A1(n5649), .A2(n5648), .A3(n5736), .ZN(n5650) );
  NAND2_X1 U7272 ( .A1(n5651), .A2(n7624), .ZN(n5771) );
  NAND2_X1 U7273 ( .A1(n7188), .A2(n9277), .ZN(n7182) );
  OR2_X1 U7274 ( .A1(n5785), .A2(n7182), .ZN(n7427) );
  NAND2_X1 U7275 ( .A1(n9740), .A2(n5653), .ZN(n5654) );
  OAI21_X1 U7276 ( .B1(n5658), .B2(n5657), .A(P1_IR_REG_31__SCAN_IN), .ZN(
        n5659) );
  MUX2_X1 U7277 ( .A(P1_IR_REG_31__SCAN_IN), .B(n5659), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n5662) );
  NAND2_X1 U7278 ( .A1(n5662), .A2(n5661), .ZN(n8094) );
  NAND2_X1 U7279 ( .A1(n5661), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5663) );
  XNOR2_X1 U7280 ( .A(n5663), .B(P1_IR_REG_26__SCAN_IN), .ZN(n6015) );
  NOR2_X1 U7281 ( .A1(n8094), .A2(n9799), .ZN(n5664) );
  NAND2_X1 U7282 ( .A1(n5665), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5667) );
  INV_X1 U7283 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5666) );
  XNOR2_X1 U7284 ( .A(n5667), .B(n5666), .ZN(n6660) );
  AND2_X1 U7285 ( .A1(n6660), .A2(P1_STATE_REG_SCAN_IN), .ZN(n5668) );
  INV_X1 U7286 ( .A(n7071), .ZN(n7195) );
  NAND2_X1 U7287 ( .A1(n9777), .A2(n7195), .ZN(n5669) );
  OR2_X1 U7288 ( .A1(n7427), .A2(n5669), .ZN(n6045) );
  NOR2_X1 U7289 ( .A1(n6660), .A2(P1_U3084), .ZN(n7758) );
  INV_X1 U7290 ( .A(P1_B_REG_SCAN_IN), .ZN(n9210) );
  AOI21_X1 U7291 ( .B1(n5784), .B2(n7758), .A(n9210), .ZN(n5670) );
  OAI21_X1 U7292 ( .B1(n6045), .B2(n9211), .A(n5670), .ZN(n5775) );
  NAND4_X1 U7293 ( .A1(n5771), .A2(n7285), .A3(n7198), .A4(n5775), .ZN(n5671)
         );
  INV_X1 U7294 ( .A(n5674), .ZN(n5740) );
  INV_X1 U7295 ( .A(n5675), .ZN(n5733) );
  INV_X1 U7296 ( .A(n9265), .ZN(n5676) );
  OR2_X1 U7297 ( .A1(n5733), .A2(n5676), .ZN(n5764) );
  INV_X1 U7298 ( .A(n5677), .ZN(n5682) );
  INV_X1 U7299 ( .A(n5678), .ZN(n5681) );
  OAI211_X1 U7300 ( .C1(n5682), .C2(n5681), .A(n5680), .B(n5679), .ZN(n5684)
         );
  INV_X1 U7301 ( .A(n9257), .ZN(n5683) );
  AOI21_X1 U7302 ( .B1(n5685), .B2(n5684), .A(n5683), .ZN(n5753) );
  NOR2_X1 U7303 ( .A1(n5686), .A2(n4873), .ZN(n5751) );
  NAND2_X1 U7304 ( .A1(n5687), .A2(n7917), .ZN(n7719) );
  NAND2_X1 U7305 ( .A1(n7719), .A2(n7848), .ZN(n7849) );
  INV_X1 U7306 ( .A(n7849), .ZN(n5688) );
  NOR2_X1 U7307 ( .A1(n5689), .A2(n5688), .ZN(n5710) );
  AND3_X1 U7308 ( .A1(n5690), .A2(n7571), .A3(n7552), .ZN(n5691) );
  NAND4_X1 U7309 ( .A1(n5710), .A2(n5691), .A3(n8110), .A4(n7857), .ZN(n5692)
         );
  OR3_X1 U7310 ( .A1(n5721), .A2(n9245), .A3(n5692), .ZN(n5749) );
  INV_X1 U7311 ( .A(n5693), .ZN(n5696) );
  INV_X1 U7312 ( .A(n7277), .ZN(n7130) );
  NAND2_X1 U7313 ( .A1(n9160), .A2(n7130), .ZN(n5695) );
  NAND3_X1 U7314 ( .A1(n5696), .A2(n7189), .A3(n5695), .ZN(n5698) );
  NAND2_X1 U7315 ( .A1(n5698), .A2(n5697), .ZN(n5699) );
  OAI22_X1 U7316 ( .A1(n7437), .A2(n5699), .B1(n8162), .B2(n7443), .ZN(n5701)
         );
  AND2_X1 U7317 ( .A1(n5701), .A2(n5700), .ZN(n5709) );
  AND2_X1 U7318 ( .A1(n5702), .A2(n7546), .ZN(n5703) );
  AND2_X1 U7319 ( .A1(n5706), .A2(n5703), .ZN(n5704) );
  AND2_X1 U7320 ( .A1(n5704), .A2(n7549), .ZN(n5743) );
  INV_X1 U7321 ( .A(n5743), .ZN(n5708) );
  NAND2_X1 U7322 ( .A1(n7549), .A2(n5706), .ZN(n5707) );
  OAI22_X1 U7323 ( .A1(n5709), .A2(n5708), .B1(n7553), .B2(n5707), .ZN(n5722)
         );
  INV_X1 U7324 ( .A(n5710), .ZN(n5714) );
  INV_X1 U7325 ( .A(n7573), .ZN(n5711) );
  NOR2_X1 U7326 ( .A1(n5712), .A2(n5711), .ZN(n5713) );
  NOR2_X1 U7327 ( .A1(n5714), .A2(n5713), .ZN(n5716) );
  OAI211_X1 U7328 ( .C1(n5717), .C2(n5716), .A(n8110), .B(n5715), .ZN(n5719)
         );
  AND3_X1 U7329 ( .A1(n5719), .A2(n5718), .A3(n9244), .ZN(n5720) );
  OR3_X1 U7330 ( .A1(n5721), .A2(n9245), .A3(n5720), .ZN(n5747) );
  OAI21_X1 U7331 ( .B1(n5749), .B2(n5722), .A(n5747), .ZN(n5723) );
  NAND2_X1 U7332 ( .A1(n5751), .A2(n5723), .ZN(n5724) );
  NAND2_X1 U7333 ( .A1(n5753), .A2(n5724), .ZN(n5726) );
  NAND2_X1 U7334 ( .A1(n5725), .A2(n9258), .ZN(n5754) );
  AOI21_X1 U7335 ( .B1(n5726), .B2(n9259), .A(n5754), .ZN(n5727) );
  OAI21_X1 U7336 ( .B1(n5727), .B2(n5756), .A(n9262), .ZN(n5728) );
  INV_X1 U7337 ( .A(n9315), .ZN(n9346) );
  NAND2_X1 U7338 ( .A1(n9527), .A2(n9346), .ZN(n9312) );
  NAND2_X1 U7339 ( .A1(n5728), .A2(n9312), .ZN(n5729) );
  OR2_X1 U7340 ( .A1(n9527), .A2(n9346), .ZN(n5759) );
  NAND2_X1 U7341 ( .A1(n5729), .A2(n5759), .ZN(n5737) );
  AND2_X1 U7342 ( .A1(n5731), .A2(n5730), .ZN(n5732) );
  OR2_X1 U7343 ( .A1(n5733), .A2(n5732), .ZN(n5735) );
  OAI211_X1 U7344 ( .C1(n5764), .C2(n5737), .A(n5762), .B(n5736), .ZN(n5739)
         );
  AOI21_X1 U7345 ( .B1(n5740), .B2(n5739), .A(n5738), .ZN(n5774) );
  NAND3_X1 U7346 ( .A1(n5774), .A2(n6051), .A3(n5775), .ZN(n5780) );
  INV_X1 U7347 ( .A(n5741), .ZN(n5745) );
  NAND2_X1 U7348 ( .A1(n7392), .A2(n5743), .ZN(n5744) );
  OAI21_X1 U7349 ( .B1(n5746), .B2(n5745), .A(n5744), .ZN(n5748) );
  OAI21_X1 U7350 ( .B1(n5749), .B2(n5748), .A(n5747), .ZN(n5750) );
  NAND2_X1 U7351 ( .A1(n5751), .A2(n5750), .ZN(n5752) );
  NAND2_X1 U7352 ( .A1(n5753), .A2(n5752), .ZN(n5755) );
  AOI21_X1 U7353 ( .B1(n5755), .B2(n9259), .A(n5754), .ZN(n5757) );
  OAI21_X1 U7354 ( .B1(n5757), .B2(n5756), .A(n9262), .ZN(n5758) );
  NAND2_X1 U7355 ( .A1(n5758), .A2(n9312), .ZN(n5760) );
  NAND2_X1 U7356 ( .A1(n5760), .A2(n5759), .ZN(n5763) );
  OAI211_X1 U7357 ( .C1(n5764), .C2(n5763), .A(n5762), .B(n5761), .ZN(n5765)
         );
  INV_X1 U7358 ( .A(n5765), .ZN(n5768) );
  INV_X1 U7359 ( .A(n5766), .ZN(n5767) );
  OAI21_X1 U7360 ( .B1(n5769), .B2(n5768), .A(n5767), .ZN(n5770) );
  NAND2_X1 U7361 ( .A1(n5771), .A2(n5770), .ZN(n5772) );
  NAND4_X1 U7362 ( .A1(n5772), .A2(n7198), .A3(n9277), .A4(n5775), .ZN(n5779)
         );
  INV_X1 U7363 ( .A(n7758), .ZN(n5773) );
  NAND2_X1 U7364 ( .A1(n5775), .A2(n5773), .ZN(n5778) );
  INV_X1 U7365 ( .A(n5774), .ZN(n5776) );
  NAND4_X1 U7366 ( .A1(n5776), .A2(n7285), .A3(n5775), .A4(n7642), .ZN(n5777)
         );
  NAND4_X1 U7367 ( .A1(n5780), .A2(n5779), .A3(n5778), .A4(n5777), .ZN(n5781)
         );
  AOI21_X1 U7368 ( .B1(n4899), .B2(n5782), .A(n5781), .ZN(P1_U3240) );
  AND2_X2 U7369 ( .A1(n7278), .A2(n5783), .ZN(n5802) );
  INV_X1 U7370 ( .A(n7278), .ZN(n5785) );
  NAND2_X1 U7371 ( .A1(n5784), .A2(n6051), .ZN(n7183) );
  OR2_X4 U7372 ( .A1(n5787), .A2(n5786), .ZN(n6003) );
  OAI22_X1 U7373 ( .A1(n9352), .A2(n5970), .B1(n9140), .B2(n6003), .ZN(n5988)
         );
  INV_X1 U7374 ( .A(n5988), .ZN(n5995) );
  OR2_X2 U7375 ( .A1(n5787), .A2(n7278), .ZN(n5971) );
  INV_X4 U7376 ( .A(n5971), .ZN(n6036) );
  NAND2_X1 U7377 ( .A1(n9533), .A2(n6036), .ZN(n5789) );
  NAND2_X1 U7378 ( .A1(n9358), .A2(n5802), .ZN(n5788) );
  NAND2_X1 U7379 ( .A1(n5789), .A2(n5788), .ZN(n5790) );
  XNOR2_X1 U7380 ( .A(n5790), .B(n7426), .ZN(n5989) );
  INV_X1 U7381 ( .A(n5989), .ZN(n5994) );
  INV_X1 U7382 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n6765) );
  OAI22_X1 U7383 ( .A1(n7345), .A2(n5971), .B1(n6765), .B2(n5783), .ZN(n5791)
         );
  INV_X1 U7384 ( .A(n5791), .ZN(n5793) );
  NAND2_X1 U7385 ( .A1(n9161), .A2(n5802), .ZN(n5792) );
  NAND2_X1 U7386 ( .A1(n5793), .A2(n5792), .ZN(n7066) );
  NAND2_X1 U7387 ( .A1(n6040), .A2(n9161), .ZN(n5797) );
  OAI22_X1 U7388 ( .A1(n7345), .A2(n5970), .B1(n6772), .B2(n5783), .ZN(n5795)
         );
  INV_X1 U7389 ( .A(n5795), .ZN(n5796) );
  NAND2_X1 U7390 ( .A1(n6036), .A2(n7277), .ZN(n5800) );
  NAND2_X1 U7391 ( .A1(n9160), .A2(n5802), .ZN(n5799) );
  NAND2_X1 U7392 ( .A1(n5800), .A2(n5799), .ZN(n5801) );
  XNOR2_X1 U7393 ( .A(n5801), .B(n7426), .ZN(n5804) );
  XNOR2_X1 U7394 ( .A(n5806), .B(n5804), .ZN(n7120) );
  CLKBUF_X3 U7395 ( .A(n5802), .Z(n6041) );
  AND2_X1 U7396 ( .A1(n7277), .A2(n6041), .ZN(n5803) );
  AOI21_X1 U7397 ( .B1(n6040), .B2(n9160), .A(n5803), .ZN(n7122) );
  NAND2_X1 U7398 ( .A1(n7120), .A2(n7122), .ZN(n7121) );
  INV_X1 U7399 ( .A(n5804), .ZN(n5805) );
  NAND2_X1 U7400 ( .A1(n5806), .A2(n5805), .ZN(n5807) );
  NAND2_X1 U7401 ( .A1(n7121), .A2(n5807), .ZN(n7164) );
  NAND2_X1 U7402 ( .A1(n9158), .A2(n5802), .ZN(n5809) );
  NAND2_X1 U7403 ( .A1(n6036), .A2(n7443), .ZN(n5808) );
  NAND2_X1 U7404 ( .A1(n5809), .A2(n5808), .ZN(n5810) );
  XNOR2_X1 U7405 ( .A(n5810), .B(n7426), .ZN(n5812) );
  AND2_X1 U7406 ( .A1(n7443), .A2(n6041), .ZN(n5811) );
  AOI21_X1 U7407 ( .B1(n6040), .B2(n9158), .A(n5811), .ZN(n5813) );
  XNOR2_X1 U7408 ( .A(n5812), .B(n5813), .ZN(n7163) );
  INV_X1 U7409 ( .A(n5812), .ZN(n5814) );
  NAND2_X1 U7410 ( .A1(n5814), .A2(n5813), .ZN(n5815) );
  OAI22_X1 U7411 ( .A1(n8179), .A2(n5970), .B1(n9952), .B2(n5971), .ZN(n5816)
         );
  XNOR2_X1 U7412 ( .A(n5816), .B(n5794), .ZN(n5817) );
  OAI22_X1 U7413 ( .A1(n8179), .A2(n6003), .B1(n9952), .B2(n5970), .ZN(n5818)
         );
  XNOR2_X1 U7414 ( .A(n5817), .B(n5818), .ZN(n8161) );
  INV_X1 U7415 ( .A(n5817), .ZN(n5819) );
  INV_X1 U7416 ( .A(n8178), .ZN(n5825) );
  NAND2_X1 U7417 ( .A1(n9156), .A2(n5802), .ZN(n5821) );
  OR2_X1 U7418 ( .A1(n9958), .A2(n5971), .ZN(n5820) );
  NAND2_X1 U7419 ( .A1(n5821), .A2(n5820), .ZN(n5822) );
  XNOR2_X1 U7420 ( .A(n5822), .B(n5794), .ZN(n8176) );
  NAND2_X1 U7421 ( .A1(n6040), .A2(n9156), .ZN(n5824) );
  NAND2_X1 U7422 ( .A1(n5186), .A2(n5802), .ZN(n5823) );
  AND2_X1 U7423 ( .A1(n5824), .A2(n5823), .ZN(n8175) );
  INV_X1 U7424 ( .A(n8176), .ZN(n5827) );
  INV_X1 U7425 ( .A(n8175), .ZN(n5826) );
  NAND2_X1 U7426 ( .A1(n5827), .A2(n5826), .ZN(n7509) );
  NAND2_X1 U7427 ( .A1(n7537), .A2(n6036), .ZN(n5828) );
  OAI21_X1 U7428 ( .B1(n7519), .B2(n5970), .A(n5828), .ZN(n5829) );
  AOI22_X1 U7429 ( .A1(n5830), .A2(n6040), .B1(n6041), .B2(n7537), .ZN(n5832)
         );
  NAND2_X1 U7430 ( .A1(n5831), .A2(n5832), .ZN(n7406) );
  INV_X1 U7431 ( .A(n5832), .ZN(n5833) );
  NAND2_X1 U7432 ( .A1(n5834), .A2(n5833), .ZN(n5835) );
  OAI22_X1 U7433 ( .A1(n7532), .A2(n5970), .B1(n9964), .B2(n5971), .ZN(n5836)
         );
  XNOR2_X1 U7434 ( .A(n5836), .B(n7426), .ZN(n7511) );
  OAI22_X1 U7435 ( .A1(n7532), .A2(n6003), .B1(n9964), .B2(n5970), .ZN(n7516)
         );
  AND2_X1 U7436 ( .A1(n7509), .A2(n5838), .ZN(n5837) );
  NAND2_X1 U7437 ( .A1(n7510), .A2(n5837), .ZN(n7405) );
  INV_X1 U7438 ( .A(n5838), .ZN(n5840) );
  OR2_X1 U7439 ( .A1(n7511), .A2(n7516), .ZN(n5839) );
  OR2_X1 U7440 ( .A1(n5840), .A2(n5839), .ZN(n7404) );
  AND2_X1 U7441 ( .A1(n7406), .A2(n7404), .ZN(n5841) );
  NAND2_X1 U7442 ( .A1(n7405), .A2(n5841), .ZN(n5853) );
  NAND2_X1 U7443 ( .A1(n5842), .A2(n6036), .ZN(n5844) );
  NAND2_X1 U7444 ( .A1(n9154), .A2(n5802), .ZN(n5843) );
  NAND2_X1 U7445 ( .A1(n5844), .A2(n5843), .ZN(n5845) );
  XNOR2_X1 U7446 ( .A(n5845), .B(n5794), .ZN(n5848) );
  NAND2_X1 U7447 ( .A1(n5842), .A2(n5802), .ZN(n5847) );
  NAND2_X1 U7448 ( .A1(n9154), .A2(n6040), .ZN(n5846) );
  AND2_X1 U7449 ( .A1(n5847), .A2(n5846), .ZN(n5849) );
  NAND2_X1 U7450 ( .A1(n5848), .A2(n5849), .ZN(n5854) );
  INV_X1 U7451 ( .A(n5848), .ZN(n5851) );
  INV_X1 U7452 ( .A(n5849), .ZN(n5850) );
  NAND2_X1 U7453 ( .A1(n5851), .A2(n5850), .ZN(n5852) );
  AND2_X1 U7454 ( .A1(n5854), .A2(n5852), .ZN(n7407) );
  NAND2_X1 U7455 ( .A1(n5853), .A2(n7407), .ZN(n7409) );
  NOR2_X1 U7456 ( .A1(n7750), .A2(n6003), .ZN(n5855) );
  AOI21_X1 U7457 ( .B1(n9981), .B2(n6041), .A(n5855), .ZN(n5859) );
  NAND2_X1 U7458 ( .A1(n9981), .A2(n6036), .ZN(n5857) );
  INV_X1 U7459 ( .A(n7750), .ZN(n9153) );
  NAND2_X1 U7460 ( .A1(n9153), .A2(n6041), .ZN(n5856) );
  NAND2_X1 U7461 ( .A1(n5857), .A2(n5856), .ZN(n5858) );
  XNOR2_X1 U7462 ( .A(n5858), .B(n7426), .ZN(n7646) );
  INV_X1 U7463 ( .A(n5859), .ZN(n5860) );
  NAND2_X1 U7464 ( .A1(n7755), .A2(n6036), .ZN(n5862) );
  NAND2_X1 U7465 ( .A1(n9152), .A2(n6041), .ZN(n5861) );
  NAND2_X1 U7466 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  XNOR2_X1 U7467 ( .A(n5863), .B(n5794), .ZN(n5865) );
  NOR2_X1 U7468 ( .A1(n7920), .A2(n6003), .ZN(n5864) );
  AOI21_X1 U7469 ( .B1(n7755), .B2(n6041), .A(n5864), .ZN(n5866) );
  NAND2_X1 U7470 ( .A1(n5865), .A2(n5866), .ZN(n7787) );
  INV_X1 U7471 ( .A(n5865), .ZN(n5868) );
  INV_X1 U7472 ( .A(n5866), .ZN(n5867) );
  NAND2_X1 U7473 ( .A1(n5868), .A2(n5867), .ZN(n5869) );
  NAND2_X1 U7474 ( .A1(n7787), .A2(n5869), .ZN(n7748) );
  INV_X1 U7475 ( .A(n7748), .ZN(n5870) );
  NAND2_X1 U7476 ( .A1(n9606), .A2(n6036), .ZN(n5872) );
  NAND2_X1 U7477 ( .A1(n9150), .A2(n6041), .ZN(n5871) );
  NAND2_X1 U7478 ( .A1(n5872), .A2(n5871), .ZN(n5873) );
  XNOR2_X1 U7479 ( .A(n5873), .B(n5794), .ZN(n7947) );
  NOR2_X1 U7480 ( .A1(n7999), .A2(n6003), .ZN(n5874) );
  AOI21_X1 U7481 ( .B1(n9606), .B2(n6041), .A(n5874), .ZN(n7946) );
  NAND2_X1 U7482 ( .A1(n7709), .A2(n6036), .ZN(n5876) );
  INV_X1 U7483 ( .A(n7724), .ZN(n9151) );
  NAND2_X1 U7484 ( .A1(n9151), .A2(n6041), .ZN(n5875) );
  NAND2_X1 U7485 ( .A1(n5876), .A2(n5875), .ZN(n5877) );
  XNOR2_X1 U7486 ( .A(n5877), .B(n5794), .ZN(n7786) );
  NOR2_X1 U7487 ( .A1(n7724), .A2(n6003), .ZN(n5878) );
  AOI21_X1 U7488 ( .B1(n7709), .B2(n6041), .A(n5878), .ZN(n5892) );
  NAND2_X1 U7489 ( .A1(n7786), .A2(n5892), .ZN(n7863) );
  NAND2_X1 U7490 ( .A1(n7863), .A2(n7787), .ZN(n5879) );
  AOI21_X1 U7491 ( .B1(n7947), .B2(n7946), .A(n5879), .ZN(n5880) );
  NAND2_X1 U7492 ( .A1(n9599), .A2(n6036), .ZN(n5882) );
  INV_X1 U7493 ( .A(n7893), .ZN(n9149) );
  NAND2_X1 U7494 ( .A1(n9149), .A2(n6041), .ZN(n5881) );
  NAND2_X1 U7495 ( .A1(n5882), .A2(n5881), .ZN(n5883) );
  XNOR2_X1 U7496 ( .A(n5883), .B(n5794), .ZN(n5885) );
  NOR2_X1 U7497 ( .A1(n7893), .A2(n6003), .ZN(n5884) );
  AOI21_X1 U7498 ( .B1(n9599), .B2(n6041), .A(n5884), .ZN(n5886) );
  NAND2_X1 U7499 ( .A1(n5885), .A2(n5886), .ZN(n5899) );
  INV_X1 U7500 ( .A(n5885), .ZN(n5888) );
  INV_X1 U7501 ( .A(n5886), .ZN(n5887) );
  NAND2_X1 U7502 ( .A1(n5888), .A2(n5887), .ZN(n5889) );
  NAND2_X1 U7503 ( .A1(n5899), .A2(n5889), .ZN(n7950) );
  INV_X1 U7504 ( .A(n7947), .ZN(n5891) );
  OAI21_X1 U7505 ( .B1(n7786), .B2(n5892), .A(n7946), .ZN(n5890) );
  NAND2_X1 U7506 ( .A1(n5891), .A2(n5890), .ZN(n5895) );
  INV_X1 U7507 ( .A(n7786), .ZN(n5893) );
  INV_X1 U7508 ( .A(n7946), .ZN(n7862) );
  INV_X1 U7509 ( .A(n5892), .ZN(n7785) );
  NAND3_X1 U7510 ( .A1(n5893), .A2(n7862), .A3(n7785), .ZN(n5894) );
  NAND2_X1 U7511 ( .A1(n5895), .A2(n5894), .ZN(n5896) );
  NOR2_X1 U7512 ( .A1(n7950), .A2(n5896), .ZN(n5897) );
  NAND2_X1 U7513 ( .A1(n9594), .A2(n6036), .ZN(n5901) );
  INV_X1 U7514 ( .A(n8125), .ZN(n9148) );
  NAND2_X1 U7515 ( .A1(n9148), .A2(n6041), .ZN(n5900) );
  NAND2_X1 U7516 ( .A1(n5901), .A2(n5900), .ZN(n5902) );
  XNOR2_X1 U7517 ( .A(n5902), .B(n7426), .ZN(n5904) );
  NOR2_X1 U7518 ( .A1(n8125), .A2(n6003), .ZN(n5903) );
  AOI21_X1 U7519 ( .B1(n9594), .B2(n6041), .A(n5903), .ZN(n5905) );
  XNOR2_X1 U7520 ( .A(n5904), .B(n5905), .ZN(n7905) );
  INV_X1 U7521 ( .A(n5904), .ZN(n5906) );
  NAND2_X1 U7522 ( .A1(n5906), .A2(n5905), .ZN(n5907) );
  NAND2_X1 U7523 ( .A1(n9590), .A2(n6036), .ZN(n5909) );
  NAND2_X1 U7524 ( .A1(n9147), .A2(n6041), .ZN(n5908) );
  NAND2_X1 U7525 ( .A1(n5909), .A2(n5908), .ZN(n5910) );
  XNOR2_X1 U7526 ( .A(n5910), .B(n5794), .ZN(n5913) );
  NAND2_X1 U7527 ( .A1(n5914), .A2(n5913), .ZN(n8121) );
  NAND2_X1 U7528 ( .A1(n9590), .A2(n6041), .ZN(n5912) );
  NAND2_X1 U7529 ( .A1(n9147), .A2(n6040), .ZN(n5911) );
  NAND2_X1 U7530 ( .A1(n5912), .A2(n5911), .ZN(n8124) );
  NOR2_X1 U7531 ( .A1(n9067), .A2(n6003), .ZN(n5916) );
  AOI21_X1 U7532 ( .B1(n9583), .B2(n6041), .A(n5916), .ZN(n9061) );
  NAND2_X1 U7533 ( .A1(n9583), .A2(n6036), .ZN(n5918) );
  INV_X1 U7534 ( .A(n9067), .ZN(n9146) );
  NAND2_X1 U7535 ( .A1(n9146), .A2(n6041), .ZN(n5917) );
  NAND2_X1 U7536 ( .A1(n5918), .A2(n5917), .ZN(n5919) );
  XNOR2_X1 U7537 ( .A(n5919), .B(n5794), .ZN(n9059) );
  NAND2_X1 U7538 ( .A1(n9580), .A2(n6036), .ZN(n5921) );
  NAND2_X1 U7539 ( .A1(n9223), .A2(n6041), .ZN(n5920) );
  NAND2_X1 U7540 ( .A1(n5921), .A2(n5920), .ZN(n5922) );
  XNOR2_X1 U7541 ( .A(n5922), .B(n7426), .ZN(n5925) );
  NAND2_X1 U7542 ( .A1(n9580), .A2(n6041), .ZN(n5924) );
  NAND2_X1 U7543 ( .A1(n9223), .A2(n6040), .ZN(n5923) );
  NAND2_X1 U7544 ( .A1(n5924), .A2(n5923), .ZN(n5926) );
  NAND2_X1 U7545 ( .A1(n5925), .A2(n5926), .ZN(n9063) );
  OAI21_X1 U7546 ( .B1(n9061), .B2(n9059), .A(n9063), .ZN(n5930) );
  INV_X1 U7547 ( .A(n5925), .ZN(n5928) );
  INV_X1 U7548 ( .A(n5926), .ZN(n5927) );
  NAND2_X1 U7549 ( .A1(n5928), .A2(n5927), .ZN(n9074) );
  NAND3_X1 U7550 ( .A1(n9063), .A2(n9061), .A3(n9059), .ZN(n5929) );
  NAND2_X1 U7551 ( .A1(n9573), .A2(n6036), .ZN(n5932) );
  OR2_X1 U7552 ( .A1(n9125), .A2(n5970), .ZN(n5931) );
  NAND2_X1 U7553 ( .A1(n5932), .A2(n5931), .ZN(n5933) );
  XNOR2_X1 U7554 ( .A(n5933), .B(n7426), .ZN(n5935) );
  NOR2_X1 U7555 ( .A1(n9125), .A2(n6003), .ZN(n5934) );
  AOI21_X1 U7556 ( .B1(n9573), .B2(n6041), .A(n5934), .ZN(n5936) );
  XNOR2_X1 U7557 ( .A(n5935), .B(n5936), .ZN(n9075) );
  INV_X1 U7558 ( .A(n5935), .ZN(n5937) );
  NAND2_X1 U7559 ( .A1(n5937), .A2(n5936), .ZN(n5938) );
  NAND2_X1 U7560 ( .A1(n9561), .A2(n6036), .ZN(n5940) );
  OR2_X1 U7561 ( .A1(n9124), .A2(n5970), .ZN(n5939) );
  NAND2_X1 U7562 ( .A1(n5940), .A2(n5939), .ZN(n5941) );
  XNOR2_X1 U7563 ( .A(n5941), .B(n7426), .ZN(n5949) );
  NAND2_X1 U7564 ( .A1(n9561), .A2(n6041), .ZN(n5943) );
  OR2_X1 U7565 ( .A1(n9124), .A2(n6003), .ZN(n5942) );
  NAND2_X1 U7566 ( .A1(n5943), .A2(n5942), .ZN(n5950) );
  NAND2_X1 U7567 ( .A1(n5949), .A2(n5950), .ZN(n9024) );
  NAND2_X1 U7568 ( .A1(n9568), .A2(n6036), .ZN(n5945) );
  INV_X1 U7569 ( .A(n9485), .ZN(n9441) );
  NAND2_X1 U7570 ( .A1(n9441), .A2(n6041), .ZN(n5944) );
  NAND2_X1 U7571 ( .A1(n5945), .A2(n5944), .ZN(n5946) );
  XNOR2_X1 U7572 ( .A(n5946), .B(n5794), .ZN(n9022) );
  NOR2_X1 U7573 ( .A1(n9485), .A2(n6003), .ZN(n5947) );
  AOI21_X1 U7574 ( .B1(n9568), .B2(n6041), .A(n5947), .ZN(n9119) );
  NAND3_X1 U7575 ( .A1(n9024), .A2(n9022), .A3(n9119), .ZN(n5953) );
  INV_X1 U7576 ( .A(n5949), .ZN(n5952) );
  INV_X1 U7577 ( .A(n5950), .ZN(n5951) );
  NAND2_X1 U7578 ( .A1(n5952), .A2(n5951), .ZN(n9094) );
  NAND2_X1 U7579 ( .A1(n9556), .A2(n6036), .ZN(n5955) );
  NAND2_X1 U7580 ( .A1(n9440), .A2(n6041), .ZN(n5954) );
  NAND2_X1 U7581 ( .A1(n5955), .A2(n5954), .ZN(n5956) );
  XNOR2_X1 U7582 ( .A(n5956), .B(n5794), .ZN(n5959) );
  INV_X1 U7583 ( .A(n5959), .ZN(n5961) );
  NOR2_X1 U7584 ( .A1(n9036), .A2(n6003), .ZN(n5957) );
  AOI21_X1 U7585 ( .B1(n9556), .B2(n6041), .A(n5957), .ZN(n5958) );
  INV_X1 U7586 ( .A(n5958), .ZN(n5960) );
  AND2_X1 U7587 ( .A1(n5959), .A2(n5958), .ZN(n5963) );
  AOI21_X1 U7588 ( .B1(n5961), .B2(n5960), .A(n5963), .ZN(n9095) );
  INV_X1 U7589 ( .A(n5963), .ZN(n5964) );
  OAI22_X1 U7590 ( .A1(n9414), .A2(n5970), .B1(n9113), .B2(n6003), .ZN(n5968)
         );
  NAND2_X1 U7591 ( .A1(n9552), .A2(n6036), .ZN(n5966) );
  NAND2_X1 U7592 ( .A1(n9419), .A2(n6041), .ZN(n5965) );
  NAND2_X1 U7593 ( .A1(n5966), .A2(n5965), .ZN(n5967) );
  XNOR2_X1 U7594 ( .A(n5967), .B(n7426), .ZN(n5969) );
  XOR2_X1 U7595 ( .A(n5968), .B(n5969), .Z(n9033) );
  AOI22_X1 U7596 ( .A1(n9546), .A2(n6041), .B1(n6040), .B2(n9402), .ZN(n5973)
         );
  NAND2_X1 U7597 ( .A1(n5974), .A2(n5973), .ZN(n9107) );
  OAI22_X1 U7598 ( .A1(n9394), .A2(n5971), .B1(n9038), .B2(n5970), .ZN(n5972)
         );
  XNOR2_X1 U7599 ( .A(n5972), .B(n7426), .ZN(n9109) );
  INV_X1 U7600 ( .A(n9013), .ZN(n5993) );
  NAND2_X1 U7601 ( .A1(n9366), .A2(n6036), .ZN(n5976) );
  NAND2_X1 U7602 ( .A1(n9374), .A2(n5802), .ZN(n5975) );
  NAND2_X1 U7603 ( .A1(n5976), .A2(n5975), .ZN(n5977) );
  XNOR2_X1 U7604 ( .A(n5977), .B(n5794), .ZN(n5985) );
  NOR2_X1 U7605 ( .A1(n9053), .A2(n6003), .ZN(n5978) );
  AOI21_X1 U7606 ( .B1(n9366), .B2(n6041), .A(n5978), .ZN(n5984) );
  NAND2_X1 U7607 ( .A1(n9541), .A2(n6036), .ZN(n5980) );
  NAND2_X1 U7608 ( .A1(n9387), .A2(n6041), .ZN(n5979) );
  NAND2_X1 U7609 ( .A1(n5980), .A2(n5979), .ZN(n5981) );
  XNOR2_X1 U7610 ( .A(n5981), .B(n5794), .ZN(n9012) );
  NOR2_X1 U7611 ( .A1(n9090), .A2(n6003), .ZN(n5982) );
  AOI21_X1 U7612 ( .B1(n9541), .B2(n6041), .A(n5982), .ZN(n9043) );
  AND2_X1 U7613 ( .A1(n9012), .A2(n9043), .ZN(n5983) );
  OR2_X1 U7614 ( .A1(n5985), .A2(n5984), .ZN(n9046) );
  OAI21_X1 U7615 ( .B1(n9012), .B2(n9043), .A(n9046), .ZN(n5987) );
  XNOR2_X1 U7616 ( .A(n5989), .B(n5988), .ZN(n9048) );
  AOI21_X2 U7617 ( .B1(n5993), .B2(n5992), .A(n5991), .ZN(n9050) );
  NAND2_X1 U7618 ( .A1(n9527), .A2(n6036), .ZN(n5997) );
  NAND2_X1 U7619 ( .A1(n9315), .A2(n5802), .ZN(n5996) );
  NAND2_X1 U7620 ( .A1(n5997), .A2(n5996), .ZN(n5998) );
  XNOR2_X1 U7621 ( .A(n5998), .B(n7426), .ZN(n6011) );
  AND2_X1 U7622 ( .A1(n9315), .A2(n6040), .ZN(n5999) );
  AOI21_X1 U7623 ( .B1(n9527), .B2(n6041), .A(n5999), .ZN(n6009) );
  XNOR2_X1 U7624 ( .A(n6011), .B(n6009), .ZN(n9136) );
  NAND2_X1 U7625 ( .A1(n9520), .A2(n6036), .ZN(n6001) );
  NAND2_X1 U7626 ( .A1(n9322), .A2(n5802), .ZN(n6000) );
  NAND2_X1 U7627 ( .A1(n6001), .A2(n6000), .ZN(n6002) );
  XNOR2_X1 U7628 ( .A(n6002), .B(n5794), .ZN(n6006) );
  INV_X1 U7629 ( .A(n6006), .ZN(n6008) );
  NOR2_X1 U7630 ( .A1(n9288), .A2(n6003), .ZN(n6004) );
  AOI21_X1 U7631 ( .B1(n9520), .B2(n6041), .A(n6004), .ZN(n6005) );
  INV_X1 U7632 ( .A(n6005), .ZN(n6007) );
  AOI21_X1 U7633 ( .B1(n6008), .B2(n6007), .A(n6044), .ZN(n9005) );
  INV_X1 U7634 ( .A(n9005), .ZN(n6012) );
  INV_X1 U7635 ( .A(n6009), .ZN(n6010) );
  NAND2_X1 U7636 ( .A1(n6014), .A2(n9210), .ZN(n6017) );
  NAND3_X1 U7637 ( .A1(n7992), .A2(P1_B_REG_SCAN_IN), .A3(n8094), .ZN(n6016)
         );
  NAND3_X1 U7638 ( .A1(n6017), .A2(n6016), .A3(n6015), .ZN(n9776) );
  NAND2_X1 U7639 ( .A1(n8094), .A2(n9799), .ZN(n6018) );
  NAND2_X1 U7640 ( .A1(n6019), .A2(n6018), .ZN(n7097) );
  NOR4_X1 U7641 ( .A1(P1_D_REG_14__SCAN_IN), .A2(P1_D_REG_15__SCAN_IN), .A3(
        P1_D_REG_17__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6023) );
  NOR4_X1 U7642 ( .A1(P1_D_REG_12__SCAN_IN), .A2(P1_D_REG_9__SCAN_IN), .A3(
        P1_D_REG_10__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n6022) );
  NOR4_X1 U7643 ( .A1(P1_D_REG_24__SCAN_IN), .A2(P1_D_REG_25__SCAN_IN), .A3(
        P1_D_REG_26__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n6021) );
  NOR4_X1 U7644 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_22__SCAN_IN), .A4(P1_D_REG_23__SCAN_IN), .ZN(n6020) );
  AND4_X1 U7645 ( .A1(n6023), .A2(n6022), .A3(n6021), .A4(n6020), .ZN(n6029)
         );
  NOR2_X1 U7646 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .ZN(
        n6027) );
  NOR4_X1 U7647 ( .A1(P1_D_REG_28__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_29__SCAN_IN), .ZN(n6026) );
  NOR4_X1 U7648 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_6__SCAN_IN), .A4(P1_D_REG_7__SCAN_IN), .ZN(n6025) );
  NOR4_X1 U7649 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_20__SCAN_IN), .A3(
        P1_D_REG_2__SCAN_IN), .A4(P1_D_REG_3__SCAN_IN), .ZN(n6024) );
  AND4_X1 U7650 ( .A1(n6027), .A2(n6026), .A3(n6025), .A4(n6024), .ZN(n6028)
         );
  NAND2_X1 U7651 ( .A1(n6029), .A2(n6028), .ZN(n7092) );
  INV_X1 U7652 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6030) );
  NOR2_X1 U7653 ( .A1(n7092), .A2(n6030), .ZN(n6031) );
  OR2_X1 U7654 ( .A1(n9776), .A2(n6031), .ZN(n6032) );
  NAND2_X1 U7655 ( .A1(n7992), .A2(n9799), .ZN(n9778) );
  NAND2_X1 U7656 ( .A1(n6032), .A2(n9778), .ZN(n7203) );
  NOR2_X1 U7657 ( .A1(n7097), .A2(n7203), .ZN(n6049) );
  NAND2_X1 U7658 ( .A1(n5784), .A2(n7624), .ZN(n7329) );
  INV_X1 U7659 ( .A(n7329), .ZN(n6033) );
  INV_X1 U7660 ( .A(n6051), .ZN(n7328) );
  NAND2_X1 U7661 ( .A1(n9777), .A2(n7194), .ZN(n6034) );
  NOR2_X1 U7662 ( .A1(n9607), .A2(n6034), .ZN(n6035) );
  NAND2_X1 U7663 ( .A1(n9514), .A2(n6036), .ZN(n6038) );
  NAND2_X1 U7664 ( .A1(n9271), .A2(n5802), .ZN(n6037) );
  NAND2_X1 U7665 ( .A1(n6038), .A2(n6037), .ZN(n6039) );
  XNOR2_X1 U7666 ( .A(n6039), .B(n5794), .ZN(n6043) );
  AOI22_X1 U7667 ( .A1(n9514), .A2(n6041), .B1(n6040), .B2(n9271), .ZN(n6042)
         );
  NAND3_X1 U7668 ( .A1(n4898), .A2(n6044), .A3(n9134), .ZN(n6062) );
  INV_X1 U7669 ( .A(n6045), .ZN(n6046) );
  NAND2_X1 U7670 ( .A1(n9777), .A2(n7071), .ZN(n6047) );
  NOR2_X1 U7671 ( .A1(n7427), .A2(n6047), .ZN(n6048) );
  INV_X1 U7672 ( .A(n9294), .ZN(n6054) );
  INV_X1 U7673 ( .A(n6049), .ZN(n6050) );
  NAND2_X1 U7674 ( .A1(n6050), .A2(n9982), .ZN(n7124) );
  NOR2_X1 U7675 ( .A1(n7329), .A2(n7642), .ZN(n7333) );
  NAND2_X1 U7676 ( .A1(n6050), .A2(n7333), .ZN(n6058) );
  OR2_X1 U7677 ( .A1(n7194), .A2(n6051), .ZN(n6056) );
  AND3_X1 U7678 ( .A1(n6056), .A2(n5783), .A3(n6660), .ZN(n6052) );
  NAND3_X1 U7679 ( .A1(n7124), .A2(n6058), .A3(n6052), .ZN(n6053) );
  AOI22_X1 U7680 ( .A1(n6054), .A2(n9137), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n6055) );
  OAI21_X1 U7681 ( .B1(n9287), .B2(n9037), .A(n6055), .ZN(n6060) );
  NAND2_X1 U7682 ( .A1(n6056), .A2(n9777), .ZN(n7204) );
  INV_X1 U7683 ( .A(n7204), .ZN(n6057) );
  NAND2_X1 U7684 ( .A1(n6058), .A2(n6057), .ZN(n7166) );
  NOR2_X1 U7685 ( .A1(n9296), .A2(n9145), .ZN(n6059) );
  AOI211_X1 U7686 ( .C1(n9016), .C2(n9322), .A(n6060), .B(n6059), .ZN(n6061)
         );
  INV_X2 U7687 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n6315) );
  INV_X2 U7688 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6104) );
  INV_X2 U7689 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6465) );
  NOR2_X1 U7690 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n6064) );
  NAND3_X1 U7691 ( .A1(n4284), .A2(n6066), .A3(n6065), .ZN(n6448) );
  INV_X1 U7692 ( .A(n6448), .ZN(n6072) );
  NAND4_X1 U7693 ( .A1(n6067), .A2(n6096), .A3(n6453), .A4(n6639), .ZN(n6641)
         );
  NOR2_X2 U7694 ( .A1(n6641), .A2(n4270), .ZN(n6071) );
  NOR2_X4 U7695 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n6156) );
  AND4_X2 U7696 ( .A1(n6156), .A2(n6070), .A3(n6069), .A4(n6068), .ZN(n6216)
         );
  INV_X1 U7697 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n6073) );
  AND2_X1 U7698 ( .A1(n6859), .A2(n6728), .ZN(n6120) );
  NAND2_X1 U7699 ( .A1(n7506), .A2(n6457), .ZN(n6077) );
  NAND2_X1 U7700 ( .A1(n6410), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n6076) );
  INV_X1 U7701 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n7629) );
  INV_X1 U7702 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n8500) );
  INV_X1 U7703 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n6344) );
  INV_X1 U7704 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n8447) );
  NAND2_X1 U7705 ( .A1(n6111), .A2(n8447), .ZN(n6080) );
  AND2_X1 U7706 ( .A1(n6364), .A2(n6080), .ZN(n8723) );
  XNOR2_X2 U7707 ( .A(n6083), .B(P2_IR_REG_30__SCAN_IN), .ZN(n8988) );
  INV_X1 U7708 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n6084) );
  NAND2_X1 U7709 ( .A1(n8723), .A2(n6435), .ZN(n6092) );
  INV_X1 U7710 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9674) );
  OR2_X2 U7711 ( .A1(n8988), .A2(n8993), .ZN(n6150) );
  INV_X4 U7712 ( .A(n6444), .ZN(n6439) );
  NAND2_X1 U7713 ( .A1(n6439), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n6089) );
  NAND2_X1 U7714 ( .A1(n6443), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6088) );
  OAI211_X1 U7715 ( .C1(n9674), .C2(n6273), .A(n6089), .B(n6088), .ZN(n6090)
         );
  INV_X1 U7716 ( .A(n6090), .ZN(n6091) );
  NAND2_X1 U7717 ( .A1(n8898), .A2(n8744), .ZN(n6599) );
  NAND2_X1 U7718 ( .A1(n7385), .A2(n6457), .ZN(n6108) );
  INV_X1 U7719 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6316) );
  NAND4_X1 U7720 ( .A1(n6094), .A2(n6093), .A3(n6316), .A4(n6315), .ZN(n6098)
         );
  NAND4_X1 U7721 ( .A1(n6095), .A2(n6096), .A3(n6239), .A4(n6317), .ZN(n6097)
         );
  NOR2_X1 U7722 ( .A1(n6098), .A2(n6097), .ZN(n6099) );
  INV_X1 U7723 ( .A(n6331), .ZN(n6100) );
  INV_X1 U7724 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6102) );
  NAND2_X1 U7725 ( .A1(n6341), .A2(n6102), .ZN(n6103) );
  NAND2_X1 U7726 ( .A1(n6103), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6105) );
  NAND2_X1 U7727 ( .A1(n6105), .A2(n6104), .ZN(n6463) );
  NAND2_X2 U7728 ( .A1(n6463), .A2(n6106), .ZN(n8637) );
  AOI22_X1 U7729 ( .A1(n7606), .A2(n6861), .B1(n6410), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n6107) );
  INV_X1 U7730 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7731 ( .A1(n6347), .A2(n6109), .ZN(n6110) );
  NAND2_X1 U7732 ( .A1(n6111), .A2(n6110), .ZN(n8749) );
  OR2_X1 U7733 ( .A1(n8749), .A2(n6421), .ZN(n6116) );
  INV_X1 U7734 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n8207) );
  NAND2_X1 U7735 ( .A1(n6439), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7736 ( .A1(n6443), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6112) );
  OAI211_X1 U7737 ( .C1(n8207), .C2(n6273), .A(n6113), .B(n6112), .ZN(n6114)
         );
  INV_X1 U7738 ( .A(n6114), .ZN(n6115) );
  NAND2_X1 U7739 ( .A1(n6116), .A2(n6115), .ZN(n8760) );
  NAND2_X1 U7740 ( .A1(n8755), .A2(n8729), .ZN(n8709) );
  NAND2_X1 U7741 ( .A1(n6599), .A2(n8709), .ZN(n6583) );
  INV_X1 U7742 ( .A(n6583), .ZN(n6360) );
  INV_X1 U7743 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6889) );
  OR2_X1 U7744 ( .A1(n6444), .A2(n6889), .ZN(n6119) );
  INV_X1 U7745 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6869) );
  OR2_X1 U7746 ( .A1(n6273), .A2(n6869), .ZN(n6118) );
  NAND2_X1 U7747 ( .A1(n6166), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n6117) );
  INV_X1 U7748 ( .A(n6743), .ZN(n6121) );
  NAND2_X1 U7749 ( .A1(n6121), .A2(n6120), .ZN(n6125) );
  INV_X1 U7750 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n6122) );
  NAND2_X1 U7751 ( .A1(n6156), .A2(n6122), .ZN(n6159) );
  NAND2_X1 U7752 ( .A1(n6159), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6123) );
  MUX2_X1 U7753 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6123), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n6124) );
  AND2_X1 U7754 ( .A1(n6124), .A2(n6179), .ZN(n6942) );
  NAND2_X1 U7755 ( .A1(n8522), .A2(n10128), .ZN(n6538) );
  INV_X1 U7756 ( .A(n7597), .ZN(n6165) );
  INV_X1 U7757 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7699) );
  INV_X1 U7758 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6886) );
  INV_X1 U7759 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6865) );
  INV_X1 U7760 ( .A(n6146), .ZN(n6134) );
  NAND2_X1 U7761 ( .A1(n6130), .A2(n6120), .ZN(n6132) );
  NAND2_X1 U7762 ( .A1(n6161), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6131) );
  NAND2_X1 U7763 ( .A1(n6166), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n6140) );
  INV_X1 U7764 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n7681) );
  OR2_X1 U7765 ( .A1(n6148), .A2(n7681), .ZN(n6139) );
  INV_X1 U7766 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6135) );
  OR2_X1 U7767 ( .A1(n6149), .A2(n6135), .ZN(n6138) );
  INV_X1 U7768 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n6136) );
  OR2_X1 U7769 ( .A1(n6150), .A2(n6136), .ZN(n6137) );
  NAND4_X2 U7770 ( .A1(n6140), .A2(n6139), .A3(n6138), .A4(n6137), .ZN(n6479)
         );
  NAND2_X1 U7771 ( .A1(n6728), .A2(SI_0_), .ZN(n6142) );
  INV_X1 U7772 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7773 ( .A1(n6142), .A2(n6141), .ZN(n6144) );
  AND2_X1 U7774 ( .A1(n6144), .A2(n6143), .ZN(n9004) );
  MUX2_X1 U7775 ( .A(n9003), .B(n9004), .S(n6859), .Z(n10117) );
  INV_X1 U7776 ( .A(n10117), .ZN(n7688) );
  NAND2_X1 U7777 ( .A1(n6513), .A2(n6477), .ZN(n6522) );
  NAND2_X1 U7778 ( .A1(n6146), .A2(n7689), .ZN(n6516) );
  AND2_X1 U7779 ( .A1(n6522), .A2(n6516), .ZN(n7239) );
  INV_X1 U7780 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n6147) );
  INV_X1 U7781 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6887) );
  INV_X1 U7782 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6864) );
  OR2_X1 U7783 ( .A1(n6150), .A2(n6864), .ZN(n6151) );
  NAND4_X1 U7784 ( .A1(n6154), .A2(n6153), .A3(n6152), .A4(n6151), .ZN(n6673)
         );
  INV_X1 U7785 ( .A(n6741), .ZN(n6155) );
  NAND2_X1 U7786 ( .A1(n6155), .A2(n6120), .ZN(n6164) );
  INV_X1 U7787 ( .A(n6156), .ZN(n6157) );
  NAND2_X1 U7788 ( .A1(n6157), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6158) );
  MUX2_X1 U7789 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6158), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n6160) );
  INV_X1 U7790 ( .A(n6888), .ZN(n8539) );
  NAND2_X1 U7791 ( .A1(n6861), .A2(n8539), .ZN(n6163) );
  NAND2_X1 U7792 ( .A1(n6161), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n6162) );
  OR2_X2 U7793 ( .A1(n6673), .A2(n7241), .ZN(n6524) );
  NAND2_X1 U7794 ( .A1(n6673), .A2(n7241), .ZN(n6515) );
  INV_X1 U7795 ( .A(n7234), .ZN(n7238) );
  NAND2_X1 U7796 ( .A1(n7239), .A2(n7238), .ZN(n7237) );
  NAND2_X1 U7797 ( .A1(n7237), .A2(n6524), .ZN(n8815) );
  NAND2_X1 U7798 ( .A1(n6165), .A2(n8815), .ZN(n8816) );
  NAND2_X1 U7799 ( .A1(n6439), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6175) );
  INV_X1 U7800 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n6167) );
  OR2_X1 U7801 ( .A1(n6388), .A2(n6167), .ZN(n6174) );
  INV_X1 U7802 ( .A(n6168), .ZN(n6188) );
  INV_X1 U7803 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n6170) );
  INV_X1 U7804 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7805 ( .A1(n6170), .A2(n6169), .ZN(n6171) );
  NAND2_X1 U7806 ( .A1(n6188), .A2(n6171), .ZN(n8429) );
  OR2_X1 U7807 ( .A1(n6421), .A2(n8429), .ZN(n6173) );
  INV_X1 U7808 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6872) );
  OR2_X1 U7809 ( .A1(n6273), .A2(n6872), .ZN(n6172) );
  NAND4_X2 U7810 ( .A1(n6175), .A2(n6174), .A3(n6173), .A4(n6172), .ZN(n10019)
         );
  NAND2_X1 U7811 ( .A1(n6724), .A2(n6120), .ZN(n6178) );
  NAND2_X1 U7812 ( .A1(n6179), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6176) );
  AOI22_X1 U7813 ( .A1(n6410), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6861), .B2(
        n6916), .ZN(n6177) );
  NAND2_X1 U7814 ( .A1(n8816), .A2(n6528), .ZN(n7731) );
  NAND2_X1 U7815 ( .A1(n6726), .A2(n6120), .ZN(n6186) );
  INV_X1 U7816 ( .A(n6179), .ZN(n6181) );
  INV_X1 U7817 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7818 ( .A1(n6181), .A2(n6180), .ZN(n6183) );
  NAND2_X1 U7819 ( .A1(n6183), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6182) );
  MUX2_X1 U7820 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6182), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n6184) );
  AOI22_X1 U7821 ( .A1(n6410), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6861), .B2(
        n6928), .ZN(n6185) );
  NAND2_X1 U7822 ( .A1(n6439), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n6194) );
  INV_X1 U7823 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n6187) );
  OR2_X1 U7824 ( .A1(n6388), .A2(n6187), .ZN(n6193) );
  INV_X1 U7825 ( .A(n6199), .ZN(n6190) );
  NAND2_X1 U7826 ( .A1(n6188), .A2(n9676), .ZN(n6189) );
  NAND2_X1 U7827 ( .A1(n6190), .A2(n6189), .ZN(n7734) );
  OR2_X1 U7828 ( .A1(n6421), .A2(n7734), .ZN(n6192) );
  INV_X1 U7829 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n6875) );
  OR2_X1 U7830 ( .A1(n6273), .A2(n6875), .ZN(n6191) );
  NAND2_X1 U7831 ( .A1(n10138), .A2(n8521), .ZN(n6537) );
  NAND2_X1 U7832 ( .A1(n10019), .A2(n7610), .ZN(n7730) );
  AND2_X1 U7833 ( .A1(n6537), .A2(n7730), .ZN(n6539) );
  NAND2_X1 U7834 ( .A1(n7731), .A2(n6539), .ZN(n6195) );
  NAND2_X1 U7835 ( .A1(n6195), .A2(n6529), .ZN(n10078) );
  NAND2_X1 U7836 ( .A1(n6731), .A2(n6457), .ZN(n6198) );
  NAND2_X1 U7837 ( .A1(n6204), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6196) );
  XNOR2_X1 U7838 ( .A(n6196), .B(P2_IR_REG_6__SCAN_IN), .ZN(n6898) );
  AOI22_X1 U7839 ( .A1(n6410), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6898), .B2(
        n6861), .ZN(n6197) );
  NAND2_X1 U7840 ( .A1(n6443), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n6203) );
  INV_X1 U7841 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10092) );
  OR2_X1 U7842 ( .A1(n6444), .A2(n10092), .ZN(n6202) );
  OAI21_X1 U7843 ( .B1(n6199), .B2(P2_REG3_REG_6__SCAN_IN), .A(n6210), .ZN(
        n10091) );
  OR2_X1 U7844 ( .A1(n6421), .A2(n10091), .ZN(n6201) );
  INV_X1 U7845 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n6878) );
  OR2_X1 U7846 ( .A1(n6273), .A2(n6878), .ZN(n6200) );
  NAND2_X1 U7847 ( .A1(n10141), .A2(n7350), .ZN(n6547) );
  NAND2_X1 U7848 ( .A1(n10078), .A2(n10087), .ZN(n10077) );
  NAND2_X1 U7849 ( .A1(n10077), .A2(n6547), .ZN(n10057) );
  NAND2_X1 U7850 ( .A1(n6737), .A2(n6457), .ZN(n6207) );
  OAI21_X1 U7851 ( .B1(n6204), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6205) );
  XNOR2_X1 U7852 ( .A(n6205), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6954) );
  AOI22_X1 U7853 ( .A1(n6954), .A2(n6861), .B1(n6410), .B2(
        P1_DATAO_REG_7__SCAN_IN), .ZN(n6206) );
  NAND2_X1 U7854 ( .A1(n6207), .A2(n6206), .ZN(n10072) );
  NAND2_X1 U7855 ( .A1(n6439), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6215) );
  INV_X1 U7856 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n6208) );
  OR2_X1 U7857 ( .A1(n6388), .A2(n6208), .ZN(n6214) );
  AND2_X1 U7858 ( .A1(n6210), .A2(n6209), .ZN(n6211) );
  OR2_X1 U7859 ( .A1(n6211), .A2(n6221), .ZN(n10070) );
  OR2_X1 U7860 ( .A1(n6421), .A2(n10070), .ZN(n6213) );
  INV_X1 U7861 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6899) );
  OR2_X1 U7862 ( .A1(n6273), .A2(n6899), .ZN(n6212) );
  OR2_X1 U7863 ( .A1(n10072), .A2(n7464), .ZN(n6549) );
  NAND2_X1 U7864 ( .A1(n10072), .A2(n7464), .ZN(n6548) );
  NAND2_X1 U7865 ( .A1(n6747), .A2(n6457), .ZN(n6219) );
  INV_X1 U7866 ( .A(n6216), .ZN(n6642) );
  NAND2_X1 U7867 ( .A1(n6642), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6217) );
  XNOR2_X1 U7868 ( .A(n6217), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7019) );
  AOI22_X1 U7869 ( .A1(n6410), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6861), .B2(
        n7019), .ZN(n6218) );
  NAND2_X1 U7870 ( .A1(n6439), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6227) );
  INV_X1 U7871 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n6220) );
  OR2_X1 U7872 ( .A1(n6388), .A2(n6220), .ZN(n6226) );
  NOR2_X1 U7873 ( .A1(n6221), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6222) );
  OR2_X1 U7874 ( .A1(n6243), .A2(n6222), .ZN(n7463) );
  OR2_X1 U7875 ( .A1(n6421), .A2(n7463), .ZN(n6225) );
  INV_X1 U7876 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6223) );
  OR2_X1 U7877 ( .A1(n6273), .A2(n6223), .ZN(n6224) );
  NAND4_X1 U7878 ( .A1(n6227), .A2(n6226), .A3(n6225), .A4(n6224), .ZN(n10061)
         );
  INV_X1 U7879 ( .A(n10061), .ZN(n7351) );
  NAND2_X1 U7880 ( .A1(n7761), .A2(n7351), .ZN(n6509) );
  NAND2_X1 U7881 ( .A1(n6756), .A2(n6457), .ZN(n6230) );
  OR2_X2 U7882 ( .A1(n6642), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U7883 ( .A1(n6450), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6228) );
  XNOR2_X1 U7884 ( .A(n6228), .B(P2_IR_REG_9__SCAN_IN), .ZN(n7031) );
  AOI22_X1 U7885 ( .A1(n6410), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6861), .B2(
        n7031), .ZN(n6229) );
  NAND2_X1 U7886 ( .A1(n6443), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6234) );
  XNOR2_X1 U7887 ( .A(n6243), .B(P2_REG3_REG_9__SCAN_IN), .ZN(n7777) );
  OR2_X1 U7888 ( .A1(n6421), .A2(n7777), .ZN(n6233) );
  INV_X1 U7889 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n7022) );
  OR2_X1 U7890 ( .A1(n6273), .A2(n7022), .ZN(n6232) );
  INV_X1 U7891 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n7032) );
  OR2_X1 U7892 ( .A1(n6444), .A2(n7032), .ZN(n6231) );
  NAND4_X1 U7893 ( .A1(n6234), .A2(n6233), .A3(n6232), .A4(n6231), .ZN(n10004)
         );
  INV_X1 U7894 ( .A(n10004), .ZN(n6235) );
  OR2_X1 U7895 ( .A1(n8957), .A2(n6235), .ZN(n6505) );
  NAND2_X1 U7896 ( .A1(n8957), .A2(n6235), .ZN(n6553) );
  NAND2_X1 U7897 ( .A1(n6505), .A2(n6553), .ZN(n7821) );
  INV_X1 U7898 ( .A(n7821), .ZN(n7766) );
  NAND2_X1 U7899 ( .A1(n7769), .A2(n7766), .ZN(n6236) );
  INV_X1 U7900 ( .A(n6450), .ZN(n6237) );
  NAND2_X1 U7901 ( .A1(n6237), .A2(n6095), .ZN(n6261) );
  AND2_X1 U7902 ( .A1(n6261), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6238) );
  NAND2_X1 U7903 ( .A1(n6238), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n6241) );
  INV_X1 U7904 ( .A(n6238), .ZN(n6240) );
  NAND2_X1 U7905 ( .A1(n6240), .A2(n6239), .ZN(n6249) );
  AOI22_X1 U7906 ( .A1(n6410), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n7153), .B2(
        n6861), .ZN(n6242) );
  NAND2_X1 U7907 ( .A1(n6443), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n6248) );
  AOI21_X1 U7908 ( .B1(n6243), .B2(P2_REG3_REG_9__SCAN_IN), .A(
        P2_REG3_REG_10__SCAN_IN), .ZN(n6244) );
  OR2_X1 U7909 ( .A1(n6253), .A2(n6244), .ZN(n10017) );
  OR2_X1 U7910 ( .A1(n6421), .A2(n10017), .ZN(n6247) );
  INV_X1 U7911 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n7025) );
  OR2_X1 U7912 ( .A1(n6273), .A2(n7025), .ZN(n6246) );
  INV_X1 U7913 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n7146) );
  OR2_X1 U7914 ( .A1(n6444), .A2(n7146), .ZN(n6245) );
  NAND2_X1 U7915 ( .A1(n6777), .A2(n6457), .ZN(n6252) );
  NAND2_X1 U7916 ( .A1(n6249), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6250) );
  XNOR2_X1 U7917 ( .A(n6250), .B(P2_IR_REG_11__SCAN_IN), .ZN(n7259) );
  AOI22_X1 U7918 ( .A1(n7259), .A2(n6861), .B1(n6410), .B2(
        P1_DATAO_REG_11__SCAN_IN), .ZN(n6251) );
  NAND2_X1 U7919 ( .A1(n6443), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6259) );
  INV_X1 U7920 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n7266) );
  OR2_X1 U7921 ( .A1(n6444), .A2(n7266), .ZN(n6258) );
  INV_X1 U7922 ( .A(n6253), .ZN(n6254) );
  INV_X1 U7923 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n7156) );
  NAND2_X1 U7924 ( .A1(n6254), .A2(n7156), .ZN(n6255) );
  NAND2_X1 U7925 ( .A1(n6270), .A2(n6255), .ZN(n10054) );
  OR2_X1 U7926 ( .A1(n6421), .A2(n10054), .ZN(n6257) );
  INV_X1 U7927 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n7150) );
  OR2_X1 U7928 ( .A1(n6273), .A2(n7150), .ZN(n6256) );
  NAND2_X1 U7929 ( .A1(n10051), .A2(n10008), .ZN(n6558) );
  AND2_X1 U7930 ( .A1(n6558), .A2(n7813), .ZN(n6260) );
  NAND2_X1 U7931 ( .A1(n7008), .A2(n6457), .ZN(n6266) );
  INV_X1 U7932 ( .A(n6261), .ZN(n6263) );
  NOR2_X1 U7933 ( .A1(P2_IR_REG_10__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n6262) );
  NAND2_X1 U7934 ( .A1(n6263), .A2(n6262), .ZN(n6279) );
  NAND2_X1 U7935 ( .A1(n6279), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6264) );
  XNOR2_X1 U7936 ( .A(n6264), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7268) );
  AOI22_X1 U7937 ( .A1(n6410), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n7268), .B2(
        n6861), .ZN(n6265) );
  NAND2_X1 U7938 ( .A1(n6439), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n6277) );
  INV_X1 U7939 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n6267) );
  OR2_X1 U7940 ( .A1(n6388), .A2(n6267), .ZN(n6276) );
  INV_X1 U7941 ( .A(n6268), .ZN(n6291) );
  INV_X1 U7942 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n6269) );
  NAND2_X1 U7943 ( .A1(n6270), .A2(n6269), .ZN(n6271) );
  NAND2_X1 U7944 ( .A1(n6291), .A2(n6271), .ZN(n7982) );
  OR2_X1 U7945 ( .A1(n6421), .A2(n7982), .ZN(n6275) );
  INV_X1 U7946 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n6272) );
  OR2_X1 U7947 ( .A1(n6273), .A2(n6272), .ZN(n6274) );
  NAND4_X1 U7948 ( .A1(n6277), .A2(n6276), .A3(n6275), .A4(n6274), .ZN(n10035)
         );
  INV_X1 U7949 ( .A(n10035), .ZN(n6278) );
  NAND2_X1 U7950 ( .A1(n8941), .A2(n6278), .ZN(n6566) );
  NAND2_X1 U7951 ( .A1(n7015), .A2(n6457), .ZN(n6282) );
  NAND2_X1 U7952 ( .A1(n6319), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U7953 ( .A1(n6287), .A2(n6315), .ZN(n6280) );
  NAND2_X1 U7954 ( .A1(n6280), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6299) );
  XNOR2_X1 U7955 ( .A(n6299), .B(P2_IR_REG_14__SCAN_IN), .ZN(n7936) );
  AOI22_X1 U7956 ( .A1(n7936), .A2(n6861), .B1(n6410), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n6281) );
  XNOR2_X1 U7957 ( .A(n6308), .B(P2_REG3_REG_14__SCAN_IN), .ZN(n8065) );
  NAND2_X1 U7958 ( .A1(n8065), .A2(n6435), .ZN(n6286) );
  INV_X1 U7959 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7935) );
  OR2_X1 U7960 ( .A1(n6444), .A2(n7935), .ZN(n6285) );
  NAND2_X1 U7961 ( .A1(n6385), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6284) );
  INV_X1 U7962 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n9711) );
  OR2_X1 U7963 ( .A1(n6388), .A2(n9711), .ZN(n6283) );
  NAND2_X1 U7964 ( .A1(n7074), .A2(n6457), .ZN(n6289) );
  XNOR2_X1 U7965 ( .A(n6287), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7382) );
  AOI22_X1 U7966 ( .A1(n7382), .A2(n6861), .B1(n6410), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7967 ( .A1(n6443), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6297) );
  INV_X1 U7968 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8051) );
  OR2_X1 U7969 ( .A1(n6444), .A2(n8051), .ZN(n6296) );
  INV_X1 U7970 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n6290) );
  NAND2_X1 U7971 ( .A1(n6291), .A2(n6290), .ZN(n6292) );
  NAND2_X1 U7972 ( .A1(n6308), .A2(n6292), .ZN(n8455) );
  OR2_X1 U7973 ( .A1(n6421), .A2(n8455), .ZN(n6295) );
  INV_X1 U7974 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n6293) );
  OR2_X1 U7975 ( .A1(n6273), .A2(n6293), .ZN(n6294) );
  NAND2_X1 U7976 ( .A1(n8934), .A2(n8068), .ZN(n8016) );
  NAND2_X1 U7977 ( .A1(n8929), .A2(n8499), .ZN(n6570) );
  NAND2_X1 U7978 ( .A1(n8016), .A2(n6570), .ZN(n6298) );
  NAND2_X1 U7979 ( .A1(n6298), .A2(n8142), .ZN(n6313) );
  NAND2_X1 U7980 ( .A1(n7090), .A2(n6457), .ZN(n6303) );
  NAND2_X1 U7981 ( .A1(n6299), .A2(n6317), .ZN(n6300) );
  NAND2_X1 U7982 ( .A1(n6300), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6301) );
  XNOR2_X1 U7983 ( .A(n6301), .B(P2_IR_REG_15__SCAN_IN), .ZN(n8188) );
  AOI22_X1 U7984 ( .A1(n8188), .A2(n6861), .B1(n6410), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n6302) );
  INV_X1 U7985 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n6304) );
  OR2_X1 U7986 ( .A1(n6444), .A2(n6304), .ZN(n6307) );
  INV_X1 U7987 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n6305) );
  OR2_X1 U7988 ( .A1(n6388), .A2(n6305), .ZN(n6306) );
  AND2_X1 U7989 ( .A1(n6307), .A2(n6306), .ZN(n6312) );
  OAI21_X1 U7990 ( .B1(n6308), .B2(n7629), .A(n8500), .ZN(n6309) );
  AND2_X1 U7991 ( .A1(n6309), .A2(n6326), .ZN(n8504) );
  NAND2_X1 U7992 ( .A1(n8504), .A2(n6435), .ZN(n6311) );
  NAND2_X1 U7993 ( .A1(n6385), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U7994 ( .A1(n8924), .A2(n8270), .ZN(n6573) );
  NAND2_X1 U7995 ( .A1(n7170), .A2(n6457), .ZN(n6325) );
  NAND3_X1 U7996 ( .A1(n6317), .A2(n6316), .A3(n6315), .ZN(n6318) );
  OAI21_X1 U7997 ( .B1(n6319), .B2(n6318), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n6320) );
  MUX2_X1 U7998 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6320), .S(
        P2_IR_REG_16__SCAN_IN), .Z(n6321) );
  NAND2_X1 U7999 ( .A1(n6321), .A2(n6331), .ZN(n8557) );
  OAI22_X1 U8000 ( .A1(n8557), .A2(n6859), .B1(n6322), .B2(n7172), .ZN(n6323)
         );
  INV_X1 U8001 ( .A(n6323), .ZN(n6324) );
  INV_X1 U8002 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n8556) );
  NAND2_X1 U8003 ( .A1(n6326), .A2(n8556), .ZN(n6327) );
  NAND2_X1 U8004 ( .A1(n6336), .A2(n6327), .ZN(n8799) );
  OR2_X1 U8005 ( .A1(n8799), .A2(n6421), .ZN(n6330) );
  AOI22_X1 U8006 ( .A1(n6439), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n6443), .B2(
        P2_REG0_REG_16__SCAN_IN), .ZN(n6329) );
  NAND2_X1 U8007 ( .A1(n6385), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n6328) );
  NAND2_X1 U8008 ( .A1(n8919), .A2(n8501), .ZN(n6579) );
  NAND2_X1 U8009 ( .A1(n7217), .A2(n6457), .ZN(n6334) );
  NAND2_X1 U8010 ( .A1(n6331), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6332) );
  XNOR2_X1 U8011 ( .A(n6332), .B(P2_IR_REG_17__SCAN_IN), .ZN(n8204) );
  AOI22_X1 U8012 ( .A1(n6410), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6861), .B2(
        n8204), .ZN(n6333) );
  INV_X1 U8013 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n6335) );
  NAND2_X1 U8014 ( .A1(n6336), .A2(n6335), .ZN(n6337) );
  NAND2_X1 U8015 ( .A1(n6345), .A2(n6337), .ZN(n8783) );
  OR2_X1 U8016 ( .A1(n8783), .A2(n6421), .ZN(n6340) );
  AOI22_X1 U8017 ( .A1(n6439), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n6443), .B2(
        P2_REG0_REG_17__SCAN_IN), .ZN(n6339) );
  NAND2_X1 U8018 ( .A1(n6385), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U8019 ( .A1(n8915), .A2(n8477), .ZN(n6500) );
  NAND2_X1 U8020 ( .A1(n8772), .A2(n6498), .ZN(n8759) );
  NAND2_X1 U8021 ( .A1(n7340), .A2(n6457), .ZN(n6343) );
  XNOR2_X1 U8022 ( .A(n6341), .B(P2_IR_REG_18__SCAN_IN), .ZN(n8202) );
  AOI22_X1 U8023 ( .A1(n6410), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6861), .B2(
        n8202), .ZN(n6342) );
  NAND2_X1 U8024 ( .A1(n6345), .A2(n6344), .ZN(n6346) );
  NAND2_X1 U8025 ( .A1(n6347), .A2(n6346), .ZN(n8481) );
  AOI22_X1 U8026 ( .A1(n6439), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n6443), .B2(
        P2_REG0_REG_18__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U8027 ( .A1(n6385), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6348) );
  OAI211_X1 U8028 ( .C1(n8481), .C2(n6421), .A(n6349), .B(n6348), .ZN(n8514)
         );
  INV_X1 U8029 ( .A(n8514), .ZN(n8743) );
  OR2_X1 U8030 ( .A1(n8909), .A2(n8743), .ZN(n6595) );
  OR2_X1 U8031 ( .A1(n8755), .A2(n8729), .ZN(n6594) );
  OAI21_X1 U8032 ( .B1(n6583), .B2(n6594), .A(n8710), .ZN(n6359) );
  NAND2_X1 U8033 ( .A1(n7620), .A2(n6457), .ZN(n6352) );
  NAND2_X1 U8034 ( .A1(n6410), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n6351) );
  XNOR2_X1 U8035 ( .A(n6364), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n8705) );
  NAND2_X1 U8036 ( .A1(n8705), .A2(n6435), .ZN(n6358) );
  INV_X1 U8037 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n6355) );
  NAND2_X1 U8038 ( .A1(n6439), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n6354) );
  NAND2_X1 U8039 ( .A1(n6443), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n6353) );
  OAI211_X1 U8040 ( .C1(n6355), .C2(n6273), .A(n6354), .B(n6353), .ZN(n6356)
         );
  INV_X1 U8041 ( .A(n6356), .ZN(n6357) );
  NAND2_X1 U8042 ( .A1(n6358), .A2(n6357), .ZN(n8513) );
  INV_X1 U8043 ( .A(n8513), .ZN(n8730) );
  XNOR2_X1 U8044 ( .A(n8893), .B(n8730), .ZN(n8711) );
  NAND2_X1 U8045 ( .A1(n7743), .A2(n6457), .ZN(n6362) );
  NAND2_X1 U8046 ( .A1(n6410), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n6361) );
  INV_X1 U8047 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n8379) );
  INV_X1 U8048 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n6363) );
  OAI21_X1 U8049 ( .B1(n6364), .B2(n8379), .A(n6363), .ZN(n6367) );
  AND2_X1 U8050 ( .A1(P2_REG3_REG_21__SCAN_IN), .A2(P2_REG3_REG_22__SCAN_IN), 
        .ZN(n6365) );
  NAND2_X1 U8051 ( .A1(n6367), .A2(n6376), .ZN(n8689) );
  OR2_X1 U8052 ( .A1(n8689), .A2(n6421), .ZN(n6373) );
  INV_X1 U8053 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n6370) );
  NAND2_X1 U8054 ( .A1(n6439), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6369) );
  NAND2_X1 U8055 ( .A1(n6443), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n6368) );
  OAI211_X1 U8056 ( .C1(n6370), .C2(n6273), .A(n6369), .B(n6368), .ZN(n6371)
         );
  INV_X1 U8057 ( .A(n6371), .ZN(n6372) );
  NAND2_X1 U8058 ( .A1(n6373), .A2(n6372), .ZN(n8715) );
  INV_X1 U8059 ( .A(n8715), .ZN(n8677) );
  INV_X1 U8060 ( .A(n6588), .ZN(n6603) );
  NAND2_X1 U8061 ( .A1(n8693), .A2(n6603), .ZN(n8674) );
  NAND2_X1 U8062 ( .A1(n7782), .A2(n6457), .ZN(n6375) );
  NAND2_X1 U8063 ( .A1(n6410), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n6374) );
  INV_X1 U8064 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9666) );
  NAND2_X1 U8065 ( .A1(n6376), .A2(n9666), .ZN(n6377) );
  NAND2_X1 U8066 ( .A1(n6394), .A2(n6377), .ZN(n8330) );
  OR2_X1 U8067 ( .A1(n8330), .A2(n6421), .ZN(n6382) );
  INV_X1 U8068 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9722) );
  NAND2_X1 U8069 ( .A1(n6439), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6379) );
  NAND2_X1 U8070 ( .A1(n6443), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6378) );
  OAI211_X1 U8071 ( .C1(n9722), .C2(n6273), .A(n6379), .B(n6378), .ZN(n6380)
         );
  INV_X1 U8072 ( .A(n6380), .ZN(n6381) );
  NAND2_X1 U8073 ( .A1(n6382), .A2(n6381), .ZN(n8658) );
  XNOR2_X1 U8074 ( .A(n8883), .B(n8658), .ZN(n8681) );
  INV_X1 U8075 ( .A(n8681), .ZN(n8675) );
  INV_X1 U8076 ( .A(n8658), .ZN(n8423) );
  AND2_X1 U8077 ( .A1(n8883), .A2(n8423), .ZN(n6591) );
  NAND2_X1 U8078 ( .A1(n7914), .A2(n6457), .ZN(n6384) );
  NAND2_X1 U8079 ( .A1(n6410), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n6383) );
  XNOR2_X1 U8080 ( .A(n6394), .B(P2_REG3_REG_24__SCAN_IN), .ZN(n8666) );
  INV_X1 U8081 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9663) );
  NAND2_X1 U8082 ( .A1(n6439), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6387) );
  NAND2_X1 U8083 ( .A1(n6385), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6386) );
  OAI211_X1 U8084 ( .C1(n6388), .C2(n9663), .A(n6387), .B(n6386), .ZN(n6389)
         );
  AOI21_X1 U8085 ( .B1(n8666), .B2(n6435), .A(n6389), .ZN(n8678) );
  NAND2_X1 U8086 ( .A1(n8667), .A2(n8678), .ZN(n6610) );
  NAND2_X1 U8087 ( .A1(n6606), .A2(n6610), .ZN(n8663) );
  NAND2_X1 U8088 ( .A1(n8091), .A2(n6457), .ZN(n6391) );
  NAND2_X1 U8089 ( .A1(n6410), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n6390) );
  NAND2_X1 U8090 ( .A1(P2_REG3_REG_25__SCAN_IN), .A2(P2_REG3_REG_24__SCAN_IN), 
        .ZN(n6392) );
  INV_X1 U8091 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n8424) );
  INV_X1 U8092 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n6393) );
  OAI21_X1 U8093 ( .B1(n6394), .B2(n8424), .A(n6393), .ZN(n6395) );
  INV_X1 U8094 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n6398) );
  NAND2_X1 U8095 ( .A1(n6439), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6397) );
  NAND2_X1 U8096 ( .A1(n6443), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6396) );
  OAI211_X1 U8097 ( .C1(n6398), .C2(n6273), .A(n6397), .B(n6396), .ZN(n6399)
         );
  AOI21_X1 U8098 ( .B1(n8650), .B2(n6435), .A(n6399), .ZN(n8661) );
  NAND2_X1 U8099 ( .A1(n8873), .A2(n8661), .ZN(n6494) );
  NAND2_X1 U8100 ( .A1(n8999), .A2(n6457), .ZN(n6401) );
  NAND2_X1 U8101 ( .A1(n6410), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n6400) );
  INV_X1 U8102 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n8491) );
  NAND2_X1 U8103 ( .A1(n6402), .A2(n8491), .ZN(n6403) );
  NAND2_X1 U8104 ( .A1(n6419), .A2(n6403), .ZN(n8639) );
  INV_X1 U8105 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n6406) );
  NAND2_X1 U8106 ( .A1(n6443), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n6405) );
  NAND2_X1 U8107 ( .A1(n6439), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6404) );
  OAI211_X1 U8108 ( .C1(n6273), .C2(n6406), .A(n6405), .B(n6404), .ZN(n6407)
         );
  INV_X1 U8109 ( .A(n6407), .ZN(n6408) );
  NAND2_X1 U8110 ( .A1(n8997), .A2(n6457), .ZN(n6412) );
  NAND2_X1 U8111 ( .A1(n6410), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n6411) );
  XNOR2_X1 U8112 ( .A(n6419), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n8621) );
  INV_X1 U8113 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n6415) );
  NAND2_X1 U8114 ( .A1(n6443), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6414) );
  NAND2_X1 U8115 ( .A1(n6439), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6413) );
  OAI211_X1 U8116 ( .C1(n6273), .C2(n6415), .A(n6414), .B(n6413), .ZN(n6416)
         );
  NAND2_X1 U8117 ( .A1(n8861), .A2(n8608), .ZN(n6618) );
  NAND2_X1 U8118 ( .A1(n9788), .A2(n6457), .ZN(n6418) );
  NAND2_X1 U8119 ( .A1(n6410), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6417) );
  INV_X1 U8120 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n8322) );
  INV_X1 U8121 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n8369) );
  OAI21_X1 U8122 ( .B1(n6419), .B2(n8322), .A(n8369), .ZN(n6420) );
  NAND2_X1 U8123 ( .A1(n6420), .A2(n6430), .ZN(n8368) );
  INV_X1 U8124 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U8125 ( .A1(n6439), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6423) );
  NAND2_X1 U8126 ( .A1(n6443), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6422) );
  OAI211_X1 U8127 ( .C1(n6424), .C2(n6273), .A(n6423), .B(n6422), .ZN(n6425)
         );
  INV_X1 U8128 ( .A(n6425), .ZN(n6426) );
  NAND2_X1 U8129 ( .A1(n8856), .A2(n8355), .ZN(n6621) );
  NAND2_X1 U8130 ( .A1(n8610), .A2(n6620), .ZN(n8222) );
  INV_X1 U8131 ( .A(n8222), .ZN(n6436) );
  NAND2_X1 U8132 ( .A1(n8992), .A2(n6457), .ZN(n6429) );
  NAND2_X1 U8133 ( .A1(n6410), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6428) );
  INV_X1 U8134 ( .A(n6430), .ZN(n8252) );
  INV_X1 U8135 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n6433) );
  NAND2_X1 U8136 ( .A1(n6443), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6432) );
  NAND2_X1 U8137 ( .A1(n6439), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6431) );
  OAI211_X1 U8138 ( .C1(n6273), .C2(n6433), .A(n6432), .B(n6431), .ZN(n6434)
         );
  AOI21_X1 U8139 ( .B1(n8252), .B2(n6435), .A(n6434), .ZN(n8607) );
  NAND2_X1 U8140 ( .A1(n8852), .A2(n8607), .ZN(n6626) );
  NAND2_X1 U8141 ( .A1(n8218), .A2(n6457), .ZN(n6438) );
  NAND2_X1 U8142 ( .A1(n6410), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n6437) );
  INV_X1 U8143 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6442) );
  NAND2_X1 U8144 ( .A1(n6439), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n6441) );
  NAND2_X1 U8145 ( .A1(n6443), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6440) );
  OAI211_X1 U8146 ( .C1(n6273), .C2(n6442), .A(n6441), .B(n6440), .ZN(n8511)
         );
  INV_X1 U8147 ( .A(n8511), .ZN(n6461) );
  NOR2_X1 U8148 ( .A1(n8847), .A2(n6461), .ZN(n6623) );
  INV_X1 U8149 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n6447) );
  NAND2_X1 U8150 ( .A1(n6443), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6446) );
  INV_X1 U8151 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n8262) );
  OR2_X1 U8152 ( .A1(n6444), .A2(n8262), .ZN(n6445) );
  OAI211_X1 U8153 ( .C1(n6273), .C2(n6447), .A(n6446), .B(n6445), .ZN(n8510)
         );
  NOR2_X2 U8155 ( .A1(n6450), .A2(n6449), .ZN(n6454) );
  INV_X1 U8156 ( .A(n6454), .ZN(n6451) );
  NAND2_X1 U8157 ( .A1(n6451), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6452) );
  MUX2_X1 U8158 ( .A(n6452), .B(P2_IR_REG_31__SCAN_IN), .S(n6453), .Z(n6455)
         );
  NAND2_X1 U8159 ( .A1(n6454), .A2(n6453), .ZN(n6466) );
  NAND2_X1 U8160 ( .A1(n6455), .A2(n6466), .ZN(n7621) );
  NAND2_X1 U8161 ( .A1(n8984), .A2(n6457), .ZN(n6459) );
  NAND2_X1 U8162 ( .A1(n6410), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n6458) );
  INV_X1 U8163 ( .A(n8510), .ZN(n6460) );
  OR2_X1 U8164 ( .A1(n8844), .A2(n6460), .ZN(n6629) );
  NAND2_X1 U8165 ( .A1(n8847), .A2(n6461), .ZN(n6628) );
  XNOR2_X1 U8166 ( .A(n6462), .B(n8637), .ZN(n6476) );
  XNOR2_X2 U8167 ( .A(n6468), .B(P2_IR_REG_22__SCAN_IN), .ZN(n6709) );
  INV_X1 U8168 ( .A(n7508), .ZN(n7608) );
  NAND2_X1 U8169 ( .A1(n7608), .A2(n4743), .ZN(n7236) );
  INV_X1 U8170 ( .A(n7236), .ZN(n6473) );
  INV_X1 U8171 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U8172 ( .A1(n6468), .A2(n6467), .ZN(n6469) );
  NAND2_X1 U8173 ( .A1(n6469), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6471) );
  INV_X1 U8174 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U8175 ( .A1(n6471), .A2(n6470), .ZN(n6638) );
  OR2_X1 U8176 ( .A1(n6471), .A2(n6470), .ZN(n6472) );
  NAND2_X1 U8177 ( .A1(n6638), .A2(n6472), .ZN(n6713) );
  NOR2_X1 U8178 ( .A1(n6713), .A2(P2_U3152), .ZN(n6637) );
  INV_X1 U8179 ( .A(n6474), .ZN(n6475) );
  NAND2_X1 U8180 ( .A1(n6476), .A2(n6475), .ZN(n6658) );
  NOR2_X1 U8181 ( .A1(n6632), .A2(n6623), .ZN(n6492) );
  INV_X1 U8182 ( .A(n8632), .ZN(n8628) );
  INV_X1 U8183 ( .A(n8694), .ZN(n8687) );
  NAND2_X1 U8184 ( .A1(n8710), .A2(n6599), .ZN(n8727) );
  NAND2_X1 U8185 ( .A1(n6497), .A2(n6579), .ZN(n8807) );
  NAND2_X1 U8186 ( .A1(n8142), .A2(n6570), .ZN(n8228) );
  NAND2_X1 U8187 ( .A1(n6565), .A2(n6566), .ZN(n8024) );
  INV_X1 U8188 ( .A(n8024), .ZN(n7878) );
  NAND2_X1 U8189 ( .A1(n6557), .A2(n6558), .ZN(n7825) );
  NAND2_X1 U8190 ( .A1(n6513), .A2(n6516), .ZN(n7231) );
  INV_X1 U8191 ( .A(n6477), .ZN(n6478) );
  NOR2_X1 U8192 ( .A1(n7231), .A2(n6478), .ZN(n7695) );
  NAND2_X1 U8193 ( .A1(n6479), .A2(n7688), .ZN(n7680) );
  NAND4_X1 U8194 ( .A1(n7238), .A2(n7608), .A3(n7695), .A4(n7680), .ZN(n6480)
         );
  NAND2_X1 U8195 ( .A1(n6529), .A2(n6537), .ZN(n7740) );
  NAND2_X1 U8196 ( .A1(n6519), .A2(n7730), .ZN(n7655) );
  NOR4_X1 U8197 ( .A1(n6480), .A2(n7597), .A3(n7740), .A4(n7655), .ZN(n6481)
         );
  NAND4_X1 U8198 ( .A1(n7766), .A2(n10064), .A3(n10087), .A4(n6481), .ZN(n6482) );
  INV_X1 U8199 ( .A(n7763), .ZN(n7668) );
  NAND3_X1 U8200 ( .A1(n8028), .A2(n7878), .A3(n6483), .ZN(n6484) );
  NAND2_X1 U8201 ( .A1(n6568), .A2(n8016), .ZN(n8037) );
  NAND4_X1 U8202 ( .A1(n8738), .A2(n8781), .A3(n8767), .A4(n6485), .ZN(n6486)
         );
  NAND4_X1 U8203 ( .A1(n8646), .A2(n8657), .A3(n6487), .A4(n8681), .ZN(n6488)
         );
  OAI22_X1 U8204 ( .A1(n6490), .A2(n4743), .B1(n7608), .B2(n7235), .ZN(n6636)
         );
  NOR2_X1 U8205 ( .A1(n8637), .A2(n7621), .ZN(n6491) );
  OAI211_X1 U8206 ( .C1(n8242), .C2(n6610), .A(n8632), .B(n6494), .ZN(n6495)
         );
  NAND2_X1 U8207 ( .A1(n6495), .A2(n6630), .ZN(n6611) );
  INV_X1 U8208 ( .A(n6496), .ZN(n6587) );
  INV_X1 U8209 ( .A(n6497), .ZN(n8773) );
  NAND2_X1 U8210 ( .A1(n8781), .A2(n8773), .ZN(n6499) );
  NAND3_X1 U8211 ( .A1(n6499), .A2(n6595), .A3(n6498), .ZN(n6502) );
  INV_X1 U8212 ( .A(n6500), .ZN(n6501) );
  MUX2_X1 U8213 ( .A(n6502), .B(n6501), .S(n6624), .Z(n6503) );
  INV_X1 U8214 ( .A(n6503), .ZN(n6580) );
  OAI21_X1 U8215 ( .B1(n7351), .B2(n7761), .A(n6505), .ZN(n6506) );
  NAND2_X1 U8216 ( .A1(n6556), .A2(n6506), .ZN(n6508) );
  NAND3_X1 U8217 ( .A1(n6508), .A2(n6557), .A3(n6507), .ZN(n6512) );
  INV_X1 U8218 ( .A(n6556), .ZN(n6510) );
  OAI211_X1 U8219 ( .C1(n6510), .C2(n6509), .A(n6558), .B(n7813), .ZN(n6511)
         );
  AND2_X1 U8220 ( .A1(n7680), .A2(n4743), .ZN(n6523) );
  INV_X1 U8221 ( .A(n6523), .ZN(n6514) );
  NAND2_X1 U8222 ( .A1(n6514), .A2(n6513), .ZN(n6517) );
  AND2_X1 U8223 ( .A1(n6516), .A2(n6515), .ZN(n6521) );
  NAND2_X1 U8224 ( .A1(n6517), .A2(n6521), .ZN(n6518) );
  NAND2_X1 U8225 ( .A1(n6518), .A2(n6524), .ZN(n6536) );
  AND2_X1 U8226 ( .A1(n6529), .A2(n6519), .ZN(n6520) );
  OAI21_X1 U8227 ( .B1(n6523), .B2(n6522), .A(n6521), .ZN(n6526) );
  AND2_X1 U8228 ( .A1(n6524), .A2(n6630), .ZN(n6525) );
  AOI21_X1 U8229 ( .B1(n6526), .B2(n6525), .A(n7597), .ZN(n6527) );
  NAND2_X1 U8230 ( .A1(n6542), .A2(n6527), .ZN(n6535) );
  INV_X1 U8231 ( .A(n6528), .ZN(n6531) );
  NAND2_X1 U8232 ( .A1(n6547), .A2(n6529), .ZN(n6530) );
  NAND2_X1 U8233 ( .A1(n6532), .A2(n6535), .ZN(n6533) );
  NAND2_X1 U8234 ( .A1(n6533), .A2(n6630), .ZN(n6534) );
  OAI21_X1 U8235 ( .B1(n6536), .B2(n6535), .A(n6534), .ZN(n6546) );
  INV_X1 U8236 ( .A(n6537), .ZN(n6541) );
  NAND2_X1 U8237 ( .A1(n6539), .A2(n6538), .ZN(n6540) );
  OAI21_X1 U8238 ( .B1(n6542), .B2(n6541), .A(n6540), .ZN(n6543) );
  AOI21_X1 U8239 ( .B1(n6543), .B2(n6545), .A(n6630), .ZN(n6544) );
  OAI21_X1 U8240 ( .B1(n6547), .B2(n6630), .A(n10064), .ZN(n6551) );
  MUX2_X1 U8241 ( .A(n6549), .B(n6548), .S(n6630), .Z(n6550) );
  OAI211_X1 U8242 ( .C1(n6552), .C2(n6551), .A(n7763), .B(n6550), .ZN(n6554)
         );
  NAND2_X1 U8243 ( .A1(n6554), .A2(n6553), .ZN(n6555) );
  NAND2_X1 U8244 ( .A1(n6565), .A2(n6557), .ZN(n6560) );
  NAND2_X1 U8245 ( .A1(n6566), .A2(n6558), .ZN(n6559) );
  MUX2_X1 U8246 ( .A(n6560), .B(n6559), .S(n6630), .Z(n6561) );
  INV_X1 U8247 ( .A(n6561), .ZN(n6562) );
  INV_X1 U8248 ( .A(n8037), .ZN(n8042) );
  MUX2_X1 U8249 ( .A(n6566), .B(n6565), .S(n6630), .Z(n6567) );
  MUX2_X1 U8250 ( .A(n8016), .B(n6568), .S(n6624), .Z(n6569) );
  INV_X1 U8251 ( .A(n8231), .ZN(n6572) );
  MUX2_X1 U8252 ( .A(n8142), .B(n6570), .S(n6624), .Z(n6571) );
  INV_X1 U8253 ( .A(n8807), .ZN(n6576) );
  MUX2_X1 U8254 ( .A(n6574), .B(n6573), .S(n6630), .Z(n6575) );
  NAND3_X1 U8255 ( .A1(n6577), .A2(n6576), .A3(n6575), .ZN(n6578) );
  INV_X1 U8256 ( .A(n6594), .ZN(n6581) );
  OR2_X1 U8257 ( .A1(n8893), .A2(n8730), .ZN(n6602) );
  NAND2_X1 U8258 ( .A1(n6588), .A2(n6630), .ZN(n6589) );
  NAND3_X1 U8259 ( .A1(n6590), .A2(n8681), .A3(n6589), .ZN(n6593) );
  NAND2_X1 U8260 ( .A1(n6591), .A2(n6630), .ZN(n6592) );
  NAND2_X1 U8261 ( .A1(n6593), .A2(n6592), .ZN(n6605) );
  NAND3_X1 U8262 ( .A1(n6596), .A2(n6595), .A3(n6594), .ZN(n6597) );
  NAND2_X1 U8263 ( .A1(n6597), .A2(n8709), .ZN(n6598) );
  NAND2_X1 U8264 ( .A1(n6598), .A2(n8710), .ZN(n6600) );
  NAND3_X1 U8265 ( .A1(n6600), .A2(n4282), .A3(n6599), .ZN(n6601) );
  NAND4_X1 U8266 ( .A1(n6603), .A2(n6624), .A3(n6602), .A4(n6601), .ZN(n6604)
         );
  OAI21_X1 U8267 ( .B1(n8423), .B2(n8883), .A(n6606), .ZN(n6607) );
  NAND2_X1 U8268 ( .A1(n6607), .A2(n6624), .ZN(n6608) );
  AOI21_X1 U8269 ( .B1(n6613), .B2(n8630), .A(n6630), .ZN(n6612) );
  AOI21_X1 U8270 ( .B1(n6614), .B2(n6613), .A(n6612), .ZN(n6616) );
  MUX2_X1 U8271 ( .A(n6618), .B(n6617), .S(n6624), .Z(n6619) );
  MUX2_X1 U8272 ( .A(n6621), .B(n6620), .S(n6630), .Z(n6622) );
  MUX2_X1 U8273 ( .A(n6626), .B(n6625), .S(n6624), .Z(n6627) );
  INV_X1 U8274 ( .A(n6629), .ZN(n6631) );
  MUX2_X1 U8275 ( .A(n6632), .B(n6631), .S(n6630), .Z(n6633) );
  INV_X1 U8276 ( .A(n6637), .ZN(n7783) );
  NAND2_X1 U8277 ( .A1(n6638), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6640) );
  OR2_X1 U8278 ( .A1(n6642), .A2(n6641), .ZN(n6643) );
  NOR2_X1 U8279 ( .A1(n6643), .A2(n6449), .ZN(n6647) );
  NOR2_X1 U8280 ( .A1(n6647), .A2(n6084), .ZN(n6644) );
  MUX2_X1 U8281 ( .A(n6084), .B(n6644), .S(P2_IR_REG_25__SCAN_IN), .Z(n6645)
         );
  INV_X1 U8282 ( .A(n6645), .ZN(n6648) );
  INV_X1 U8283 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n6646) );
  NAND2_X1 U8284 ( .A1(n6647), .A2(n6646), .ZN(n6649) );
  NAND2_X1 U8285 ( .A1(n6648), .A2(n6649), .ZN(n8092) );
  NAND2_X1 U8286 ( .A1(n6649), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6650) );
  MUX2_X1 U8287 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6650), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n6651) );
  INV_X1 U8288 ( .A(n10102), .ZN(n6711) );
  XNOR2_X1 U8289 ( .A(n6652), .B(P2_IR_REG_27__SCAN_IN), .ZN(n8223) );
  NAND2_X1 U8290 ( .A1(n6653), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6654) );
  XNOR2_X1 U8291 ( .A(n6654), .B(n4766), .ZN(n6891) );
  INV_X1 U8292 ( .A(n6891), .ZN(n6655) );
  NAND4_X1 U8293 ( .A1(n6711), .A2(n4247), .A3(n8223), .A4(n10058), .ZN(n6656)
         );
  OAI211_X1 U8294 ( .C1(n6709), .C2(n7783), .A(n6656), .B(P2_B_REG_SCAN_IN), 
        .ZN(n6657) );
  INV_X1 U8295 ( .A(n6856), .ZN(n6659) );
  NAND2_X2 U8296 ( .A1(n6659), .A2(n10111), .ZN(n8518) );
  INV_X1 U8297 ( .A(n6660), .ZN(n6661) );
  OR2_X1 U8298 ( .A1(n7194), .A2(n6661), .ZN(n6662) );
  NAND2_X1 U8299 ( .A1(n6783), .A2(n6663), .ZN(n6770) );
  NAND2_X1 U8300 ( .A1(n6770), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  NOR2_X2 U8301 ( .A1(n6760), .A2(P1_U3084), .ZN(P1_U4006) );
  NAND2_X1 U8302 ( .A1(n7508), .A2(n4743), .ZN(n7604) );
  INV_X4 U8303 ( .A(n8306), .ZN(n8356) );
  XNOR2_X1 U8304 ( .A(n4810), .B(n8356), .ZN(n6664) );
  AND2_X1 U8305 ( .A1(n8310), .A2(n8521), .ZN(n6665) );
  NAND2_X1 U8306 ( .A1(n6664), .A2(n6665), .ZN(n7297) );
  INV_X1 U8307 ( .A(n6664), .ZN(n7294) );
  INV_X1 U8308 ( .A(n6665), .ZN(n6666) );
  NAND2_X1 U8309 ( .A1(n7294), .A2(n6666), .ZN(n6667) );
  NAND2_X1 U8310 ( .A1(n7297), .A2(n6667), .ZN(n6707) );
  NAND2_X1 U8311 ( .A1(n8523), .A2(n8310), .ZN(n6671) );
  INV_X1 U8312 ( .A(n8306), .ZN(n6674) );
  XNOR2_X1 U8313 ( .A(n6674), .B(n6133), .ZN(n6669) );
  XNOR2_X1 U8314 ( .A(n6671), .B(n6669), .ZN(n7211) );
  OR2_X1 U8315 ( .A1(n7698), .A2(n8354), .ZN(n7250) );
  NAND2_X1 U8316 ( .A1(n8306), .A2(n7688), .ZN(n6668) );
  AND2_X1 U8317 ( .A1(n7250), .A2(n6668), .ZN(n7212) );
  INV_X1 U8318 ( .A(n6669), .ZN(n6670) );
  NAND2_X1 U8319 ( .A1(n6671), .A2(n6670), .ZN(n6672) );
  NAND2_X1 U8320 ( .A1(n6673), .A2(n8310), .ZN(n6675) );
  XNOR2_X1 U8321 ( .A(n6674), .B(n7241), .ZN(n10020) );
  NAND2_X1 U8322 ( .A1(n6675), .A2(n10020), .ZN(n6676) );
  NAND2_X1 U8323 ( .A1(n6677), .A2(n6676), .ZN(n7177) );
  XNOR2_X1 U8324 ( .A(n10128), .B(n8356), .ZN(n8438) );
  NAND2_X1 U8325 ( .A1(n8522), .A2(n8310), .ZN(n6678) );
  OR2_X1 U8326 ( .A1(n8438), .A2(n6678), .ZN(n6680) );
  NAND2_X1 U8327 ( .A1(n6678), .A2(n8438), .ZN(n6679) );
  XNOR2_X1 U8328 ( .A(n7610), .B(n8306), .ZN(n6682) );
  NAND2_X1 U8329 ( .A1(n10019), .A2(n8310), .ZN(n6683) );
  XNOR2_X1 U8330 ( .A(n6682), .B(n6683), .ZN(n8437) );
  AND2_X1 U8331 ( .A1(n8437), .A2(n6680), .ZN(n6681) );
  INV_X1 U8332 ( .A(n6682), .ZN(n6684) );
  NAND2_X1 U8333 ( .A1(n6684), .A2(n6683), .ZN(n6685) );
  NAND2_X1 U8334 ( .A1(n8435), .A2(n6685), .ZN(n6706) );
  NOR4_X1 U8335 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_2__SCAN_IN), .A3(
        P2_D_REG_3__SCAN_IN), .A4(P2_D_REG_4__SCAN_IN), .ZN(n6694) );
  INV_X1 U8336 ( .A(P2_D_REG_10__SCAN_IN), .ZN(n10106) );
  INV_X1 U8337 ( .A(P2_D_REG_27__SCAN_IN), .ZN(n10104) );
  INV_X1 U8338 ( .A(P2_D_REG_28__SCAN_IN), .ZN(n10103) );
  INV_X1 U8339 ( .A(P2_D_REG_15__SCAN_IN), .ZN(n10105) );
  NAND4_X1 U8340 ( .A1(n10106), .A2(n10104), .A3(n10103), .A4(n10105), .ZN(
        n6691) );
  NOR4_X1 U8341 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_17__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_19__SCAN_IN), .ZN(n6689) );
  NOR4_X1 U8342 ( .A1(P2_D_REG_13__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_14__SCAN_IN), .ZN(n6688) );
  NOR4_X1 U8343 ( .A1(P2_D_REG_24__SCAN_IN), .A2(P2_D_REG_25__SCAN_IN), .A3(
        P2_D_REG_26__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n6687) );
  NOR4_X1 U8344 ( .A1(P2_D_REG_20__SCAN_IN), .A2(P2_D_REG_21__SCAN_IN), .A3(
        P2_D_REG_22__SCAN_IN), .A4(P2_D_REG_23__SCAN_IN), .ZN(n6686) );
  NAND4_X1 U8345 ( .A1(n6689), .A2(n6688), .A3(n6687), .A4(n6686), .ZN(n6690)
         );
  NOR4_X1 U8346 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n6691), .A4(n6690), .ZN(n6693) );
  NOR4_X1 U8347 ( .A1(P2_D_REG_5__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n6692) );
  NAND3_X1 U8348 ( .A1(n6694), .A2(n6693), .A3(n6692), .ZN(n6698) );
  INV_X1 U8349 ( .A(n9002), .ZN(n6697) );
  XNOR2_X1 U8350 ( .A(n7915), .B(P2_B_REG_SCAN_IN), .ZN(n6695) );
  NAND2_X1 U8351 ( .A1(n8092), .A2(n6695), .ZN(n6696) );
  NAND2_X1 U8352 ( .A1(n6698), .A2(n10101), .ZN(n7224) );
  INV_X1 U8353 ( .A(n7224), .ZN(n6700) );
  INV_X1 U8354 ( .A(n10101), .ZN(n6699) );
  NAND2_X1 U8355 ( .A1(n8092), .A2(n9002), .ZN(n10114) );
  OAI21_X1 U8356 ( .B1(P2_D_REG_1__SCAN_IN), .B2(n6699), .A(n10114), .ZN(n7226) );
  NOR2_X1 U8357 ( .A1(n6700), .A2(n7226), .ZN(n7602) );
  AND2_X1 U8358 ( .A1(n7915), .A2(n9002), .ZN(n10110) );
  INV_X1 U8359 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10109) );
  NAND2_X1 U8360 ( .A1(n7602), .A2(n7600), .ZN(n8362) );
  INV_X1 U8361 ( .A(n6855), .ZN(n7228) );
  NAND3_X1 U8362 ( .A1(n6711), .A2(n7228), .A3(n10159), .ZN(n8363) );
  INV_X1 U8363 ( .A(n6707), .ZN(n6703) );
  INV_X1 U8364 ( .A(n7299), .ZN(n6705) );
  AOI211_X1 U8365 ( .C1(n6707), .C2(n6706), .A(n10010), .B(n6705), .ZN(n6721)
         );
  NAND2_X1 U8366 ( .A1(n6711), .A2(n4247), .ZN(n6708) );
  NAND2_X1 U8367 ( .A1(n8493), .A2(n10058), .ZN(n10038) );
  INV_X1 U8368 ( .A(n10019), .ZN(n8822) );
  NOR2_X1 U8369 ( .A1(n10038), .A2(n8822), .ZN(n6720) );
  NAND2_X1 U8370 ( .A1(n6855), .A2(n6891), .ZN(n8823) );
  NAND2_X1 U8371 ( .A1(n8493), .A2(n10060), .ZN(n10007) );
  INV_X1 U8372 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9676) );
  OAI22_X1 U8373 ( .A1(n10007), .A2(n7350), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9676), .ZN(n6719) );
  NOR2_X1 U8374 ( .A1(n6709), .A2(n8637), .ZN(n6710) );
  INV_X1 U8375 ( .A(n7222), .ZN(n7603) );
  NAND2_X1 U8376 ( .A1(n8362), .A2(n7603), .ZN(n6716) );
  NAND2_X1 U8377 ( .A1(n6716), .A2(n6711), .ZN(n7174) );
  AND2_X1 U8378 ( .A1(n6712), .A2(n6855), .ZN(n7221) );
  INV_X1 U8379 ( .A(n7221), .ZN(n6714) );
  AND3_X1 U8380 ( .A1(n6714), .A2(n6713), .A3(n6856), .ZN(n6715) );
  NAND2_X1 U8381 ( .A1(n6716), .A2(n6715), .ZN(n6717) );
  OAI22_X1 U8382 ( .A1(n8486), .A2(n10138), .B1(n10055), .B2(n7734), .ZN(n6718) );
  OR4_X1 U8383 ( .A1(n6721), .A2(n6720), .A3(n6719), .A4(n6718), .ZN(P2_U3229)
         );
  NAND2_X1 U8384 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_STATE_REG_SCAN_IN), .ZN(
        n6763) );
  OAI21_X1 U8385 ( .B1(n6722), .B2(P1_STATE_REG_SCAN_IN), .A(n6763), .ZN(
        P1_U3353) );
  AND2_X1 U8386 ( .A1(n6728), .A2(P2_U3152), .ZN(n8994) );
  NOR2_X1 U8387 ( .A1(n6728), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8989) );
  OAI222_X1 U8388 ( .A1(n6888), .A2(P2_U3152), .B1(n4249), .B2(n6741), .C1(
        n9633), .C2(n9000), .ZN(P2_U3356) );
  INV_X1 U8389 ( .A(n6942), .ZN(n6953) );
  OAI222_X1 U8390 ( .A1(n9000), .A2(n6723), .B1(n4249), .B2(n6743), .C1(
        P2_U3152), .C2(n6953), .ZN(P2_U3355) );
  INV_X1 U8391 ( .A(n6724), .ZN(n6730) );
  INV_X1 U8392 ( .A(n6916), .ZN(n6927) );
  OAI222_X1 U8393 ( .A1(n9000), .A2(n6725), .B1(n4249), .B2(n6730), .C1(
        P2_U3152), .C2(n6927), .ZN(P2_U3354) );
  INV_X1 U8394 ( .A(n6726), .ZN(n6745) );
  INV_X1 U8395 ( .A(n6928), .ZN(n6941) );
  OAI222_X1 U8396 ( .A1(n9000), .A2(n6727), .B1(n4249), .B2(n6745), .C1(
        P2_U3152), .C2(n6941), .ZN(P2_U3353) );
  NAND2_X1 U8397 ( .A1(n6728), .A2(P1_U3084), .ZN(n9787) );
  INV_X1 U8398 ( .A(n9787), .ZN(n9793) );
  AOI22_X1 U8399 ( .A1(n7063), .A2(P1_STATE_REG_SCAN_IN), .B1(n9793), .B2(
        P2_DATAO_REG_4__SCAN_IN), .ZN(n6729) );
  OAI21_X1 U8400 ( .B1(n6730), .B2(n9798), .A(n6729), .ZN(P1_U3349) );
  INV_X1 U8401 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6732) );
  INV_X1 U8402 ( .A(n6731), .ZN(n6736) );
  INV_X1 U8403 ( .A(n6898), .ZN(n6910) );
  OAI222_X1 U8404 ( .A1(n9000), .A2(n6732), .B1(n4249), .B2(n6736), .C1(
        P2_U3152), .C2(n6910), .ZN(P2_U3352) );
  INV_X1 U8405 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6734) );
  INV_X1 U8406 ( .A(n7097), .ZN(n7283) );
  NAND2_X1 U8407 ( .A1(n7283), .A2(n9777), .ZN(n6733) );
  OAI21_X1 U8408 ( .B1(n9777), .B2(n6734), .A(n6733), .ZN(P1_U3441) );
  AOI22_X1 U8409 ( .A1(n7141), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n9793), .ZN(n6735) );
  OAI21_X1 U8410 ( .B1(n6736), .B2(n9798), .A(n6735), .ZN(P1_U3347) );
  INV_X1 U8411 ( .A(n6737), .ZN(n6739) );
  AOI22_X1 U8412 ( .A1(n9163), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n9793), .ZN(n6738) );
  OAI21_X1 U8413 ( .B1(n6739), .B2(n9798), .A(n6738), .ZN(P1_U3346) );
  INV_X1 U8414 ( .A(n6954), .ZN(n6967) );
  OAI222_X1 U8415 ( .A1(n9000), .A2(n4380), .B1(n4249), .B2(n6739), .C1(
        P2_U3152), .C2(n6967), .ZN(P2_U3351) );
  INV_X1 U8416 ( .A(n7087), .ZN(n6742) );
  OAI222_X1 U8417 ( .A1(n6742), .A2(P1_U3084), .B1(n9798), .B2(n6741), .C1(
        n6740), .C2(n9787), .ZN(P1_U3351) );
  INV_X1 U8418 ( .A(n6795), .ZN(n6973) );
  OAI222_X1 U8419 ( .A1(n9787), .A2(n6744), .B1(n9798), .B2(n6743), .C1(
        P1_U3084), .C2(n6973), .ZN(P1_U3350) );
  OAI222_X1 U8420 ( .A1(n9787), .A2(n6746), .B1(n9798), .B2(n6745), .C1(
        P1_U3084), .C2(n6815), .ZN(P1_U3348) );
  INV_X1 U8421 ( .A(n6747), .ZN(n6749) );
  INV_X1 U8422 ( .A(n7019), .ZN(n7030) );
  OAI222_X1 U8423 ( .A1(n9000), .A2(n6748), .B1(n4249), .B2(n6749), .C1(
        P2_U3152), .C2(n7030), .ZN(P2_U3350) );
  INV_X1 U8424 ( .A(n6822), .ZN(n6847) );
  OAI222_X1 U8425 ( .A1(n9787), .A2(n6750), .B1(n9798), .B2(n6749), .C1(
        P1_U3084), .C2(n6847), .ZN(P1_U3345) );
  OAI21_X1 U8426 ( .B1(n10102), .B2(n7228), .A(n6859), .ZN(n6752) );
  NAND2_X1 U8427 ( .A1(n10102), .A2(n7783), .ZN(n6751) );
  NAND2_X1 U8428 ( .A1(n6752), .A2(n6751), .ZN(n8217) );
  NOR2_X1 U8429 ( .A1(n8587), .A2(P2_U3966), .ZN(P2_U3151) );
  NAND2_X1 U8430 ( .A1(n6479), .A2(P2_U3966), .ZN(n6753) );
  OAI21_X1 U8431 ( .B1(n5142), .B2(P2_U3966), .A(n6753), .ZN(P2_U3552) );
  NAND2_X1 U8432 ( .A1(n9213), .A2(P1_U4006), .ZN(n6754) );
  OAI21_X1 U8433 ( .B1(P1_U4006), .B2(n5060), .A(n6754), .ZN(P1_U3586) );
  MUX2_X1 U8434 ( .A(n6780), .B(n10039), .S(P2_U3966), .Z(n6755) );
  INV_X1 U8435 ( .A(n6755), .ZN(P2_U3562) );
  INV_X1 U8436 ( .A(n6756), .ZN(n6759) );
  INV_X1 U8437 ( .A(n6824), .ZN(n7108) );
  OAI222_X1 U8438 ( .A1(n9787), .A2(n6757), .B1(n9798), .B2(n6759), .C1(n7108), 
        .C2(P1_U3084), .ZN(P1_U3344) );
  INV_X1 U8439 ( .A(n7031), .ZN(n7040) );
  OAI222_X1 U8440 ( .A1(P2_U3152), .A2(n7040), .B1(n4249), .B2(n6759), .C1(
        n6758), .C2(n9000), .ZN(P2_U3349) );
  INV_X1 U8441 ( .A(n6760), .ZN(n7070) );
  INV_X1 U8442 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6776) );
  NOR2_X1 U8443 ( .A1(n7071), .A2(P1_U3084), .ZN(n9789) );
  INV_X1 U8444 ( .A(n9211), .ZN(n6761) );
  NAND2_X1 U8445 ( .A1(n6761), .A2(n7344), .ZN(n6762) );
  NAND2_X1 U8446 ( .A1(n9789), .A2(n6762), .ZN(n6764) );
  NAND2_X1 U8447 ( .A1(n6764), .A2(n6763), .ZN(n7069) );
  AND2_X1 U8448 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(
        n7064) );
  OAI21_X1 U8449 ( .B1(n7064), .B2(n9211), .A(n7195), .ZN(n6768) );
  INV_X1 U8450 ( .A(n6764), .ZN(n6767) );
  NOR2_X1 U8451 ( .A1(n6765), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n6766) );
  AOI22_X1 U8452 ( .A1(n7069), .A2(n6768), .B1(n6767), .B2(n6766), .ZN(n6769)
         );
  NOR2_X1 U8453 ( .A1(n6770), .A2(n6769), .ZN(n6774) );
  AND2_X1 U8454 ( .A1(n9789), .A2(n9211), .ZN(n6771) );
  NOR3_X1 U8455 ( .A1(n9934), .A2(P1_REG1_REG_0__SCAN_IN), .A3(n6772), .ZN(
        n6773) );
  AOI211_X1 U8456 ( .C1(P1_REG3_REG_0__SCAN_IN), .C2(P1_U3084), .A(n6774), .B(
        n6773), .ZN(n6775) );
  OAI21_X1 U8457 ( .B1(n9877), .B2(n6776), .A(n6775), .ZN(P1_U3241) );
  INV_X1 U8458 ( .A(n6777), .ZN(n6837) );
  AOI22_X1 U8459 ( .A1(n9187), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n9793), .ZN(n6778) );
  OAI21_X1 U8460 ( .B1(n6837), .B2(n9798), .A(n6778), .ZN(P1_U3342) );
  INV_X1 U8461 ( .A(n6779), .ZN(n6782) );
  INV_X1 U8462 ( .A(n6993), .ZN(n6831) );
  OAI222_X1 U8463 ( .A1(n9787), .A2(n6780), .B1(n9798), .B2(n6782), .C1(n6831), 
        .C2(P1_U3084), .ZN(P1_U3343) );
  INV_X1 U8464 ( .A(n7153), .ZN(n7147) );
  OAI222_X1 U8465 ( .A1(P2_U3152), .A2(n7147), .B1(n4249), .B2(n6782), .C1(
        n6781), .C2(n9000), .ZN(P2_U3348) );
  INV_X1 U8466 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6805) );
  NOR2_X1 U8467 ( .A1(n9211), .A2(P1_U3084), .ZN(n9792) );
  INV_X1 U8468 ( .A(n6846), .ZN(n9201) );
  NAND2_X1 U8469 ( .A1(n6980), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6784) );
  NAND2_X1 U8470 ( .A1(n6988), .A2(n6784), .ZN(n7082) );
  XNOR2_X1 U8471 ( .A(n7087), .B(n6785), .ZN(n7083) );
  NAND2_X1 U8472 ( .A1(n7082), .A2(n7083), .ZN(n7081) );
  NAND2_X1 U8473 ( .A1(n7087), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6786) );
  NAND2_X1 U8474 ( .A1(n7081), .A2(n6786), .ZN(n6976) );
  XNOR2_X1 U8475 ( .A(n6795), .B(n6787), .ZN(n6977) );
  NAND2_X1 U8476 ( .A1(n6976), .A2(n6977), .ZN(n6975) );
  NAND2_X1 U8477 ( .A1(n6795), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6788) );
  NAND2_X1 U8478 ( .A1(n6975), .A2(n6788), .ZN(n7058) );
  XNOR2_X1 U8479 ( .A(n7063), .B(P1_REG2_REG_4__SCAN_IN), .ZN(n7057) );
  OR2_X1 U8480 ( .A1(n7058), .A2(n7057), .ZN(n7060) );
  OR2_X1 U8481 ( .A1(n7063), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6789) );
  NAND2_X1 U8482 ( .A1(n7060), .A2(n6789), .ZN(n6807) );
  XNOR2_X1 U8483 ( .A(n6815), .B(P1_REG2_REG_5__SCAN_IN), .ZN(n6806) );
  XNOR2_X1 U8484 ( .A(n6807), .B(n6806), .ZN(n6803) );
  NAND2_X1 U8485 ( .A1(n6846), .A2(n7071), .ZN(n9923) );
  AND2_X1 U8486 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7517) );
  INV_X1 U8487 ( .A(n7517), .ZN(n6801) );
  XNOR2_X1 U8488 ( .A(n6815), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n6799) );
  INV_X1 U8489 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n7209) );
  MUX2_X1 U8490 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n7209), .S(n6980), .Z(n6981)
         );
  AND2_X1 U8491 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(
        n6790) );
  NAND2_X1 U8492 ( .A1(n6981), .A2(n6790), .ZN(n6982) );
  NAND2_X1 U8493 ( .A1(n6980), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6791) );
  NAND2_X1 U8494 ( .A1(n6982), .A2(n6791), .ZN(n7077) );
  INV_X1 U8495 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6792) );
  XNOR2_X1 U8496 ( .A(n7087), .B(n6792), .ZN(n7078) );
  NAND2_X1 U8497 ( .A1(n7077), .A2(n7078), .ZN(n7076) );
  NAND2_X1 U8498 ( .A1(n7087), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6793) );
  NAND2_X1 U8499 ( .A1(n7076), .A2(n6793), .ZN(n6969) );
  INV_X1 U8500 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6794) );
  XNOR2_X1 U8501 ( .A(n6795), .B(n6794), .ZN(n6970) );
  NAND2_X1 U8502 ( .A1(n6969), .A2(n6970), .ZN(n6968) );
  NAND2_X1 U8503 ( .A1(n6795), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6796) );
  NAND2_X1 U8504 ( .A1(n6968), .A2(n6796), .ZN(n7053) );
  XNOR2_X1 U8505 ( .A(n7063), .B(P1_REG1_REG_4__SCAN_IN), .ZN(n7054) );
  OR2_X1 U8506 ( .A1(n7063), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6797) );
  AND2_X1 U8507 ( .A1(n7051), .A2(n6797), .ZN(n6798) );
  NAND2_X1 U8508 ( .A1(n6798), .A2(n6799), .ZN(n6818) );
  OAI211_X1 U8509 ( .C1(n6799), .C2(n6798), .A(n9911), .B(n6818), .ZN(n6800)
         );
  OAI211_X1 U8510 ( .C1(n9923), .C2(n6815), .A(n6801), .B(n6800), .ZN(n6802)
         );
  AOI21_X1 U8511 ( .B1(n9929), .B2(n6803), .A(n6802), .ZN(n6804) );
  OAI21_X1 U8512 ( .B1(n9877), .B2(n6805), .A(n6804), .ZN(P1_U3246) );
  NAND2_X1 U8513 ( .A1(n6807), .A2(n6806), .ZN(n6809) );
  NAND2_X1 U8514 ( .A1(n6815), .A2(n7431), .ZN(n6808) );
  NAND2_X1 U8515 ( .A1(n6809), .A2(n6808), .ZN(n7137) );
  XNOR2_X1 U8516 ( .A(n7141), .B(P1_REG2_REG_6__SCAN_IN), .ZN(n7138) );
  NAND2_X1 U8517 ( .A1(n7141), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n6810) );
  XNOR2_X1 U8518 ( .A(n9163), .B(n7484), .ZN(n9170) );
  OAI21_X1 U8519 ( .B1(n7561), .B2(n6847), .A(n6845), .ZN(n6811) );
  NAND2_X1 U8520 ( .A1(n6847), .A2(n7561), .ZN(n6850) );
  NAND2_X1 U8521 ( .A1(n6811), .A2(n6850), .ZN(n7112) );
  MUX2_X1 U8522 ( .A(n7577), .B(P1_REG2_REG_9__SCAN_IN), .S(n6824), .Z(n7111)
         );
  NAND2_X1 U8523 ( .A1(n6824), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6813) );
  MUX2_X1 U8524 ( .A(n7926), .B(P1_REG2_REG_10__SCAN_IN), .S(n6993), .Z(n6812)
         );
  AOI21_X1 U8525 ( .B1(n7109), .B2(n6813), .A(n6812), .ZN(n6992) );
  NAND3_X1 U8526 ( .A1(n7109), .A2(n6813), .A3(n6812), .ZN(n6814) );
  NAND2_X1 U8527 ( .A1(n6814), .A2(n9929), .ZN(n6835) );
  INV_X1 U8528 ( .A(n6815), .ZN(n6816) );
  NAND2_X1 U8529 ( .A1(n6816), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6817) );
  NAND2_X1 U8530 ( .A1(n6818), .A2(n6817), .ZN(n7133) );
  MUX2_X1 U8531 ( .A(n5213), .B(P1_REG1_REG_6__SCAN_IN), .S(n7141), .Z(n7134)
         );
  OR2_X1 U8532 ( .A1(n7141), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n6819) );
  XNOR2_X1 U8533 ( .A(n9163), .B(n6820), .ZN(n9166) );
  NAND2_X1 U8534 ( .A1(n9165), .A2(n9166), .ZN(n9164) );
  OR2_X1 U8535 ( .A1(n9163), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6821) );
  NAND2_X1 U8536 ( .A1(n9164), .A2(n6821), .ZN(n6839) );
  INV_X1 U8537 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10001) );
  OR2_X1 U8538 ( .A1(n6847), .A2(n10001), .ZN(n6838) );
  NOR2_X1 U8539 ( .A1(n6822), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6840) );
  AOI21_X1 U8540 ( .B1(n6839), .B2(n6838), .A(n6840), .ZN(n7105) );
  MUX2_X1 U8541 ( .A(n6823), .B(P1_REG1_REG_9__SCAN_IN), .S(n6824), .Z(n7104)
         );
  NOR2_X1 U8542 ( .A1(n6824), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n6828) );
  INV_X1 U8543 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6825) );
  NAND2_X1 U8544 ( .A1(n6831), .A2(n6825), .ZN(n7001) );
  NAND2_X1 U8545 ( .A1(n6993), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6826) );
  AND2_X1 U8546 ( .A1(n7001), .A2(n6826), .ZN(n6827) );
  INV_X1 U8547 ( .A(n7002), .ZN(n6830) );
  NOR3_X1 U8548 ( .A1(n7103), .A2(n6828), .A3(n6827), .ZN(n6829) );
  OAI21_X1 U8549 ( .B1(n6830), .B2(n6829), .A(n9911), .ZN(n6834) );
  INV_X1 U8550 ( .A(n9877), .ZN(n9927) );
  NAND2_X1 U8551 ( .A1(P1_U3084), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7792) );
  OAI21_X1 U8552 ( .B1(n9923), .B2(n6831), .A(n7792), .ZN(n6832) );
  AOI21_X1 U8553 ( .B1(n9927), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n6832), .ZN(
        n6833) );
  OAI211_X1 U8554 ( .C1(n6992), .C2(n6835), .A(n6834), .B(n6833), .ZN(P1_U3251) );
  INV_X1 U8555 ( .A(n7259), .ZN(n7267) );
  OAI222_X1 U8556 ( .A1(P2_U3152), .A2(n7267), .B1(n4249), .B2(n6837), .C1(
        n6836), .C2(n9000), .ZN(P2_U3347) );
  INV_X1 U8557 ( .A(n6839), .ZN(n6843) );
  INV_X1 U8558 ( .A(n6838), .ZN(n6842) );
  AOI21_X1 U8559 ( .B1(n6840), .B2(n6839), .A(n7105), .ZN(n6841) );
  AOI21_X1 U8560 ( .B1(n6843), .B2(n6842), .A(n6841), .ZN(n6854) );
  NOR2_X1 U8561 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6844), .ZN(n7649) );
  INV_X1 U8562 ( .A(n6845), .ZN(n6851) );
  NAND3_X1 U8563 ( .A1(n6851), .A2(P1_REG2_REG_8__SCAN_IN), .A3(n6846), .ZN(
        n6848) );
  AOI21_X1 U8564 ( .B1(n6848), .B2(n9923), .A(n6847), .ZN(n6849) );
  AOI211_X1 U8565 ( .C1(n9927), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n7649), .B(
        n6849), .ZN(n6853) );
  OAI211_X1 U8566 ( .C1(n6851), .C2(n6850), .A(n7112), .B(n9929), .ZN(n6852)
         );
  OAI211_X1 U8567 ( .C1(n6854), .C2(n9934), .A(n6853), .B(n6852), .ZN(P1_U3249) );
  NOR2_X1 U8568 ( .A1(n10102), .A2(n6855), .ZN(n6858) );
  OR2_X1 U8569 ( .A1(n6891), .A2(P2_U3152), .ZN(n8995) );
  OAI21_X1 U8570 ( .B1(n6856), .B2(n8995), .A(n7783), .ZN(n6857) );
  OR2_X1 U8571 ( .A1(n6858), .A2(n6857), .ZN(n6863) );
  NAND2_X1 U8572 ( .A1(n6863), .A2(n6859), .ZN(n6860) );
  NAND2_X1 U8573 ( .A1(n6860), .A2(n8518), .ZN(n6893) );
  NAND2_X1 U8574 ( .A1(P2_U3152), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n7293) );
  INV_X1 U8575 ( .A(n7293), .ZN(n6885) );
  NOR2_X1 U8576 ( .A1(n6861), .A2(n8223), .ZN(n6862) );
  MUX2_X1 U8577 ( .A(n6864), .B(P2_REG1_REG_2__SCAN_IN), .S(n6888), .Z(n8544)
         );
  MUX2_X1 U8578 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6865), .S(n8527), .Z(n6867)
         );
  AND2_X1 U8579 ( .A1(n9003), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6866) );
  NAND2_X1 U8580 ( .A1(n6867), .A2(n6866), .ZN(n8531) );
  NAND2_X1 U8581 ( .A1(n8527), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6868) );
  NAND2_X1 U8582 ( .A1(n8531), .A2(n6868), .ZN(n8543) );
  NAND2_X1 U8583 ( .A1(n8544), .A2(n8543), .ZN(n8541) );
  NAND2_X1 U8584 ( .A1(n8539), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6943) );
  NAND2_X1 U8585 ( .A1(n8541), .A2(n6943), .ZN(n6871) );
  MUX2_X1 U8586 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6869), .S(n6942), .Z(n6870)
         );
  NAND2_X1 U8587 ( .A1(n6871), .A2(n6870), .ZN(n6946) );
  NAND2_X1 U8588 ( .A1(n6942), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6918) );
  NAND2_X1 U8589 ( .A1(n6946), .A2(n6918), .ZN(n6874) );
  MUX2_X1 U8590 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6872), .S(n6916), .Z(n6873)
         );
  NAND2_X1 U8591 ( .A1(n6874), .A2(n6873), .ZN(n6930) );
  NAND2_X1 U8592 ( .A1(n6916), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6929) );
  NAND2_X1 U8593 ( .A1(n6930), .A2(n6929), .ZN(n6877) );
  MUX2_X1 U8594 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n6875), .S(n6928), .Z(n6876)
         );
  NAND2_X1 U8595 ( .A1(n6877), .A2(n6876), .ZN(n6933) );
  NAND2_X1 U8596 ( .A1(n6928), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n6882) );
  NAND2_X1 U8597 ( .A1(n6933), .A2(n6882), .ZN(n6880) );
  MUX2_X1 U8598 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n6878), .S(n6898), .Z(n6879)
         );
  NAND2_X1 U8599 ( .A1(n6880), .A2(n6879), .ZN(n6957) );
  MUX2_X1 U8600 ( .A(n6878), .B(P2_REG1_REG_6__SCAN_IN), .S(n6898), .Z(n6881)
         );
  NAND3_X1 U8601 ( .A1(n6933), .A2(n6882), .A3(n6881), .ZN(n6883) );
  AND3_X1 U8602 ( .A1(n8542), .A2(n6957), .A3(n6883), .ZN(n6884) );
  AOI211_X1 U8603 ( .C1(n8587), .C2(P2_ADDR_REG_6__SCAN_IN), .A(n6885), .B(
        n6884), .ZN(n6897) );
  XOR2_X1 U8604 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n6898), .Z(n6895) );
  INV_X1 U8605 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n6890) );
  INV_X1 U8606 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7612) );
  XOR2_X1 U8607 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6942), .Z(n6950) );
  INV_X1 U8608 ( .A(n8527), .ZN(n8157) );
  AND2_X1 U8609 ( .A1(n9003), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8525) );
  OAI21_X1 U8610 ( .B1(n6886), .B2(n8157), .A(n8524), .ZN(n8537) );
  XNOR2_X1 U8611 ( .A(n6888), .B(P2_REG2_REG_2__SCAN_IN), .ZN(n8538) );
  NAND2_X1 U8612 ( .A1(n8537), .A2(n8538), .ZN(n8536) );
  OAI21_X1 U8613 ( .B1(n6888), .B2(n6887), .A(n8536), .ZN(n6949) );
  XOR2_X1 U8614 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n6916), .Z(n6924) );
  XOR2_X1 U8615 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n6928), .Z(n6938) );
  OAI21_X1 U8616 ( .B1(n6941), .B2(n6890), .A(n6936), .ZN(n6894) );
  INV_X1 U8617 ( .A(n8223), .ZN(n8998) );
  NOR2_X1 U8618 ( .A1(n8998), .A2(n6891), .ZN(n6892) );
  NAND2_X1 U8619 ( .A1(n6893), .A2(n6892), .ZN(n8564) );
  OAI211_X1 U8620 ( .C1(n6895), .C2(n6894), .A(n8593), .B(n6909), .ZN(n6896)
         );
  OAI211_X1 U8621 ( .C1(n8590), .C2(n6910), .A(n6897), .B(n6896), .ZN(P2_U3251) );
  INV_X1 U8622 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n7465) );
  NOR2_X1 U8623 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7465), .ZN(n6908) );
  NAND2_X1 U8624 ( .A1(n6898), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n6956) );
  NAND2_X1 U8625 ( .A1(n6957), .A2(n6956), .ZN(n6901) );
  MUX2_X1 U8626 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6899), .S(n6954), .Z(n6900)
         );
  NAND2_X1 U8627 ( .A1(n6901), .A2(n6900), .ZN(n6959) );
  NAND2_X1 U8628 ( .A1(n6954), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6905) );
  NAND2_X1 U8629 ( .A1(n6959), .A2(n6905), .ZN(n6903) );
  MUX2_X1 U8630 ( .A(n6223), .B(P2_REG1_REG_8__SCAN_IN), .S(n7019), .Z(n6904)
         );
  INV_X1 U8631 ( .A(n6904), .ZN(n6902) );
  NAND2_X1 U8632 ( .A1(n6903), .A2(n6902), .ZN(n7021) );
  NAND3_X1 U8633 ( .A1(n6959), .A2(n6905), .A3(n6904), .ZN(n6906) );
  AND3_X1 U8634 ( .A1(n8542), .A2(n7021), .A3(n6906), .ZN(n6907) );
  AOI211_X1 U8635 ( .C1(n8587), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n6908), .B(
        n6907), .ZN(n6915) );
  XOR2_X1 U8636 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n7019), .Z(n6913) );
  INV_X1 U8637 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6911) );
  XOR2_X1 U8638 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n6954), .Z(n6964) );
  NAND2_X1 U8639 ( .A1(n6912), .A2(n6913), .ZN(n7028) );
  OAI211_X1 U8640 ( .C1(n6913), .C2(n6912), .A(n8593), .B(n7028), .ZN(n6914)
         );
  OAI211_X1 U8641 ( .C1(n8590), .C2(n7030), .A(n6915), .B(n6914), .ZN(P2_U3253) );
  NAND2_X1 U8642 ( .A1(P2_U3152), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n8430) );
  INV_X1 U8643 ( .A(n8430), .ZN(n6921) );
  MUX2_X1 U8644 ( .A(n6872), .B(P2_REG1_REG_4__SCAN_IN), .S(n6916), .Z(n6917)
         );
  NAND3_X1 U8645 ( .A1(n6946), .A2(n6918), .A3(n6917), .ZN(n6919) );
  AND3_X1 U8646 ( .A1(n8542), .A2(n6930), .A3(n6919), .ZN(n6920) );
  AOI211_X1 U8647 ( .C1(n8587), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n6921), .B(
        n6920), .ZN(n6926) );
  OAI211_X1 U8648 ( .C1(n6924), .C2(n6923), .A(n8593), .B(n6922), .ZN(n6925)
         );
  OAI211_X1 U8649 ( .C1(n8590), .C2(n6927), .A(n6926), .B(n6925), .ZN(P2_U3249) );
  NOR2_X1 U8650 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9676), .ZN(n6935) );
  MUX2_X1 U8651 ( .A(n6875), .B(P2_REG1_REG_5__SCAN_IN), .S(n6928), .Z(n6931)
         );
  NAND3_X1 U8652 ( .A1(n6931), .A2(n6930), .A3(n6929), .ZN(n6932) );
  AND3_X1 U8653 ( .A1(n8542), .A2(n6933), .A3(n6932), .ZN(n6934) );
  AOI211_X1 U8654 ( .C1(n8587), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n6935), .B(
        n6934), .ZN(n6940) );
  OAI211_X1 U8655 ( .C1(n6938), .C2(n6937), .A(n8593), .B(n6936), .ZN(n6939)
         );
  OAI211_X1 U8656 ( .C1(n8590), .C2(n6941), .A(n6940), .B(n6939), .ZN(P2_U3250) );
  AND2_X1 U8657 ( .A1(P2_U3152), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n10018) );
  MUX2_X1 U8658 ( .A(n6869), .B(P2_REG1_REG_3__SCAN_IN), .S(n6942), .Z(n6944)
         );
  NAND3_X1 U8659 ( .A1(n6944), .A2(n8541), .A3(n6943), .ZN(n6945) );
  AND3_X1 U8660 ( .A1(n8542), .A2(n6946), .A3(n6945), .ZN(n6947) );
  AOI211_X1 U8661 ( .C1(n8587), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n10018), .B(
        n6947), .ZN(n6952) );
  OAI211_X1 U8662 ( .C1(n6950), .C2(n6949), .A(n8593), .B(n6948), .ZN(n6951)
         );
  OAI211_X1 U8663 ( .C1(n8590), .C2(n6953), .A(n6952), .B(n6951), .ZN(P2_U3248) );
  NOR2_X1 U8664 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6209), .ZN(n6961) );
  MUX2_X1 U8665 ( .A(n6899), .B(P2_REG1_REG_7__SCAN_IN), .S(n6954), .Z(n6955)
         );
  NAND3_X1 U8666 ( .A1(n6957), .A2(n6956), .A3(n6955), .ZN(n6958) );
  AND3_X1 U8667 ( .A1(n8542), .A2(n6959), .A3(n6958), .ZN(n6960) );
  AOI211_X1 U8668 ( .C1(n8587), .C2(P2_ADDR_REG_7__SCAN_IN), .A(n6961), .B(
        n6960), .ZN(n6966) );
  OAI211_X1 U8669 ( .C1(n6964), .C2(n6963), .A(n8593), .B(n6962), .ZN(n6965)
         );
  OAI211_X1 U8670 ( .C1(n8590), .C2(n6967), .A(n6966), .B(n6965), .ZN(P2_U3252) );
  AND2_X1 U8671 ( .A1(P1_U3084), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n8164) );
  INV_X1 U8672 ( .A(n8164), .ZN(n6972) );
  OAI211_X1 U8673 ( .C1(n6970), .C2(n6969), .A(n9911), .B(n6968), .ZN(n6971)
         );
  OAI211_X1 U8674 ( .C1(n9923), .C2(n6973), .A(n6972), .B(n6971), .ZN(n6974)
         );
  INV_X1 U8675 ( .A(n6974), .ZN(n6979) );
  OAI211_X1 U8676 ( .C1(n6977), .C2(n6976), .A(n9929), .B(n6975), .ZN(n6978)
         );
  OAI211_X1 U8677 ( .C1(n9807), .C2(n9877), .A(n6979), .B(n6978), .ZN(P1_U3244) );
  INV_X1 U8678 ( .A(n6980), .ZN(n8154) );
  NOR2_X1 U8679 ( .A1(n9923), .A2(n8154), .ZN(n6987) );
  NAND2_X1 U8680 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n6985) );
  INV_X1 U8681 ( .A(n6981), .ZN(n6984) );
  INV_X1 U8682 ( .A(n6982), .ZN(n6983) );
  AOI211_X1 U8683 ( .C1(n6985), .C2(n6984), .A(n6983), .B(n9934), .ZN(n6986)
         );
  AOI211_X1 U8684 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(P1_U3084), .A(n6987), .B(
        n6986), .ZN(n6991) );
  OAI211_X1 U8685 ( .C1(n6989), .C2(n7064), .A(n9929), .B(n6988), .ZN(n6990)
         );
  OAI211_X1 U8686 ( .C1(n9668), .C2(n9877), .A(n6991), .B(n6990), .ZN(P1_U3242) );
  MUX2_X1 U8687 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n7727), .S(n9187), .Z(n6995)
         );
  OAI21_X1 U8688 ( .B1(n6995), .B2(n6994), .A(n9177), .ZN(n6999) );
  INV_X1 U8689 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6997) );
  INV_X1 U8690 ( .A(n9923), .ZN(n9886) );
  NAND2_X1 U8691 ( .A1(n9886), .A2(n9187), .ZN(n6996) );
  NAND2_X1 U8692 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7867) );
  OAI211_X1 U8693 ( .C1(n6997), .C2(n9877), .A(n6996), .B(n7867), .ZN(n6998)
         );
  AOI21_X1 U8694 ( .B1(n6999), .B2(n9929), .A(n6998), .ZN(n7007) );
  XNOR2_X1 U8695 ( .A(n9187), .B(n7000), .ZN(n7004) );
  NAND2_X1 U8696 ( .A1(n7002), .A2(n7001), .ZN(n7003) );
  OAI21_X1 U8697 ( .B1(n7004), .B2(n7003), .A(n9186), .ZN(n7005) );
  NAND2_X1 U8698 ( .A1(n7005), .A2(n9911), .ZN(n7006) );
  NAND2_X1 U8699 ( .A1(n7007), .A2(n7006), .ZN(P1_U3252) );
  INV_X1 U8700 ( .A(n7008), .ZN(n7049) );
  AOI22_X1 U8701 ( .A1(n9839), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n9793), .ZN(n7009) );
  OAI21_X1 U8702 ( .B1(n7049), .B2(n9798), .A(n7009), .ZN(P1_U3341) );
  OAI211_X1 U8703 ( .C1(P2_REG1_REG_0__SCAN_IN), .C2(n8584), .A(n8590), .B(
        n9003), .ZN(n7010) );
  AOI21_X1 U8704 ( .B1(n8593), .B2(n6135), .A(n7010), .ZN(n7014) );
  AOI21_X1 U8705 ( .B1(n8542), .B2(P2_REG1_REG_0__SCAN_IN), .A(n9003), .ZN(
        n7013) );
  AOI22_X1 U8706 ( .A1(n8587), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n7012) );
  NAND3_X1 U8707 ( .A1(n7010), .A2(n8593), .A3(P2_REG2_REG_0__SCAN_IN), .ZN(
        n7011) );
  OAI211_X1 U8708 ( .C1(n7014), .C2(n7013), .A(n7012), .B(n7011), .ZN(P2_U3245) );
  INV_X1 U8709 ( .A(n7936), .ZN(n7934) );
  INV_X1 U8710 ( .A(n7015), .ZN(n7017) );
  OAI222_X1 U8711 ( .A1(P2_U3152), .A2(n7934), .B1(n4249), .B2(n7017), .C1(
        n7016), .C2(n9000), .ZN(P2_U3344) );
  INV_X1 U8712 ( .A(n9191), .ZN(n9874) );
  OAI222_X1 U8713 ( .A1(n9787), .A2(n7018), .B1(n9798), .B2(n7017), .C1(n9874), 
        .C2(P1_U3084), .ZN(P1_U3339) );
  NAND2_X1 U8714 ( .A1(n7019), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7020) );
  NAND2_X1 U8715 ( .A1(n7021), .A2(n7020), .ZN(n7039) );
  XNOR2_X1 U8716 ( .A(n7031), .B(n7022), .ZN(n7038) );
  NAND2_X1 U8717 ( .A1(n7039), .A2(n7038), .ZN(n7024) );
  NAND2_X1 U8718 ( .A1(n7031), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7023) );
  NAND2_X1 U8719 ( .A1(n7024), .A2(n7023), .ZN(n7152) );
  XNOR2_X1 U8720 ( .A(n7153), .B(n7025), .ZN(n7151) );
  XNOR2_X1 U8721 ( .A(n7152), .B(n7151), .ZN(n7037) );
  NAND2_X1 U8722 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3152), .ZN(n10005) );
  INV_X1 U8723 ( .A(n10005), .ZN(n7027) );
  NOR2_X1 U8724 ( .A1(n8590), .A2(n7147), .ZN(n7026) );
  AOI211_X1 U8725 ( .C1(n8587), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n7027), .B(
        n7026), .ZN(n7036) );
  INV_X1 U8726 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n7029) );
  MUX2_X1 U8727 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n7032), .S(n7031), .Z(n7044)
         );
  XOR2_X1 U8728 ( .A(n7153), .B(P2_REG2_REG_10__SCAN_IN), .Z(n7033) );
  OAI211_X1 U8729 ( .C1(n7034), .C2(n7033), .A(n7145), .B(n8593), .ZN(n7035)
         );
  OAI211_X1 U8730 ( .C1(n7037), .C2(n8584), .A(n7036), .B(n7035), .ZN(P2_U3255) );
  XNOR2_X1 U8731 ( .A(n7039), .B(n7038), .ZN(n7048) );
  AND2_X1 U8732 ( .A1(P2_U3152), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n7042) );
  NOR2_X1 U8733 ( .A1(n8590), .A2(n7040), .ZN(n7041) );
  AOI211_X1 U8734 ( .C1(n8587), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n7042), .B(
        n7041), .ZN(n7047) );
  OAI211_X1 U8735 ( .C1(n7045), .C2(n7044), .A(n7043), .B(n8593), .ZN(n7046)
         );
  OAI211_X1 U8736 ( .C1(n7048), .C2(n8584), .A(n7047), .B(n7046), .ZN(P2_U3254) );
  INV_X1 U8737 ( .A(n7268), .ZN(n7369) );
  OAI222_X1 U8738 ( .A1(n9000), .A2(n7050), .B1(n4249), .B2(n7049), .C1(
        P2_U3152), .C2(n7369), .ZN(P2_U3346) );
  INV_X1 U8739 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9806) );
  INV_X1 U8740 ( .A(n7051), .ZN(n7052) );
  AOI21_X1 U8741 ( .B1(n7054), .B2(n7053), .A(n7052), .ZN(n7056) );
  INV_X1 U8742 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9662) );
  NOR2_X1 U8743 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9662), .ZN(n8181) );
  INV_X1 U8744 ( .A(n8181), .ZN(n7055) );
  OAI21_X1 U8745 ( .B1(n9934), .B2(n7056), .A(n7055), .ZN(n7062) );
  NAND2_X1 U8746 ( .A1(n7058), .A2(n7057), .ZN(n7059) );
  INV_X1 U8747 ( .A(n9929), .ZN(n9863) );
  AOI21_X1 U8748 ( .B1(n7060), .B2(n7059), .A(n9863), .ZN(n7061) );
  AOI211_X1 U8749 ( .C1(n9886), .C2(n7063), .A(n7062), .B(n7061), .ZN(n7073)
         );
  INV_X1 U8750 ( .A(n7064), .ZN(n7068) );
  OAI21_X1 U8751 ( .B1(n7067), .B2(n7066), .A(n7065), .ZN(n8170) );
  MUX2_X1 U8752 ( .A(n7068), .B(n8170), .S(n9211), .Z(n7072) );
  OAI211_X1 U8753 ( .C1(n7072), .C2(n7071), .A(n7070), .B(n7069), .ZN(n7089)
         );
  OAI211_X1 U8754 ( .C1(n9806), .C2(n9877), .A(n7073), .B(n7089), .ZN(P1_U3245) );
  INV_X1 U8755 ( .A(n7074), .ZN(n7117) );
  AOI22_X1 U8756 ( .A1(n9856), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n9793), .ZN(n7075) );
  OAI21_X1 U8757 ( .B1(n7117), .B2(n9798), .A(n7075), .ZN(P1_U3340) );
  OAI211_X1 U8758 ( .C1(n7078), .C2(n7077), .A(n9911), .B(n7076), .ZN(n7080)
         );
  NAND2_X1 U8759 ( .A1(P1_U3084), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7079) );
  NAND2_X1 U8760 ( .A1(n7080), .A2(n7079), .ZN(n7086) );
  OAI211_X1 U8761 ( .C1(n7083), .C2(n7082), .A(n9929), .B(n7081), .ZN(n7084)
         );
  INV_X1 U8762 ( .A(n7084), .ZN(n7085) );
  AOI211_X1 U8763 ( .C1(n9886), .C2(n7087), .A(n7086), .B(n7085), .ZN(n7088)
         );
  OAI211_X1 U8764 ( .C1(n9808), .C2(n9877), .A(n7089), .B(n7088), .ZN(P1_U3243) );
  INV_X1 U8765 ( .A(n7090), .ZN(n7118) );
  AOI22_X1 U8766 ( .A1(n9885), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n9793), .ZN(n7091) );
  OAI21_X1 U8767 ( .B1(n7118), .B2(n9798), .A(n7091), .ZN(P1_U3338) );
  INV_X1 U8768 ( .A(n7092), .ZN(n7094) );
  OAI21_X1 U8769 ( .B1(n9776), .B2(P1_D_REG_0__SCAN_IN), .A(n9778), .ZN(n7093)
         );
  OAI21_X1 U8770 ( .B1(n7094), .B2(n9776), .A(n7093), .ZN(n7095) );
  NOR2_X1 U8771 ( .A1(n7095), .A2(n7204), .ZN(n7284) );
  OR2_X1 U8772 ( .A1(n9602), .A2(n7189), .ZN(n7098) );
  NAND2_X1 U8773 ( .A1(n7427), .A2(n7329), .ZN(n7099) );
  OAI22_X1 U8774 ( .A1(n7100), .A2(n7099), .B1(n4640), .B2(n9484), .ZN(n7348)
         );
  INV_X1 U8775 ( .A(n7348), .ZN(n7101) );
  OAI21_X1 U8776 ( .B1(n7345), .B2(n7329), .A(n7101), .ZN(n9613) );
  NAND2_X1 U8777 ( .A1(n9613), .A2(n9991), .ZN(n7102) );
  OAI21_X1 U8778 ( .B1(n9991), .B2(n5137), .A(n7102), .ZN(P1_U3454) );
  NAND2_X1 U8779 ( .A1(P1_U3084), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7749) );
  AOI21_X1 U8780 ( .B1(n7105), .B2(n7104), .A(n7103), .ZN(n7106) );
  OR2_X1 U8781 ( .A1(n7106), .A2(n9934), .ZN(n7107) );
  OAI211_X1 U8782 ( .C1(n9923), .C2(n7108), .A(n7749), .B(n7107), .ZN(n7114)
         );
  INV_X1 U8783 ( .A(n7109), .ZN(n7110) );
  AOI211_X1 U8784 ( .C1(n7112), .C2(n7111), .A(n9863), .B(n7110), .ZN(n7113)
         );
  AOI211_X1 U8785 ( .C1(n9927), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n7114), .B(
        n7113), .ZN(n7115) );
  INV_X1 U8786 ( .A(n7115), .ZN(P1_U3250) );
  INV_X1 U8787 ( .A(n7382), .ZN(n7626) );
  OAI222_X1 U8788 ( .A1(P2_U3152), .A2(n7626), .B1(n4249), .B2(n7117), .C1(
        n7116), .C2(n9000), .ZN(P2_U3345) );
  INV_X1 U8789 ( .A(n8188), .ZN(n8195) );
  OAI222_X1 U8790 ( .A1(n9000), .A2(n7119), .B1(n4249), .B2(n7118), .C1(
        P2_U3152), .C2(n8195), .ZN(P2_U3343) );
  OAI21_X1 U8791 ( .B1(n7122), .B2(n7120), .A(n7121), .ZN(n7123) );
  NAND2_X1 U8792 ( .A1(n7123), .A2(n9134), .ZN(n7129) );
  INV_X1 U8793 ( .A(n7166), .ZN(n7125) );
  NAND2_X1 U8794 ( .A1(n7125), .A2(n7124), .ZN(n8172) );
  INV_X1 U8795 ( .A(n9161), .ZN(n7126) );
  OAI22_X1 U8796 ( .A1(n8162), .A2(n9037), .B1(n9139), .B2(n7126), .ZN(n7127)
         );
  AOI21_X1 U8797 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n8172), .A(n7127), .ZN(
        n7128) );
  OAI211_X1 U8798 ( .C1(n7130), .C2(n9145), .A(n7129), .B(n7128), .ZN(P1_U3220) );
  INV_X1 U8799 ( .A(n7131), .ZN(n7132) );
  AOI21_X1 U8800 ( .B1(n7134), .B2(n7133), .A(n7132), .ZN(n7144) );
  NAND2_X1 U8801 ( .A1(P1_U3084), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7588) );
  INV_X1 U8802 ( .A(n7588), .ZN(n7140) );
  INV_X1 U8803 ( .A(n7135), .ZN(n7136) );
  AOI211_X1 U8804 ( .C1(n7138), .C2(n7137), .A(n7136), .B(n9863), .ZN(n7139)
         );
  AOI211_X1 U8805 ( .C1(n9886), .C2(n7141), .A(n7140), .B(n7139), .ZN(n7143)
         );
  NAND2_X1 U8806 ( .A1(n9927), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n7142) );
  OAI211_X1 U8807 ( .C1(n7144), .C2(n9934), .A(n7143), .B(n7142), .ZN(P1_U3247) );
  XNOR2_X1 U8808 ( .A(n7259), .B(P2_REG2_REG_11__SCAN_IN), .ZN(n7149) );
  OAI21_X1 U8809 ( .B1(n7147), .B2(n7146), .A(n7145), .ZN(n7148) );
  AOI21_X1 U8810 ( .B1(n7149), .B2(n7148), .A(n7265), .ZN(n7162) );
  XNOR2_X1 U8811 ( .A(n7259), .B(n7150), .ZN(n7257) );
  NAND2_X1 U8812 ( .A1(n7152), .A2(n7151), .ZN(n7155) );
  NAND2_X1 U8813 ( .A1(n7153), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7154) );
  NAND2_X1 U8814 ( .A1(n7155), .A2(n7154), .ZN(n7258) );
  XOR2_X1 U8815 ( .A(n7257), .B(n7258), .Z(n7160) );
  NOR2_X1 U8816 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7156), .ZN(n7157) );
  AOI21_X1 U8817 ( .B1(n8587), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n7157), .ZN(
        n7158) );
  OAI21_X1 U8818 ( .B1(n8590), .B2(n7267), .A(n7158), .ZN(n7159) );
  AOI21_X1 U8819 ( .B1(n7160), .B2(n8542), .A(n7159), .ZN(n7161) );
  OAI21_X1 U8820 ( .B1(n7162), .B2(n8564), .A(n7161), .ZN(P2_U3256) );
  XOR2_X1 U8821 ( .A(n7164), .B(n7163), .Z(n7169) );
  NAND2_X1 U8822 ( .A1(n9607), .A2(n7443), .ZN(n9947) );
  AOI22_X1 U8823 ( .A1(n9016), .A2(n9160), .B1(n9142), .B2(n9157), .ZN(n7165)
         );
  OAI21_X1 U8824 ( .B1(n7166), .B2(n9947), .A(n7165), .ZN(n7167) );
  AOI21_X1 U8825 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n8172), .A(n7167), .ZN(
        n7168) );
  OAI21_X1 U8826 ( .B1(n7169), .B2(n9132), .A(n7168), .ZN(P1_U3235) );
  INV_X1 U8827 ( .A(n7170), .ZN(n7173) );
  INV_X1 U8828 ( .A(n9185), .ZN(n9895) );
  OAI222_X1 U8829 ( .A1(n9787), .A2(n7171), .B1(n9798), .B2(n7173), .C1(n9895), 
        .C2(P1_U3084), .ZN(P1_U3337) );
  OAI222_X1 U8830 ( .A1(P2_U3152), .A2(n8557), .B1(n4249), .B2(n7173), .C1(
        n7172), .C2(n9000), .ZN(P2_U3342) );
  OR2_X1 U8831 ( .A1(n7174), .A2(n7221), .ZN(n7252) );
  OAI22_X1 U8832 ( .A1(n6134), .A2(n10038), .B1(n10007), .B2(n6127), .ZN(n7175) );
  AOI21_X1 U8833 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(n7252), .A(n7175), .ZN(
        n7181) );
  INV_X1 U8834 ( .A(n7176), .ZN(n10023) );
  AOI211_X1 U8835 ( .C1(n7178), .C2(n7177), .A(n10023), .B(n10010), .ZN(n7179)
         );
  INV_X1 U8836 ( .A(n7179), .ZN(n7180) );
  OAI211_X1 U8837 ( .C1(n7241), .C2(n8486), .A(n7181), .B(n7180), .ZN(P2_U3239) );
  OR2_X1 U8838 ( .A1(n7182), .A2(n7278), .ZN(n7185) );
  OR2_X1 U8839 ( .A1(n7183), .A2(n7624), .ZN(n7184) );
  AND2_X1 U8840 ( .A1(n7185), .A2(n7184), .ZN(n7924) );
  NAND2_X1 U8841 ( .A1(n7924), .A2(n9602), .ZN(n9979) );
  INV_X1 U8842 ( .A(n7345), .ZN(n8171) );
  NAND2_X1 U8843 ( .A1(n9161), .A2(n8171), .ZN(n7186) );
  NAND2_X1 U8844 ( .A1(n7187), .A2(n7186), .ZN(n7307) );
  OAI21_X1 U8845 ( .B1(n7187), .B2(n7186), .A(n7307), .ZN(n7279) );
  INV_X1 U8846 ( .A(n7279), .ZN(n7201) );
  NAND2_X1 U8847 ( .A1(n7188), .A2(n7285), .ZN(n7191) );
  NAND2_X1 U8848 ( .A1(n7189), .A2(n7198), .ZN(n7190) );
  XNOR2_X1 U8849 ( .A(n7193), .B(n7192), .ZN(n7197) );
  INV_X1 U8850 ( .A(n7194), .ZN(n7196) );
  AOI222_X1 U8851 ( .A1(n9454), .A2(n7197), .B1(n9161), .B2(n9451), .C1(n9158), 
        .C2(n9449), .ZN(n7282) );
  NOR2_X1 U8852 ( .A1(n8171), .A2(n7277), .ZN(n7331) );
  INV_X1 U8853 ( .A(n7331), .ZN(n7444) );
  AND2_X1 U8854 ( .A1(n8171), .A2(n7277), .ZN(n7305) );
  NOR2_X1 U8855 ( .A1(n7305), .A2(n9984), .ZN(n7199) );
  AND2_X1 U8856 ( .A1(n7444), .A2(n7199), .ZN(n7287) );
  AOI21_X1 U8857 ( .B1(n9607), .B2(n7277), .A(n7287), .ZN(n7200) );
  OAI211_X1 U8858 ( .C1(n9611), .C2(n7201), .A(n7282), .B(n7200), .ZN(n7207)
         );
  NAND2_X1 U8859 ( .A1(n7207), .A2(n9991), .ZN(n7202) );
  OAI21_X1 U8860 ( .B1(n9991), .B2(n5129), .A(n7202), .ZN(P1_U3457) );
  NOR2_X1 U8861 ( .A1(n7204), .A2(n7203), .ZN(n7205) );
  AND2_X2 U8862 ( .A1(n7206), .A2(n7205), .ZN(n10003) );
  NAND2_X1 U8863 ( .A1(n7207), .A2(n10003), .ZN(n7208) );
  OAI21_X1 U8864 ( .B1(n10003), .B2(n7209), .A(n7208), .ZN(P1_U3524) );
  INV_X1 U8865 ( .A(n7252), .ZN(n7216) );
  INV_X1 U8866 ( .A(n10007), .ZN(n10036) );
  AOI22_X1 U8867 ( .A1(n10029), .A2(n6479), .B1(n10036), .B2(n6673), .ZN(n7215) );
  OAI21_X1 U8868 ( .B1(n7212), .B2(n7211), .A(n7210), .ZN(n7213) );
  AOI22_X1 U8869 ( .A1(n10052), .A2(n6133), .B1(n10043), .B2(n7213), .ZN(n7214) );
  OAI211_X1 U8870 ( .C1(n7216), .C2(n7699), .A(n7215), .B(n7214), .ZN(P2_U3224) );
  INV_X1 U8871 ( .A(n8204), .ZN(n8574) );
  INV_X1 U8872 ( .A(n7217), .ZN(n7219) );
  OAI222_X1 U8873 ( .A1(P2_U3152), .A2(n8574), .B1(n4249), .B2(n7219), .C1(
        n7218), .C2(n9000), .ZN(P2_U3341) );
  INV_X1 U8874 ( .A(n9184), .ZN(n9907) );
  OAI222_X1 U8875 ( .A1(n9787), .A2(n7220), .B1(n9798), .B2(n7219), .C1(n9907), 
        .C2(P1_U3084), .ZN(P1_U3336) );
  NOR2_X1 U8876 ( .A1(n7599), .A2(n7222), .ZN(n7223) );
  AND2_X1 U8877 ( .A1(n7224), .A2(n7223), .ZN(n7225) );
  INV_X1 U8878 ( .A(n7600), .ZN(n7227) );
  INV_X1 U8879 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n7246) );
  NAND2_X1 U8880 ( .A1(n7604), .A2(n7744), .ZN(n7230) );
  AND2_X1 U8881 ( .A1(n7228), .A2(n8637), .ZN(n7229) );
  NAND2_X1 U8882 ( .A1(n7230), .A2(n7229), .ZN(n10157) );
  INV_X1 U8883 ( .A(n8903), .ZN(n10158) );
  NAND2_X1 U8884 ( .A1(n7231), .A2(n7698), .ZN(n7697) );
  OR2_X1 U8885 ( .A1(n6146), .A2(n6133), .ZN(n7232) );
  NAND2_X1 U8886 ( .A1(n7697), .A2(n7232), .ZN(n7233) );
  NAND2_X1 U8887 ( .A1(n7233), .A2(n7234), .ZN(n7596) );
  OAI21_X1 U8888 ( .B1(n7233), .B2(n7234), .A(n7596), .ZN(n8835) );
  INV_X1 U8889 ( .A(n8835), .ZN(n7244) );
  OAI21_X1 U8890 ( .B1(n7239), .B2(n7238), .A(n7237), .ZN(n7240) );
  AOI222_X1 U8891 ( .A1(n10080), .A2(n7240), .B1(n8522), .B2(n10060), .C1(
        n8523), .C2(n10058), .ZN(n8839) );
  INV_X1 U8892 ( .A(n7241), .ZN(n8834) );
  NAND2_X1 U8893 ( .A1(n7508), .A2(n10116), .ZN(n10149) );
  OAI21_X1 U8894 ( .B1(n4890), .B2(n7241), .A(n8950), .ZN(n7242) );
  NOR2_X1 U8895 ( .A1(n7242), .A2(n8826), .ZN(n8837) );
  AOI21_X1 U8896 ( .B1(n8958), .B2(n8834), .A(n8837), .ZN(n7243) );
  OAI211_X1 U8897 ( .C1(n8949), .C2(n7244), .A(n8839), .B(n7243), .ZN(n7248)
         );
  NAND2_X1 U8898 ( .A1(n7248), .A2(n10166), .ZN(n7245) );
  OAI21_X1 U8899 ( .B1(n10166), .B2(n7246), .A(n7245), .ZN(P2_U3457) );
  AND2_X2 U8900 ( .A1(n7247), .A2(n7600), .ZN(n10176) );
  NAND2_X1 U8901 ( .A1(n7248), .A2(n10176), .ZN(n7249) );
  OAI21_X1 U8902 ( .B1(n10176), .B2(n6864), .A(n7249), .ZN(P2_U3522) );
  NAND2_X1 U8903 ( .A1(n10043), .A2(n8310), .ZN(n10026) );
  OAI22_X1 U8904 ( .A1(n10026), .A2(n6145), .B1(n10010), .B2(n7688), .ZN(n7251) );
  AOI22_X1 U8905 ( .A1(n7251), .A2(n7250), .B1(n10052), .B2(n10117), .ZN(n7254) );
  AOI22_X1 U8906 ( .A1(n10036), .A2(n8523), .B1(P2_REG3_REG_0__SCAN_IN), .B2(
        n7252), .ZN(n7253) );
  NAND2_X1 U8907 ( .A1(n7254), .A2(n7253), .ZN(P2_U3234) );
  NAND2_X1 U8908 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n8518), .ZN(n7255) );
  OAI21_X1 U8909 ( .B1(n8608), .B2(n8518), .A(n7255), .ZN(P2_U3579) );
  OR2_X1 U8910 ( .A1(n7268), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7377) );
  NAND2_X1 U8911 ( .A1(n7268), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n7256) );
  NAND2_X1 U8912 ( .A1(n7377), .A2(n7256), .ZN(n7264) );
  NAND2_X1 U8913 ( .A1(n7258), .A2(n7257), .ZN(n7261) );
  NAND2_X1 U8914 ( .A1(n7259), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n7260) );
  NAND2_X1 U8915 ( .A1(n7261), .A2(n7260), .ZN(n7263) );
  INV_X1 U8916 ( .A(n7378), .ZN(n7262) );
  AOI21_X1 U8917 ( .B1(n7264), .B2(n7263), .A(n7262), .ZN(n7275) );
  XOR2_X1 U8918 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7268), .Z(n7269) );
  OAI211_X1 U8919 ( .C1(n7270), .C2(n7269), .A(n7367), .B(n8593), .ZN(n7274)
         );
  NAND2_X1 U8920 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7979) );
  INV_X1 U8921 ( .A(n7979), .ZN(n7272) );
  NOR2_X1 U8922 ( .A1(n8590), .A2(n7369), .ZN(n7271) );
  AOI211_X1 U8923 ( .C1(n8587), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n7272), .B(
        n7271), .ZN(n7273) );
  OAI211_X1 U8924 ( .C1(n7275), .C2(n8584), .A(n7274), .B(n7273), .ZN(P2_U3257) );
  NAND2_X1 U8925 ( .A1(n9777), .A2(n7624), .ZN(n7276) );
  INV_X1 U8926 ( .A(n9460), .ZN(n9472) );
  AOI22_X1 U8927 ( .A1(n9472), .A2(P1_REG3_REG_1__SCAN_IN), .B1(n7333), .B2(
        n7277), .ZN(n7281) );
  AND2_X1 U8928 ( .A1(n7278), .A2(n7285), .ZN(n7327) );
  INV_X1 U8929 ( .A(n7924), .ZN(n7996) );
  OAI21_X1 U8930 ( .B1(n7327), .B2(n7996), .A(n7279), .ZN(n7280) );
  AND3_X1 U8931 ( .A1(n7282), .A2(n7281), .A3(n7280), .ZN(n7289) );
  NAND2_X1 U8932 ( .A1(n7284), .A2(n7283), .ZN(n7286) );
  NOR2_X1 U8933 ( .A1(n7286), .A2(n7285), .ZN(n9410) );
  AOI22_X1 U8934 ( .A1(n9410), .A2(n7287), .B1(n4246), .B2(
        P1_REG2_REG_1__SCAN_IN), .ZN(n7288) );
  OAI21_X1 U8935 ( .B1(n7289), .B2(n4246), .A(n7288), .ZN(P1_U3290) );
  OR2_X1 U8936 ( .A1(n7464), .A2(n8823), .ZN(n7291) );
  NAND2_X1 U8937 ( .A1(n8521), .A2(n10058), .ZN(n7290) );
  NAND2_X1 U8938 ( .A1(n7291), .A2(n7290), .ZN(n10079) );
  NAND2_X1 U8939 ( .A1(n8493), .A2(n10079), .ZN(n7292) );
  OAI211_X1 U8940 ( .C1(n10055), .C2(n10091), .A(n7293), .B(n7292), .ZN(n7296)
         );
  INV_X1 U8941 ( .A(n8521), .ZN(n8431) );
  XNOR2_X1 U8942 ( .A(n10141), .B(n8306), .ZN(n7356) );
  NOR2_X1 U8943 ( .A1(n7350), .A2(n8354), .ZN(n7354) );
  XNOR2_X1 U8944 ( .A(n7356), .B(n7354), .ZN(n7300) );
  NOR4_X1 U8945 ( .A1(n10026), .A2(n8431), .A3(n7294), .A4(n7300), .ZN(n7295)
         );
  AOI211_X1 U8946 ( .C1(n10052), .C2(n10141), .A(n7296), .B(n7295), .ZN(n7303)
         );
  AND2_X1 U8947 ( .A1(n7300), .A2(n7297), .ZN(n7298) );
  OAI21_X1 U8948 ( .B1(n7300), .B2(n7299), .A(n7358), .ZN(n7301) );
  NAND2_X1 U8949 ( .A1(n7301), .A2(n10043), .ZN(n7302) );
  NAND2_X1 U8950 ( .A1(n7303), .A2(n7302), .ZN(P2_U3241) );
  NAND2_X1 U8951 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n8518), .ZN(n7304) );
  OAI21_X1 U8952 ( .B1(n8607), .B2(n8518), .A(n7304), .ZN(P2_U3581) );
  AND2_X1 U8953 ( .A1(n7305), .A2(n9161), .ZN(n7306) );
  AOI21_X1 U8954 ( .B1(n7307), .B2(n9160), .A(n7306), .ZN(n7419) );
  NAND2_X1 U8955 ( .A1(n7419), .A2(n7442), .ZN(n7441) );
  NAND2_X1 U8956 ( .A1(n8162), .A2(n7447), .ZN(n7310) );
  NAND2_X1 U8957 ( .A1(n7441), .A2(n7310), .ZN(n7390) );
  NAND2_X1 U8958 ( .A1(n7390), .A2(n7391), .ZN(n7389) );
  NAND2_X1 U8959 ( .A1(n7308), .A2(n7546), .ZN(n7320) );
  NOR2_X1 U8960 ( .A1(n7320), .A2(n7313), .ZN(n7309) );
  NAND2_X1 U8961 ( .A1(n7389), .A2(n7309), .ZN(n7318) );
  INV_X1 U8962 ( .A(n7313), .ZN(n7311) );
  NAND2_X1 U8963 ( .A1(n7311), .A2(n7310), .ZN(n7420) );
  INV_X1 U8964 ( .A(n7420), .ZN(n7312) );
  NAND2_X1 U8965 ( .A1(n7441), .A2(n7312), .ZN(n7316) );
  NAND2_X1 U8966 ( .A1(n7314), .A2(n7311), .ZN(n7315) );
  NAND2_X1 U8967 ( .A1(n7316), .A2(n7421), .ZN(n7317) );
  NAND2_X1 U8968 ( .A1(n7318), .A2(n7317), .ZN(n9961) );
  NAND2_X1 U8969 ( .A1(n9961), .A2(n7996), .ZN(n7326) );
  OAI22_X1 U8970 ( .A1(n8179), .A2(n9482), .B1(n7532), .B2(n9484), .ZN(n7319)
         );
  INV_X1 U8971 ( .A(n7319), .ZN(n7325) );
  INV_X1 U8972 ( .A(n7546), .ZN(n7322) );
  AOI21_X1 U8973 ( .B1(n7555), .B2(n7320), .A(n9479), .ZN(n7321) );
  OAI21_X1 U8974 ( .B1(n7323), .B2(n7322), .A(n7321), .ZN(n7324) );
  AND3_X1 U8975 ( .A1(n7326), .A2(n7325), .A3(n7324), .ZN(n9963) );
  AND2_X1 U8976 ( .A1(n9463), .A2(n7327), .ZN(n7900) );
  NOR2_X1 U8977 ( .A1(n7329), .A2(n7328), .ZN(n7330) );
  INV_X1 U8978 ( .A(n9491), .ZN(n9369) );
  AND2_X1 U8979 ( .A1(n7396), .A2(n5186), .ZN(n7332) );
  OR2_X1 U8980 ( .A1(n7332), .A2(n7429), .ZN(n9959) );
  INV_X1 U8981 ( .A(n8184), .ZN(n7334) );
  OAI22_X1 U8982 ( .A1(n9463), .A2(n7335), .B1(n7334), .B2(n9460), .ZN(n7336)
         );
  AOI21_X1 U8983 ( .B1(n9365), .B2(n5186), .A(n7336), .ZN(n7337) );
  OAI21_X1 U8984 ( .B1(n9369), .B2(n9959), .A(n7337), .ZN(n7338) );
  AOI21_X1 U8985 ( .B1(n9961), .B2(n7900), .A(n7338), .ZN(n7339) );
  OAI21_X1 U8986 ( .B1(n9963), .B2(n4246), .A(n7339), .ZN(P1_U3287) );
  INV_X1 U8987 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7341) );
  INV_X1 U8988 ( .A(n7340), .ZN(n7342) );
  OAI222_X1 U8989 ( .A1(n9000), .A2(n7341), .B1(n4249), .B2(n7342), .C1(
        P2_U3152), .C2(n4516), .ZN(P2_U3340) );
  INV_X1 U8990 ( .A(n9183), .ZN(n9924) );
  OAI222_X1 U8991 ( .A1(n9787), .A2(n9732), .B1(n9798), .B2(n7342), .C1(
        P1_U3084), .C2(n9924), .ZN(P1_U3335) );
  INV_X1 U8992 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n7343) );
  OAI22_X1 U8993 ( .A1(n9463), .A2(n7344), .B1(n7343), .B2(n9460), .ZN(n7347)
         );
  AOI21_X1 U8994 ( .B1(n9475), .B2(n9369), .A(n7345), .ZN(n7346) );
  AOI211_X1 U8995 ( .C1(n9463), .C2(n7348), .A(n7347), .B(n7346), .ZN(n7349)
         );
  INV_X1 U8996 ( .A(n7349), .ZN(P1_U3291) );
  INV_X1 U8997 ( .A(n7350), .ZN(n10059) );
  OAI22_X1 U8998 ( .A1(n10007), .A2(n7351), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6209), .ZN(n7353) );
  INV_X1 U8999 ( .A(n10072), .ZN(n10148) );
  OAI22_X1 U9000 ( .A1(n8486), .A2(n10148), .B1(n10055), .B2(n10070), .ZN(
        n7352) );
  AOI211_X1 U9001 ( .C1(n10029), .C2(n10059), .A(n7353), .B(n7352), .ZN(n7366)
         );
  INV_X1 U9002 ( .A(n7354), .ZN(n7355) );
  NAND2_X1 U9003 ( .A1(n7356), .A2(n7355), .ZN(n7357) );
  XNOR2_X1 U9004 ( .A(n10072), .B(n8356), .ZN(n7359) );
  NOR2_X1 U9005 ( .A1(n7464), .A2(n8354), .ZN(n7360) );
  NAND2_X1 U9006 ( .A1(n7359), .A2(n7360), .ZN(n7457) );
  INV_X1 U9007 ( .A(n7359), .ZN(n7456) );
  INV_X1 U9008 ( .A(n7360), .ZN(n7361) );
  NAND2_X1 U9009 ( .A1(n7456), .A2(n7361), .ZN(n7362) );
  AND2_X1 U9010 ( .A1(n7457), .A2(n7362), .ZN(n7363) );
  OAI211_X1 U9011 ( .C1(n7364), .C2(n7363), .A(n7458), .B(n10043), .ZN(n7365)
         );
  NAND2_X1 U9012 ( .A1(n7366), .A2(n7365), .ZN(P2_U3215) );
  XNOR2_X1 U9013 ( .A(n7382), .B(P2_REG2_REG_13__SCAN_IN), .ZN(n7371) );
  INV_X1 U9014 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7368) );
  AOI21_X1 U9015 ( .B1(n7371), .B2(n7370), .A(n7625), .ZN(n7384) );
  INV_X1 U9016 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7372) );
  NAND2_X1 U9017 ( .A1(P2_U3152), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n8452) );
  OAI21_X1 U9018 ( .B1(n8217), .B2(n7372), .A(n8452), .ZN(n7381) );
  NAND2_X1 U9019 ( .A1(n7378), .A2(n7377), .ZN(n7375) );
  OR2_X1 U9020 ( .A1(n7382), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7632) );
  NAND2_X1 U9021 ( .A1(n7382), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n7373) );
  NAND2_X1 U9022 ( .A1(n7632), .A2(n7373), .ZN(n7376) );
  INV_X1 U9023 ( .A(n7376), .ZN(n7374) );
  NAND2_X1 U9024 ( .A1(n7375), .A2(n7374), .ZN(n7633) );
  NAND3_X1 U9025 ( .A1(n7378), .A2(n7377), .A3(n7376), .ZN(n7379) );
  AOI21_X1 U9026 ( .B1(n7633), .B2(n7379), .A(n8584), .ZN(n7380) );
  AOI211_X1 U9027 ( .C1(n8540), .C2(n7382), .A(n7381), .B(n7380), .ZN(n7383)
         );
  OAI21_X1 U9028 ( .B1(n7384), .B2(n8564), .A(n7383), .ZN(P2_U3258) );
  INV_X1 U9029 ( .A(n7385), .ZN(n7387) );
  OAI222_X1 U9030 ( .A1(n9787), .A2(n7386), .B1(n9798), .B2(n7387), .C1(n9277), 
        .C2(P1_U3084), .ZN(P1_U3334) );
  OAI222_X1 U9031 ( .A1(n9000), .A2(n7388), .B1(n4249), .B2(n7387), .C1(
        P2_U3152), .C2(n8637), .ZN(P2_U3339) );
  OAI21_X1 U9032 ( .B1(n7390), .B2(n7391), .A(n7389), .ZN(n9956) );
  INV_X1 U9033 ( .A(n9956), .ZN(n7403) );
  INV_X1 U9034 ( .A(n7900), .ZN(n8015) );
  XNOR2_X1 U9035 ( .A(n7392), .B(n7391), .ZN(n7395) );
  NAND2_X1 U9036 ( .A1(n9956), .A2(n7996), .ZN(n7394) );
  AOI22_X1 U9037 ( .A1(n9451), .A2(n9158), .B1(n9156), .B2(n9449), .ZN(n7393)
         );
  OAI211_X1 U9038 ( .C1(n9479), .C2(n7395), .A(n7394), .B(n7393), .ZN(n9954)
         );
  NAND2_X1 U9039 ( .A1(n9954), .A2(n9463), .ZN(n7402) );
  INV_X1 U9040 ( .A(n9944), .ZN(n7397) );
  OAI21_X1 U9041 ( .B1(n7397), .B2(n9952), .A(n7396), .ZN(n9953) );
  AOI22_X1 U9042 ( .A1(n4246), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n9472), .B2(
        n8167), .ZN(n7398) );
  OAI21_X1 U9043 ( .B1(n9369), .B2(n9953), .A(n7398), .ZN(n7399) );
  AOI21_X1 U9044 ( .B1(n9365), .B2(n7400), .A(n7399), .ZN(n7401) );
  OAI211_X1 U9045 ( .C1(n7403), .C2(n8015), .A(n7402), .B(n7401), .ZN(P1_U3288) );
  NAND2_X1 U9046 ( .A1(n7405), .A2(n7404), .ZN(n7586) );
  INV_X1 U9047 ( .A(n7406), .ZN(n7408) );
  NOR3_X1 U9048 ( .A1(n7586), .A2(n7408), .A3(n7407), .ZN(n7411) );
  INV_X1 U9049 ( .A(n7409), .ZN(n7410) );
  OAI21_X1 U9050 ( .B1(n7411), .B2(n7410), .A(n9134), .ZN(n7416) );
  INV_X1 U9051 ( .A(n7483), .ZN(n7414) );
  AND2_X1 U9052 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9162) );
  AOI21_X1 U9053 ( .B1(n9016), .B2(n5830), .A(n9162), .ZN(n7412) );
  OAI21_X1 U9054 ( .B1(n9037), .B2(n7750), .A(n7412), .ZN(n7413) );
  AOI21_X1 U9055 ( .B1(n7414), .B2(n9137), .A(n7413), .ZN(n7415) );
  OAI211_X1 U9056 ( .C1(n7482), .C2(n9145), .A(n7416), .B(n7415), .ZN(P1_U3211) );
  OAI21_X1 U9057 ( .B1(n7474), .B2(n4332), .A(n7417), .ZN(n7418) );
  AOI222_X1 U9058 ( .A1(n9454), .A2(n7418), .B1(n5830), .B2(n9449), .C1(n9156), 
        .C2(n9451), .ZN(n9966) );
  NAND3_X1 U9059 ( .A1(n7421), .A2(n7442), .A3(n7419), .ZN(n7424) );
  NAND2_X1 U9060 ( .A1(n7421), .A2(n7420), .ZN(n7423) );
  OR2_X1 U9061 ( .A1(n5186), .A2(n9156), .ZN(n7422) );
  NAND3_X1 U9062 ( .A1(n7424), .A2(n7423), .A3(n7422), .ZN(n7473) );
  OR2_X1 U9063 ( .A1(n7473), .A2(n7474), .ZN(n7526) );
  INV_X1 U9064 ( .A(n7526), .ZN(n7425) );
  AOI21_X1 U9065 ( .B1(n7474), .B2(n7473), .A(n7425), .ZN(n9969) );
  AND2_X1 U9066 ( .A1(n7427), .A2(n7426), .ZN(n7428) );
  NAND2_X1 U9067 ( .A1(n9463), .A2(n7428), .ZN(n9493) );
  INV_X1 U9068 ( .A(n9493), .ZN(n9467) );
  NOR2_X1 U9069 ( .A1(n7429), .A2(n9964), .ZN(n7430) );
  OR2_X1 U9070 ( .A1(n7533), .A2(n7430), .ZN(n9965) );
  OAI22_X1 U9071 ( .A1(n9463), .A2(n7431), .B1(n7520), .B2(n9460), .ZN(n7432)
         );
  AOI21_X1 U9072 ( .B1(n9365), .B2(n5207), .A(n7432), .ZN(n7433) );
  OAI21_X1 U9073 ( .B1(n9965), .B2(n9369), .A(n7433), .ZN(n7434) );
  AOI21_X1 U9074 ( .B1(n9969), .B2(n9467), .A(n7434), .ZN(n7435) );
  OAI21_X1 U9075 ( .B1(n9966), .B2(n4246), .A(n7435), .ZN(P1_U3286) );
  XNOR2_X1 U9076 ( .A(n7437), .B(n7436), .ZN(n7438) );
  NAND2_X1 U9077 ( .A1(n7438), .A2(n9454), .ZN(n7440) );
  AOI22_X1 U9078 ( .A1(n9157), .A2(n9449), .B1(n9451), .B2(n9160), .ZN(n7439)
         );
  NAND2_X1 U9079 ( .A1(n7440), .A2(n7439), .ZN(n9949) );
  INV_X1 U9080 ( .A(n9949), .ZN(n7450) );
  OAI21_X1 U9081 ( .B1(n7419), .B2(n7442), .A(n7441), .ZN(n9951) );
  AOI22_X1 U9082 ( .A1(n4246), .A2(P1_REG2_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(n9472), .ZN(n7446) );
  NAND2_X1 U9083 ( .A1(n7444), .A2(n7443), .ZN(n9946) );
  NAND3_X1 U9084 ( .A1(n9491), .A2(n9944), .A3(n9946), .ZN(n7445) );
  OAI211_X1 U9085 ( .C1(n9475), .C2(n7447), .A(n7446), .B(n7445), .ZN(n7448)
         );
  AOI21_X1 U9086 ( .B1(n9467), .B2(n9951), .A(n7448), .ZN(n7449) );
  OAI21_X1 U9087 ( .B1(n4246), .B2(n7450), .A(n7449), .ZN(P1_U3289) );
  INV_X1 U9088 ( .A(n7761), .ZN(n10160) );
  XNOR2_X1 U9089 ( .A(n7761), .B(n8356), .ZN(n7493) );
  AND2_X1 U9090 ( .A1(n8310), .A2(n10061), .ZN(n7451) );
  NAND2_X1 U9091 ( .A1(n7493), .A2(n7451), .ZN(n7490) );
  INV_X1 U9092 ( .A(n7493), .ZN(n7453) );
  INV_X1 U9093 ( .A(n7451), .ZN(n7452) );
  NAND2_X1 U9094 ( .A1(n7453), .A2(n7452), .ZN(n7454) );
  AND2_X1 U9095 ( .A1(n7490), .A2(n7454), .ZN(n7459) );
  INV_X1 U9096 ( .A(n7459), .ZN(n7455) );
  AOI21_X1 U9097 ( .B1(n7458), .B2(n7455), .A(n10010), .ZN(n7462) );
  NOR3_X1 U9098 ( .A1(n10026), .A2(n7464), .A3(n7456), .ZN(n7461) );
  OAI21_X1 U9099 ( .B1(n7462), .B2(n7461), .A(n7492), .ZN(n7468) );
  INV_X1 U9100 ( .A(n7463), .ZN(n7665) );
  INV_X1 U9101 ( .A(n7464), .ZN(n8520) );
  AOI22_X1 U9102 ( .A1(n8520), .A2(n10058), .B1(n10060), .B2(n10004), .ZN(
        n7670) );
  OAI22_X1 U9103 ( .A1(n8386), .A2(n7670), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7465), .ZN(n7466) );
  AOI21_X1 U9104 ( .B1(n8505), .B2(n7665), .A(n7466), .ZN(n7467) );
  OAI211_X1 U9105 ( .C1(n10160), .C2(n8486), .A(n7468), .B(n7467), .ZN(
        P2_U3223) );
  INV_X2 U9106 ( .A(P1_U4006), .ZN(n9159) );
  NAND2_X1 U9107 ( .A1(n9159), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n7469) );
  OAI21_X1 U9108 ( .B1(n9287), .B2(n9159), .A(n7469), .ZN(P1_U3584) );
  OAI21_X1 U9109 ( .B1(n4332), .B2(n7547), .A(n7549), .ZN(n7470) );
  XNOR2_X1 U9110 ( .A(n7470), .B(n7550), .ZN(n7471) );
  OAI222_X1 U9111 ( .A1(n9484), .A2(n7750), .B1(n9482), .B2(n7519), .C1(n9479), 
        .C2(n7471), .ZN(n9976) );
  INV_X1 U9112 ( .A(n9976), .ZN(n7489) );
  NAND2_X1 U9113 ( .A1(n9155), .A2(n5207), .ZN(n7525) );
  NAND2_X1 U9114 ( .A1(n7473), .A2(n7472), .ZN(n7478) );
  NAND3_X1 U9115 ( .A1(n7474), .A2(n7529), .A3(n7525), .ZN(n7476) );
  NAND2_X1 U9116 ( .A1(n7519), .A2(n9971), .ZN(n7475) );
  AND2_X1 U9117 ( .A1(n7476), .A2(n7475), .ZN(n7477) );
  NAND2_X1 U9118 ( .A1(n7478), .A2(n7477), .ZN(n7479) );
  INV_X1 U9119 ( .A(n7550), .ZN(n7480) );
  OAI21_X1 U9120 ( .B1(n7479), .B2(n7480), .A(n7542), .ZN(n9978) );
  OAI211_X1 U9121 ( .C1(n4750), .C2(n7482), .A(n9945), .B(n7562), .ZN(n9975)
         );
  INV_X1 U9122 ( .A(n9410), .ZN(n7534) );
  OAI22_X1 U9123 ( .A1(n9463), .A2(n7484), .B1(n7483), .B2(n9460), .ZN(n7485)
         );
  AOI21_X1 U9124 ( .B1(n9365), .B2(n5842), .A(n7485), .ZN(n7486) );
  OAI21_X1 U9125 ( .B1(n9975), .B2(n7534), .A(n7486), .ZN(n7487) );
  AOI21_X1 U9126 ( .B1(n9467), .B2(n9978), .A(n7487), .ZN(n7488) );
  OAI21_X1 U9127 ( .B1(n7489), .B2(n4246), .A(n7488), .ZN(P1_U3284) );
  XNOR2_X1 U9128 ( .A(n8957), .B(n8356), .ZN(n7966) );
  NAND2_X1 U9129 ( .A1(n10004), .A2(n8310), .ZN(n7967) );
  XNOR2_X1 U9130 ( .A(n7966), .B(n7967), .ZN(n7501) );
  AND2_X1 U9131 ( .A1(n7501), .A2(n7490), .ZN(n7491) );
  OAI21_X1 U9132 ( .B1(n7501), .B2(n7492), .A(n7970), .ZN(n7504) );
  INV_X1 U9133 ( .A(n10026), .ZN(n10042) );
  NAND3_X1 U9134 ( .A1(n10042), .A2(n10061), .A3(n7493), .ZN(n7502) );
  INV_X1 U9135 ( .A(n7777), .ZN(n7498) );
  OR2_X1 U9136 ( .A1(n10039), .A2(n8823), .ZN(n7495) );
  NAND2_X1 U9137 ( .A1(n10061), .A2(n10058), .ZN(n7494) );
  AND2_X1 U9138 ( .A1(n7495), .A2(n7494), .ZN(n7771) );
  INV_X1 U9139 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7496) );
  OAI22_X1 U9140 ( .A1(n8386), .A2(n7771), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n7496), .ZN(n7497) );
  AOI21_X1 U9141 ( .B1(n8505), .B2(n7498), .A(n7497), .ZN(n7500) );
  NAND2_X1 U9142 ( .A1(n10052), .A2(n8957), .ZN(n7499) );
  OAI211_X1 U9143 ( .C1(n7502), .C2(n7501), .A(n7500), .B(n7499), .ZN(n7503)
         );
  AOI21_X1 U9144 ( .B1(n7504), .B2(n10043), .A(n7503), .ZN(n7505) );
  INV_X1 U9145 ( .A(n7505), .ZN(P2_U3233) );
  INV_X1 U9146 ( .A(n7506), .ZN(n7641) );
  OAI222_X1 U9147 ( .A1(n7508), .A2(P2_U3152), .B1(n4249), .B2(n7641), .C1(
        n7507), .C2(n9000), .ZN(P2_U3338) );
  NAND2_X1 U9148 ( .A1(n7510), .A2(n7509), .ZN(n7512) );
  INV_X1 U9149 ( .A(n7512), .ZN(n7514) );
  INV_X1 U9150 ( .A(n7511), .ZN(n7513) );
  OR2_X1 U9151 ( .A1(n7512), .A2(n7511), .ZN(n7582) );
  OAI21_X1 U9152 ( .B1(n7514), .B2(n7513), .A(n7582), .ZN(n7515) );
  NOR2_X1 U9153 ( .A1(n7515), .A2(n7516), .ZN(n7585) );
  AOI21_X1 U9154 ( .B1(n7516), .B2(n7515), .A(n7585), .ZN(n7524) );
  AOI21_X1 U9155 ( .B1(n9016), .B2(n9156), .A(n7517), .ZN(n7518) );
  OAI21_X1 U9156 ( .B1(n9037), .B2(n7519), .A(n7518), .ZN(n7522) );
  NOR2_X1 U9157 ( .A1(n9128), .A2(n7520), .ZN(n7521) );
  AOI211_X1 U9158 ( .C1(n9130), .C2(n5207), .A(n7522), .B(n7521), .ZN(n7523)
         );
  OAI21_X1 U9159 ( .B1(n7524), .B2(n9132), .A(n7523), .ZN(P1_U3225) );
  NAND2_X1 U9160 ( .A1(n7526), .A2(n7525), .ZN(n7528) );
  XNOR2_X1 U9161 ( .A(n7528), .B(n7527), .ZN(n9974) );
  INV_X1 U9162 ( .A(n9974), .ZN(n7540) );
  XNOR2_X1 U9163 ( .A(n7530), .B(n7529), .ZN(n7531) );
  OAI222_X1 U9164 ( .A1(n9484), .A2(n7589), .B1(n9482), .B2(n7532), .C1(n7531), 
        .C2(n9479), .ZN(n9972) );
  NAND2_X1 U9165 ( .A1(n9972), .A2(n9463), .ZN(n7539) );
  OAI22_X1 U9166 ( .A1(n9463), .A2(n5208), .B1(n7590), .B2(n9460), .ZN(n7536)
         );
  OAI211_X1 U9167 ( .C1(n7533), .C2(n9971), .A(n9945), .B(n7481), .ZN(n9970)
         );
  NOR2_X1 U9168 ( .A1(n9970), .A2(n7534), .ZN(n7535) );
  AOI211_X1 U9169 ( .C1(n9365), .C2(n7537), .A(n7536), .B(n7535), .ZN(n7538)
         );
  OAI211_X1 U9170 ( .C1(n9493), .C2(n7540), .A(n7539), .B(n7538), .ZN(P1_U3285) );
  OR2_X1 U9171 ( .A1(n5842), .A2(n9154), .ZN(n7541) );
  NAND2_X1 U9172 ( .A1(n7544), .A2(n7557), .ZN(n7545) );
  INV_X1 U9173 ( .A(n9988), .ZN(n7568) );
  NAND2_X1 U9174 ( .A1(n7551), .A2(n7552), .ZN(n7556) );
  NAND2_X1 U9175 ( .A1(n7553), .A2(n7552), .ZN(n7554) );
  NAND2_X1 U9176 ( .A1(n7556), .A2(n4298), .ZN(n7572) );
  XNOR2_X1 U9177 ( .A(n7572), .B(n7557), .ZN(n7560) );
  OAI22_X1 U9178 ( .A1(n7589), .A2(n9482), .B1(n7920), .B2(n9484), .ZN(n7558)
         );
  AOI21_X1 U9179 ( .B1(n9988), .B2(n7996), .A(n7558), .ZN(n7559) );
  OAI21_X1 U9180 ( .B1(n9479), .B2(n7560), .A(n7559), .ZN(n9986) );
  NAND2_X1 U9181 ( .A1(n9986), .A2(n9463), .ZN(n7567) );
  OAI22_X1 U9182 ( .A1(n9463), .A2(n7561), .B1(n7647), .B2(n9460), .ZN(n7565)
         );
  AND2_X1 U9183 ( .A1(n7562), .A2(n9981), .ZN(n7563) );
  OR2_X1 U9184 ( .A1(n7563), .A2(n7578), .ZN(n9985) );
  NOR2_X1 U9185 ( .A1(n9985), .A2(n9369), .ZN(n7564) );
  AOI211_X1 U9186 ( .C1(n9365), .C2(n9981), .A(n7565), .B(n7564), .ZN(n7566)
         );
  OAI211_X1 U9187 ( .C1(n7568), .C2(n8015), .A(n7567), .B(n7566), .ZN(P1_U3283) );
  NAND2_X1 U9188 ( .A1(n9981), .A2(n9153), .ZN(n7569) );
  XNOR2_X1 U9189 ( .A(n7706), .B(n7574), .ZN(n7677) );
  NAND2_X1 U9190 ( .A1(n7718), .A2(n7573), .ZN(n7575) );
  XNOR2_X1 U9191 ( .A(n7575), .B(n7574), .ZN(n7576) );
  AOI222_X1 U9192 ( .A1(n9454), .A2(n7576), .B1(n9153), .B2(n9451), .C1(n9151), 
        .C2(n9449), .ZN(n7676) );
  MUX2_X1 U9193 ( .A(n7577), .B(n7676), .S(n9463), .Z(n7581) );
  AOI21_X1 U9194 ( .B1(n7755), .B2(n4751), .A(n7927), .ZN(n7674) );
  OAI22_X1 U9195 ( .A1(n9475), .A2(n4245), .B1(n9460), .B2(n7753), .ZN(n7579)
         );
  AOI21_X1 U9196 ( .B1(n7674), .B2(n9491), .A(n7579), .ZN(n7580) );
  OAI211_X1 U9197 ( .C1(n7677), .C2(n9493), .A(n7581), .B(n7580), .ZN(P1_U3282) );
  INV_X1 U9198 ( .A(n7582), .ZN(n7583) );
  NOR3_X1 U9199 ( .A1(n7585), .A2(n7584), .A3(n7583), .ZN(n7587) );
  OAI21_X1 U9200 ( .B1(n7587), .B2(n7586), .A(n9134), .ZN(n7594) );
  OAI21_X1 U9201 ( .B1(n9037), .B2(n7589), .A(n7588), .ZN(n7592) );
  NOR2_X1 U9202 ( .A1(n9128), .A2(n7590), .ZN(n7591) );
  AOI211_X1 U9203 ( .C1(n9016), .C2(n9155), .A(n7592), .B(n7591), .ZN(n7593)
         );
  OAI211_X1 U9204 ( .C1(n9971), .C2(n9145), .A(n7594), .B(n7593), .ZN(P1_U3237) );
  OR2_X1 U9205 ( .A1(n6673), .A2(n8834), .ZN(n7595) );
  NAND2_X1 U9206 ( .A1(n8825), .A2(n7597), .ZN(n8824) );
  OR2_X1 U9207 ( .A1(n8522), .A2(n6126), .ZN(n7598) );
  NAND2_X1 U9208 ( .A1(n8824), .A2(n7598), .ZN(n7656) );
  XNOR2_X1 U9209 ( .A(n7656), .B(n7655), .ZN(n10135) );
  INV_X1 U9210 ( .A(n10135), .ZN(n7619) );
  NOR2_X1 U9211 ( .A1(n7600), .A2(n7599), .ZN(n7601) );
  NAND2_X1 U9212 ( .A1(n7602), .A2(n7601), .ZN(n7607) );
  OR2_X1 U9213 ( .A1(n7604), .A2(n8637), .ZN(n7768) );
  AND2_X1 U9214 ( .A1(n10157), .A2(n7768), .ZN(n7605) );
  NOR2_X1 U9215 ( .A1(n7607), .A2(n7606), .ZN(n8838) );
  INV_X1 U9216 ( .A(n8813), .ZN(n10074) );
  NAND2_X1 U9217 ( .A1(n7608), .A2(n10116), .ZN(n7609) );
  NAND2_X1 U9218 ( .A1(n10074), .A2(n8803), .ZN(n7703) );
  XNOR2_X1 U9219 ( .A(n8828), .B(n8434), .ZN(n7611) );
  OAI22_X1 U9220 ( .A1(n7611), .A2(n10149), .B1(n7610), .B2(n10159), .ZN(
        n10134) );
  OAI22_X1 U9221 ( .A1(n10093), .A2(n7612), .B1(n8429), .B2(n10090), .ZN(n7613) );
  AOI21_X1 U9222 ( .B1(n7703), .B2(n10134), .A(n7613), .ZN(n7618) );
  INV_X1 U9223 ( .A(n10058), .ZN(n8821) );
  NAND2_X1 U9224 ( .A1(n8816), .A2(n7614), .ZN(n7615) );
  XNOR2_X1 U9225 ( .A(n7615), .B(n7655), .ZN(n7616) );
  OAI222_X1 U9226 ( .A1(n8823), .A2(n8431), .B1(n8821), .B2(n6127), .C1(n7616), 
        .C2(n8820), .ZN(n10133) );
  NAND2_X1 U9227 ( .A1(n10133), .A2(n10093), .ZN(n7617) );
  OAI211_X1 U9228 ( .C1(n7619), .C2(n8790), .A(n7618), .B(n7617), .ZN(P2_U3292) );
  INV_X1 U9229 ( .A(n7620), .ZN(n7623) );
  OAI222_X1 U9230 ( .A1(n9000), .A2(n7622), .B1(n4249), .B2(n7623), .C1(n7621), 
        .C2(P2_U3152), .ZN(P2_U3337) );
  OAI222_X1 U9231 ( .A1(P1_U3084), .A2(n7624), .B1(n9798), .B2(n7623), .C1(
        n9755), .C2(n9787), .ZN(P1_U3332) );
  MUX2_X1 U9232 ( .A(n7935), .B(P2_REG2_REG_14__SCAN_IN), .S(n7936), .Z(n7628)
         );
  AOI21_X1 U9233 ( .B1(n7628), .B2(n7627), .A(n7933), .ZN(n7639) );
  NOR2_X1 U9234 ( .A1(n7629), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8064) );
  NOR2_X1 U9235 ( .A1(n8217), .A2(n4346), .ZN(n7630) );
  AOI211_X1 U9236 ( .C1(n8540), .C2(n7936), .A(n8064), .B(n7630), .ZN(n7638)
         );
  INV_X1 U9237 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n7631) );
  XNOR2_X1 U9238 ( .A(n7936), .B(n7631), .ZN(n7635) );
  NAND2_X1 U9239 ( .A1(n7633), .A2(n7632), .ZN(n7634) );
  NAND2_X1 U9240 ( .A1(n7634), .A2(n7635), .ZN(n7938) );
  OAI21_X1 U9241 ( .B1(n7635), .B2(n7634), .A(n7938), .ZN(n7636) );
  NAND2_X1 U9242 ( .A1(n7636), .A2(n8542), .ZN(n7637) );
  OAI211_X1 U9243 ( .C1(n7639), .C2(n8564), .A(n7638), .B(n7637), .ZN(P2_U3259) );
  OAI222_X1 U9244 ( .A1(P1_U3084), .A2(n7642), .B1(n9798), .B2(n7641), .C1(
        n7640), .C2(n9787), .ZN(P1_U3333) );
  NAND2_X1 U9245 ( .A1(n7644), .A2(n7643), .ZN(n7645) );
  XOR2_X1 U9246 ( .A(n7646), .B(n7645), .Z(n7654) );
  INV_X1 U9247 ( .A(n7647), .ZN(n7648) );
  NAND2_X1 U9248 ( .A1(n9137), .A2(n7648), .ZN(n7651) );
  AOI21_X1 U9249 ( .B1(n9016), .B2(n9154), .A(n7649), .ZN(n7650) );
  OAI211_X1 U9250 ( .C1(n7920), .C2(n9037), .A(n7651), .B(n7650), .ZN(n7652)
         );
  AOI21_X1 U9251 ( .B1(n9130), .B2(n9981), .A(n7652), .ZN(n7653) );
  OAI21_X1 U9252 ( .B1(n7654), .B2(n9132), .A(n7653), .ZN(P1_U3219) );
  NAND2_X1 U9253 ( .A1(n7656), .A2(n7655), .ZN(n7658) );
  OR2_X1 U9254 ( .A1(n10019), .A2(n8434), .ZN(n7657) );
  NAND2_X1 U9255 ( .A1(n8521), .A2(n7739), .ZN(n10082) );
  NAND2_X1 U9256 ( .A1(n10141), .A2(n10059), .ZN(n7659) );
  AND2_X1 U9257 ( .A1(n10082), .A2(n7659), .ZN(n7663) );
  INV_X1 U9258 ( .A(n7659), .ZN(n7662) );
  OR2_X1 U9259 ( .A1(n7739), .A2(n8521), .ZN(n10084) );
  AND2_X1 U9260 ( .A1(n7660), .A2(n10084), .ZN(n7661) );
  OR2_X2 U9261 ( .A1(n10063), .A2(n10064), .ZN(n10065) );
  OR2_X1 U9262 ( .A1(n10072), .A2(n8520), .ZN(n7664) );
  XNOR2_X1 U9263 ( .A(n7763), .B(n7764), .ZN(n10156) );
  AOI211_X1 U9264 ( .C1(n7761), .C2(n10069), .A(n10149), .B(n7775), .ZN(n10162) );
  INV_X1 U9265 ( .A(n10090), .ZN(n8800) );
  AOI22_X1 U9266 ( .A1(n8836), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n7665), .B2(
        n8800), .ZN(n7666) );
  OAI21_X1 U9267 ( .B1(n8803), .B2(n10160), .A(n7666), .ZN(n7667) );
  AOI21_X1 U9268 ( .B1(n10162), .B2(n8838), .A(n7667), .ZN(n7673) );
  XNOR2_X1 U9269 ( .A(n7669), .B(n7668), .ZN(n7671) );
  OAI21_X1 U9270 ( .B1(n7671), .B2(n8820), .A(n7670), .ZN(n10161) );
  NAND2_X1 U9271 ( .A1(n10161), .A2(n10093), .ZN(n7672) );
  OAI211_X1 U9272 ( .C1(n10156), .C2(n8790), .A(n7673), .B(n7672), .ZN(
        P2_U3288) );
  INV_X1 U9273 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n7679) );
  AOI22_X1 U9274 ( .A1(n7674), .A2(n9945), .B1(n9607), .B2(n7755), .ZN(n7675)
         );
  OAI211_X1 U9275 ( .C1(n9611), .C2(n7677), .A(n7676), .B(n7675), .ZN(n7686)
         );
  NAND2_X1 U9276 ( .A1(n7686), .A2(n9991), .ZN(n7678) );
  OAI21_X1 U9277 ( .B1(n9991), .B2(n7679), .A(n7678), .ZN(P1_U3481) );
  INV_X1 U9278 ( .A(n7703), .ZN(n7685) );
  NAND2_X1 U9279 ( .A1(n6477), .A2(n7680), .ZN(n10118) );
  AOI22_X1 U9280 ( .A1(n10118), .A2(n10080), .B1(n10060), .B2(n8523), .ZN(
        n10120) );
  OAI22_X1 U9281 ( .A1(n8717), .A2(n10120), .B1(n7681), .B2(n10090), .ZN(n7683) );
  NOR2_X1 U9282 ( .A1(n10093), .A2(n6135), .ZN(n7682) );
  AOI211_X1 U9283 ( .C1(n10099), .C2(n10118), .A(n7683), .B(n7682), .ZN(n7684)
         );
  OAI21_X1 U9284 ( .B1(n7685), .B2(n7688), .A(n7684), .ZN(P2_U3296) );
  NAND2_X1 U9285 ( .A1(n7686), .A2(n10003), .ZN(n7687) );
  OAI21_X1 U9286 ( .B1(n10003), .B2(n6823), .A(n7687), .ZN(P1_U3532) );
  OAI21_X1 U9287 ( .B1(n7689), .B2(n7688), .A(n8950), .ZN(n7690) );
  OR2_X1 U9288 ( .A1(n7690), .A2(n4890), .ZN(n7692) );
  NAND2_X1 U9289 ( .A1(n8958), .A2(n6133), .ZN(n7691) );
  NAND2_X1 U9290 ( .A1(n7692), .A2(n7691), .ZN(n10123) );
  INV_X1 U9291 ( .A(n7231), .ZN(n7693) );
  OAI21_X1 U9292 ( .B1(n7693), .B2(n6477), .A(n10080), .ZN(n7696) );
  AOI22_X1 U9293 ( .A1(n10058), .A2(n6479), .B1(n6673), .B2(n10060), .ZN(n7694) );
  OAI21_X1 U9294 ( .B1(n7696), .B2(n7695), .A(n7694), .ZN(n10122) );
  MUX2_X1 U9295 ( .A(n10122), .B(P2_REG2_REG_1__SCAN_IN), .S(n8717), .Z(n7702)
         );
  OAI21_X1 U9296 ( .B1(n7231), .B2(n7698), .A(n7697), .ZN(n10124) );
  INV_X1 U9297 ( .A(n10124), .ZN(n7700) );
  OAI22_X1 U9298 ( .A1(n8790), .A2(n7700), .B1(n7699), .B2(n10090), .ZN(n7701)
         );
  AOI211_X1 U9299 ( .C1(n7703), .C2(n10123), .A(n7702), .B(n7701), .ZN(n7704)
         );
  INV_X1 U9300 ( .A(n7704), .ZN(P2_U3295) );
  AND2_X1 U9301 ( .A1(n7755), .A2(n9152), .ZN(n7705) );
  NAND2_X1 U9302 ( .A1(n7916), .A2(n7919), .ZN(n7707) );
  OR2_X1 U9303 ( .A1(n7709), .A2(n9151), .ZN(n7838) );
  NAND2_X1 U9304 ( .A1(n7707), .A2(n7838), .ZN(n7708) );
  XNOR2_X1 U9305 ( .A(n7708), .B(n7850), .ZN(n9612) );
  NAND2_X1 U9306 ( .A1(n7710), .A2(n7959), .ZN(n7713) );
  NAND2_X1 U9307 ( .A1(n7713), .A2(n9606), .ZN(n7714) );
  AND2_X1 U9308 ( .A1(n8006), .A2(n7714), .ZN(n9608) );
  NAND2_X1 U9309 ( .A1(n9606), .A2(n9365), .ZN(n7715) );
  OAI21_X1 U9310 ( .B1(n9460), .B2(n7868), .A(n7715), .ZN(n7716) );
  AOI21_X1 U9311 ( .B1(n9608), .B2(n9491), .A(n7716), .ZN(n7729) );
  INV_X1 U9312 ( .A(n7719), .ZN(n7720) );
  NAND2_X1 U9313 ( .A1(n7721), .A2(n7848), .ZN(n7723) );
  INV_X1 U9314 ( .A(n7850), .ZN(n7722) );
  XNOR2_X1 U9315 ( .A(n7723), .B(n7722), .ZN(n7726) );
  OAI22_X1 U9316 ( .A1(n7893), .A2(n9484), .B1(n7724), .B2(n9482), .ZN(n7725)
         );
  AOI21_X1 U9317 ( .B1(n7726), .B2(n9454), .A(n7725), .ZN(n9610) );
  MUX2_X1 U9318 ( .A(n7727), .B(n9610), .S(n9463), .Z(n7728) );
  OAI211_X1 U9319 ( .C1(n9612), .C2(n9493), .A(n7729), .B(n7728), .ZN(P1_U3280) );
  NAND2_X1 U9320 ( .A1(n7731), .A2(n7730), .ZN(n7732) );
  XNOR2_X1 U9321 ( .A(n7732), .B(n7740), .ZN(n7733) );
  AOI222_X1 U9322 ( .A1(n10080), .A2(n7733), .B1(n10059), .B2(n10060), .C1(
        n10019), .C2(n10058), .ZN(n10137) );
  OAI22_X1 U9323 ( .A1(n10093), .A2(n6890), .B1(n7734), .B2(n10090), .ZN(n7738) );
  INV_X1 U9324 ( .A(n8838), .ZN(n10097) );
  OAI211_X1 U9325 ( .C1(n7736), .C2(n10138), .A(n7735), .B(n8950), .ZN(n10136)
         );
  NOR2_X1 U9326 ( .A1(n10097), .A2(n10136), .ZN(n7737) );
  AOI211_X1 U9327 ( .C1(n10095), .C2(n7739), .A(n7738), .B(n7737), .ZN(n7742)
         );
  XNOR2_X1 U9328 ( .A(n10083), .B(n7740), .ZN(n10140) );
  NAND2_X1 U9329 ( .A1(n10140), .A2(n10099), .ZN(n7741) );
  OAI211_X1 U9330 ( .C1(n8717), .C2(n10137), .A(n7742), .B(n7741), .ZN(
        P2_U3291) );
  INV_X1 U9331 ( .A(n7743), .ZN(n8158) );
  OAI222_X1 U9332 ( .A1(n9000), .A2(n7745), .B1(n4249), .B2(n8158), .C1(n7744), 
        .C2(P2_U3152), .ZN(P2_U3336) );
  INV_X1 U9333 ( .A(n7788), .ZN(n7746) );
  AOI21_X1 U9334 ( .B1(n7748), .B2(n7747), .A(n7746), .ZN(n7757) );
  OAI21_X1 U9335 ( .B1(n9139), .B2(n7750), .A(n7749), .ZN(n7751) );
  AOI21_X1 U9336 ( .B1(n9142), .B2(n9151), .A(n7751), .ZN(n7752) );
  OAI21_X1 U9337 ( .B1(n7753), .B2(n9128), .A(n7752), .ZN(n7754) );
  AOI21_X1 U9338 ( .B1(n9130), .B2(n7755), .A(n7754), .ZN(n7756) );
  OAI21_X1 U9339 ( .B1(n7757), .B2(n9132), .A(n7756), .ZN(P1_U3229) );
  INV_X1 U9340 ( .A(n7782), .ZN(n7760) );
  AOI21_X1 U9341 ( .B1(P2_DATAO_REG_23__SCAN_IN), .B2(n9793), .A(n7758), .ZN(
        n7759) );
  OAI21_X1 U9342 ( .B1(n7760), .B2(n9798), .A(n7759), .ZN(P1_U3330) );
  NAND2_X1 U9343 ( .A1(n7761), .A2(n10061), .ZN(n7762) );
  INV_X1 U9344 ( .A(n7818), .ZN(n7765) );
  NAND2_X1 U9345 ( .A1(n7765), .A2(n7821), .ZN(n7797) );
  NAND2_X1 U9346 ( .A1(n7818), .A2(n7766), .ZN(n7767) );
  NAND2_X1 U9347 ( .A1(n7797), .A2(n7767), .ZN(n7770) );
  INV_X1 U9348 ( .A(n7770), .ZN(n8961) );
  OR2_X1 U9349 ( .A1(n8717), .A2(n7768), .ZN(n8810) );
  XNOR2_X1 U9350 ( .A(n7769), .B(n7821), .ZN(n7773) );
  INV_X1 U9351 ( .A(n10157), .ZN(n8805) );
  NAND2_X1 U9352 ( .A1(n7770), .A2(n8805), .ZN(n7772) );
  OAI211_X1 U9353 ( .C1(n8820), .C2(n7773), .A(n7772), .B(n7771), .ZN(n8955)
         );
  MUX2_X1 U9354 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n8955), .S(n10093), .Z(n7774)
         );
  INV_X1 U9355 ( .A(n7774), .ZN(n7781) );
  INV_X1 U9356 ( .A(n7775), .ZN(n7776) );
  INV_X1 U9357 ( .A(n8957), .ZN(n7778) );
  AOI211_X1 U9358 ( .C1(n8957), .C2(n7776), .A(n10149), .B(n7803), .ZN(n8956)
         );
  OAI22_X1 U9359 ( .A1(n8803), .A2(n7778), .B1(n7777), .B2(n10090), .ZN(n7779)
         );
  AOI21_X1 U9360 ( .B1(n8956), .B2(n8838), .A(n7779), .ZN(n7780) );
  OAI211_X1 U9361 ( .C1(n8961), .C2(n8810), .A(n7781), .B(n7780), .ZN(P2_U3287) );
  NAND2_X1 U9362 ( .A1(n7782), .A2(n8994), .ZN(n7784) );
  OAI211_X1 U9363 ( .C1(n9750), .C2(n9000), .A(n7784), .B(n7783), .ZN(P2_U3335) );
  XNOR2_X1 U9364 ( .A(n7786), .B(n7785), .ZN(n7790) );
  NAND2_X1 U9365 ( .A1(n7788), .A2(n7787), .ZN(n7789) );
  NAND2_X1 U9366 ( .A1(n7789), .A2(n7790), .ZN(n7864) );
  OAI21_X1 U9367 ( .B1(n7790), .B2(n7789), .A(n7864), .ZN(n7791) );
  NAND2_X1 U9368 ( .A1(n7791), .A2(n9134), .ZN(n7796) );
  OAI21_X1 U9369 ( .B1(n9037), .B2(n7999), .A(n7792), .ZN(n7794) );
  NOR2_X1 U9370 ( .A1(n9128), .A2(n7928), .ZN(n7793) );
  AOI211_X1 U9371 ( .C1(n9016), .C2(n9152), .A(n7794), .B(n7793), .ZN(n7795)
         );
  OAI211_X1 U9372 ( .C1(n7959), .C2(n9145), .A(n7796), .B(n7795), .ZN(P1_U3215) );
  OR2_X1 U9373 ( .A1(n8957), .A2(n10004), .ZN(n7819) );
  NAND2_X1 U9374 ( .A1(n7797), .A2(n7819), .ZN(n7798) );
  XNOR2_X1 U9375 ( .A(n7798), .B(n7823), .ZN(n7809) );
  XNOR2_X1 U9376 ( .A(n7799), .B(n7823), .ZN(n7801) );
  INV_X1 U9377 ( .A(n10008), .ZN(n8519) );
  AOI22_X1 U9378 ( .A1(n8519), .A2(n10060), .B1(n10058), .B2(n10004), .ZN(
        n7800) );
  OAI21_X1 U9379 ( .B1(n7801), .B2(n8820), .A(n7800), .ZN(n7802) );
  AOI21_X1 U9380 ( .B1(n7809), .B2(n8805), .A(n7802), .ZN(n8953) );
  INV_X1 U9381 ( .A(n7803), .ZN(n7805) );
  INV_X1 U9382 ( .A(n10015), .ZN(n7808) );
  INV_X1 U9383 ( .A(n7827), .ZN(n7804) );
  AOI21_X1 U9384 ( .B1(n10015), .B2(n7805), .A(n7804), .ZN(n8951) );
  INV_X1 U9385 ( .A(n10017), .ZN(n7806) );
  AOI22_X1 U9386 ( .A1(n8717), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7806), .B2(
        n8800), .ZN(n7807) );
  OAI21_X1 U9387 ( .B1(n8803), .B2(n7808), .A(n7807), .ZN(n7811) );
  INV_X1 U9388 ( .A(n7809), .ZN(n8954) );
  NOR2_X1 U9389 ( .A1(n8954), .A2(n8810), .ZN(n7810) );
  AOI211_X1 U9390 ( .C1(n8951), .C2(n8813), .A(n7811), .B(n7810), .ZN(n7812)
         );
  OAI21_X1 U9391 ( .B1(n8836), .B2(n8953), .A(n7812), .ZN(P2_U3286) );
  NAND2_X1 U9392 ( .A1(n7814), .A2(n7813), .ZN(n7815) );
  XOR2_X1 U9393 ( .A(n7825), .B(n7815), .Z(n7816) );
  INV_X1 U9394 ( .A(n10039), .ZN(n10040) );
  AOI222_X1 U9395 ( .A1(n10080), .A2(n7816), .B1(n10035), .B2(n10060), .C1(
        n10040), .C2(n10058), .ZN(n8947) );
  OAI21_X1 U9396 ( .B1(n10054), .B2(n10090), .A(n8947), .ZN(n7832) );
  INV_X1 U9397 ( .A(n7819), .ZN(n7820) );
  NOR2_X1 U9398 ( .A1(n7821), .A2(n7820), .ZN(n7822) );
  AOI22_X1 U9399 ( .A1(n7823), .A2(n7822), .B1(n10040), .B2(n10015), .ZN(n7824) );
  OAI21_X1 U9400 ( .B1(n7826), .B2(n7825), .A(n7876), .ZN(n8948) );
  AOI22_X1 U9401 ( .A1(n10095), .A2(n10051), .B1(n8717), .B2(
        P2_REG2_REG_11__SCAN_IN), .ZN(n7830) );
  NAND2_X1 U9402 ( .A1(n7827), .A2(n10051), .ZN(n7828) );
  AND2_X1 U9403 ( .A1(n7881), .A2(n7828), .ZN(n8945) );
  NAND2_X1 U9404 ( .A1(n8945), .A2(n8813), .ZN(n7829) );
  OAI211_X1 U9405 ( .C1(n8948), .C2(n8790), .A(n7830), .B(n7829), .ZN(n7831)
         );
  AOI21_X1 U9406 ( .B1(n7832), .B2(n10093), .A(n7831), .ZN(n7833) );
  INV_X1 U9407 ( .A(n7833), .ZN(P2_U3285) );
  NAND2_X1 U9408 ( .A1(n9606), .A2(n9150), .ZN(n7836) );
  AND2_X1 U9409 ( .A1(n7919), .A2(n7836), .ZN(n7834) );
  NAND2_X1 U9410 ( .A1(n7835), .A2(n7834), .ZN(n7994) );
  INV_X1 U9411 ( .A(n7836), .ZN(n7840) );
  OR2_X1 U9412 ( .A1(n9606), .A2(n9150), .ZN(n7837) );
  AND2_X1 U9413 ( .A1(n7838), .A2(n7837), .ZN(n7839) );
  NAND2_X1 U9414 ( .A1(n7994), .A2(n7841), .ZN(n7843) );
  NAND2_X1 U9415 ( .A1(n9599), .A2(n9149), .ZN(n7842) );
  NAND2_X1 U9416 ( .A1(n9594), .A2(n9148), .ZN(n7844) );
  XNOR2_X1 U9417 ( .A(n8098), .B(n8108), .ZN(n9592) );
  INV_X1 U9418 ( .A(n9590), .ZN(n7846) );
  OR2_X1 U9419 ( .A1(n7896), .A2(n7846), .ZN(n7845) );
  AND3_X1 U9420 ( .A1(n8133), .A2(n9945), .A3(n7845), .ZN(n9589) );
  INV_X1 U9421 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9178) );
  OAI22_X1 U9422 ( .A1(n7846), .A2(n9475), .B1(n9463), .B2(n9178), .ZN(n7847)
         );
  AOI21_X1 U9423 ( .B1(n9589), .B2(n9410), .A(n7847), .ZN(n7861) );
  INV_X1 U9424 ( .A(n7890), .ZN(n7855) );
  XNOR2_X1 U9425 ( .A(n8109), .B(n8108), .ZN(n7858) );
  OAI222_X1 U9426 ( .A1(n9482), .A2(n8125), .B1(n9484), .B2(n9067), .C1(n9479), 
        .C2(n7858), .ZN(n9588) );
  NOR2_X1 U9427 ( .A1(n9460), .A2(n8128), .ZN(n7859) );
  OAI21_X1 U9428 ( .B1(n9588), .B2(n7859), .A(n9463), .ZN(n7860) );
  OAI211_X1 U9429 ( .C1(n9592), .C2(n9493), .A(n7861), .B(n7860), .ZN(P1_U3277) );
  AND2_X1 U9430 ( .A1(n7864), .A2(n7863), .ZN(n7866) );
  XNOR2_X1 U9431 ( .A(n7947), .B(n7862), .ZN(n7865) );
  NAND3_X1 U9432 ( .A1(n7864), .A2(n7865), .A3(n7863), .ZN(n7945) );
  OAI211_X1 U9433 ( .C1(n7866), .C2(n7865), .A(n9134), .B(n7945), .ZN(n7872)
         );
  OAI21_X1 U9434 ( .B1(n9037), .B2(n7893), .A(n7867), .ZN(n7870) );
  NOR2_X1 U9435 ( .A1(n9128), .A2(n7868), .ZN(n7869) );
  AOI211_X1 U9436 ( .C1(n9016), .C2(n9151), .A(n7870), .B(n7869), .ZN(n7871)
         );
  OAI211_X1 U9437 ( .C1(n7711), .C2(n9145), .A(n7872), .B(n7871), .ZN(P1_U3234) );
  XNOR2_X1 U9438 ( .A(n7873), .B(n8024), .ZN(n7874) );
  INV_X1 U9439 ( .A(n8068), .ZN(n8517) );
  AOI222_X1 U9440 ( .A1(n10080), .A2(n7874), .B1(n8519), .B2(n10058), .C1(
        n8517), .C2(n10060), .ZN(n8943) );
  NAND2_X1 U9441 ( .A1(n10051), .A2(n8519), .ZN(n7875) );
  INV_X1 U9442 ( .A(n8036), .ZN(n7877) );
  AOI21_X1 U9443 ( .B1(n7878), .B2(n8022), .A(n7877), .ZN(n8944) );
  NAND2_X1 U9444 ( .A1(n8717), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n7879) );
  OAI21_X1 U9445 ( .B1(n10090), .B2(n7982), .A(n7879), .ZN(n7880) );
  AOI21_X1 U9446 ( .B1(n8941), .B2(n10095), .A(n7880), .ZN(n7885) );
  NAND2_X1 U9447 ( .A1(n8941), .A2(n7881), .ZN(n7882) );
  NAND2_X1 U9448 ( .A1(n7882), .A2(n8950), .ZN(n7883) );
  NOR2_X1 U9449 ( .A1(n8048), .A2(n7883), .ZN(n8940) );
  NAND2_X1 U9450 ( .A1(n8940), .A2(n8838), .ZN(n7884) );
  OAI211_X1 U9451 ( .C1(n8944), .C2(n8790), .A(n7885), .B(n7884), .ZN(n7886)
         );
  INV_X1 U9452 ( .A(n7886), .ZN(n7887) );
  OAI21_X1 U9453 ( .B1(n8836), .B2(n8943), .A(n7887), .ZN(P2_U3284) );
  XOR2_X1 U9454 ( .A(n7888), .B(n7890), .Z(n9593) );
  NAND2_X1 U9455 ( .A1(n7889), .A2(n7890), .ZN(n7891) );
  AOI21_X1 U9456 ( .B1(n7892), .B2(n7891), .A(n9479), .ZN(n7895) );
  OAI22_X1 U9457 ( .A1(n7907), .A2(n9484), .B1(n7893), .B2(n9482), .ZN(n7894)
         );
  AOI211_X1 U9458 ( .C1(n9593), .C2(n7996), .A(n7895), .B(n7894), .ZN(n9597)
         );
  AOI21_X1 U9459 ( .B1(n9594), .B2(n8007), .A(n7896), .ZN(n9595) );
  INV_X1 U9460 ( .A(n9594), .ZN(n7913) );
  NOR2_X1 U9461 ( .A1(n7913), .A2(n9475), .ZN(n7899) );
  INV_X1 U9462 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7897) );
  OAI22_X1 U9463 ( .A1(n9463), .A2(n7897), .B1(n7908), .B2(n9460), .ZN(n7898)
         );
  AOI211_X1 U9464 ( .C1(n9595), .C2(n9491), .A(n7899), .B(n7898), .ZN(n7902)
         );
  NAND2_X1 U9465 ( .A1(n9593), .A2(n7900), .ZN(n7901) );
  OAI211_X1 U9466 ( .C1(n9597), .C2(n4246), .A(n7902), .B(n7901), .ZN(P1_U3278) );
  OAI21_X1 U9467 ( .B1(n7905), .B2(n7904), .A(n7903), .ZN(n7906) );
  NAND2_X1 U9468 ( .A1(n7906), .A2(n9134), .ZN(n7912) );
  NAND2_X1 U9469 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n9859) );
  OAI21_X1 U9470 ( .B1(n9037), .B2(n7907), .A(n9859), .ZN(n7910) );
  NOR2_X1 U9471 ( .A1(n9128), .A2(n7908), .ZN(n7909) );
  AOI211_X1 U9472 ( .C1(n9016), .C2(n9149), .A(n7910), .B(n7909), .ZN(n7911)
         );
  OAI211_X1 U9473 ( .C1(n7913), .C2(n9145), .A(n7912), .B(n7911), .ZN(P1_U3232) );
  INV_X1 U9474 ( .A(n7914), .ZN(n7991) );
  OAI222_X1 U9475 ( .A1(n7915), .A2(P2_U3152), .B1(n4249), .B2(n7991), .C1(
        n9646), .C2(n9000), .ZN(P2_U3334) );
  XOR2_X1 U9476 ( .A(n7916), .B(n7919), .Z(n7957) );
  XOR2_X1 U9477 ( .A(n7919), .B(n7918), .Z(n7922) );
  OAI22_X1 U9478 ( .A1(n7999), .A2(n9484), .B1(n7920), .B2(n9482), .ZN(n7921)
         );
  AOI21_X1 U9479 ( .B1(n7922), .B2(n9454), .A(n7921), .ZN(n7923) );
  OAI21_X1 U9480 ( .B1(n7957), .B2(n7924), .A(n7923), .ZN(n7960) );
  INV_X1 U9481 ( .A(n7960), .ZN(n7925) );
  MUX2_X1 U9482 ( .A(n7926), .B(n7925), .S(n9463), .Z(n7932) );
  OAI211_X1 U9483 ( .C1(n7927), .C2(n7959), .A(n9945), .B(n7713), .ZN(n7958)
         );
  INV_X1 U9484 ( .A(n7958), .ZN(n7930) );
  OAI22_X1 U9485 ( .A1(n7959), .A2(n9475), .B1(n9460), .B2(n7928), .ZN(n7929)
         );
  AOI21_X1 U9486 ( .B1(n7930), .B2(n9410), .A(n7929), .ZN(n7931) );
  OAI211_X1 U9487 ( .C1(n7957), .C2(n8015), .A(n7932), .B(n7931), .ZN(P1_U3281) );
  XNOR2_X1 U9488 ( .A(n8187), .B(n6304), .ZN(n7944) );
  OR2_X1 U9489 ( .A1(n7936), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n7937) );
  NAND2_X1 U9490 ( .A1(n7938), .A2(n7937), .ZN(n8196) );
  XNOR2_X1 U9491 ( .A(n8196), .B(n8188), .ZN(n8194) );
  XOR2_X1 U9492 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8194), .Z(n7942) );
  AND2_X1 U9493 ( .A1(P2_U3152), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n7939) );
  AOI21_X1 U9494 ( .B1(n8587), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n7939), .ZN(
        n7940) );
  OAI21_X1 U9495 ( .B1(n8590), .B2(n8195), .A(n7940), .ZN(n7941) );
  AOI21_X1 U9496 ( .B1(n7942), .B2(n8542), .A(n7941), .ZN(n7943) );
  OAI21_X1 U9497 ( .B1(n7944), .B2(n8564), .A(n7943), .ZN(P2_U3260) );
  OAI21_X1 U9498 ( .B1(n7947), .B2(n7946), .A(n7945), .ZN(n7951) );
  INV_X1 U9499 ( .A(n7948), .ZN(n7949) );
  AOI21_X1 U9500 ( .B1(n7951), .B2(n7950), .A(n7949), .ZN(n7956) );
  NAND2_X1 U9501 ( .A1(P1_U3084), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n9842) );
  OAI21_X1 U9502 ( .B1(n9037), .B2(n8125), .A(n9842), .ZN(n7952) );
  AOI21_X1 U9503 ( .B1(n9016), .B2(n9150), .A(n7952), .ZN(n7953) );
  OAI21_X1 U9504 ( .B1(n8009), .B2(n9128), .A(n7953), .ZN(n7954) );
  AOI21_X1 U9505 ( .B1(n9599), .B2(n9130), .A(n7954), .ZN(n7955) );
  OAI21_X1 U9506 ( .B1(n7956), .B2(n9132), .A(n7955), .ZN(P1_U3222) );
  INV_X1 U9507 ( .A(n9602), .ZN(n9989) );
  INV_X1 U9508 ( .A(n7957), .ZN(n7962) );
  OAI21_X1 U9509 ( .B1(n7959), .B2(n9982), .A(n7958), .ZN(n7961) );
  AOI211_X1 U9510 ( .C1(n9989), .C2(n7962), .A(n7961), .B(n7960), .ZN(n7965)
         );
  NAND2_X1 U9511 ( .A1(n10000), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7963) );
  OAI21_X1 U9512 ( .B1(n7965), .B2(n10000), .A(n7963), .ZN(P1_U3533) );
  NAND2_X1 U9513 ( .A1(n9990), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n7964) );
  OAI21_X1 U9514 ( .B1(n7965), .B2(n9990), .A(n7964), .ZN(P1_U3484) );
  INV_X1 U9515 ( .A(n7966), .ZN(n7968) );
  NAND2_X1 U9516 ( .A1(n7968), .A2(n7967), .ZN(n7969) );
  XNOR2_X1 U9517 ( .A(n10015), .B(n8356), .ZN(n10041) );
  NOR2_X1 U9518 ( .A1(n10039), .A2(n8354), .ZN(n7971) );
  NAND2_X1 U9519 ( .A1(n10041), .A2(n7971), .ZN(n7975) );
  INV_X1 U9520 ( .A(n10041), .ZN(n7973) );
  INV_X1 U9521 ( .A(n7971), .ZN(n7972) );
  NAND2_X1 U9522 ( .A1(n7973), .A2(n7972), .ZN(n7974) );
  NAND2_X1 U9523 ( .A1(n7975), .A2(n7974), .ZN(n10012) );
  NAND2_X1 U9524 ( .A1(n10009), .A2(n7975), .ZN(n7978) );
  XNOR2_X1 U9525 ( .A(n10051), .B(n8356), .ZN(n8076) );
  NOR2_X1 U9526 ( .A1(n10008), .A2(n8354), .ZN(n8075) );
  NAND2_X1 U9527 ( .A1(n8076), .A2(n8075), .ZN(n8070) );
  INV_X1 U9528 ( .A(n8076), .ZN(n7983) );
  INV_X1 U9529 ( .A(n8075), .ZN(n7976) );
  NAND2_X1 U9530 ( .A1(n7983), .A2(n7976), .ZN(n7977) );
  AND2_X1 U9531 ( .A1(n8070), .A2(n7977), .ZN(n10044) );
  NAND2_X1 U9532 ( .A1(n7978), .A2(n10044), .ZN(n8085) );
  XNOR2_X1 U9533 ( .A(n8941), .B(n8356), .ZN(n8072) );
  NAND2_X1 U9534 ( .A1(n10035), .A2(n8310), .ZN(n8073) );
  XNOR2_X1 U9535 ( .A(n8072), .B(n8073), .ZN(n7985) );
  NAND3_X1 U9536 ( .A1(n8085), .A2(n8070), .A3(n7985), .ZN(n8058) );
  OAI21_X1 U9537 ( .B1(n10038), .B2(n10008), .A(n7979), .ZN(n7980) );
  AOI21_X1 U9538 ( .B1(n10036), .B2(n8517), .A(n7980), .ZN(n7981) );
  OAI21_X1 U9539 ( .B1(n7982), .B2(n10055), .A(n7981), .ZN(n7988) );
  INV_X1 U9540 ( .A(n8085), .ZN(n10046) );
  NOR3_X1 U9541 ( .A1(n7983), .A2(n10008), .A3(n10026), .ZN(n7984) );
  AOI21_X1 U9542 ( .B1(n10046), .B2(n10043), .A(n7984), .ZN(n7986) );
  NOR2_X1 U9543 ( .A1(n7986), .A2(n7985), .ZN(n7987) );
  AOI211_X1 U9544 ( .C1(n10052), .C2(n8941), .A(n7988), .B(n7987), .ZN(n7989)
         );
  OAI21_X1 U9545 ( .B1(n10010), .B2(n8058), .A(n7989), .ZN(P2_U3226) );
  OAI222_X1 U9546 ( .A1(P1_U3084), .A2(n7992), .B1(n9798), .B2(n7991), .C1(
        n7990), .C2(n9787), .ZN(P1_U3329) );
  AND2_X1 U9547 ( .A1(n7994), .A2(n7993), .ZN(n7995) );
  XNOR2_X1 U9548 ( .A(n7995), .B(n4444), .ZN(n9603) );
  INV_X1 U9549 ( .A(n9603), .ZN(n7997) );
  NAND2_X1 U9550 ( .A1(n7997), .A2(n7996), .ZN(n8003) );
  XNOR2_X1 U9551 ( .A(n7998), .B(n4444), .ZN(n8001) );
  OAI22_X1 U9552 ( .A1(n8125), .A2(n9484), .B1(n7999), .B2(n9482), .ZN(n8000)
         );
  AOI21_X1 U9553 ( .B1(n8001), .B2(n9454), .A(n8000), .ZN(n8002) );
  NAND2_X1 U9554 ( .A1(n8003), .A2(n8002), .ZN(n9604) );
  INV_X1 U9555 ( .A(n9604), .ZN(n8005) );
  MUX2_X1 U9556 ( .A(n8005), .B(n8004), .S(n4246), .Z(n8014) );
  AOI21_X1 U9557 ( .B1(n8006), .B2(n9599), .A(n9984), .ZN(n8008) );
  NAND2_X1 U9558 ( .A1(n8008), .A2(n8007), .ZN(n9600) );
  INV_X1 U9559 ( .A(n9600), .ZN(n8012) );
  INV_X1 U9560 ( .A(n9599), .ZN(n8010) );
  OAI22_X1 U9561 ( .A1(n8010), .A2(n9475), .B1(n9460), .B2(n8009), .ZN(n8011)
         );
  AOI21_X1 U9562 ( .B1(n8012), .B2(n9410), .A(n8011), .ZN(n8013) );
  OAI211_X1 U9563 ( .C1(n9603), .C2(n8015), .A(n8014), .B(n8013), .ZN(P1_U3279) );
  NAND2_X1 U9564 ( .A1(n8041), .A2(n8042), .ZN(n8040) );
  NAND3_X1 U9565 ( .A1(n8040), .A2(n8028), .A3(n8016), .ZN(n8143) );
  INV_X1 U9566 ( .A(n8143), .ZN(n8018) );
  AOI21_X1 U9567 ( .B1(n8040), .B2(n8016), .A(n8028), .ZN(n8017) );
  NOR3_X1 U9568 ( .A1(n8018), .A2(n8017), .A3(n8820), .ZN(n8020) );
  OAI22_X1 U9569 ( .A1(n8270), .A2(n8823), .B1(n8068), .B2(n8821), .ZN(n8019)
         );
  NOR2_X1 U9570 ( .A1(n8020), .A2(n8019), .ZN(n8932) );
  OR2_X1 U9571 ( .A1(n8941), .A2(n10035), .ZN(n8035) );
  INV_X1 U9572 ( .A(n8035), .ZN(n8023) );
  NOR2_X1 U9573 ( .A1(n8024), .A2(n8023), .ZN(n8025) );
  AOI22_X1 U9574 ( .A1(n8037), .A2(n8025), .B1(n8934), .B2(n8517), .ZN(n8026)
         );
  NOR2_X1 U9575 ( .A1(n8233), .A2(n8028), .ZN(n8149) );
  AOI21_X1 U9576 ( .B1(n8028), .B2(n8233), .A(n8149), .ZN(n8933) );
  INV_X1 U9577 ( .A(n8933), .ZN(n8033) );
  INV_X1 U9578 ( .A(n8934), .ZN(n8052) );
  NAND2_X1 U9579 ( .A1(n8049), .A2(n8929), .ZN(n8029) );
  AND2_X1 U9580 ( .A1(n8147), .A2(n8029), .ZN(n8930) );
  NAND2_X1 U9581 ( .A1(n8930), .A2(n8813), .ZN(n8031) );
  AOI22_X1 U9582 ( .A1(n8836), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n8065), .B2(
        n8800), .ZN(n8030) );
  OAI211_X1 U9583 ( .C1(n4801), .C2(n8803), .A(n8031), .B(n8030), .ZN(n8032)
         );
  AOI21_X1 U9584 ( .B1(n8033), .B2(n10099), .A(n8032), .ZN(n8034) );
  OAI21_X1 U9585 ( .B1(n8836), .B2(n8932), .A(n8034), .ZN(P2_U3282) );
  NAND2_X1 U9586 ( .A1(n8036), .A2(n8035), .ZN(n8038) );
  XNOR2_X1 U9587 ( .A(n8038), .B(n8037), .ZN(n8039) );
  INV_X1 U9588 ( .A(n8039), .ZN(n8937) );
  NAND2_X1 U9589 ( .A1(n8039), .A2(n8805), .ZN(n8047) );
  OAI21_X1 U9590 ( .B1(n8042), .B2(n8041), .A(n8040), .ZN(n8045) );
  NAND2_X1 U9591 ( .A1(n10035), .A2(n10058), .ZN(n8043) );
  OAI21_X1 U9592 ( .B1(n8499), .B2(n8823), .A(n8043), .ZN(n8044) );
  AOI21_X1 U9593 ( .B1(n8045), .B2(n10080), .A(n8044), .ZN(n8046) );
  NAND2_X1 U9594 ( .A1(n8047), .A2(n8046), .ZN(n8939) );
  NAND2_X1 U9595 ( .A1(n8939), .A2(n10093), .ZN(n8056) );
  OR2_X1 U9596 ( .A1(n8052), .A2(n8048), .ZN(n8050) );
  AND2_X1 U9597 ( .A1(n8050), .A2(n8049), .ZN(n8935) );
  OAI22_X1 U9598 ( .A1(n10093), .A2(n8051), .B1(n8455), .B2(n10090), .ZN(n8054) );
  NOR2_X1 U9599 ( .A1(n8052), .A2(n8803), .ZN(n8053) );
  AOI211_X1 U9600 ( .C1(n8935), .C2(n8813), .A(n8054), .B(n8053), .ZN(n8055)
         );
  OAI211_X1 U9601 ( .C1(n8937), .C2(n8810), .A(n8056), .B(n8055), .ZN(P2_U3283) );
  INV_X1 U9602 ( .A(n8072), .ZN(n8057) );
  NAND2_X1 U9603 ( .A1(n8057), .A2(n8073), .ZN(n8069) );
  NAND2_X1 U9604 ( .A1(n8058), .A2(n8069), .ZN(n8457) );
  XNOR2_X1 U9605 ( .A(n8934), .B(n8306), .ZN(n8062) );
  OR2_X1 U9606 ( .A1(n8068), .A2(n8354), .ZN(n8059) );
  NAND2_X1 U9607 ( .A1(n8062), .A2(n8059), .ZN(n8080) );
  INV_X1 U9608 ( .A(n8062), .ZN(n8061) );
  INV_X1 U9609 ( .A(n8059), .ZN(n8060) );
  NAND2_X1 U9610 ( .A1(n8061), .A2(n8060), .ZN(n8081) );
  NAND2_X1 U9611 ( .A1(n8080), .A2(n8081), .ZN(n8458) );
  NOR2_X1 U9612 ( .A1(n8457), .A2(n8458), .ZN(n8456) );
  NOR3_X1 U9613 ( .A1(n8062), .A2(n8068), .A3(n10026), .ZN(n8063) );
  AOI21_X1 U9614 ( .B1(n8456), .B2(n10043), .A(n8063), .ZN(n8090) );
  XNOR2_X1 U9615 ( .A(n8929), .B(n8306), .ZN(n8267) );
  NOR2_X1 U9616 ( .A1(n8499), .A2(n8354), .ZN(n8265) );
  XNOR2_X1 U9617 ( .A(n8267), .B(n8265), .ZN(n8089) );
  INV_X1 U9618 ( .A(n8270), .ZN(n8794) );
  AOI21_X1 U9619 ( .B1(n10036), .B2(n8794), .A(n8064), .ZN(n8067) );
  NAND2_X1 U9620 ( .A1(n8505), .A2(n8065), .ZN(n8066) );
  OAI211_X1 U9621 ( .C1(n8068), .C2(n10038), .A(n8067), .B(n8066), .ZN(n8087)
         );
  NAND2_X1 U9622 ( .A1(n8080), .A2(n8069), .ZN(n8084) );
  NAND2_X1 U9623 ( .A1(n8070), .A2(n8073), .ZN(n8071) );
  NAND2_X1 U9624 ( .A1(n8072), .A2(n8071), .ZN(n8078) );
  INV_X1 U9625 ( .A(n8073), .ZN(n8074) );
  NAND3_X1 U9626 ( .A1(n8076), .A2(n8075), .A3(n8074), .ZN(n8077) );
  NAND2_X1 U9627 ( .A1(n8078), .A2(n8077), .ZN(n8079) );
  NAND2_X1 U9628 ( .A1(n8080), .A2(n8079), .ZN(n8082) );
  AND3_X1 U9629 ( .A1(n8082), .A2(n8089), .A3(n8081), .ZN(n8083) );
  NOR2_X1 U9630 ( .A1(n8269), .A2(n10010), .ZN(n8086) );
  AOI211_X1 U9631 ( .C1(n10052), .C2(n8929), .A(n8087), .B(n8086), .ZN(n8088)
         );
  OAI21_X1 U9632 ( .B1(n8090), .B2(n8089), .A(n8088), .ZN(P2_U3217) );
  INV_X1 U9633 ( .A(n8091), .ZN(n8095) );
  OAI222_X1 U9634 ( .A1(n9000), .A2(n8093), .B1(n4249), .B2(n8095), .C1(n8092), 
        .C2(P2_U3152), .ZN(P2_U3333) );
  OAI222_X1 U9635 ( .A1(n9787), .A2(n8096), .B1(n9798), .B2(n8095), .C1(
        P1_U3084), .C2(n8094), .ZN(P1_U3328) );
  AND2_X1 U9636 ( .A1(n9590), .A2(n9147), .ZN(n8097) );
  NOR2_X1 U9637 ( .A1(n9583), .A2(n9146), .ZN(n8099) );
  NAND2_X1 U9638 ( .A1(n9583), .A2(n9146), .ZN(n8100) );
  XNOR2_X1 U9639 ( .A(n9222), .B(n9221), .ZN(n9582) );
  NAND2_X1 U9640 ( .A1(n4756), .A2(n9580), .ZN(n8102) );
  NAND2_X1 U9641 ( .A1(n8102), .A2(n9945), .ZN(n8103) );
  NOR2_X1 U9642 ( .A1(n9208), .A2(n8103), .ZN(n9579) );
  INV_X1 U9643 ( .A(n9580), .ZN(n8104) );
  NOR2_X1 U9644 ( .A1(n8104), .A2(n9475), .ZN(n8106) );
  INV_X1 U9645 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n9640) );
  OAI22_X1 U9646 ( .A1(n9463), .A2(n9640), .B1(n9070), .B2(n9460), .ZN(n8105)
         );
  AOI211_X1 U9647 ( .C1(n9579), .C2(n9410), .A(n8106), .B(n8105), .ZN(n8113)
         );
  XNOR2_X1 U9648 ( .A(n9246), .B(n9221), .ZN(n8111) );
  OAI222_X1 U9649 ( .A1(n9484), .A2(n9125), .B1(n9482), .B2(n9067), .C1(n8111), 
        .C2(n9479), .ZN(n9578) );
  NAND2_X1 U9650 ( .A1(n9578), .A2(n9463), .ZN(n8112) );
  OAI211_X1 U9651 ( .C1(n9582), .C2(n9493), .A(n8113), .B(n8112), .ZN(P1_U3275) );
  INV_X1 U9652 ( .A(n9059), .ZN(n9057) );
  XNOR2_X1 U9653 ( .A(n9057), .B(n9061), .ZN(n8114) );
  XNOR2_X1 U9654 ( .A(n9058), .B(n8114), .ZN(n8120) );
  NAND2_X1 U9655 ( .A1(n9137), .A2(n8134), .ZN(n8117) );
  NOR2_X1 U9656 ( .A1(n8115), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9884) );
  AOI21_X1 U9657 ( .B1(n9016), .B2(n9147), .A(n9884), .ZN(n8116) );
  OAI211_X1 U9658 ( .C1(n9483), .C2(n9037), .A(n8117), .B(n8116), .ZN(n8118)
         );
  AOI21_X1 U9659 ( .B1(n9583), .B2(n9130), .A(n8118), .ZN(n8119) );
  OAI21_X1 U9660 ( .B1(n8120), .B2(n9132), .A(n8119), .ZN(P1_U3239) );
  NAND2_X1 U9661 ( .A1(n8122), .A2(n8121), .ZN(n8123) );
  XOR2_X1 U9662 ( .A(n8124), .B(n8123), .Z(n8131) );
  NAND2_X1 U9663 ( .A1(P1_U3084), .A2(P1_REG3_REG_14__SCAN_IN), .ZN(n9876) );
  OAI21_X1 U9664 ( .B1(n9139), .B2(n8125), .A(n9876), .ZN(n8126) );
  AOI21_X1 U9665 ( .B1(n9142), .B2(n9146), .A(n8126), .ZN(n8127) );
  OAI21_X1 U9666 ( .B1(n8128), .B2(n9128), .A(n8127), .ZN(n8129) );
  AOI21_X1 U9667 ( .B1(n9590), .B2(n9130), .A(n8129), .ZN(n8130) );
  OAI21_X1 U9668 ( .B1(n8131), .B2(n9132), .A(n8130), .ZN(P1_U3213) );
  XNOR2_X1 U9669 ( .A(n8132), .B(n4268), .ZN(n9587) );
  AOI21_X1 U9670 ( .B1(n9583), .B2(n8133), .A(n8101), .ZN(n9584) );
  AOI22_X1 U9671 ( .A1(n4246), .A2(P1_REG2_REG_15__SCAN_IN), .B1(n8134), .B2(
        n9472), .ZN(n8135) );
  OAI21_X1 U9672 ( .B1(n4753), .B2(n9475), .A(n8135), .ZN(n8140) );
  OAI21_X1 U9673 ( .B1(n8137), .B2(n4268), .A(n8136), .ZN(n8138) );
  AOI222_X1 U9674 ( .A1(n9454), .A2(n8138), .B1(n9147), .B2(n9451), .C1(n9223), 
        .C2(n9449), .ZN(n9586) );
  NOR2_X1 U9675 ( .A1(n9586), .A2(n4246), .ZN(n8139) );
  AOI211_X1 U9676 ( .C1(n9584), .C2(n9491), .A(n8140), .B(n8139), .ZN(n8141)
         );
  OAI21_X1 U9677 ( .B1(n9587), .B2(n9493), .A(n8141), .ZN(P1_U3276) );
  NAND2_X1 U9678 ( .A1(n8143), .A2(n8142), .ZN(n8144) );
  XNOR2_X1 U9679 ( .A(n8144), .B(n8231), .ZN(n8145) );
  INV_X1 U9680 ( .A(n8501), .ZN(n8515) );
  INV_X1 U9681 ( .A(n8499), .ZN(n8516) );
  AOI222_X1 U9682 ( .A1(n10080), .A2(n8145), .B1(n8515), .B2(n10060), .C1(
        n8516), .C2(n10058), .ZN(n8927) );
  INV_X1 U9683 ( .A(n8798), .ZN(n8146) );
  AOI21_X1 U9684 ( .B1(n8924), .B2(n8147), .A(n8146), .ZN(n8925) );
  AOI22_X1 U9685 ( .A1(n8717), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8504), .B2(
        n8800), .ZN(n8148) );
  OAI21_X1 U9686 ( .B1(n4477), .B2(n8803), .A(n8148), .ZN(n8152) );
  NOR2_X1 U9687 ( .A1(n8929), .A2(n8516), .ZN(n8230) );
  NOR2_X1 U9688 ( .A1(n8149), .A2(n8230), .ZN(n8150) );
  XNOR2_X1 U9689 ( .A(n8150), .B(n8231), .ZN(n8928) );
  NOR2_X1 U9690 ( .A1(n8928), .A2(n8790), .ZN(n8151) );
  AOI211_X1 U9691 ( .C1(n8925), .C2(n8813), .A(n8152), .B(n8151), .ZN(n8153)
         );
  OAI21_X1 U9692 ( .B1(n8836), .B2(n8927), .A(n8153), .ZN(P2_U3281) );
  INV_X1 U9693 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n9637) );
  OAI222_X1 U9694 ( .A1(P1_U3084), .A2(n8154), .B1(n9798), .B2(n8156), .C1(
        n9637), .C2(n9787), .ZN(P1_U3352) );
  INV_X1 U9695 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8155) );
  OAI222_X1 U9696 ( .A1(n8157), .A2(P2_U3152), .B1(n4249), .B2(n8156), .C1(
        n8155), .C2(n9000), .ZN(P2_U3357) );
  OAI222_X1 U9697 ( .A1(n9787), .A2(n8159), .B1(n9798), .B2(n8158), .C1(n5784), 
        .C2(P1_U3084), .ZN(P1_U3331) );
  XOR2_X1 U9698 ( .A(n8161), .B(n8160), .Z(n8169) );
  NOR2_X1 U9699 ( .A1(n9139), .A2(n8162), .ZN(n8163) );
  AOI211_X1 U9700 ( .C1(n9142), .C2(n9156), .A(n8164), .B(n8163), .ZN(n8165)
         );
  OAI21_X1 U9701 ( .B1(n9952), .B2(n9145), .A(n8165), .ZN(n8166) );
  AOI21_X1 U9702 ( .B1(n9137), .B2(n8167), .A(n8166), .ZN(n8168) );
  OAI21_X1 U9703 ( .B1(n8169), .B2(n9132), .A(n8168), .ZN(P1_U3216) );
  AOI22_X1 U9704 ( .A1(n9130), .A2(n8171), .B1(n8170), .B2(n9134), .ZN(n8174)
         );
  AOI22_X1 U9705 ( .A1(n8172), .A2(P1_REG3_REG_0__SCAN_IN), .B1(n9142), .B2(
        n9160), .ZN(n8173) );
  NAND2_X1 U9706 ( .A1(n8174), .A2(n8173), .ZN(P1_U3230) );
  XNOR2_X1 U9707 ( .A(n8176), .B(n8175), .ZN(n8177) );
  XNOR2_X1 U9708 ( .A(n8178), .B(n8177), .ZN(n8186) );
  NOR2_X1 U9709 ( .A1(n9139), .A2(n8179), .ZN(n8180) );
  AOI211_X1 U9710 ( .C1(n9142), .C2(n9155), .A(n8181), .B(n8180), .ZN(n8182)
         );
  OAI21_X1 U9711 ( .B1(n9958), .B2(n9145), .A(n8182), .ZN(n8183) );
  AOI21_X1 U9712 ( .B1(n8184), .B2(n9137), .A(n8183), .ZN(n8185) );
  OAI21_X1 U9713 ( .B1(n8186), .B2(n9132), .A(n8185), .ZN(P1_U3228) );
  INV_X1 U9714 ( .A(n8557), .ZN(n8190) );
  OAI22_X1 U9715 ( .A1(n8189), .A2(n8188), .B1(P2_REG2_REG_15__SCAN_IN), .B2(
        n8187), .ZN(n8553) );
  XOR2_X1 U9716 ( .A(n8557), .B(P2_REG2_REG_16__SCAN_IN), .Z(n8554) );
  NOR2_X1 U9717 ( .A1(n8553), .A2(n8554), .ZN(n8552) );
  XNOR2_X1 U9718 ( .A(n8204), .B(P2_REG2_REG_17__SCAN_IN), .ZN(n8565) );
  INV_X1 U9719 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8579) );
  NAND2_X1 U9720 ( .A1(n8580), .A2(n8579), .ZN(n8578) );
  NAND2_X1 U9721 ( .A1(n8191), .A2(n4516), .ZN(n8192) );
  NAND2_X1 U9722 ( .A1(n8578), .A2(n8192), .ZN(n8193) );
  XNOR2_X1 U9723 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n8193), .ZN(n8213) );
  NAND2_X1 U9724 ( .A1(n8194), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n8198) );
  OR2_X1 U9725 ( .A1(n8196), .A2(n8195), .ZN(n8197) );
  NAND2_X1 U9726 ( .A1(n8198), .A2(n8197), .ZN(n8550) );
  INV_X1 U9727 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n8199) );
  XNOR2_X1 U9728 ( .A(n8557), .B(n8199), .ZN(n8551) );
  NAND2_X1 U9729 ( .A1(n8557), .A2(n8199), .ZN(n8569) );
  INV_X1 U9730 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n8200) );
  XNOR2_X1 U9731 ( .A(n8204), .B(n8200), .ZN(n8568) );
  AND2_X1 U9732 ( .A1(n8569), .A2(n8568), .ZN(n8201) );
  NAND2_X1 U9733 ( .A1(n8570), .A2(n8201), .ZN(n8567) );
  OR2_X1 U9734 ( .A1(n8202), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8206) );
  NAND2_X1 U9735 ( .A1(n8202), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8203) );
  NAND2_X1 U9736 ( .A1(n8206), .A2(n8203), .ZN(n8581) );
  AND2_X1 U9737 ( .A1(n8204), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8582) );
  NOR2_X1 U9738 ( .A1(n8581), .A2(n8582), .ZN(n8205) );
  NAND2_X1 U9739 ( .A1(n8567), .A2(n8205), .ZN(n8585) );
  NAND2_X1 U9740 ( .A1(n8585), .A2(n8206), .ZN(n8208) );
  XNOR2_X1 U9741 ( .A(n8208), .B(n8207), .ZN(n8211) );
  AOI21_X1 U9742 ( .B1(n8211), .B2(n8542), .A(n8540), .ZN(n8209) );
  OAI21_X1 U9743 ( .B1(n8213), .B2(n8564), .A(n8209), .ZN(n8210) );
  INV_X1 U9744 ( .A(n8210), .ZN(n8215) );
  INV_X1 U9745 ( .A(n8211), .ZN(n8212) );
  AOI22_X1 U9746 ( .A1(n8213), .A2(n8593), .B1(n8212), .B2(n8542), .ZN(n8214)
         );
  NAND2_X1 U9747 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n8339) );
  OAI211_X1 U9748 ( .C1(n4796), .C2(n8217), .A(n8216), .B(n8339), .ZN(P2_U3264) );
  INV_X1 U9749 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n8220) );
  INV_X1 U9750 ( .A(n8218), .ZN(n8991) );
  OAI222_X1 U9751 ( .A1(n9787), .A2(n8220), .B1(n9798), .B2(n8991), .C1(n8219), 
        .C2(P1_U3084), .ZN(P1_U3323) );
  AND2_X1 U9752 ( .A1(n8223), .A2(P2_B_REG_SCAN_IN), .ZN(n8224) );
  NOR2_X1 U9753 ( .A1(n8823), .A2(n8224), .ZN(n8261) );
  NOR2_X1 U9754 ( .A1(n8924), .A2(n8794), .ZN(n8229) );
  AOI21_X1 U9755 ( .B1(n8231), .B2(n8230), .A(n8229), .ZN(n8232) );
  NAND2_X1 U9756 ( .A1(n8919), .A2(n8515), .ZN(n8234) );
  NAND2_X1 U9757 ( .A1(n8806), .A2(n8234), .ZN(n8780) );
  INV_X1 U9758 ( .A(n8780), .ZN(n8236) );
  INV_X1 U9759 ( .A(n8477), .ZN(n8795) );
  OR2_X1 U9760 ( .A1(n8915), .A2(n8795), .ZN(n8237) );
  NAND2_X1 U9761 ( .A1(n8909), .A2(n8514), .ZN(n8239) );
  NOR2_X1 U9762 ( .A1(n8909), .A2(n8514), .ZN(n8238) );
  INV_X1 U9763 ( .A(n8744), .ZN(n8714) );
  INV_X1 U9764 ( .A(n8678), .ZN(n8512) );
  NAND2_X1 U9765 ( .A1(n8662), .A2(n8241), .ZN(n8643) );
  INV_X1 U9766 ( .A(n8873), .ZN(n8653) );
  XNOR2_X1 U9767 ( .A(n8245), .B(n8244), .ZN(n8855) );
  INV_X1 U9768 ( .A(n8855), .ZN(n8257) );
  INV_X1 U9769 ( .A(n8852), .ZN(n8255) );
  INV_X1 U9770 ( .A(n8915), .ZN(n8785) );
  AOI21_X1 U9771 ( .B1(n8852), .B2(n8601), .A(n10149), .ZN(n8248) );
  INV_X1 U9772 ( .A(n8248), .ZN(n8251) );
  INV_X1 U9773 ( .A(n8596), .ZN(n8250) );
  NOR2_X1 U9774 ( .A1(n8251), .A2(n8250), .ZN(n8851) );
  NAND2_X1 U9775 ( .A1(n8851), .A2(n8838), .ZN(n8254) );
  AOI22_X1 U9776 ( .A1(n8252), .A2(n8800), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n8717), .ZN(n8253) );
  OAI211_X1 U9777 ( .C1(n8255), .C2(n8803), .A(n8254), .B(n8253), .ZN(n8256)
         );
  AOI21_X1 U9778 ( .B1(n8257), .B2(n10099), .A(n8256), .ZN(n8258) );
  OAI21_X1 U9779 ( .B1(n8854), .B2(n8717), .A(n8258), .ZN(P2_U3267) );
  NAND2_X1 U9780 ( .A1(n8510), .A2(n8261), .ZN(n8849) );
  NOR2_X1 U9781 ( .A1(n8836), .A2(n8849), .ZN(n8597) );
  NOR2_X1 U9782 ( .A1(n10093), .A2(n8262), .ZN(n8263) );
  AOI211_X1 U9783 ( .C1(n8844), .C2(n10095), .A(n8597), .B(n8263), .ZN(n8264)
         );
  OAI21_X1 U9784 ( .B1(n8846), .B2(n10074), .A(n8264), .ZN(P2_U3265) );
  XNOR2_X1 U9785 ( .A(n8861), .B(n8306), .ZN(n8348) );
  NOR2_X1 U9786 ( .A1(n8608), .A2(n8354), .ZN(n8349) );
  XNOR2_X1 U9787 ( .A(n8348), .B(n8349), .ZN(n8352) );
  INV_X1 U9788 ( .A(n8265), .ZN(n8266) );
  NAND2_X1 U9789 ( .A1(n8267), .A2(n8266), .ZN(n8268) );
  XNOR2_X1 U9790 ( .A(n8919), .B(n8356), .ZN(n8402) );
  NOR2_X1 U9791 ( .A1(n8501), .A2(n8354), .ZN(n8273) );
  NOR2_X1 U9792 ( .A1(n8270), .A2(n8354), .ZN(n8398) );
  XNOR2_X1 U9793 ( .A(n8924), .B(n8356), .ZN(n8397) );
  OAI22_X1 U9794 ( .A1(n8402), .A2(n8273), .B1(n8398), .B2(n8397), .ZN(n8271)
         );
  INV_X1 U9795 ( .A(n8397), .ZN(n8400) );
  INV_X1 U9796 ( .A(n8398), .ZN(n8272) );
  INV_X1 U9797 ( .A(n8273), .ZN(n8401) );
  OAI21_X1 U9798 ( .B1(n8400), .B2(n8272), .A(n8401), .ZN(n8275) );
  AND3_X1 U9799 ( .A1(n8397), .A2(n8398), .A3(n8273), .ZN(n8274) );
  AOI21_X1 U9800 ( .B1(n8402), .B2(n8275), .A(n8274), .ZN(n8276) );
  XNOR2_X1 U9801 ( .A(n8915), .B(n8356), .ZN(n8277) );
  NOR2_X1 U9802 ( .A1(n8477), .A2(n8354), .ZN(n8278) );
  NAND2_X1 U9803 ( .A1(n8277), .A2(n8278), .ZN(n8281) );
  INV_X1 U9804 ( .A(n8277), .ZN(n8478) );
  INV_X1 U9805 ( .A(n8278), .ZN(n8279) );
  NAND2_X1 U9806 ( .A1(n8478), .A2(n8279), .ZN(n8280) );
  AND2_X1 U9807 ( .A1(n8281), .A2(n8280), .ZN(n8411) );
  XNOR2_X1 U9808 ( .A(n8909), .B(n8356), .ZN(n8282) );
  AND2_X1 U9809 ( .A1(n8514), .A2(n8310), .ZN(n8283) );
  NAND2_X1 U9810 ( .A1(n8282), .A2(n8283), .ZN(n8287) );
  INV_X1 U9811 ( .A(n8282), .ZN(n8342) );
  INV_X1 U9812 ( .A(n8283), .ZN(n8284) );
  NAND2_X1 U9813 ( .A1(n8342), .A2(n8284), .ZN(n8285) );
  AND2_X1 U9814 ( .A1(n8287), .A2(n8285), .ZN(n8474) );
  NAND2_X1 U9815 ( .A1(n8286), .A2(n8474), .ZN(n8336) );
  XNOR2_X1 U9816 ( .A(n8755), .B(n8356), .ZN(n8288) );
  NAND2_X1 U9817 ( .A1(n8760), .A2(n8310), .ZN(n8289) );
  XNOR2_X1 U9818 ( .A(n8288), .B(n8289), .ZN(n8343) );
  NAND3_X1 U9819 ( .A1(n8336), .A2(n8343), .A3(n8287), .ZN(n8337) );
  INV_X1 U9820 ( .A(n8288), .ZN(n8290) );
  NAND2_X1 U9821 ( .A1(n8290), .A2(n8289), .ZN(n8291) );
  XNOR2_X1 U9822 ( .A(n8898), .B(n8356), .ZN(n8292) );
  NOR2_X1 U9823 ( .A1(n8744), .A2(n8354), .ZN(n8293) );
  NAND2_X1 U9824 ( .A1(n8292), .A2(n8293), .ZN(n8296) );
  INV_X1 U9825 ( .A(n8292), .ZN(n8375) );
  INV_X1 U9826 ( .A(n8293), .ZN(n8294) );
  NAND2_X1 U9827 ( .A1(n8375), .A2(n8294), .ZN(n8295) );
  NAND2_X1 U9828 ( .A1(n8296), .A2(n8295), .ZN(n8443) );
  XNOR2_X1 U9829 ( .A(n8893), .B(n8356), .ZN(n8299) );
  NAND2_X1 U9830 ( .A1(n8513), .A2(n8310), .ZN(n8297) );
  XNOR2_X1 U9831 ( .A(n8299), .B(n8297), .ZN(n8373) );
  XNOR2_X1 U9832 ( .A(n8692), .B(n8306), .ZN(n8301) );
  AND2_X1 U9833 ( .A1(n8715), .A2(n8310), .ZN(n8302) );
  INV_X1 U9834 ( .A(n8297), .ZN(n8298) );
  AND2_X1 U9835 ( .A1(n8299), .A2(n8298), .ZN(n8464) );
  AOI21_X1 U9836 ( .B1(n8301), .B2(n8302), .A(n8464), .ZN(n8300) );
  INV_X1 U9837 ( .A(n8301), .ZN(n8466) );
  INV_X1 U9838 ( .A(n8302), .ZN(n8470) );
  NAND2_X1 U9839 ( .A1(n8466), .A2(n8470), .ZN(n8303) );
  NAND2_X1 U9840 ( .A1(n8304), .A2(n8303), .ZN(n8309) );
  INV_X1 U9841 ( .A(n8309), .ZN(n8305) );
  XNOR2_X1 U9842 ( .A(n8883), .B(n8356), .ZN(n8308) );
  XNOR2_X1 U9843 ( .A(n8667), .B(n8306), .ZN(n8418) );
  OR2_X1 U9844 ( .A1(n8678), .A2(n8354), .ZN(n8421) );
  NAND2_X1 U9845 ( .A1(n8418), .A2(n8421), .ZN(n8307) );
  NAND2_X1 U9846 ( .A1(n8416), .A2(n8307), .ZN(n8314) );
  NAND2_X1 U9847 ( .A1(n8658), .A2(n8310), .ZN(n8327) );
  AOI21_X1 U9848 ( .B1(n8418), .B2(n8678), .A(n8327), .ZN(n8311) );
  XNOR2_X1 U9849 ( .A(n8873), .B(n8356), .ZN(n8388) );
  NOR2_X1 U9850 ( .A1(n8661), .A2(n8354), .ZN(n8315) );
  AND2_X1 U9851 ( .A1(n8388), .A2(n8315), .ZN(n8387) );
  INV_X1 U9852 ( .A(n8388), .ZN(n8317) );
  INV_X1 U9853 ( .A(n8315), .ZN(n8316) );
  NAND2_X1 U9854 ( .A1(n8317), .A2(n8316), .ZN(n8390) );
  XNOR2_X1 U9855 ( .A(n8867), .B(n8356), .ZN(n8319) );
  NOR2_X1 U9856 ( .A1(n8321), .A2(n8354), .ZN(n8318) );
  XNOR2_X1 U9857 ( .A(n8319), .B(n8318), .ZN(n8487) );
  XOR2_X1 U9858 ( .A(n8352), .B(n8353), .Z(n8320) );
  NAND2_X1 U9859 ( .A1(n8320), .A2(n10043), .ZN(n8326) );
  NOR2_X1 U9860 ( .A1(n8321), .A2(n10038), .ZN(n8324) );
  OAI22_X1 U9861 ( .A1(n8355), .A2(n10007), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8322), .ZN(n8323) );
  AOI211_X1 U9862 ( .C1(n8505), .C2(n8621), .A(n8324), .B(n8323), .ZN(n8325)
         );
  OAI211_X1 U9863 ( .C1(n8624), .C2(n8486), .A(n8326), .B(n8325), .ZN(P2_U3216) );
  INV_X1 U9864 ( .A(n8329), .ZN(n8328) );
  NOR2_X1 U9865 ( .A1(n8328), .A2(n8327), .ZN(n8417) );
  AOI22_X1 U9866 ( .A1(n8329), .A2(n10043), .B1(n10042), .B2(n8658), .ZN(n8335) );
  INV_X1 U9867 ( .A(n8330), .ZN(n8682) );
  NOR2_X1 U9868 ( .A1(n10038), .A2(n8677), .ZN(n8332) );
  OAI22_X1 U9869 ( .A1(n8678), .A2(n10007), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9666), .ZN(n8331) );
  AOI211_X1 U9870 ( .C1(n8505), .C2(n8682), .A(n8332), .B(n8331), .ZN(n8334)
         );
  NAND2_X1 U9871 ( .A1(n8883), .A2(n10052), .ZN(n8333) );
  OAI211_X1 U9872 ( .C1(n8417), .C2(n8335), .A(n8334), .B(n8333), .ZN(P2_U3218) );
  OAI21_X1 U9873 ( .B1(n8336), .B2(n8343), .A(n8337), .ZN(n8338) );
  NAND2_X1 U9874 ( .A1(n8338), .A2(n10043), .ZN(n8347) );
  NOR2_X1 U9875 ( .A1(n10055), .A2(n8749), .ZN(n8341) );
  OAI21_X1 U9876 ( .B1(n10007), .B2(n8744), .A(n8339), .ZN(n8340) );
  AOI211_X1 U9877 ( .C1(n8755), .C2(n10052), .A(n8341), .B(n8340), .ZN(n8346)
         );
  NOR3_X1 U9878 ( .A1(n8343), .A2(n8342), .A3(n10026), .ZN(n8344) );
  OAI21_X1 U9879 ( .B1(n8344), .B2(n10029), .A(n8514), .ZN(n8345) );
  NAND3_X1 U9880 ( .A1(n8347), .A2(n8346), .A3(n8345), .ZN(P2_U3221) );
  INV_X1 U9881 ( .A(n8348), .ZN(n8350) );
  AND2_X1 U9882 ( .A1(n8350), .A2(n8349), .ZN(n8351) );
  NOR2_X1 U9883 ( .A1(n8355), .A2(n8354), .ZN(n8357) );
  XNOR2_X1 U9884 ( .A(n8357), .B(n8356), .ZN(n8360) );
  NOR3_X1 U9885 ( .A1(n4823), .A2(n8958), .A3(n8360), .ZN(n8358) );
  AOI21_X1 U9886 ( .B1(n8360), .B2(n4823), .A(n8358), .ZN(n8366) );
  NAND3_X1 U9887 ( .A1(n8856), .A2(n8360), .A3(n10159), .ZN(n8359) );
  OAI21_X1 U9888 ( .B1(n8856), .B2(n8360), .A(n8359), .ZN(n8361) );
  NAND2_X1 U9889 ( .A1(n8367), .A2(n8361), .ZN(n8365) );
  OAI22_X1 U9890 ( .A1(n4823), .A2(n8486), .B1(n8363), .B2(n8362), .ZN(n8364)
         );
  OAI211_X1 U9891 ( .C1(n8367), .C2(n8366), .A(n8365), .B(n8364), .ZN(n8372)
         );
  INV_X1 U9892 ( .A(n8368), .ZN(n8602) );
  OAI22_X1 U9893 ( .A1(n8607), .A2(n10007), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8369), .ZN(n8370) );
  AOI21_X1 U9894 ( .B1(n8602), .B2(n8505), .A(n8370), .ZN(n8371) );
  OAI211_X1 U9895 ( .C1(n8608), .C2(n10038), .A(n8372), .B(n8371), .ZN(
        P2_U3222) );
  INV_X1 U9896 ( .A(n8373), .ZN(n8374) );
  AOI21_X1 U9897 ( .B1(n8445), .B2(n8374), .A(n10010), .ZN(n8378) );
  NOR3_X1 U9898 ( .A1(n8375), .A2(n8744), .A3(n10026), .ZN(n8377) );
  OAI21_X1 U9899 ( .B1(n8378), .B2(n8377), .A(n8376), .ZN(n8383) );
  NOR2_X1 U9900 ( .A1(n10038), .A2(n8744), .ZN(n8381) );
  OAI22_X1 U9901 ( .A1(n10007), .A2(n8677), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8379), .ZN(n8380) );
  AOI211_X1 U9902 ( .C1(n8505), .C2(n8705), .A(n8381), .B(n8380), .ZN(n8382)
         );
  OAI211_X1 U9903 ( .C1(n8707), .C2(n8486), .A(n8383), .B(n8382), .ZN(P2_U3225) );
  NOR2_X1 U9904 ( .A1(n8678), .A2(n8821), .ZN(n8384) );
  AOI21_X1 U9905 ( .B1(n8615), .B2(n10060), .A(n8384), .ZN(n8647) );
  AOI22_X1 U9906 ( .A1(n8505), .A2(n8650), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3152), .ZN(n8385) );
  OAI21_X1 U9907 ( .B1(n8647), .B2(n8386), .A(n8385), .ZN(n8395) );
  NOR3_X1 U9908 ( .A1(n8387), .A2(n4720), .A3(n10010), .ZN(n8393) );
  NAND3_X1 U9909 ( .A1(n8388), .A2(n10042), .A3(n4846), .ZN(n8389) );
  OAI21_X1 U9910 ( .B1(n8390), .B2(n10010), .A(n8389), .ZN(n8392) );
  MUX2_X1 U9911 ( .A(n8393), .B(n8392), .S(n8391), .Z(n8394) );
  AOI211_X1 U9912 ( .C1(n10052), .C2(n8873), .A(n8395), .B(n8394), .ZN(n8396)
         );
  INV_X1 U9913 ( .A(n8396), .ZN(P2_U3227) );
  XNOR2_X1 U9914 ( .A(n4363), .B(n8397), .ZN(n8497) );
  NAND2_X1 U9915 ( .A1(n8497), .A2(n8398), .ZN(n8498) );
  OAI21_X1 U9916 ( .B1(n8400), .B2(n4363), .A(n8498), .ZN(n8404) );
  XNOR2_X1 U9917 ( .A(n8402), .B(n8401), .ZN(n8403) );
  XNOR2_X1 U9918 ( .A(n8404), .B(n8403), .ZN(n8409) );
  OAI22_X1 U9919 ( .A1(n10007), .A2(n8477), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8556), .ZN(n8405) );
  AOI21_X1 U9920 ( .B1(n10029), .B2(n8794), .A(n8405), .ZN(n8406) );
  OAI21_X1 U9921 ( .B1(n8799), .B2(n10055), .A(n8406), .ZN(n8407) );
  AOI21_X1 U9922 ( .B1(n8919), .B2(n10052), .A(n8407), .ZN(n8408) );
  OAI21_X1 U9923 ( .B1(n8409), .B2(n10010), .A(n8408), .ZN(P2_U3228) );
  OAI211_X1 U9924 ( .C1(n8411), .C2(n8410), .A(n8476), .B(n10043), .ZN(n8415)
         );
  OAI22_X1 U9925 ( .A1(n8743), .A2(n8823), .B1(n8501), .B2(n8821), .ZN(n8776)
         );
  AOI22_X1 U9926 ( .A1(n8493), .A2(n8776), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n8412) );
  OAI21_X1 U9927 ( .B1(n8783), .B2(n10055), .A(n8412), .ZN(n8413) );
  AOI21_X1 U9928 ( .B1(n8915), .B2(n10052), .A(n8413), .ZN(n8414) );
  NAND2_X1 U9929 ( .A1(n8415), .A2(n8414), .ZN(P2_U3230) );
  NOR2_X1 U9930 ( .A1(n8417), .A2(n8416), .ZN(n8419) );
  XNOR2_X1 U9931 ( .A(n8419), .B(n8418), .ZN(n8422) );
  OAI22_X1 U9932 ( .A1(n8422), .A2(n10010), .B1(n8678), .B2(n10026), .ZN(n8420) );
  OAI21_X1 U9933 ( .B1(n8422), .B2(n8421), .A(n8420), .ZN(n8428) );
  NOR2_X1 U9934 ( .A1(n8423), .A2(n10038), .ZN(n8426) );
  OAI22_X1 U9935 ( .A1(n8661), .A2(n10007), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8424), .ZN(n8425) );
  AOI211_X1 U9936 ( .C1(n8505), .C2(n8666), .A(n8426), .B(n8425), .ZN(n8427)
         );
  OAI211_X1 U9937 ( .C1(n8877), .C2(n8486), .A(n8428), .B(n8427), .ZN(P2_U3231) );
  NOR2_X1 U9938 ( .A1(n10055), .A2(n8429), .ZN(n8433) );
  OAI21_X1 U9939 ( .B1(n10007), .B2(n8431), .A(n8430), .ZN(n8432) );
  AOI211_X1 U9940 ( .C1(n10052), .C2(n8434), .A(n8433), .B(n8432), .ZN(n8442)
         );
  OAI21_X1 U9941 ( .B1(n8437), .B2(n10027), .A(n8435), .ZN(n8436) );
  NAND2_X1 U9942 ( .A1(n8436), .A2(n10043), .ZN(n8441) );
  NOR3_X1 U9943 ( .A1(n10026), .A2(n8438), .A3(n8437), .ZN(n8439) );
  OAI21_X1 U9944 ( .B1(n8439), .B2(n10029), .A(n8522), .ZN(n8440) );
  NAND3_X1 U9945 ( .A1(n8442), .A2(n8441), .A3(n8440), .ZN(P2_U3232) );
  INV_X1 U9946 ( .A(n8898), .ZN(n8725) );
  AOI21_X1 U9947 ( .B1(n8444), .B2(n8443), .A(n10010), .ZN(n8446) );
  NAND2_X1 U9948 ( .A1(n8446), .A2(n8445), .ZN(n8451) );
  NOR2_X1 U9949 ( .A1(n10038), .A2(n8729), .ZN(n8449) );
  OAI22_X1 U9950 ( .A1(n10007), .A2(n8730), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8447), .ZN(n8448) );
  AOI211_X1 U9951 ( .C1(n8505), .C2(n8723), .A(n8449), .B(n8448), .ZN(n8450)
         );
  OAI211_X1 U9952 ( .C1(n8725), .C2(n8486), .A(n8451), .B(n8450), .ZN(P2_U3235) );
  OAI21_X1 U9953 ( .B1(n10007), .B2(n8499), .A(n8452), .ZN(n8453) );
  AOI21_X1 U9954 ( .B1(n10029), .B2(n10035), .A(n8453), .ZN(n8454) );
  OAI21_X1 U9955 ( .B1(n8455), .B2(n10055), .A(n8454), .ZN(n8460) );
  AOI211_X1 U9956 ( .C1(n8458), .C2(n8457), .A(n10010), .B(n8456), .ZN(n8459)
         );
  AOI211_X1 U9957 ( .C1(n10052), .C2(n8934), .A(n8460), .B(n8459), .ZN(n8461)
         );
  INV_X1 U9958 ( .A(n8461), .ZN(P2_U3236) );
  AOI22_X1 U9959 ( .A1(n8658), .A2(n10060), .B1(n10058), .B2(n8513), .ZN(n8696) );
  INV_X1 U9960 ( .A(n8696), .ZN(n8462) );
  AOI22_X1 U9961 ( .A1(n8462), .A2(n8493), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3152), .ZN(n8463) );
  OAI21_X1 U9962 ( .B1(n8689), .B2(n10055), .A(n8463), .ZN(n8469) );
  INV_X1 U9963 ( .A(n8464), .ZN(n8465) );
  NAND2_X1 U9964 ( .A1(n8376), .A2(n8465), .ZN(n8467) );
  XNOR2_X1 U9965 ( .A(n8467), .B(n8466), .ZN(n8471) );
  NOR3_X1 U9966 ( .A1(n8471), .A2(n8677), .A3(n10026), .ZN(n8468) );
  AOI211_X1 U9967 ( .C1(n10052), .C2(n8888), .A(n8469), .B(n8468), .ZN(n8473)
         );
  NAND3_X1 U9968 ( .A1(n8471), .A2(n10043), .A3(n8470), .ZN(n8472) );
  NAND2_X1 U9969 ( .A1(n8473), .A2(n8472), .ZN(P2_U3237) );
  INV_X1 U9970 ( .A(n8909), .ZN(n8766) );
  INV_X1 U9971 ( .A(n8474), .ZN(n8475) );
  AOI21_X1 U9972 ( .B1(n8476), .B2(n8475), .A(n10010), .ZN(n8480) );
  NOR3_X1 U9973 ( .A1(n8478), .A2(n8477), .A3(n10026), .ZN(n8479) );
  OAI21_X1 U9974 ( .B1(n8480), .B2(n8479), .A(n8336), .ZN(n8485) );
  INV_X1 U9975 ( .A(n8481), .ZN(n8764) );
  NAND2_X1 U9976 ( .A1(n10029), .A2(n8795), .ZN(n8482) );
  NAND2_X1 U9977 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n8589) );
  OAI211_X1 U9978 ( .C1(n8729), .C2(n10007), .A(n8482), .B(n8589), .ZN(n8483)
         );
  AOI21_X1 U9979 ( .B1(n8764), .B2(n8505), .A(n8483), .ZN(n8484) );
  OAI211_X1 U9980 ( .C1(n8766), .C2(n8486), .A(n8485), .B(n8484), .ZN(P2_U3240) );
  XNOR2_X1 U9981 ( .A(n8488), .B(n8487), .ZN(n8496) );
  OR2_X1 U9982 ( .A1(n8608), .A2(n8823), .ZN(n8490) );
  OR2_X1 U9983 ( .A1(n8661), .A2(n8821), .ZN(n8489) );
  NAND2_X1 U9984 ( .A1(n8490), .A2(n8489), .ZN(n8634) );
  OAI22_X1 U9985 ( .A1(n8639), .A2(n10055), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8491), .ZN(n8492) );
  AOI21_X1 U9986 ( .B1(n8634), .B2(n8493), .A(n8492), .ZN(n8495) );
  NAND2_X1 U9987 ( .A1(n8867), .A2(n10052), .ZN(n8494) );
  OAI211_X1 U9988 ( .C1(n8496), .C2(n10010), .A(n8495), .B(n8494), .ZN(
        P2_U3242) );
  AOI22_X1 U9989 ( .A1(n8497), .A2(n10043), .B1(n10042), .B2(n8794), .ZN(n8509) );
  INV_X1 U9990 ( .A(n8498), .ZN(n8508) );
  NOR2_X1 U9991 ( .A1(n10038), .A2(n8499), .ZN(n8503) );
  OAI22_X1 U9992 ( .A1(n10007), .A2(n8501), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8500), .ZN(n8502) );
  AOI211_X1 U9993 ( .C1(n8505), .C2(n8504), .A(n8503), .B(n8502), .ZN(n8507)
         );
  NAND2_X1 U9994 ( .A1(n8924), .A2(n10052), .ZN(n8506) );
  OAI211_X1 U9995 ( .C1(n8509), .C2(n8508), .A(n8507), .B(n8506), .ZN(P2_U3243) );
  MUX2_X1 U9996 ( .A(n8510), .B(P2_DATAO_REG_31__SCAN_IN), .S(n8518), .Z(
        P2_U3583) );
  MUX2_X1 U9997 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8511), .S(P2_U3966), .Z(
        P2_U3582) );
  MUX2_X1 U9998 ( .A(n8616), .B(P2_DATAO_REG_28__SCAN_IN), .S(n8518), .Z(
        P2_U3580) );
  MUX2_X1 U9999 ( .A(n8615), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8518), .Z(
        P2_U3578) );
  MUX2_X1 U10000 ( .A(n4846), .B(P2_DATAO_REG_25__SCAN_IN), .S(n8518), .Z(
        P2_U3577) );
  MUX2_X1 U10001 ( .A(n8512), .B(P2_DATAO_REG_24__SCAN_IN), .S(n8518), .Z(
        P2_U3576) );
  MUX2_X1 U10002 ( .A(n8658), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8518), .Z(
        P2_U3575) );
  MUX2_X1 U10003 ( .A(n8715), .B(P2_DATAO_REG_22__SCAN_IN), .S(n8518), .Z(
        P2_U3574) );
  MUX2_X1 U10004 ( .A(n8513), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8518), .Z(
        P2_U3573) );
  MUX2_X1 U10005 ( .A(n8714), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8518), .Z(
        P2_U3572) );
  MUX2_X1 U10006 ( .A(n8760), .B(P2_DATAO_REG_19__SCAN_IN), .S(n8518), .Z(
        P2_U3571) );
  MUX2_X1 U10007 ( .A(n8514), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8518), .Z(
        P2_U3570) );
  MUX2_X1 U10008 ( .A(n8795), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8518), .Z(
        P2_U3569) );
  MUX2_X1 U10009 ( .A(n8515), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8518), .Z(
        P2_U3568) );
  MUX2_X1 U10010 ( .A(n8794), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8518), .Z(
        P2_U3567) );
  MUX2_X1 U10011 ( .A(n8516), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8518), .Z(
        P2_U3566) );
  MUX2_X1 U10012 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8517), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10013 ( .A(n10035), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8518), .Z(
        P2_U3564) );
  MUX2_X1 U10014 ( .A(n8519), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8518), .Z(
        P2_U3563) );
  MUX2_X1 U10015 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n10004), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10016 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n10061), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U10017 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n8520), .S(P2_U3966), .Z(
        P2_U3559) );
  MUX2_X1 U10018 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n10059), .S(P2_U3966), .Z(
        P2_U3558) );
  MUX2_X1 U10019 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n8521), .S(P2_U3966), .Z(
        P2_U3557) );
  MUX2_X1 U10020 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n10019), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U10021 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n8522), .S(P2_U3966), .Z(
        P2_U3555) );
  MUX2_X1 U10022 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n6673), .S(P2_U3966), .Z(
        P2_U3554) );
  MUX2_X1 U10023 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n8523), .S(P2_U3966), .Z(
        P2_U3553) );
  OAI211_X1 U10024 ( .C1(n8526), .C2(n8525), .A(n8593), .B(n8524), .ZN(n8535)
         );
  AOI22_X1 U10025 ( .A1(n8587), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n8534) );
  NAND2_X1 U10026 ( .A1(n8540), .A2(n8527), .ZN(n8533) );
  INV_X1 U10027 ( .A(n9003), .ZN(n8529) );
  MUX2_X1 U10028 ( .A(n6865), .B(P2_REG1_REG_1__SCAN_IN), .S(n8527), .Z(n8528)
         );
  OAI21_X1 U10029 ( .B1(n6136), .B2(n8529), .A(n8528), .ZN(n8530) );
  NAND3_X1 U10030 ( .A1(n8542), .A2(n8531), .A3(n8530), .ZN(n8532) );
  NAND4_X1 U10031 ( .A1(n8535), .A2(n8534), .A3(n8533), .A4(n8532), .ZN(
        P2_U3246) );
  OAI211_X1 U10032 ( .C1(n8538), .C2(n8537), .A(n8593), .B(n8536), .ZN(n8548)
         );
  AOI22_X1 U10033 ( .A1(n8587), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n8547) );
  NAND2_X1 U10034 ( .A1(n8540), .A2(n8539), .ZN(n8546) );
  OAI211_X1 U10035 ( .C1(n8544), .C2(n8543), .A(n8542), .B(n8541), .ZN(n8545)
         );
  NAND4_X1 U10036 ( .A1(n8548), .A2(n8547), .A3(n8546), .A4(n8545), .ZN(
        P2_U3247) );
  INV_X1 U10037 ( .A(n8570), .ZN(n8549) );
  AOI21_X1 U10038 ( .B1(n8551), .B2(n8550), .A(n8549), .ZN(n8562) );
  AOI211_X1 U10039 ( .C1(n8554), .C2(n8553), .A(n8564), .B(n8552), .ZN(n8555)
         );
  INV_X1 U10040 ( .A(n8555), .ZN(n8561) );
  NOR2_X1 U10041 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8556), .ZN(n8559) );
  NOR2_X1 U10042 ( .A1(n8590), .A2(n8557), .ZN(n8558) );
  AOI211_X1 U10043 ( .C1(n8587), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n8559), .B(
        n8558), .ZN(n8560) );
  OAI211_X1 U10044 ( .C1(n8562), .C2(n8584), .A(n8561), .B(n8560), .ZN(
        P2_U3261) );
  AOI211_X1 U10045 ( .C1(n8566), .C2(n8565), .A(n8564), .B(n8563), .ZN(n8577)
         );
  INV_X1 U10046 ( .A(n8567), .ZN(n8583) );
  AOI21_X1 U10047 ( .B1(n8570), .B2(n8569), .A(n8568), .ZN(n8571) );
  NOR3_X1 U10048 ( .A1(n8583), .A2(n8571), .A3(n8584), .ZN(n8576) );
  AND2_X1 U10049 ( .A1(P2_U3152), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n8572) );
  AOI21_X1 U10050 ( .B1(n8587), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n8572), .ZN(
        n8573) );
  OAI21_X1 U10051 ( .B1(n8590), .B2(n8574), .A(n8573), .ZN(n8575) );
  OR3_X1 U10052 ( .A1(n8577), .A2(n8576), .A3(n8575), .ZN(P2_U3262) );
  OAI21_X1 U10053 ( .B1(n8580), .B2(n8579), .A(n8578), .ZN(n8594) );
  OAI21_X1 U10054 ( .B1(n8583), .B2(n8582), .A(n8581), .ZN(n8586) );
  AOI21_X1 U10055 ( .B1(n8586), .B2(n8585), .A(n8584), .ZN(n8592) );
  NAND2_X1 U10056 ( .A1(n8587), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n8588) );
  OAI211_X1 U10057 ( .C1(n8590), .C2(n4516), .A(n8589), .B(n8588), .ZN(n8591)
         );
  AOI211_X1 U10058 ( .C1(n8594), .C2(n8593), .A(n8592), .B(n8591), .ZN(n8595)
         );
  INV_X1 U10059 ( .A(n8595), .ZN(P2_U3263) );
  XNOR2_X1 U10060 ( .A(n8596), .B(n8847), .ZN(n8850) );
  AOI21_X1 U10061 ( .B1(n8836), .B2(P2_REG2_REG_30__SCAN_IN), .A(n8597), .ZN(
        n8599) );
  NAND2_X1 U10062 ( .A1(n8847), .A2(n10095), .ZN(n8598) );
  OAI211_X1 U10063 ( .C1(n8850), .C2(n10074), .A(n8599), .B(n8598), .ZN(
        P2_U3266) );
  XNOR2_X1 U10064 ( .A(n8600), .B(n8605), .ZN(n8860) );
  AOI21_X1 U10065 ( .B1(n8856), .B2(n8619), .A(n8249), .ZN(n8857) );
  AOI22_X1 U10066 ( .A1(n8602), .A2(n8800), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n8717), .ZN(n8603) );
  OAI21_X1 U10067 ( .B1(n4823), .B2(n8803), .A(n8603), .ZN(n8613) );
  INV_X1 U10068 ( .A(n8604), .ZN(n8606) );
  AOI21_X1 U10069 ( .B1(n8606), .B2(n8605), .A(n8820), .ZN(n8611) );
  OAI22_X1 U10070 ( .A1(n8608), .A2(n8821), .B1(n8607), .B2(n8823), .ZN(n8609)
         );
  AOI21_X1 U10071 ( .B1(n8611), .B2(n8610), .A(n8609), .ZN(n8859) );
  NOR2_X1 U10072 ( .A1(n8859), .A2(n8717), .ZN(n8612) );
  AOI211_X1 U10073 ( .C1(n8813), .C2(n8857), .A(n8613), .B(n8612), .ZN(n8614)
         );
  OAI21_X1 U10074 ( .B1(n8860), .B2(n8790), .A(n8614), .ZN(P2_U3268) );
  XOR2_X1 U10075 ( .A(n8618), .B(n8617), .Z(n8865) );
  INV_X1 U10076 ( .A(n8865), .ZN(n8626) );
  OR2_X1 U10077 ( .A1(n8624), .A2(n8636), .ZN(n8620) );
  AND2_X1 U10078 ( .A1(n8620), .A2(n8619), .ZN(n8862) );
  NAND2_X1 U10079 ( .A1(n8862), .A2(n8813), .ZN(n8623) );
  AOI22_X1 U10080 ( .A1(n8621), .A2(n8800), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n8717), .ZN(n8622) );
  OAI211_X1 U10081 ( .C1(n8624), .C2(n8803), .A(n8623), .B(n8622), .ZN(n8625)
         );
  AOI21_X1 U10082 ( .B1(n8626), .B2(n10099), .A(n8625), .ZN(n8627) );
  OAI21_X1 U10083 ( .B1(n8717), .B2(n8864), .A(n8627), .ZN(P2_U3269) );
  XNOR2_X1 U10084 ( .A(n8629), .B(n8628), .ZN(n8870) );
  AOI22_X1 U10085 ( .A1(n8867), .A2(n10095), .B1(n8836), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n8642) );
  AND2_X1 U10086 ( .A1(n8644), .A2(n8630), .ZN(n8633) );
  OAI21_X1 U10087 ( .B1(n8633), .B2(n8632), .A(n8631), .ZN(n8635) );
  AOI21_X1 U10088 ( .B1(n8635), .B2(n10080), .A(n8634), .ZN(n8869) );
  AOI211_X1 U10089 ( .C1(n8867), .C2(n8649), .A(n10149), .B(n8636), .ZN(n8866)
         );
  NAND2_X1 U10090 ( .A1(n8866), .A2(n8637), .ZN(n8638) );
  OAI211_X1 U10091 ( .C1(n10090), .C2(n8639), .A(n8869), .B(n8638), .ZN(n8640)
         );
  NAND2_X1 U10092 ( .A1(n8640), .A2(n10093), .ZN(n8641) );
  OAI211_X1 U10093 ( .C1(n8870), .C2(n8790), .A(n8642), .B(n8641), .ZN(
        P2_U3270) );
  XNOR2_X1 U10094 ( .A(n8643), .B(n8646), .ZN(n8875) );
  OAI211_X1 U10095 ( .C1(n8646), .C2(n8645), .A(n8644), .B(n10080), .ZN(n8648)
         );
  NAND2_X1 U10096 ( .A1(n8648), .A2(n8647), .ZN(n8871) );
  AOI211_X1 U10097 ( .C1(n8873), .C2(n8665), .A(n10149), .B(n8247), .ZN(n8872)
         );
  NAND2_X1 U10098 ( .A1(n8872), .A2(n8838), .ZN(n8652) );
  AOI22_X1 U10099 ( .A1(n8650), .A2(n8800), .B1(P2_REG2_REG_25__SCAN_IN), .B2(
        n8717), .ZN(n8651) );
  OAI211_X1 U10100 ( .C1(n8653), .C2(n8803), .A(n8652), .B(n8651), .ZN(n8654)
         );
  AOI21_X1 U10101 ( .B1(n8871), .B2(n10093), .A(n8654), .ZN(n8655) );
  OAI21_X1 U10102 ( .B1(n8875), .B2(n8790), .A(n8655), .ZN(P2_U3271) );
  NAND2_X1 U10103 ( .A1(n8658), .A2(n10058), .ZN(n8659) );
  OAI211_X1 U10104 ( .C1(n8661), .C2(n8823), .A(n8660), .B(n8659), .ZN(n8879)
         );
  INV_X1 U10105 ( .A(n8879), .ZN(n8672) );
  OAI21_X1 U10106 ( .B1(n8664), .B2(n8663), .A(n8662), .ZN(n8880) );
  OAI211_X1 U10107 ( .C1(n8877), .C2(n4254), .A(n8950), .B(n8665), .ZN(n8876)
         );
  AOI22_X1 U10108 ( .A1(n8666), .A2(n8800), .B1(n8717), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U10109 ( .A1(n8667), .A2(n10095), .ZN(n8668) );
  OAI211_X1 U10110 ( .C1(n8876), .C2(n10097), .A(n8669), .B(n8668), .ZN(n8670)
         );
  AOI21_X1 U10111 ( .B1(n8880), .B2(n10099), .A(n8670), .ZN(n8671) );
  OAI21_X1 U10112 ( .B1(n8836), .B2(n8672), .A(n8671), .ZN(P2_U3272) );
  AOI21_X1 U10113 ( .B1(n8675), .B2(n8674), .A(n8673), .ZN(n8676) );
  OAI222_X1 U10114 ( .A1(n8823), .A2(n8678), .B1(n8821), .B2(n8677), .C1(n8820), .C2(n8676), .ZN(n8679) );
  INV_X1 U10115 ( .A(n8679), .ZN(n8886) );
  AOI21_X1 U10116 ( .B1(n8681), .B2(n8680), .A(n4305), .ZN(n8882) );
  AOI21_X1 U10117 ( .B1(n8883), .B2(n4466), .A(n4254), .ZN(n8884) );
  NAND2_X1 U10118 ( .A1(n8884), .A2(n8813), .ZN(n8684) );
  AOI22_X1 U10119 ( .A1(P2_REG2_REG_23__SCAN_IN), .A2(n8836), .B1(n8682), .B2(
        n8800), .ZN(n8683) );
  OAI211_X1 U10120 ( .C1(n4800), .C2(n8803), .A(n8684), .B(n8683), .ZN(n8685)
         );
  AOI21_X1 U10121 ( .B1(n8882), .B2(n10099), .A(n8685), .ZN(n8686) );
  OAI21_X1 U10122 ( .B1(n8886), .B2(n8717), .A(n8686), .ZN(P2_U3273) );
  XNOR2_X1 U10123 ( .A(n8688), .B(n8687), .ZN(n8892) );
  AOI21_X1 U10124 ( .B1(n8888), .B2(n8702), .A(n8246), .ZN(n8889) );
  INV_X1 U10125 ( .A(n8689), .ZN(n8690) );
  AOI22_X1 U10126 ( .A1(n8836), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n8690), .B2(
        n8800), .ZN(n8691) );
  OAI21_X1 U10127 ( .B1(n8692), .B2(n8803), .A(n8691), .ZN(n8699) );
  OAI211_X1 U10128 ( .C1(n8695), .C2(n8694), .A(n8693), .B(n10080), .ZN(n8697)
         );
  NOR2_X1 U10129 ( .A1(n8891), .A2(n8717), .ZN(n8698) );
  AOI211_X1 U10130 ( .C1(n8889), .C2(n8813), .A(n8699), .B(n8698), .ZN(n8700)
         );
  OAI21_X1 U10131 ( .B1(n8892), .B2(n8790), .A(n8700), .ZN(P2_U3274) );
  XOR2_X1 U10132 ( .A(n8711), .B(n8701), .Z(n8897) );
  INV_X1 U10133 ( .A(n8722), .ZN(n8704) );
  INV_X1 U10134 ( .A(n8702), .ZN(n8703) );
  AOI21_X1 U10135 ( .B1(n8893), .B2(n8704), .A(n8703), .ZN(n8894) );
  AOI22_X1 U10136 ( .A1(n8836), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n8705), .B2(
        n8800), .ZN(n8706) );
  OAI21_X1 U10137 ( .B1(n8707), .B2(n8803), .A(n8706), .ZN(n8719) );
  INV_X1 U10138 ( .A(n8738), .ZN(n8740) );
  NOR2_X1 U10139 ( .A1(n8708), .A2(n8740), .ZN(n8742) );
  INV_X1 U10140 ( .A(n8709), .ZN(n8728) );
  NOR3_X1 U10141 ( .A1(n8742), .A2(n8728), .A3(n8727), .ZN(n8726) );
  INV_X1 U10142 ( .A(n8710), .ZN(n8712) );
  OAI21_X1 U10143 ( .B1(n8726), .B2(n8712), .A(n8711), .ZN(n8713) );
  NAND2_X1 U10144 ( .A1(n8713), .A2(n4291), .ZN(n8716) );
  AOI222_X1 U10145 ( .A1(n10080), .A2(n8716), .B1(n8715), .B2(n10060), .C1(
        n8714), .C2(n10058), .ZN(n8896) );
  NOR2_X1 U10146 ( .A1(n8896), .A2(n8717), .ZN(n8718) );
  AOI211_X1 U10147 ( .C1(n8894), .C2(n8813), .A(n8719), .B(n8718), .ZN(n8720)
         );
  OAI21_X1 U10148 ( .B1(n8897), .B2(n8790), .A(n8720), .ZN(P2_U3275) );
  XNOR2_X1 U10149 ( .A(n8721), .B(n8727), .ZN(n8902) );
  AOI21_X1 U10150 ( .B1(n8898), .B2(n8751), .A(n8722), .ZN(n8899) );
  AOI22_X1 U10151 ( .A1(n8836), .A2(P2_REG2_REG_20__SCAN_IN), .B1(n8723), .B2(
        n8800), .ZN(n8724) );
  OAI21_X1 U10152 ( .B1(n8725), .B2(n8803), .A(n8724), .ZN(n8735) );
  NOR2_X1 U10153 ( .A1(n8726), .A2(n8820), .ZN(n8733) );
  OAI21_X1 U10154 ( .B1(n8742), .B2(n8728), .A(n8727), .ZN(n8732) );
  OAI22_X1 U10155 ( .A1(n8730), .A2(n8823), .B1(n8729), .B2(n8821), .ZN(n8731)
         );
  AOI21_X1 U10156 ( .B1(n8733), .B2(n8732), .A(n8731), .ZN(n8901) );
  NOR2_X1 U10157 ( .A1(n8901), .A2(n8836), .ZN(n8734) );
  AOI211_X1 U10158 ( .C1(n8899), .C2(n8813), .A(n8735), .B(n8734), .ZN(n8736)
         );
  OAI21_X1 U10159 ( .B1(n8790), .B2(n8902), .A(n8736), .ZN(P2_U3276) );
  XNOR2_X1 U10160 ( .A(n8739), .B(n8738), .ZN(n8904) );
  INV_X1 U10161 ( .A(n8904), .ZN(n8758) );
  NAND2_X1 U10162 ( .A1(n8904), .A2(n8805), .ZN(n8748) );
  AND2_X1 U10163 ( .A1(n8708), .A2(n8740), .ZN(n8741) );
  OR2_X1 U10164 ( .A1(n8742), .A2(n8741), .ZN(n8746) );
  OAI22_X1 U10165 ( .A1(n8744), .A2(n8823), .B1(n8743), .B2(n8821), .ZN(n8745)
         );
  AOI21_X1 U10166 ( .B1(n8746), .B2(n10080), .A(n8745), .ZN(n8747) );
  NAND2_X1 U10167 ( .A1(n8748), .A2(n8747), .ZN(n8908) );
  NAND2_X1 U10168 ( .A1(n8908), .A2(n10093), .ZN(n8757) );
  INV_X1 U10169 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n8750) );
  OAI22_X1 U10170 ( .A1(n10093), .A2(n8750), .B1(n8749), .B2(n10090), .ZN(
        n8754) );
  AOI21_X1 U10171 ( .B1(n8755), .B2(n8762), .A(n10149), .ZN(n8752) );
  NAND2_X1 U10172 ( .A1(n8752), .A2(n8751), .ZN(n8905) );
  NOR2_X1 U10173 ( .A1(n8905), .A2(n10097), .ZN(n8753) );
  AOI211_X1 U10174 ( .C1(n10095), .C2(n8755), .A(n8754), .B(n8753), .ZN(n8756)
         );
  OAI211_X1 U10175 ( .C1(n8758), .C2(n8810), .A(n8757), .B(n8756), .ZN(
        P2_U3277) );
  XOR2_X1 U10176 ( .A(n8759), .B(n8767), .Z(n8761) );
  AOI222_X1 U10177 ( .A1(n10080), .A2(n8761), .B1(n8760), .B2(n10060), .C1(
        n8795), .C2(n10058), .ZN(n8912) );
  INV_X1 U10178 ( .A(n8762), .ZN(n8763) );
  AOI21_X1 U10179 ( .B1(n8909), .B2(n8787), .A(n8763), .ZN(n8910) );
  AOI22_X1 U10180 ( .A1(n8717), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n8764), .B2(
        n8800), .ZN(n8765) );
  OAI21_X1 U10181 ( .B1(n8766), .B2(n8803), .A(n8765), .ZN(n8770) );
  XNOR2_X1 U10182 ( .A(n8768), .B(n8767), .ZN(n8913) );
  NOR2_X1 U10183 ( .A1(n8913), .A2(n8790), .ZN(n8769) );
  AOI211_X1 U10184 ( .C1(n8910), .C2(n8813), .A(n8770), .B(n8769), .ZN(n8771)
         );
  OAI21_X1 U10185 ( .B1(n8836), .B2(n8912), .A(n8771), .ZN(P2_U3278) );
  NOR2_X1 U10186 ( .A1(n8781), .A2(n8773), .ZN(n8774) );
  AOI21_X1 U10187 ( .B1(n8775), .B2(n8774), .A(n8820), .ZN(n8777) );
  AOI21_X1 U10188 ( .B1(n8772), .B2(n8777), .A(n8776), .ZN(n8917) );
  INV_X1 U10189 ( .A(n8778), .ZN(n8779) );
  AOI21_X1 U10190 ( .B1(n8781), .B2(n8780), .A(n8779), .ZN(n8918) );
  NAND2_X1 U10191 ( .A1(n8717), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n8782) );
  OAI21_X1 U10192 ( .B1(n10090), .B2(n8783), .A(n8782), .ZN(n8784) );
  AOI21_X1 U10193 ( .B1(n8915), .B2(n10095), .A(n8784), .ZN(n8789) );
  OR2_X1 U10194 ( .A1(n8797), .A2(n8785), .ZN(n8786) );
  AND3_X1 U10195 ( .A1(n8787), .A2(n8950), .A3(n8786), .ZN(n8914) );
  NAND2_X1 U10196 ( .A1(n8914), .A2(n8838), .ZN(n8788) );
  OAI211_X1 U10197 ( .C1(n8918), .C2(n8790), .A(n8789), .B(n8788), .ZN(n8791)
         );
  INV_X1 U10198 ( .A(n8791), .ZN(n8792) );
  OAI21_X1 U10199 ( .B1(n8836), .B2(n8917), .A(n8792), .ZN(P2_U3279) );
  XNOR2_X1 U10200 ( .A(n8793), .B(n8807), .ZN(n8796) );
  AOI222_X1 U10201 ( .A1(n10080), .A2(n8796), .B1(n8795), .B2(n10060), .C1(
        n8794), .C2(n10058), .ZN(n8922) );
  AOI21_X1 U10202 ( .B1(n8919), .B2(n8798), .A(n8797), .ZN(n8920) );
  INV_X1 U10203 ( .A(n8919), .ZN(n8804) );
  INV_X1 U10204 ( .A(n8799), .ZN(n8801) );
  AOI22_X1 U10205 ( .A1(n8717), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n8801), .B2(
        n8800), .ZN(n8802) );
  OAI21_X1 U10206 ( .B1(n8804), .B2(n8803), .A(n8802), .ZN(n8812) );
  NAND2_X1 U10207 ( .A1(n10093), .A2(n8805), .ZN(n8809) );
  OAI21_X1 U10208 ( .B1(n8808), .B2(n8807), .A(n8806), .ZN(n8923) );
  AOI21_X1 U10209 ( .B1(n8810), .B2(n8809), .A(n8923), .ZN(n8811) );
  AOI211_X1 U10210 ( .C1(n8920), .C2(n8813), .A(n8812), .B(n8811), .ZN(n8814)
         );
  OAI21_X1 U10211 ( .B1(n8836), .B2(n8922), .A(n8814), .ZN(P2_U3280) );
  INV_X1 U10212 ( .A(n6673), .ZN(n10021) );
  INV_X1 U10213 ( .A(n8815), .ZN(n8818) );
  INV_X1 U10214 ( .A(n8816), .ZN(n8817) );
  AOI21_X1 U10215 ( .B1(n8818), .B2(n7597), .A(n8817), .ZN(n8819) );
  OAI222_X1 U10216 ( .A1(n8823), .A2(n8822), .B1(n8821), .B2(n10021), .C1(
        n8820), .C2(n8819), .ZN(n10129) );
  NAND2_X1 U10217 ( .A1(n10129), .A2(n10093), .ZN(n8833) );
  OAI21_X1 U10218 ( .B1(n8825), .B2(n7597), .A(n8824), .ZN(n10131) );
  AOI22_X1 U10219 ( .A1(n10099), .A2(n10131), .B1(n10095), .B2(n6126), .ZN(
        n8832) );
  OR2_X1 U10220 ( .A1(n8826), .A2(n10128), .ZN(n8827) );
  AND3_X1 U10221 ( .A1(n8828), .A2(n8827), .A3(n8950), .ZN(n10126) );
  NOR2_X1 U10222 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(n10090), .ZN(n8829) );
  AOI21_X1 U10223 ( .B1(n8838), .B2(n10126), .A(n8829), .ZN(n8831) );
  NAND2_X1 U10224 ( .A1(n8836), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n8830) );
  NAND4_X1 U10225 ( .A1(n8833), .A2(n8832), .A3(n8831), .A4(n8830), .ZN(
        P2_U3293) );
  AOI22_X1 U10226 ( .A1(n10099), .A2(n8835), .B1(n10095), .B2(n8834), .ZN(
        n8843) );
  AOI22_X1 U10227 ( .A1(n8838), .A2(n8837), .B1(n8836), .B2(
        P2_REG2_REG_2__SCAN_IN), .ZN(n8842) );
  OAI21_X1 U10228 ( .B1(n6147), .B2(n10090), .A(n8839), .ZN(n8840) );
  NAND2_X1 U10229 ( .A1(n8840), .A2(n10093), .ZN(n8841) );
  NAND3_X1 U10230 ( .A1(n8843), .A2(n8842), .A3(n8841), .ZN(P2_U3294) );
  NAND2_X1 U10231 ( .A1(n8844), .A2(n8958), .ZN(n8845) );
  NAND2_X1 U10232 ( .A1(n8847), .A2(n8958), .ZN(n8848) );
  OAI211_X1 U10233 ( .C1(n8850), .C2(n10149), .A(n8849), .B(n8848), .ZN(n8962)
         );
  MUX2_X1 U10234 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n8962), .S(n10176), .Z(
        P2_U3550) );
  AOI21_X1 U10235 ( .B1(n8958), .B2(n8852), .A(n8851), .ZN(n8853) );
  OAI211_X1 U10236 ( .C1(n8855), .C2(n8949), .A(n8854), .B(n8853), .ZN(n8963)
         );
  MUX2_X1 U10237 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n8963), .S(n10176), .Z(
        P2_U3549) );
  AOI22_X1 U10238 ( .A1(n8857), .A2(n8950), .B1(n8958), .B2(n8856), .ZN(n8858)
         );
  OAI211_X1 U10239 ( .C1(n8860), .C2(n8949), .A(n8859), .B(n8858), .ZN(n8964)
         );
  MUX2_X1 U10240 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n8964), .S(n10176), .Z(
        P2_U3548) );
  AOI22_X1 U10241 ( .A1(n8862), .A2(n8950), .B1(n8958), .B2(n8861), .ZN(n8863)
         );
  OAI211_X1 U10242 ( .C1(n8865), .C2(n8949), .A(n8864), .B(n8863), .ZN(n8965)
         );
  MUX2_X1 U10243 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n8965), .S(n10176), .Z(
        P2_U3547) );
  AOI21_X1 U10244 ( .B1(n8958), .B2(n8867), .A(n8866), .ZN(n8868) );
  OAI211_X1 U10245 ( .C1(n8870), .C2(n8949), .A(n8869), .B(n8868), .ZN(n8966)
         );
  MUX2_X1 U10246 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n8966), .S(n10176), .Z(
        P2_U3546) );
  AOI211_X1 U10247 ( .C1(n8958), .C2(n8873), .A(n8872), .B(n8871), .ZN(n8874)
         );
  OAI21_X1 U10248 ( .B1(n8875), .B2(n8949), .A(n8874), .ZN(n8967) );
  MUX2_X1 U10249 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n8967), .S(n10176), .Z(
        P2_U3545) );
  OAI21_X1 U10250 ( .B1(n8877), .B2(n10159), .A(n8876), .ZN(n8878) );
  INV_X1 U10251 ( .A(n8881), .ZN(n8968) );
  MUX2_X1 U10252 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n8968), .S(n10176), .Z(
        P2_U3544) );
  INV_X1 U10253 ( .A(n8882), .ZN(n8887) );
  AOI22_X1 U10254 ( .A1(n8884), .A2(n8950), .B1(n8958), .B2(n8883), .ZN(n8885)
         );
  OAI211_X1 U10255 ( .C1(n8887), .C2(n8949), .A(n8886), .B(n8885), .ZN(n8969)
         );
  MUX2_X1 U10256 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n8969), .S(n10176), .Z(
        P2_U3543) );
  AOI22_X1 U10257 ( .A1(n8889), .A2(n8950), .B1(n8958), .B2(n8888), .ZN(n8890)
         );
  OAI211_X1 U10258 ( .C1(n8892), .C2(n8949), .A(n8891), .B(n8890), .ZN(n8970)
         );
  MUX2_X1 U10259 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n8970), .S(n10176), .Z(
        P2_U3542) );
  AOI22_X1 U10260 ( .A1(n8894), .A2(n8950), .B1(n8958), .B2(n8893), .ZN(n8895)
         );
  OAI211_X1 U10261 ( .C1(n8949), .C2(n8897), .A(n8896), .B(n8895), .ZN(n8971)
         );
  MUX2_X1 U10262 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n8971), .S(n10176), .Z(
        P2_U3541) );
  AOI22_X1 U10263 ( .A1(n8899), .A2(n8950), .B1(n8958), .B2(n8898), .ZN(n8900)
         );
  OAI211_X1 U10264 ( .C1(n8949), .C2(n8902), .A(n8901), .B(n8900), .ZN(n8972)
         );
  MUX2_X1 U10265 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n8972), .S(n10176), .Z(
        P2_U3540) );
  NAND2_X1 U10266 ( .A1(n8904), .A2(n8903), .ZN(n8906) );
  OAI211_X1 U10267 ( .C1(n4824), .C2(n10159), .A(n8906), .B(n8905), .ZN(n8907)
         );
  MUX2_X1 U10268 ( .A(n8973), .B(P2_REG1_REG_19__SCAN_IN), .S(n10174), .Z(
        P2_U3539) );
  AOI22_X1 U10269 ( .A1(n8910), .A2(n8950), .B1(n8958), .B2(n8909), .ZN(n8911)
         );
  OAI211_X1 U10270 ( .C1(n8949), .C2(n8913), .A(n8912), .B(n8911), .ZN(n8974)
         );
  MUX2_X1 U10271 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n8974), .S(n10176), .Z(
        P2_U3538) );
  AOI21_X1 U10272 ( .B1(n8958), .B2(n8915), .A(n8914), .ZN(n8916) );
  OAI211_X1 U10273 ( .C1(n8918), .C2(n8949), .A(n8917), .B(n8916), .ZN(n8975)
         );
  MUX2_X1 U10274 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n8975), .S(n10176), .Z(
        P2_U3537) );
  AOI22_X1 U10275 ( .A1(n8920), .A2(n8950), .B1(n8958), .B2(n8919), .ZN(n8921)
         );
  OAI211_X1 U10276 ( .C1(n8949), .C2(n8923), .A(n8922), .B(n8921), .ZN(n8976)
         );
  MUX2_X1 U10277 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n8976), .S(n10176), .Z(
        P2_U3536) );
  AOI22_X1 U10278 ( .A1(n8925), .A2(n8950), .B1(n8958), .B2(n8924), .ZN(n8926)
         );
  OAI211_X1 U10279 ( .C1(n8949), .C2(n8928), .A(n8927), .B(n8926), .ZN(n8977)
         );
  MUX2_X1 U10280 ( .A(P2_REG1_REG_15__SCAN_IN), .B(n8977), .S(n10176), .Z(
        P2_U3535) );
  AOI22_X1 U10281 ( .A1(n8930), .A2(n8950), .B1(n8958), .B2(n8929), .ZN(n8931)
         );
  OAI211_X1 U10282 ( .C1(n8933), .C2(n8949), .A(n8932), .B(n8931), .ZN(n8978)
         );
  MUX2_X1 U10283 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n8978), .S(n10176), .Z(
        P2_U3534) );
  AOI22_X1 U10284 ( .A1(n8935), .A2(n8950), .B1(n8958), .B2(n8934), .ZN(n8936)
         );
  OAI21_X1 U10285 ( .B1(n8937), .B2(n10158), .A(n8936), .ZN(n8938) );
  OR2_X1 U10286 ( .A1(n8939), .A2(n8938), .ZN(n8979) );
  MUX2_X1 U10287 ( .A(P2_REG1_REG_13__SCAN_IN), .B(n8979), .S(n10176), .Z(
        P2_U3533) );
  AOI21_X1 U10288 ( .B1(n8958), .B2(n8941), .A(n8940), .ZN(n8942) );
  OAI211_X1 U10289 ( .C1(n8944), .C2(n8949), .A(n8943), .B(n8942), .ZN(n8980)
         );
  MUX2_X1 U10290 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n8980), .S(n10176), .Z(
        P2_U3532) );
  AOI22_X1 U10291 ( .A1(n8945), .A2(n8950), .B1(n8958), .B2(n10051), .ZN(n8946) );
  OAI211_X1 U10292 ( .C1(n8949), .C2(n8948), .A(n8947), .B(n8946), .ZN(n8981)
         );
  MUX2_X1 U10293 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n8981), .S(n10176), .Z(
        P2_U3531) );
  AOI22_X1 U10294 ( .A1(n8951), .A2(n8950), .B1(n8958), .B2(n10015), .ZN(n8952) );
  OAI211_X1 U10295 ( .C1(n8954), .C2(n10158), .A(n8953), .B(n8952), .ZN(n8982)
         );
  MUX2_X1 U10296 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n8982), .S(n10176), .Z(
        P2_U3530) );
  INV_X1 U10297 ( .A(n8955), .ZN(n8960) );
  AOI21_X1 U10298 ( .B1(n8958), .B2(n8957), .A(n8956), .ZN(n8959) );
  OAI211_X1 U10299 ( .C1(n8961), .C2(n10158), .A(n8960), .B(n8959), .ZN(n8983)
         );
  MUX2_X1 U10300 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n8983), .S(n10176), .Z(
        P2_U3529) );
  MUX2_X1 U10301 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n8962), .S(n10166), .Z(
        P2_U3518) );
  MUX2_X1 U10302 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n8963), .S(n10166), .Z(
        P2_U3517) );
  MUX2_X1 U10303 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n8964), .S(n10166), .Z(
        P2_U3516) );
  MUX2_X1 U10304 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n8965), .S(n10166), .Z(
        P2_U3515) );
  MUX2_X1 U10305 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n8966), .S(n10166), .Z(
        P2_U3514) );
  MUX2_X1 U10306 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n8967), .S(n10166), .Z(
        P2_U3513) );
  MUX2_X1 U10307 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n8968), .S(n10166), .Z(
        P2_U3512) );
  MUX2_X1 U10308 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n8969), .S(n10166), .Z(
        P2_U3511) );
  MUX2_X1 U10309 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n8970), .S(n10166), .Z(
        P2_U3510) );
  MUX2_X1 U10310 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n8971), .S(n10166), .Z(
        P2_U3509) );
  MUX2_X1 U10311 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n8972), .S(n10166), .Z(
        P2_U3508) );
  MUX2_X1 U10312 ( .A(n8973), .B(P2_REG0_REG_19__SCAN_IN), .S(n10165), .Z(
        P2_U3507) );
  MUX2_X1 U10313 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n8974), .S(n10166), .Z(
        P2_U3505) );
  MUX2_X1 U10314 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n8975), .S(n10166), .Z(
        P2_U3502) );
  MUX2_X1 U10315 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n8976), .S(n10166), .Z(
        P2_U3499) );
  MUX2_X1 U10316 ( .A(P2_REG0_REG_15__SCAN_IN), .B(n8977), .S(n10166), .Z(
        P2_U3496) );
  MUX2_X1 U10317 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8978), .S(n10166), .Z(
        P2_U3493) );
  MUX2_X1 U10318 ( .A(n8979), .B(P2_REG0_REG_13__SCAN_IN), .S(n10165), .Z(
        P2_U3490) );
  MUX2_X1 U10319 ( .A(P2_REG0_REG_12__SCAN_IN), .B(n8980), .S(n10166), .Z(
        P2_U3487) );
  MUX2_X1 U10320 ( .A(P2_REG0_REG_11__SCAN_IN), .B(n8981), .S(n10166), .Z(
        P2_U3484) );
  MUX2_X1 U10321 ( .A(P2_REG0_REG_10__SCAN_IN), .B(n8982), .S(n10166), .Z(
        P2_U3481) );
  MUX2_X1 U10322 ( .A(P2_REG0_REG_9__SCAN_IN), .B(n8983), .S(n10166), .Z(
        P2_U3478) );
  INV_X1 U10323 ( .A(n8984), .ZN(n9783) );
  NOR4_X1 U10324 ( .A1(n8985), .A2(P2_IR_REG_30__SCAN_IN), .A3(n6084), .A4(
        P2_U3152), .ZN(n8986) );
  AOI21_X1 U10325 ( .B1(n8989), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n8986), .ZN(
        n8987) );
  OAI21_X1 U10326 ( .B1(n9783), .B2(n4249), .A(n8987), .ZN(P2_U3327) );
  AOI22_X1 U10327 ( .A1(n8988), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_30__SCAN_IN), .B2(n8989), .ZN(n8990) );
  OAI21_X1 U10328 ( .B1(n8991), .B2(n4249), .A(n8990), .ZN(P2_U3328) );
  INV_X1 U10329 ( .A(n8992), .ZN(n9784) );
  OAI222_X1 U10330 ( .A1(n9000), .A2(n9665), .B1(n4249), .B2(n9784), .C1(n8993), .C2(P2_U3152), .ZN(P2_U3329) );
  NAND2_X1 U10331 ( .A1(n9788), .A2(n8994), .ZN(n8996) );
  OAI211_X1 U10332 ( .C1(n9000), .C2(n9757), .A(n8996), .B(n8995), .ZN(
        P2_U3330) );
  INV_X1 U10333 ( .A(n8997), .ZN(n9795) );
  OAI222_X1 U10334 ( .A1(n8998), .A2(P2_U3152), .B1(n4249), .B2(n9795), .C1(
        n9733), .C2(n9000), .ZN(P2_U3331) );
  INV_X1 U10335 ( .A(n8999), .ZN(n9797) );
  OAI222_X1 U10336 ( .A1(n9002), .A2(P2_U3152), .B1(n4249), .B2(n9797), .C1(
        n9001), .C2(n9000), .ZN(P2_U3332) );
  MUX2_X1 U10337 ( .A(n9004), .B(n9003), .S(P2_STATE_REG_SCAN_IN), .Z(P2_U3358) );
  NAND2_X1 U10338 ( .A1(n9315), .A2(n9016), .ZN(n9007) );
  NAND2_X1 U10339 ( .A1(n9307), .A2(n9137), .ZN(n9006) );
  OAI211_X1 U10340 ( .C1(P1_STATE_REG_SCAN_IN), .C2(n9008), .A(n9007), .B(
        n9006), .ZN(n9009) );
  AOI21_X1 U10341 ( .B1(n9271), .B2(n9142), .A(n9009), .ZN(n9010) );
  OAI211_X1 U10342 ( .C1(n4371), .C2(n9145), .A(n9011), .B(n9010), .ZN(
        P1_U3212) );
  OR2_X1 U10343 ( .A1(n9013), .A2(n9012), .ZN(n9085) );
  NAND2_X1 U10344 ( .A1(n9013), .A2(n9012), .ZN(n9045) );
  NAND2_X1 U10345 ( .A1(n9085), .A2(n9045), .ZN(n9014) );
  XNOR2_X1 U10346 ( .A(n9014), .B(n9043), .ZN(n9021) );
  INV_X1 U10347 ( .A(n9015), .ZN(n9378) );
  AOI22_X1 U10348 ( .A1(n9378), .A2(n9137), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9018) );
  NAND2_X1 U10349 ( .A1(n9402), .A2(n9016), .ZN(n9017) );
  OAI211_X1 U10350 ( .C1(n9053), .C2(n9037), .A(n9018), .B(n9017), .ZN(n9019)
         );
  AOI21_X1 U10351 ( .B1(n9541), .B2(n9130), .A(n9019), .ZN(n9020) );
  OAI21_X1 U10352 ( .B1(n9021), .B2(n9132), .A(n9020), .ZN(P1_U3214) );
  INV_X1 U10353 ( .A(n9561), .ZN(n9435) );
  OR2_X1 U10354 ( .A1(n9023), .A2(n9022), .ZN(n9120) );
  NAND2_X1 U10355 ( .A1(n9120), .A2(n9119), .ZN(n9118) );
  NAND2_X1 U10356 ( .A1(n9023), .A2(n9022), .ZN(n9122) );
  NAND2_X1 U10357 ( .A1(n9024), .A2(n9094), .ZN(n9025) );
  AOI21_X1 U10358 ( .B1(n9118), .B2(n9122), .A(n9025), .ZN(n9097) );
  AND3_X1 U10359 ( .A1(n9118), .A2(n9122), .A3(n9025), .ZN(n9026) );
  OAI21_X1 U10360 ( .B1(n9097), .B2(n9026), .A(n9134), .ZN(n9030) );
  NAND2_X1 U10361 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9205) );
  OAI21_X1 U10362 ( .B1(n9485), .B2(n9139), .A(n9205), .ZN(n9028) );
  NOR2_X1 U10363 ( .A1(n9128), .A2(n9443), .ZN(n9027) );
  AOI211_X1 U10364 ( .C1(n9142), .C2(n9440), .A(n9028), .B(n9027), .ZN(n9029)
         );
  OAI211_X1 U10365 ( .C1(n9435), .C2(n9145), .A(n9030), .B(n9029), .ZN(
        P1_U3217) );
  OAI21_X1 U10366 ( .B1(n9033), .B2(n9032), .A(n9031), .ZN(n9034) );
  NAND2_X1 U10367 ( .A1(n9034), .A2(n9134), .ZN(n9042) );
  OAI22_X1 U10368 ( .A1(n9036), .A2(n9139), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9035), .ZN(n9040) );
  NOR2_X1 U10369 ( .A1(n9038), .A2(n9037), .ZN(n9039) );
  AOI211_X1 U10370 ( .C1(n9137), .C2(n9411), .A(n9040), .B(n9039), .ZN(n9041)
         );
  OAI211_X1 U10371 ( .C1(n9414), .C2(n9145), .A(n9042), .B(n9041), .ZN(
        P1_U3221) );
  INV_X1 U10372 ( .A(n9043), .ZN(n9044) );
  NAND2_X1 U10373 ( .A1(n9045), .A2(n9044), .ZN(n9086) );
  AND2_X1 U10374 ( .A1(n9047), .A2(n9046), .ZN(n9084) );
  NAND3_X1 U10375 ( .A1(n9086), .A2(n9084), .A3(n9085), .ZN(n9083) );
  AND3_X1 U10376 ( .A1(n9083), .A2(n9048), .A3(n9047), .ZN(n9049) );
  INV_X1 U10377 ( .A(n9051), .ZN(n9349) );
  AOI22_X1 U10378 ( .A1(n9349), .A2(n9137), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9052) );
  OAI21_X1 U10379 ( .B1(n9053), .B2(n9139), .A(n9052), .ZN(n9054) );
  AOI21_X1 U10380 ( .B1(n9142), .B2(n9315), .A(n9054), .ZN(n9055) );
  OAI211_X1 U10381 ( .C1(n9352), .C2(n9145), .A(n9056), .B(n9055), .ZN(
        P1_U3223) );
  NOR2_X1 U10382 ( .A1(n9058), .A2(n9057), .ZN(n9062) );
  INV_X1 U10383 ( .A(n9058), .ZN(n9060) );
  OAI22_X1 U10384 ( .A1(n9062), .A2(n9061), .B1(n9060), .B2(n9059), .ZN(n9065)
         );
  NAND2_X1 U10385 ( .A1(n9063), .A2(n9074), .ZN(n9064) );
  NOR2_X1 U10386 ( .A1(n9065), .A2(n9064), .ZN(n9077) );
  AOI21_X1 U10387 ( .B1(n9065), .B2(n9064), .A(n9077), .ZN(n9073) );
  INV_X1 U10388 ( .A(n9125), .ZN(n9452) );
  AND2_X1 U10389 ( .A1(P1_U3084), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n9897) );
  NOR2_X1 U10390 ( .A1(n9139), .A2(n9067), .ZN(n9068) );
  AOI211_X1 U10391 ( .C1(n9142), .C2(n9452), .A(n9897), .B(n9068), .ZN(n9069)
         );
  OAI21_X1 U10392 ( .B1(n9070), .B2(n9128), .A(n9069), .ZN(n9071) );
  AOI21_X1 U10393 ( .B1(n9580), .B2(n9130), .A(n9071), .ZN(n9072) );
  OAI21_X1 U10394 ( .B1(n9073), .B2(n9132), .A(n9072), .ZN(P1_U3224) );
  INV_X1 U10395 ( .A(n9573), .ZN(n9476) );
  INV_X1 U10396 ( .A(n9074), .ZN(n9076) );
  NOR3_X1 U10397 ( .A1(n9077), .A2(n9076), .A3(n9075), .ZN(n9078) );
  OAI21_X1 U10398 ( .B1(n9078), .B2(n4312), .A(n9134), .ZN(n9082) );
  NOR2_X1 U10399 ( .A1(n9730), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9909) );
  AOI21_X1 U10400 ( .B1(n9441), .B2(n9142), .A(n9909), .ZN(n9079) );
  OAI21_X1 U10401 ( .B1(n9483), .B2(n9139), .A(n9079), .ZN(n9080) );
  AOI21_X1 U10402 ( .B1(n9473), .B2(n9137), .A(n9080), .ZN(n9081) );
  OAI211_X1 U10403 ( .C1(n9476), .C2(n9145), .A(n9082), .B(n9081), .ZN(
        P1_U3226) );
  INV_X1 U10404 ( .A(n9083), .ZN(n9088) );
  AOI21_X1 U10405 ( .B1(n9086), .B2(n9085), .A(n9084), .ZN(n9087) );
  OAI21_X1 U10406 ( .B1(n9088), .B2(n9087), .A(n9134), .ZN(n9093) );
  AOI22_X1 U10407 ( .A1(n9364), .A2(n9137), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9089) );
  OAI21_X1 U10408 ( .B1(n9090), .B2(n9139), .A(n9089), .ZN(n9091) );
  AOI21_X1 U10409 ( .B1(n9358), .B2(n9142), .A(n9091), .ZN(n9092) );
  OAI211_X1 U10410 ( .C1(n4757), .C2(n9145), .A(n9093), .B(n9092), .ZN(
        P1_U3227) );
  INV_X1 U10411 ( .A(n9556), .ZN(n9426) );
  INV_X1 U10412 ( .A(n9094), .ZN(n9096) );
  NOR3_X1 U10413 ( .A1(n9097), .A2(n9096), .A3(n9095), .ZN(n9100) );
  INV_X1 U10414 ( .A(n9098), .ZN(n9099) );
  OAI21_X1 U10415 ( .B1(n9100), .B2(n9099), .A(n9134), .ZN(n9105) );
  OAI22_X1 U10416 ( .A1(n9124), .A2(n9139), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9101), .ZN(n9103) );
  NOR2_X1 U10417 ( .A1(n9128), .A2(n9423), .ZN(n9102) );
  AOI211_X1 U10418 ( .C1(n9419), .C2(n9142), .A(n9103), .B(n9102), .ZN(n9104)
         );
  OAI211_X1 U10419 ( .C1(n9426), .C2(n9145), .A(n9105), .B(n9104), .ZN(
        P1_U3231) );
  INV_X1 U10420 ( .A(n9106), .ZN(n9108) );
  NAND2_X1 U10421 ( .A1(n9108), .A2(n9107), .ZN(n9110) );
  XNOR2_X1 U10422 ( .A(n9110), .B(n9109), .ZN(n9111) );
  NAND2_X1 U10423 ( .A1(n9111), .A2(n9134), .ZN(n9117) );
  NOR2_X1 U10424 ( .A1(n9391), .A2(n9128), .ZN(n9115) );
  OAI22_X1 U10425 ( .A1(n9113), .A2(n9139), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n9112), .ZN(n9114) );
  AOI211_X1 U10426 ( .C1(n9387), .C2(n9142), .A(n9115), .B(n9114), .ZN(n9116)
         );
  OAI211_X1 U10427 ( .C1(n9394), .C2(n9145), .A(n9117), .B(n9116), .ZN(
        P1_U3233) );
  INV_X1 U10428 ( .A(n9118), .ZN(n9123) );
  AOI21_X1 U10429 ( .B1(n9120), .B2(n9122), .A(n9119), .ZN(n9121) );
  AOI21_X1 U10430 ( .B1(n9123), .B2(n9122), .A(n9121), .ZN(n9133) );
  NOR2_X1 U10431 ( .A1(n9712), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9926) );
  NOR2_X1 U10432 ( .A1(n9139), .A2(n9125), .ZN(n9126) );
  AOI211_X1 U10433 ( .C1(n9450), .C2(n9142), .A(n9926), .B(n9126), .ZN(n9127)
         );
  OAI21_X1 U10434 ( .B1(n9461), .B2(n9128), .A(n9127), .ZN(n9129) );
  AOI21_X1 U10435 ( .B1(n9568), .B2(n9130), .A(n9129), .ZN(n9131) );
  OAI21_X1 U10436 ( .B1(n9133), .B2(n9132), .A(n9131), .ZN(P1_U3236) );
  INV_X1 U10437 ( .A(n9527), .ZN(n9331) );
  OAI211_X1 U10438 ( .C1(n4265), .C2(n9136), .A(n9135), .B(n9134), .ZN(n9144)
         );
  AOI22_X1 U10439 ( .A1(n9329), .A2(n9137), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9138) );
  OAI21_X1 U10440 ( .B1(n9140), .B2(n9139), .A(n9138), .ZN(n9141) );
  AOI21_X1 U10441 ( .B1(n9322), .B2(n9142), .A(n9141), .ZN(n9143) );
  OAI211_X1 U10442 ( .C1(n9331), .C2(n9145), .A(n9144), .B(n9143), .ZN(
        P1_U3238) );
  MUX2_X1 U10443 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9268), .S(P1_U4006), .Z(
        P1_U3585) );
  MUX2_X1 U10444 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n9271), .S(P1_U4006), .Z(
        P1_U3583) );
  MUX2_X1 U10445 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9322), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10446 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9315), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10447 ( .A(n9358), .B(P1_DATAO_REG_25__SCAN_IN), .S(n9159), .Z(
        P1_U3580) );
  MUX2_X1 U10448 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9374), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10449 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n9387), .S(P1_U4006), .Z(
        P1_U3578) );
  MUX2_X1 U10450 ( .A(n9402), .B(P1_DATAO_REG_22__SCAN_IN), .S(n9159), .Z(
        P1_U3577) );
  MUX2_X1 U10451 ( .A(n9419), .B(P1_DATAO_REG_21__SCAN_IN), .S(n9159), .Z(
        P1_U3576) );
  MUX2_X1 U10452 ( .A(n9440), .B(P1_DATAO_REG_20__SCAN_IN), .S(n9159), .Z(
        P1_U3575) );
  MUX2_X1 U10453 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9450), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10454 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9441), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10455 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9452), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10456 ( .A(n9223), .B(P1_DATAO_REG_16__SCAN_IN), .S(n9159), .Z(
        P1_U3571) );
  MUX2_X1 U10457 ( .A(n9146), .B(P1_DATAO_REG_15__SCAN_IN), .S(n9159), .Z(
        P1_U3570) );
  MUX2_X1 U10458 ( .A(n9147), .B(P1_DATAO_REG_14__SCAN_IN), .S(n9159), .Z(
        P1_U3569) );
  MUX2_X1 U10459 ( .A(n9148), .B(P1_DATAO_REG_13__SCAN_IN), .S(n9159), .Z(
        P1_U3568) );
  MUX2_X1 U10460 ( .A(n9149), .B(P1_DATAO_REG_12__SCAN_IN), .S(n9159), .Z(
        P1_U3567) );
  MUX2_X1 U10461 ( .A(n9150), .B(P1_DATAO_REG_11__SCAN_IN), .S(n9159), .Z(
        P1_U3566) );
  MUX2_X1 U10462 ( .A(n9151), .B(P1_DATAO_REG_10__SCAN_IN), .S(n9159), .Z(
        P1_U3565) );
  MUX2_X1 U10463 ( .A(n9152), .B(P1_DATAO_REG_9__SCAN_IN), .S(n9159), .Z(
        P1_U3564) );
  MUX2_X1 U10464 ( .A(n9153), .B(P1_DATAO_REG_8__SCAN_IN), .S(n9159), .Z(
        P1_U3563) );
  MUX2_X1 U10465 ( .A(n9154), .B(P1_DATAO_REG_7__SCAN_IN), .S(n9159), .Z(
        P1_U3562) );
  MUX2_X1 U10466 ( .A(n5830), .B(P1_DATAO_REG_6__SCAN_IN), .S(n9159), .Z(
        P1_U3561) );
  MUX2_X1 U10467 ( .A(n9155), .B(P1_DATAO_REG_5__SCAN_IN), .S(n9159), .Z(
        P1_U3560) );
  MUX2_X1 U10468 ( .A(n9156), .B(P1_DATAO_REG_4__SCAN_IN), .S(n9159), .Z(
        P1_U3559) );
  MUX2_X1 U10469 ( .A(n9157), .B(P1_DATAO_REG_3__SCAN_IN), .S(n9159), .Z(
        P1_U3558) );
  MUX2_X1 U10470 ( .A(n9158), .B(P1_DATAO_REG_2__SCAN_IN), .S(n9159), .Z(
        P1_U3557) );
  MUX2_X1 U10471 ( .A(n9160), .B(P1_DATAO_REG_1__SCAN_IN), .S(n9159), .Z(
        P1_U3556) );
  MUX2_X1 U10472 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9161), .S(P1_U4006), .Z(
        P1_U3555) );
  NAND2_X1 U10473 ( .A1(n9927), .A2(P1_ADDR_REG_7__SCAN_IN), .ZN(n9175) );
  AOI21_X1 U10474 ( .B1(n9886), .B2(n9163), .A(n9162), .ZN(n9174) );
  OAI21_X1 U10475 ( .B1(n9166), .B2(n9165), .A(n9164), .ZN(n9167) );
  NAND2_X1 U10476 ( .A1(n9167), .A2(n9911), .ZN(n9173) );
  OAI21_X1 U10477 ( .B1(n9170), .B2(n9169), .A(n9168), .ZN(n9171) );
  NAND2_X1 U10478 ( .A1(n9929), .A2(n9171), .ZN(n9172) );
  NAND4_X1 U10479 ( .A1(n9175), .A2(n9174), .A3(n9173), .A4(n9172), .ZN(
        P1_U3248) );
  MUX2_X1 U10480 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n9462), .S(n9183), .Z(n9930) );
  NAND2_X1 U10481 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n9184), .ZN(n9181) );
  MUX2_X1 U10482 ( .A(n5423), .B(P1_REG2_REG_17__SCAN_IN), .S(n9184), .Z(n9176) );
  INV_X1 U10483 ( .A(n9176), .ZN(n9916) );
  MUX2_X1 U10484 ( .A(P1_REG2_REG_16__SCAN_IN), .B(n9640), .S(n9185), .Z(n9902) );
  MUX2_X1 U10485 ( .A(n8004), .B(P1_REG2_REG_12__SCAN_IN), .S(n9839), .Z(n9847) );
  AOI21_X1 U10486 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n9839), .A(n9845), .ZN(
        n9865) );
  MUX2_X1 U10487 ( .A(n7897), .B(P1_REG2_REG_13__SCAN_IN), .S(n9856), .Z(n9864) );
  NOR2_X1 U10488 ( .A1(n9865), .A2(n9864), .ZN(n9862) );
  NAND2_X1 U10489 ( .A1(n9885), .A2(n9179), .ZN(n9180) );
  NAND2_X1 U10490 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n9890), .ZN(n9889) );
  NAND2_X1 U10491 ( .A1(n9180), .A2(n9889), .ZN(n9903) );
  NAND2_X1 U10492 ( .A1(n9902), .A2(n9903), .ZN(n9901) );
  OAI21_X1 U10493 ( .B1(n9895), .B2(n9640), .A(n9901), .ZN(n9915) );
  NAND2_X1 U10494 ( .A1(n9916), .A2(n9915), .ZN(n9914) );
  NAND2_X1 U10495 ( .A1(n9181), .A2(n9914), .ZN(n9931) );
  NAND2_X1 U10496 ( .A1(n9930), .A2(n9931), .ZN(n9928) );
  OAI21_X1 U10497 ( .B1(n9462), .B2(n9924), .A(n9928), .ZN(n9182) );
  INV_X1 U10498 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9197) );
  AOI22_X1 U10499 ( .A1(n9183), .A2(n9197), .B1(P1_REG1_REG_18__SCAN_IN), .B2(
        n9924), .ZN(n9922) );
  INV_X1 U10500 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9196) );
  AOI22_X1 U10501 ( .A1(P1_REG1_REG_17__SCAN_IN), .A2(n9184), .B1(n9907), .B2(
        n9196), .ZN(n9913) );
  INV_X1 U10502 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n9195) );
  AOI22_X1 U10503 ( .A1(P1_REG1_REG_16__SCAN_IN), .A2(n9185), .B1(n9895), .B2(
        n9195), .ZN(n9900) );
  XNOR2_X1 U10504 ( .A(n9839), .B(n9188), .ZN(n9836) );
  NAND2_X1 U10505 ( .A1(n9837), .A2(n9836), .ZN(n9835) );
  XNOR2_X1 U10506 ( .A(n9856), .B(n9189), .ZN(n9853) );
  NAND2_X1 U10507 ( .A1(n9854), .A2(n9853), .ZN(n9852) );
  OAI21_X1 U10508 ( .B1(n9856), .B2(P1_REG1_REG_13__SCAN_IN), .A(n9852), .ZN(
        n9872) );
  XNOR2_X1 U10509 ( .A(n9191), .B(n9190), .ZN(n9871) );
  INV_X1 U10510 ( .A(n9193), .ZN(n9192) );
  NAND2_X1 U10511 ( .A1(n9192), .A2(n9885), .ZN(n9194) );
  XNOR2_X1 U10512 ( .A(n9193), .B(n9885), .ZN(n9888) );
  NAND2_X1 U10513 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n9888), .ZN(n9887) );
  NAND2_X1 U10514 ( .A1(n9194), .A2(n9887), .ZN(n9899) );
  NAND2_X1 U10515 ( .A1(n9900), .A2(n9899), .ZN(n9898) );
  OAI21_X1 U10516 ( .B1(n9895), .B2(n9195), .A(n9898), .ZN(n9912) );
  NAND2_X1 U10517 ( .A1(n9913), .A2(n9912), .ZN(n9910) );
  OAI21_X1 U10518 ( .B1(n9907), .B2(n9196), .A(n9910), .ZN(n9921) );
  NOR2_X1 U10519 ( .A1(n9922), .A2(n9921), .ZN(n9920) );
  XOR2_X1 U10520 ( .A(n9198), .B(P1_REG1_REG_19__SCAN_IN), .Z(n9202) );
  INV_X1 U10521 ( .A(n9202), .ZN(n9199) );
  NAND2_X1 U10522 ( .A1(n9199), .A2(n9911), .ZN(n9200) );
  AOI22_X1 U10523 ( .A1(n9203), .A2(n9929), .B1(n9911), .B2(n9202), .ZN(n9204)
         );
  OAI211_X1 U10524 ( .C1(n9207), .C2(n9877), .A(n9206), .B(n9205), .ZN(
        P1_U3260) );
  INV_X1 U10525 ( .A(n9568), .ZN(n9459) );
  NAND2_X1 U10526 ( .A1(n9455), .A2(n9459), .ZN(n9456) );
  AND2_X2 U10527 ( .A1(n9407), .A2(n9414), .ZN(n9408) );
  XOR2_X1 U10528 ( .A(n9216), .B(n9496), .Z(n9494) );
  NAND2_X1 U10529 ( .A1(n9494), .A2(n9491), .ZN(n9215) );
  NOR2_X1 U10530 ( .A1(n9211), .A2(n9210), .ZN(n9212) );
  NOR2_X1 U10531 ( .A1(n9484), .A2(n9212), .ZN(n9269) );
  NAND2_X1 U10532 ( .A1(n9269), .A2(n9213), .ZN(n9499) );
  NOR2_X1 U10533 ( .A1(n4246), .A2(n9499), .ZN(n9218) );
  AOI21_X1 U10534 ( .B1(n4246), .B2(P1_REG2_REG_31__SCAN_IN), .A(n9218), .ZN(
        n9214) );
  OAI211_X1 U10535 ( .C1(n9475), .C2(n9496), .A(n9215), .B(n9214), .ZN(
        P1_U3261) );
  INV_X1 U10536 ( .A(n9217), .ZN(n9501) );
  INV_X1 U10537 ( .A(n9216), .ZN(n9498) );
  NAND2_X1 U10538 ( .A1(n9217), .A2(n9275), .ZN(n9497) );
  NAND3_X1 U10539 ( .A1(n9498), .A2(n9491), .A3(n9497), .ZN(n9220) );
  AOI21_X1 U10540 ( .B1(n4246), .B2(P1_REG2_REG_30__SCAN_IN), .A(n9218), .ZN(
        n9219) );
  OAI211_X1 U10541 ( .C1(n9501), .C2(n9475), .A(n9220), .B(n9219), .ZN(
        P1_U3262) );
  NAND2_X1 U10542 ( .A1(n9222), .A2(n9221), .ZN(n9225) );
  NAND2_X1 U10543 ( .A1(n9580), .A2(n9223), .ZN(n9224) );
  AND2_X1 U10544 ( .A1(n9573), .A2(n9452), .ZN(n9227) );
  OR2_X1 U10545 ( .A1(n9573), .A2(n9452), .ZN(n9226) );
  NAND2_X1 U10546 ( .A1(n9561), .A2(n9450), .ZN(n9228) );
  NAND2_X1 U10547 ( .A1(n9229), .A2(n9228), .ZN(n9428) );
  INV_X1 U10548 ( .A(n9428), .ZN(n9231) );
  AOI21_X2 U10549 ( .B1(n9231), .B2(n4264), .A(n9230), .ZN(n9406) );
  NAND2_X1 U10550 ( .A1(n9552), .A2(n9419), .ZN(n9232) );
  OR2_X1 U10551 ( .A1(n9546), .A2(n9402), .ZN(n9233) );
  AND2_X1 U10552 ( .A1(n9541), .A2(n9387), .ZN(n9235) );
  OAI21_X1 U10553 ( .B1(n9381), .B2(n9235), .A(n9234), .ZN(n9337) );
  NAND2_X1 U10554 ( .A1(n9366), .A2(n9374), .ZN(n9338) );
  NAND3_X1 U10555 ( .A1(n9340), .A2(n9356), .A3(n9338), .ZN(n9236) );
  OAI21_X1 U10556 ( .B1(n9358), .B2(n9533), .A(n9236), .ZN(n9237) );
  OR2_X1 U10557 ( .A1(n9520), .A2(n9322), .ZN(n9242) );
  NAND2_X1 U10558 ( .A1(n9514), .A2(n9271), .ZN(n9507) );
  NAND2_X1 U10559 ( .A1(n9502), .A2(n9507), .ZN(n9243) );
  XNOR2_X1 U10560 ( .A(n9243), .B(n9508), .ZN(n9283) );
  INV_X1 U10561 ( .A(n9248), .ZN(n9249) );
  NAND2_X1 U10562 ( .A1(n9400), .A2(n9255), .ZN(n9386) );
  INV_X1 U10563 ( .A(n9260), .ZN(n9341) );
  NOR2_X1 U10564 ( .A1(n9340), .A2(n9341), .ZN(n9261) );
  NAND2_X1 U10565 ( .A1(n9313), .A2(n9265), .ZN(n9286) );
  NAND2_X1 U10566 ( .A1(n9286), .A2(n9285), .ZN(n9284) );
  NAND2_X1 U10567 ( .A1(n9284), .A2(n9266), .ZN(n9267) );
  XNOR2_X1 U10568 ( .A(n9267), .B(n9508), .ZN(n9274) );
  AOI21_X2 U10569 ( .B1(n9274), .B2(n9454), .A(n9273), .ZN(n9513) );
  AOI21_X1 U10570 ( .B1(n9511), .B2(n9297), .A(n9984), .ZN(n9276) );
  AND2_X2 U10571 ( .A1(n9276), .A2(n9275), .ZN(n9510) );
  NAND2_X1 U10572 ( .A1(n9510), .A2(n9277), .ZN(n9278) );
  OAI211_X1 U10573 ( .C1(n9279), .C2(n9460), .A(n9513), .B(n9278), .ZN(n9280)
         );
  NAND2_X1 U10574 ( .A1(n9280), .A2(n9463), .ZN(n9282) );
  AOI22_X1 U10575 ( .A1(n9511), .A2(n9365), .B1(n4246), .B2(
        P1_REG2_REG_29__SCAN_IN), .ZN(n9281) );
  OAI211_X1 U10576 ( .C1(n9493), .C2(n9283), .A(n9282), .B(n9281), .ZN(
        P1_U3355) );
  OAI211_X1 U10577 ( .C1(n9286), .C2(n9285), .A(n9284), .B(n9454), .ZN(n9291)
         );
  OAI22_X1 U10578 ( .A1(n9288), .A2(n9482), .B1(n9287), .B2(n9484), .ZN(n9289)
         );
  INV_X1 U10579 ( .A(n9289), .ZN(n9290) );
  OAI22_X1 U10580 ( .A1(n9294), .A2(n9460), .B1(n9293), .B2(n9463), .ZN(n9295)
         );
  AOI21_X1 U10581 ( .B1(n9514), .B2(n9365), .A(n9295), .ZN(n9300) );
  OR2_X1 U10582 ( .A1(n9296), .A2(n9306), .ZN(n9298) );
  AND2_X1 U10583 ( .A1(n9298), .A2(n9297), .ZN(n9515) );
  NAND2_X1 U10584 ( .A1(n9515), .A2(n9491), .ZN(n9299) );
  OAI211_X1 U10585 ( .C1(n9518), .C2(n9493), .A(n9300), .B(n9299), .ZN(n9301)
         );
  INV_X1 U10586 ( .A(n9301), .ZN(n9302) );
  OAI21_X1 U10587 ( .B1(n4246), .B2(n9517), .A(n9302), .ZN(P1_U3263) );
  XOR2_X1 U10588 ( .A(n9314), .B(n9303), .Z(n9524) );
  NAND2_X1 U10589 ( .A1(n9520), .A2(n9328), .ZN(n9304) );
  NAND2_X1 U10590 ( .A1(n9304), .A2(n9945), .ZN(n9305) );
  NOR2_X1 U10591 ( .A1(n9306), .A2(n9305), .ZN(n9519) );
  NAND2_X1 U10592 ( .A1(n9520), .A2(n9365), .ZN(n9309) );
  AOI22_X1 U10593 ( .A1(n9307), .A2(n9472), .B1(P1_REG2_REG_27__SCAN_IN), .B2(
        n4246), .ZN(n9308) );
  NAND2_X1 U10594 ( .A1(n9309), .A2(n9308), .ZN(n9310) );
  AOI21_X1 U10595 ( .B1(n9519), .B2(n9410), .A(n9310), .ZN(n9320) );
  OAI211_X1 U10596 ( .C1(n4327), .C2(n9314), .A(n9313), .B(n9454), .ZN(n9317)
         );
  NAND2_X1 U10597 ( .A1(n9315), .A2(n9451), .ZN(n9316) );
  NAND2_X1 U10598 ( .A1(n9523), .A2(n9463), .ZN(n9319) );
  OAI211_X1 U10599 ( .C1(n9524), .C2(n9493), .A(n9320), .B(n9319), .ZN(
        P1_U3264) );
  NAND2_X1 U10600 ( .A1(n9358), .A2(n9451), .ZN(n9323) );
  AOI211_X1 U10601 ( .C1(n9527), .C2(n9327), .A(n9984), .B(n9209), .ZN(n9526)
         );
  AOI22_X1 U10602 ( .A1(n9329), .A2(n9472), .B1(P1_REG2_REG_26__SCAN_IN), .B2(
        n4246), .ZN(n9330) );
  OAI21_X1 U10603 ( .B1(n9331), .B2(n9475), .A(n9330), .ZN(n9335) );
  XNOR2_X1 U10604 ( .A(n9333), .B(n9332), .ZN(n9530) );
  NOR2_X1 U10605 ( .A1(n9530), .A2(n9493), .ZN(n9334) );
  AOI211_X1 U10606 ( .C1(n9410), .C2(n9526), .A(n9335), .B(n9334), .ZN(n9336)
         );
  OAI21_X1 U10607 ( .B1(n4246), .B2(n9529), .A(n9336), .ZN(P1_U3265) );
  INV_X1 U10608 ( .A(n9337), .ZN(n9361) );
  NAND2_X1 U10609 ( .A1(n9361), .A2(n9360), .ZN(n9359) );
  NAND2_X1 U10610 ( .A1(n9359), .A2(n9338), .ZN(n9339) );
  XNOR2_X1 U10611 ( .A(n9339), .B(n9340), .ZN(n9535) );
  OAI21_X1 U10612 ( .B1(n9342), .B2(n9341), .A(n9340), .ZN(n9344) );
  NAND2_X1 U10613 ( .A1(n9374), .A2(n9451), .ZN(n9345) );
  INV_X1 U10614 ( .A(n9363), .ZN(n9348) );
  INV_X1 U10615 ( .A(n9327), .ZN(n9347) );
  AOI211_X1 U10616 ( .C1(n9533), .C2(n9348), .A(n9984), .B(n9347), .ZN(n9532)
         );
  NAND2_X1 U10617 ( .A1(n9532), .A2(n9410), .ZN(n9351) );
  AOI22_X1 U10618 ( .A1(n9349), .A2(n9472), .B1(P1_REG2_REG_25__SCAN_IN), .B2(
        n4246), .ZN(n9350) );
  OAI211_X1 U10619 ( .C1(n9352), .C2(n9475), .A(n9351), .B(n9350), .ZN(n9353)
         );
  AOI21_X1 U10620 ( .B1(n9531), .B2(n9463), .A(n9353), .ZN(n9354) );
  OAI21_X1 U10621 ( .B1(n9535), .B2(n9493), .A(n9354), .ZN(P1_U3266) );
  OAI21_X1 U10622 ( .B1(n9361), .B2(n9360), .A(n9359), .ZN(n9540) );
  INV_X1 U10623 ( .A(n9540), .ZN(n9371) );
  AND2_X1 U10624 ( .A1(n9377), .A2(n9366), .ZN(n9362) );
  OR2_X1 U10625 ( .A1(n9363), .A2(n9362), .ZN(n9536) );
  AOI22_X1 U10626 ( .A1(n9364), .A2(n9472), .B1(P1_REG2_REG_24__SCAN_IN), .B2(
        n4246), .ZN(n9368) );
  NAND2_X1 U10627 ( .A1(n9366), .A2(n9365), .ZN(n9367) );
  OAI211_X1 U10628 ( .C1(n9536), .C2(n9369), .A(n9368), .B(n9367), .ZN(n9370)
         );
  AOI21_X1 U10629 ( .B1(n9371), .B2(n9467), .A(n9370), .ZN(n9372) );
  OAI21_X1 U10630 ( .B1(n4246), .B2(n9539), .A(n9372), .ZN(P1_U3267) );
  XOR2_X1 U10631 ( .A(n9373), .B(n9382), .Z(n9375) );
  AOI222_X1 U10632 ( .A1(n9454), .A2(n9375), .B1(n9374), .B2(n9449), .C1(n9402), .C2(n9451), .ZN(n9544) );
  NAND2_X1 U10633 ( .A1(n9390), .A2(n9541), .ZN(n9376) );
  AND2_X1 U10634 ( .A1(n9377), .A2(n9376), .ZN(n9542) );
  INV_X1 U10635 ( .A(n9541), .ZN(n9380) );
  AOI22_X1 U10636 ( .A1(n9378), .A2(n9472), .B1(P1_REG2_REG_23__SCAN_IN), .B2(
        n4246), .ZN(n9379) );
  OAI21_X1 U10637 ( .B1(n9380), .B2(n9475), .A(n9379), .ZN(n9384) );
  XOR2_X1 U10638 ( .A(n9381), .B(n9382), .Z(n9545) );
  NOR2_X1 U10639 ( .A1(n9545), .A2(n9493), .ZN(n9383) );
  AOI211_X1 U10640 ( .C1(n9542), .C2(n9491), .A(n9384), .B(n9383), .ZN(n9385)
         );
  OAI21_X1 U10641 ( .B1(n4246), .B2(n9544), .A(n9385), .ZN(P1_U3268) );
  XNOR2_X1 U10642 ( .A(n9386), .B(n9396), .ZN(n9388) );
  AOI222_X1 U10643 ( .A1(n9454), .A2(n9388), .B1(n9387), .B2(n9449), .C1(n9419), .C2(n9451), .ZN(n9549) );
  OR2_X1 U10644 ( .A1(n9408), .A2(n9394), .ZN(n9389) );
  AND2_X1 U10645 ( .A1(n9390), .A2(n9389), .ZN(n9547) );
  INV_X1 U10646 ( .A(n9391), .ZN(n9392) );
  AOI22_X1 U10647 ( .A1(n9392), .A2(n9472), .B1(P1_REG2_REG_22__SCAN_IN), .B2(
        n4246), .ZN(n9393) );
  OAI21_X1 U10648 ( .B1(n9394), .B2(n9475), .A(n9393), .ZN(n9398) );
  XOR2_X1 U10649 ( .A(n9396), .B(n9395), .Z(n9550) );
  NOR2_X1 U10650 ( .A1(n9550), .A2(n9493), .ZN(n9397) );
  AOI211_X1 U10651 ( .C1(n9547), .C2(n9491), .A(n9398), .B(n9397), .ZN(n9399)
         );
  OAI21_X1 U10652 ( .B1(n4246), .B2(n9549), .A(n9399), .ZN(P1_U3269) );
  OAI21_X1 U10653 ( .B1(n9401), .B2(n9254), .A(n9400), .ZN(n9403) );
  AOI222_X1 U10654 ( .A1(n9454), .A2(n9403), .B1(n9402), .B2(n9449), .C1(n9440), .C2(n9451), .ZN(n9554) );
  OAI21_X1 U10655 ( .B1(n9406), .B2(n9405), .A(n9404), .ZN(n9555) );
  INV_X1 U10656 ( .A(n9555), .ZN(n9416) );
  OAI21_X1 U10657 ( .B1(n9407), .B2(n9414), .A(n9945), .ZN(n9409) );
  NOR2_X1 U10658 ( .A1(n9409), .A2(n9408), .ZN(n9551) );
  NAND2_X1 U10659 ( .A1(n9551), .A2(n9410), .ZN(n9413) );
  AOI22_X1 U10660 ( .A1(n9411), .A2(n9472), .B1(P1_REG2_REG_21__SCAN_IN), .B2(
        n4246), .ZN(n9412) );
  OAI211_X1 U10661 ( .C1(n9414), .C2(n9475), .A(n9413), .B(n9412), .ZN(n9415)
         );
  AOI21_X1 U10662 ( .B1(n9416), .B2(n9467), .A(n9415), .ZN(n9417) );
  OAI21_X1 U10663 ( .B1(n4246), .B2(n9554), .A(n9417), .ZN(P1_U3270) );
  XOR2_X1 U10664 ( .A(n9418), .B(n9427), .Z(n9420) );
  AOI222_X1 U10665 ( .A1(n9454), .A2(n9420), .B1(n9419), .B2(n9449), .C1(n9450), .C2(n9451), .ZN(n9559) );
  INV_X1 U10666 ( .A(n9421), .ZN(n9434) );
  AND2_X1 U10667 ( .A1(n9434), .A2(n9556), .ZN(n9422) );
  NOR2_X1 U10668 ( .A1(n9407), .A2(n9422), .ZN(n9557) );
  INV_X1 U10669 ( .A(n9423), .ZN(n9424) );
  AOI22_X1 U10670 ( .A1(n9424), .A2(n9472), .B1(n4246), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9425) );
  OAI21_X1 U10671 ( .B1(n9426), .B2(n9475), .A(n9425), .ZN(n9430) );
  XNOR2_X1 U10672 ( .A(n9428), .B(n9427), .ZN(n9560) );
  NOR2_X1 U10673 ( .A1(n9560), .A2(n9493), .ZN(n9429) );
  AOI211_X1 U10674 ( .C1(n9557), .C2(n9491), .A(n9430), .B(n9429), .ZN(n9431)
         );
  OAI21_X1 U10675 ( .B1(n4246), .B2(n9559), .A(n9431), .ZN(P1_U3271) );
  XOR2_X1 U10676 ( .A(n9432), .B(n9439), .Z(n9565) );
  NAND2_X1 U10677 ( .A1(n9456), .A2(n9561), .ZN(n9433) );
  AND2_X1 U10678 ( .A1(n9434), .A2(n9433), .ZN(n9562) );
  OAI22_X1 U10679 ( .A1(n9435), .A2(n9475), .B1(n9463), .B2(n4526), .ZN(n9436)
         );
  AOI21_X1 U10680 ( .B1(n9562), .B2(n9491), .A(n9436), .ZN(n9446) );
  OAI21_X1 U10681 ( .B1(n9439), .B2(n9438), .A(n9437), .ZN(n9442) );
  AOI222_X1 U10682 ( .A1(n9454), .A2(n9442), .B1(n9441), .B2(n9451), .C1(n9440), .C2(n9449), .ZN(n9564) );
  OAI21_X1 U10683 ( .B1(n9443), .B2(n9460), .A(n9564), .ZN(n9444) );
  NAND2_X1 U10684 ( .A1(n9444), .A2(n9463), .ZN(n9445) );
  OAI211_X1 U10685 ( .C1(n9565), .C2(n9493), .A(n9446), .B(n9445), .ZN(
        P1_U3272) );
  OAI21_X1 U10686 ( .B1(n9448), .B2(n9249), .A(n9447), .ZN(n9453) );
  AOI222_X1 U10687 ( .A1(n9454), .A2(n9453), .B1(n9452), .B2(n9451), .C1(n9450), .C2(n9449), .ZN(n9571) );
  INV_X1 U10688 ( .A(n9455), .ZN(n9458) );
  INV_X1 U10689 ( .A(n9456), .ZN(n9457) );
  AOI21_X1 U10690 ( .B1(n9568), .B2(n9458), .A(n9457), .ZN(n9569) );
  NOR2_X1 U10691 ( .A1(n9459), .A2(n9475), .ZN(n9465) );
  OAI22_X1 U10692 ( .A1(n9463), .A2(n9462), .B1(n9461), .B2(n9460), .ZN(n9464)
         );
  AOI211_X1 U10693 ( .C1(n9569), .C2(n9491), .A(n9465), .B(n9464), .ZN(n9469)
         );
  NAND2_X1 U10694 ( .A1(n9466), .A2(n9249), .ZN(n9566) );
  NAND3_X1 U10695 ( .A1(n9567), .A2(n9566), .A3(n9467), .ZN(n9468) );
  OAI211_X1 U10696 ( .C1(n9571), .C2(n4246), .A(n9469), .B(n9468), .ZN(
        P1_U3273) );
  XOR2_X1 U10697 ( .A(n4356), .B(n9478), .Z(n9577) );
  INV_X1 U10698 ( .A(n9208), .ZN(n9471) );
  AOI21_X1 U10699 ( .B1(n9573), .B2(n9471), .A(n9455), .ZN(n9574) );
  AOI22_X1 U10700 ( .A1(n4246), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9473), .B2(
        n9472), .ZN(n9474) );
  OAI21_X1 U10701 ( .B1(n9476), .B2(n9475), .A(n9474), .ZN(n9490) );
  INV_X1 U10702 ( .A(n9477), .ZN(n9481) );
  INV_X1 U10703 ( .A(n9478), .ZN(n9480) );
  AOI21_X1 U10704 ( .B1(n9481), .B2(n9480), .A(n9479), .ZN(n9488) );
  OAI22_X1 U10705 ( .A1(n9485), .A2(n9484), .B1(n9483), .B2(n9482), .ZN(n9486)
         );
  AOI21_X1 U10706 ( .B1(n9488), .B2(n9487), .A(n9486), .ZN(n9576) );
  NOR2_X1 U10707 ( .A1(n9576), .A2(n4246), .ZN(n9489) );
  AOI211_X1 U10708 ( .C1(n9574), .C2(n9491), .A(n9490), .B(n9489), .ZN(n9492)
         );
  OAI21_X1 U10709 ( .B1(n9493), .B2(n9577), .A(n9492), .ZN(P1_U3274) );
  NAND2_X1 U10710 ( .A1(n9494), .A2(n9945), .ZN(n9495) );
  OAI211_X1 U10711 ( .C1(n9982), .C2(n9496), .A(n9495), .B(n9499), .ZN(n9614)
         );
  MUX2_X1 U10712 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n9614), .S(n10003), .Z(
        P1_U3554) );
  NAND3_X1 U10713 ( .A1(n9498), .A2(n9945), .A3(n9497), .ZN(n9500) );
  OAI211_X1 U10714 ( .C1(n9501), .C2(n9982), .A(n9500), .B(n9499), .ZN(n9615)
         );
  MUX2_X1 U10715 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n9615), .S(n10003), .Z(
        P1_U3553) );
  NAND4_X1 U10716 ( .A1(n9502), .A2(n9508), .A3(n9979), .A4(n9507), .ZN(n9506)
         );
  INV_X1 U10717 ( .A(n9508), .ZN(n9503) );
  NAND3_X1 U10718 ( .A1(n9504), .A2(n9503), .A3(n9979), .ZN(n9505) );
  NOR3_X1 U10719 ( .A1(n9508), .A2(n9611), .A3(n9507), .ZN(n9509) );
  MUX2_X1 U10720 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n9616), .S(n10003), .Z(
        P1_U3552) );
  AOI22_X1 U10721 ( .A1(n9515), .A2(n9945), .B1(n9607), .B2(n9514), .ZN(n9516)
         );
  OAI211_X1 U10722 ( .C1(n9518), .C2(n9611), .A(n9517), .B(n9516), .ZN(n9617)
         );
  MUX2_X1 U10723 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n9617), .S(n10003), .Z(
        P1_U3551) );
  MUX2_X1 U10724 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n9618), .S(n10003), .Z(
        P1_U3550) );
  AOI21_X1 U10725 ( .B1(n9607), .B2(n9527), .A(n9526), .ZN(n9528) );
  OAI211_X1 U10726 ( .C1(n9611), .C2(n9530), .A(n9529), .B(n9528), .ZN(n9619)
         );
  MUX2_X1 U10727 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n9619), .S(n10003), .Z(
        P1_U3549) );
  AOI211_X1 U10728 ( .C1(n9607), .C2(n9533), .A(n9532), .B(n9531), .ZN(n9534)
         );
  OAI21_X1 U10729 ( .B1(n9611), .B2(n9535), .A(n9534), .ZN(n9620) );
  MUX2_X1 U10730 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n9620), .S(n10003), .Z(
        P1_U3548) );
  OAI22_X1 U10731 ( .A1(n9536), .A2(n9984), .B1(n4757), .B2(n9982), .ZN(n9537)
         );
  INV_X1 U10732 ( .A(n9537), .ZN(n9538) );
  OAI211_X1 U10733 ( .C1(n9540), .C2(n9611), .A(n9539), .B(n9538), .ZN(n9621)
         );
  MUX2_X1 U10734 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n9621), .S(n10003), .Z(
        P1_U3547) );
  AOI22_X1 U10735 ( .A1(n9542), .A2(n9945), .B1(n9607), .B2(n9541), .ZN(n9543)
         );
  OAI211_X1 U10736 ( .C1(n9545), .C2(n9611), .A(n9544), .B(n9543), .ZN(n9622)
         );
  MUX2_X1 U10737 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n9622), .S(n10003), .Z(
        P1_U3546) );
  AOI22_X1 U10738 ( .A1(n9547), .A2(n9945), .B1(n9607), .B2(n9546), .ZN(n9548)
         );
  OAI211_X1 U10739 ( .C1(n9550), .C2(n9611), .A(n9549), .B(n9548), .ZN(n9623)
         );
  MUX2_X1 U10740 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n9623), .S(n10003), .Z(
        P1_U3545) );
  AOI21_X1 U10741 ( .B1(n9607), .B2(n9552), .A(n9551), .ZN(n9553) );
  OAI211_X1 U10742 ( .C1(n9555), .C2(n9611), .A(n9554), .B(n9553), .ZN(n9624)
         );
  MUX2_X1 U10743 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n9624), .S(n10003), .Z(
        P1_U3544) );
  AOI22_X1 U10744 ( .A1(n9557), .A2(n9945), .B1(n9607), .B2(n9556), .ZN(n9558)
         );
  OAI211_X1 U10745 ( .C1(n9611), .C2(n9560), .A(n9559), .B(n9558), .ZN(n9625)
         );
  MUX2_X1 U10746 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n9625), .S(n10003), .Z(
        P1_U3543) );
  AOI22_X1 U10747 ( .A1(n9562), .A2(n9945), .B1(n9607), .B2(n9561), .ZN(n9563)
         );
  OAI211_X1 U10748 ( .C1(n9565), .C2(n9611), .A(n9564), .B(n9563), .ZN(n9626)
         );
  MUX2_X1 U10749 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n9626), .S(n10003), .Z(
        P1_U3542) );
  NAND3_X1 U10750 ( .A1(n9567), .A2(n9979), .A3(n9566), .ZN(n9572) );
  AOI22_X1 U10751 ( .A1(n9569), .A2(n9945), .B1(n9607), .B2(n9568), .ZN(n9570)
         );
  NAND3_X1 U10752 ( .A1(n9572), .A2(n9571), .A3(n9570), .ZN(n9627) );
  MUX2_X1 U10753 ( .A(n9627), .B(P1_REG1_REG_18__SCAN_IN), .S(n10000), .Z(
        P1_U3541) );
  AOI22_X1 U10754 ( .A1(n9574), .A2(n9945), .B1(n9607), .B2(n9573), .ZN(n9575)
         );
  OAI211_X1 U10755 ( .C1(n9577), .C2(n9611), .A(n9576), .B(n9575), .ZN(n9628)
         );
  MUX2_X1 U10756 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n9628), .S(n10003), .Z(
        P1_U3540) );
  AOI211_X1 U10757 ( .C1(n9607), .C2(n9580), .A(n9579), .B(n9578), .ZN(n9581)
         );
  OAI21_X1 U10758 ( .B1(n9611), .B2(n9582), .A(n9581), .ZN(n9629) );
  MUX2_X1 U10759 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9629), .S(n10003), .Z(
        P1_U3539) );
  AOI22_X1 U10760 ( .A1(n9584), .A2(n9945), .B1(n9607), .B2(n9583), .ZN(n9585)
         );
  OAI211_X1 U10761 ( .C1(n9587), .C2(n9611), .A(n9586), .B(n9585), .ZN(n9630)
         );
  MUX2_X1 U10762 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n9630), .S(n10003), .Z(
        P1_U3538) );
  AOI211_X1 U10763 ( .C1(n9607), .C2(n9590), .A(n9589), .B(n9588), .ZN(n9591)
         );
  OAI21_X1 U10764 ( .B1(n9611), .B2(n9592), .A(n9591), .ZN(n9772) );
  MUX2_X1 U10765 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n9772), .S(n10003), .Z(
        P1_U3537) );
  INV_X1 U10766 ( .A(n9593), .ZN(n9598) );
  AOI22_X1 U10767 ( .A1(n9595), .A2(n9945), .B1(n9607), .B2(n9594), .ZN(n9596)
         );
  OAI211_X1 U10768 ( .C1(n9602), .C2(n9598), .A(n9597), .B(n9596), .ZN(n9773)
         );
  MUX2_X1 U10769 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n9773), .S(n10003), .Z(
        P1_U3536) );
  NAND2_X1 U10770 ( .A1(n9599), .A2(n9607), .ZN(n9601) );
  OAI211_X1 U10771 ( .C1(n9603), .C2(n9602), .A(n9601), .B(n9600), .ZN(n9605)
         );
  MUX2_X1 U10772 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n9774), .S(n10003), .Z(
        P1_U3535) );
  AOI22_X1 U10773 ( .A1(n9608), .A2(n9945), .B1(n9607), .B2(n9606), .ZN(n9609)
         );
  OAI211_X1 U10774 ( .C1(n9612), .C2(n9611), .A(n9610), .B(n9609), .ZN(n9775)
         );
  MUX2_X1 U10775 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n9775), .S(n10003), .Z(
        P1_U3534) );
  MUX2_X1 U10776 ( .A(P1_REG1_REG_0__SCAN_IN), .B(n9613), .S(n10003), .Z(
        P1_U3523) );
  MUX2_X1 U10777 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n9614), .S(n9991), .Z(
        P1_U3522) );
  MUX2_X1 U10778 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n9615), .S(n9991), .Z(
        P1_U3521) );
  MUX2_X1 U10779 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n9616), .S(n9991), .Z(
        P1_U3520) );
  MUX2_X1 U10780 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n9617), .S(n9991), .Z(
        P1_U3519) );
  MUX2_X1 U10781 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n9619), .S(n9991), .Z(
        P1_U3517) );
  MUX2_X1 U10782 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n9620), .S(n9991), .Z(
        P1_U3516) );
  MUX2_X1 U10783 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n9621), .S(n9991), .Z(
        P1_U3515) );
  MUX2_X1 U10784 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n9622), .S(n9991), .Z(
        P1_U3514) );
  MUX2_X1 U10785 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n9623), .S(n9991), .Z(
        P1_U3513) );
  MUX2_X1 U10786 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n9624), .S(n9991), .Z(
        P1_U3512) );
  MUX2_X1 U10787 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n9625), .S(n9991), .Z(
        P1_U3511) );
  MUX2_X1 U10788 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n9626), .S(n9991), .Z(
        P1_U3510) );
  MUX2_X1 U10789 ( .A(n9627), .B(P1_REG0_REG_18__SCAN_IN), .S(n9990), .Z(
        P1_U3508) );
  MUX2_X1 U10790 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n9628), .S(n9991), .Z(
        P1_U3505) );
  MUX2_X1 U10791 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n9629), .S(n9991), .Z(
        P1_U3502) );
  MUX2_X1 U10792 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n9630), .S(n9991), .Z(n9771) );
  INV_X1 U10793 ( .A(P1_D_REG_11__SCAN_IN), .ZN(n9940) );
  NOR4_X1 U10794 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(P1_REG0_REG_7__SCAN_IN), 
        .A3(P2_ADDR_REG_17__SCAN_IN), .A4(n9940), .ZN(n9631) );
  INV_X1 U10795 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n9805) );
  NAND4_X1 U10796 ( .A1(P1_REG1_REG_6__SCAN_IN), .A2(P1_ADDR_REG_1__SCAN_IN), 
        .A3(n9631), .A4(n9805), .ZN(n9650) );
  NOR4_X1 U10797 ( .A1(n9633), .A2(n9632), .A3(P1_DATAO_REG_7__SCAN_IN), .A4(
        P2_REG3_REG_4__SCAN_IN), .ZN(n9639) );
  NAND4_X1 U10798 ( .A1(P2_REG0_REG_14__SCAN_IN), .A2(n9712), .A3(n9717), .A4(
        n9674), .ZN(n9636) );
  NAND4_X1 U10799 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(P1_REG2_REG_28__SCAN_IN), .A3(n9634), .A4(n9676), .ZN(n9635) );
  NOR4_X1 U10800 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(n9636), .A3(n9635), .A4(
        P2_REG2_REG_14__SCAN_IN), .ZN(n9638) );
  NAND4_X1 U10801 ( .A1(n9639), .A2(n9638), .A3(n9733), .A4(n9637), .ZN(n9649)
         );
  NOR4_X1 U10802 ( .A1(n9680), .A2(n9640), .A3(P1_REG0_REG_25__SCAN_IN), .A4(
        P1_REG0_REG_13__SCAN_IN), .ZN(n9645) );
  NOR4_X1 U10803 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .A3(
        P1_IR_REG_25__SCAN_IN), .A4(P1_REG3_REG_26__SCAN_IN), .ZN(n9644) );
  NAND4_X1 U10804 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(P2_IR_REG_17__SCAN_IN), 
        .A3(P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_6__SCAN_IN), .ZN(n9642) );
  NAND4_X1 U10805 ( .A1(P1_REG0_REG_2__SCAN_IN), .A2(P2_D_REG_28__SCAN_IN), 
        .A3(P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n9641) );
  NOR2_X1 U10806 ( .A1(n9642), .A2(n9641), .ZN(n9643) );
  NAND3_X1 U10807 ( .A1(n9645), .A2(n9644), .A3(n9643), .ZN(n9648) );
  NAND4_X1 U10808 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), 
        .A3(P2_REG0_REG_24__SCAN_IN), .A4(n9646), .ZN(n9647) );
  NOR4_X1 U10809 ( .A1(n9650), .A2(n9649), .A3(n9648), .A4(n9647), .ZN(n9657)
         );
  NOR4_X1 U10810 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_REG0_REG_10__SCAN_IN), 
        .A3(n9750), .A4(n5567), .ZN(n9656) );
  NAND3_X1 U10811 ( .A1(P2_REG3_REG_23__SCAN_IN), .A2(P2_WR_REG_SCAN_IN), .A3(
        n9665), .ZN(n9653) );
  INV_X1 U10812 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n9725) );
  NAND4_X1 U10813 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(P1_REG3_REG_6__SCAN_IN), 
        .A3(P2_REG2_REG_9__SCAN_IN), .A4(n9725), .ZN(n9652) );
  NAND4_X1 U10814 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .A3(P2_REG1_REG_23__SCAN_IN), .A4(P1_DATAO_REG_30__SCAN_IN), .ZN(n9651) );
  NOR4_X1 U10815 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n9653), .A3(n9652), .A4(n9651), .ZN(n9655) );
  NOR4_X1 U10816 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P2_DATAO_REG_21__SCAN_IN), 
        .A3(P2_DATAO_REG_28__SCAN_IN), .A4(n10104), .ZN(n9654) );
  NAND4_X1 U10817 ( .A1(n9657), .A2(n9656), .A3(n9655), .A4(n9654), .ZN(n9658)
         );
  AND2_X1 U10818 ( .A1(n9658), .A2(n9740), .ZN(n9769) );
  INV_X1 U10819 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n9660) );
  AOI22_X1 U10820 ( .A1(n10106), .A2(keyinput18), .B1(keyinput17), .B2(n9660), 
        .ZN(n9659) );
  OAI221_X1 U10821 ( .B1(n10106), .B2(keyinput18), .C1(n9660), .C2(keyinput17), 
        .A(n9659), .ZN(n9672) );
  AOI22_X1 U10822 ( .A1(n9663), .A2(keyinput9), .B1(n9662), .B2(keyinput50), 
        .ZN(n9661) );
  OAI221_X1 U10823 ( .B1(n9663), .B2(keyinput9), .C1(n9662), .C2(keyinput50), 
        .A(n9661), .ZN(n9671) );
  AOI22_X1 U10824 ( .A1(n9666), .A2(keyinput54), .B1(keyinput27), .B2(n9665), 
        .ZN(n9664) );
  OAI221_X1 U10825 ( .B1(n9666), .B2(keyinput54), .C1(n9665), .C2(keyinput27), 
        .A(n9664), .ZN(n9670) );
  INV_X1 U10826 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n9668) );
  INV_X1 U10827 ( .A(P1_D_REG_8__SCAN_IN), .ZN(n9941) );
  AOI22_X1 U10828 ( .A1(n9668), .A2(keyinput63), .B1(n9941), .B2(keyinput56), 
        .ZN(n9667) );
  OAI221_X1 U10829 ( .B1(n9668), .B2(keyinput63), .C1(n9941), .C2(keyinput56), 
        .A(n9667), .ZN(n9669) );
  NOR4_X1 U10830 ( .A1(n9672), .A2(n9671), .A3(n9670), .A4(n9669), .ZN(n9768)
         );
  AOI22_X1 U10831 ( .A1(n9674), .A2(keyinput3), .B1(n5567), .B2(keyinput8), 
        .ZN(n9673) );
  OAI221_X1 U10832 ( .B1(n9674), .B2(keyinput3), .C1(n5567), .C2(keyinput8), 
        .A(n9673), .ZN(n9678) );
  AOI22_X1 U10833 ( .A1(n9676), .A2(keyinput12), .B1(n9293), .B2(keyinput34), 
        .ZN(n9675) );
  OAI221_X1 U10834 ( .B1(n9676), .B2(keyinput12), .C1(n9293), .C2(keyinput34), 
        .A(n9675), .ZN(n9677) );
  NOR2_X1 U10835 ( .A1(n9678), .A2(n9677), .ZN(n9708) );
  AOI22_X1 U10836 ( .A1(n9640), .A2(keyinput1), .B1(n9680), .B2(keyinput16), 
        .ZN(n9679) );
  OAI221_X1 U10837 ( .B1(n9640), .B2(keyinput1), .C1(n9680), .C2(keyinput16), 
        .A(n9679), .ZN(n9684) );
  AOI22_X1 U10838 ( .A1(n9940), .A2(keyinput30), .B1(keyinput32), .B2(n9682), 
        .ZN(n9681) );
  OAI221_X1 U10839 ( .B1(n9940), .B2(keyinput30), .C1(n9682), .C2(keyinput32), 
        .A(n9681), .ZN(n9683) );
  NOR2_X1 U10840 ( .A1(n9684), .A2(n9683), .ZN(n9707) );
  XNOR2_X1 U10841 ( .A(SI_9_), .B(keyinput5), .ZN(n9688) );
  XNOR2_X1 U10842 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(keyinput2), .ZN(n9687) );
  XNOR2_X1 U10843 ( .A(P1_IR_REG_25__SCAN_IN), .B(keyinput37), .ZN(n9686) );
  XNOR2_X1 U10844 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(keyinput25), .ZN(n9685)
         );
  NAND4_X1 U10845 ( .A1(n9688), .A2(n9687), .A3(n9686), .A4(n9685), .ZN(n9694)
         );
  XNOR2_X1 U10846 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput22), .ZN(n9692) );
  XNOR2_X1 U10847 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(keyinput62), .ZN(n9691) );
  XNOR2_X1 U10848 ( .A(P1_REG3_REG_6__SCAN_IN), .B(keyinput29), .ZN(n9690) );
  XNOR2_X1 U10849 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(keyinput60), .ZN(n9689)
         );
  NAND4_X1 U10850 ( .A1(n9692), .A2(n9691), .A3(n9690), .A4(n9689), .ZN(n9693)
         );
  NOR2_X1 U10851 ( .A1(n9694), .A2(n9693), .ZN(n9706) );
  XNOR2_X1 U10852 ( .A(P1_REG3_REG_26__SCAN_IN), .B(keyinput45), .ZN(n9698) );
  XNOR2_X1 U10853 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(keyinput59), .ZN(n9697) );
  XNOR2_X1 U10854 ( .A(keyinput42), .B(P2_REG2_REG_9__SCAN_IN), .ZN(n9696) );
  XNOR2_X1 U10855 ( .A(keyinput26), .B(P2_REG2_REG_14__SCAN_IN), .ZN(n9695) );
  NAND4_X1 U10856 ( .A1(n9698), .A2(n9697), .A3(n9696), .A4(n9695), .ZN(n9704)
         );
  XNOR2_X1 U10857 ( .A(keyinput36), .B(P2_D_REG_28__SCAN_IN), .ZN(n9702) );
  XNOR2_X1 U10858 ( .A(keyinput47), .B(P1_REG0_REG_2__SCAN_IN), .ZN(n9701) );
  XNOR2_X1 U10859 ( .A(keyinput24), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n9700) );
  INV_X1 U10860 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n9980) );
  XNOR2_X1 U10861 ( .A(keyinput58), .B(P1_REG0_REG_7__SCAN_IN), .ZN(n9699) );
  NAND4_X1 U10862 ( .A1(n9702), .A2(n9701), .A3(n9700), .A4(n9699), .ZN(n9703)
         );
  NOR2_X1 U10863 ( .A1(n9704), .A2(n9703), .ZN(n9705) );
  AND4_X1 U10864 ( .A1(n9708), .A2(n9707), .A3(n9706), .A4(n9705), .ZN(n9715)
         );
  INV_X1 U10865 ( .A(P1_D_REG_16__SCAN_IN), .ZN(n9939) );
  INV_X1 U10866 ( .A(P1_D_REG_20__SCAN_IN), .ZN(n9938) );
  OAI22_X1 U10867 ( .A1(n9939), .A2(keyinput53), .B1(n9938), .B2(keyinput21), 
        .ZN(n9709) );
  AOI221_X1 U10868 ( .B1(n9939), .B2(keyinput53), .C1(keyinput21), .C2(n9938), 
        .A(n9709), .ZN(n9714) );
  OAI22_X1 U10869 ( .A1(n9712), .A2(keyinput43), .B1(n9711), .B2(keyinput14), 
        .ZN(n9710) );
  AOI221_X1 U10870 ( .B1(n9712), .B2(keyinput43), .C1(keyinput14), .C2(n9711), 
        .A(n9710), .ZN(n9713) );
  NAND3_X1 U10871 ( .A1(n9715), .A2(n9714), .A3(n9713), .ZN(n9766) );
  INV_X1 U10872 ( .A(P1_D_REG_29__SCAN_IN), .ZN(n9936) );
  OAI22_X1 U10873 ( .A1(n9936), .A2(keyinput61), .B1(n9717), .B2(keyinput41), 
        .ZN(n9716) );
  AOI221_X1 U10874 ( .B1(n9936), .B2(keyinput61), .C1(keyinput41), .C2(n9717), 
        .A(n9716), .ZN(n9718) );
  INV_X1 U10875 ( .A(n9718), .ZN(n9765) );
  INV_X1 U10876 ( .A(P2_WR_REG_SCAN_IN), .ZN(n9834) );
  AOI22_X1 U10877 ( .A1(n9834), .A2(keyinput40), .B1(n9462), .B2(keyinput55), 
        .ZN(n9719) );
  OAI221_X1 U10878 ( .B1(n9834), .B2(keyinput40), .C1(n9462), .C2(keyinput55), 
        .A(n9719), .ZN(n9728) );
  AOI22_X1 U10879 ( .A1(n9722), .A2(keyinput10), .B1(n9721), .B2(keyinput6), 
        .ZN(n9720) );
  OAI221_X1 U10880 ( .B1(n9722), .B2(keyinput10), .C1(n9721), .C2(keyinput6), 
        .A(n9720), .ZN(n9727) );
  AOI22_X1 U10881 ( .A1(n9725), .A2(keyinput15), .B1(n9724), .B2(keyinput31), 
        .ZN(n9723) );
  OAI221_X1 U10882 ( .B1(n9725), .B2(keyinput15), .C1(n9724), .C2(keyinput31), 
        .A(n9723), .ZN(n9726) );
  NOR3_X1 U10883 ( .A1(n9728), .A2(n9727), .A3(n9726), .ZN(n9763) );
  INV_X1 U10884 ( .A(P1_D_REG_27__SCAN_IN), .ZN(n9937) );
  AOI22_X1 U10885 ( .A1(n9937), .A2(keyinput20), .B1(keyinput57), .B2(n9730), 
        .ZN(n9729) );
  OAI221_X1 U10886 ( .B1(n9937), .B2(keyinput20), .C1(n9730), .C2(keyinput57), 
        .A(n9729), .ZN(n9735) );
  AOI22_X1 U10887 ( .A1(n9733), .A2(keyinput35), .B1(keyinput49), .B2(n9732), 
        .ZN(n9731) );
  OAI221_X1 U10888 ( .B1(n9733), .B2(keyinput35), .C1(n9732), .C2(keyinput49), 
        .A(n9731), .ZN(n9734) );
  NOR2_X1 U10889 ( .A1(n9735), .A2(n9734), .ZN(n9748) );
  XNOR2_X1 U10890 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(keyinput28), .ZN(n9739) );
  XNOR2_X1 U10891 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput11), .ZN(n9738) );
  XNOR2_X1 U10892 ( .A(P1_REG0_REG_10__SCAN_IN), .B(keyinput33), .ZN(n9737) );
  XNOR2_X1 U10893 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput48), .ZN(n9736) );
  NAND4_X1 U10894 ( .A1(n9739), .A2(n9738), .A3(n9737), .A4(n9736), .ZN(n9746)
         );
  XNOR2_X1 U10895 ( .A(P2_IR_REG_17__SCAN_IN), .B(keyinput52), .ZN(n9744) );
  XNOR2_X1 U10896 ( .A(SI_22_), .B(keyinput0), .ZN(n9743) );
  XNOR2_X1 U10897 ( .A(P2_IR_REG_21__SCAN_IN), .B(keyinput23), .ZN(n9742) );
  NAND2_X1 U10898 ( .A1(n9740), .A2(keyinput44), .ZN(n9741) );
  NAND4_X1 U10899 ( .A1(n9744), .A2(n9743), .A3(n9742), .A4(n9741), .ZN(n9745)
         );
  NOR2_X1 U10900 ( .A1(n9746), .A2(n9745), .ZN(n9747) );
  AND2_X1 U10901 ( .A1(n9748), .A2(n9747), .ZN(n9762) );
  INV_X1 U10902 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10216) );
  AOI22_X1 U10903 ( .A1(n9750), .A2(keyinput13), .B1(keyinput51), .B2(n10216), 
        .ZN(n9749) );
  OAI221_X1 U10904 ( .B1(n9750), .B2(keyinput13), .C1(n10216), .C2(keyinput51), 
        .A(n9749), .ZN(n9753) );
  INV_X1 U10905 ( .A(P2_D_REG_6__SCAN_IN), .ZN(n10107) );
  AOI22_X1 U10906 ( .A1(n10105), .A2(keyinput19), .B1(keyinput7), .B2(n10107), 
        .ZN(n9751) );
  OAI221_X1 U10907 ( .B1(n10105), .B2(keyinput19), .C1(n10107), .C2(keyinput7), 
        .A(n9751), .ZN(n9752) );
  NOR2_X1 U10908 ( .A1(n9753), .A2(n9752), .ZN(n9761) );
  AOI22_X1 U10909 ( .A1(n9755), .A2(keyinput38), .B1(keyinput4), .B2(n10104), 
        .ZN(n9754) );
  OAI221_X1 U10910 ( .B1(n9755), .B2(keyinput38), .C1(n10104), .C2(keyinput4), 
        .A(n9754), .ZN(n9759) );
  AOI22_X1 U10911 ( .A1(n9757), .A2(keyinput46), .B1(keyinput39), .B2(n5213), 
        .ZN(n9756) );
  OAI221_X1 U10912 ( .B1(n9757), .B2(keyinput46), .C1(n5213), .C2(keyinput39), 
        .A(n9756), .ZN(n9758) );
  NOR2_X1 U10913 ( .A1(n9759), .A2(n9758), .ZN(n9760) );
  NAND4_X1 U10914 ( .A1(n9763), .A2(n9762), .A3(n9761), .A4(n9760), .ZN(n9764)
         );
  NOR3_X1 U10915 ( .A1(n9766), .A2(n9765), .A3(n9764), .ZN(n9767) );
  OAI211_X1 U10916 ( .C1(n9769), .C2(keyinput44), .A(n9768), .B(n9767), .ZN(
        n9770) );
  XNOR2_X1 U10917 ( .A(n9771), .B(n9770), .ZN(P1_U3499) );
  MUX2_X1 U10918 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n9772), .S(n9991), .Z(
        P1_U3496) );
  MUX2_X1 U10919 ( .A(P1_REG0_REG_13__SCAN_IN), .B(n9773), .S(n9991), .Z(
        P1_U3493) );
  MUX2_X1 U10920 ( .A(n9774), .B(P1_REG0_REG_12__SCAN_IN), .S(n9990), .Z(
        P1_U3490) );
  MUX2_X1 U10921 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n9775), .S(n9991), .Z(
        P1_U3487) );
  MUX2_X1 U10922 ( .A(P1_D_REG_0__SCAN_IN), .B(n9778), .S(n9942), .Z(P1_U3440)
         );
  NOR4_X1 U10923 ( .A1(n9780), .A2(P1_IR_REG_30__SCAN_IN), .A3(n9779), .A4(
        P1_U3084), .ZN(n9781) );
  AOI21_X1 U10924 ( .B1(n9793), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n9781), .ZN(
        n9782) );
  OAI21_X1 U10925 ( .B1(n9783), .B2(n9798), .A(n9782), .ZN(P1_U3322) );
  OAI222_X1 U10926 ( .A1(n9787), .A2(n9786), .B1(P1_U3084), .B2(n9785), .C1(
        n9798), .C2(n9784), .ZN(P1_U3324) );
  INV_X1 U10927 ( .A(n9788), .ZN(n9791) );
  AOI21_X1 U10928 ( .B1(n9793), .B2(P2_DATAO_REG_28__SCAN_IN), .A(n9789), .ZN(
        n9790) );
  OAI21_X1 U10929 ( .B1(n9791), .B2(n9798), .A(n9790), .ZN(P1_U3325) );
  AOI21_X1 U10930 ( .B1(n9793), .B2(P2_DATAO_REG_27__SCAN_IN), .A(n9792), .ZN(
        n9794) );
  OAI21_X1 U10931 ( .B1(n9795), .B2(n9798), .A(n9794), .ZN(P1_U3326) );
  OAI222_X1 U10932 ( .A1(P1_U3084), .A2(n9799), .B1(n9798), .B2(n9797), .C1(
        n9796), .C2(n9787), .ZN(P1_U3327) );
  INV_X1 U10933 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n10212) );
  NOR2_X1 U10934 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n9800) );
  AOI21_X1 U10935 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n9800), .ZN(n10184) );
  NOR2_X1 U10936 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n9801) );
  AOI21_X1 U10937 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n9801), .ZN(n10187) );
  NOR2_X1 U10938 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n9802) );
  AOI21_X1 U10939 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n9802), .ZN(n10190) );
  NOR2_X1 U10940 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n9803) );
  AOI21_X1 U10941 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n9803), .ZN(n10193) );
  NOR2_X1 U10942 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n9804) );
  AOI21_X1 U10943 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n9804), .ZN(n10196) );
  NOR2_X1 U10944 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(P1_ADDR_REG_4__SCAN_IN), 
        .ZN(n9813) );
  AOI22_X1 U10945 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n9806), .B1(
        P1_ADDR_REG_4__SCAN_IN), .B2(n9805), .ZN(n10224) );
  NAND2_X1 U10946 ( .A1(P1_ADDR_REG_3__SCAN_IN), .A2(P2_ADDR_REG_3__SCAN_IN), 
        .ZN(n9811) );
  XNOR2_X1 U10947 ( .A(n9807), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(n10222) );
  NAND2_X1 U10948 ( .A1(P2_ADDR_REG_2__SCAN_IN), .A2(P1_ADDR_REG_2__SCAN_IN), 
        .ZN(n9810) );
  XNOR2_X1 U10949 ( .A(P2_ADDR_REG_2__SCAN_IN), .B(n9808), .ZN(n10220) );
  AOI21_X1 U10950 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(P2_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10177) );
  NAND3_X1 U10951 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .A3(P2_ADDR_REG_0__SCAN_IN), .ZN(n10179) );
  NAND2_X1 U10952 ( .A1(n10220), .A2(n10219), .ZN(n9809) );
  NAND2_X1 U10953 ( .A1(n9810), .A2(n9809), .ZN(n10221) );
  NOR2_X1 U10954 ( .A1(n10224), .A2(n10223), .ZN(n9812) );
  NOR2_X1 U10955 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n9814), .ZN(n10208) );
  NAND2_X1 U10956 ( .A1(n9816), .A2(P1_ADDR_REG_6__SCAN_IN), .ZN(n9818) );
  NAND2_X1 U10957 ( .A1(n10206), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n9817) );
  NAND2_X1 U10958 ( .A1(n9818), .A2(n9817), .ZN(n9819) );
  NAND2_X1 U10959 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n9819), .ZN(n9821) );
  NAND2_X1 U10960 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10218), .ZN(n9820) );
  NAND2_X1 U10961 ( .A1(n9821), .A2(n9820), .ZN(n9822) );
  NAND2_X1 U10962 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n9822), .ZN(n9825) );
  INV_X1 U10963 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n9823) );
  XNOR2_X1 U10964 ( .A(n9823), .B(n9822), .ZN(n10217) );
  NAND2_X1 U10965 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10217), .ZN(n9824) );
  AND2_X1 U10966 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n9826), .ZN(n9827) );
  NAND2_X1 U10967 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n9828) );
  OAI21_X1 U10968 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n9828), .ZN(n10204) );
  NAND2_X1 U10969 ( .A1(P1_ADDR_REG_11__SCAN_IN), .A2(P2_ADDR_REG_11__SCAN_IN), 
        .ZN(n9829) );
  OAI21_X1 U10970 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n9829), .ZN(n10201) );
  NOR2_X1 U10971 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n9830) );
  AOI21_X1 U10972 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n9830), .ZN(n10198) );
  NAND2_X1 U10973 ( .A1(n10199), .A2(n10198), .ZN(n10197) );
  NAND2_X1 U10974 ( .A1(n10196), .A2(n10195), .ZN(n10194) );
  NAND2_X1 U10975 ( .A1(n10193), .A2(n10192), .ZN(n10191) );
  OAI21_X1 U10976 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10188), .ZN(n10186) );
  NAND2_X1 U10977 ( .A1(n10187), .A2(n10186), .ZN(n10185) );
  OAI21_X1 U10978 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10185), .ZN(n10183) );
  NAND2_X1 U10979 ( .A1(n10184), .A2(n10183), .ZN(n10182) );
  NOR2_X1 U10980 ( .A1(n10212), .A2(n10211), .ZN(n9831) );
  NAND2_X1 U10981 ( .A1(n10212), .A2(n10211), .ZN(n10210) );
  XNOR2_X1 U10982 ( .A(n4796), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n9832) );
  XNOR2_X1 U10983 ( .A(n9833), .B(n9832), .ZN(ADD_1071_U4) );
  XOR2_X1 U10984 ( .A(n9834), .B(P1_WR_REG_SCAN_IN), .Z(U123) );
  XNOR2_X1 U10985 ( .A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .ZN(U126) );
  OAI21_X1 U10986 ( .B1(n9837), .B2(n9836), .A(n9835), .ZN(n9838) );
  INV_X1 U10987 ( .A(n9838), .ZN(n9851) );
  INV_X1 U10988 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n9843) );
  INV_X1 U10989 ( .A(n9839), .ZN(n9840) );
  OR2_X1 U10990 ( .A1(n9923), .A2(n9840), .ZN(n9841) );
  OAI211_X1 U10991 ( .C1(n9877), .C2(n9843), .A(n9842), .B(n9841), .ZN(n9844)
         );
  INV_X1 U10992 ( .A(n9844), .ZN(n9850) );
  AOI211_X1 U10993 ( .C1(n9847), .C2(n9846), .A(n9863), .B(n9845), .ZN(n9848)
         );
  INV_X1 U10994 ( .A(n9848), .ZN(n9849) );
  OAI211_X1 U10995 ( .C1(n9851), .C2(n9934), .A(n9850), .B(n9849), .ZN(
        P1_U3253) );
  OAI21_X1 U10996 ( .B1(n9854), .B2(n9853), .A(n9852), .ZN(n9855) );
  INV_X1 U10997 ( .A(n9855), .ZN(n9869) );
  INV_X1 U10998 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n9860) );
  INV_X1 U10999 ( .A(n9856), .ZN(n9857) );
  OR2_X1 U11000 ( .A1(n9923), .A2(n9857), .ZN(n9858) );
  OAI211_X1 U11001 ( .C1(n9877), .C2(n9860), .A(n9859), .B(n9858), .ZN(n9861)
         );
  INV_X1 U11002 ( .A(n9861), .ZN(n9868) );
  AOI211_X1 U11003 ( .C1(n9865), .C2(n9864), .A(n9863), .B(n9862), .ZN(n9866)
         );
  INV_X1 U11004 ( .A(n9866), .ZN(n9867) );
  OAI211_X1 U11005 ( .C1(n9869), .C2(n9934), .A(n9868), .B(n9867), .ZN(
        P1_U3254) );
  OAI21_X1 U11006 ( .B1(n9872), .B2(n9871), .A(n9870), .ZN(n9873) );
  INV_X1 U11007 ( .A(n9873), .ZN(n9883) );
  OR2_X1 U11008 ( .A1(n9923), .A2(n9874), .ZN(n9875) );
  OAI211_X1 U11009 ( .C1(n9877), .C2(n4345), .A(n9876), .B(n9875), .ZN(n9878)
         );
  INV_X1 U11010 ( .A(n9878), .ZN(n9882) );
  XNOR2_X1 U11011 ( .A(n9879), .B(P1_REG2_REG_14__SCAN_IN), .ZN(n9880) );
  NAND2_X1 U11012 ( .A1(n9880), .A2(n9929), .ZN(n9881) );
  OAI211_X1 U11013 ( .C1(n9883), .C2(n9934), .A(n9882), .B(n9881), .ZN(
        P1_U3255) );
  AOI21_X1 U11014 ( .B1(n9886), .B2(n9885), .A(n9884), .ZN(n9894) );
  OAI211_X1 U11015 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n9888), .A(n9911), .B(
        n9887), .ZN(n9893) );
  NAND2_X1 U11016 ( .A1(n9927), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n9892) );
  OAI211_X1 U11017 ( .C1(n9890), .C2(P1_REG2_REG_15__SCAN_IN), .A(n9929), .B(
        n9889), .ZN(n9891) );
  NAND4_X1 U11018 ( .A1(n9894), .A2(n9893), .A3(n9892), .A4(n9891), .ZN(
        P1_U3256) );
  NOR2_X1 U11019 ( .A1(n9923), .A2(n9895), .ZN(n9896) );
  AOI211_X1 U11020 ( .C1(n9927), .C2(P1_ADDR_REG_16__SCAN_IN), .A(n9897), .B(
        n9896), .ZN(n9906) );
  OAI211_X1 U11021 ( .C1(n9900), .C2(n9899), .A(n9911), .B(n9898), .ZN(n9905)
         );
  OAI211_X1 U11022 ( .C1(n9903), .C2(n9902), .A(n9929), .B(n9901), .ZN(n9904)
         );
  NAND3_X1 U11023 ( .A1(n9906), .A2(n9905), .A3(n9904), .ZN(P1_U3257) );
  NOR2_X1 U11024 ( .A1(n9923), .A2(n9907), .ZN(n9908) );
  AOI211_X1 U11025 ( .C1(n9927), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n9909), .B(
        n9908), .ZN(n9919) );
  OAI211_X1 U11026 ( .C1(n9913), .C2(n9912), .A(n9911), .B(n9910), .ZN(n9918)
         );
  OAI211_X1 U11027 ( .C1(n9916), .C2(n9915), .A(n9914), .B(n9929), .ZN(n9917)
         );
  NAND3_X1 U11028 ( .A1(n9919), .A2(n9918), .A3(n9917), .ZN(P1_U3258) );
  AOI21_X1 U11029 ( .B1(n9922), .B2(n9921), .A(n9920), .ZN(n9935) );
  NOR2_X1 U11030 ( .A1(n9924), .A2(n9923), .ZN(n9925) );
  AOI211_X1 U11031 ( .C1(n9927), .C2(P1_ADDR_REG_18__SCAN_IN), .A(n9926), .B(
        n9925), .ZN(n9933) );
  OAI211_X1 U11032 ( .C1(n9931), .C2(n9930), .A(n9929), .B(n9928), .ZN(n9932)
         );
  OAI211_X1 U11033 ( .C1(n9935), .C2(n9934), .A(n9933), .B(n9932), .ZN(
        P1_U3259) );
  AND2_X1 U11034 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n9943), .ZN(P1_U3292) );
  AND2_X1 U11035 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n9943), .ZN(P1_U3293) );
  NOR2_X1 U11036 ( .A1(n9942), .A2(n9936), .ZN(P1_U3294) );
  AND2_X1 U11037 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n9943), .ZN(P1_U3295) );
  NOR2_X1 U11038 ( .A1(n9942), .A2(n9937), .ZN(P1_U3296) );
  AND2_X1 U11039 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n9943), .ZN(P1_U3297) );
  AND2_X1 U11040 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n9943), .ZN(P1_U3298) );
  AND2_X1 U11041 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n9943), .ZN(P1_U3299) );
  AND2_X1 U11042 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n9943), .ZN(P1_U3300) );
  AND2_X1 U11043 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n9943), .ZN(P1_U3301) );
  AND2_X1 U11044 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n9943), .ZN(P1_U3302) );
  NOR2_X1 U11045 ( .A1(n9942), .A2(n9938), .ZN(P1_U3303) );
  AND2_X1 U11046 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n9943), .ZN(P1_U3304) );
  AND2_X1 U11047 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n9943), .ZN(P1_U3305) );
  AND2_X1 U11048 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n9943), .ZN(P1_U3306) );
  NOR2_X1 U11049 ( .A1(n9942), .A2(n9939), .ZN(P1_U3307) );
  AND2_X1 U11050 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n9943), .ZN(P1_U3308) );
  AND2_X1 U11051 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n9943), .ZN(P1_U3309) );
  AND2_X1 U11052 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n9943), .ZN(P1_U3310) );
  AND2_X1 U11053 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n9943), .ZN(P1_U3311) );
  NOR2_X1 U11054 ( .A1(n9942), .A2(n9940), .ZN(P1_U3312) );
  AND2_X1 U11055 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n9943), .ZN(P1_U3313) );
  AND2_X1 U11056 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n9943), .ZN(P1_U3314) );
  NOR2_X1 U11057 ( .A1(n9942), .A2(n9941), .ZN(P1_U3315) );
  AND2_X1 U11058 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n9943), .ZN(P1_U3316) );
  AND2_X1 U11059 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n9943), .ZN(P1_U3317) );
  AND2_X1 U11060 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n9943), .ZN(P1_U3318) );
  AND2_X1 U11061 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n9943), .ZN(P1_U3319) );
  AND2_X1 U11062 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n9943), .ZN(P1_U3320) );
  AND2_X1 U11063 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n9943), .ZN(P1_U3321) );
  NAND3_X1 U11064 ( .A1(n9946), .A2(n9945), .A3(n9944), .ZN(n9948) );
  NAND2_X1 U11065 ( .A1(n9948), .A2(n9947), .ZN(n9950) );
  AOI211_X1 U11066 ( .C1(n9979), .C2(n9951), .A(n9950), .B(n9949), .ZN(n9992)
         );
  AOI22_X1 U11067 ( .A1(n9991), .A2(n9992), .B1(n5145), .B2(n9990), .ZN(
        P1_U3460) );
  OAI22_X1 U11068 ( .A1(n9953), .A2(n9984), .B1(n9952), .B2(n9982), .ZN(n9955)
         );
  AOI211_X1 U11069 ( .C1(n9989), .C2(n9956), .A(n9955), .B(n9954), .ZN(n9993)
         );
  INV_X1 U11070 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9957) );
  AOI22_X1 U11071 ( .A1(n9991), .A2(n9993), .B1(n9957), .B2(n9990), .ZN(
        P1_U3463) );
  OAI22_X1 U11072 ( .A1(n9959), .A2(n9984), .B1(n9958), .B2(n9982), .ZN(n9960)
         );
  AOI21_X1 U11073 ( .B1(n9961), .B2(n9989), .A(n9960), .ZN(n9962) );
  AND2_X1 U11074 ( .A1(n9963), .A2(n9962), .ZN(n9995) );
  AOI22_X1 U11075 ( .A1(n9991), .A2(n9995), .B1(n5179), .B2(n9990), .ZN(
        P1_U3466) );
  OAI22_X1 U11076 ( .A1(n9965), .A2(n9984), .B1(n9964), .B2(n9982), .ZN(n9968)
         );
  INV_X1 U11077 ( .A(n9966), .ZN(n9967) );
  AOI211_X1 U11078 ( .C1(n9969), .C2(n9979), .A(n9968), .B(n9967), .ZN(n9997)
         );
  AOI22_X1 U11079 ( .A1(n9991), .A2(n9997), .B1(n5187), .B2(n9990), .ZN(
        P1_U3469) );
  OAI21_X1 U11080 ( .B1(n9971), .B2(n9982), .A(n9970), .ZN(n9973) );
  AOI211_X1 U11081 ( .C1(n9974), .C2(n9979), .A(n9973), .B(n9972), .ZN(n9998)
         );
  AOI22_X1 U11082 ( .A1(n9991), .A2(n9998), .B1(n5209), .B2(n9990), .ZN(
        P1_U3472) );
  OAI21_X1 U11083 ( .B1(n7482), .B2(n9982), .A(n9975), .ZN(n9977) );
  AOI211_X1 U11084 ( .C1(n9979), .C2(n9978), .A(n9977), .B(n9976), .ZN(n9999)
         );
  AOI22_X1 U11085 ( .A1(n9991), .A2(n9999), .B1(n9980), .B2(n9990), .ZN(
        P1_U3475) );
  INV_X1 U11086 ( .A(n9981), .ZN(n9983) );
  OAI22_X1 U11087 ( .A1(n9985), .A2(n9984), .B1(n9983), .B2(n9982), .ZN(n9987)
         );
  AOI211_X1 U11088 ( .C1(n9989), .C2(n9988), .A(n9987), .B(n9986), .ZN(n10002)
         );
  AOI22_X1 U11089 ( .A1(n9991), .A2(n10002), .B1(n5253), .B2(n9990), .ZN(
        P1_U3478) );
  AOI22_X1 U11090 ( .A1(n10003), .A2(n9992), .B1(n6792), .B2(n10000), .ZN(
        P1_U3525) );
  AOI22_X1 U11091 ( .A1(n10003), .A2(n9993), .B1(n6794), .B2(n10000), .ZN(
        P1_U3526) );
  INV_X1 U11092 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n9994) );
  AOI22_X1 U11093 ( .A1(n10003), .A2(n9995), .B1(n9994), .B2(n10000), .ZN(
        P1_U3527) );
  INV_X1 U11094 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n9996) );
  AOI22_X1 U11095 ( .A1(n10003), .A2(n9997), .B1(n9996), .B2(n10000), .ZN(
        P1_U3528) );
  AOI22_X1 U11096 ( .A1(n10003), .A2(n9998), .B1(n5213), .B2(n10000), .ZN(
        P1_U3529) );
  AOI22_X1 U11097 ( .A1(n10003), .A2(n9999), .B1(n6820), .B2(n10000), .ZN(
        P1_U3530) );
  AOI22_X1 U11098 ( .A1(n10003), .A2(n10002), .B1(n10001), .B2(n10000), .ZN(
        P1_U3531) );
  NAND2_X1 U11099 ( .A1(n10029), .A2(n10004), .ZN(n10006) );
  OAI211_X1 U11100 ( .C1(n10008), .C2(n10007), .A(n10006), .B(n10005), .ZN(
        n10014) );
  INV_X1 U11101 ( .A(n10009), .ZN(n10045) );
  AOI211_X1 U11102 ( .C1(n10012), .C2(n10011), .A(n10010), .B(n10045), .ZN(
        n10013) );
  AOI211_X1 U11103 ( .C1(n10052), .C2(n10015), .A(n10014), .B(n10013), .ZN(
        n10016) );
  OAI21_X1 U11104 ( .B1(n10055), .B2(n10017), .A(n10016), .ZN(P2_U3219) );
  AOI21_X1 U11105 ( .B1(n10036), .B2(n10019), .A(n10018), .ZN(n10033) );
  OR2_X1 U11106 ( .A1(n10021), .A2(n10020), .ZN(n10025) );
  OAI21_X1 U11107 ( .B1(n10023), .B2(n10022), .A(n10043), .ZN(n10024) );
  OAI21_X1 U11108 ( .B1(n10026), .B2(n10025), .A(n10024), .ZN(n10028) );
  NAND2_X1 U11109 ( .A1(n10028), .A2(n10027), .ZN(n10032) );
  NAND2_X1 U11110 ( .A1(n10052), .A2(n6126), .ZN(n10031) );
  NAND2_X1 U11111 ( .A1(n10029), .A2(n6673), .ZN(n10030) );
  AND4_X1 U11112 ( .A1(n10033), .A2(n10032), .A3(n10031), .A4(n10030), .ZN(
        n10034) );
  OAI21_X1 U11113 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n10055), .A(n10034), .ZN(
        P2_U3220) );
  AOI22_X1 U11114 ( .A1(n10036), .A2(n10035), .B1(P2_REG3_REG_11__SCAN_IN), 
        .B2(P2_U3152), .ZN(n10037) );
  OAI21_X1 U11115 ( .B1(n10039), .B2(n10038), .A(n10037), .ZN(n10050) );
  NAND3_X1 U11116 ( .A1(n10042), .A2(n10041), .A3(n10040), .ZN(n10048) );
  OAI21_X1 U11117 ( .B1(n10045), .B2(n10044), .A(n10043), .ZN(n10047) );
  AOI21_X1 U11118 ( .B1(n10048), .B2(n10047), .A(n10046), .ZN(n10049) );
  AOI211_X1 U11119 ( .C1(n10052), .C2(n10051), .A(n10050), .B(n10049), .ZN(
        n10053) );
  OAI21_X1 U11120 ( .B1(n10055), .B2(n10054), .A(n10053), .ZN(P2_U3238) );
  OAI21_X1 U11121 ( .B1(n10064), .B2(n10057), .A(n10056), .ZN(n10062) );
  AOI222_X1 U11122 ( .A1(n10080), .A2(n10062), .B1(n10061), .B2(n10060), .C1(
        n10059), .C2(n10058), .ZN(n10151) );
  INV_X1 U11123 ( .A(n10063), .ZN(n10067) );
  INV_X1 U11124 ( .A(n10064), .ZN(n10066) );
  OAI21_X1 U11125 ( .B1(n10067), .B2(n10066), .A(n10065), .ZN(n10154) );
  NAND2_X1 U11126 ( .A1(n10088), .A2(n10072), .ZN(n10068) );
  NAND2_X1 U11127 ( .A1(n10069), .A2(n10068), .ZN(n10150) );
  OAI22_X1 U11128 ( .A1(n10093), .A2(n6911), .B1(n10070), .B2(n10090), .ZN(
        n10071) );
  AOI21_X1 U11129 ( .B1(n10095), .B2(n10072), .A(n10071), .ZN(n10073) );
  OAI21_X1 U11130 ( .B1(n10074), .B2(n10150), .A(n10073), .ZN(n10075) );
  AOI21_X1 U11131 ( .B1(n10154), .B2(n10099), .A(n10075), .ZN(n10076) );
  OAI21_X1 U11132 ( .B1(n8717), .B2(n10151), .A(n10076), .ZN(P2_U3289) );
  OAI21_X1 U11133 ( .B1(n10087), .B2(n10078), .A(n10077), .ZN(n10081) );
  AOI21_X1 U11134 ( .B1(n10081), .B2(n10080), .A(n10079), .ZN(n10143) );
  NAND2_X1 U11135 ( .A1(n10083), .A2(n10082), .ZN(n10085) );
  NAND2_X1 U11136 ( .A1(n10085), .A2(n10084), .ZN(n10086) );
  XOR2_X1 U11137 ( .A(n10087), .B(n10086), .Z(n10146) );
  AOI21_X1 U11138 ( .B1(n7735), .B2(n10141), .A(n10149), .ZN(n10089) );
  NAND2_X1 U11139 ( .A1(n10089), .A2(n10088), .ZN(n10142) );
  OAI22_X1 U11140 ( .A1(n10093), .A2(n10092), .B1(n10091), .B2(n10090), .ZN(
        n10094) );
  AOI21_X1 U11141 ( .B1(n10095), .B2(n10141), .A(n10094), .ZN(n10096) );
  OAI21_X1 U11142 ( .B1(n10097), .B2(n10142), .A(n10096), .ZN(n10098) );
  AOI21_X1 U11143 ( .B1(n10146), .B2(n10099), .A(n10098), .ZN(n10100) );
  OAI21_X1 U11144 ( .B1(n8717), .B2(n10143), .A(n10100), .ZN(P2_U3290) );
  AND2_X1 U11145 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10108), .ZN(P2_U3297) );
  AND2_X1 U11146 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10108), .ZN(P2_U3298) );
  AND2_X1 U11147 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10108), .ZN(P2_U3299) );
  NOR2_X1 U11148 ( .A1(n10112), .A2(n10103), .ZN(P2_U3300) );
  NOR2_X1 U11149 ( .A1(n10112), .A2(n10104), .ZN(P2_U3301) );
  AND2_X1 U11150 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10108), .ZN(P2_U3302) );
  AND2_X1 U11151 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10108), .ZN(P2_U3303) );
  AND2_X1 U11152 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10108), .ZN(P2_U3304) );
  AND2_X1 U11153 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10108), .ZN(P2_U3305) );
  AND2_X1 U11154 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10108), .ZN(P2_U3306) );
  AND2_X1 U11155 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10108), .ZN(P2_U3307) );
  AND2_X1 U11156 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10108), .ZN(P2_U3308) );
  AND2_X1 U11157 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10108), .ZN(P2_U3309) );
  AND2_X1 U11158 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10108), .ZN(P2_U3310) );
  AND2_X1 U11159 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10108), .ZN(P2_U3311) );
  AND2_X1 U11160 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10108), .ZN(P2_U3312) );
  NOR2_X1 U11161 ( .A1(n10112), .A2(n10105), .ZN(P2_U3313) );
  AND2_X1 U11162 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10108), .ZN(P2_U3314) );
  AND2_X1 U11163 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10108), .ZN(P2_U3315) );
  AND2_X1 U11164 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10108), .ZN(P2_U3316) );
  AND2_X1 U11165 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10108), .ZN(P2_U3317) );
  NOR2_X1 U11166 ( .A1(n10112), .A2(n10106), .ZN(P2_U3318) );
  AND2_X1 U11167 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10108), .ZN(P2_U3319) );
  AND2_X1 U11168 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10108), .ZN(P2_U3320) );
  AND2_X1 U11169 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10108), .ZN(P2_U3321) );
  NOR2_X1 U11170 ( .A1(n10112), .A2(n10107), .ZN(P2_U3322) );
  AND2_X1 U11171 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10108), .ZN(P2_U3323) );
  AND2_X1 U11172 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10108), .ZN(P2_U3324) );
  AND2_X1 U11173 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10108), .ZN(P2_U3325) );
  AND2_X1 U11174 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10108), .ZN(P2_U3326) );
  AOI22_X1 U11175 ( .A1(n10110), .A2(n10111), .B1(n10109), .B2(n10108), .ZN(
        P2_U3437) );
  INV_X1 U11176 ( .A(n10111), .ZN(n10113) );
  OAI22_X1 U11177 ( .A1(n10114), .A2(n10113), .B1(P2_D_REG_1__SCAN_IN), .B2(
        n10112), .ZN(n10115) );
  INV_X1 U11178 ( .A(n10115), .ZN(P2_U3438) );
  AOI22_X1 U11179 ( .A1(n10118), .A2(n10155), .B1(n10117), .B2(n10116), .ZN(
        n10119) );
  AND2_X1 U11180 ( .A1(n10120), .A2(n10119), .ZN(n10167) );
  INV_X1 U11181 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n10121) );
  AOI22_X1 U11182 ( .A1(n10166), .A2(n10167), .B1(n10121), .B2(n10165), .ZN(
        P2_U3451) );
  AOI211_X1 U11183 ( .C1(n10155), .C2(n10124), .A(n10123), .B(n10122), .ZN(
        n10168) );
  INV_X1 U11184 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10125) );
  AOI22_X1 U11185 ( .A1(n10166), .A2(n10168), .B1(n10125), .B2(n10165), .ZN(
        P2_U3454) );
  INV_X1 U11186 ( .A(n10126), .ZN(n10127) );
  OAI21_X1 U11187 ( .B1(n10128), .B2(n10159), .A(n10127), .ZN(n10130) );
  AOI211_X1 U11188 ( .C1(n10155), .C2(n10131), .A(n10130), .B(n10129), .ZN(
        n10169) );
  INV_X1 U11189 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n10132) );
  AOI22_X1 U11190 ( .A1(n10166), .A2(n10169), .B1(n10132), .B2(n10165), .ZN(
        P2_U3460) );
  AOI211_X1 U11191 ( .C1(n10155), .C2(n10135), .A(n10134), .B(n10133), .ZN(
        n10170) );
  AOI22_X1 U11192 ( .A1(n10166), .A2(n10170), .B1(n6167), .B2(n10165), .ZN(
        P2_U3463) );
  OAI211_X1 U11193 ( .C1(n10138), .C2(n10159), .A(n10137), .B(n10136), .ZN(
        n10139) );
  AOI21_X1 U11194 ( .B1(n10155), .B2(n10140), .A(n10139), .ZN(n10171) );
  AOI22_X1 U11195 ( .A1(n10166), .A2(n10171), .B1(n6187), .B2(n10165), .ZN(
        P2_U3466) );
  INV_X1 U11196 ( .A(n10141), .ZN(n10144) );
  OAI211_X1 U11197 ( .C1(n10144), .C2(n10159), .A(n10143), .B(n10142), .ZN(
        n10145) );
  AOI21_X1 U11198 ( .B1(n10146), .B2(n10155), .A(n10145), .ZN(n10172) );
  INV_X1 U11199 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10147) );
  AOI22_X1 U11200 ( .A1(n10166), .A2(n10172), .B1(n10147), .B2(n10165), .ZN(
        P2_U3469) );
  OAI22_X1 U11201 ( .A1(n10150), .A2(n10149), .B1(n10148), .B2(n10159), .ZN(
        n10153) );
  INV_X1 U11202 ( .A(n10151), .ZN(n10152) );
  AOI211_X1 U11203 ( .C1(n10155), .C2(n10154), .A(n10153), .B(n10152), .ZN(
        n10173) );
  AOI22_X1 U11204 ( .A1(n10166), .A2(n10173), .B1(n6208), .B2(n10165), .ZN(
        P2_U3472) );
  AOI21_X1 U11205 ( .B1(n10158), .B2(n10157), .A(n10156), .ZN(n10164) );
  NOR2_X1 U11206 ( .A1(n10160), .A2(n10159), .ZN(n10163) );
  NOR4_X1 U11207 ( .A1(n10164), .A2(n10163), .A3(n10162), .A4(n10161), .ZN(
        n10175) );
  AOI22_X1 U11208 ( .A1(n10166), .A2(n10175), .B1(n6220), .B2(n10165), .ZN(
        P2_U3475) );
  AOI22_X1 U11209 ( .A1(n10176), .A2(n10167), .B1(n6136), .B2(n10174), .ZN(
        P2_U3520) );
  AOI22_X1 U11210 ( .A1(n10176), .A2(n10168), .B1(n6865), .B2(n10174), .ZN(
        P2_U3521) );
  AOI22_X1 U11211 ( .A1(n10176), .A2(n10169), .B1(n6869), .B2(n10174), .ZN(
        P2_U3523) );
  AOI22_X1 U11212 ( .A1(n10176), .A2(n10170), .B1(n6872), .B2(n10174), .ZN(
        P2_U3524) );
  AOI22_X1 U11213 ( .A1(n10176), .A2(n10171), .B1(n6875), .B2(n10174), .ZN(
        P2_U3525) );
  AOI22_X1 U11214 ( .A1(n10176), .A2(n10172), .B1(n6878), .B2(n10174), .ZN(
        P2_U3526) );
  AOI22_X1 U11215 ( .A1(n10176), .A2(n10173), .B1(n6899), .B2(n10174), .ZN(
        P2_U3527) );
  AOI22_X1 U11216 ( .A1(n10176), .A2(n10175), .B1(n6223), .B2(n10174), .ZN(
        P2_U3528) );
  INV_X1 U11217 ( .A(n10177), .ZN(n10178) );
  NAND2_X1 U11218 ( .A1(n10179), .A2(n10178), .ZN(n10180) );
  XOR2_X1 U11219 ( .A(n10181), .B(n10180), .Z(ADD_1071_U5) );
  XOR2_X1 U11220 ( .A(P1_ADDR_REG_0__SCAN_IN), .B(P2_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  OAI21_X1 U11221 ( .B1(n10184), .B2(n10183), .A(n10182), .ZN(ADD_1071_U56) );
  OAI21_X1 U11222 ( .B1(n10187), .B2(n10186), .A(n10185), .ZN(ADD_1071_U57) );
  OAI21_X1 U11223 ( .B1(n10190), .B2(n10189), .A(n10188), .ZN(ADD_1071_U58) );
  OAI21_X1 U11224 ( .B1(n10193), .B2(n10192), .A(n10191), .ZN(ADD_1071_U59) );
  OAI21_X1 U11225 ( .B1(n10196), .B2(n10195), .A(n10194), .ZN(ADD_1071_U60) );
  OAI21_X1 U11226 ( .B1(n10199), .B2(n10198), .A(n10197), .ZN(ADD_1071_U61) );
  AOI21_X1 U11227 ( .B1(n10202), .B2(n10201), .A(n10200), .ZN(ADD_1071_U62) );
  AOI21_X1 U11228 ( .B1(n10205), .B2(n10204), .A(n10203), .ZN(ADD_1071_U63) );
  XOR2_X1 U11229 ( .A(n10206), .B(P2_ADDR_REG_6__SCAN_IN), .Z(ADD_1071_U50) );
  NOR2_X1 U11230 ( .A1(n10208), .A2(n10207), .ZN(n10209) );
  XOR2_X1 U11231 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n10209), .Z(ADD_1071_U51) );
  OAI21_X1 U11232 ( .B1(n10212), .B2(n10211), .A(n10210), .ZN(n10213) );
  XNOR2_X1 U11233 ( .A(n10213), .B(P1_ADDR_REG_18__SCAN_IN), .ZN(ADD_1071_U55)
         );
  AOI21_X1 U11234 ( .B1(n10216), .B2(n10215), .A(n10214), .ZN(ADD_1071_U47) );
  XOR2_X1 U11235 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10217), .Z(ADD_1071_U48) );
  XOR2_X1 U11236 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10218), .Z(ADD_1071_U49) );
  XOR2_X1 U11237 ( .A(n10220), .B(n10219), .Z(ADD_1071_U54) );
  XOR2_X1 U11238 ( .A(n10222), .B(n10221), .Z(ADD_1071_U53) );
  XNOR2_X1 U11239 ( .A(n10224), .B(n10223), .ZN(ADD_1071_U52) );
  NAND2_X1 U4752 ( .A1(n6859), .A2(n4440), .ZN(n6322) );
  CLKBUF_X2 U4757 ( .A(n6120), .Z(n6457) );
  CLKBUF_X1 U5550 ( .A(n6448), .Z(n6449) );
  CLKBUF_X1 U8154 ( .A(n8399), .Z(n4363) );
endmodule

