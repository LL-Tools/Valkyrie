

module b15_C_AntiSAT_k_128_7 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757;

  NAND2_X1 U34510 ( .A1(n5509), .A2(n5060), .ZN(n4351) );
  CLKBUF_X2 U34520 ( .A(n3207), .Z(n3814) );
  INV_X1 U34530 ( .A(n5060), .ZN(n5467) );
  BUF_X1 U3454 ( .A(n3919), .Z(n4006) );
  CLKBUF_X2 U34550 ( .A(n3939), .Z(n3956) );
  CLKBUF_X2 U34560 ( .A(n3280), .Z(n3822) );
  CLKBUF_X2 U3458 ( .A(n3136), .Z(n3748) );
  CLKBUF_X2 U34590 ( .A(n3134), .Z(n3815) );
  CLKBUF_X2 U34600 ( .A(n3125), .Z(n3823) );
  BUF_X2 U34610 ( .A(n3182), .Z(n5063) );
  AND2_X2 U34620 ( .A1(n4109), .A2(n4070), .ZN(n3128) );
  AND2_X2 U34630 ( .A1(n4067), .A2(n4068), .ZN(n3281) );
  CLKBUF_X1 U34640 ( .A(n6098), .Z(n3003) );
  NOR2_X1 U34650 ( .A1(n5067), .A2(n5066), .ZN(n6098) );
  CLKBUF_X2 U3466 ( .A(n3180), .Z(n4164) );
  INV_X1 U3467 ( .A(n3555), .ZN(n5424) );
  AND2_X1 U34680 ( .A1(n4183), .A2(n4230), .ZN(n3357) );
  CLKBUF_X2 U34690 ( .A(n3223), .Z(n3776) );
  XNOR2_X1 U34700 ( .A(n3271), .B(n3270), .ZN(n4103) );
  INV_X1 U34710 ( .A(n5445), .ZN(n5495) );
  AND2_X2 U34720 ( .A1(n4112), .A2(n3153), .ZN(n5060) );
  INV_X1 U34730 ( .A(n6038), .ZN(n6073) );
  NAND2_X1 U34740 ( .A1(n4351), .A2(n3916), .ZN(n4190) );
  INV_X1 U3475 ( .A(n6108), .ZN(n6094) );
  AND2_X4 U3476 ( .A1(n3041), .A2(n4070), .ZN(n3017) );
  AND2_X2 U3477 ( .A1(n3035), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4068)
         );
  AND2_X2 U3478 ( .A1(n3153), .A2(n3155), .ZN(n3182) );
  NAND2_X2 U3479 ( .A1(n4816), .A2(n4815), .ZN(n4827) );
  NAND2_X2 U3480 ( .A1(n4762), .A2(n4761), .ZN(n4816) );
  NAND4_X4 U3481 ( .A1(n3098), .A2(n3097), .A3(n3096), .A4(n3095), .ZN(n3153)
         );
  AND4_X2 U3482 ( .A1(n3082), .A2(n3081), .A3(n3080), .A4(n3079), .ZN(n3098)
         );
  NAND2_X4 U3483 ( .A1(n3068), .A2(n3067), .ZN(n3163) );
  AND2_X4 U3484 ( .A1(n3019), .A2(n3077), .ZN(n3142) );
  NAND2_X2 U3485 ( .A1(n3159), .A2(n3158), .ZN(n4064) );
  NAND2_X2 U3486 ( .A1(n3048), .A2(n3047), .ZN(n3157) );
  AND4_X2 U3487 ( .A1(n3046), .A2(n3045), .A3(n3044), .A4(n3043), .ZN(n3047)
         );
  NAND2_X2 U3488 ( .A1(n3058), .A2(n3057), .ZN(n3161) );
  AND4_X2 U3489 ( .A1(n3056), .A2(n3055), .A3(n3054), .A4(n3053), .ZN(n3057)
         );
  AND4_X2 U3490 ( .A1(n3052), .A2(n3051), .A3(n3050), .A4(n3049), .ZN(n3058)
         );
  AND2_X2 U3491 ( .A1(n5625), .A2(n5626), .ZN(n5598) );
  OAI22_X2 U3492 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n5605), .B1(n5620), .B2(n5599), .ZN(n5600) );
  OAI21_X2 U3493 ( .B1(n5891), .B2(INSTADDRPOINTER_REG_21__SCAN_IN), .A(n5624), 
        .ZN(n5620) );
  INV_X2 U3494 ( .A(n5598), .ZN(n5624) );
  NAND2_X1 U3495 ( .A1(n6191), .A2(n4272), .ZN(n4280) );
  NAND2_X1 U3496 ( .A1(n6193), .A2(n6192), .ZN(n6191) );
  NOR2_X2 U3497 ( .A1(n5384), .A2(n4395), .ZN(n6287) );
  AND2_X1 U3498 ( .A1(n4184), .A2(n3356), .ZN(n4227) );
  NAND2_X1 U3499 ( .A1(n4156), .A2(n4508), .ZN(n4173) );
  AND2_X2 U3500 ( .A1(n3898), .A2(n3897), .ZN(n4506) );
  AND2_X1 U3501 ( .A1(n3119), .A2(n4162), .ZN(n3178) );
  INV_X2 U3502 ( .A(n3153), .ZN(n3180) );
  CLKBUF_X2 U3503 ( .A(n3127), .Z(n3817) );
  CLKBUF_X2 U3504 ( .A(n3128), .Z(n3813) );
  CLKBUF_X1 U3505 ( .A(n5582), .Z(n3006) );
  CLKBUF_X1 U3506 ( .A(n5416), .Z(n5417) );
  AOI21_X1 U3507 ( .B1(n5632), .B2(n5631), .A(n5597), .ZN(n5625) );
  AOI211_X1 U3508 ( .C1(n6177), .C2(n5578), .A(n5577), .B(n5576), .ZN(n5579)
         );
  CLKBUF_X1 U3509 ( .A(n5356), .Z(n5315) );
  INV_X1 U3510 ( .A(n3010), .ZN(n5098) );
  NOR2_X2 U3511 ( .A1(n5545), .A2(n5536), .ZN(n5537) );
  AND2_X1 U3512 ( .A1(n5721), .A2(n5398), .ZN(n5715) );
  AND2_X1 U3513 ( .A1(n5604), .A2(n5770), .ZN(n5721) );
  NAND2_X1 U3514 ( .A1(n3401), .A2(n3400), .ZN(n4646) );
  NOR2_X1 U3515 ( .A1(n5952), .A2(n5953), .ZN(n5934) );
  NOR2_X1 U3516 ( .A1(n3787), .A2(n5564), .ZN(n3788) );
  INV_X1 U3517 ( .A(n4472), .ZN(n3015) );
  NOR2_X1 U3518 ( .A1(n4324), .A2(n4471), .ZN(n6376) );
  NAND2_X2 U3519 ( .A1(n6123), .A2(n3163), .ZN(n6118) );
  NAND2_X1 U3520 ( .A1(n3329), .A2(n3328), .ZN(n4545) );
  NAND2_X2 U3521 ( .A1(n3253), .A2(n3029), .ZN(n4140) );
  XNOR2_X1 U3522 ( .A(n3296), .B(n3295), .ZN(n3305) );
  NAND2_X1 U3523 ( .A1(n3938), .A2(n3937), .ZN(n4780) );
  XNOR2_X1 U3524 ( .A(n4445), .B(n4547), .ZN(n4054) );
  INV_X1 U3525 ( .A(n4368), .ZN(n3938) );
  OR2_X1 U3526 ( .A1(n3309), .A2(n3308), .ZN(n4445) );
  NOR2_X1 U3527 ( .A1(n3641), .A2(n5633), .ZN(n3642) );
  AND2_X1 U3528 ( .A1(n3249), .A2(n3251), .ZN(n3250) );
  AOI21_X1 U3529 ( .B1(n3272), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n3168), 
        .ZN(n3166) );
  INV_X1 U3530 ( .A(n4367), .ZN(n3937) );
  AND2_X1 U3531 ( .A1(n3928), .A2(n3927), .ZN(n4354) );
  AND3_X1 U3532 ( .A1(n3217), .A2(n3216), .A3(n3215), .ZN(n3259) );
  NOR2_X2 U3533 ( .A1(n3186), .A2(n4319), .ZN(n4037) );
  CLKBUF_X1 U3534 ( .A(n3186), .Z(n3843) );
  AND3_X1 U3535 ( .A1(n3178), .A2(n3123), .A3(n4088), .ZN(n3147) );
  AND2_X1 U3536 ( .A1(n3174), .A2(n5063), .ZN(n4089) );
  NOR2_X1 U3537 ( .A1(n3441), .A2(n6690), .ZN(n3489) );
  NOR2_X1 U3538 ( .A1(n4319), .A2(n3160), .ZN(n3901) );
  NAND2_X1 U3539 ( .A1(n3179), .A2(n3157), .ZN(n3484) );
  CLKBUF_X1 U3540 ( .A(n3155), .Z(n4144) );
  CLKBUF_X1 U3541 ( .A(n3161), .Z(n3162) );
  OR2_X1 U3542 ( .A1(n3214), .A2(n3213), .ZN(n4823) );
  INV_X1 U3543 ( .A(n3161), .ZN(n3179) );
  AND2_X1 U3544 ( .A1(n3024), .A2(n3031), .ZN(n4146) );
  AND4_X1 U3545 ( .A1(n3040), .A2(n3039), .A3(n3038), .A4(n3037), .ZN(n3048)
         );
  AND4_X1 U3546 ( .A1(n3066), .A2(n3065), .A3(n3064), .A4(n3063), .ZN(n3067)
         );
  AND4_X1 U3547 ( .A1(n3076), .A2(n3075), .A3(n3074), .A4(n3073), .ZN(n3077)
         );
  INV_X2 U3548 ( .A(n5679), .ZN(n6205) );
  AND4_X1 U3549 ( .A1(n3090), .A2(n3089), .A3(n3088), .A4(n3087), .ZN(n3096)
         );
  AND4_X1 U3550 ( .A1(n3086), .A2(n3085), .A3(n3084), .A4(n3083), .ZN(n3097)
         );
  BUF_X2 U3551 ( .A(n3126), .Z(n3824) );
  BUF_X2 U3552 ( .A(n3135), .Z(n3816) );
  BUF_X2 U3553 ( .A(n3281), .Z(n3004) );
  NOR2_X1 U3554 ( .A1(n3351), .A2(n3350), .ZN(n3349) );
  CLKBUF_X1 U3555 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n4073) );
  NOR2_X2 U3556 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n4551) );
  AND2_X2 U3557 ( .A1(n5329), .A2(n5070), .ZN(n6108) );
  CLKBUF_X1 U3558 ( .A(n6185), .Z(n3005) );
  NAND2_X1 U3559 ( .A1(n5416), .A2(n5373), .ZN(n5582) );
  NAND2_X1 U3560 ( .A1(n4733), .A2(n4264), .ZN(n6193) );
  NAND2_X1 U3561 ( .A1(n5372), .A2(n5371), .ZN(n5416) );
  AND2_X2 U3562 ( .A1(n4936), .A2(n5038), .ZN(n5037) );
  CLKBUF_X1 U3563 ( .A(n4742), .Z(n3007) );
  AND2_X1 U3564 ( .A1(n5037), .A2(n3611), .ZN(n3008) );
  AND2_X1 U3565 ( .A1(n5037), .A2(n3611), .ZN(n5201) );
  AND4_X1 U3566 ( .A1(n3062), .A2(n3061), .A3(n3060), .A4(n3059), .ZN(n3068)
         );
  AND2_X1 U3567 ( .A1(n4255), .A2(n4254), .ZN(n4734) );
  AOI21_X1 U3568 ( .B1(n4253), .B2(n4753), .A(n4252), .ZN(n6200) );
  AND2_X4 U3570 ( .A1(n4109), .A2(n4458), .ZN(n3133) );
  AOI22_X2 U3571 ( .A1(n3136), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3106) );
  XNOR2_X2 U3572 ( .A(n3916), .B(n4174), .ZN(n5509) );
  NAND2_X2 U3573 ( .A1(n3304), .A2(n4185), .ZN(n4183) );
  NAND2_X1 U3574 ( .A1(n4826), .A2(n4827), .ZN(n3009) );
  NAND2_X1 U3575 ( .A1(n4827), .A2(n4826), .ZN(n4931) );
  NOR2_X2 U3576 ( .A1(n3380), .A2(n3379), .ZN(n3403) );
  NAND2_X1 U3577 ( .A1(n3360), .A2(n3359), .ZN(n3380) );
  NAND2_X1 U3578 ( .A1(n3954), .A2(n3953), .ZN(n5109) );
  NAND2_X1 U3579 ( .A1(n3967), .A2(n3966), .ZN(n5930) );
  NAND2_X2 U3580 ( .A1(n5531), .A2(n5522), .ZN(n5524) );
  AND2_X2 U3581 ( .A1(n5537), .A2(n5529), .ZN(n5531) );
  AND2_X2 U3582 ( .A1(n4067), .A2(n4458), .ZN(n3223) );
  AND2_X4 U3583 ( .A1(n3041), .A2(n3042), .ZN(n3127) );
  INV_X2 U3584 ( .A(n4009), .ZN(n5204) );
  AND2_X2 U3585 ( .A1(n5044), .A2(n5043), .ZN(n3010) );
  NAND2_X1 U3586 ( .A1(n3009), .A2(n4930), .ZN(n3011) );
  CLKBUF_X1 U3587 ( .A(n5607), .Z(n3012) );
  OAI21_X1 U3588 ( .B1(n5274), .B2(n5273), .A(n5272), .ZN(n3013) );
  AOI21_X1 U3589 ( .B1(n3267), .B2(n3266), .A(n3265), .ZN(n3014) );
  OAI21_X1 U3590 ( .B1(n5274), .B2(n5273), .A(n5272), .ZN(n5312) );
  AOI21_X1 U3591 ( .B1(n3267), .B2(n3266), .A(n3265), .ZN(n3306) );
  XNOR2_X1 U3592 ( .A(n3297), .B(n3305), .ZN(n4253) );
  NOR2_X2 U3593 ( .A1(n4937), .A2(n4938), .ZN(n4936) );
  AND2_X1 U3594 ( .A1(n4070), .A2(n4067), .ZN(n3016) );
  NAND2_X2 U3595 ( .A1(n3268), .A2(n3170), .ZN(n3271) );
  OR2_X2 U3596 ( .A1(n5731), .A2(n5543), .ZN(n5545) );
  NOR2_X2 U3597 ( .A1(n5582), .A2(n5891), .ZN(n5561) );
  OR2_X4 U3598 ( .A1(n3108), .A2(n3107), .ZN(n4112) );
  NOR3_X4 U3599 ( .A1(n5445), .A2(n5442), .A3(n3023), .ZN(n4019) );
  OR2_X4 U3600 ( .A1(n5524), .A2(n5496), .ZN(n5445) );
  OAI21_X1 U3601 ( .B1(n4157), .B2(n3165), .A(STATE2_REG_0__SCAN_IN), .ZN(
        n3167) );
  OAI21_X1 U3602 ( .B1(n4034), .B2(n3164), .A(n4170), .ZN(n3165) );
  CLKBUF_X1 U3603 ( .A(n3282), .Z(n3222) );
  CLKBUF_X1 U3604 ( .A(n3228), .Z(n3799) );
  AND2_X1 U3605 ( .A1(n4055), .A2(n3121), .ZN(n3123) );
  XNOR2_X1 U3606 ( .A(n4821), .B(n3405), .ZN(n4754) );
  INV_X1 U3607 ( .A(n4220), .ZN(n3376) );
  INV_X1 U3608 ( .A(n4219), .ZN(n3377) );
  OR2_X1 U3609 ( .A1(n4216), .A2(n4187), .ZN(n4184) );
  NAND2_X1 U3610 ( .A1(n3403), .A2(n3402), .ZN(n4821) );
  NAND2_X1 U3611 ( .A1(n3923), .A2(n3922), .ZN(n4191) );
  NAND2_X1 U3612 ( .A1(n3263), .A2(n3260), .ZN(n3218) );
  AOI21_X1 U3613 ( .B1(n3243), .B2(n3251), .A(n4817), .ZN(n3266) );
  OR2_X1 U3614 ( .A1(n4372), .A2(n4034), .ZN(n4051) );
  OR2_X1 U3615 ( .A1(n4506), .A2(n6443), .ZN(n4372) );
  NOR2_X2 U3616 ( .A1(n5451), .A2(n5453), .ZN(n5452) );
  NAND2_X1 U3617 ( .A1(n3726), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3764)
         );
  BUF_X1 U3618 ( .A(n5037), .Z(n5139) );
  NAND2_X1 U3619 ( .A1(n4356), .A2(n4222), .ZN(n4368) );
  NOR2_X2 U3620 ( .A1(n4361), .A2(n4354), .ZN(n4356) );
  NOR2_X1 U3621 ( .A1(n5940), .A2(n5961), .ZN(n5384) );
  OR2_X1 U3622 ( .A1(n4173), .A2(n4161), .ZN(n6212) );
  AOI21_X1 U3623 ( .B1(n4295), .B2(n5050), .A(n3294), .ZN(n3296) );
  INV_X1 U3624 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n5050) );
  NAND2_X1 U3625 ( .A1(n5514), .A2(n6086), .ZN(n5475) );
  NAND2_X1 U3626 ( .A1(n5058), .A2(n5329), .ZN(n6038) );
  OR2_X1 U3627 ( .A1(n5346), .A2(n5546), .ZN(n4022) );
  AND2_X2 U3628 ( .A1(n3905), .A2(n4508), .ZN(n6123) );
  XNOR2_X1 U3629 ( .A(n5452), .B(n3841), .ZN(n5380) );
  INV_X1 U3630 ( .A(n5422), .ZN(n3841) );
  NAND2_X1 U3631 ( .A1(n6421), .A2(n4508), .ZN(n6181) );
  CLKBUF_X1 U3632 ( .A(n4292), .Z(n5778) );
  NOR2_X1 U3633 ( .A1(n3874), .A2(n3884), .ZN(n3883) );
  OR2_X1 U3634 ( .A1(n3326), .A2(n3325), .ZN(n4266) );
  NAND2_X1 U3635 ( .A1(n3900), .A2(n3078), .ZN(n3156) );
  AND2_X1 U3636 ( .A1(n3163), .A2(n3142), .ZN(n3078) );
  CLKBUF_X1 U3637 ( .A(n3208), .Z(n3287) );
  OR2_X1 U3638 ( .A1(n3370), .A2(n3369), .ZN(n4745) );
  OR2_X1 U3639 ( .A1(n3340), .A2(n3339), .ZN(n4744) );
  OR2_X1 U3640 ( .A1(n3201), .A2(n3200), .ZN(n4248) );
  OR2_X1 U3641 ( .A1(n3235), .A2(n3234), .ZN(n4247) );
  AND2_X1 U3642 ( .A1(n5071), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3869) );
  INV_X1 U3643 ( .A(n3856), .ZN(n3890) );
  AOI21_X1 U3644 ( .B1(n3484), .B2(n3160), .A(n5433), .ZN(n3144) );
  AOI22_X1 U3645 ( .A1(n3128), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3126), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3056) );
  AND2_X1 U3646 ( .A1(n3316), .A2(n3315), .ZN(n3874) );
  NAND2_X1 U3647 ( .A1(n4112), .A2(n3180), .ZN(n4055) );
  NAND2_X1 U3648 ( .A1(n5492), .A2(n5494), .ZN(n5451) );
  OR2_X1 U3649 ( .A1(n3688), .A2(n5838), .ZN(n3689) );
  INV_X1 U3650 ( .A(n5589), .ZN(n5371) );
  OR2_X1 U3651 ( .A1(n5657), .A2(n5357), .ZN(n5645) );
  AND2_X1 U3652 ( .A1(n5363), .A2(n5658), .ZN(n5367) );
  OR2_X1 U3653 ( .A1(n5647), .A2(n5362), .ZN(n5657) );
  AND2_X1 U3654 ( .A1(n5163), .A2(n5938), .ZN(n5362) );
  NAND2_X1 U3656 ( .A1(n3160), .A2(n4146), .ZN(n4236) );
  INV_X1 U3657 ( .A(n4818), .ZN(n4753) );
  AOI22_X1 U3658 ( .A1(n3127), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3223), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3073) );
  NAND2_X1 U3659 ( .A1(n4164), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3315) );
  NAND2_X1 U3660 ( .A1(n4308), .A2(n3869), .ZN(n3856) );
  NOR2_X1 U3661 ( .A1(n3293), .A2(n3292), .ZN(n4257) );
  NAND2_X1 U3662 ( .A1(n3278), .A2(n3277), .ZN(n3307) );
  NAND2_X1 U3663 ( .A1(n3272), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3278) );
  BUF_X1 U3664 ( .A(n3268), .Z(n3269) );
  NAND2_X1 U3665 ( .A1(n3250), .A2(n3252), .ZN(n3253) );
  OAI21_X1 U3666 ( .B1(n6555), .B2(n6429), .A(n6438), .ZN(n4301) );
  INV_X1 U3667 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n4787) );
  OR2_X1 U3668 ( .A1(n3521), .A2(n5295), .ZN(n3506) );
  NAND2_X1 U3669 ( .A1(n5329), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5067) );
  INV_X1 U3670 ( .A(n5067), .ZN(n5473) );
  BUF_X1 U3671 ( .A(n5451), .Z(n5493) );
  AND2_X1 U3672 ( .A1(n3725), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3726)
         );
  AND2_X1 U3673 ( .A1(n3729), .A2(n3728), .ZN(n5535) );
  NOR2_X1 U3674 ( .A1(n3689), .A2(n5609), .ZN(n3725) );
  AND2_X2 U3675 ( .A1(n5201), .A2(n5202), .ZN(n5265) );
  INV_X1 U3676 ( .A(n3605), .ZN(n3606) );
  NAND2_X1 U3677 ( .A1(n3607), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3641)
         );
  AND2_X1 U3678 ( .A1(n3502), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3587)
         );
  NAND2_X1 U3679 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n3587), .ZN(n3605)
         );
  AND2_X1 U3680 ( .A1(n5177), .A2(n5137), .ZN(n5281) );
  OR2_X1 U3681 ( .A1(n5288), .A2(n5289), .ZN(n5286) );
  NAND2_X1 U3682 ( .A1(n3489), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3556)
         );
  OR2_X1 U3683 ( .A1(n3440), .A2(n6043), .ZN(n3441) );
  NAND2_X1 U3684 ( .A1(n4844), .A2(n3439), .ZN(n4937) );
  NOR2_X1 U3685 ( .A1(n3419), .A2(n5151), .ZN(n3423) );
  AOI21_X1 U3686 ( .B1(n4754), .B2(n3567), .A(n3408), .ZN(n4647) );
  NOR2_X1 U3687 ( .A1(n3394), .A2(n5117), .ZN(n3395) );
  INV_X1 U3688 ( .A(n4364), .ZN(n3400) );
  INV_X1 U3689 ( .A(n4218), .ZN(n3401) );
  AOI21_X1 U3690 ( .B1(n4273), .B2(n3567), .A(n3375), .ZN(n4220) );
  NAND2_X1 U3691 ( .A1(n3349), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3394)
         );
  INV_X1 U3692 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3351) );
  NAND2_X1 U3693 ( .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n3350) );
  NAND2_X1 U3694 ( .A1(n3248), .A2(n3247), .ZN(n4214) );
  NAND2_X1 U3695 ( .A1(n5730), .A2(n5729), .ZN(n5731) );
  OR2_X1 U3696 ( .A1(n5362), .A2(n5648), .ZN(n5658) );
  INV_X1 U3697 ( .A(n5293), .ZN(n3967) );
  OR2_X1 U3698 ( .A1(n5163), .A2(n5952), .ZN(n5668) );
  NOR2_X1 U3699 ( .A1(n5163), .A2(n6223), .ZN(n5273) );
  INV_X1 U3700 ( .A(n4846), .ZN(n3954) );
  INV_X1 U3701 ( .A(n5163), .ZN(n5891) );
  OR2_X1 U3702 ( .A1(n5163), .A2(n6225), .ZN(n5043) );
  NAND2_X1 U3703 ( .A1(n3925), .A2(n3027), .ZN(n4361) );
  INV_X1 U3704 ( .A(n4190), .ZN(n3925) );
  OR2_X1 U3705 ( .A1(n4173), .A2(n4452), .ZN(n5944) );
  AND2_X1 U3706 ( .A1(n3264), .A2(n3263), .ZN(n3265) );
  INV_X1 U3707 ( .A(n6103), .ZN(n5223) );
  OR2_X1 U3708 ( .A1(n4786), .A2(n5778), .ZN(n4784) );
  OR2_X1 U3709 ( .A1(n4784), .A2(n4892), .ZN(n4617) );
  CLKBUF_X1 U3710 ( .A(n3153), .Z(n5071) );
  BUF_X1 U3711 ( .A(n3157), .Z(n4329) );
  NAND2_X1 U3712 ( .A1(n4052), .A2(n4051), .ZN(n6549) );
  INV_X1 U3713 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n5117) );
  NAND2_X1 U3714 ( .A1(n5329), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6078) );
  CLKBUF_X1 U3715 ( .A(n4103), .Z(n4104) );
  CLKBUF_X1 U3716 ( .A(n3254), .Z(n3255) );
  INV_X1 U3717 ( .A(n3163), .ZN(n5433) );
  INV_X1 U3718 ( .A(n5867), .ZN(n6128) );
  AND2_X1 U3719 ( .A1(n5432), .A2(n5157), .ZN(n6131) );
  INV_X2 U3720 ( .A(n5432), .ZN(n6130) );
  AND2_X1 U3721 ( .A1(n5432), .A2(n4210), .ZN(n5301) );
  INV_X1 U3722 ( .A(n5301), .ZN(n5088) );
  AND2_X1 U3723 ( .A1(n4375), .A2(n6431), .ZN(n6162) );
  CLKBUF_X1 U3724 ( .A(n6160), .Z(n6552) );
  INV_X1 U3725 ( .A(n4374), .ZN(n6173) );
  NAND2_X1 U3726 ( .A1(n4115), .A2(n4114), .ZN(n6172) );
  INV_X1 U3727 ( .A(n6172), .ZN(n4199) );
  OR2_X1 U3728 ( .A1(n5056), .A2(n5350), .ZN(n5057) );
  AND2_X1 U3729 ( .A1(n5902), .A2(n5901), .ZN(n6124) );
  AND2_X1 U3730 ( .A1(n6181), .A2(n4510), .ZN(n6199) );
  INV_X1 U3731 ( .A(n6199), .ZN(n5651) );
  OR2_X1 U3732 ( .A1(n5726), .A2(n5394), .ZN(n5703) );
  INV_X1 U3733 ( .A(n6260), .ZN(n6216) );
  INV_X1 U3734 ( .A(n5906), .ZN(n6284) );
  INV_X1 U3735 ( .A(n6216), .ZN(n6277) );
  INV_X1 U3736 ( .A(n6212), .ZN(n6280) );
  INV_X1 U3737 ( .A(n6217), .ZN(n6279) );
  INV_X1 U3738 ( .A(n5944), .ZN(n5961) );
  CLKBUF_X1 U3739 ( .A(n4295), .Z(n5328) );
  CLKBUF_X1 U3740 ( .A(n4054), .Z(n6103) );
  INV_X1 U3741 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6718) );
  CLKBUF_X1 U3742 ( .A(n5005), .Z(n6298) );
  OR2_X1 U3743 ( .A1(n4580), .A2(n5004), .ZN(n6366) );
  INV_X1 U3744 ( .A(n4959), .ZN(n6375) );
  INV_X1 U3745 ( .A(n4977), .ZN(n6329) );
  INV_X1 U3746 ( .A(n4954), .ZN(n6381) );
  INV_X1 U3747 ( .A(n4987), .ZN(n6339) );
  INV_X1 U3748 ( .A(n4964), .ZN(n6389) );
  INV_X1 U3749 ( .A(n4981), .ZN(n6356) );
  INV_X1 U3750 ( .A(n4478), .ZN(n4541) );
  INV_X1 U3751 ( .A(n5407), .ZN(n6438) );
  INV_X1 U3752 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6532) );
  OAI211_X1 U3753 ( .C1(n5480), .C2(n5479), .A(n3021), .B(n5478), .ZN(n5481)
         );
  AND2_X1 U3754 ( .A1(n4022), .A2(n4021), .ZN(n4023) );
  NAND2_X1 U3755 ( .A1(n5380), .A2(n3906), .ZN(n4024) );
  INV_X1 U3756 ( .A(n4112), .ZN(n3155) );
  OR2_X1 U3757 ( .A1(n3152), .A2(n3153), .ZN(n3018) );
  INV_X1 U3758 ( .A(n3160), .ZN(n3907) );
  NAND2_X1 U3759 ( .A1(n5265), .A2(n5264), .ZN(n5263) );
  NAND2_X2 U3760 ( .A1(n4821), .A2(n4820), .ZN(n5163) );
  AND4_X1 U3761 ( .A1(n3072), .A2(n3071), .A3(n3070), .A4(n3069), .ZN(n3019)
         );
  BUF_X1 U3762 ( .A(n4256), .Z(n3348) );
  NOR2_X2 U3763 ( .A1(n5528), .A2(n5520), .ZN(n5492) );
  INV_X1 U3764 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3256) );
  NAND2_X1 U3765 ( .A1(n3357), .A2(n4227), .ZN(n4219) );
  NAND2_X1 U3766 ( .A1(n5050), .A2(n4301), .ZN(n4471) );
  NOR2_X2 U3767 ( .A1(n6560), .A2(STATE_REG_2__SCAN_IN), .ZN(n6514) );
  AND2_X4 U3768 ( .A1(n4070), .A2(n4067), .ZN(n3207) );
  NAND2_X1 U3769 ( .A1(n5932), .A2(n5142), .ZN(n5141) );
  NAND2_X1 U3770 ( .A1(n4006), .A2(n3956), .ZN(n5468) );
  AOI22_X1 U3771 ( .A1(n3282), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3228), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3103) );
  AND2_X1 U3772 ( .A1(n3006), .A2(n5437), .ZN(n5438) );
  NAND2_X1 U3773 ( .A1(n5098), .A2(n3032), .ZN(n5161) );
  INV_X1 U3774 ( .A(n5305), .ZN(n5611) );
  AOI22_X1 U3775 ( .A1(n3281), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3074) );
  AOI21_X1 U3776 ( .B1(n5439), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5374), 
        .ZN(n5376) );
  XNOR2_X1 U3777 ( .A(n3267), .B(n3266), .ZN(n4233) );
  OR2_X1 U3778 ( .A1(n3168), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3020)
         );
  OR3_X1 U3779 ( .A1(n5462), .A2(REIP_REG_31__SCAN_IN), .A3(n6519), .ZN(n3021)
         );
  OR2_X1 U3780 ( .A1(n5462), .A2(REIP_REG_30__SCAN_IN), .ZN(n3022) );
  AND2_X1 U3781 ( .A1(n5060), .A2(n6724), .ZN(n3023) );
  AND2_X2 U3782 ( .A1(n4105), .A2(n4458), .ZN(n3228) );
  AND4_X1 U3783 ( .A1(n3132), .A2(n3131), .A3(n3130), .A4(n3129), .ZN(n3024)
         );
  NOR2_X1 U3784 ( .A1(n5645), .A2(n5358), .ZN(n3025) );
  OR2_X1 U3785 ( .A1(n5468), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3026)
         );
  AND2_X1 U3786 ( .A1(n3924), .A2(n4191), .ZN(n3027) );
  INV_X1 U3787 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5375) );
  OR2_X1 U3788 ( .A1(n5346), .A2(n6100), .ZN(n3028) );
  OR2_X1 U3789 ( .A1(n3252), .A2(n3251), .ZN(n3029) );
  OR2_X1 U3790 ( .A1(n5468), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3030)
         );
  AND4_X1 U3791 ( .A1(n3140), .A2(n3139), .A3(n3138), .A4(n3137), .ZN(n3031)
         );
  AND2_X1 U3792 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3032) );
  INV_X1 U3793 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5099) );
  NOR2_X1 U3794 ( .A1(n5352), .A2(n5351), .ZN(n3033) );
  OAI22_X1 U3795 ( .A1(n3881), .A2(n3880), .B1(n3872), .B2(n3882), .ZN(n3877)
         );
  OR2_X1 U3796 ( .A1(n3874), .A2(n4144), .ZN(n3867) );
  OR2_X1 U3797 ( .A1(n3864), .A2(n5055), .ZN(n3882) );
  AND2_X1 U3798 ( .A1(n6406), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3868)
         );
  INV_X1 U3799 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3035) );
  AOI22_X1 U3800 ( .A1(n3136), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3071) );
  OAI211_X1 U3801 ( .C1(n3484), .C2(n4308), .A(n3163), .B(n3900), .ZN(n4057)
         );
  AOI22_X1 U3802 ( .A1(n3207), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3053) );
  AND2_X1 U3803 ( .A1(n3189), .A2(n3188), .ZN(n3190) );
  INV_X1 U3804 ( .A(n4266), .ZN(n4259) );
  OAI21_X1 U3805 ( .B1(n3890), .B2(n4027), .A(n3889), .ZN(n3891) );
  NAND2_X1 U3806 ( .A1(n3142), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3316) );
  OR2_X1 U3807 ( .A1(n5163), .A2(n5360), .ZN(n5363) );
  OR2_X1 U3808 ( .A1(n3855), .A2(n3854), .ZN(n4032) );
  AND2_X1 U3809 ( .A1(n5204), .A2(n5060), .ZN(n3932) );
  NAND2_X1 U3810 ( .A1(n4112), .A2(n3160), .ZN(n3939) );
  AND4_X1 U3811 ( .A1(n3094), .A2(n3093), .A3(n3092), .A4(n3091), .ZN(n3095)
         );
  INV_X1 U3812 ( .A(n3244), .ZN(n3555) );
  NAND2_X1 U3813 ( .A1(n3393), .A2(n3392), .ZN(n4743) );
  AND2_X1 U3814 ( .A1(n5769), .A2(n5367), .ZN(n5364) );
  INV_X1 U3815 ( .A(n3932), .ZN(n3991) );
  XNOR2_X1 U3816 ( .A(n3380), .B(n3378), .ZN(n4273) );
  INV_X1 U3817 ( .A(n4025), .ZN(n4026) );
  INV_X1 U3818 ( .A(n5610), .ZN(n3693) );
  MUX2_X1 U3819 ( .A(n3991), .B(n4006), .S(EBX_REG_2__SCAN_IN), .Z(n3923) );
  OR2_X1 U3820 ( .A1(n3764), .A2(n5583), .ZN(n3765) );
  AND2_X1 U3821 ( .A1(n5138), .A2(n3590), .ZN(n5123) );
  AOI21_X1 U3822 ( .B1(n4743), .B2(n3567), .A(n3399), .ZN(n4364) );
  NAND2_X1 U3823 ( .A1(n5607), .A2(n5367), .ZN(n5638) );
  AND2_X1 U3824 ( .A1(n5361), .A2(n5668), .ZN(n5648) );
  NOR2_X1 U3825 ( .A1(n5107), .A2(n5106), .ZN(n3953) );
  AND2_X1 U3826 ( .A1(n3936), .A2(n3935), .ZN(n4367) );
  BUF_X1 U3827 ( .A(n4233), .Z(n4292) );
  AND2_X1 U3828 ( .A1(n4302), .A2(n4301), .ZN(n4340) );
  INV_X1 U3829 ( .A(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n5151) );
  AND2_X1 U3830 ( .A1(n3180), .A2(n3155), .ZN(n5055) );
  INV_X1 U3831 ( .A(n5292), .ZN(n3966) );
  OR2_X1 U3832 ( .A1(n3765), .A2(n5575), .ZN(n3787) );
  NOR2_X1 U3833 ( .A1(n6019), .A2(n3506), .ZN(n3502) );
  NOR2_X1 U3834 ( .A1(n3556), .A2(n5166), .ZN(n3536) );
  INV_X1 U3835 ( .A(n4843), .ZN(n3439) );
  OR2_X1 U3836 ( .A1(n5607), .A2(n5769), .ZN(n5594) );
  CLKBUF_X1 U3837 ( .A(n4771), .Z(n4778) );
  OR2_X1 U3838 ( .A1(n4173), .A2(n4172), .ZN(n6217) );
  OR2_X1 U3839 ( .A1(n6424), .A2(n4464), .ZN(n4466) );
  NAND2_X1 U3840 ( .A1(n3314), .A2(n3313), .ZN(n4547) );
  INV_X1 U3841 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4946) );
  NAND2_X1 U3842 ( .A1(n3642), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3688)
         );
  AND2_X1 U3843 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n3606), .ZN(n3607)
         );
  OR2_X1 U3844 ( .A1(n6549), .A2(n5054), .ZN(n5329) );
  INV_X1 U3845 ( .A(n6078), .ZN(n6097) );
  INV_X1 U3846 ( .A(n6118), .ZN(n3906) );
  INV_X1 U3847 ( .A(n5546), .ZN(n6563) );
  INV_X1 U3848 ( .A(n5829), .ZN(n5874) );
  INV_X1 U3849 ( .A(n4206), .ZN(n6168) );
  INV_X1 U3850 ( .A(n4051), .ZN(n4115) );
  OR2_X1 U3851 ( .A1(n5175), .A2(n5174), .ZN(n5288) );
  INV_X1 U3852 ( .A(n6210), .ZN(n6177) );
  NAND2_X1 U3853 ( .A1(n3395), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3419)
         );
  NOR2_X1 U3854 ( .A1(n4507), .A2(n4506), .ZN(n6421) );
  NAND2_X1 U3855 ( .A1(n5595), .A2(n5594), .ZN(n5632) );
  AND2_X1 U3856 ( .A1(n5091), .A2(n5050), .ZN(n6260) );
  INV_X1 U3857 ( .A(n4471), .ZN(n4612) );
  NOR2_X1 U3858 ( .A1(n3149), .A2(n4506), .ZN(n5407) );
  INV_X1 U3859 ( .A(n4344), .ZN(n4926) );
  NOR2_X1 U3860 ( .A1(n4893), .A2(n4892), .ZN(n4989) );
  INV_X1 U3861 ( .A(n6313), .ZN(n6359) );
  INV_X1 U3862 ( .A(n4617), .ZN(n4810) );
  INV_X1 U3863 ( .A(n4477), .ZN(n6386) );
  INV_X1 U3864 ( .A(n4969), .ZN(n6311) );
  INV_X1 U3865 ( .A(n4973), .ZN(n6345) );
  INV_X1 U3866 ( .A(n4140), .ZN(n4892) );
  INV_X1 U3867 ( .A(n4664), .ZN(n4695) );
  NOR2_X1 U3868 ( .A1(n4519), .A2(n4947), .ZN(n4669) );
  INV_X1 U3869 ( .A(n3003), .ZN(n6065) );
  INV_X1 U3870 ( .A(n6086), .ZN(n6100) );
  AND2_X1 U3871 ( .A1(n5059), .A2(n6038), .ZN(n6105) );
  AND2_X1 U3872 ( .A1(n6566), .A2(n6565), .ZN(n6757) );
  NAND2_X1 U3873 ( .A1(n6123), .A2(n5433), .ZN(n5546) );
  INV_X1 U3874 ( .A(n5380), .ZN(n5550) );
  NAND2_X1 U3875 ( .A1(n4207), .A2(n4206), .ZN(n5432) );
  NAND2_X1 U3876 ( .A1(n5432), .A2(n4209), .ZN(n5867) );
  OR2_X1 U3877 ( .A1(n6162), .A2(n6552), .ZN(n6145) );
  INV_X1 U3878 ( .A(n6162), .ZN(n6166) );
  NAND2_X1 U3879 ( .A1(n4115), .A2(n4144), .ZN(n4374) );
  NAND2_X1 U3880 ( .A1(n4115), .A2(n4113), .ZN(n4206) );
  OR2_X1 U3881 ( .A1(n5126), .A2(n5190), .ZN(n5656) );
  OR2_X1 U3882 ( .A1(n6199), .A2(n4721), .ZN(n6210) );
  AND2_X1 U3883 ( .A1(n5383), .A2(n4835), .ZN(n6251) );
  OR2_X1 U3884 ( .A1(n4173), .A2(n4160), .ZN(n5906) );
  INV_X1 U3885 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6406) );
  AND2_X1 U3886 ( .A1(n4298), .A2(n4297), .ZN(n4349) );
  NAND2_X1 U3887 ( .A1(n4590), .A2(n4892), .ZN(n5257) );
  INV_X1 U3888 ( .A(n6369), .ZN(n4579) );
  OR2_X1 U3889 ( .A1(n4784), .A2(n4140), .ZN(n4887) );
  OR2_X1 U3890 ( .A1(n4786), .A2(n4947), .ZN(n6395) );
  NOR2_X1 U3891 ( .A1(n4476), .A2(n4475), .ZN(n4504) );
  OR2_X1 U3892 ( .A1(n4518), .A2(n4892), .ZN(n4664) );
  NAND2_X1 U3893 ( .A1(n4024), .A2(n4023), .ZN(U2829) );
  INV_X1 U3894 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3034) );
  AND2_X4 U3895 ( .A1(n3034), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4070)
         );
  NOR2_X4 U3896 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4105) );
  AND2_X2 U3897 ( .A1(n4070), .A2(n4105), .ZN(n3125) );
  AND2_X4 U3898 ( .A1(n3256), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3041)
         );
  NOR2_X4 U3899 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3042) );
  AOI22_X1 U3900 ( .A1(n3125), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3040) );
  INV_X1 U3901 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3036) );
  AND2_X2 U3902 ( .A1(n3036), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4109)
         );
  AND2_X2 U3903 ( .A1(n4068), .A2(n4109), .ZN(n3136) );
  AOI22_X1 U3904 ( .A1(n3136), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3017), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3039) );
  AND2_X4 U3905 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4067) );
  AND2_X2 U3906 ( .A1(n3042), .A2(n4105), .ZN(n3135) );
  AOI22_X1 U3907 ( .A1(n3281), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3038) );
  AND2_X4 U3908 ( .A1(n3041), .A2(n4068), .ZN(n3282) );
  AND2_X2 U3909 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4458) );
  AOI22_X1 U3910 ( .A1(n3282), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3228), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3037) );
  AND2_X4 U3911 ( .A1(n3041), .A2(n4458), .ZN(n3280) );
  AOI22_X1 U3912 ( .A1(n3133), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3046) );
  AND2_X2 U3913 ( .A1(n4109), .A2(n3042), .ZN(n3134) );
  AOI22_X1 U3914 ( .A1(n3134), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3016), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3045) );
  AND2_X2 U3915 ( .A1(n4068), .A2(n4105), .ZN(n3126) );
  AND2_X4 U3916 ( .A1(n3042), .A2(n4067), .ZN(n3208) );
  AOI22_X1 U3917 ( .A1(n3126), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3044) );
  AOI22_X1 U3918 ( .A1(n3128), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3223), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3043) );
  INV_X2 U3919 ( .A(n3157), .ZN(n3120) );
  AOI22_X1 U3920 ( .A1(n3134), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3052) );
  AOI22_X1 U3921 ( .A1(n3136), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3051) );
  AOI22_X1 U3922 ( .A1(n3281), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3050) );
  AOI22_X1 U3923 ( .A1(n3282), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3228), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3049) );
  AOI22_X1 U3924 ( .A1(n3127), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3223), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3055) );
  AOI22_X1 U3925 ( .A1(n3017), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3125), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3054) );
  NAND2_X2 U3926 ( .A1(n3120), .A2(n3161), .ZN(n3900) );
  AOI22_X1 U3927 ( .A1(n3134), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3062) );
  AOI22_X1 U3928 ( .A1(n3281), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3061) );
  AOI22_X1 U3929 ( .A1(n3136), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3060) );
  AOI22_X1 U3930 ( .A1(n3282), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3228), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3059) );
  AOI22_X1 U3931 ( .A1(n3017), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3125), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3066) );
  AOI22_X1 U3932 ( .A1(n3128), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3126), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3065) );
  AOI22_X1 U3933 ( .A1(n3207), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3064) );
  AOI22_X1 U3934 ( .A1(n3127), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3223), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3063) );
  AOI22_X1 U3935 ( .A1(n3128), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3017), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3072) );
  AOI22_X1 U3936 ( .A1(n3282), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3070) );
  AOI22_X1 U3937 ( .A1(n3280), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3228), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3069) );
  AOI22_X1 U3938 ( .A1(n3126), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3125), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3076) );
  AOI22_X1 U3939 ( .A1(n3134), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3075) );
  NAND2_X1 U3940 ( .A1(n3136), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3082) );
  NAND2_X1 U3941 ( .A1(n3134), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3081) );
  NAND2_X1 U3942 ( .A1(n3279), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3080)
         );
  NAND2_X1 U3943 ( .A1(n3280), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3079)
         );
  NAND2_X1 U3944 ( .A1(n3207), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3086) );
  NAND2_X1 U3945 ( .A1(n3017), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3085) );
  NAND2_X1 U3946 ( .A1(n3125), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3084) );
  NAND2_X1 U3947 ( .A1(n3208), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3083) );
  NAND2_X1 U3948 ( .A1(n3126), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3090) );
  NAND2_X1 U3949 ( .A1(n3128), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3089) );
  NAND2_X1 U3950 ( .A1(n3127), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3088) );
  NAND2_X1 U3951 ( .A1(n3223), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3087)
         );
  NAND2_X1 U3952 ( .A1(n3281), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3094)
         );
  NAND2_X1 U3953 ( .A1(n3282), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3093)
         );
  NAND2_X1 U3954 ( .A1(n3135), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3092) );
  NAND2_X1 U3955 ( .A1(n3228), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3091)
         );
  AOI22_X1 U3956 ( .A1(n3128), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3126), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3102) );
  AOI22_X1 U3957 ( .A1(n3017), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3125), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3101) );
  AOI22_X1 U3958 ( .A1(n3207), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3100) );
  AOI22_X1 U3959 ( .A1(n3127), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3223), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3099) );
  NAND4_X1 U3960 ( .A1(n3102), .A2(n3101), .A3(n3100), .A4(n3099), .ZN(n3108)
         );
  AOI22_X1 U3961 ( .A1(n3134), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3105) );
  AOI22_X1 U3962 ( .A1(n3281), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3104) );
  NAND4_X1 U3963 ( .A1(n3106), .A2(n3105), .A3(n3104), .A4(n3103), .ZN(n3107)
         );
  NAND2_X1 U3964 ( .A1(n3156), .A2(n3182), .ZN(n3119) );
  NAND2_X1 U3965 ( .A1(n3142), .A2(n3157), .ZN(n3152) );
  AOI22_X1 U3966 ( .A1(n3126), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3125), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3112) );
  AOI22_X1 U3967 ( .A1(n3127), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3223), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3111) );
  AOI22_X1 U3968 ( .A1(n3280), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3207), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3110) );
  AOI22_X1 U3969 ( .A1(n3281), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n3109) );
  NAND4_X1 U3970 ( .A1(n3112), .A2(n3111), .A3(n3110), .A4(n3109), .ZN(n3118)
         );
  AOI22_X1 U3971 ( .A1(n3128), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3017), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3116) );
  AOI22_X1 U3972 ( .A1(n3136), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3115) );
  AOI22_X1 U3973 ( .A1(n3135), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3228), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3114) );
  AOI22_X1 U3974 ( .A1(n3134), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3113) );
  NAND4_X1 U3975 ( .A1(n3116), .A2(n3115), .A3(n3114), .A4(n3113), .ZN(n3117)
         );
  OR2_X2 U3976 ( .A1(n3118), .A2(n3117), .ZN(n3160) );
  OR2_X2 U3977 ( .A1(n3152), .A2(n3939), .ZN(n4162) );
  INV_X1 U3978 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6462) );
  XNOR2_X1 U3979 ( .A(n6462), .B(STATE_REG_2__SCAN_IN), .ZN(n4048) );
  OAI21_X1 U3980 ( .B1(n4048), .B2(n4112), .A(n3120), .ZN(n3121) );
  AND2_X1 U3981 ( .A1(n3484), .A2(n3153), .ZN(n3122) );
  NAND2_X1 U3982 ( .A1(n3122), .A2(n3156), .ZN(n4088) );
  INV_X2 U3983 ( .A(n3142), .ZN(n4308) );
  INV_X1 U3984 ( .A(n4057), .ZN(n3124) );
  NAND2_X1 U3985 ( .A1(n3124), .A2(n3160), .ZN(n3186) );
  AOI22_X1 U3986 ( .A1(n3281), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3282), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3132) );
  AOI22_X1 U3987 ( .A1(n3126), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3125), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3131) );
  AOI22_X1 U3988 ( .A1(n3128), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3130) );
  AOI22_X1 U3989 ( .A1(n3280), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3228), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3129) );
  AOI22_X1 U3990 ( .A1(n3134), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3133), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3140) );
  AOI22_X1 U3991 ( .A1(n3136), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3135), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3139) );
  AOI22_X1 U3992 ( .A1(n3207), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3208), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3138) );
  AOI22_X1 U3993 ( .A1(n3017), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3223), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3137) );
  INV_X2 U3994 ( .A(n4146), .ZN(n4319) );
  MUX2_X1 U3995 ( .A(n3142), .B(n4146), .S(n3161), .Z(n3141) );
  NAND2_X1 U3996 ( .A1(n3141), .A2(n3900), .ZN(n3146) );
  NAND2_X1 U3997 ( .A1(n3900), .A2(n3142), .ZN(n3143) );
  NAND2_X1 U3998 ( .A1(n3143), .A2(n4319), .ZN(n3145) );
  NAND3_X1 U3999 ( .A1(n3146), .A2(n3145), .A3(n3144), .ZN(n3154) );
  NAND2_X1 U4000 ( .A1(n3154), .A2(n5055), .ZN(n3177) );
  NAND3_X1 U4001 ( .A1(n3147), .A2(n4037), .A3(n3177), .ZN(n3148) );
  AND2_X2 U4002 ( .A1(n3148), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3272) );
  INV_X1 U4003 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n3149) );
  NAND2_X1 U4004 ( .A1(n6532), .A2(n3149), .ZN(n6539) );
  NOR2_X1 U4005 ( .A1(n6539), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4509) );
  XNOR2_X1 U4006 ( .A(n6406), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6305)
         );
  NAND2_X1 U4007 ( .A1(n4509), .A2(n6305), .ZN(n3151) );
  AND2_X1 U4008 ( .A1(n6532), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3904) );
  INV_X1 U4009 ( .A(n3904), .ZN(n3276) );
  NAND2_X1 U4010 ( .A1(n3276), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3150) );
  NAND2_X1 U4011 ( .A1(n3151), .A2(n3150), .ZN(n3168) );
  NOR2_X2 U4012 ( .A1(n3154), .A2(n3018), .ZN(n4025) );
  NAND2_X1 U4013 ( .A1(n4025), .A2(n4144), .ZN(n4063) );
  INV_X1 U4014 ( .A(n3156), .ZN(n3159) );
  NOR2_X1 U4015 ( .A1(n4236), .A2(n4329), .ZN(n3158) );
  NOR2_X2 U4016 ( .A1(n4064), .A2(n4164), .ZN(n4040) );
  NAND2_X1 U4017 ( .A1(n4040), .A2(n4112), .ZN(n4081) );
  NAND2_X1 U4018 ( .A1(n4063), .A2(n4081), .ZN(n4157) );
  INV_X1 U4019 ( .A(n4040), .ZN(n4034) );
  INV_X1 U4020 ( .A(n4048), .ZN(n3164) );
  NAND3_X1 U4021 ( .A1(n3901), .A2(n5055), .A3(n3120), .ZN(n4065) );
  NAND2_X1 U4022 ( .A1(n3162), .A2(n3163), .ZN(n5156) );
  OR2_X2 U4023 ( .A1(n4065), .A2(n5156), .ZN(n4170) );
  NAND2_X1 U4024 ( .A1(n3166), .A2(n3167), .ZN(n3268) );
  INV_X1 U4025 ( .A(n3167), .ZN(n3169) );
  NAND2_X1 U4026 ( .A1(n3169), .A2(n3020), .ZN(n3170) );
  NAND2_X1 U4027 ( .A1(n3272), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3173) );
  MUX2_X1 U4028 ( .A(n3276), .B(n4509), .S(n6406), .Z(n3171) );
  INV_X1 U4029 ( .A(n3171), .ZN(n3172) );
  NAND2_X1 U4030 ( .A1(n3173), .A2(n3172), .ZN(n3221) );
  INV_X1 U4031 ( .A(n3484), .ZN(n3174) );
  INV_X1 U4032 ( .A(n4055), .ZN(n5069) );
  AND2_X1 U4033 ( .A1(n3152), .A2(n5069), .ZN(n3175) );
  NOR2_X1 U4034 ( .A1(n4089), .A2(n3175), .ZN(n3176) );
  AND2_X1 U4035 ( .A1(n3177), .A2(n3176), .ZN(n4062) );
  INV_X1 U4036 ( .A(n3178), .ZN(n3185) );
  AND4_X1 U4037 ( .A1(n3179), .A2(n3180), .A3(n4308), .A4(n3163), .ZN(n3181)
         );
  NAND2_X1 U4038 ( .A1(n3181), .A2(n3901), .ZN(n4450) );
  OR2_X1 U4039 ( .A1(n6539), .A2(n5050), .ZN(n6444) );
  AOI21_X1 U4040 ( .B1(n4319), .B2(n3153), .A(n6444), .ZN(n3183) );
  NAND2_X1 U4041 ( .A1(n3182), .A2(n3907), .ZN(n3993) );
  NAND3_X1 U4042 ( .A1(n4450), .A2(n3183), .A3(n3993), .ZN(n3184) );
  NOR2_X1 U4043 ( .A1(n3185), .A2(n3184), .ZN(n3189) );
  AND2_X1 U4044 ( .A1(n3484), .A2(n4308), .ZN(n3187) );
  OAI21_X1 U4045 ( .B1(n3843), .B2(n3187), .A(n4112), .ZN(n3188) );
  NAND2_X1 U4046 ( .A1(n4062), .A2(n3190), .ZN(n3219) );
  AND2_X2 U4047 ( .A1(n3221), .A2(n3219), .ZN(n3270) );
  NAND2_X1 U4048 ( .A1(n4103), .A2(n5050), .ZN(n3263) );
  AOI22_X1 U4049 ( .A1(n3748), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3279), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3194) );
  AOI22_X1 U4050 ( .A1(n3824), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3127), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3193) );
  AOI22_X1 U4051 ( .A1(n3280), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3192) );
  BUF_X1 U4052 ( .A(n3208), .Z(n3229) );
  AOI22_X1 U4053 ( .A1(n3794), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3191) );
  NAND4_X1 U4054 ( .A1(n3194), .A2(n3193), .A3(n3192), .A4(n3191), .ZN(n3201)
         );
  BUF_X1 U4055 ( .A(n3282), .Z(n3195) );
  AOI22_X1 U4056 ( .A1(n3004), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3199) );
  AOI22_X1 U4057 ( .A1(n3207), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3125), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3198) );
  BUF_X1 U4058 ( .A(n3228), .Z(n3771) );
  AOI22_X1 U4059 ( .A1(n3134), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3197) );
  AOI22_X1 U4060 ( .A1(n3128), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3196) );
  NAND4_X1 U4061 ( .A1(n3199), .A2(n3198), .A3(n3197), .A4(n3196), .ZN(n3200)
         );
  INV_X1 U4062 ( .A(n4248), .ZN(n3202) );
  OR2_X1 U4063 ( .A1(n3316), .A2(n3202), .ZN(n3260) );
  INV_X1 U4064 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4328) );
  OR2_X1 U4065 ( .A1(n3856), .A2(n4328), .ZN(n3217) );
  OR2_X1 U4066 ( .A1(n3315), .A2(n3202), .ZN(n3216) );
  AOI22_X1 U4067 ( .A1(n3815), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3279), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3206) );
  AOI22_X1 U4068 ( .A1(n3748), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3280), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3205) );
  AOI22_X1 U4069 ( .A1(n3004), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3204) );
  AOI22_X1 U4070 ( .A1(n3222), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3203) );
  NAND4_X1 U4071 ( .A1(n3206), .A2(n3205), .A3(n3204), .A4(n3203), .ZN(n3214)
         );
  AOI22_X1 U4072 ( .A1(n3128), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3212) );
  AOI22_X1 U4073 ( .A1(n3017), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3211) );
  AOI22_X1 U4074 ( .A1(n3207), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3210) );
  AOI22_X1 U4075 ( .A1(n3127), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3209) );
  NAND4_X1 U4076 ( .A1(n3212), .A2(n3211), .A3(n3210), .A4(n3209), .ZN(n3213)
         );
  OR2_X1 U4077 ( .A1(n3316), .A2(n4823), .ZN(n3215) );
  XNOR2_X2 U4078 ( .A(n3218), .B(n3259), .ZN(n3267) );
  INV_X1 U4079 ( .A(n3219), .ZN(n3220) );
  XNOR2_X1 U4080 ( .A(n3221), .B(n3220), .ZN(n3254) );
  NAND2_X1 U4081 ( .A1(n3254), .A2(n5050), .ZN(n3249) );
  NAND2_X1 U4082 ( .A1(n3142), .A2(n4823), .ZN(n3242) );
  INV_X1 U4083 ( .A(n4823), .ZN(n3404) );
  NAND2_X1 U4084 ( .A1(n3142), .A2(n3404), .ZN(n3236) );
  AOI22_X1 U4085 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n3279), .B1(n3280), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3227) );
  AOI22_X1 U4086 ( .A1(n3134), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3125), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3226) );
  AOI22_X1 U4087 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3222), .B1(n3816), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3225) );
  AOI22_X1 U4088 ( .A1(n3824), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3224) );
  NAND4_X1 U4089 ( .A1(n3227), .A2(n3226), .A3(n3225), .A4(n3224), .ZN(n3235)
         );
  AOI22_X1 U4090 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n3748), .B1(n3207), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3233) );
  AOI22_X1 U4091 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n3128), .B1(n3127), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3232) );
  AOI22_X1 U4092 ( .A1(n3004), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3231) );
  AOI22_X1 U4093 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n3017), .B1(n3229), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3230) );
  NAND4_X1 U4094 ( .A1(n3233), .A2(n3232), .A3(n3231), .A4(n3230), .ZN(n3234)
         );
  MUX2_X1 U4095 ( .A(n3242), .B(n3236), .S(n4247), .Z(n3237) );
  INV_X1 U4096 ( .A(n3237), .ZN(n3238) );
  NAND2_X1 U4097 ( .A1(n3238), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3252) );
  NAND2_X1 U4098 ( .A1(n3249), .A2(n3252), .ZN(n3243) );
  AOI21_X1 U4099 ( .B1(n4164), .B2(n4247), .A(n5050), .ZN(n3239) );
  AND2_X1 U4100 ( .A1(n3239), .A2(n3242), .ZN(n3241) );
  INV_X1 U4101 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4307) );
  OR2_X1 U4102 ( .A1(n3856), .A2(n4307), .ZN(n3240) );
  NAND2_X1 U4103 ( .A1(n3241), .A2(n3240), .ZN(n3251) );
  NOR2_X1 U4104 ( .A1(n3242), .A2(n5050), .ZN(n4817) );
  INV_X2 U4105 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6433) );
  NOR2_X2 U4106 ( .A1(n3162), .A2(n6433), .ZN(n3567) );
  NAND2_X1 U4107 ( .A1(n4292), .A2(n3567), .ZN(n3248) );
  NOR2_X1 U4108 ( .A1(n5156), .A2(n6433), .ZN(n3299) );
  NAND2_X1 U4109 ( .A1(n3299), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3246) );
  NOR2_X1 U4110 ( .A1(n3163), .A2(n6433), .ZN(n3244) );
  AOI22_X1 U4111 ( .A1(n5424), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6433), .ZN(n3245) );
  AND2_X1 U4112 ( .A1(n3246), .A2(n3245), .ZN(n3247) );
  AOI21_X1 U4113 ( .B1(n4892), .B2(n3179), .A(n6433), .ZN(n4225) );
  OR2_X1 U4114 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n3810) );
  INV_X1 U4115 ( .A(n3810), .ZN(n5051) );
  INV_X1 U4116 ( .A(n3299), .ZN(n3354) );
  AOI22_X1 U4117 ( .A1(n5424), .A2(EAX_REG_0__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n6433), .ZN(n3257) );
  OAI21_X1 U4118 ( .B1(n3256), .B2(n3354), .A(n3257), .ZN(n3258) );
  AOI21_X1 U4119 ( .B1(n3255), .B2(n3567), .A(n3258), .ZN(n4226) );
  MUX2_X1 U4120 ( .A(n4225), .B(n5051), .S(n4226), .Z(n4213) );
  AND2_X2 U4121 ( .A1(n4214), .A2(n4213), .ZN(n4216) );
  INV_X1 U4122 ( .A(n3259), .ZN(n3262) );
  INV_X1 U4123 ( .A(n3260), .ZN(n3261) );
  NOR2_X1 U4124 ( .A1(n3262), .A2(n3261), .ZN(n3264) );
  INV_X1 U4125 ( .A(n3306), .ZN(n3297) );
  OAI21_X2 U4126 ( .B1(n3271), .B2(n3270), .A(n3269), .ZN(n3309) );
  AND2_X1 U4127 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3273) );
  NAND2_X1 U4128 ( .A1(n3273), .A2(n4946), .ZN(n4995) );
  INV_X1 U4129 ( .A(n3273), .ZN(n3274) );
  NAND2_X1 U4130 ( .A1(n3274), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3275) );
  NAND2_X1 U4131 ( .A1(n4995), .A2(n3275), .ZN(n4300) );
  AOI22_X1 U4132 ( .A1(n4509), .A2(n4300), .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n3276), .ZN(n3277) );
  XNOR2_X1 U4133 ( .A(n3309), .B(n3307), .ZN(n4295) );
  BUF_X1 U4134 ( .A(n3279), .Z(n3825) );
  AOI22_X1 U4135 ( .A1(n3815), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3286) );
  AOI22_X1 U4136 ( .A1(n3748), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3285) );
  AOI22_X1 U4137 ( .A1(n3004), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3284) );
  AOI22_X1 U4138 ( .A1(n3195), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3283) );
  NAND4_X1 U4139 ( .A1(n3286), .A2(n3285), .A3(n3284), .A4(n3283), .ZN(n3293)
         );
  AOI22_X1 U4140 ( .A1(n3813), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3291) );
  AOI22_X1 U4141 ( .A1(n3794), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3290) );
  AOI22_X1 U4142 ( .A1(n3207), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3289) );
  AOI22_X1 U4143 ( .A1(n3817), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3288) );
  NAND4_X1 U4144 ( .A1(n3291), .A2(n3290), .A3(n3289), .A4(n3288), .ZN(n3292)
         );
  NOR2_X1 U4145 ( .A1(n3316), .A2(n4257), .ZN(n3294) );
  INV_X1 U4146 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4323) );
  OAI22_X1 U4147 ( .A1(n3856), .A2(n4323), .B1(n3315), .B2(n4257), .ZN(n3295)
         );
  NAND2_X1 U4148 ( .A1(n4253), .A2(n3567), .ZN(n3298) );
  NAND2_X1 U4149 ( .A1(n6433), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3372) );
  NAND2_X1 U4150 ( .A1(n3298), .A2(n3372), .ZN(n4187) );
  NAND2_X1 U4151 ( .A1(n4216), .A2(n4187), .ZN(n3304) );
  NAND2_X1 U4152 ( .A1(n3299), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3303) );
  INV_X1 U4153 ( .A(PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5330) );
  OAI21_X1 U4154 ( .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_1__SCAN_IN), .A(n3350), .ZN(n6209) );
  NAND2_X1 U4155 ( .A1(n5051), .A2(n6209), .ZN(n3300) );
  OAI21_X1 U4156 ( .B1(n5330), .B2(n3372), .A(n3300), .ZN(n3301) );
  AOI21_X1 U4157 ( .B1(n5424), .B2(EAX_REG_2__SCAN_IN), .A(n3301), .ZN(n3302)
         );
  AND2_X1 U4158 ( .A1(n3303), .A2(n3302), .ZN(n4185) );
  NAND2_X1 U4159 ( .A1(n3014), .A2(n3305), .ZN(n3347) );
  INV_X1 U4160 ( .A(n3347), .ZN(n3330) );
  INV_X1 U4161 ( .A(n3307), .ZN(n3308) );
  NAND2_X1 U4162 ( .A1(n3272), .A2(n4073), .ZN(n3314) );
  INV_X1 U4163 ( .A(n4509), .ZN(n3311) );
  AND3_X1 U4164 ( .A1(n6718), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6310) );
  NAND2_X1 U4165 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6310), .ZN(n6365) );
  NAND2_X1 U4166 ( .A1(n6718), .A2(n6365), .ZN(n3310) );
  NOR3_X1 U4167 ( .A1(n6718), .A2(n4946), .A3(n4787), .ZN(n4662) );
  NAND2_X1 U4168 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4662), .ZN(n4440) );
  NAND2_X1 U4169 ( .A1(n3310), .A2(n4440), .ZN(n4470) );
  OAI22_X1 U4170 ( .A1(n3311), .A2(n4470), .B1(n3904), .B2(n6718), .ZN(n3312)
         );
  INV_X1 U4171 ( .A(n3312), .ZN(n3313) );
  NAND2_X1 U4172 ( .A1(n4054), .A2(n5050), .ZN(n3329) );
  AOI22_X1 U4173 ( .A1(n3748), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3320) );
  AOI22_X1 U4174 ( .A1(n3195), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4175 ( .A1(n3207), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4176 ( .A1(n3817), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3317) );
  NAND4_X1 U4177 ( .A1(n3320), .A2(n3319), .A3(n3318), .A4(n3317), .ZN(n3326)
         );
  AOI22_X1 U4178 ( .A1(n3813), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3324) );
  AOI22_X1 U4179 ( .A1(n3794), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3323) );
  AOI22_X1 U4180 ( .A1(n3004), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3322) );
  AOI22_X1 U4181 ( .A1(n3815), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3321) );
  NAND4_X1 U4182 ( .A1(n3324), .A2(n3323), .A3(n3322), .A4(n3321), .ZN(n3325)
         );
  INV_X1 U4183 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4318) );
  OAI22_X1 U4184 ( .A1(n3874), .A2(n4259), .B1(n4318), .B2(n3856), .ZN(n3327)
         );
  INV_X1 U4185 ( .A(n3327), .ZN(n3328) );
  NAND2_X1 U4186 ( .A1(n3330), .A2(n4545), .ZN(n3358) );
  AOI22_X1 U4187 ( .A1(n3815), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4188 ( .A1(n3748), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3333) );
  AOI22_X1 U4189 ( .A1(n3004), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3332) );
  AOI22_X1 U4190 ( .A1(n3195), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3331) );
  NAND4_X1 U4191 ( .A1(n3334), .A2(n3333), .A3(n3332), .A4(n3331), .ZN(n3340)
         );
  AOI22_X1 U4192 ( .A1(n3813), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4193 ( .A1(n3794), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3337) );
  AOI22_X1 U4194 ( .A1(n3207), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4195 ( .A1(n3817), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3335) );
  NAND4_X1 U4196 ( .A1(n3338), .A2(n3337), .A3(n3336), .A4(n3335), .ZN(n3339)
         );
  INV_X1 U4197 ( .A(n4744), .ZN(n3341) );
  INV_X1 U4198 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4313) );
  OAI22_X1 U4199 ( .A1(n3874), .A2(n3341), .B1(n4313), .B2(n3856), .ZN(n3359)
         );
  XNOR2_X1 U4200 ( .A(n3358), .B(n3359), .ZN(n4265) );
  NAND2_X1 U4201 ( .A1(n4265), .A2(n3567), .ZN(n3346) );
  INV_X1 U4202 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4203 ( .A1(n5424), .A2(EAX_REG_4__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n6433), .ZN(n3342) );
  OAI21_X1 U4204 ( .B1(n3851), .B2(n3354), .A(n3342), .ZN(n3344) );
  OAI21_X1 U4205 ( .B1(n3349), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n3394), 
        .ZN(n6198) );
  AND2_X1 U4206 ( .A1(n6198), .A2(n5051), .ZN(n3343) );
  AOI21_X1 U4207 ( .B1(n3344), .B2(n3810), .A(n3343), .ZN(n3345) );
  NAND2_X1 U4208 ( .A1(n3346), .A2(n3345), .ZN(n4230) );
  XNOR2_X1 U4209 ( .A(n3347), .B(n4545), .ZN(n4256) );
  INV_X1 U4210 ( .A(n4073), .ZN(n4101) );
  AOI21_X1 U4211 ( .B1(n3351), .B2(n3350), .A(n3349), .ZN(n6109) );
  OAI22_X1 U4212 ( .A1(n6109), .A2(n3810), .B1(n3372), .B2(n3351), .ZN(n3352)
         );
  AOI21_X1 U4213 ( .B1(n5424), .B2(EAX_REG_3__SCAN_IN), .A(n3352), .ZN(n3353)
         );
  OAI21_X1 U4214 ( .B1(n3354), .B2(n4101), .A(n3353), .ZN(n3355) );
  AOI21_X1 U4215 ( .B1(n3348), .B2(n3567), .A(n3355), .ZN(n4229) );
  INV_X1 U4216 ( .A(n4229), .ZN(n3356) );
  INV_X1 U4217 ( .A(n3358), .ZN(n3360) );
  AOI22_X1 U4218 ( .A1(n3815), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4219 ( .A1(n3813), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4220 ( .A1(n3794), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4221 ( .A1(n3817), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3361) );
  NAND4_X1 U4222 ( .A1(n3364), .A2(n3363), .A3(n3362), .A4(n3361), .ZN(n3370)
         );
  AOI22_X1 U4223 ( .A1(n3748), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4224 ( .A1(n3004), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4225 ( .A1(n3195), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4226 ( .A1(n3814), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3365) );
  NAND4_X1 U4227 ( .A1(n3368), .A2(n3367), .A3(n3366), .A4(n3365), .ZN(n3369)
         );
  INV_X1 U4228 ( .A(n4745), .ZN(n3371) );
  INV_X1 U4229 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4334) );
  OAI22_X1 U4230 ( .A1(n3874), .A2(n3371), .B1(n4334), .B2(n3856), .ZN(n3378)
         );
  XOR2_X1 U4231 ( .A(n5117), .B(n3394), .Z(n5114) );
  NAND2_X1 U4232 ( .A1(n3244), .A2(EAX_REG_5__SCAN_IN), .ZN(n3374) );
  INV_X1 U4233 ( .A(n3372), .ZN(n5423) );
  NAND2_X1 U4234 ( .A1(n5423), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3373)
         );
  OAI211_X1 U4235 ( .C1(n5114), .C2(n3810), .A(n3374), .B(n3373), .ZN(n3375)
         );
  NAND2_X1 U4236 ( .A1(n3377), .A2(n3376), .ZN(n4218) );
  INV_X1 U4237 ( .A(n3378), .ZN(n3379) );
  INV_X1 U4238 ( .A(n3403), .ZN(n3393) );
  AOI22_X1 U4239 ( .A1(n3815), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3384) );
  AOI22_X1 U4240 ( .A1(n3748), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3383) );
  AOI22_X1 U4241 ( .A1(n3004), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4242 ( .A1(n3195), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3381) );
  NAND4_X1 U4243 ( .A1(n3384), .A2(n3383), .A3(n3382), .A4(n3381), .ZN(n3390)
         );
  AOI22_X1 U4244 ( .A1(n3813), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3388) );
  AOI22_X1 U4245 ( .A1(n3794), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U4246 ( .A1(n3814), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4247 ( .A1(n3817), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3385) );
  NAND4_X1 U4248 ( .A1(n3388), .A2(n3387), .A3(n3386), .A4(n3385), .ZN(n3389)
         );
  OR2_X1 U4249 ( .A1(n3390), .A2(n3389), .ZN(n4756) );
  INV_X1 U4250 ( .A(n4756), .ZN(n3391) );
  INV_X1 U4251 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4338) );
  OAI22_X1 U4252 ( .A1(n3874), .A2(n3391), .B1(n3856), .B2(n4338), .ZN(n3402)
         );
  INV_X1 U4253 ( .A(n3402), .ZN(n3392) );
  OAI21_X1 U4254 ( .B1(n3395), .B2(PHYADDRPOINTER_REG_6__SCAN_IN), .A(n3419), 
        .ZN(n6190) );
  INV_X1 U4255 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3397) );
  INV_X1 U4256 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3396) );
  OAI22_X1 U4257 ( .A1(n3555), .A2(n3397), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n3396), .ZN(n3398) );
  MUX2_X1 U4258 ( .A(n6190), .B(n3398), .S(n3810), .Z(n3399) );
  INV_X1 U4259 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4348) );
  OAI22_X1 U4260 ( .A1(n3874), .A2(n3404), .B1(n4348), .B2(n3856), .ZN(n3405)
         );
  XOR2_X1 U4261 ( .A(n5151), .B(n3419), .Z(n4763) );
  NAND2_X1 U4262 ( .A1(n5423), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3407)
         );
  NAND2_X1 U4263 ( .A1(n3244), .A2(EAX_REG_7__SCAN_IN), .ZN(n3406) );
  OAI211_X1 U4264 ( .C1(n4763), .C2(n3810), .A(n3407), .B(n3406), .ZN(n3408)
         );
  NOR2_X2 U4265 ( .A1(n4646), .A2(n4647), .ZN(n4769) );
  AOI22_X1 U4266 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3195), .B1(n3815), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3412) );
  AOI22_X1 U4267 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n3824), .B1(n3814), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3411) );
  AOI22_X1 U4268 ( .A1(n3004), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3410) );
  AOI22_X1 U4269 ( .A1(n3817), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3409) );
  NAND4_X1 U4270 ( .A1(n3412), .A2(n3411), .A3(n3410), .A4(n3409), .ZN(n3418)
         );
  AOI22_X1 U4271 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3748), .B1(n3825), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4272 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n3813), .B1(n3823), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3415) );
  AOI22_X1 U4273 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n3822), .B1(n3771), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3414) );
  AOI22_X1 U4274 ( .A1(n3794), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3413) );
  NAND4_X1 U4275 ( .A1(n3416), .A2(n3415), .A3(n3414), .A4(n3413), .ZN(n3417)
         );
  NOR2_X1 U4276 ( .A1(n3418), .A2(n3417), .ZN(n3422) );
  INV_X1 U4277 ( .A(n3567), .ZN(n3472) );
  XNOR2_X1 U4278 ( .A(n3423), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6058) );
  NAND2_X1 U4279 ( .A1(n6058), .A2(n5051), .ZN(n3421) );
  AOI22_X1 U4280 ( .A1(n5424), .A2(EAX_REG_8__SCAN_IN), .B1(n5423), .B2(
        PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3420) );
  OAI211_X1 U4281 ( .C1(n3422), .C2(n3472), .A(n3421), .B(n3420), .ZN(n4768)
         );
  NAND2_X1 U4282 ( .A1(n4769), .A2(n4768), .ZN(n4767) );
  INV_X1 U4283 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n6043) );
  NAND2_X1 U4284 ( .A1(PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n3423), .ZN(n3440)
         );
  XOR2_X1 U4285 ( .A(n6043), .B(n3440), .Z(n6046) );
  INV_X1 U4286 ( .A(n6046), .ZN(n3438) );
  AOI22_X1 U4287 ( .A1(n3748), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3427) );
  AOI22_X1 U4288 ( .A1(n3813), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4289 ( .A1(n3195), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4290 ( .A1(n3815), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3424) );
  NAND4_X1 U4291 ( .A1(n3427), .A2(n3426), .A3(n3425), .A4(n3424), .ZN(n3433)
         );
  AOI22_X1 U4292 ( .A1(n3822), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3814), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3431) );
  AOI22_X1 U4293 ( .A1(n3824), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3430) );
  AOI22_X1 U4294 ( .A1(n3004), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4295 ( .A1(n3817), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3428) );
  NAND4_X1 U4296 ( .A1(n3431), .A2(n3430), .A3(n3429), .A4(n3428), .ZN(n3432)
         );
  OAI21_X1 U4297 ( .B1(n3433), .B2(n3432), .A(n3567), .ZN(n3436) );
  NAND2_X1 U4298 ( .A1(n3244), .A2(EAX_REG_9__SCAN_IN), .ZN(n3435) );
  NAND2_X1 U4299 ( .A1(n5423), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3434)
         );
  NAND3_X1 U4300 ( .A1(n3436), .A2(n3435), .A3(n3434), .ZN(n3437) );
  AOI21_X1 U4301 ( .B1(n3438), .B2(n5051), .A(n3437), .ZN(n4843) );
  INV_X1 U4302 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n6690) );
  NAND2_X1 U4303 ( .A1(n3441), .A2(n6690), .ZN(n3443) );
  INV_X1 U4304 ( .A(n3489), .ZN(n3442) );
  NAND2_X1 U4305 ( .A1(n3443), .A2(n3442), .ZN(n6037) );
  AOI22_X1 U4306 ( .A1(n3748), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3447) );
  AOI22_X1 U4307 ( .A1(n3815), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3814), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3446) );
  AOI22_X1 U4308 ( .A1(n3824), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3445) );
  AOI22_X1 U4309 ( .A1(n3817), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3444) );
  NAND4_X1 U4310 ( .A1(n3447), .A2(n3446), .A3(n3445), .A4(n3444), .ZN(n3453)
         );
  AOI22_X1 U4311 ( .A1(n3825), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4312 ( .A1(n3813), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4313 ( .A1(n3004), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3449) );
  AOI22_X1 U4314 ( .A1(n3195), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3448) );
  NAND4_X1 U4315 ( .A1(n3451), .A2(n3450), .A3(n3449), .A4(n3448), .ZN(n3452)
         );
  OAI21_X1 U4316 ( .B1(n3453), .B2(n3452), .A(n3567), .ZN(n3456) );
  NAND2_X1 U4317 ( .A1(n3244), .A2(EAX_REG_10__SCAN_IN), .ZN(n3455) );
  NAND2_X1 U4318 ( .A1(n5423), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3454)
         );
  NAND3_X1 U4319 ( .A1(n3456), .A2(n3455), .A3(n3454), .ZN(n3457) );
  AOI21_X1 U4320 ( .B1(n6037), .B2(n5051), .A(n3457), .ZN(n4938) );
  AOI22_X1 U4321 ( .A1(n3748), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3461) );
  AOI22_X1 U4322 ( .A1(n3815), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3460) );
  AOI22_X1 U4323 ( .A1(n3824), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3459) );
  AOI22_X1 U4324 ( .A1(n3004), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3458) );
  NAND4_X1 U4325 ( .A1(n3461), .A2(n3460), .A3(n3459), .A4(n3458), .ZN(n3467)
         );
  AOI22_X1 U4326 ( .A1(n3279), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3814), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3465) );
  AOI22_X1 U4327 ( .A1(n3822), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4328 ( .A1(n3794), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3463) );
  AOI22_X1 U4329 ( .A1(n3813), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3462) );
  NAND4_X1 U4330 ( .A1(n3465), .A2(n3464), .A3(n3463), .A4(n3462), .ZN(n3466)
         );
  NOR2_X1 U4331 ( .A1(n3467), .A2(n3466), .ZN(n3471) );
  XOR2_X1 U4332 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n3489), .Z(n6176) );
  INV_X1 U4333 ( .A(n6176), .ZN(n3468) );
  AOI22_X1 U4334 ( .A1(n5423), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .B1(n5051), 
        .B2(n3468), .ZN(n3470) );
  NAND2_X1 U4335 ( .A1(n3244), .A2(EAX_REG_11__SCAN_IN), .ZN(n3469) );
  OAI211_X1 U4336 ( .C1(n3472), .C2(n3471), .A(n3470), .B(n3469), .ZN(n5038)
         );
  AOI22_X1 U4337 ( .A1(n3748), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3476) );
  AOI22_X1 U4338 ( .A1(n3195), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3475) );
  AOI22_X1 U4339 ( .A1(n3814), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3474) );
  AOI22_X1 U4340 ( .A1(n3825), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3473) );
  NAND4_X1 U4341 ( .A1(n3476), .A2(n3475), .A3(n3474), .A4(n3473), .ZN(n3486)
         );
  AOI22_X1 U4342 ( .A1(n3004), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3482) );
  AOI22_X1 U4343 ( .A1(n3823), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3481) );
  NAND2_X1 U4344 ( .A1(n3822), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3478) );
  NAND2_X1 U4345 ( .A1(n3776), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3477) );
  AND3_X1 U4346 ( .A1(n3478), .A2(n3810), .A3(n3477), .ZN(n3480) );
  AOI22_X1 U4347 ( .A1(n3813), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3479) );
  NAND4_X1 U4348 ( .A1(n3482), .A2(n3481), .A3(n3480), .A4(n3479), .ZN(n3485)
         );
  NAND2_X1 U4349 ( .A1(n4308), .A2(n3163), .ZN(n3483) );
  OR2_X1 U4350 ( .A1(n3484), .A2(n3483), .ZN(n4038) );
  NOR2_X1 U4351 ( .A1(n4038), .A2(n4319), .ZN(n6401) );
  NAND2_X1 U4352 ( .A1(n6401), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3834) );
  NAND2_X1 U4353 ( .A1(n3834), .A2(n3810), .ZN(n3657) );
  OAI21_X1 U4354 ( .B1(n3486), .B2(n3485), .A(n3657), .ZN(n3488) );
  AOI22_X1 U4355 ( .A1(n5424), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6433), .ZN(n3487) );
  NAND2_X1 U4356 ( .A1(n3488), .A2(n3487), .ZN(n3491) );
  INV_X1 U4357 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n6019) );
  INV_X1 U4358 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5166) );
  NAND2_X1 U4359 ( .A1(n3536), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3521)
         );
  INV_X1 U4360 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n5295) );
  XNOR2_X1 U4361 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n3605), .ZN(n5653)
         );
  NAND2_X1 U4362 ( .A1(n5051), .A2(n5653), .ZN(n3490) );
  NAND2_X1 U4363 ( .A1(n3491), .A2(n3490), .ZN(n5124) );
  INV_X1 U4364 ( .A(n5124), .ZN(n3591) );
  AOI22_X1 U4365 ( .A1(n3195), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3495) );
  AOI22_X1 U4366 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n3825), .B1(n3815), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3494) );
  AOI22_X1 U4367 ( .A1(n3813), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3493) );
  AOI22_X1 U4368 ( .A1(n3004), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3492) );
  NAND4_X1 U4369 ( .A1(n3495), .A2(n3494), .A3(n3493), .A4(n3492), .ZN(n3501)
         );
  AOI22_X1 U4370 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n3824), .B1(n3794), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3499) );
  AOI22_X1 U4371 ( .A1(n3748), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3498) );
  AOI22_X1 U4372 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n3814), .B1(n3229), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3497) );
  AOI22_X1 U4373 ( .A1(n3817), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3496) );
  NAND4_X1 U4374 ( .A1(n3499), .A2(n3498), .A3(n3497), .A4(n3496), .ZN(n3500)
         );
  NOR2_X1 U4375 ( .A1(n3501), .A2(n3500), .ZN(n3505) );
  XNOR2_X1 U4376 ( .A(n3502), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6012)
         );
  NAND2_X1 U4377 ( .A1(n6012), .A2(n5051), .ZN(n3504) );
  AOI22_X1 U4378 ( .A1(n5424), .A2(EAX_REG_16__SCAN_IN), .B1(n5423), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3503) );
  OAI211_X1 U4379 ( .C1(n3505), .C2(n3834), .A(n3504), .B(n3503), .ZN(n5140)
         );
  XOR2_X1 U4380 ( .A(n6019), .B(n3506), .Z(n6023) );
  INV_X1 U4381 ( .A(n6023), .ZN(n5675) );
  AOI22_X1 U4382 ( .A1(n3748), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3510) );
  AOI22_X1 U4383 ( .A1(n3815), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3814), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3509) );
  AOI22_X1 U4384 ( .A1(n3824), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3508) );
  AOI22_X1 U4385 ( .A1(n3004), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3507) );
  NAND4_X1 U4386 ( .A1(n3510), .A2(n3509), .A3(n3508), .A4(n3507), .ZN(n3516)
         );
  AOI22_X1 U4387 ( .A1(n3813), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4388 ( .A1(n3822), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4389 ( .A1(n3825), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3512) );
  AOI22_X1 U4390 ( .A1(n3817), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3511) );
  NAND4_X1 U4391 ( .A1(n3514), .A2(n3513), .A3(n3512), .A4(n3511), .ZN(n3515)
         );
  OAI21_X1 U4392 ( .B1(n3516), .B2(n3515), .A(n3567), .ZN(n3519) );
  NAND2_X1 U4393 ( .A1(n5424), .A2(EAX_REG_15__SCAN_IN), .ZN(n3518) );
  NAND2_X1 U4394 ( .A1(n5423), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3517)
         );
  NAND3_X1 U4395 ( .A1(n3519), .A2(n3518), .A3(n3517), .ZN(n3520) );
  AOI21_X1 U4396 ( .B1(n5675), .B2(n5051), .A(n3520), .ZN(n5282) );
  XNOR2_X1 U4397 ( .A(n3521), .B(n5295), .ZN(n5319) );
  AOI22_X1 U4398 ( .A1(n3748), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3815), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3525) );
  AOI22_X1 U4399 ( .A1(n3813), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3524) );
  AOI22_X1 U4400 ( .A1(n3822), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3523) );
  AOI22_X1 U4401 ( .A1(n3817), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3522) );
  NAND4_X1 U4402 ( .A1(n3525), .A2(n3524), .A3(n3523), .A4(n3522), .ZN(n3531)
         );
  AOI22_X1 U4403 ( .A1(n3004), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3529) );
  AOI22_X1 U4404 ( .A1(n3794), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3528) );
  AOI22_X1 U4405 ( .A1(n3825), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3527) );
  AOI22_X1 U4406 ( .A1(n3814), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3526) );
  NAND4_X1 U4407 ( .A1(n3529), .A2(n3528), .A3(n3527), .A4(n3526), .ZN(n3530)
         );
  OAI21_X1 U4408 ( .B1(n3531), .B2(n3530), .A(n3567), .ZN(n3534) );
  NAND2_X1 U4409 ( .A1(n5424), .A2(EAX_REG_14__SCAN_IN), .ZN(n3533) );
  NAND2_X1 U4410 ( .A1(n5423), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3532)
         );
  NAND3_X1 U4411 ( .A1(n3534), .A2(n3533), .A3(n3532), .ZN(n3535) );
  AOI21_X1 U4412 ( .B1(n5319), .B2(n5051), .A(n3535), .ZN(n5289) );
  OR2_X1 U4413 ( .A1(n5282), .A2(n5289), .ZN(n3552) );
  XOR2_X1 U4414 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .B(n3536), .Z(n5277) );
  INV_X1 U4415 ( .A(n5277), .ZN(n3551) );
  AOI22_X1 U4416 ( .A1(n3004), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4417 ( .A1(n3748), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3814), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3539) );
  AOI22_X1 U4418 ( .A1(n3823), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4419 ( .A1(n3817), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3537) );
  NAND4_X1 U4420 ( .A1(n3540), .A2(n3539), .A3(n3538), .A4(n3537), .ZN(n3546)
         );
  AOI22_X1 U4421 ( .A1(n3815), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3544) );
  AOI22_X1 U4422 ( .A1(n3813), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3543) );
  AOI22_X1 U4423 ( .A1(n3825), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4424 ( .A1(n3816), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3541) );
  NAND4_X1 U4425 ( .A1(n3544), .A2(n3543), .A3(n3542), .A4(n3541), .ZN(n3545)
         );
  OAI21_X1 U4426 ( .B1(n3546), .B2(n3545), .A(n3567), .ZN(n3549) );
  NAND2_X1 U4427 ( .A1(n3244), .A2(EAX_REG_13__SCAN_IN), .ZN(n3548) );
  NAND2_X1 U4428 ( .A1(n5423), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n3547)
         );
  NAND3_X1 U4429 ( .A1(n3549), .A2(n3548), .A3(n3547), .ZN(n3550) );
  AOI21_X1 U4430 ( .B1(n3551), .B2(n5051), .A(n3550), .ZN(n5174) );
  NOR2_X1 U4431 ( .A1(n3552), .A2(n5174), .ZN(n5137) );
  AND2_X1 U4432 ( .A1(n5140), .A2(n5137), .ZN(n3572) );
  INV_X1 U4433 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5090) );
  AOI21_X1 U4434 ( .B1(STATEBS16_REG_SCAN_IN), .B2(n5166), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3553) );
  INV_X1 U4435 ( .A(n3553), .ZN(n3554) );
  OAI21_X1 U4436 ( .B1(n3555), .B2(n5090), .A(n3554), .ZN(n3558) );
  XNOR2_X1 U4437 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3556), .ZN(n5168)
         );
  NAND2_X1 U4438 ( .A1(n5051), .A2(n5168), .ZN(n3557) );
  NAND2_X1 U4439 ( .A1(n3558), .A2(n3557), .ZN(n3571) );
  AOI22_X1 U4440 ( .A1(n3815), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4441 ( .A1(n3794), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3814), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4442 ( .A1(n3824), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4443 ( .A1(n3195), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3559) );
  NAND4_X1 U4444 ( .A1(n3562), .A2(n3561), .A3(n3560), .A4(n3559), .ZN(n3569)
         );
  AOI22_X1 U4445 ( .A1(n3748), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3279), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4446 ( .A1(n3004), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4447 ( .A1(n3823), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4448 ( .A1(n3813), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3563) );
  NAND4_X1 U4449 ( .A1(n3566), .A2(n3565), .A3(n3564), .A4(n3563), .ZN(n3568)
         );
  OAI21_X1 U4450 ( .B1(n3569), .B2(n3568), .A(n3567), .ZN(n3570) );
  NAND2_X1 U4451 ( .A1(n3571), .A2(n3570), .ZN(n5081) );
  AND2_X1 U4452 ( .A1(n3572), .A2(n5081), .ZN(n5138) );
  AOI22_X1 U4453 ( .A1(n3748), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3576) );
  AOI22_X1 U4454 ( .A1(n3824), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3575) );
  AOI22_X1 U4455 ( .A1(n3195), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3574) );
  AOI22_X1 U4456 ( .A1(n3817), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3573) );
  NAND4_X1 U4457 ( .A1(n3576), .A2(n3575), .A3(n3574), .A4(n3573), .ZN(n3582)
         );
  AOI22_X1 U4458 ( .A1(n3279), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3580) );
  AOI22_X1 U4459 ( .A1(n3815), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3814), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3579) );
  AOI22_X1 U4460 ( .A1(n3004), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3578) );
  AOI22_X1 U4461 ( .A1(n3813), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3577) );
  NAND4_X1 U4462 ( .A1(n3580), .A2(n3579), .A3(n3578), .A4(n3577), .ZN(n3581)
         );
  NOR2_X1 U4463 ( .A1(n3582), .A2(n3581), .ZN(n3586) );
  INV_X1 U4464 ( .A(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3583) );
  OAI21_X1 U4465 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n3583), .A(n3810), .ZN(
        n3584) );
  AOI21_X1 U4466 ( .B1(n3244), .B2(EAX_REG_17__SCAN_IN), .A(n3584), .ZN(n3585)
         );
  OAI21_X1 U4467 ( .B1(n3834), .B2(n3586), .A(n3585), .ZN(n3589) );
  OAI21_X1 U4468 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3587), .A(n3605), 
        .ZN(n6003) );
  OR2_X1 U4469 ( .A1(n3810), .A2(n6003), .ZN(n3588) );
  NAND2_X1 U4470 ( .A1(n3589), .A2(n3588), .ZN(n5899) );
  INV_X1 U4471 ( .A(n5899), .ZN(n3590) );
  AND2_X1 U4472 ( .A1(n3591), .A2(n5123), .ZN(n5125) );
  AOI22_X1 U4473 ( .A1(n3748), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3595) );
  AOI22_X1 U4474 ( .A1(n3815), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3279), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3594) );
  AOI22_X1 U4475 ( .A1(n3814), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3593) );
  AOI22_X1 U4476 ( .A1(n3004), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3592) );
  NAND4_X1 U4477 ( .A1(n3595), .A2(n3594), .A3(n3593), .A4(n3592), .ZN(n3601)
         );
  AOI22_X1 U4478 ( .A1(n3813), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3599) );
  AOI22_X1 U4479 ( .A1(n3822), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3598) );
  AOI22_X1 U4480 ( .A1(n3794), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4481 ( .A1(n3817), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3596) );
  NAND4_X1 U4482 ( .A1(n3599), .A2(n3598), .A3(n3597), .A4(n3596), .ZN(n3600)
         );
  NOR2_X1 U4483 ( .A1(n3601), .A2(n3600), .ZN(n3602) );
  OR2_X1 U4484 ( .A1(n3834), .A2(n3602), .ZN(n3610) );
  NAND2_X1 U4485 ( .A1(n6433), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n3603)
         );
  NAND2_X1 U4486 ( .A1(n3810), .A2(n3603), .ZN(n3604) );
  AOI21_X1 U4487 ( .B1(n3244), .B2(EAX_REG_19__SCAN_IN), .A(n3604), .ZN(n3609)
         );
  OAI21_X1 U4488 ( .B1(n3607), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n3641), 
        .ZN(n5862) );
  NOR2_X1 U4489 ( .A1(n5862), .A2(n3810), .ZN(n3608) );
  AOI21_X1 U4490 ( .B1(n3610), .B2(n3609), .A(n3608), .ZN(n5189) );
  AND2_X1 U4491 ( .A1(n5125), .A2(n5189), .ZN(n3611) );
  AOI22_X1 U4492 ( .A1(n3815), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3813), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3617) );
  NAND2_X1 U4493 ( .A1(n3748), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3613)
         );
  NAND2_X1 U4494 ( .A1(n3817), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3612) );
  AND3_X1 U4495 ( .A1(n3613), .A2(n3612), .A3(n3810), .ZN(n3616) );
  AOI22_X1 U4496 ( .A1(n3004), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3615) );
  AOI22_X1 U4497 ( .A1(n3814), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3614) );
  NAND4_X1 U4498 ( .A1(n3617), .A2(n3616), .A3(n3615), .A4(n3614), .ZN(n3623)
         );
  AOI22_X1 U4499 ( .A1(n3825), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3621) );
  AOI22_X1 U4500 ( .A1(n3824), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3620) );
  AOI22_X1 U4501 ( .A1(n3222), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3619) );
  AOI22_X1 U4502 ( .A1(n3794), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3618) );
  NAND4_X1 U4503 ( .A1(n3621), .A2(n3620), .A3(n3619), .A4(n3618), .ZN(n3622)
         );
  OR2_X1 U4504 ( .A1(n3623), .A2(n3622), .ZN(n3624) );
  NAND2_X1 U4505 ( .A1(n3657), .A2(n3624), .ZN(n3627) );
  AOI22_X1 U4506 ( .A1(n5424), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6433), .ZN(n3626) );
  XNOR2_X1 U4507 ( .A(n3641), .B(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5636)
         );
  AND2_X1 U4508 ( .A1(n5636), .A2(n5051), .ZN(n3625) );
  AOI21_X1 U4509 ( .B1(n3627), .B2(n3626), .A(n3625), .ZN(n5202) );
  AOI22_X1 U4510 ( .A1(n3748), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3631) );
  AOI22_X1 U4511 ( .A1(n3825), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3814), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3630) );
  AOI22_X1 U4512 ( .A1(n3794), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3629) );
  AOI22_X1 U4513 ( .A1(n3824), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3628) );
  NAND4_X1 U4514 ( .A1(n3631), .A2(n3630), .A3(n3629), .A4(n3628), .ZN(n3637)
         );
  AOI22_X1 U4515 ( .A1(n3813), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3635) );
  AOI22_X1 U4516 ( .A1(n3004), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3634) );
  AOI22_X1 U4517 ( .A1(n3822), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3633) );
  AOI22_X1 U4518 ( .A1(n3815), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3632) );
  NAND4_X1 U4519 ( .A1(n3635), .A2(n3634), .A3(n3633), .A4(n3632), .ZN(n3636)
         );
  NOR2_X1 U4520 ( .A1(n3637), .A2(n3636), .ZN(n3638) );
  OR2_X1 U4521 ( .A1(n3834), .A2(n3638), .ZN(n3646) );
  INV_X1 U4522 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6743) );
  OAI21_X1 U4523 ( .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n6743), .A(n6433), 
        .ZN(n3639) );
  INV_X1 U4524 ( .A(n3639), .ZN(n3640) );
  AOI21_X1 U4525 ( .B1(n3244), .B2(EAX_REG_21__SCAN_IN), .A(n3640), .ZN(n3645)
         );
  INV_X1 U4526 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5633) );
  OR2_X1 U4527 ( .A1(n3642), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n3643)
         );
  NAND2_X1 U4528 ( .A1(n3688), .A2(n3643), .ZN(n5852) );
  NOR2_X1 U4529 ( .A1(n5852), .A2(n3810), .ZN(n3644) );
  AOI21_X1 U4530 ( .B1(n3646), .B2(n3645), .A(n3644), .ZN(n5264) );
  AOI22_X1 U4531 ( .A1(n3815), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3650) );
  AOI22_X1 U4532 ( .A1(n3195), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3813), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3649) );
  AOI22_X1 U4533 ( .A1(n3823), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3648) );
  AOI22_X1 U4534 ( .A1(n3794), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3647) );
  NAND4_X1 U4535 ( .A1(n3650), .A2(n3649), .A3(n3648), .A4(n3647), .ZN(n3659)
         );
  AOI22_X1 U4536 ( .A1(n3748), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3656) );
  AOI22_X1 U4537 ( .A1(n3814), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3655) );
  NAND2_X1 U4538 ( .A1(n3280), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3652) );
  NAND2_X1 U4539 ( .A1(n3776), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3651) );
  AND3_X1 U4540 ( .A1(n3652), .A2(n3810), .A3(n3651), .ZN(n3654) );
  AOI22_X1 U4541 ( .A1(n3825), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3653) );
  NAND4_X1 U4542 ( .A1(n3656), .A2(n3655), .A3(n3654), .A4(n3653), .ZN(n3658)
         );
  OAI21_X1 U4543 ( .B1(n3659), .B2(n3658), .A(n3657), .ZN(n3662) );
  INV_X1 U4544 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5838) );
  NOR2_X1 U4545 ( .A1(n5838), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3660) );
  AOI21_X1 U4546 ( .B1(n3244), .B2(EAX_REG_22__SCAN_IN), .A(n3660), .ZN(n3661)
         );
  NAND2_X1 U4547 ( .A1(n3662), .A2(n3661), .ZN(n3664) );
  XNOR2_X1 U4548 ( .A(n3688), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5835)
         );
  NAND2_X1 U4549 ( .A1(n5835), .A2(n5051), .ZN(n3663) );
  NAND2_X1 U4550 ( .A1(n3664), .A2(n3663), .ZN(n5306) );
  NOR2_X2 U4551 ( .A1(n5263), .A2(n5306), .ZN(n5305) );
  AOI22_X1 U4552 ( .A1(n3004), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3668) );
  AOI22_X1 U4553 ( .A1(n3748), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3667) );
  AOI22_X1 U4554 ( .A1(n3825), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3666) );
  AOI22_X1 U4555 ( .A1(n3824), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3665) );
  NAND4_X1 U4556 ( .A1(n3668), .A2(n3667), .A3(n3666), .A4(n3665), .ZN(n3674)
         );
  AOI22_X1 U4557 ( .A1(n3815), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3814), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3672) );
  AOI22_X1 U4558 ( .A1(n3816), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3671) );
  AOI22_X1 U4559 ( .A1(n3794), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3670) );
  AOI22_X1 U4560 ( .A1(n3813), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3669) );
  NAND4_X1 U4561 ( .A1(n3672), .A2(n3671), .A3(n3670), .A4(n3669), .ZN(n3673)
         );
  NOR2_X1 U4562 ( .A1(n3674), .A2(n3673), .ZN(n3694) );
  AOI22_X1 U4563 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n3825), .B1(n3822), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3678) );
  AOI22_X1 U4564 ( .A1(n3815), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3814), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3677) );
  AOI22_X1 U4565 ( .A1(n3823), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3676) );
  AOI22_X1 U4566 ( .A1(n3813), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3675) );
  NAND4_X1 U4567 ( .A1(n3678), .A2(n3677), .A3(n3676), .A4(n3675), .ZN(n3684)
         );
  AOI22_X1 U4568 ( .A1(n3748), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3682) );
  AOI22_X1 U4569 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n3824), .B1(n3817), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3681) );
  AOI22_X1 U4570 ( .A1(n3004), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3680) );
  AOI22_X1 U4571 ( .A1(n3222), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3679) );
  NAND4_X1 U4572 ( .A1(n3682), .A2(n3681), .A3(n3680), .A4(n3679), .ZN(n3683)
         );
  NOR2_X1 U4573 ( .A1(n3684), .A2(n3683), .ZN(n3695) );
  XNOR2_X1 U4574 ( .A(n3694), .B(n3695), .ZN(n3687) );
  INV_X1 U4575 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5609) );
  OAI21_X1 U4576 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5609), .A(n3810), .ZN(
        n3685) );
  AOI21_X1 U4577 ( .B1(n3244), .B2(EAX_REG_23__SCAN_IN), .A(n3685), .ZN(n3686)
         );
  OAI21_X1 U4578 ( .B1(n3834), .B2(n3687), .A(n3686), .ZN(n3692) );
  AND2_X1 U4579 ( .A1(n3689), .A2(n5609), .ZN(n3690) );
  OR2_X1 U4580 ( .A1(n3690), .A2(n3725), .ZN(n5826) );
  INV_X1 U4581 ( .A(n5826), .ZN(n5616) );
  NAND2_X1 U4582 ( .A1(n5616), .A2(n5051), .ZN(n3691) );
  NAND2_X1 U4583 ( .A1(n3692), .A2(n3691), .ZN(n5610) );
  AND2_X2 U4584 ( .A1(n5305), .A2(n3693), .ZN(n5612) );
  OR2_X1 U4585 ( .A1(n3695), .A2(n3694), .ZN(n3711) );
  AOI22_X1 U4586 ( .A1(n3824), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3699) );
  AOI22_X1 U4587 ( .A1(n3222), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3698) );
  AOI22_X1 U4588 ( .A1(n3823), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3697) );
  AOI22_X1 U4589 ( .A1(n3816), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3696) );
  NAND4_X1 U4590 ( .A1(n3699), .A2(n3698), .A3(n3697), .A4(n3696), .ZN(n3705)
         );
  AOI22_X1 U4591 ( .A1(n3815), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3813), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3703) );
  AOI22_X1 U4592 ( .A1(n3748), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3004), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3702) );
  AOI22_X1 U4593 ( .A1(n3822), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3701) );
  AOI22_X1 U4594 ( .A1(n3814), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3700) );
  NAND4_X1 U4595 ( .A1(n3703), .A2(n3702), .A3(n3701), .A4(n3700), .ZN(n3704)
         );
  NOR2_X1 U4596 ( .A1(n3705), .A2(n3704), .ZN(n3710) );
  XNOR2_X1 U4597 ( .A(n3711), .B(n3710), .ZN(n3709) );
  AOI22_X1 U4598 ( .A1(n5424), .A2(EAX_REG_24__SCAN_IN), .B1(n5423), .B2(
        PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n3707) );
  XNOR2_X1 U4599 ( .A(n3725), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5813)
         );
  NAND2_X1 U4600 ( .A1(n5813), .A2(n5051), .ZN(n3706) );
  AND2_X1 U4601 ( .A1(n3707), .A2(n3706), .ZN(n3708) );
  OAI21_X1 U4602 ( .B1(n3834), .B2(n3709), .A(n3708), .ZN(n5539) );
  AND2_X2 U4603 ( .A1(n5612), .A2(n5539), .ZN(n5540) );
  NOR2_X1 U4604 ( .A1(n3711), .A2(n3710), .ZN(n3730) );
  AOI22_X1 U4605 ( .A1(n3748), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3715) );
  AOI22_X1 U4606 ( .A1(n3824), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3714) );
  AOI22_X1 U4607 ( .A1(n3825), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3814), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3713) );
  AOI22_X1 U4608 ( .A1(n3817), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3712) );
  NAND4_X1 U4609 ( .A1(n3715), .A2(n3714), .A3(n3713), .A4(n3712), .ZN(n3721)
         );
  AOI22_X1 U4610 ( .A1(n3813), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3719) );
  AOI22_X1 U4611 ( .A1(n3004), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3718) );
  AOI22_X1 U4612 ( .A1(n3822), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3717) );
  AOI22_X1 U4613 ( .A1(n3815), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3716) );
  NAND4_X1 U4614 ( .A1(n3719), .A2(n3718), .A3(n3717), .A4(n3716), .ZN(n3720)
         );
  OR2_X1 U4615 ( .A1(n3721), .A2(n3720), .ZN(n3731) );
  XNOR2_X1 U4616 ( .A(n3730), .B(n3731), .ZN(n3724) );
  INV_X1 U4617 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5802) );
  AOI21_X1 U4618 ( .B1(n5802), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3722) );
  AOI21_X1 U4619 ( .B1(n5424), .B2(EAX_REG_25__SCAN_IN), .A(n3722), .ZN(n3723)
         );
  OAI21_X1 U4620 ( .B1(n3724), .B2(n3834), .A(n3723), .ZN(n3729) );
  OR2_X1 U4621 ( .A1(n3726), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n3727)
         );
  AND2_X1 U4622 ( .A1(n3764), .A2(n3727), .ZN(n5804) );
  NAND2_X1 U4623 ( .A1(n5804), .A2(n5051), .ZN(n3728) );
  NAND2_X2 U4624 ( .A1(n5540), .A2(n5535), .ZN(n5534) );
  AND2_X1 U4625 ( .A1(n3731), .A2(n3730), .ZN(n3760) );
  AOI22_X1 U4626 ( .A1(n3815), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3735) );
  AOI22_X1 U4627 ( .A1(n3748), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3734) );
  AOI22_X1 U4628 ( .A1(n3004), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3733) );
  AOI22_X1 U4629 ( .A1(n3222), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3732) );
  NAND4_X1 U4630 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n3741)
         );
  AOI22_X1 U4631 ( .A1(n3813), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3739) );
  AOI22_X1 U4632 ( .A1(n3794), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3738) );
  AOI22_X1 U4633 ( .A1(n3814), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3737) );
  AOI22_X1 U4634 ( .A1(n3817), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3736) );
  NAND4_X1 U4635 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3740)
         );
  OR2_X1 U4636 ( .A1(n3741), .A2(n3740), .ZN(n3759) );
  XNOR2_X1 U4637 ( .A(n3760), .B(n3759), .ZN(n3744) );
  INV_X1 U4638 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5583) );
  OAI21_X1 U4639 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5583), .A(n3810), .ZN(
        n3742) );
  AOI21_X1 U4640 ( .B1(n5424), .B2(EAX_REG_26__SCAN_IN), .A(n3742), .ZN(n3743)
         );
  OAI21_X1 U4641 ( .B1(n3744), .B2(n3834), .A(n3743), .ZN(n3746) );
  XNOR2_X1 U4642 ( .A(n3764), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5792)
         );
  NAND2_X1 U4643 ( .A1(n5792), .A2(n5051), .ZN(n3745) );
  NAND2_X1 U4644 ( .A1(n3746), .A2(n3745), .ZN(n5526) );
  NOR2_X2 U4645 ( .A1(n5534), .A2(n5526), .ZN(n3747) );
  INV_X1 U4646 ( .A(n3747), .ZN(n5528) );
  AOI22_X1 U4647 ( .A1(n3004), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3752) );
  AOI22_X1 U4648 ( .A1(n3279), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3814), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3751) );
  AOI22_X1 U4649 ( .A1(n3748), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3750) );
  AOI22_X1 U4650 ( .A1(n3823), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3749) );
  NAND4_X1 U4651 ( .A1(n3752), .A2(n3751), .A3(n3750), .A4(n3749), .ZN(n3758)
         );
  AOI22_X1 U4652 ( .A1(n3813), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3756) );
  AOI22_X1 U4653 ( .A1(n3815), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3755) );
  AOI22_X1 U4654 ( .A1(n3822), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3754) );
  AOI22_X1 U4655 ( .A1(n3817), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3753) );
  NAND4_X1 U4656 ( .A1(n3756), .A2(n3755), .A3(n3754), .A4(n3753), .ZN(n3757)
         );
  NOR2_X1 U4657 ( .A1(n3758), .A2(n3757), .ZN(n3770) );
  NAND2_X1 U4658 ( .A1(n3760), .A2(n3759), .ZN(n3769) );
  XNOR2_X1 U4659 ( .A(n3770), .B(n3769), .ZN(n3763) );
  INV_X1 U4660 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5575) );
  AOI21_X1 U4661 ( .B1(n5575), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3761) );
  AOI21_X1 U4662 ( .B1(n5424), .B2(EAX_REG_27__SCAN_IN), .A(n3761), .ZN(n3762)
         );
  OAI21_X1 U4663 ( .B1(n3763), .B2(n3834), .A(n3762), .ZN(n3768) );
  NAND2_X1 U4664 ( .A1(n3765), .A2(n5575), .ZN(n3766) );
  NAND2_X1 U4665 ( .A1(n3787), .A2(n3766), .ZN(n5785) );
  INV_X1 U4666 ( .A(n5785), .ZN(n5578) );
  NAND2_X1 U4667 ( .A1(n5578), .A2(n5051), .ZN(n3767) );
  NAND2_X1 U4668 ( .A1(n3768), .A2(n3767), .ZN(n5520) );
  XNOR2_X1 U4669 ( .A(n3787), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5566)
         );
  INV_X1 U4670 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5564) );
  OAI21_X1 U4671 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5564), .A(n3810), .ZN(
        n3785) );
  NOR2_X1 U4672 ( .A1(n3770), .A2(n3769), .ZN(n3793) );
  AOI22_X1 U4673 ( .A1(n3815), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3775) );
  AOI22_X1 U4674 ( .A1(n3748), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3774) );
  AOI22_X1 U4675 ( .A1(n3004), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3773) );
  AOI22_X1 U4676 ( .A1(n3222), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3771), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3772) );
  NAND4_X1 U4677 ( .A1(n3775), .A2(n3774), .A3(n3773), .A4(n3772), .ZN(n3782)
         );
  AOI22_X1 U4678 ( .A1(n3813), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3824), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3780) );
  AOI22_X1 U4679 ( .A1(n3794), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U4680 ( .A1(n3814), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3778) );
  AOI22_X1 U4681 ( .A1(n3817), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3777) );
  NAND4_X1 U4682 ( .A1(n3780), .A2(n3779), .A3(n3778), .A4(n3777), .ZN(n3781)
         );
  OR2_X1 U4683 ( .A1(n3782), .A2(n3781), .ZN(n3792) );
  XNOR2_X1 U4684 ( .A(n3793), .B(n3792), .ZN(n3783) );
  NOR2_X1 U4685 ( .A1(n3783), .A2(n3834), .ZN(n3784) );
  AOI211_X1 U4686 ( .C1(n5424), .C2(EAX_REG_28__SCAN_IN), .A(n3785), .B(n3784), 
        .ZN(n3786) );
  AOI21_X1 U4687 ( .B1(n5051), .B2(n5566), .A(n3786), .ZN(n5494) );
  NAND2_X1 U4688 ( .A1(n3788), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5056)
         );
  INV_X1 U4689 ( .A(n3788), .ZN(n3790) );
  INV_X1 U4690 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n3789) );
  NAND2_X1 U4691 ( .A1(n3790), .A2(n3789), .ZN(n3791) );
  NAND2_X1 U4692 ( .A1(n5056), .A2(n3791), .ZN(n5485) );
  NAND2_X1 U4693 ( .A1(n3793), .A2(n3792), .ZN(n3811) );
  AOI22_X1 U4694 ( .A1(n3222), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3825), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U4695 ( .A1(n3824), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3797) );
  AOI22_X1 U4696 ( .A1(n3815), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3814), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3796) );
  AOI22_X1 U4697 ( .A1(n3813), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3795) );
  NAND4_X1 U4698 ( .A1(n3798), .A2(n3797), .A3(n3796), .A4(n3795), .ZN(n3805)
         );
  AOI22_X1 U4699 ( .A1(n3823), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3817), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3803) );
  AOI22_X1 U4700 ( .A1(n3004), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3816), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3802) );
  AOI22_X1 U4701 ( .A1(n3822), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3801) );
  AOI22_X1 U4702 ( .A1(n3748), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3229), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3800) );
  NAND4_X1 U4703 ( .A1(n3803), .A2(n3802), .A3(n3801), .A4(n3800), .ZN(n3804)
         );
  NOR2_X1 U4704 ( .A1(n3805), .A2(n3804), .ZN(n3812) );
  XNOR2_X1 U4705 ( .A(n3811), .B(n3812), .ZN(n3808) );
  NAND2_X1 U4706 ( .A1(n5424), .A2(EAX_REG_29__SCAN_IN), .ZN(n3807) );
  OAI21_X1 U4707 ( .B1(n6743), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n6433), 
        .ZN(n3806) );
  OAI211_X1 U4708 ( .C1(n3808), .C2(n3834), .A(n3807), .B(n3806), .ZN(n3809)
         );
  OAI21_X1 U4709 ( .B1(n3810), .B2(n5485), .A(n3809), .ZN(n5453) );
  NOR2_X1 U4710 ( .A1(n3812), .A2(n3811), .ZN(n3833) );
  AOI22_X1 U4711 ( .A1(n3813), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3794), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3821) );
  AOI22_X1 U4712 ( .A1(n3815), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3814), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3820) );
  AOI22_X1 U4713 ( .A1(n3816), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3799), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3819) );
  AOI22_X1 U4714 ( .A1(n3817), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3776), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3818) );
  NAND4_X1 U4715 ( .A1(n3821), .A2(n3820), .A3(n3819), .A4(n3818), .ZN(n3831)
         );
  AOI22_X1 U4716 ( .A1(n3004), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3222), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4717 ( .A1(n3748), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3822), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3828) );
  AOI22_X1 U4718 ( .A1(n3824), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3823), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4719 ( .A1(n3825), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3287), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3826) );
  NAND4_X1 U4720 ( .A1(n3829), .A2(n3828), .A3(n3827), .A4(n3826), .ZN(n3830)
         );
  NOR2_X1 U4721 ( .A1(n3831), .A2(n3830), .ZN(n3832) );
  XNOR2_X1 U4722 ( .A(n3833), .B(n3832), .ZN(n3836) );
  INV_X1 U4723 ( .A(n3834), .ZN(n3835) );
  NAND2_X1 U4724 ( .A1(n3836), .A2(n3835), .ZN(n3840) );
  INV_X1 U4725 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5350) );
  AOI21_X1 U4726 ( .B1(n5350), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n3837) );
  AOI21_X1 U4727 ( .B1(n5424), .B2(EAX_REG_30__SCAN_IN), .A(n3837), .ZN(n3839)
         );
  XNOR2_X1 U4728 ( .A(n5056), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5349)
         );
  AND2_X1 U4729 ( .A1(n5349), .A2(n5051), .ZN(n3838) );
  AOI21_X1 U4730 ( .B1(n3840), .B2(n3839), .A(n3838), .ZN(n5422) );
  NAND3_X1 U4731 ( .A1(n6401), .A2(n4112), .A3(n4055), .ZN(n3842) );
  OR2_X1 U4732 ( .A1(n3843), .A2(n3842), .ZN(n4161) );
  INV_X1 U4733 ( .A(n4161), .ZN(n3899) );
  NAND2_X1 U4734 ( .A1(n4329), .A2(n4112), .ZN(n4818) );
  NOR2_X1 U4735 ( .A1(n3856), .A2(n4818), .ZN(n3875) );
  XNOR2_X1 U4736 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3865) );
  NAND2_X1 U4737 ( .A1(n3868), .A2(n3865), .ZN(n3845) );
  NAND2_X1 U4738 ( .A1(n4787), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3844) );
  NAND2_X1 U4739 ( .A1(n3845), .A2(n3844), .ZN(n3863) );
  XNOR2_X1 U4740 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3861) );
  NAND2_X1 U4741 ( .A1(n3863), .A2(n3861), .ZN(n3847) );
  NAND2_X1 U4742 ( .A1(n4946), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3846) );
  NAND2_X1 U4743 ( .A1(n3847), .A2(n3846), .ZN(n3860) );
  XNOR2_X1 U4744 ( .A(n4073), .B(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3858)
         );
  NAND2_X1 U4745 ( .A1(n3860), .A2(n3858), .ZN(n3849) );
  NAND2_X1 U4746 ( .A1(n6718), .A2(n4073), .ZN(n3848) );
  NAND2_X1 U4747 ( .A1(n3849), .A2(n3848), .ZN(n3855) );
  INV_X1 U4748 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6293) );
  AND2_X1 U4749 ( .A1(n6293), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3850)
         );
  OR2_X1 U4750 ( .A1(n3855), .A2(n3850), .ZN(n3852) );
  NAND2_X1 U4751 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3851), .ZN(n3854) );
  NAND2_X1 U4752 ( .A1(n3852), .A2(n3854), .ZN(n4031) );
  INV_X1 U4753 ( .A(n4031), .ZN(n3853) );
  NAND2_X1 U4754 ( .A1(n3875), .A2(n3853), .ZN(n3898) );
  OR2_X1 U4755 ( .A1(n3874), .A2(n4031), .ZN(n3896) );
  AOI21_X1 U4756 ( .B1(n3874), .B2(n4753), .A(n4032), .ZN(n3893) );
  INV_X1 U4757 ( .A(n4032), .ZN(n3857) );
  AOI22_X1 U4758 ( .A1(n3857), .A2(n3890), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n5050), .ZN(n3892) );
  INV_X1 U4759 ( .A(n3858), .ZN(n3859) );
  XNOR2_X1 U4760 ( .A(n3860), .B(n3859), .ZN(n4027) );
  INV_X1 U4761 ( .A(n3861), .ZN(n3862) );
  XNOR2_X1 U4762 ( .A(n3863), .B(n3862), .ZN(n4028) );
  INV_X1 U4763 ( .A(n4028), .ZN(n3884) );
  INV_X1 U4764 ( .A(n3883), .ZN(n3888) );
  AND2_X1 U4765 ( .A1(n4144), .A2(n4329), .ZN(n3864) );
  INV_X1 U4766 ( .A(n3882), .ZN(n3887) );
  INV_X1 U4767 ( .A(n3865), .ZN(n3866) );
  XNOR2_X1 U4768 ( .A(n3866), .B(n3868), .ZN(n4029) );
  AND2_X1 U4769 ( .A1(n4029), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3881) );
  NAND2_X1 U4770 ( .A1(n3867), .A2(n4329), .ZN(n3880) );
  AOI21_X1 U4771 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n3256), .A(n3868), 
        .ZN(n3871) );
  INV_X1 U4772 ( .A(n3871), .ZN(n3873) );
  INV_X1 U4773 ( .A(n3869), .ZN(n3870) );
  AOI21_X1 U4774 ( .B1(n3871), .B2(n3152), .A(n3870), .ZN(n3872) );
  NOR3_X1 U4775 ( .A1(n3874), .A2(n3873), .A3(n3877), .ZN(n3879) );
  INV_X1 U4776 ( .A(n3875), .ZN(n3876) );
  AOI21_X1 U4777 ( .B1(n4029), .B2(n3877), .A(n3876), .ZN(n3878) );
  AOI211_X1 U4778 ( .C1(n3881), .C2(n3880), .A(n3879), .B(n3878), .ZN(n3886)
         );
  AOI211_X1 U4779 ( .C1(n3890), .C2(n3884), .A(n3883), .B(n3882), .ZN(n3885)
         );
  OAI222_X1 U4780 ( .A1(n3888), .A2(n3887), .B1(n4818), .B2(n4027), .C1(n3886), 
        .C2(n3885), .ZN(n3889) );
  AOI222_X1 U4781 ( .A1(n3893), .A2(n3892), .B1(n3893), .B2(n3891), .C1(n3892), 
        .C2(n3891), .ZN(n3894) );
  INV_X1 U4782 ( .A(n3894), .ZN(n3895) );
  NAND2_X1 U4783 ( .A1(n3896), .A2(n3895), .ZN(n3897) );
  NAND2_X1 U4784 ( .A1(n3899), .A2(n4506), .ZN(n4094) );
  INV_X1 U4785 ( .A(n3900), .ZN(n3902) );
  NOR2_X1 U4786 ( .A1(n4308), .A2(n3163), .ZN(n4202) );
  NAND4_X1 U4787 ( .A1(n3902), .A2(n3901), .A3(n5060), .A4(n4202), .ZN(n3903)
         );
  NAND2_X1 U4788 ( .A1(n4094), .A2(n3903), .ZN(n3905) );
  AND2_X1 U4789 ( .A1(n3904), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4508) );
  CLKBUF_X3 U4790 ( .A(n3939), .Z(n4009) );
  INV_X1 U4791 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3908) );
  NAND2_X1 U4792 ( .A1(n3932), .A2(n3908), .ZN(n3912) );
  NAND2_X1 U4793 ( .A1(n3907), .A2(n3153), .ZN(n3919) );
  INV_X1 U4794 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4281) );
  NAND2_X1 U4795 ( .A1(n3919), .A2(n4281), .ZN(n3910) );
  NAND2_X1 U4796 ( .A1(n5060), .A2(n3908), .ZN(n3909) );
  NAND3_X1 U4797 ( .A1(n3910), .A2(n3956), .A3(n3909), .ZN(n3911) );
  NAND2_X1 U4798 ( .A1(n3912), .A2(n3911), .ZN(n3916) );
  NAND2_X1 U4799 ( .A1(n3919), .A2(EBX_REG_0__SCAN_IN), .ZN(n3915) );
  INV_X1 U4800 ( .A(EBX_REG_0__SCAN_IN), .ZN(n3913) );
  NAND2_X1 U4801 ( .A1(n3956), .A2(n3913), .ZN(n3914) );
  NAND2_X1 U4802 ( .A1(n3915), .A2(n3914), .ZN(n4174) );
  NAND2_X1 U4805 ( .A1(n5060), .A2(n4009), .ZN(n4001) );
  MUX2_X1 U4806 ( .A(n4001), .B(n4009), .S(EBX_REG_3__SCAN_IN), .Z(n3920) );
  OAI21_X1 U4807 ( .B1(INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n5468), .A(n3920), 
        .ZN(n4359) );
  INV_X1 U4808 ( .A(n4359), .ZN(n3924) );
  NAND2_X1 U4809 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n5467), .ZN(n3921)
         );
  AND2_X1 U4810 ( .A1(n3993), .A2(n3921), .ZN(n3922) );
  MUX2_X1 U4811 ( .A(n3991), .B(n4006), .S(EBX_REG_4__SCAN_IN), .Z(n3928) );
  NAND2_X1 U4812 ( .A1(n5467), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3926)
         );
  AND2_X1 U4813 ( .A1(n3993), .A2(n3926), .ZN(n3927) );
  MUX2_X1 U4814 ( .A(n4001), .B(n3956), .S(EBX_REG_5__SCAN_IN), .Z(n3929) );
  INV_X1 U4815 ( .A(n3929), .ZN(n3931) );
  NOR2_X1 U4816 ( .A1(n5468), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3930)
         );
  NOR2_X1 U4817 ( .A1(n3931), .A2(n3930), .ZN(n4222) );
  INV_X1 U4818 ( .A(EBX_REG_6__SCAN_IN), .ZN(n6066) );
  NAND2_X1 U4819 ( .A1(n4004), .A2(n6066), .ZN(n3936) );
  INV_X1 U4820 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n6256) );
  NAND2_X1 U4821 ( .A1(n4006), .A2(n6256), .ZN(n3934) );
  NAND2_X1 U4822 ( .A1(n5060), .A2(n6066), .ZN(n3933) );
  NAND3_X1 U4823 ( .A1(n3934), .A2(n3956), .A3(n3933), .ZN(n3935) );
  MUX2_X1 U4824 ( .A(n4001), .B(n3956), .S(EBX_REG_7__SCAN_IN), .Z(n3940) );
  NAND2_X1 U4825 ( .A1(n3030), .A2(n3940), .ZN(n4779) );
  NOR2_X2 U4826 ( .A1(n4780), .A2(n4779), .ZN(n4771) );
  INV_X1 U4827 ( .A(EBX_REG_8__SCAN_IN), .ZN(n6056) );
  NAND2_X1 U4828 ( .A1(n4004), .A2(n6056), .ZN(n3944) );
  INV_X1 U4829 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4836) );
  NAND2_X1 U4830 ( .A1(n4006), .A2(n4836), .ZN(n3942) );
  NAND2_X1 U4831 ( .A1(n5060), .A2(n6056), .ZN(n3941) );
  NAND3_X1 U4832 ( .A1(n3942), .A2(n3956), .A3(n3941), .ZN(n3943) );
  NAND2_X1 U4833 ( .A1(n3944), .A2(n3943), .ZN(n4772) );
  AND2_X2 U4834 ( .A1(n4771), .A2(n4772), .ZN(n4848) );
  MUX2_X1 U4835 ( .A(n4001), .B(n4009), .S(EBX_REG_9__SCAN_IN), .Z(n3945) );
  INV_X1 U4836 ( .A(n3945), .ZN(n3947) );
  NOR2_X1 U4837 ( .A1(n5468), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n3946)
         );
  NOR2_X1 U4838 ( .A1(n3947), .A2(n3946), .ZN(n4847) );
  NAND2_X1 U4839 ( .A1(n4848), .A2(n4847), .ZN(n4846) );
  MUX2_X1 U4840 ( .A(n3991), .B(n4006), .S(EBX_REG_10__SCAN_IN), .Z(n3950) );
  NAND2_X1 U4841 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n5467), .ZN(n3948) );
  AND2_X1 U4842 ( .A1(n3993), .A2(n3948), .ZN(n3949) );
  NAND2_X1 U4843 ( .A1(n3950), .A2(n3949), .ZN(n4941) );
  INV_X1 U4844 ( .A(n4941), .ZN(n5107) );
  NAND2_X1 U4845 ( .A1(n3956), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3951) );
  OAI211_X1 U4846 ( .C1(n5467), .C2(EBX_REG_11__SCAN_IN), .A(n4006), .B(n3951), 
        .ZN(n3952) );
  OAI21_X1 U4847 ( .B1(n4001), .B2(EBX_REG_11__SCAN_IN), .A(n3952), .ZN(n5106)
         );
  INV_X1 U4848 ( .A(EBX_REG_12__SCAN_IN), .ZN(n6719) );
  NAND2_X1 U4849 ( .A1(n4004), .A2(n6719), .ZN(n3959) );
  INV_X1 U4850 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6223) );
  NAND2_X1 U4851 ( .A1(n4006), .A2(n6223), .ZN(n3957) );
  NAND2_X1 U4852 ( .A1(n5060), .A2(n6719), .ZN(n3955) );
  NAND3_X1 U4853 ( .A1(n3957), .A2(n3956), .A3(n3955), .ZN(n3958) );
  AND2_X1 U4854 ( .A1(n3959), .A2(n3958), .ZN(n5083) );
  NOR2_X2 U4855 ( .A1(n5109), .A2(n5083), .ZN(n5179) );
  INV_X1 U4856 ( .A(n4001), .ZN(n5444) );
  INV_X1 U4857 ( .A(EBX_REG_13__SCAN_IN), .ZN(n6695) );
  NAND2_X1 U4858 ( .A1(n5444), .A2(n6695), .ZN(n3962) );
  NAND2_X1 U4859 ( .A1(n3956), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3960) );
  OAI211_X1 U4860 ( .C1(n5467), .C2(EBX_REG_13__SCAN_IN), .A(n4006), .B(n3960), 
        .ZN(n3961) );
  AND2_X1 U4861 ( .A1(n3962), .A2(n3961), .ZN(n5178) );
  NAND2_X1 U4862 ( .A1(n5179), .A2(n5178), .ZN(n5293) );
  MUX2_X1 U4863 ( .A(n3991), .B(n4006), .S(EBX_REG_14__SCAN_IN), .Z(n3965) );
  NAND2_X1 U4864 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5467), .ZN(n3963) );
  AND2_X1 U4865 ( .A1(n3993), .A2(n3963), .ZN(n3964) );
  AND2_X1 U4866 ( .A1(n3965), .A2(n3964), .ZN(n5292) );
  NAND2_X1 U4867 ( .A1(n4009), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3968) );
  OAI211_X1 U4868 ( .C1(n5467), .C2(EBX_REG_15__SCAN_IN), .A(n4006), .B(n3968), 
        .ZN(n3969) );
  OAI21_X1 U4869 ( .B1(n4001), .B2(EBX_REG_15__SCAN_IN), .A(n3969), .ZN(n5929)
         );
  NOR2_X2 U4870 ( .A1(n5930), .A2(n5929), .ZN(n5932) );
  MUX2_X1 U4871 ( .A(n3991), .B(n4006), .S(EBX_REG_16__SCAN_IN), .Z(n3972) );
  NAND2_X1 U4872 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n5467), .ZN(n3970) );
  AND2_X1 U4873 ( .A1(n3993), .A2(n3970), .ZN(n3971) );
  NAND2_X1 U4874 ( .A1(n3972), .A2(n3971), .ZN(n5142) );
  NAND2_X1 U4875 ( .A1(n3956), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3973) );
  OAI211_X1 U4876 ( .C1(n5467), .C2(EBX_REG_17__SCAN_IN), .A(n4006), .B(n3973), 
        .ZN(n3974) );
  OAI21_X1 U4877 ( .B1(n4001), .B2(EBX_REG_17__SCAN_IN), .A(n3974), .ZN(n5914)
         );
  OR2_X2 U4878 ( .A1(n5141), .A2(n5914), .ZN(n5916) );
  INV_X1 U4879 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5197) );
  NAND2_X1 U4880 ( .A1(n4004), .A2(n5197), .ZN(n3978) );
  INV_X1 U4881 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U4882 ( .A1(n4006), .A2(n5769), .ZN(n3976) );
  NAND2_X1 U4883 ( .A1(n5060), .A2(n5197), .ZN(n3975) );
  NAND3_X1 U4884 ( .A1(n3976), .A2(n3956), .A3(n3975), .ZN(n3977) );
  AND2_X1 U4885 ( .A1(n3978), .A2(n3977), .ZN(n5193) );
  OR2_X2 U4886 ( .A1(n5916), .A2(n5193), .ZN(n5203) );
  OR2_X1 U4887 ( .A1(n5468), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3979)
         );
  INV_X1 U4888 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U4889 ( .A1(n5060), .A2(n5173), .ZN(n5129) );
  AND2_X1 U4890 ( .A1(n3979), .A2(n5129), .ZN(n5205) );
  OAI22_X1 U4891 ( .A1(n5468), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n5467), .ZN(n5207) );
  NAND2_X1 U4892 ( .A1(n5205), .A2(n5207), .ZN(n3981) );
  NAND2_X1 U4893 ( .A1(n5204), .A2(EBX_REG_20__SCAN_IN), .ZN(n3980) );
  OAI211_X1 U4894 ( .C1(n5205), .C2(n5204), .A(n3981), .B(n3980), .ZN(n3982)
         );
  NOR2_X2 U4895 ( .A1(n5203), .A2(n3982), .ZN(n5266) );
  MUX2_X1 U4896 ( .A(n4001), .B(n3956), .S(EBX_REG_21__SCAN_IN), .Z(n3983) );
  OAI21_X1 U4897 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5468), .A(n3983), 
        .ZN(n5268) );
  INV_X1 U4898 ( .A(n5268), .ZN(n3984) );
  AND2_X2 U4899 ( .A1(n5266), .A2(n3984), .ZN(n5267) );
  MUX2_X1 U4900 ( .A(n3991), .B(n4006), .S(EBX_REG_22__SCAN_IN), .Z(n3987) );
  NAND2_X1 U4901 ( .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n5467), .ZN(n3985) );
  AND2_X1 U4902 ( .A1(n3993), .A2(n3985), .ZN(n3986) );
  NAND2_X1 U4903 ( .A1(n3987), .A2(n3986), .ZN(n5308) );
  AND2_X2 U4904 ( .A1(n5267), .A2(n5308), .ZN(n5730) );
  INV_X1 U4905 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5865) );
  NAND2_X1 U4906 ( .A1(n5444), .A2(n5865), .ZN(n3990) );
  NAND2_X1 U4907 ( .A1(n4009), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3988) );
  OAI211_X1 U4908 ( .C1(n5467), .C2(EBX_REG_23__SCAN_IN), .A(n4006), .B(n3988), 
        .ZN(n3989) );
  AND2_X1 U4909 ( .A1(n3990), .A2(n3989), .ZN(n5729) );
  MUX2_X1 U4910 ( .A(n3991), .B(n4006), .S(EBX_REG_24__SCAN_IN), .Z(n3995) );
  NAND2_X1 U4911 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n5467), .ZN(n3992) );
  AND2_X1 U4912 ( .A1(n3993), .A2(n3992), .ZN(n3994) );
  AND2_X1 U4913 ( .A1(n3995), .A2(n3994), .ZN(n5543) );
  MUX2_X1 U4914 ( .A(n4001), .B(n3956), .S(EBX_REG_25__SCAN_IN), .Z(n3996) );
  NAND2_X1 U4915 ( .A1(n3026), .A2(n3996), .ZN(n5536) );
  INV_X1 U4916 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6704) );
  NAND2_X1 U4917 ( .A1(n4004), .A2(n6704), .ZN(n4000) );
  INV_X1 U4918 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5580) );
  NAND2_X1 U4919 ( .A1(n4006), .A2(n5580), .ZN(n3998) );
  NAND2_X1 U4920 ( .A1(n5060), .A2(n6704), .ZN(n3997) );
  NAND3_X1 U4921 ( .A1(n3998), .A2(n3956), .A3(n3997), .ZN(n3999) );
  NAND2_X1 U4922 ( .A1(n4000), .A2(n3999), .ZN(n5529) );
  MUX2_X1 U4923 ( .A(n4001), .B(n4009), .S(EBX_REG_27__SCAN_IN), .Z(n4002) );
  OAI21_X1 U4924 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5468), .A(n4002), 
        .ZN(n4003) );
  INV_X1 U4925 ( .A(n4003), .ZN(n5522) );
  INV_X1 U4926 ( .A(EBX_REG_28__SCAN_IN), .ZN(n4007) );
  NAND2_X1 U4927 ( .A1(n4004), .A2(n4007), .ZN(n4012) );
  INV_X1 U4928 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4005) );
  NAND2_X1 U4929 ( .A1(n4006), .A2(n4005), .ZN(n4010) );
  NAND2_X1 U4930 ( .A1(n5060), .A2(n4007), .ZN(n4008) );
  NAND3_X1 U4931 ( .A1(n4010), .A2(n4009), .A3(n4008), .ZN(n4011) );
  AND2_X1 U4932 ( .A1(n4012), .A2(n4011), .ZN(n5496) );
  NOR2_X1 U4933 ( .A1(n5468), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5442)
         );
  INV_X1 U4934 ( .A(EBX_REG_29__SCAN_IN), .ZN(n6724) );
  NAND2_X1 U4935 ( .A1(n5468), .A2(EBX_REG_30__SCAN_IN), .ZN(n4014) );
  NAND2_X1 U4936 ( .A1(n5467), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4013) );
  NAND2_X1 U4937 ( .A1(n4014), .A2(n4013), .ZN(n4016) );
  INV_X1 U4938 ( .A(n4016), .ZN(n5464) );
  OAI21_X1 U4939 ( .B1(n5495), .B2(n4009), .A(n5464), .ZN(n4018) );
  INV_X1 U4940 ( .A(n4019), .ZN(n4015) );
  NAND2_X1 U4941 ( .A1(n4015), .A2(n4009), .ZN(n5466) );
  OAI211_X1 U4942 ( .C1(n4019), .C2(n5445), .A(n5466), .B(n4016), .ZN(n4017)
         );
  OAI21_X1 U4943 ( .B1(n4019), .B2(n4018), .A(n4017), .ZN(n5346) );
  INV_X1 U4944 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4020) );
  OR2_X1 U4945 ( .A1(n6123), .A2(n4020), .ZN(n4021) );
  NAND3_X1 U4946 ( .A1(n4029), .A2(n4028), .A3(n4027), .ZN(n4030) );
  NAND2_X1 U4947 ( .A1(n4031), .A2(n4030), .ZN(n4033) );
  AND2_X1 U4948 ( .A1(n4033), .A2(n4032), .ZN(n4085) );
  NOR2_X1 U4949 ( .A1(n4026), .A2(n4085), .ZN(n4044) );
  NAND2_X1 U4950 ( .A1(n4044), .A2(n4508), .ZN(n4052) );
  INV_X1 U4951 ( .A(n4508), .ZN(n6443) );
  INV_X1 U4952 ( .A(n6549), .ZN(n4036) );
  OR2_X1 U4953 ( .A1(n5063), .A2(n5069), .ZN(n4049) );
  AND2_X1 U4954 ( .A1(n4551), .A2(n6532), .ZN(n5091) );
  OAI21_X1 U4955 ( .B1(n5091), .B2(READREQUEST_REG_SCAN_IN), .A(n4036), .ZN(
        n4035) );
  OAI21_X1 U4956 ( .B1(n4036), .B2(n4049), .A(n4035), .ZN(U3474) );
  NAND2_X1 U4957 ( .A1(n4038), .A2(n4164), .ZN(n4039) );
  NAND2_X1 U4958 ( .A1(n4037), .A2(n4039), .ZN(n4091) );
  INV_X1 U4959 ( .A(n5055), .ZN(n4045) );
  OR2_X1 U4960 ( .A1(n4091), .A2(n4045), .ZN(n4084) );
  OR2_X1 U4961 ( .A1(n4091), .A2(n3152), .ZN(n4507) );
  NAND2_X1 U4962 ( .A1(n4084), .A2(n4507), .ZN(n4159) );
  OR2_X1 U4963 ( .A1(n4159), .A2(n4040), .ZN(n4043) );
  INV_X1 U4964 ( .A(n4085), .ZN(n4041) );
  OAI22_X1 U4965 ( .A1(n4161), .A2(n4506), .B1(n4026), .B2(n4041), .ZN(n4042)
         );
  AOI21_X1 U4966 ( .B1(n4043), .B2(n4506), .A(n4042), .ZN(n6423) );
  OR2_X1 U4967 ( .A1(n4044), .A2(n4040), .ZN(n4047) );
  NAND2_X1 U4968 ( .A1(n4506), .A2(n4045), .ZN(n4046) );
  NAND2_X1 U4969 ( .A1(n4047), .A2(n4046), .ZN(n5971) );
  INV_X1 U4970 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6463) );
  NAND2_X1 U4971 ( .A1(n4048), .A2(n6463), .ZN(n6461) );
  AOI21_X1 U4972 ( .B1(n4049), .B2(n6461), .A(READY_N), .ZN(n6553) );
  NOR2_X1 U4973 ( .A1(n5971), .A2(n6553), .ZN(n6418) );
  OR2_X1 U4974 ( .A1(n6418), .A2(n6443), .ZN(n5976) );
  NAND2_X1 U4975 ( .A1(n5976), .A2(MORE_REG_SCAN_IN), .ZN(n4050) );
  OAI21_X1 U4976 ( .B1(n6423), .B2(n5976), .A(n4050), .ZN(U3471) );
  AOI211_X1 U4977 ( .C1(MEMORYFETCH_REG_SCAN_IN), .C2(n4052), .A(n5091), .B(
        n4115), .ZN(n4053) );
  INV_X1 U4978 ( .A(n4053), .ZN(U2788) );
  OAI21_X1 U4979 ( .B1(n5156), .B2(n5071), .A(n4319), .ZN(n4060) );
  OR2_X1 U4980 ( .A1(n4055), .A2(n4319), .ZN(n4093) );
  INV_X1 U4981 ( .A(n4093), .ZN(n4056) );
  OAI21_X1 U4982 ( .B1(n4056), .B2(n5468), .A(n4236), .ZN(n4059) );
  NAND2_X1 U4983 ( .A1(n4057), .A2(n5204), .ZN(n4058) );
  AND4_X1 U4984 ( .A1(n4088), .A2(n4060), .A3(n4059), .A4(n4058), .ZN(n4061)
         );
  AND2_X1 U4985 ( .A1(n4062), .A2(n4061), .ZN(n4167) );
  AND4_X1 U4986 ( .A1(n4162), .A2(n4063), .A3(n4064), .A4(n4065), .ZN(n4066)
         );
  NAND2_X1 U4987 ( .A1(n4167), .A2(n4066), .ZN(n6400) );
  NAND2_X1 U4988 ( .A1(n6103), .A2(n6400), .ZN(n4079) );
  MUX2_X1 U4989 ( .A(n4068), .B(n4101), .S(n4067), .Z(n4069) );
  NAND2_X1 U4990 ( .A1(n4084), .A2(n4161), .ZN(n4455) );
  OAI21_X1 U4991 ( .B1(n4070), .B2(n4069), .A(n4455), .ZN(n4077) );
  NAND2_X1 U4992 ( .A1(n4112), .A2(n4025), .ZN(n4452) );
  INV_X1 U4993 ( .A(n4452), .ZN(n6405) );
  NAND2_X1 U4994 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4071) );
  INV_X1 U4995 ( .A(n4071), .ZN(n4072) );
  MUX2_X1 U4996 ( .A(n4072), .B(n4071), .S(n4073), .Z(n4075) );
  INV_X1 U4997 ( .A(n4450), .ZN(n4163) );
  AOI21_X1 U4998 ( .B1(n4067), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n4073), 
        .ZN(n4074) );
  NOR2_X1 U4999 ( .A1(n3776), .A2(n4074), .ZN(n4080) );
  AOI22_X1 U5000 ( .A1(n6405), .A2(n4075), .B1(n4163), .B2(n4080), .ZN(n4076)
         );
  AND2_X1 U5001 ( .A1(n4077), .A2(n4076), .ZN(n4078) );
  NAND2_X1 U5002 ( .A1(n4079), .A2(n4078), .ZN(n6397) );
  INV_X1 U5003 ( .A(n6539), .ZN(n5967) );
  AOI22_X1 U5004 ( .A1(n6397), .A2(n5967), .B1(n4080), .B2(n5407), .ZN(n4100)
         );
  NAND2_X1 U5005 ( .A1(n4452), .A2(n4064), .ZN(n4083) );
  INV_X1 U5006 ( .A(n6461), .ZN(n6431) );
  INV_X1 U5007 ( .A(n4081), .ZN(n4082) );
  AOI21_X1 U5008 ( .B1(n4083), .B2(n6431), .A(n4082), .ZN(n4098) );
  OR2_X1 U5009 ( .A1(n4506), .A2(READY_N), .ZN(n4097) );
  OR2_X1 U5010 ( .A1(n4084), .A2(n4506), .ZN(n4087) );
  INV_X1 U5011 ( .A(n4063), .ZN(n5966) );
  NOR2_X1 U5012 ( .A1(READY_N), .A2(n4085), .ZN(n4148) );
  NAND2_X1 U5013 ( .A1(n5966), .A2(n4148), .ZN(n4086) );
  NAND2_X1 U5014 ( .A1(n4087), .A2(n4086), .ZN(n4205) );
  INV_X1 U5015 ( .A(n4205), .ZN(n4096) );
  INV_X1 U5016 ( .A(n4088), .ZN(n4090) );
  OR3_X1 U5017 ( .A1(n4091), .A2(n4090), .A3(n4089), .ZN(n4092) );
  NAND2_X1 U5018 ( .A1(n4092), .A2(n4026), .ZN(n4155) );
  AND3_X1 U5019 ( .A1(n4155), .A2(n4094), .A3(n4093), .ZN(n4095) );
  OAI211_X1 U5020 ( .C1(n4098), .C2(n4097), .A(n4096), .B(n4095), .ZN(n6398)
         );
  INV_X1 U5021 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5977) );
  NOR2_X1 U5022 ( .A1(n6433), .A2(n6532), .ZN(n6429) );
  NAND2_X1 U5023 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6429), .ZN(n6527) );
  NOR2_X1 U5024 ( .A1(n5977), .A2(n6527), .ZN(n4099) );
  AOI21_X1 U5025 ( .B1(n4508), .B2(n6398), .A(n4099), .ZN(n5969) );
  NAND2_X1 U5026 ( .A1(n5050), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6528) );
  NAND2_X1 U5027 ( .A1(n5969), .A2(n6528), .ZN(n6537) );
  MUX2_X1 U5028 ( .A(n4101), .B(n4100), .S(n6537), .Z(n4102) );
  INV_X1 U5029 ( .A(n4102), .ZN(U3456) );
  NAND2_X1 U5030 ( .A1(n4104), .A2(n6400), .ZN(n4108) );
  INV_X1 U5031 ( .A(n4105), .ZN(n4106) );
  INV_X1 U5032 ( .A(n4067), .ZN(n5405) );
  NAND3_X1 U5033 ( .A1(n6401), .A2(n4106), .A3(n5405), .ZN(n4107) );
  OAI211_X1 U5034 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n4452), .A(n4108), .B(n4107), .ZN(n6408) );
  INV_X1 U5035 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4168) );
  NOR2_X1 U5036 ( .A1(n6532), .A2(n4168), .ZN(n5406) );
  INV_X1 U5037 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5685) );
  AOI22_X1 U5038 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5685), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n4281), .ZN(n5410) );
  AOI222_X1 U5039 ( .A1(n6408), .A2(n5967), .B1(n5406), .B2(n5410), .C1(n4109), 
        .C2(n5407), .ZN(n4111) );
  INV_X1 U5040 ( .A(n6537), .ZN(n5412) );
  NOR2_X1 U5041 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6438), .ZN(n6530)
         );
  OAI21_X1 U5042 ( .B1(n5412), .B2(n6530), .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), 
        .ZN(n4110) );
  OAI21_X1 U5043 ( .B1(n4111), .B2(n5412), .A(n4110), .ZN(U3460) );
  INV_X1 U5044 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6142) );
  INV_X1 U5045 ( .A(READY_N), .ZN(n6551) );
  AND2_X1 U5046 ( .A1(n4112), .A2(n6551), .ZN(n4113) );
  NAND2_X1 U5047 ( .A1(n6168), .A2(DATAI_13_), .ZN(n4125) );
  INV_X1 U5048 ( .A(n5063), .ZN(n6554) );
  NAND2_X1 U5049 ( .A1(n6554), .A2(READY_N), .ZN(n4114) );
  NAND2_X1 U5050 ( .A1(n6172), .A2(LWORD_REG_13__SCAN_IN), .ZN(n4116) );
  OAI211_X1 U5051 ( .C1(n6142), .C2(n4374), .A(n4125), .B(n4116), .ZN(U2952)
         );
  NAND2_X1 U5052 ( .A1(n6168), .A2(DATAI_12_), .ZN(n4124) );
  NAND2_X1 U5053 ( .A1(n6172), .A2(LWORD_REG_12__SCAN_IN), .ZN(n4117) );
  OAI211_X1 U5054 ( .C1(n5090), .C2(n4374), .A(n4124), .B(n4117), .ZN(U2951)
         );
  INV_X1 U5055 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6150) );
  NAND2_X1 U5056 ( .A1(n6168), .A2(DATAI_8_), .ZN(n4121) );
  NAND2_X1 U5057 ( .A1(n6172), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4118) );
  OAI211_X1 U5058 ( .C1(n6150), .C2(n4374), .A(n4121), .B(n4118), .ZN(U2947)
         );
  INV_X1 U5059 ( .A(EAX_REG_26__SCAN_IN), .ZN(n6733) );
  NAND2_X1 U5060 ( .A1(n6168), .A2(DATAI_10_), .ZN(n4179) );
  NAND2_X1 U5061 ( .A1(n6172), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4119) );
  OAI211_X1 U5062 ( .C1(n6733), .C2(n4374), .A(n4179), .B(n4119), .ZN(U2934)
         );
  INV_X1 U5063 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4381) );
  NAND2_X1 U5064 ( .A1(n6172), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4120) );
  OAI211_X1 U5065 ( .C1(n4381), .C2(n4374), .A(n4121), .B(n4120), .ZN(U2932)
         );
  INV_X1 U5066 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4386) );
  NAND2_X1 U5067 ( .A1(n6168), .A2(DATAI_11_), .ZN(n6170) );
  NAND2_X1 U5068 ( .A1(n6172), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4122) );
  OAI211_X1 U5069 ( .C1(n4374), .C2(n4386), .A(n6170), .B(n4122), .ZN(U2935)
         );
  INV_X1 U5070 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4390) );
  NAND2_X1 U5071 ( .A1(n6172), .A2(UWORD_REG_12__SCAN_IN), .ZN(n4123) );
  OAI211_X1 U5072 ( .C1(n4390), .C2(n4374), .A(n4124), .B(n4123), .ZN(U2936)
         );
  AOI22_X1 U5073 ( .A1(n6173), .A2(EAX_REG_29__SCAN_IN), .B1(
        UWORD_REG_13__SCAN_IN), .B2(n6172), .ZN(n4126) );
  NAND2_X1 U5074 ( .A1(n4126), .A2(n4125), .ZN(U2937) );
  AOI22_X1 U5075 ( .A1(n6173), .A2(EAX_REG_23__SCAN_IN), .B1(
        UWORD_REG_7__SCAN_IN), .B2(n6172), .ZN(n4127) );
  INV_X1 U5076 ( .A(DATAI_7_), .ZN(n4339) );
  OR2_X1 U5077 ( .A1(n4206), .A2(n4339), .ZN(n4128) );
  NAND2_X1 U5078 ( .A1(n4127), .A2(n4128), .ZN(U2931) );
  AOI22_X1 U5079 ( .A1(n6173), .A2(EAX_REG_7__SCAN_IN), .B1(
        LWORD_REG_7__SCAN_IN), .B2(n6172), .ZN(n4129) );
  NAND2_X1 U5080 ( .A1(n4129), .A2(n4128), .ZN(U2946) );
  AOI22_X1 U5081 ( .A1(n6173), .A2(EAX_REG_22__SCAN_IN), .B1(
        UWORD_REG_6__SCAN_IN), .B2(n6172), .ZN(n4130) );
  NAND2_X1 U5082 ( .A1(n6168), .A2(DATAI_6_), .ZN(n4131) );
  NAND2_X1 U5083 ( .A1(n4130), .A2(n4131), .ZN(U2930) );
  AOI22_X1 U5084 ( .A1(n6173), .A2(EAX_REG_6__SCAN_IN), .B1(
        LWORD_REG_6__SCAN_IN), .B2(n6172), .ZN(n4132) );
  NAND2_X1 U5085 ( .A1(n4132), .A2(n4131), .ZN(U2945) );
  AOI22_X1 U5086 ( .A1(n6173), .A2(EAX_REG_25__SCAN_IN), .B1(
        UWORD_REG_9__SCAN_IN), .B2(n6172), .ZN(n4133) );
  NAND2_X1 U5087 ( .A1(n6168), .A2(DATAI_9_), .ZN(n4181) );
  NAND2_X1 U5088 ( .A1(n4133), .A2(n4181), .ZN(U2933) );
  INV_X1 U5089 ( .A(DATAI_0_), .ZN(n4299) );
  AOI22_X1 U5090 ( .A1(n6173), .A2(EAX_REG_0__SCAN_IN), .B1(
        LWORD_REG_0__SCAN_IN), .B2(n6172), .ZN(n4134) );
  OAI21_X1 U5091 ( .B1(n4299), .B2(n4206), .A(n4134), .ZN(U2939) );
  INV_X1 U5092 ( .A(DATAI_1_), .ZN(n4324) );
  AOI22_X1 U5093 ( .A1(n6173), .A2(EAX_REG_1__SCAN_IN), .B1(
        LWORD_REG_1__SCAN_IN), .B2(n6172), .ZN(n4135) );
  OAI21_X1 U5094 ( .B1(n4324), .B2(n4206), .A(n4135), .ZN(U2940) );
  INV_X1 U5095 ( .A(DATAI_5_), .ZN(n6569) );
  AOI22_X1 U5096 ( .A1(n6173), .A2(EAX_REG_5__SCAN_IN), .B1(
        LWORD_REG_5__SCAN_IN), .B2(n6172), .ZN(n4136) );
  OAI21_X1 U5097 ( .B1(n6569), .B2(n4206), .A(n4136), .ZN(U2944) );
  INV_X1 U5098 ( .A(DATAI_3_), .ZN(n4314) );
  AOI22_X1 U5099 ( .A1(n6173), .A2(EAX_REG_3__SCAN_IN), .B1(
        LWORD_REG_3__SCAN_IN), .B2(n6172), .ZN(n4137) );
  OAI21_X1 U5100 ( .B1(n4314), .B2(n4206), .A(n4137), .ZN(U2942) );
  AOI22_X1 U5101 ( .A1(n6173), .A2(EAX_REG_2__SCAN_IN), .B1(
        LWORD_REG_2__SCAN_IN), .B2(n6172), .ZN(n4138) );
  OAI21_X1 U5102 ( .B1(n4201), .B2(n4206), .A(n4138), .ZN(U2941) );
  INV_X1 U5103 ( .A(DATAI_4_), .ZN(n6721) );
  AOI22_X1 U5104 ( .A1(n6173), .A2(EAX_REG_4__SCAN_IN), .B1(
        LWORD_REG_4__SCAN_IN), .B2(n6172), .ZN(n4139) );
  OAI21_X1 U5105 ( .B1(n6721), .B2(n4206), .A(n4139), .ZN(U2943) );
  NAND2_X1 U5106 ( .A1(n4140), .A2(n4753), .ZN(n4143) );
  INV_X1 U5107 ( .A(n4247), .ZN(n4234) );
  NAND2_X1 U5108 ( .A1(n4164), .A2(n3160), .ZN(n4250) );
  INV_X1 U5109 ( .A(n4250), .ZN(n4141) );
  AOI21_X1 U5110 ( .B1(n4234), .B2(n5063), .A(n4141), .ZN(n4142) );
  NAND2_X1 U5111 ( .A1(n4143), .A2(n4142), .ZN(n4243) );
  XNOR2_X1 U5112 ( .A(n4243), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4505)
         );
  NAND2_X1 U5113 ( .A1(n4144), .A2(n6461), .ZN(n5073) );
  NAND2_X1 U5114 ( .A1(n5073), .A2(n6551), .ZN(n4145) );
  OAI211_X1 U5115 ( .C1(n4064), .C2(n4145), .A(n5071), .B(n5156), .ZN(n4147)
         );
  NAND2_X1 U5116 ( .A1(n4147), .A2(n4146), .ZN(n4151) );
  NAND2_X1 U5117 ( .A1(n4112), .A2(n6461), .ZN(n4149) );
  NAND3_X1 U5118 ( .A1(n4149), .A2(n4148), .A3(n4319), .ZN(n4150) );
  OAI21_X1 U5119 ( .B1(n4151), .B2(n4506), .A(n4150), .ZN(n4152) );
  INV_X1 U5120 ( .A(n4152), .ZN(n4154) );
  NAND3_X1 U5121 ( .A1(n4506), .A2(n6401), .A3(n4112), .ZN(n4153) );
  NAND3_X1 U5122 ( .A1(n4155), .A2(n4154), .A3(n4153), .ZN(n4156) );
  NOR2_X1 U5123 ( .A1(n4170), .A2(n3142), .ZN(n4158) );
  NOR3_X1 U5124 ( .A1(n4159), .A2(n4158), .A3(n4157), .ZN(n4160) );
  INV_X1 U5125 ( .A(n4162), .ZN(n4165) );
  AOI21_X1 U5126 ( .B1(n4165), .B2(n4164), .A(n4163), .ZN(n4166) );
  AOI21_X1 U5127 ( .B1(n4167), .B2(n4166), .A(n4173), .ZN(n5940) );
  AOI22_X1 U5128 ( .A1(n5940), .A2(n4168), .B1(n4173), .B2(n6216), .ZN(n5383)
         );
  OAI21_X1 U5129 ( .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n6212), .A(n5383), 
        .ZN(n4396) );
  NOR2_X1 U5130 ( .A1(n6280), .A2(n5940), .ZN(n5946) );
  INV_X1 U5131 ( .A(n5946), .ZN(n4169) );
  OAI22_X1 U5132 ( .A1(n4396), .A2(n5961), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n4169), .ZN(n4177) );
  OR2_X1 U5133 ( .A1(n4064), .A2(n6554), .ZN(n6428) );
  OAI21_X1 U5134 ( .B1(n4170), .B2(n4308), .A(n6428), .ZN(n4171) );
  INV_X1 U5135 ( .A(n4171), .ZN(n4172) );
  OR2_X1 U5136 ( .A1(n5468), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4175)
         );
  AND2_X1 U5137 ( .A1(n4175), .A2(n4174), .ZN(n5068) );
  AND2_X1 U5138 ( .A1(n6277), .A2(REIP_REG_0__SCAN_IN), .ZN(n4515) );
  AOI21_X1 U5139 ( .B1(n6279), .B2(n5068), .A(n4515), .ZN(n4176) );
  OAI211_X1 U5140 ( .C1(n4505), .C2(n5906), .A(n4177), .B(n4176), .ZN(U3018)
         );
  INV_X1 U5141 ( .A(LWORD_REG_10__SCAN_IN), .ZN(n6591) );
  NAND2_X1 U5142 ( .A1(n6173), .A2(EAX_REG_10__SCAN_IN), .ZN(n4178) );
  OAI211_X1 U5143 ( .C1(n4199), .C2(n6591), .A(n4179), .B(n4178), .ZN(U2949)
         );
  INV_X1 U5144 ( .A(LWORD_REG_9__SCAN_IN), .ZN(n6725) );
  NAND2_X1 U5145 ( .A1(n6173), .A2(EAX_REG_9__SCAN_IN), .ZN(n4180) );
  OAI211_X1 U5146 ( .C1(n4199), .C2(n6725), .A(n4181), .B(n4180), .ZN(U2948)
         );
  AOI222_X1 U5147 ( .A1(n6172), .A2(UWORD_REG_5__SCAN_IN), .B1(n6168), .B2(
        DATAI_5_), .C1(EAX_REG_21__SCAN_IN), .C2(n6173), .ZN(n4182) );
  INV_X1 U5148 ( .A(n4182), .ZN(U2929) );
  NAND2_X1 U5149 ( .A1(n4183), .A2(n4184), .ZN(n4228) );
  INV_X1 U5150 ( .A(n4228), .ZN(n4189) );
  INV_X1 U5151 ( .A(n4185), .ZN(n4186) );
  NOR3_X1 U5152 ( .A1(n4187), .A2(n4216), .A3(n4186), .ZN(n4188) );
  NOR2_X1 U5153 ( .A1(n4189), .A2(n4188), .ZN(n6206) );
  INV_X1 U5154 ( .A(n6206), .ZN(n4212) );
  INV_X1 U5155 ( .A(EBX_REG_2__SCAN_IN), .ZN(n4192) );
  INV_X1 U5156 ( .A(n4191), .ZN(n4360) );
  XNOR2_X1 U5157 ( .A(n4190), .B(n4360), .ZN(n6276) );
  OAI222_X1 U5158 ( .A1(n6118), .A2(n4212), .B1(n4192), .B2(n6123), .C1(n5546), 
        .C2(n6276), .ZN(U2857) );
  INV_X1 U5159 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n4193) );
  INV_X1 U5160 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4405) );
  OAI222_X1 U5161 ( .A1(n4324), .A2(n4206), .B1(n4193), .B2(n4199), .C1(n4374), 
        .C2(n4405), .ZN(U2925) );
  INV_X1 U5162 ( .A(UWORD_REG_4__SCAN_IN), .ZN(n4194) );
  INV_X1 U5163 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4379) );
  OAI222_X1 U5164 ( .A1(n6721), .A2(n4206), .B1(n4194), .B2(n4199), .C1(n4374), 
        .C2(n4379), .ZN(U2928) );
  INV_X1 U5165 ( .A(DATAI_15_), .ZN(n4196) );
  INV_X1 U5166 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4195) );
  INV_X1 U5167 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6139) );
  OAI222_X1 U5168 ( .A1(n4196), .A2(n4206), .B1(n4195), .B2(n4199), .C1(n4374), 
        .C2(n6139), .ZN(U2954) );
  INV_X1 U5169 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n4197) );
  INV_X1 U5170 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4384) );
  OAI222_X1 U5171 ( .A1(n4314), .A2(n4206), .B1(n4197), .B2(n4199), .C1(n4374), 
        .C2(n4384), .ZN(U2927) );
  INV_X1 U5172 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n4198) );
  INV_X1 U5173 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4403) );
  OAI222_X1 U5174 ( .A1(n4299), .A2(n4206), .B1(n4198), .B2(n4199), .C1(n4374), 
        .C2(n4403), .ZN(U2924) );
  INV_X1 U5175 ( .A(DATAI_2_), .ZN(n4201) );
  INV_X1 U5176 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n4200) );
  INV_X1 U5177 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4388) );
  OAI222_X1 U5178 ( .A1(n4201), .A2(n4206), .B1(n4200), .B2(n4199), .C1(n4374), 
        .C2(n4388), .ZN(U2926) );
  NAND2_X1 U5179 ( .A1(n4202), .A2(n3162), .ZN(n4203) );
  NOR2_X1 U5180 ( .A1(n4065), .A2(n4203), .ZN(n4204) );
  OAI21_X1 U5181 ( .B1(n4205), .B2(n4204), .A(n4508), .ZN(n4207) );
  AND2_X1 U5182 ( .A1(n3120), .A2(n3163), .ZN(n5157) );
  INV_X1 U5183 ( .A(n5157), .ZN(n4208) );
  AND2_X1 U5184 ( .A1(n4208), .A2(n5156), .ZN(n4209) );
  INV_X1 U5185 ( .A(n4209), .ZN(n4210) );
  AOI22_X1 U5186 ( .A1(n5301), .A2(DATAI_2_), .B1(n6130), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n4211) );
  OAI21_X1 U5187 ( .B1(n4212), .B2(n5867), .A(n4211), .ZN(U2889) );
  NOR2_X1 U5188 ( .A1(n4214), .A2(n4213), .ZN(n4215) );
  NOR2_X1 U5189 ( .A1(n4216), .A2(n4215), .ZN(n5504) );
  INV_X1 U5190 ( .A(n5504), .ZN(n4353) );
  AOI22_X1 U5191 ( .A1(n5301), .A2(DATAI_1_), .B1(n6130), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n4217) );
  OAI21_X1 U5192 ( .B1(n4353), .B2(n5867), .A(n4217), .ZN(U2890) );
  CLKBUF_X1 U5193 ( .A(n4218), .Z(n4365) );
  NAND2_X1 U5194 ( .A1(n4219), .A2(n4220), .ZN(n4221) );
  NAND2_X1 U5195 ( .A1(n4365), .A2(n4221), .ZN(n5122) );
  INV_X1 U5196 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4224) );
  OR2_X1 U5197 ( .A1(n4356), .A2(n4222), .ZN(n4223) );
  NAND2_X1 U5198 ( .A1(n4368), .A2(n4223), .ZN(n5116) );
  OAI222_X1 U5199 ( .A1(n5122), .A2(n6118), .B1(n6123), .B2(n4224), .C1(n5116), 
        .C2(n5546), .ZN(U2854) );
  XOR2_X1 U5200 ( .A(n4226), .B(n4225), .Z(n5080) );
  INV_X1 U5201 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6167) );
  OAI222_X1 U5202 ( .A1(n5867), .A2(n5080), .B1(n5088), .B2(n4299), .C1(n5432), 
        .C2(n6167), .ZN(U2891) );
  INV_X1 U5203 ( .A(EAX_REG_5__SCAN_IN), .ZN(n6155) );
  OAI222_X1 U5204 ( .A1(n5122), .A2(n5867), .B1(n5088), .B2(n6569), .C1(n5432), 
        .C2(n6155), .ZN(U2886) );
  AND2_X1 U5205 ( .A1(n4183), .A2(n4227), .ZN(n4231) );
  AOI21_X1 U5206 ( .B1(n4229), .B2(n4228), .A(n4231), .ZN(n4738) );
  INV_X1 U5207 ( .A(n4738), .ZN(n6106) );
  INV_X1 U5208 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6159) );
  OAI222_X1 U5209 ( .A1(n6106), .A2(n5867), .B1(n5088), .B2(n4314), .C1(n5432), 
        .C2(n6159), .ZN(U2888) );
  OR2_X1 U5210 ( .A1(n4231), .A2(n4230), .ZN(n4232) );
  AND2_X1 U5211 ( .A1(n4219), .A2(n4232), .ZN(n6195) );
  INV_X1 U5212 ( .A(n6195), .ZN(n4358) );
  INV_X1 U5213 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6157) );
  OAI222_X1 U5214 ( .A1(n4358), .A2(n5867), .B1(n5088), .B2(n6721), .C1(n5432), 
        .C2(n6157), .ZN(U2887) );
  NAND2_X1 U5215 ( .A1(n4233), .A2(n4753), .ZN(n4240) );
  XNOR2_X1 U5216 ( .A(n4234), .B(n4248), .ZN(n4235) );
  NAND2_X1 U5217 ( .A1(n4235), .A2(n5063), .ZN(n4238) );
  NOR2_X1 U5218 ( .A1(n4236), .A2(n3120), .ZN(n4237) );
  AND2_X1 U5219 ( .A1(n4238), .A2(n4237), .ZN(n4239) );
  NAND2_X1 U5220 ( .A1(n4240), .A2(n4239), .ZN(n4393) );
  NAND2_X1 U5221 ( .A1(n4243), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4241)
         );
  NAND2_X1 U5222 ( .A1(n4241), .A2(n4281), .ZN(n4244) );
  AND2_X1 U5223 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4242) );
  NAND2_X1 U5224 ( .A1(n4243), .A2(n4242), .ZN(n4245) );
  AND2_X1 U5225 ( .A1(n4244), .A2(n4245), .ZN(n4394) );
  INV_X1 U5226 ( .A(n4245), .ZN(n4246) );
  AOI21_X2 U5227 ( .B1(n4393), .B2(n4394), .A(n4246), .ZN(n6202) );
  INV_X1 U5228 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6286) );
  NAND2_X1 U5229 ( .A1(n4248), .A2(n4247), .ZN(n4258) );
  XNOR2_X1 U5230 ( .A(n4258), .B(n4257), .ZN(n4249) );
  NAND2_X1 U5231 ( .A1(n4249), .A2(n5063), .ZN(n4251) );
  NAND2_X1 U5232 ( .A1(n4251), .A2(n4250), .ZN(n4252) );
  OAI21_X1 U5233 ( .B1(n6202), .B2(n6286), .A(n6200), .ZN(n4255) );
  NAND2_X1 U5234 ( .A1(n6202), .A2(n6286), .ZN(n4254) );
  NAND2_X1 U5235 ( .A1(n4256), .A2(n4753), .ZN(n4262) );
  NAND2_X1 U5236 ( .A1(n4258), .A2(n4257), .ZN(n4267) );
  XNOR2_X1 U5237 ( .A(n4267), .B(n4259), .ZN(n4260) );
  NAND2_X1 U5238 ( .A1(n4260), .A2(n5063), .ZN(n4261) );
  NAND2_X1 U5239 ( .A1(n4262), .A2(n4261), .ZN(n4263) );
  INV_X1 U5240 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6274) );
  XNOR2_X1 U5241 ( .A(n4263), .B(n6274), .ZN(n4732) );
  NAND2_X1 U5242 ( .A1(n4734), .A2(n4732), .ZN(n4733) );
  NAND2_X1 U5243 ( .A1(n4263), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4264)
         );
  NAND2_X1 U5244 ( .A1(n4265), .A2(n4753), .ZN(n4270) );
  NAND2_X1 U5245 ( .A1(n4267), .A2(n4266), .ZN(n4747) );
  XNOR2_X1 U5246 ( .A(n4747), .B(n4744), .ZN(n4268) );
  NAND2_X1 U5247 ( .A1(n4268), .A2(n5063), .ZN(n4269) );
  NAND2_X1 U5248 ( .A1(n4270), .A2(n4269), .ZN(n4271) );
  INV_X1 U5249 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n6265) );
  XNOR2_X1 U5250 ( .A(n4271), .B(n6265), .ZN(n6192) );
  NAND2_X1 U5251 ( .A1(n4271), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n4272)
         );
  NAND2_X1 U5252 ( .A1(n4273), .A2(n4753), .ZN(n4278) );
  INV_X1 U5253 ( .A(n4747), .ZN(n4274) );
  NAND2_X1 U5254 ( .A1(n4274), .A2(n4744), .ZN(n4275) );
  XNOR2_X1 U5255 ( .A(n4275), .B(n4745), .ZN(n4276) );
  NAND2_X1 U5256 ( .A1(n4276), .A2(n5063), .ZN(n4277) );
  NAND2_X1 U5257 ( .A1(n4278), .A2(n4277), .ZN(n4740) );
  INV_X1 U5258 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4284) );
  XNOR2_X1 U5259 ( .A(n4740), .B(n4284), .ZN(n4279) );
  NAND2_X1 U5260 ( .A1(n4280), .A2(n4279), .ZN(n4742) );
  OAI21_X1 U5261 ( .B1(n4280), .B2(n4279), .A(n3007), .ZN(n4731) );
  AOI21_X1 U5262 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n6282) );
  NAND2_X1 U5263 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n6262) );
  NOR2_X1 U5264 ( .A1(n6282), .A2(n6262), .ZN(n4832) );
  NOR2_X1 U5265 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5961), .ZN(n4395)
         );
  NOR2_X1 U5266 ( .A1(n6286), .A2(n4281), .ZN(n6281) );
  INV_X1 U5267 ( .A(n6281), .ZN(n4282) );
  NOR2_X1 U5268 ( .A1(n6262), .A2(n4282), .ZN(n4833) );
  AOI22_X1 U5269 ( .A1(n6280), .A2(n4832), .B1(n6287), .B2(n4833), .ZN(n4285)
         );
  NAND2_X1 U5270 ( .A1(n6212), .A2(n5384), .ZN(n5921) );
  NAND2_X1 U5271 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4832), .ZN(n4283)
         );
  OAI21_X1 U5272 ( .B1(n5384), .B2(n6281), .A(n5383), .ZN(n6285) );
  AOI21_X1 U5273 ( .B1(n5921), .B2(n4283), .A(n6285), .ZN(n6255) );
  AOI21_X1 U5274 ( .B1(n4285), .B2(n4284), .A(n6255), .ZN(n4287) );
  INV_X1 U5275 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6479) );
  OAI22_X1 U5276 ( .A1(n5116), .A2(n6217), .B1(n6479), .B2(n6216), .ZN(n4286)
         );
  NOR2_X1 U5277 ( .A1(n4287), .A2(n4286), .ZN(n4288) );
  OAI21_X1 U5278 ( .B1(n5906), .B2(n4731), .A(n4288), .ZN(U3013) );
  NAND3_X1 U5279 ( .A1(n6718), .A2(n4946), .A3(n4787), .ZN(n4895) );
  NOR2_X1 U5280 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4895), .ZN(n4342)
         );
  INV_X1 U5281 ( .A(n4342), .ZN(n4291) );
  AND2_X1 U5282 ( .A1(n4300), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6306) );
  INV_X1 U5283 ( .A(n4470), .ZN(n4289) );
  OR2_X1 U5284 ( .A1(n6305), .A2(n4289), .ZN(n5224) );
  INV_X1 U5285 ( .A(n5224), .ZN(n4290) );
  NOR2_X1 U5286 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATE2_REG_1__SCAN_IN), .ZN(
        n6555) );
  OAI21_X1 U5287 ( .B1(n4290), .B2(n6433), .A(n4612), .ZN(n5221) );
  AOI211_X1 U5288 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4291), .A(n6306), .B(
        n5221), .ZN(n4298) );
  INV_X1 U5289 ( .A(n3348), .ZN(n4294) );
  INV_X1 U5290 ( .A(n5778), .ZN(n4293) );
  INV_X1 U5291 ( .A(n4253), .ZN(n4472) );
  NAND3_X1 U5292 ( .A1(n4294), .A2(n4293), .A3(n4472), .ZN(n4893) );
  INV_X1 U5293 ( .A(n4893), .ZN(n4888) );
  NAND2_X1 U5294 ( .A1(n4888), .A2(n4892), .ZN(n4344) );
  NAND2_X1 U5295 ( .A1(n3015), .A2(n4545), .ZN(n4519) );
  NAND2_X1 U5296 ( .A1(n5778), .A2(n4140), .ZN(n5004) );
  NOR2_X1 U5297 ( .A1(n4519), .A2(n5004), .ZN(n4416) );
  OAI21_X1 U5298 ( .B1(n4926), .B2(n4416), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4296) );
  OR2_X1 U5299 ( .A1(n4104), .A2(n5328), .ZN(n4857) );
  OR2_X1 U5300 ( .A1(n4857), .A2(n6103), .ZN(n4890) );
  NAND3_X1 U5301 ( .A1(n4296), .A2(n4551), .A3(n4890), .ZN(n4297) );
  NOR2_X1 U5302 ( .A1(n4299), .A2(n4471), .ZN(n6312) );
  INV_X1 U5303 ( .A(n4551), .ZN(n5000) );
  NOR2_X1 U5304 ( .A1(n4300), .A2(n6433), .ZN(n6316) );
  INV_X1 U5305 ( .A(n6316), .ZN(n4944) );
  OAI22_X1 U5306 ( .A1(n4890), .A2(n5000), .B1(n4944), .B2(n5224), .ZN(n4346)
         );
  AND2_X1 U5307 ( .A1(n5050), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5052) );
  NAND2_X1 U5308 ( .A1(n5052), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6451) );
  OR2_X1 U5309 ( .A1(n6451), .A2(n5000), .ZN(n5679) );
  NAND2_X1 U5310 ( .A1(n6205), .A2(DATAI_16_), .ZN(n6324) );
  INV_X1 U5311 ( .A(n6528), .ZN(n4302) );
  NAND2_X1 U5312 ( .A1(n4340), .A2(n5071), .ZN(n4969) );
  INV_X1 U5313 ( .A(DATAI_24_), .ZN(n4303) );
  NOR2_X1 U5314 ( .A1(n5679), .A2(n4303), .ZN(n6321) );
  AOI22_X1 U5315 ( .A1(n6311), .A2(n4342), .B1(n6321), .B2(n4416), .ZN(n4304)
         );
  OAI21_X1 U5316 ( .B1(n6324), .B2(n4344), .A(n4304), .ZN(n4305) );
  AOI21_X1 U5317 ( .B1(n6312), .B2(n4346), .A(n4305), .ZN(n4306) );
  OAI21_X1 U5318 ( .B1(n4349), .B2(n4307), .A(n4306), .ZN(U3020) );
  NOR2_X1 U5319 ( .A1(n6721), .A2(n4471), .ZN(n6340) );
  NAND2_X1 U5320 ( .A1(n6205), .A2(DATAI_20_), .ZN(n6344) );
  NAND2_X1 U5321 ( .A1(n4340), .A2(n4308), .ZN(n4987) );
  INV_X1 U5322 ( .A(DATAI_28_), .ZN(n4309) );
  NOR2_X1 U5323 ( .A1(n5679), .A2(n4309), .ZN(n6341) );
  AOI22_X1 U5324 ( .A1(n6339), .A2(n4342), .B1(n6341), .B2(n4416), .ZN(n4310)
         );
  OAI21_X1 U5325 ( .B1(n6344), .B2(n4344), .A(n4310), .ZN(n4311) );
  AOI21_X1 U5326 ( .B1(n6340), .B2(n4346), .A(n4311), .ZN(n4312) );
  OAI21_X1 U5327 ( .B1(n4349), .B2(n4313), .A(n4312), .ZN(U3024) );
  NOR2_X1 U5328 ( .A1(n4314), .A2(n4471), .ZN(n6382) );
  NAND2_X1 U5329 ( .A1(n6205), .A2(DATAI_19_), .ZN(n6338) );
  NAND2_X1 U5330 ( .A1(n4340), .A2(n3160), .ZN(n4954) );
  NAND2_X1 U5331 ( .A1(n6205), .A2(DATAI_27_), .ZN(n6385) );
  INV_X1 U5332 ( .A(n6385), .ZN(n6335) );
  AOI22_X1 U5333 ( .A1(n6381), .A2(n4342), .B1(n6335), .B2(n4416), .ZN(n4315)
         );
  OAI21_X1 U5334 ( .B1(n6338), .B2(n4344), .A(n4315), .ZN(n4316) );
  AOI21_X1 U5335 ( .B1(n6382), .B2(n4346), .A(n4316), .ZN(n4317) );
  OAI21_X1 U5336 ( .B1(n4349), .B2(n4318), .A(n4317), .ZN(U3023) );
  NOR2_X1 U5337 ( .A1(n4201), .A2(n4471), .ZN(n6330) );
  NAND2_X1 U5338 ( .A1(n6205), .A2(DATAI_18_), .ZN(n6334) );
  NAND2_X1 U5339 ( .A1(n4340), .A2(n4319), .ZN(n4977) );
  INV_X1 U5340 ( .A(DATAI_26_), .ZN(n6740) );
  NOR2_X1 U5341 ( .A1(n5679), .A2(n6740), .ZN(n6331) );
  AOI22_X1 U5342 ( .A1(n6329), .A2(n4342), .B1(n6331), .B2(n4416), .ZN(n4320)
         );
  OAI21_X1 U5343 ( .B1(n6334), .B2(n4344), .A(n4320), .ZN(n4321) );
  AOI21_X1 U5344 ( .B1(n6330), .B2(n4346), .A(n4321), .ZN(n4322) );
  OAI21_X1 U5345 ( .B1(n4349), .B2(n4323), .A(n4322), .ZN(U3022) );
  NAND2_X1 U5346 ( .A1(n6205), .A2(DATAI_17_), .ZN(n6328) );
  NAND2_X1 U5347 ( .A1(n4340), .A2(n4112), .ZN(n4959) );
  NAND2_X1 U5348 ( .A1(n6205), .A2(DATAI_25_), .ZN(n6379) );
  INV_X1 U5349 ( .A(n6379), .ZN(n6325) );
  AOI22_X1 U5350 ( .A1(n6375), .A2(n4342), .B1(n6325), .B2(n4416), .ZN(n4325)
         );
  OAI21_X1 U5351 ( .B1(n6328), .B2(n4344), .A(n4325), .ZN(n4326) );
  AOI21_X1 U5352 ( .B1(n6376), .B2(n4346), .A(n4326), .ZN(n4327) );
  OAI21_X1 U5353 ( .B1(n4349), .B2(n4328), .A(n4327), .ZN(U3021) );
  NOR2_X1 U5354 ( .A1(n6569), .A2(n4471), .ZN(n6346) );
  NAND2_X1 U5355 ( .A1(n6205), .A2(DATAI_21_), .ZN(n6350) );
  NAND2_X1 U5356 ( .A1(n4340), .A2(n4329), .ZN(n4973) );
  INV_X1 U5357 ( .A(DATAI_29_), .ZN(n4330) );
  NOR2_X1 U5358 ( .A1(n5679), .A2(n4330), .ZN(n6347) );
  AOI22_X1 U5359 ( .A1(n6345), .A2(n4342), .B1(n6347), .B2(n4416), .ZN(n4331)
         );
  OAI21_X1 U5360 ( .B1(n6350), .B2(n4344), .A(n4331), .ZN(n4332) );
  AOI21_X1 U5361 ( .B1(n6346), .B2(n4346), .A(n4332), .ZN(n4333) );
  OAI21_X1 U5362 ( .B1(n4349), .B2(n4334), .A(n4333), .ZN(U3025) );
  INV_X1 U5363 ( .A(DATAI_6_), .ZN(n6593) );
  NOR2_X1 U5364 ( .A1(n6593), .A2(n4471), .ZN(n6391) );
  NAND2_X1 U5365 ( .A1(n6205), .A2(DATAI_22_), .ZN(n6354) );
  NAND2_X1 U5366 ( .A1(n4340), .A2(n3162), .ZN(n4964) );
  NAND2_X1 U5367 ( .A1(n6205), .A2(DATAI_30_), .ZN(n6396) );
  INV_X1 U5368 ( .A(n6396), .ZN(n6351) );
  AOI22_X1 U5369 ( .A1(n6389), .A2(n4342), .B1(n6351), .B2(n4416), .ZN(n4335)
         );
  OAI21_X1 U5370 ( .B1(n6354), .B2(n4344), .A(n4335), .ZN(n4336) );
  AOI21_X1 U5371 ( .B1(n6391), .B2(n4346), .A(n4336), .ZN(n4337) );
  OAI21_X1 U5372 ( .B1(n4349), .B2(n4338), .A(n4337), .ZN(U3026) );
  NOR2_X1 U5373 ( .A1(n4339), .A2(n4471), .ZN(n6358) );
  NAND2_X1 U5374 ( .A1(n6205), .A2(DATAI_23_), .ZN(n6364) );
  NAND2_X1 U5375 ( .A1(n4340), .A2(n3163), .ZN(n4981) );
  INV_X1 U5376 ( .A(DATAI_31_), .ZN(n4341) );
  NOR2_X1 U5377 ( .A1(n5679), .A2(n4341), .ZN(n6360) );
  AOI22_X1 U5378 ( .A1(n6356), .A2(n4342), .B1(n6360), .B2(n4416), .ZN(n4343)
         );
  OAI21_X1 U5379 ( .B1(n6364), .B2(n4344), .A(n4343), .ZN(n4345) );
  AOI21_X1 U5380 ( .B1(n6358), .B2(n4346), .A(n4345), .ZN(n4347) );
  OAI21_X1 U5381 ( .B1(n4349), .B2(n4348), .A(n4347), .ZN(U3027) );
  INV_X1 U5382 ( .A(n6123), .ZN(n6562) );
  AOI22_X1 U5383 ( .A1(n6563), .A2(n5068), .B1(EBX_REG_0__SCAN_IN), .B2(n6562), 
        .ZN(n4350) );
  OAI21_X1 U5384 ( .B1(n5080), .B2(n6118), .A(n4350), .ZN(U2859) );
  OAI21_X1 U5385 ( .B1(n5509), .B2(n5060), .A(n4351), .ZN(n4399) );
  AOI22_X1 U5386 ( .A1(n6563), .A2(n4399), .B1(EBX_REG_1__SCAN_IN), .B2(n6562), 
        .ZN(n4352) );
  OAI21_X1 U5387 ( .B1(n4353), .B2(n6118), .A(n4352), .ZN(U2858) );
  AND2_X1 U5388 ( .A1(n4361), .A2(n4354), .ZN(n4355) );
  NOR2_X1 U5389 ( .A1(n4356), .A2(n4355), .ZN(n6259) );
  AOI22_X1 U5390 ( .A1(n6259), .A2(n6563), .B1(EBX_REG_4__SCAN_IN), .B2(n6562), 
        .ZN(n4357) );
  OAI21_X1 U5391 ( .B1(n4358), .B2(n6118), .A(n4357), .ZN(U2855) );
  OAI21_X1 U5392 ( .B1(n4190), .B2(n4360), .A(n4359), .ZN(n4362) );
  NAND2_X1 U5393 ( .A1(n4362), .A2(n4361), .ZN(n6266) );
  INV_X1 U5394 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4363) );
  OAI222_X1 U5395 ( .A1(n6266), .A2(n5546), .B1(n4363), .B2(n6123), .C1(n6106), 
        .C2(n6118), .ZN(U2856) );
  NAND2_X1 U5396 ( .A1(n4365), .A2(n4364), .ZN(n4366) );
  AND2_X1 U5397 ( .A1(n4646), .A2(n4366), .ZN(n6187) );
  INV_X1 U5398 ( .A(n6187), .ZN(n4407) );
  NAND2_X1 U5399 ( .A1(n4368), .A2(n4367), .ZN(n4369) );
  AND2_X1 U5400 ( .A1(n4780), .A2(n4369), .ZN(n6253) );
  NOR2_X1 U5401 ( .A1(n6123), .A2(n6066), .ZN(n4370) );
  AOI21_X1 U5402 ( .B1(n6253), .B2(n6563), .A(n4370), .ZN(n4371) );
  OAI21_X1 U5403 ( .B1(n4407), .B2(n6118), .A(n4371), .ZN(U2853) );
  INV_X1 U5404 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4377) );
  OR2_X1 U5405 ( .A1(n4452), .A2(n4372), .ZN(n4373) );
  NAND2_X1 U5406 ( .A1(n4374), .A2(n4373), .ZN(n4375) );
  NAND2_X1 U5407 ( .A1(n6162), .A2(n5071), .ZN(n6134) );
  NAND2_X1 U5408 ( .A1(n6429), .A2(n5050), .ZN(n6148) );
  INV_X1 U5409 ( .A(n6148), .ZN(n6160) );
  AOI22_X1 U5410 ( .A1(n6160), .A2(UWORD_REG_7__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4376) );
  OAI21_X1 U5411 ( .B1(n4377), .B2(n6134), .A(n4376), .ZN(U2900) );
  AOI22_X1 U5412 ( .A1(n6160), .A2(UWORD_REG_4__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4378) );
  OAI21_X1 U5413 ( .B1(n4379), .B2(n6134), .A(n4378), .ZN(U2903) );
  AOI22_X1 U5414 ( .A1(n6160), .A2(UWORD_REG_8__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4380) );
  OAI21_X1 U5415 ( .B1(n4381), .B2(n6134), .A(n4380), .ZN(U2899) );
  INV_X1 U5416 ( .A(EAX_REG_25__SCAN_IN), .ZN(n6573) );
  AOI22_X1 U5417 ( .A1(n6160), .A2(UWORD_REG_9__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4382) );
  OAI21_X1 U5418 ( .B1(n6573), .B2(n6134), .A(n4382), .ZN(U2898) );
  AOI22_X1 U5419 ( .A1(n6160), .A2(UWORD_REG_3__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4383) );
  OAI21_X1 U5420 ( .B1(n4384), .B2(n6134), .A(n4383), .ZN(U2904) );
  AOI22_X1 U5421 ( .A1(UWORD_REG_11__SCAN_IN), .A2(n6160), .B1(n6163), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4385) );
  OAI21_X1 U5422 ( .B1(n4386), .B2(n6134), .A(n4385), .ZN(U2896) );
  AOI22_X1 U5423 ( .A1(n6160), .A2(UWORD_REG_2__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4387) );
  OAI21_X1 U5424 ( .B1(n4388), .B2(n6134), .A(n4387), .ZN(U2905) );
  AOI22_X1 U5425 ( .A1(n6160), .A2(UWORD_REG_12__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_28__SCAN_IN), .ZN(n4389) );
  OAI21_X1 U5426 ( .B1(n4390), .B2(n6134), .A(n4389), .ZN(U2895) );
  INV_X1 U5427 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4392) );
  AOI22_X1 U5428 ( .A1(n6160), .A2(UWORD_REG_5__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_21__SCAN_IN), .ZN(n4391) );
  OAI21_X1 U5429 ( .B1(n4392), .B2(n6134), .A(n4391), .ZN(U2902) );
  XNOR2_X1 U5430 ( .A(n4394), .B(n4393), .ZN(n4725) );
  INV_X1 U5431 ( .A(n5921), .ZN(n6228) );
  NOR2_X1 U5432 ( .A1(n4395), .A2(n6228), .ZN(n4397) );
  MUX2_X1 U5433 ( .A(n4397), .B(n4396), .S(INSTADDRPOINTER_REG_1__SCAN_IN), 
        .Z(n4398) );
  INV_X1 U5434 ( .A(n4398), .ZN(n4401) );
  AOI22_X1 U5435 ( .A1(n6279), .A2(n4399), .B1(n6260), .B2(REIP_REG_1__SCAN_IN), .ZN(n4400) );
  OAI211_X1 U5436 ( .C1(n4725), .C2(n5906), .A(n4401), .B(n4400), .ZN(U3017)
         );
  AOI22_X1 U5437 ( .A1(n6552), .A2(UWORD_REG_0__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4402) );
  OAI21_X1 U5438 ( .B1(n4403), .B2(n6134), .A(n4402), .ZN(U2907) );
  AOI22_X1 U5439 ( .A1(n6552), .A2(UWORD_REG_1__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4404) );
  OAI21_X1 U5440 ( .B1(n4405), .B2(n6134), .A(n4404), .ZN(U2906) );
  AOI22_X1 U5441 ( .A1(n6552), .A2(UWORD_REG_10__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4406) );
  OAI21_X1 U5442 ( .B1(n6733), .B2(n6134), .A(n4406), .ZN(U2897) );
  OAI222_X1 U5443 ( .A1(n4407), .A2(n5867), .B1(n5088), .B2(n6593), .C1(n5432), 
        .C2(n3397), .ZN(U2885) );
  INV_X1 U5444 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4409) );
  INV_X2 U5445 ( .A(n6145), .ZN(n6163) );
  AOI22_X1 U5446 ( .A1(n6552), .A2(UWORD_REG_13__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4408) );
  OAI21_X1 U5447 ( .B1(n4409), .B2(n6134), .A(n4408), .ZN(U2894) );
  AND2_X1 U5448 ( .A1(n6103), .A2(n3255), .ZN(n4789) );
  NAND2_X1 U5449 ( .A1(n5328), .A2(n4104), .ZN(n6308) );
  INV_X1 U5450 ( .A(n6308), .ZN(n4660) );
  INV_X1 U5451 ( .A(n4440), .ZN(n4410) );
  AOI21_X1 U5452 ( .B1(n4789), .B2(n4660), .A(n4410), .ZN(n4413) );
  INV_X1 U5453 ( .A(n4413), .ZN(n4411) );
  AOI22_X1 U5454 ( .A1(n4411), .A2(n4551), .B1(n4662), .B2(
        STATE2_REG_2__SCAN_IN), .ZN(n4444) );
  INV_X1 U5455 ( .A(n6312), .ZN(n5017) );
  AOI21_X1 U5456 ( .B1(n6406), .B2(STATE2_REG_3__SCAN_IN), .A(n4471), .ZN(
        n4899) );
  INV_X1 U5457 ( .A(n4519), .ZN(n4412) );
  AOI21_X1 U5458 ( .B1(n4412), .B2(n5778), .A(n5679), .ZN(n4414) );
  AND2_X1 U5459 ( .A1(n4551), .A2(n6743), .ZN(n4657) );
  OAI21_X1 U5460 ( .B1(n4414), .B2(n4657), .A(n4413), .ZN(n4415) );
  OAI211_X1 U5461 ( .C1(n4662), .C2(n4551), .A(n4899), .B(n4415), .ZN(n4438)
         );
  NAND2_X1 U5462 ( .A1(n4438), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n4419)
         );
  NAND2_X1 U5463 ( .A1(n5778), .A2(n4892), .ZN(n4947) );
  INV_X1 U5464 ( .A(n4416), .ZN(n4439) );
  OAI22_X1 U5465 ( .A1(n4969), .A2(n4440), .B1(n6324), .B2(n4439), .ZN(n4417)
         );
  AOI21_X1 U5466 ( .B1(n6321), .B2(n4669), .A(n4417), .ZN(n4418) );
  OAI211_X1 U5467 ( .C1(n4444), .C2(n5017), .A(n4419), .B(n4418), .ZN(U3140)
         );
  INV_X1 U5468 ( .A(n6376), .ZN(n4963) );
  NAND2_X1 U5469 ( .A1(n4438), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4422)
         );
  OAI22_X1 U5470 ( .A1(n4959), .A2(n4440), .B1(n6328), .B2(n4439), .ZN(n4420)
         );
  AOI21_X1 U5471 ( .B1(n6325), .B2(n4669), .A(n4420), .ZN(n4421) );
  OAI211_X1 U5472 ( .C1(n4444), .C2(n4963), .A(n4422), .B(n4421), .ZN(U3141)
         );
  INV_X1 U5473 ( .A(n6382), .ZN(n4958) );
  NAND2_X1 U5474 ( .A1(n4438), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4425)
         );
  OAI22_X1 U5475 ( .A1(n4954), .A2(n4440), .B1(n6338), .B2(n4439), .ZN(n4423)
         );
  AOI21_X1 U5476 ( .B1(n6335), .B2(n4669), .A(n4423), .ZN(n4424) );
  OAI211_X1 U5477 ( .C1(n4444), .C2(n4958), .A(n4425), .B(n4424), .ZN(U3143)
         );
  INV_X1 U5478 ( .A(n6340), .ZN(n5023) );
  NAND2_X1 U5479 ( .A1(n4438), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4428)
         );
  OAI22_X1 U5480 ( .A1(n4987), .A2(n4440), .B1(n6344), .B2(n4439), .ZN(n4426)
         );
  AOI21_X1 U5481 ( .B1(n6341), .B2(n4669), .A(n4426), .ZN(n4427) );
  OAI211_X1 U5482 ( .C1(n4444), .C2(n5023), .A(n4428), .B(n4427), .ZN(U3144)
         );
  INV_X1 U5483 ( .A(n6391), .ZN(n4968) );
  NAND2_X1 U5484 ( .A1(n4438), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4431)
         );
  OAI22_X1 U5485 ( .A1(n4964), .A2(n4440), .B1(n6354), .B2(n4439), .ZN(n4429)
         );
  AOI21_X1 U5486 ( .B1(n6351), .B2(n4669), .A(n4429), .ZN(n4430) );
  OAI211_X1 U5487 ( .C1(n4444), .C2(n4968), .A(n4431), .B(n4430), .ZN(U3146)
         );
  INV_X1 U5488 ( .A(n6346), .ZN(n5011) );
  NAND2_X1 U5489 ( .A1(n4438), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4434)
         );
  OAI22_X1 U5490 ( .A1(n4973), .A2(n4440), .B1(n6350), .B2(n4439), .ZN(n4432)
         );
  AOI21_X1 U5491 ( .B1(n6347), .B2(n4669), .A(n4432), .ZN(n4433) );
  OAI211_X1 U5492 ( .C1(n4444), .C2(n5011), .A(n4434), .B(n4433), .ZN(U3145)
         );
  INV_X1 U5493 ( .A(n6330), .ZN(n5029) );
  NAND2_X1 U5494 ( .A1(n4438), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4437)
         );
  OAI22_X1 U5495 ( .A1(n4977), .A2(n4440), .B1(n6334), .B2(n4439), .ZN(n4435)
         );
  AOI21_X1 U5496 ( .B1(n6331), .B2(n4669), .A(n4435), .ZN(n4436) );
  OAI211_X1 U5497 ( .C1(n4444), .C2(n5029), .A(n4437), .B(n4436), .ZN(U3142)
         );
  INV_X1 U5498 ( .A(n6358), .ZN(n5035) );
  NAND2_X1 U5499 ( .A1(n4438), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4443)
         );
  OAI22_X1 U5500 ( .A1(n4981), .A2(n4440), .B1(n6364), .B2(n4439), .ZN(n4441)
         );
  AOI21_X1 U5501 ( .B1(n6360), .B2(n4669), .A(n4441), .ZN(n4442) );
  OAI211_X1 U5502 ( .C1(n4444), .C2(n5035), .A(n4443), .B(n4442), .ZN(U3147)
         );
  INV_X1 U5503 ( .A(n4547), .ZN(n4583) );
  OR2_X1 U5504 ( .A1(n4445), .A2(n4583), .ZN(n4446) );
  XNOR2_X1 U5505 ( .A(n4446), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6082)
         );
  NOR2_X1 U5506 ( .A1(n4063), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4449) );
  NAND2_X1 U5507 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5977), .ZN(n4447) );
  OAI21_X1 U5508 ( .B1(n6398), .B2(STATE2_REG_1__SCAN_IN), .A(n4447), .ZN(
        n4460) );
  AND2_X1 U5509 ( .A1(n4460), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4448)
         );
  AOI21_X1 U5510 ( .B1(n6082), .B2(n4449), .A(n4448), .ZN(n4463) );
  NAND2_X1 U5511 ( .A1(n5328), .A2(n6400), .ZN(n4457) );
  XNOR2_X1 U5512 ( .A(n4067), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4454)
         );
  XNOR2_X1 U5513 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4451) );
  OAI22_X1 U5514 ( .A1(n4452), .A2(n4451), .B1(n4450), .B2(n4454), .ZN(n4453)
         );
  AOI21_X1 U5515 ( .B1(n4455), .B2(n4454), .A(n4453), .ZN(n4456) );
  NAND2_X1 U5516 ( .A1(n4457), .A2(n4456), .ZN(n6399) );
  NAND4_X1 U5517 ( .A1(n6397), .A2(n6532), .A3(n6399), .A4(n6398), .ZN(n4462)
         );
  CLKBUF_X1 U5518 ( .A(n4458), .Z(n4459) );
  NAND2_X1 U5519 ( .A1(n4460), .A2(n4459), .ZN(n4461) );
  AND3_X1 U5520 ( .A1(n4463), .A2(n4462), .A3(n4461), .ZN(n6424) );
  AND2_X1 U5521 ( .A1(n4463), .A2(n4105), .ZN(n4464) );
  AOI21_X1 U5522 ( .B1(n4466), .B2(n5977), .A(n6527), .ZN(n4465) );
  NOR2_X1 U5523 ( .A1(n4612), .A2(n4465), .ZN(n5782) );
  INV_X1 U5524 ( .A(n5782), .ZN(n6292) );
  NAND2_X1 U5525 ( .A1(n4466), .A2(n6429), .ZN(n6434) );
  INV_X1 U5526 ( .A(n6434), .ZN(n4468) );
  INV_X1 U5527 ( .A(n3255), .ZN(n6404) );
  NAND2_X1 U5528 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n3149), .ZN(n5324) );
  INV_X1 U5529 ( .A(n5324), .ZN(n5781) );
  OAI22_X1 U5530 ( .A1(n4892), .A2(n5000), .B1(n6404), .B2(n5781), .ZN(n4467)
         );
  OAI21_X1 U5531 ( .B1(n4468), .B2(n4467), .A(n6292), .ZN(n4469) );
  OAI21_X1 U5532 ( .B1(n6292), .B2(n6406), .A(n4469), .ZN(U3465) );
  NAND3_X1 U5533 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n4787), .ZN(n4522) );
  NOR2_X1 U5534 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4522), .ZN(n4499)
         );
  OR2_X1 U5535 ( .A1(n6305), .A2(n4470), .ZN(n4856) );
  AOI21_X1 U5536 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n4856), .A(n4471), .ZN(
        n4853) );
  OAI211_X1 U5537 ( .C1(n3149), .C2(n4499), .A(n4853), .B(n4944), .ZN(n4476)
         );
  NAND2_X1 U5538 ( .A1(n3348), .A2(n4472), .ZN(n4786) );
  INV_X1 U5539 ( .A(n4786), .ZN(n4651) );
  INV_X1 U5540 ( .A(n5004), .ZN(n4473) );
  NAND2_X1 U5541 ( .A1(n4651), .A2(n4473), .ZN(n4477) );
  OR2_X1 U5542 ( .A1(n4519), .A2(n5778), .ZN(n4518) );
  OR2_X1 U5543 ( .A1(n4518), .A2(n4140), .ZN(n4478) );
  NAND3_X1 U5544 ( .A1(n4477), .A2(n4551), .A3(n4478), .ZN(n4474) );
  INV_X1 U5545 ( .A(n4657), .ZN(n5217) );
  INV_X1 U5546 ( .A(n4104), .ZN(n5780) );
  AND2_X1 U5547 ( .A1(n5328), .A2(n5780), .ZN(n4584) );
  AOI22_X1 U5548 ( .A1(n4474), .A2(n5217), .B1(n4584), .B2(n4547), .ZN(n4475)
         );
  INV_X1 U5549 ( .A(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4481) );
  AOI22_X1 U5550 ( .A1(n6381), .A2(n4499), .B1(n6335), .B2(n6386), .ZN(n4480)
         );
  NOR2_X1 U5551 ( .A1(n5223), .A2(n5000), .ZN(n4661) );
  INV_X1 U5552 ( .A(n4661), .ZN(n4858) );
  INV_X1 U5553 ( .A(n4584), .ZN(n5226) );
  INV_X1 U5554 ( .A(n6306), .ZN(n5225) );
  OAI22_X1 U5555 ( .A1(n4858), .A2(n5226), .B1(n4856), .B2(n5225), .ZN(n4500)
         );
  INV_X1 U5556 ( .A(n6338), .ZN(n6380) );
  AOI22_X1 U5557 ( .A1(n6382), .A2(n4500), .B1(n6380), .B2(n4541), .ZN(n4479)
         );
  OAI211_X1 U5558 ( .C1(n4504), .C2(n4481), .A(n4480), .B(n4479), .ZN(U3119)
         );
  INV_X1 U5559 ( .A(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4484) );
  AOI22_X1 U5560 ( .A1(n6339), .A2(n4499), .B1(n6341), .B2(n6386), .ZN(n4483)
         );
  INV_X1 U5561 ( .A(n6344), .ZN(n5018) );
  AOI22_X1 U5562 ( .A1(n6340), .A2(n4500), .B1(n5018), .B2(n4541), .ZN(n4482)
         );
  OAI211_X1 U5563 ( .C1(n4504), .C2(n4484), .A(n4483), .B(n4482), .ZN(U3120)
         );
  INV_X1 U5564 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4487) );
  AOI22_X1 U5565 ( .A1(n6329), .A2(n4499), .B1(n6331), .B2(n6386), .ZN(n4486)
         );
  INV_X1 U5566 ( .A(n6334), .ZN(n5024) );
  AOI22_X1 U5567 ( .A1(n6330), .A2(n4500), .B1(n5024), .B2(n4541), .ZN(n4485)
         );
  OAI211_X1 U5568 ( .C1(n4504), .C2(n4487), .A(n4486), .B(n4485), .ZN(U3118)
         );
  AOI22_X1 U5569 ( .A1(n6389), .A2(n4499), .B1(n6351), .B2(n6386), .ZN(n4489)
         );
  INV_X1 U5570 ( .A(n6354), .ZN(n6387) );
  AOI22_X1 U5571 ( .A1(n6391), .A2(n4500), .B1(n6387), .B2(n4541), .ZN(n4488)
         );
  OAI211_X1 U5572 ( .C1(n4504), .C2(n6602), .A(n4489), .B(n4488), .ZN(U3122)
         );
  INV_X1 U5573 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4492) );
  AOI22_X1 U5574 ( .A1(n6311), .A2(n4499), .B1(n6321), .B2(n6386), .ZN(n4491)
         );
  INV_X1 U5575 ( .A(n6324), .ZN(n5012) );
  AOI22_X1 U5576 ( .A1(n6312), .A2(n4500), .B1(n5012), .B2(n4541), .ZN(n4490)
         );
  OAI211_X1 U5577 ( .C1(n4504), .C2(n4492), .A(n4491), .B(n4490), .ZN(U3116)
         );
  INV_X1 U5578 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4495) );
  AOI22_X1 U5579 ( .A1(n6345), .A2(n4499), .B1(n6347), .B2(n6386), .ZN(n4494)
         );
  INV_X1 U5580 ( .A(n6350), .ZN(n5006) );
  AOI22_X1 U5581 ( .A1(n6346), .A2(n4500), .B1(n5006), .B2(n4541), .ZN(n4493)
         );
  OAI211_X1 U5582 ( .C1(n4504), .C2(n4495), .A(n4494), .B(n4493), .ZN(U3121)
         );
  INV_X1 U5583 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4498) );
  AOI22_X1 U5584 ( .A1(n6356), .A2(n4499), .B1(n6360), .B2(n6386), .ZN(n4497)
         );
  INV_X1 U5585 ( .A(n6364), .ZN(n5030) );
  AOI22_X1 U5586 ( .A1(n6358), .A2(n4500), .B1(n5030), .B2(n4541), .ZN(n4496)
         );
  OAI211_X1 U5587 ( .C1(n4504), .C2(n4498), .A(n4497), .B(n4496), .ZN(U3123)
         );
  INV_X1 U5588 ( .A(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4503) );
  AOI22_X1 U5589 ( .A1(n6375), .A2(n4499), .B1(n6325), .B2(n6386), .ZN(n4502)
         );
  INV_X1 U5590 ( .A(n6328), .ZN(n6374) );
  AOI22_X1 U5591 ( .A1(n6376), .A2(n4500), .B1(n6374), .B2(n4541), .ZN(n4501)
         );
  OAI211_X1 U5592 ( .C1(n4504), .C2(n4503), .A(n4502), .B(n4501), .ZN(U3117)
         );
  INV_X1 U5593 ( .A(n4505), .ZN(n4516) );
  INV_X1 U5594 ( .A(n6181), .ZN(n6204) );
  OR2_X1 U5595 ( .A1(n4509), .A2(n4551), .ZN(n6550) );
  NAND2_X1 U5596 ( .A1(n6550), .A2(n5050), .ZN(n4510) );
  NAND2_X1 U5597 ( .A1(n5050), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4512) );
  NAND2_X1 U5598 ( .A1(n6743), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4511) );
  AND2_X1 U5599 ( .A1(n4512), .A2(n4511), .ZN(n4721) );
  INV_X1 U5600 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n4513) );
  AOI21_X1 U5601 ( .B1(n5651), .B2(n4721), .A(n4513), .ZN(n4514) );
  AOI211_X1 U5602 ( .C1(n4516), .C2(n6204), .A(n4515), .B(n4514), .ZN(n4517)
         );
  OAI21_X1 U5603 ( .B1(n5080), .B2(n5679), .A(n4517), .ZN(U2986) );
  NOR2_X1 U5604 ( .A1(n6406), .A2(n4522), .ZN(n4542) );
  AOI21_X1 U5605 ( .B1(n4789), .B2(n4584), .A(n4542), .ZN(n4524) );
  OR2_X1 U5606 ( .A1(n5778), .A2(n6743), .ZN(n4785) );
  NOR2_X1 U5607 ( .A1(n4519), .A2(n4785), .ZN(n4652) );
  NOR2_X1 U5608 ( .A1(n4652), .A2(n5000), .ZN(n4521) );
  AOI22_X1 U5609 ( .A1(n4524), .A2(n4521), .B1(n5000), .B2(n4522), .ZN(n4520)
         );
  NAND2_X1 U5610 ( .A1(n4899), .A2(n4520), .ZN(n4540) );
  INV_X1 U5611 ( .A(n4521), .ZN(n4523) );
  OAI22_X1 U5612 ( .A1(n4524), .A2(n4523), .B1(n6433), .B2(n4522), .ZN(n4539)
         );
  AOI22_X1 U5613 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4540), .B1(n6382), 
        .B2(n4539), .ZN(n4526) );
  AOI22_X1 U5614 ( .A1(n6381), .A2(n4542), .B1(n6335), .B2(n4541), .ZN(n4525)
         );
  OAI211_X1 U5615 ( .C1(n6338), .C2(n4664), .A(n4526), .B(n4525), .ZN(U3127)
         );
  AOI22_X1 U5616 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4540), .B1(n6340), 
        .B2(n4539), .ZN(n4528) );
  AOI22_X1 U5617 ( .A1(n6339), .A2(n4542), .B1(n6341), .B2(n4541), .ZN(n4527)
         );
  OAI211_X1 U5618 ( .C1(n6344), .C2(n4664), .A(n4528), .B(n4527), .ZN(U3128)
         );
  AOI22_X1 U5619 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4540), .B1(n6346), 
        .B2(n4539), .ZN(n4530) );
  AOI22_X1 U5620 ( .A1(n6345), .A2(n4542), .B1(n6347), .B2(n4541), .ZN(n4529)
         );
  OAI211_X1 U5621 ( .C1(n6350), .C2(n4664), .A(n4530), .B(n4529), .ZN(U3129)
         );
  AOI22_X1 U5622 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4540), .B1(n6358), 
        .B2(n4539), .ZN(n4532) );
  AOI22_X1 U5623 ( .A1(n6356), .A2(n4542), .B1(n6360), .B2(n4541), .ZN(n4531)
         );
  OAI211_X1 U5624 ( .C1(n6364), .C2(n4664), .A(n4532), .B(n4531), .ZN(U3131)
         );
  AOI22_X1 U5625 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4540), .B1(n6391), 
        .B2(n4539), .ZN(n4534) );
  AOI22_X1 U5626 ( .A1(n6389), .A2(n4542), .B1(n6351), .B2(n4541), .ZN(n4533)
         );
  OAI211_X1 U5627 ( .C1(n6354), .C2(n4664), .A(n4534), .B(n4533), .ZN(U3130)
         );
  AOI22_X1 U5628 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4540), .B1(n6312), 
        .B2(n4539), .ZN(n4536) );
  AOI22_X1 U5629 ( .A1(n6311), .A2(n4542), .B1(n6321), .B2(n4541), .ZN(n4535)
         );
  OAI211_X1 U5630 ( .C1(n6324), .C2(n4664), .A(n4536), .B(n4535), .ZN(U3124)
         );
  AOI22_X1 U5631 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4540), .B1(n6330), 
        .B2(n4539), .ZN(n4538) );
  AOI22_X1 U5632 ( .A1(n6329), .A2(n4542), .B1(n6331), .B2(n4541), .ZN(n4537)
         );
  OAI211_X1 U5633 ( .C1(n6334), .C2(n4664), .A(n4538), .B(n4537), .ZN(U3126)
         );
  AOI22_X1 U5634 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4540), .B1(n6376), 
        .B2(n4539), .ZN(n4544) );
  AOI22_X1 U5635 ( .A1(n6375), .A2(n4542), .B1(n6325), .B2(n4541), .ZN(n4543)
         );
  OAI211_X1 U5636 ( .C1(n6328), .C2(n4664), .A(n4544), .B(n4543), .ZN(U3125)
         );
  INV_X1 U5637 ( .A(n4545), .ZN(n4546) );
  NAND2_X1 U5638 ( .A1(n3015), .A2(n4546), .ZN(n4580) );
  NAND2_X1 U5639 ( .A1(n5778), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5777) );
  OR2_X1 U5640 ( .A1(n4580), .A2(n5777), .ZN(n4649) );
  NAND2_X1 U5641 ( .A1(n4649), .A2(n4551), .ZN(n4552) );
  OR2_X1 U5642 ( .A1(n6308), .A2(n4547), .ZN(n6314) );
  OR2_X1 U5643 ( .A1(n6314), .A2(n6404), .ZN(n4548) );
  AND2_X1 U5644 ( .A1(n4548), .A2(n6365), .ZN(n4553) );
  OR2_X1 U5645 ( .A1(n4552), .A2(n4553), .ZN(n4550) );
  NAND2_X1 U5646 ( .A1(STATE2_REG_2__SCAN_IN), .A2(n6310), .ZN(n4549) );
  NAND2_X1 U5647 ( .A1(n4550), .A2(n4549), .ZN(n6369) );
  INV_X1 U5648 ( .A(n4552), .ZN(n4554) );
  NAND2_X1 U5649 ( .A1(n4554), .A2(n4553), .ZN(n4555) );
  OAI211_X1 U5650 ( .C1(n6310), .C2(n4551), .A(n4899), .B(n4555), .ZN(n6370)
         );
  NAND2_X1 U5651 ( .A1(n6370), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4559) );
  INV_X1 U5652 ( .A(n4580), .ZN(n4582) );
  INV_X1 U5653 ( .A(n4947), .ZN(n4556) );
  NAND2_X1 U5654 ( .A1(n4582), .A2(n4556), .ZN(n6373) );
  INV_X1 U5655 ( .A(n6373), .ZN(n4576) );
  OAI22_X1 U5656 ( .A1(n4954), .A2(n6365), .B1(n6338), .B2(n6366), .ZN(n4557)
         );
  AOI21_X1 U5657 ( .B1(n6335), .B2(n4576), .A(n4557), .ZN(n4558) );
  OAI211_X1 U5658 ( .C1(n4579), .C2(n4958), .A(n4559), .B(n4558), .ZN(U3079)
         );
  NAND2_X1 U5659 ( .A1(n6370), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4562) );
  OAI22_X1 U5660 ( .A1(n4969), .A2(n6365), .B1(n6324), .B2(n6366), .ZN(n4560)
         );
  AOI21_X1 U5661 ( .B1(n6321), .B2(n4576), .A(n4560), .ZN(n4561) );
  OAI211_X1 U5662 ( .C1(n4579), .C2(n5017), .A(n4562), .B(n4561), .ZN(U3076)
         );
  NAND2_X1 U5663 ( .A1(n6370), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4565) );
  OAI22_X1 U5664 ( .A1(n4987), .A2(n6365), .B1(n6344), .B2(n6366), .ZN(n4563)
         );
  AOI21_X1 U5665 ( .B1(n6341), .B2(n4576), .A(n4563), .ZN(n4564) );
  OAI211_X1 U5666 ( .C1(n4579), .C2(n5023), .A(n4565), .B(n4564), .ZN(U3080)
         );
  NAND2_X1 U5667 ( .A1(n6370), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4568) );
  OAI22_X1 U5668 ( .A1(n4977), .A2(n6365), .B1(n6334), .B2(n6366), .ZN(n4566)
         );
  AOI21_X1 U5669 ( .B1(n6331), .B2(n4576), .A(n4566), .ZN(n4567) );
  OAI211_X1 U5670 ( .C1(n4579), .C2(n5029), .A(n4568), .B(n4567), .ZN(U3078)
         );
  NAND2_X1 U5671 ( .A1(n6370), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4571) );
  OAI22_X1 U5672 ( .A1(n4973), .A2(n6365), .B1(n6350), .B2(n6366), .ZN(n4569)
         );
  AOI21_X1 U5673 ( .B1(n6347), .B2(n4576), .A(n4569), .ZN(n4570) );
  OAI211_X1 U5674 ( .C1(n4579), .C2(n5011), .A(n4571), .B(n4570), .ZN(U3081)
         );
  NAND2_X1 U5675 ( .A1(n6370), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4574) );
  OAI22_X1 U5676 ( .A1(n4981), .A2(n6365), .B1(n6364), .B2(n6366), .ZN(n4572)
         );
  AOI21_X1 U5677 ( .B1(n6360), .B2(n4576), .A(n4572), .ZN(n4573) );
  OAI211_X1 U5678 ( .C1(n4579), .C2(n5035), .A(n4574), .B(n4573), .ZN(U3083)
         );
  NAND2_X1 U5679 ( .A1(n6370), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4578) );
  OAI22_X1 U5680 ( .A1(n4964), .A2(n6365), .B1(n6354), .B2(n6366), .ZN(n4575)
         );
  AOI21_X1 U5681 ( .B1(n6351), .B2(n4576), .A(n4575), .ZN(n4577) );
  OAI211_X1 U5682 ( .C1(n4579), .C2(n4968), .A(n4578), .B(n4577), .ZN(U3082)
         );
  INV_X1 U5683 ( .A(n6321), .ZN(n5014) );
  NOR2_X1 U5684 ( .A1(n4580), .A2(n5778), .ZN(n4590) );
  INV_X1 U5685 ( .A(n4785), .ZN(n4581) );
  AOI21_X1 U5686 ( .B1(n4582), .B2(n4581), .A(n5000), .ZN(n4587) );
  INV_X1 U5687 ( .A(n4587), .ZN(n4585) );
  AND2_X1 U5688 ( .A1(n4584), .A2(n4583), .ZN(n5216) );
  NAND3_X1 U5689 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6718), .A3(n4787), .ZN(n5219) );
  NOR2_X1 U5690 ( .A1(n6406), .A2(n5219), .ZN(n4607) );
  AOI21_X1 U5691 ( .B1(n5216), .B2(n3255), .A(n4607), .ZN(n4586) );
  OAI22_X1 U5692 ( .A1(n4585), .A2(n4586), .B1(n5219), .B2(n6433), .ZN(n4606)
         );
  INV_X1 U5693 ( .A(n5219), .ZN(n4589) );
  NAND2_X1 U5694 ( .A1(n4587), .A2(n4586), .ZN(n4588) );
  OAI211_X1 U5695 ( .C1(n4551), .C2(n4589), .A(n4588), .B(n4899), .ZN(n4605)
         );
  AOI22_X1 U5696 ( .A1(n6312), .A2(n4606), .B1(INSTQUEUE_REG_5__0__SCAN_IN), 
        .B2(n4605), .ZN(n4592) );
  NAND2_X1 U5697 ( .A1(n4590), .A2(n4140), .ZN(n6313) );
  AOI22_X1 U5698 ( .A1(n6311), .A2(n4607), .B1(n5012), .B2(n6359), .ZN(n4591)
         );
  OAI211_X1 U5699 ( .C1(n5014), .C2(n5257), .A(n4592), .B(n4591), .ZN(U3060)
         );
  AOI22_X1 U5700 ( .A1(n6382), .A2(n4606), .B1(INSTQUEUE_REG_5__3__SCAN_IN), 
        .B2(n4605), .ZN(n4594) );
  AOI22_X1 U5701 ( .A1(n6381), .A2(n4607), .B1(n6380), .B2(n6359), .ZN(n4593)
         );
  OAI211_X1 U5702 ( .C1(n6385), .C2(n5257), .A(n4594), .B(n4593), .ZN(U3063)
         );
  AOI22_X1 U5703 ( .A1(n6376), .A2(n4606), .B1(INSTQUEUE_REG_5__1__SCAN_IN), 
        .B2(n4605), .ZN(n4596) );
  AOI22_X1 U5704 ( .A1(n6375), .A2(n4607), .B1(n6374), .B2(n6359), .ZN(n4595)
         );
  OAI211_X1 U5705 ( .C1(n6379), .C2(n5257), .A(n4596), .B(n4595), .ZN(U3061)
         );
  INV_X1 U5706 ( .A(n6347), .ZN(n5008) );
  AOI22_X1 U5707 ( .A1(n6346), .A2(n4606), .B1(INSTQUEUE_REG_5__5__SCAN_IN), 
        .B2(n4605), .ZN(n4598) );
  AOI22_X1 U5708 ( .A1(n6345), .A2(n4607), .B1(n5006), .B2(n6359), .ZN(n4597)
         );
  OAI211_X1 U5709 ( .C1(n5008), .C2(n5257), .A(n4598), .B(n4597), .ZN(U3065)
         );
  INV_X1 U5710 ( .A(n6360), .ZN(n5032) );
  AOI22_X1 U5711 ( .A1(n6358), .A2(n4606), .B1(INSTQUEUE_REG_5__7__SCAN_IN), 
        .B2(n4605), .ZN(n4600) );
  AOI22_X1 U5712 ( .A1(n6356), .A2(n4607), .B1(n5030), .B2(n6359), .ZN(n4599)
         );
  OAI211_X1 U5713 ( .C1(n5032), .C2(n5257), .A(n4600), .B(n4599), .ZN(U3067)
         );
  AOI22_X1 U5714 ( .A1(n6391), .A2(n4606), .B1(INSTQUEUE_REG_5__6__SCAN_IN), 
        .B2(n4605), .ZN(n4602) );
  AOI22_X1 U5715 ( .A1(n6389), .A2(n4607), .B1(n6387), .B2(n6359), .ZN(n4601)
         );
  OAI211_X1 U5716 ( .C1(n6396), .C2(n5257), .A(n4602), .B(n4601), .ZN(U3066)
         );
  INV_X1 U5717 ( .A(n6331), .ZN(n5026) );
  AOI22_X1 U5718 ( .A1(n6330), .A2(n4606), .B1(INSTQUEUE_REG_5__2__SCAN_IN), 
        .B2(n4605), .ZN(n4604) );
  AOI22_X1 U5719 ( .A1(n6329), .A2(n4607), .B1(n5024), .B2(n6359), .ZN(n4603)
         );
  OAI211_X1 U5720 ( .C1(n5026), .C2(n5257), .A(n4604), .B(n4603), .ZN(U3062)
         );
  INV_X1 U5721 ( .A(n6341), .ZN(n5020) );
  AOI22_X1 U5722 ( .A1(n6340), .A2(n4606), .B1(INSTQUEUE_REG_5__4__SCAN_IN), 
        .B2(n4605), .ZN(n4609) );
  AOI22_X1 U5723 ( .A1(n6339), .A2(n4607), .B1(n5018), .B2(n6359), .ZN(n4608)
         );
  OAI211_X1 U5724 ( .C1(n5020), .C2(n5257), .A(n4609), .B(n4608), .ZN(U3064)
         );
  NAND2_X1 U5725 ( .A1(n4617), .A2(n6395), .ZN(n4610) );
  AOI21_X1 U5726 ( .B1(n4610), .B2(STATEBS16_REG_SCAN_IN), .A(n5000), .ZN(
        n4615) );
  NOR2_X1 U5727 ( .A1(n5328), .A2(n5780), .ZN(n4943) );
  AND2_X1 U5728 ( .A1(n4943), .A2(n6103), .ZN(n4699) );
  NOR2_X1 U5729 ( .A1(n4944), .A2(n6718), .ZN(n4611) );
  AOI22_X1 U5730 ( .A1(n4615), .A2(n4699), .B1(n6305), .B2(n4611), .ZN(n4645)
         );
  OAI21_X1 U5731 ( .B1(n6305), .B2(n6433), .A(n4612), .ZN(n6315) );
  NOR2_X1 U5732 ( .A1(n6306), .A2(n6315), .ZN(n4951) );
  INV_X1 U5733 ( .A(n4699), .ZN(n4614) );
  NAND3_X1 U5734 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n4946), .ZN(n4701) );
  NOR2_X1 U5735 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4701), .ZN(n4618)
         );
  NOR2_X1 U5736 ( .A1(n4618), .A2(n3149), .ZN(n4613) );
  AOI21_X1 U5737 ( .B1(n4615), .B2(n4614), .A(n4613), .ZN(n4616) );
  OAI211_X1 U5738 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6433), .A(n4951), .B(n4616), .ZN(n4640) );
  NAND2_X1 U5739 ( .A1(n4640), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4621)
         );
  INV_X1 U5740 ( .A(n4618), .ZN(n4641) );
  OAI22_X1 U5741 ( .A1(n4973), .A2(n4641), .B1(n6395), .B2(n6350), .ZN(n4619)
         );
  AOI21_X1 U5742 ( .B1(n4810), .B2(n6347), .A(n4619), .ZN(n4620) );
  OAI211_X1 U5743 ( .C1(n4645), .C2(n5011), .A(n4621), .B(n4620), .ZN(U3105)
         );
  NAND2_X1 U5744 ( .A1(n4640), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4624)
         );
  OAI22_X1 U5745 ( .A1(n4987), .A2(n4641), .B1(n6395), .B2(n6344), .ZN(n4622)
         );
  AOI21_X1 U5746 ( .B1(n4810), .B2(n6341), .A(n4622), .ZN(n4623) );
  OAI211_X1 U5747 ( .C1(n4645), .C2(n5023), .A(n4624), .B(n4623), .ZN(U3104)
         );
  NAND2_X1 U5748 ( .A1(n4640), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4627)
         );
  OAI22_X1 U5749 ( .A1(n4969), .A2(n4641), .B1(n6395), .B2(n6324), .ZN(n4625)
         );
  AOI21_X1 U5750 ( .B1(n4810), .B2(n6321), .A(n4625), .ZN(n4626) );
  OAI211_X1 U5751 ( .C1(n4645), .C2(n5017), .A(n4627), .B(n4626), .ZN(U3100)
         );
  NAND2_X1 U5752 ( .A1(n4640), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4630)
         );
  OAI22_X1 U5753 ( .A1(n4964), .A2(n4641), .B1(n6395), .B2(n6354), .ZN(n4628)
         );
  AOI21_X1 U5754 ( .B1(n4810), .B2(n6351), .A(n4628), .ZN(n4629) );
  OAI211_X1 U5755 ( .C1(n4645), .C2(n4968), .A(n4630), .B(n4629), .ZN(U3106)
         );
  NAND2_X1 U5756 ( .A1(n4640), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4633)
         );
  OAI22_X1 U5757 ( .A1(n4981), .A2(n4641), .B1(n6395), .B2(n6364), .ZN(n4631)
         );
  AOI21_X1 U5758 ( .B1(n4810), .B2(n6360), .A(n4631), .ZN(n4632) );
  OAI211_X1 U5759 ( .C1(n4645), .C2(n5035), .A(n4633), .B(n4632), .ZN(U3107)
         );
  NAND2_X1 U5760 ( .A1(n4640), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4636)
         );
  OAI22_X1 U5761 ( .A1(n4977), .A2(n4641), .B1(n6395), .B2(n6334), .ZN(n4634)
         );
  AOI21_X1 U5762 ( .B1(n4810), .B2(n6331), .A(n4634), .ZN(n4635) );
  OAI211_X1 U5763 ( .C1(n4645), .C2(n5029), .A(n4636), .B(n4635), .ZN(U3102)
         );
  NAND2_X1 U5764 ( .A1(n4640), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4639)
         );
  OAI22_X1 U5765 ( .A1(n4959), .A2(n4641), .B1(n6395), .B2(n6328), .ZN(n4637)
         );
  AOI21_X1 U5766 ( .B1(n4810), .B2(n6325), .A(n4637), .ZN(n4638) );
  OAI211_X1 U5767 ( .C1(n4645), .C2(n4963), .A(n4639), .B(n4638), .ZN(U3101)
         );
  NAND2_X1 U5768 ( .A1(n4640), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4644)
         );
  OAI22_X1 U5769 ( .A1(n4954), .A2(n4641), .B1(n6395), .B2(n6338), .ZN(n4642)
         );
  AOI21_X1 U5770 ( .B1(n4810), .B2(n6335), .A(n4642), .ZN(n4643) );
  OAI211_X1 U5771 ( .C1(n4645), .C2(n4958), .A(n4644), .B(n4643), .ZN(U3103)
         );
  XOR2_X1 U5772 ( .A(n4647), .B(n4646), .Z(n5154) );
  INV_X1 U5773 ( .A(n5154), .ZN(n4782) );
  AOI22_X1 U5774 ( .A1(n5301), .A2(DATAI_7_), .B1(n6130), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n4648) );
  OAI21_X1 U5775 ( .B1(n4782), .B2(n5867), .A(n4648), .ZN(U2884) );
  NAND2_X1 U5776 ( .A1(n6103), .A2(n5324), .ZN(n4655) );
  INV_X1 U5777 ( .A(n4649), .ZN(n4650) );
  NOR3_X1 U5778 ( .A1(n4652), .A2(n4651), .A3(n4650), .ZN(n4653) );
  NOR2_X1 U5779 ( .A1(n4653), .A2(n5000), .ZN(n4993) );
  NOR2_X1 U5780 ( .A1(n5782), .A2(n4993), .ZN(n4654) );
  NAND2_X1 U5781 ( .A1(n4655), .A2(n4654), .ZN(n4656) );
  AOI21_X1 U5782 ( .B1(n3348), .B2(n4657), .A(n4656), .ZN(n4658) );
  AOI21_X1 U5783 ( .B1(n5782), .B2(n6718), .A(n4658), .ZN(U3462) );
  NOR2_X1 U5784 ( .A1(n5225), .A2(n6718), .ZN(n4659) );
  AOI22_X1 U5785 ( .A1(n4661), .A2(n4660), .B1(n6305), .B2(n4659), .ZN(n4698)
         );
  INV_X1 U5786 ( .A(n4662), .ZN(n4663) );
  NOR2_X1 U5787 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4663), .ZN(n4668)
         );
  NOR3_X1 U5788 ( .A1(n6315), .A2(n6718), .A3(n6316), .ZN(n4667) );
  OAI21_X1 U5789 ( .B1(n4695), .B2(n4669), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n4665) );
  NAND3_X1 U5790 ( .A1(n6308), .A2(n4551), .A3(n4665), .ZN(n4666) );
  OAI211_X1 U5791 ( .C1(n4668), .C2(n3149), .A(n4667), .B(n4666), .ZN(n4691)
         );
  NAND2_X1 U5792 ( .A1(n4691), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4672)
         );
  INV_X1 U5793 ( .A(n4668), .ZN(n4693) );
  INV_X1 U5794 ( .A(n4669), .ZN(n4692) );
  OAI22_X1 U5795 ( .A1(n4954), .A2(n4693), .B1(n6338), .B2(n4692), .ZN(n4670)
         );
  AOI21_X1 U5796 ( .B1(n6335), .B2(n4695), .A(n4670), .ZN(n4671) );
  OAI211_X1 U5797 ( .C1(n4698), .C2(n4958), .A(n4672), .B(n4671), .ZN(U3135)
         );
  NAND2_X1 U5798 ( .A1(n4691), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4675)
         );
  OAI22_X1 U5799 ( .A1(n4964), .A2(n4693), .B1(n6354), .B2(n4692), .ZN(n4673)
         );
  AOI21_X1 U5800 ( .B1(n6351), .B2(n4695), .A(n4673), .ZN(n4674) );
  OAI211_X1 U5801 ( .C1(n4698), .C2(n4968), .A(n4675), .B(n4674), .ZN(U3138)
         );
  NAND2_X1 U5802 ( .A1(n4691), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4678)
         );
  OAI22_X1 U5803 ( .A1(n4987), .A2(n4693), .B1(n6344), .B2(n4692), .ZN(n4676)
         );
  AOI21_X1 U5804 ( .B1(n6341), .B2(n4695), .A(n4676), .ZN(n4677) );
  OAI211_X1 U5805 ( .C1(n4698), .C2(n5023), .A(n4678), .B(n4677), .ZN(U3136)
         );
  NAND2_X1 U5806 ( .A1(n4691), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4681)
         );
  OAI22_X1 U5807 ( .A1(n4973), .A2(n4693), .B1(n6350), .B2(n4692), .ZN(n4679)
         );
  AOI21_X1 U5808 ( .B1(n6347), .B2(n4695), .A(n4679), .ZN(n4680) );
  OAI211_X1 U5809 ( .C1(n4698), .C2(n5011), .A(n4681), .B(n4680), .ZN(U3137)
         );
  NAND2_X1 U5810 ( .A1(n4691), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4684)
         );
  OAI22_X1 U5811 ( .A1(n4977), .A2(n4693), .B1(n6334), .B2(n4692), .ZN(n4682)
         );
  AOI21_X1 U5812 ( .B1(n6331), .B2(n4695), .A(n4682), .ZN(n4683) );
  OAI211_X1 U5813 ( .C1(n4698), .C2(n5029), .A(n4684), .B(n4683), .ZN(U3134)
         );
  NAND2_X1 U5814 ( .A1(n4691), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4687)
         );
  OAI22_X1 U5815 ( .A1(n4959), .A2(n4693), .B1(n6328), .B2(n4692), .ZN(n4685)
         );
  AOI21_X1 U5816 ( .B1(n6325), .B2(n4695), .A(n4685), .ZN(n4686) );
  OAI211_X1 U5817 ( .C1(n4698), .C2(n4963), .A(n4687), .B(n4686), .ZN(U3133)
         );
  NAND2_X1 U5818 ( .A1(n4691), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4690)
         );
  OAI22_X1 U5819 ( .A1(n4981), .A2(n4693), .B1(n6364), .B2(n4692), .ZN(n4688)
         );
  AOI21_X1 U5820 ( .B1(n6360), .B2(n4695), .A(n4688), .ZN(n4689) );
  OAI211_X1 U5821 ( .C1(n4698), .C2(n5035), .A(n4690), .B(n4689), .ZN(U3139)
         );
  NAND2_X1 U5822 ( .A1(n4691), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4697)
         );
  OAI22_X1 U5823 ( .A1(n4969), .A2(n4693), .B1(n6324), .B2(n4692), .ZN(n4694)
         );
  AOI21_X1 U5824 ( .B1(n6321), .B2(n4695), .A(n4694), .ZN(n4696) );
  OAI211_X1 U5825 ( .C1(n4698), .C2(n5017), .A(n4697), .B(n4696), .ZN(U3132)
         );
  OAI21_X1 U5826 ( .B1(n4786), .B2(n5777), .A(n4551), .ZN(n4704) );
  NOR2_X1 U5827 ( .A1(n4995), .A2(n6718), .ZN(n6388) );
  AOI21_X1 U5828 ( .B1(n4699), .B2(n3255), .A(n6388), .ZN(n4700) );
  OAI22_X1 U5829 ( .A1(n4704), .A2(n4700), .B1(n4701), .B2(n6433), .ZN(n6390)
         );
  INV_X1 U5830 ( .A(n6390), .ZN(n4720) );
  INV_X1 U5831 ( .A(n4700), .ZN(n4703) );
  INV_X1 U5832 ( .A(n4899), .ZN(n4998) );
  AOI21_X1 U5833 ( .B1(n5000), .B2(n4701), .A(n4998), .ZN(n4702) );
  OAI21_X1 U5834 ( .B1(n4704), .B2(n4703), .A(n4702), .ZN(n6392) );
  AOI22_X1 U5835 ( .A1(n6339), .A2(n6388), .B1(n5018), .B2(n6386), .ZN(n4705)
         );
  OAI21_X1 U5836 ( .B1(n6395), .B2(n5020), .A(n4705), .ZN(n4706) );
  AOI21_X1 U5837 ( .B1(INSTQUEUE_REG_11__4__SCAN_IN), .B2(n6392), .A(n4706), 
        .ZN(n4707) );
  OAI21_X1 U5838 ( .B1(n4720), .B2(n5023), .A(n4707), .ZN(U3112) );
  AOI22_X1 U5839 ( .A1(n6329), .A2(n6388), .B1(n5024), .B2(n6386), .ZN(n4708)
         );
  OAI21_X1 U5840 ( .B1(n6395), .B2(n5026), .A(n4708), .ZN(n4709) );
  AOI21_X1 U5841 ( .B1(INSTQUEUE_REG_11__2__SCAN_IN), .B2(n6392), .A(n4709), 
        .ZN(n4710) );
  OAI21_X1 U5842 ( .B1(n4720), .B2(n5029), .A(n4710), .ZN(U3110) );
  AOI22_X1 U5843 ( .A1(n6311), .A2(n6388), .B1(n5012), .B2(n6386), .ZN(n4711)
         );
  OAI21_X1 U5844 ( .B1(n6395), .B2(n5014), .A(n4711), .ZN(n4712) );
  AOI21_X1 U5845 ( .B1(INSTQUEUE_REG_11__0__SCAN_IN), .B2(n6392), .A(n4712), 
        .ZN(n4713) );
  OAI21_X1 U5846 ( .B1(n4720), .B2(n5017), .A(n4713), .ZN(U3108) );
  AOI22_X1 U5847 ( .A1(n6356), .A2(n6388), .B1(n5030), .B2(n6386), .ZN(n4714)
         );
  OAI21_X1 U5848 ( .B1(n6395), .B2(n5032), .A(n4714), .ZN(n4715) );
  AOI21_X1 U5849 ( .B1(INSTQUEUE_REG_11__7__SCAN_IN), .B2(n6392), .A(n4715), 
        .ZN(n4716) );
  OAI21_X1 U5850 ( .B1(n4720), .B2(n5035), .A(n4716), .ZN(U3115) );
  AOI22_X1 U5851 ( .A1(n6345), .A2(n6388), .B1(n5006), .B2(n6386), .ZN(n4717)
         );
  OAI21_X1 U5852 ( .B1(n6395), .B2(n5008), .A(n4717), .ZN(n4718) );
  AOI21_X1 U5853 ( .B1(INSTQUEUE_REG_11__5__SCAN_IN), .B2(n6392), .A(n4718), 
        .ZN(n4719) );
  OAI21_X1 U5854 ( .B1(n4720), .B2(n5011), .A(n4719), .ZN(U3113) );
  AOI22_X1 U5855 ( .A1(n6199), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n6260), 
        .B2(REIP_REG_1__SCAN_IN), .ZN(n4722) );
  OAI21_X1 U5856 ( .B1(n6210), .B2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4722), 
        .ZN(n4723) );
  AOI21_X1 U5857 ( .B1(n5504), .B2(n6205), .A(n4723), .ZN(n4724) );
  OAI21_X1 U5858 ( .B1(n4725), .B2(n6181), .A(n4724), .ZN(U2985) );
  INV_X1 U5859 ( .A(n5122), .ZN(n4729) );
  INV_X1 U5860 ( .A(n5114), .ZN(n4727) );
  AOI22_X1 U5861 ( .A1(n6199), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .B1(n6260), 
        .B2(REIP_REG_5__SCAN_IN), .ZN(n4726) );
  OAI21_X1 U5862 ( .B1(n6210), .B2(n4727), .A(n4726), .ZN(n4728) );
  AOI21_X1 U5863 ( .B1(n4729), .B2(n6205), .A(n4728), .ZN(n4730) );
  OAI21_X1 U5864 ( .B1(n4731), .B2(n6181), .A(n4730), .ZN(U2981) );
  OAI21_X1 U5865 ( .B1(n4732), .B2(n4734), .A(n4733), .ZN(n6269) );
  INV_X1 U5866 ( .A(n6109), .ZN(n4736) );
  AND2_X1 U5867 ( .A1(n6260), .A2(REIP_REG_3__SCAN_IN), .ZN(n6267) );
  AOI21_X1 U5868 ( .B1(n6199), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n6267), 
        .ZN(n4735) );
  OAI21_X1 U5869 ( .B1(n6210), .B2(n4736), .A(n4735), .ZN(n4737) );
  AOI21_X1 U5870 ( .B1(n4738), .B2(n6205), .A(n4737), .ZN(n4739) );
  OAI21_X1 U5871 ( .B1(n6181), .B2(n6269), .A(n4739), .ZN(U2983) );
  NAND2_X1 U5872 ( .A1(n4740), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4741)
         );
  NAND2_X1 U5873 ( .A1(n4742), .A2(n4741), .ZN(n6185) );
  NAND3_X1 U5874 ( .A1(n4821), .A2(n4753), .A3(n4743), .ZN(n4750) );
  NAND2_X1 U5875 ( .A1(n4745), .A2(n4744), .ZN(n4746) );
  OR2_X1 U5876 ( .A1(n4747), .A2(n4746), .ZN(n4755) );
  XNOR2_X1 U5877 ( .A(n4755), .B(n4756), .ZN(n4748) );
  NAND2_X1 U5878 ( .A1(n4748), .A2(n5063), .ZN(n4749) );
  NAND2_X1 U5879 ( .A1(n4750), .A2(n4749), .ZN(n4751) );
  XNOR2_X1 U5880 ( .A(n4751), .B(n6256), .ZN(n6184) );
  NAND2_X1 U5881 ( .A1(n6185), .A2(n6184), .ZN(n6183) );
  NAND2_X1 U5882 ( .A1(n4751), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4752)
         );
  NAND2_X1 U5883 ( .A1(n6183), .A2(n4752), .ZN(n4762) );
  NAND2_X1 U5884 ( .A1(n4754), .A2(n4753), .ZN(n4760) );
  INV_X1 U5885 ( .A(n4755), .ZN(n4757) );
  NAND2_X1 U5886 ( .A1(n4757), .A2(n4756), .ZN(n4822) );
  XNOR2_X1 U5887 ( .A(n4822), .B(n4823), .ZN(n4758) );
  NAND2_X1 U5888 ( .A1(n4758), .A2(n5063), .ZN(n4759) );
  NAND2_X1 U5889 ( .A1(n4760), .A2(n4759), .ZN(n4814) );
  INV_X1 U5890 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6250) );
  XNOR2_X1 U5891 ( .A(n4814), .B(n6250), .ZN(n4761) );
  OAI21_X1 U5892 ( .B1(n4762), .B2(n4761), .A(n4816), .ZN(n6245) );
  INV_X1 U5893 ( .A(n4763), .ZN(n5149) );
  NAND2_X1 U5894 ( .A1(n6260), .A2(REIP_REG_7__SCAN_IN), .ZN(n6242) );
  NAND2_X1 U5895 ( .A1(n6199), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4764)
         );
  OAI211_X1 U5896 ( .C1(n6210), .C2(n5149), .A(n6242), .B(n4764), .ZN(n4765)
         );
  AOI21_X1 U5897 ( .B1(n5154), .B2(n6205), .A(n4765), .ZN(n4766) );
  OAI21_X1 U5898 ( .B1(n6245), .B2(n6181), .A(n4766), .ZN(U2979) );
  OR2_X1 U5899 ( .A1(n4769), .A2(n4768), .ZN(n4770) );
  AND2_X1 U5900 ( .A1(n4767), .A2(n4770), .ZN(n6060) );
  NOR2_X1 U5901 ( .A1(n4778), .A2(n4772), .ZN(n4773) );
  OR2_X1 U5902 ( .A1(n4848), .A2(n4773), .ZN(n6055) );
  OAI22_X1 U5903 ( .A1(n6055), .A2(n5546), .B1(n6056), .B2(n6123), .ZN(n4774)
         );
  AOI21_X1 U5904 ( .B1(n6060), .B2(n3906), .A(n4774), .ZN(n4775) );
  INV_X1 U5905 ( .A(n4775), .ZN(U2851) );
  INV_X1 U5906 ( .A(n6060), .ZN(n4777) );
  AOI22_X1 U5907 ( .A1(n5301), .A2(DATAI_8_), .B1(n6130), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4776) );
  OAI21_X1 U5908 ( .B1(n4777), .B2(n5867), .A(n4776), .ZN(U2883) );
  AOI21_X1 U5909 ( .B1(n4780), .B2(n4779), .A(n4778), .ZN(n6244) );
  INV_X1 U5910 ( .A(n6244), .ZN(n4783) );
  INV_X1 U5911 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4781) );
  OAI222_X1 U5912 ( .A1(n4783), .A2(n5546), .B1(n6118), .B2(n4782), .C1(n4781), 
        .C2(n6123), .ZN(U2852) );
  OAI21_X1 U5913 ( .B1(n4786), .B2(n4785), .A(n4551), .ZN(n4792) );
  INV_X1 U5914 ( .A(n4857), .ZN(n4788) );
  NAND3_X1 U5915 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n4946), .A3(n4787), .ZN(n4850) );
  NOR2_X1 U5916 ( .A1(n6406), .A2(n4850), .ZN(n4811) );
  AOI21_X1 U5917 ( .B1(n4789), .B2(n4788), .A(n4811), .ZN(n4793) );
  INV_X1 U5918 ( .A(n4793), .ZN(n4791) );
  AOI21_X1 U5919 ( .B1(n5000), .B2(n4850), .A(n4998), .ZN(n4790) );
  OAI21_X1 U5920 ( .B1(n4792), .B2(n4791), .A(n4790), .ZN(n4809) );
  OAI22_X1 U5921 ( .A1(n4793), .A2(n4792), .B1(n6433), .B2(n4850), .ZN(n4808)
         );
  AOI22_X1 U5922 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4809), .B1(n6346), 
        .B2(n4808), .ZN(n4795) );
  AOI22_X1 U5923 ( .A1(n6345), .A2(n4811), .B1(n4810), .B2(n5006), .ZN(n4794)
         );
  OAI211_X1 U5924 ( .C1(n5008), .C2(n4887), .A(n4795), .B(n4794), .ZN(U3097)
         );
  AOI22_X1 U5925 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4809), .B1(n6340), 
        .B2(n4808), .ZN(n4797) );
  AOI22_X1 U5926 ( .A1(n6339), .A2(n4811), .B1(n4810), .B2(n5018), .ZN(n4796)
         );
  OAI211_X1 U5927 ( .C1(n5020), .C2(n4887), .A(n4797), .B(n4796), .ZN(U3096)
         );
  AOI22_X1 U5928 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4809), .B1(n6358), 
        .B2(n4808), .ZN(n4799) );
  AOI22_X1 U5929 ( .A1(n6356), .A2(n4811), .B1(n4810), .B2(n5030), .ZN(n4798)
         );
  OAI211_X1 U5930 ( .C1(n5032), .C2(n4887), .A(n4799), .B(n4798), .ZN(U3099)
         );
  AOI22_X1 U5931 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4809), .B1(n6391), 
        .B2(n4808), .ZN(n4801) );
  AOI22_X1 U5932 ( .A1(n6389), .A2(n4811), .B1(n4810), .B2(n6387), .ZN(n4800)
         );
  OAI211_X1 U5933 ( .C1(n6396), .C2(n4887), .A(n4801), .B(n4800), .ZN(U3098)
         );
  AOI22_X1 U5934 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4809), .B1(n6312), 
        .B2(n4808), .ZN(n4803) );
  AOI22_X1 U5935 ( .A1(n6311), .A2(n4811), .B1(n4810), .B2(n5012), .ZN(n4802)
         );
  OAI211_X1 U5936 ( .C1(n5014), .C2(n4887), .A(n4803), .B(n4802), .ZN(U3092)
         );
  AOI22_X1 U5937 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4809), .B1(n6376), 
        .B2(n4808), .ZN(n4805) );
  AOI22_X1 U5938 ( .A1(n6375), .A2(n4811), .B1(n4810), .B2(n6374), .ZN(n4804)
         );
  OAI211_X1 U5939 ( .C1(n6379), .C2(n4887), .A(n4805), .B(n4804), .ZN(U3093)
         );
  AOI22_X1 U5940 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4809), .B1(n6330), 
        .B2(n4808), .ZN(n4807) );
  AOI22_X1 U5941 ( .A1(n6329), .A2(n4811), .B1(n4810), .B2(n5024), .ZN(n4806)
         );
  OAI211_X1 U5942 ( .C1(n5026), .C2(n4887), .A(n4807), .B(n4806), .ZN(U3094)
         );
  AOI22_X1 U5943 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4809), .B1(n6382), 
        .B2(n4808), .ZN(n4813) );
  AOI22_X1 U5944 ( .A1(n6381), .A2(n4811), .B1(n4810), .B2(n6380), .ZN(n4812)
         );
  OAI211_X1 U5945 ( .C1(n6385), .C2(n4887), .A(n4813), .B(n4812), .ZN(U3095)
         );
  NAND2_X1 U5946 ( .A1(n4814), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4815)
         );
  INV_X1 U5947 ( .A(n4817), .ZN(n4819) );
  NOR2_X1 U5948 ( .A1(n4819), .A2(n4818), .ZN(n4820) );
  INV_X1 U5949 ( .A(n4822), .ZN(n4824) );
  NAND3_X1 U5950 ( .A1(n4824), .A2(n5063), .A3(n4823), .ZN(n4825) );
  NAND2_X1 U5951 ( .A1(n5163), .A2(n4825), .ZN(n4929) );
  XNOR2_X1 U5952 ( .A(n4929), .B(n4836), .ZN(n4826) );
  OAI21_X1 U5953 ( .B1(n4827), .B2(n4826), .A(n3009), .ZN(n4842) );
  AND2_X1 U5954 ( .A1(n6277), .A2(REIP_REG_8__SCAN_IN), .ZN(n4839) );
  AOI21_X1 U5955 ( .B1(n6199), .B2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n4839), 
        .ZN(n4828) );
  OAI21_X1 U5956 ( .B1(n6210), .B2(n6058), .A(n4828), .ZN(n4829) );
  AOI21_X1 U5957 ( .B1(n6060), .B2(n6205), .A(n4829), .ZN(n4830) );
  OAI21_X1 U5958 ( .B1(n4842), .B2(n6181), .A(n4830), .ZN(U2978) );
  INV_X1 U5959 ( .A(n6055), .ZN(n4840) );
  NOR2_X1 U5960 ( .A1(n4836), .A2(n6250), .ZN(n6229) );
  AOI21_X1 U5961 ( .B1(n6287), .B2(n6281), .A(n6280), .ZN(n6261) );
  INV_X1 U5962 ( .A(n6261), .ZN(n4831) );
  NAND3_X1 U5963 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4832), .A3(n4831), 
        .ZN(n6257) );
  NOR2_X1 U5964 ( .A1(n6256), .A2(n6257), .ZN(n6247) );
  OAI21_X1 U5965 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n6247), .ZN(n4837) );
  NAND3_X1 U5966 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n4832), .ZN(n5103) );
  INV_X1 U5967 ( .A(n5384), .ZN(n4834) );
  NAND3_X1 U5968 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n4833), .ZN(n5104) );
  AOI22_X1 U5969 ( .A1(n6280), .A2(n5103), .B1(n4834), .B2(n5104), .ZN(n4835)
         );
  OAI22_X1 U5970 ( .A1(n6229), .A2(n4837), .B1(n6251), .B2(n4836), .ZN(n4838)
         );
  AOI211_X1 U5971 ( .C1(n6279), .C2(n4840), .A(n4839), .B(n4838), .ZN(n4841)
         );
  OAI21_X1 U5972 ( .B1(n5906), .B2(n4842), .A(n4841), .ZN(U3010) );
  INV_X1 U5973 ( .A(n4767), .ZN(n4844) );
  OAI21_X1 U5974 ( .B1(n4844), .B2(n3439), .A(n4937), .ZN(n6045) );
  AOI22_X1 U5975 ( .A1(n5301), .A2(DATAI_9_), .B1(n6130), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n4845) );
  OAI21_X1 U5976 ( .B1(n6045), .B2(n5867), .A(n4845), .ZN(U2882) );
  INV_X1 U5977 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4849) );
  CLKBUF_X1 U5978 ( .A(n4846), .Z(n5108) );
  OAI21_X1 U5979 ( .B1(n4848), .B2(n4847), .A(n5108), .ZN(n6048) );
  OAI222_X1 U5980 ( .A1(n6045), .A2(n6118), .B1(n4849), .B2(n6123), .C1(n5546), 
        .C2(n6048), .ZN(U2850) );
  AOI21_X1 U5981 ( .B1(n4887), .B2(n6366), .A(n6743), .ZN(n4855) );
  OAI21_X1 U5982 ( .B1(n5223), .B2(n4857), .A(n4551), .ZN(n4854) );
  NOR2_X1 U5983 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4850), .ZN(n4859)
         );
  OAI21_X1 U5984 ( .B1(n3149), .B2(n4859), .A(n5225), .ZN(n4851) );
  INV_X1 U5985 ( .A(n4851), .ZN(n4852) );
  OAI211_X1 U5986 ( .C1(n4855), .C2(n4854), .A(n4853), .B(n4852), .ZN(n4881)
         );
  NAND2_X1 U5987 ( .A1(n4881), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4862) );
  OAI22_X1 U5988 ( .A1(n4858), .A2(n4857), .B1(n4944), .B2(n4856), .ZN(n4884)
         );
  INV_X1 U5989 ( .A(n4859), .ZN(n4882) );
  OAI22_X1 U5990 ( .A1(n4969), .A2(n4882), .B1(n5014), .B2(n6366), .ZN(n4860)
         );
  AOI21_X1 U5991 ( .B1(n6312), .B2(n4884), .A(n4860), .ZN(n4861) );
  OAI211_X1 U5992 ( .C1(n4887), .C2(n6324), .A(n4862), .B(n4861), .ZN(U3084)
         );
  NAND2_X1 U5993 ( .A1(n4881), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4865) );
  OAI22_X1 U5994 ( .A1(n4959), .A2(n4882), .B1(n6379), .B2(n6366), .ZN(n4863)
         );
  AOI21_X1 U5995 ( .B1(n6376), .B2(n4884), .A(n4863), .ZN(n4864) );
  OAI211_X1 U5996 ( .C1(n4887), .C2(n6328), .A(n4865), .B(n4864), .ZN(U3085)
         );
  NAND2_X1 U5997 ( .A1(n4881), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4868) );
  OAI22_X1 U5998 ( .A1(n4964), .A2(n4882), .B1(n6396), .B2(n6366), .ZN(n4866)
         );
  AOI21_X1 U5999 ( .B1(n6391), .B2(n4884), .A(n4866), .ZN(n4867) );
  OAI211_X1 U6000 ( .C1(n4887), .C2(n6354), .A(n4868), .B(n4867), .ZN(U3090)
         );
  NAND2_X1 U6001 ( .A1(n4881), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4871) );
  OAI22_X1 U6002 ( .A1(n4987), .A2(n4882), .B1(n5020), .B2(n6366), .ZN(n4869)
         );
  AOI21_X1 U6003 ( .B1(n6340), .B2(n4884), .A(n4869), .ZN(n4870) );
  OAI211_X1 U6004 ( .C1(n4887), .C2(n6344), .A(n4871), .B(n4870), .ZN(U3088)
         );
  NAND2_X1 U6005 ( .A1(n4881), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4874) );
  OAI22_X1 U6006 ( .A1(n4981), .A2(n4882), .B1(n5032), .B2(n6366), .ZN(n4872)
         );
  AOI21_X1 U6007 ( .B1(n6358), .B2(n4884), .A(n4872), .ZN(n4873) );
  OAI211_X1 U6008 ( .C1(n4887), .C2(n6364), .A(n4874), .B(n4873), .ZN(U3091)
         );
  NAND2_X1 U6009 ( .A1(n4881), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4877) );
  OAI22_X1 U6010 ( .A1(n4977), .A2(n4882), .B1(n5026), .B2(n6366), .ZN(n4875)
         );
  AOI21_X1 U6011 ( .B1(n6330), .B2(n4884), .A(n4875), .ZN(n4876) );
  OAI211_X1 U6012 ( .C1(n4887), .C2(n6334), .A(n4877), .B(n4876), .ZN(U3086)
         );
  NAND2_X1 U6013 ( .A1(n4881), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4880) );
  OAI22_X1 U6014 ( .A1(n4973), .A2(n4882), .B1(n5008), .B2(n6366), .ZN(n4878)
         );
  AOI21_X1 U6015 ( .B1(n6346), .B2(n4884), .A(n4878), .ZN(n4879) );
  OAI211_X1 U6016 ( .C1(n4887), .C2(n6350), .A(n4880), .B(n4879), .ZN(U3089)
         );
  NAND2_X1 U6017 ( .A1(n4881), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4886) );
  OAI22_X1 U6018 ( .A1(n4954), .A2(n4882), .B1(n6385), .B2(n6366), .ZN(n4883)
         );
  AOI21_X1 U6019 ( .B1(n6382), .B2(n4884), .A(n4883), .ZN(n4885) );
  OAI211_X1 U6020 ( .C1(n4887), .C2(n6338), .A(n4886), .B(n4885), .ZN(U3087)
         );
  OAI21_X1 U6021 ( .B1(n4888), .B2(n5000), .A(n5217), .ZN(n4896) );
  NOR2_X1 U6022 ( .A1(n6406), .A2(n4895), .ZN(n4922) );
  INV_X1 U6023 ( .A(n4922), .ZN(n4889) );
  OAI21_X1 U6024 ( .B1(n4890), .B2(n6404), .A(n4889), .ZN(n4894) );
  INV_X1 U6025 ( .A(n4895), .ZN(n4891) );
  AOI22_X1 U6026 ( .A1(n4896), .A2(n4894), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4891), .ZN(n4928) );
  INV_X1 U6027 ( .A(n4989), .ZN(n4924) );
  INV_X1 U6028 ( .A(n4894), .ZN(n4897) );
  AOI22_X1 U6029 ( .A1(n4897), .A2(n4896), .B1(n4895), .B2(n5000), .ZN(n4898)
         );
  NAND2_X1 U6030 ( .A1(n4899), .A2(n4898), .ZN(n4921) );
  AOI22_X1 U6031 ( .A1(n6375), .A2(n4922), .B1(INSTQUEUE_REG_1__1__SCAN_IN), 
        .B2(n4921), .ZN(n4900) );
  OAI21_X1 U6032 ( .B1(n6328), .B2(n4924), .A(n4900), .ZN(n4901) );
  AOI21_X1 U6033 ( .B1(n6325), .B2(n4926), .A(n4901), .ZN(n4902) );
  OAI21_X1 U6034 ( .B1(n4928), .B2(n4963), .A(n4902), .ZN(U3029) );
  AOI22_X1 U6035 ( .A1(n6356), .A2(n4922), .B1(INSTQUEUE_REG_1__7__SCAN_IN), 
        .B2(n4921), .ZN(n4903) );
  OAI21_X1 U6036 ( .B1(n6364), .B2(n4924), .A(n4903), .ZN(n4904) );
  AOI21_X1 U6037 ( .B1(n6360), .B2(n4926), .A(n4904), .ZN(n4905) );
  OAI21_X1 U6038 ( .B1(n4928), .B2(n5035), .A(n4905), .ZN(U3035) );
  AOI22_X1 U6039 ( .A1(n6389), .A2(n4922), .B1(INSTQUEUE_REG_1__6__SCAN_IN), 
        .B2(n4921), .ZN(n4906) );
  OAI21_X1 U6040 ( .B1(n6354), .B2(n4924), .A(n4906), .ZN(n4907) );
  AOI21_X1 U6041 ( .B1(n6351), .B2(n4926), .A(n4907), .ZN(n4908) );
  OAI21_X1 U6042 ( .B1(n4928), .B2(n4968), .A(n4908), .ZN(U3034) );
  AOI22_X1 U6043 ( .A1(n6381), .A2(n4922), .B1(INSTQUEUE_REG_1__3__SCAN_IN), 
        .B2(n4921), .ZN(n4909) );
  OAI21_X1 U6044 ( .B1(n6338), .B2(n4924), .A(n4909), .ZN(n4910) );
  AOI21_X1 U6045 ( .B1(n6335), .B2(n4926), .A(n4910), .ZN(n4911) );
  OAI21_X1 U6046 ( .B1(n4928), .B2(n4958), .A(n4911), .ZN(U3031) );
  AOI22_X1 U6047 ( .A1(n6311), .A2(n4922), .B1(INSTQUEUE_REG_1__0__SCAN_IN), 
        .B2(n4921), .ZN(n4912) );
  OAI21_X1 U6048 ( .B1(n6324), .B2(n4924), .A(n4912), .ZN(n4913) );
  AOI21_X1 U6049 ( .B1(n6321), .B2(n4926), .A(n4913), .ZN(n4914) );
  OAI21_X1 U6050 ( .B1(n4928), .B2(n5017), .A(n4914), .ZN(U3028) );
  AOI22_X1 U6051 ( .A1(n6339), .A2(n4922), .B1(INSTQUEUE_REG_1__4__SCAN_IN), 
        .B2(n4921), .ZN(n4915) );
  OAI21_X1 U6052 ( .B1(n6344), .B2(n4924), .A(n4915), .ZN(n4916) );
  AOI21_X1 U6053 ( .B1(n6341), .B2(n4926), .A(n4916), .ZN(n4917) );
  OAI21_X1 U6054 ( .B1(n4928), .B2(n5023), .A(n4917), .ZN(U3032) );
  AOI22_X1 U6055 ( .A1(n6329), .A2(n4922), .B1(INSTQUEUE_REG_1__2__SCAN_IN), 
        .B2(n4921), .ZN(n4918) );
  OAI21_X1 U6056 ( .B1(n6334), .B2(n4924), .A(n4918), .ZN(n4919) );
  AOI21_X1 U6057 ( .B1(n6331), .B2(n4926), .A(n4919), .ZN(n4920) );
  OAI21_X1 U6058 ( .B1(n4928), .B2(n5029), .A(n4920), .ZN(U3030) );
  AOI22_X1 U6059 ( .A1(n6345), .A2(n4922), .B1(INSTQUEUE_REG_1__5__SCAN_IN), 
        .B2(n4921), .ZN(n4923) );
  OAI21_X1 U6060 ( .B1(n6350), .B2(n4924), .A(n4923), .ZN(n4925) );
  AOI21_X1 U6061 ( .B1(n6347), .B2(n4926), .A(n4925), .ZN(n4927) );
  OAI21_X1 U6062 ( .B1(n4928), .B2(n5011), .A(n4927), .ZN(U3033) );
  NAND2_X1 U6063 ( .A1(n4929), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n4930)
         );
  NAND2_X1 U6064 ( .A1(n4931), .A2(n4930), .ZN(n5042) );
  INV_X1 U6065 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U6066 ( .A1(n5163), .A2(n6225), .ZN(n5041) );
  NAND2_X1 U6067 ( .A1(n5043), .A2(n5041), .ZN(n4932) );
  XNOR2_X1 U6068 ( .A(n3011), .B(n4932), .ZN(n6238) );
  NAND2_X1 U6069 ( .A1(n6238), .A2(n6204), .ZN(n4935) );
  NAND2_X1 U6070 ( .A1(n6260), .A2(REIP_REG_9__SCAN_IN), .ZN(n6234) );
  OAI21_X1 U6071 ( .B1(n5651), .B2(n6043), .A(n6234), .ZN(n4933) );
  AOI21_X1 U6072 ( .B1(n6177), .B2(n6046), .A(n4933), .ZN(n4934) );
  OAI211_X1 U6073 ( .C1(n5679), .C2(n6045), .A(n4935), .B(n4934), .ZN(U2977)
         );
  AOI21_X1 U6074 ( .B1(n4938), .B2(n4937), .A(n4936), .ZN(n4939) );
  INV_X1 U6075 ( .A(n4939), .ZN(n6039) );
  AOI22_X1 U6076 ( .A1(n5301), .A2(DATAI_10_), .B1(n6130), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4940) );
  OAI21_X1 U6077 ( .B1(n6039), .B2(n5867), .A(n4940), .ZN(U2881) );
  XNOR2_X1 U6078 ( .A(n5108), .B(n4941), .ZN(n6227) );
  AOI22_X1 U6079 ( .A1(n6227), .A2(n6563), .B1(EBX_REG_10__SCAN_IN), .B2(n6562), .ZN(n4942) );
  OAI21_X1 U6080 ( .B1(n6039), .B2(n6118), .A(n4942), .ZN(U2849) );
  AND2_X1 U6081 ( .A1(n4943), .A2(n5223), .ZN(n4996) );
  NOR2_X1 U6082 ( .A1(n4944), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4945)
         );
  AOI22_X1 U6083 ( .A1(n4996), .A2(n4551), .B1(n6305), .B2(n4945), .ZN(n4992)
         );
  NAND3_X1 U6084 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n6718), .A3(n4946), .ZN(n4999) );
  NOR2_X1 U6085 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4999), .ZN(n4953)
         );
  OR3_X1 U6086 ( .A1(n3348), .A2(n3015), .A3(n4947), .ZN(n6304) );
  INV_X1 U6087 ( .A(n6304), .ZN(n4948) );
  OAI21_X1 U6088 ( .B1(n4989), .B2(n4948), .A(n5217), .ZN(n4950) );
  INV_X1 U6089 ( .A(n4996), .ZN(n4949) );
  NAND2_X1 U6090 ( .A1(n4950), .A2(n4949), .ZN(n4952) );
  OAI221_X1 U6091 ( .B1(n4953), .B2(n3149), .C1(n4953), .C2(n4952), .A(n4951), 
        .ZN(n4985) );
  NAND2_X1 U6092 ( .A1(n4985), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4957) );
  INV_X1 U6093 ( .A(n4953), .ZN(n4986) );
  OAI22_X1 U6094 ( .A1(n4954), .A2(n4986), .B1(n6338), .B2(n6304), .ZN(n4955)
         );
  AOI21_X1 U6095 ( .B1(n6335), .B2(n4989), .A(n4955), .ZN(n4956) );
  OAI211_X1 U6096 ( .C1(n4992), .C2(n4958), .A(n4957), .B(n4956), .ZN(U3039)
         );
  NAND2_X1 U6097 ( .A1(n4985), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4962) );
  OAI22_X1 U6098 ( .A1(n4959), .A2(n4986), .B1(n6328), .B2(n6304), .ZN(n4960)
         );
  AOI21_X1 U6099 ( .B1(n6325), .B2(n4989), .A(n4960), .ZN(n4961) );
  OAI211_X1 U6100 ( .C1(n4992), .C2(n4963), .A(n4962), .B(n4961), .ZN(U3037)
         );
  NAND2_X1 U6101 ( .A1(n4985), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4967) );
  OAI22_X1 U6102 ( .A1(n4964), .A2(n4986), .B1(n6354), .B2(n6304), .ZN(n4965)
         );
  AOI21_X1 U6103 ( .B1(n6351), .B2(n4989), .A(n4965), .ZN(n4966) );
  OAI211_X1 U6104 ( .C1(n4992), .C2(n4968), .A(n4967), .B(n4966), .ZN(U3042)
         );
  NAND2_X1 U6105 ( .A1(n4985), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4972) );
  OAI22_X1 U6106 ( .A1(n4969), .A2(n4986), .B1(n6324), .B2(n6304), .ZN(n4970)
         );
  AOI21_X1 U6107 ( .B1(n6321), .B2(n4989), .A(n4970), .ZN(n4971) );
  OAI211_X1 U6108 ( .C1(n4992), .C2(n5017), .A(n4972), .B(n4971), .ZN(U3036)
         );
  NAND2_X1 U6109 ( .A1(n4985), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4976) );
  OAI22_X1 U6110 ( .A1(n4973), .A2(n4986), .B1(n6350), .B2(n6304), .ZN(n4974)
         );
  AOI21_X1 U6111 ( .B1(n6347), .B2(n4989), .A(n4974), .ZN(n4975) );
  OAI211_X1 U6112 ( .C1(n4992), .C2(n5011), .A(n4976), .B(n4975), .ZN(U3041)
         );
  NAND2_X1 U6113 ( .A1(n4985), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4980) );
  OAI22_X1 U6114 ( .A1(n4977), .A2(n4986), .B1(n6334), .B2(n6304), .ZN(n4978)
         );
  AOI21_X1 U6115 ( .B1(n6331), .B2(n4989), .A(n4978), .ZN(n4979) );
  OAI211_X1 U6116 ( .C1(n4992), .C2(n5029), .A(n4980), .B(n4979), .ZN(U3038)
         );
  NAND2_X1 U6117 ( .A1(n4985), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4984) );
  OAI22_X1 U6118 ( .A1(n4981), .A2(n4986), .B1(n6364), .B2(n6304), .ZN(n4982)
         );
  AOI21_X1 U6119 ( .B1(n6360), .B2(n4989), .A(n4982), .ZN(n4983) );
  OAI211_X1 U6120 ( .C1(n4992), .C2(n5035), .A(n4984), .B(n4983), .ZN(U3043)
         );
  NAND2_X1 U6121 ( .A1(n4985), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4991) );
  OAI22_X1 U6122 ( .A1(n4987), .A2(n4986), .B1(n6344), .B2(n6304), .ZN(n4988)
         );
  AOI21_X1 U6123 ( .B1(n6341), .B2(n4989), .A(n4988), .ZN(n4990) );
  OAI211_X1 U6124 ( .C1(n4992), .C2(n5023), .A(n4991), .B(n4990), .ZN(U3040)
         );
  OR2_X1 U6125 ( .A1(n3015), .A2(n5777), .ZN(n4994) );
  AOI21_X1 U6126 ( .B1(n4551), .B2(n4994), .A(n4993), .ZN(n5003) );
  NOR2_X1 U6127 ( .A1(n4995), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6299)
         );
  AOI21_X1 U6128 ( .B1(n4996), .B2(n3255), .A(n6299), .ZN(n4997) );
  OAI22_X1 U6129 ( .A1(n5003), .A2(n4997), .B1(n4999), .B2(n6433), .ZN(n6300)
         );
  INV_X1 U6130 ( .A(n6300), .ZN(n5036) );
  INV_X1 U6131 ( .A(n4997), .ZN(n5002) );
  AOI21_X1 U6132 ( .B1(n5000), .B2(n4999), .A(n4998), .ZN(n5001) );
  OAI21_X1 U6133 ( .B1(n5003), .B2(n5002), .A(n5001), .ZN(n6301) );
  NOR3_X1 U6134 ( .A1(n3348), .A2(n3015), .A3(n5004), .ZN(n5005) );
  AOI22_X1 U6135 ( .A1(n6345), .A2(n6299), .B1(n5006), .B2(n6298), .ZN(n5007)
         );
  OAI21_X1 U6136 ( .B1(n5008), .B2(n6304), .A(n5007), .ZN(n5009) );
  AOI21_X1 U6137 ( .B1(n6301), .B2(INSTQUEUE_REG_3__5__SCAN_IN), .A(n5009), 
        .ZN(n5010) );
  OAI21_X1 U6138 ( .B1(n5036), .B2(n5011), .A(n5010), .ZN(U3049) );
  AOI22_X1 U6139 ( .A1(n6311), .A2(n6299), .B1(n5012), .B2(n6298), .ZN(n5013)
         );
  OAI21_X1 U6140 ( .B1(n5014), .B2(n6304), .A(n5013), .ZN(n5015) );
  AOI21_X1 U6141 ( .B1(n6301), .B2(INSTQUEUE_REG_3__0__SCAN_IN), .A(n5015), 
        .ZN(n5016) );
  OAI21_X1 U6142 ( .B1(n5036), .B2(n5017), .A(n5016), .ZN(U3044) );
  AOI22_X1 U6143 ( .A1(n6339), .A2(n6299), .B1(n5018), .B2(n6298), .ZN(n5019)
         );
  OAI21_X1 U6144 ( .B1(n5020), .B2(n6304), .A(n5019), .ZN(n5021) );
  AOI21_X1 U6145 ( .B1(n6301), .B2(INSTQUEUE_REG_3__4__SCAN_IN), .A(n5021), 
        .ZN(n5022) );
  OAI21_X1 U6146 ( .B1(n5036), .B2(n5023), .A(n5022), .ZN(U3048) );
  AOI22_X1 U6147 ( .A1(n6329), .A2(n6299), .B1(n5024), .B2(n6298), .ZN(n5025)
         );
  OAI21_X1 U6148 ( .B1(n5026), .B2(n6304), .A(n5025), .ZN(n5027) );
  AOI21_X1 U6149 ( .B1(n6301), .B2(INSTQUEUE_REG_3__2__SCAN_IN), .A(n5027), 
        .ZN(n5028) );
  OAI21_X1 U6150 ( .B1(n5036), .B2(n5029), .A(n5028), .ZN(U3046) );
  AOI22_X1 U6151 ( .A1(n6356), .A2(n6299), .B1(n5030), .B2(n6298), .ZN(n5031)
         );
  OAI21_X1 U6152 ( .B1(n5032), .B2(n6304), .A(n5031), .ZN(n5033) );
  AOI21_X1 U6153 ( .B1(n6301), .B2(INSTQUEUE_REG_3__7__SCAN_IN), .A(n5033), 
        .ZN(n5034) );
  OAI21_X1 U6154 ( .B1(n5036), .B2(n5035), .A(n5034), .ZN(U3051) );
  NOR2_X1 U6155 ( .A1(n4936), .A2(n5038), .ZN(n5039) );
  OR2_X1 U6156 ( .A1(n5139), .A2(n5039), .ZN(n6119) );
  AOI22_X1 U6157 ( .A1(n5301), .A2(DATAI_11_), .B1(n6130), .B2(
        EAX_REG_11__SCAN_IN), .ZN(n5040) );
  OAI21_X1 U6158 ( .B1(n6119), .B2(n5867), .A(n5040), .ZN(U2880) );
  NAND2_X1 U6159 ( .A1(n5042), .A2(n5041), .ZN(n5044) );
  XNOR2_X1 U6160 ( .A(n5891), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5045)
         );
  XNOR2_X1 U6161 ( .A(n5098), .B(n5045), .ZN(n6230) );
  NAND2_X1 U6162 ( .A1(n6230), .A2(n6204), .ZN(n5049) );
  INV_X1 U6163 ( .A(REIP_REG_10__SCAN_IN), .ZN(n5046) );
  NOR2_X1 U6164 ( .A1(n6216), .A2(n5046), .ZN(n6226) );
  NOR2_X1 U6165 ( .A1(n6210), .A2(n6037), .ZN(n5047) );
  AOI211_X1 U6166 ( .C1(n6199), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n6226), 
        .B(n5047), .ZN(n5048) );
  OAI211_X1 U6167 ( .C1(n5679), .C2(n6039), .A(n5049), .B(n5048), .ZN(U2976)
         );
  INV_X1 U6168 ( .A(n6555), .ZN(n6439) );
  NOR3_X1 U6169 ( .A1(n5050), .A2(n3149), .A3(n6439), .ZN(n6435) );
  AND2_X1 U6170 ( .A1(n5052), .A2(n5051), .ZN(n6447) );
  OR2_X1 U6171 ( .A1(n6277), .A2(n6447), .ZN(n5053) );
  OR2_X1 U6172 ( .A1(n6435), .A2(n5053), .ZN(n5054) );
  NAND2_X1 U6173 ( .A1(n5473), .A2(n5055), .ZN(n5059) );
  INV_X1 U6174 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5476) );
  XNOR2_X1 U6175 ( .A(n5057), .B(n5476), .ZN(n5429) );
  NOR2_X1 U6176 ( .A1(n5429), .A2(n6532), .ZN(n5058) );
  NOR2_X1 U6177 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .ZN(n5072) );
  INV_X1 U6178 ( .A(n5072), .ZN(n6427) );
  NAND3_X1 U6179 ( .A1(n5060), .A2(EBX_REG_31__SCAN_IN), .A3(n6427), .ZN(n5061) );
  NOR2_X2 U6180 ( .A1(n5067), .A2(n5061), .ZN(n6086) );
  OR2_X1 U6181 ( .A1(n6461), .A2(n6427), .ZN(n5062) );
  AND2_X1 U6182 ( .A1(n5063), .A2(n5062), .ZN(n5472) );
  NOR2_X1 U6183 ( .A1(n5072), .A2(EBX_REG_31__SCAN_IN), .ZN(n5064) );
  AND2_X1 U6184 ( .A1(n5071), .A2(n5064), .ZN(n5065) );
  NOR2_X1 U6185 ( .A1(n5472), .A2(n5065), .ZN(n5066) );
  AOI22_X1 U6186 ( .A1(n5068), .A2(n6086), .B1(n3003), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n5078) );
  NAND2_X1 U6187 ( .A1(n5473), .A2(n5069), .ZN(n6088) );
  INV_X1 U6188 ( .A(n6088), .ZN(n6102) );
  NAND2_X1 U6189 ( .A1(n6102), .A2(n3255), .ZN(n5077) );
  AND2_X1 U6190 ( .A1(n5429), .A2(STATE2_REG_1__SCAN_IN), .ZN(n5070) );
  OAI21_X1 U6191 ( .B1(n6097), .B2(n6108), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5076) );
  AND3_X1 U6192 ( .A1(n5073), .A2(n5072), .A3(n5071), .ZN(n5074) );
  NAND2_X2 U6193 ( .A1(n5473), .A2(n5074), .ZN(n6084) );
  NAND2_X1 U6194 ( .A1(n6084), .A2(n5329), .ZN(n6076) );
  NAND2_X1 U6195 ( .A1(n6076), .A2(REIP_REG_0__SCAN_IN), .ZN(n5075) );
  AND4_X1 U6196 ( .A1(n5078), .A2(n5077), .A3(n5076), .A4(n5075), .ZN(n5079)
         );
  OAI21_X1 U6197 ( .B1(n5080), .B2(n6105), .A(n5079), .ZN(U2827) );
  NAND2_X1 U6198 ( .A1(n5139), .A2(n5081), .ZN(n5175) );
  OR2_X1 U6199 ( .A1(n5139), .A2(n5081), .ZN(n5082) );
  NAND2_X1 U6200 ( .A1(n5175), .A2(n5082), .ZN(n5171) );
  INV_X1 U6201 ( .A(n5179), .ZN(n5085) );
  NAND2_X1 U6202 ( .A1(n5109), .A2(n5083), .ZN(n5084) );
  NAND2_X1 U6203 ( .A1(n5085), .A2(n5084), .ZN(n6218) );
  OAI22_X1 U6204 ( .A1(n6218), .A2(n5546), .B1(n6719), .B2(n6123), .ZN(n5086)
         );
  INV_X1 U6205 ( .A(n5086), .ZN(n5087) );
  OAI21_X1 U6206 ( .B1(n5171), .B2(n6118), .A(n5087), .ZN(U2847) );
  INV_X1 U6207 ( .A(DATAI_12_), .ZN(n5089) );
  OAI222_X1 U6208 ( .A1(n5171), .A2(n5867), .B1(n5432), .B2(n5090), .C1(n5089), 
        .C2(n5088), .ZN(U2879) );
  NAND2_X1 U6209 ( .A1(n5329), .A2(n5091), .ZN(n6070) );
  INV_X1 U6210 ( .A(n6070), .ZN(n6081) );
  INV_X1 U6211 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6491) );
  NAND3_X1 U6212 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .ZN(n5093) );
  INV_X1 U6213 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6484) );
  INV_X1 U6214 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6477) );
  NAND3_X1 U6215 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_3__SCAN_IN), .A3(
        REIP_REG_2__SCAN_IN), .ZN(n6083) );
  OR2_X1 U6216 ( .A1(n6477), .A2(n6083), .ZN(n5113) );
  NOR2_X1 U6217 ( .A1(n6479), .A2(n5113), .ZN(n5145) );
  NAND2_X1 U6218 ( .A1(REIP_REG_6__SCAN_IN), .A2(n5145), .ZN(n5146) );
  NOR2_X1 U6219 ( .A1(n6484), .A2(n5146), .ZN(n6053) );
  NAND2_X1 U6220 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6053), .ZN(n6026) );
  INV_X1 U6221 ( .A(n6026), .ZN(n6034) );
  NAND2_X1 U6222 ( .A1(n6034), .A2(n5329), .ZN(n6033) );
  OAI21_X1 U6223 ( .B1(n5093), .B2(n6033), .A(n6076), .ZN(n6031) );
  OAI22_X1 U6224 ( .A1(n5166), .A2(n6078), .B1(n6491), .B2(n6031), .ZN(n5092)
         );
  AOI211_X1 U6225 ( .C1(n3003), .C2(EBX_REG_12__SCAN_IN), .A(n6081), .B(n5092), 
        .ZN(n5095) );
  NOR2_X1 U6226 ( .A1(n6026), .A2(n5093), .ZN(n5127) );
  INV_X1 U6227 ( .A(n5127), .ZN(n5094) );
  NOR2_X1 U6228 ( .A1(n6084), .A2(n5094), .ZN(n6005) );
  NAND2_X1 U6229 ( .A1(n6005), .A2(n6491), .ZN(n5184) );
  OAI211_X1 U6230 ( .C1(n6218), .C2(n6100), .A(n5095), .B(n5184), .ZN(n5096)
         );
  AOI21_X1 U6231 ( .B1(n6108), .B2(n5168), .A(n5096), .ZN(n5097) );
  OAI21_X1 U6232 ( .B1(n6038), .B2(n5171), .A(n5097), .ZN(U2815) );
  NAND2_X1 U6233 ( .A1(n3010), .A2(n5099), .ZN(n5160) );
  AOI22_X1 U6234 ( .A1(n5160), .A2(n5891), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n5098), .ZN(n5101) );
  XNOR2_X1 U6235 ( .A(n5891), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5100)
         );
  XNOR2_X1 U6236 ( .A(n5101), .B(n5100), .ZN(n6182) );
  NAND3_X1 U6237 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n6229), .ZN(n5105) );
  INV_X1 U6238 ( .A(n5105), .ZN(n5102) );
  OAI21_X1 U6239 ( .B1(n5102), .B2(n6228), .A(n6251), .ZN(n6214) );
  NOR2_X1 U6240 ( .A1(n5103), .A2(n5105), .ZN(n5386) );
  NAND2_X1 U6241 ( .A1(n6280), .A2(n5386), .ZN(n5943) );
  NOR2_X1 U6242 ( .A1(n5105), .A2(n5104), .ZN(n5960) );
  NAND2_X1 U6243 ( .A1(n6287), .A2(n5960), .ZN(n6213) );
  NAND2_X1 U6244 ( .A1(n5943), .A2(n6213), .ZN(n6211) );
  INV_X1 U6245 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5382) );
  AOI22_X1 U6246 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6214), .B1(n6211), .B2(n5382), .ZN(n5112) );
  OAI21_X1 U6247 ( .B1(n5108), .B2(n5107), .A(n5106), .ZN(n5110) );
  AND2_X1 U6248 ( .A1(n5110), .A2(n5109), .ZN(n6116) );
  AOI22_X1 U6249 ( .A1(n6116), .A2(n6279), .B1(n6260), .B2(
        REIP_REG_11__SCAN_IN), .ZN(n5111) );
  OAI211_X1 U6250 ( .C1(n6182), .C2(n5906), .A(n5112), .B(n5111), .ZN(U3007)
         );
  OAI21_X1 U6251 ( .B1(n6084), .B2(n5145), .A(n5329), .ZN(n6069) );
  OAI21_X1 U6252 ( .B1(n6084), .B2(n5113), .A(n6479), .ZN(n5120) );
  AOI21_X1 U6253 ( .B1(n6108), .B2(n5114), .A(n6081), .ZN(n5115) );
  OAI21_X1 U6254 ( .B1(n6065), .B2(n4224), .A(n5115), .ZN(n5119) );
  OAI22_X1 U6255 ( .A1(n5117), .A2(n6078), .B1(n6100), .B2(n5116), .ZN(n5118)
         );
  AOI211_X1 U6256 ( .C1(n6069), .C2(n5120), .A(n5119), .B(n5118), .ZN(n5121)
         );
  OAI21_X1 U6257 ( .B1(n6105), .B2(n5122), .A(n5121), .ZN(U2822) );
  NAND2_X1 U6258 ( .A1(n5139), .A2(n5123), .ZN(n5902) );
  AND2_X1 U6259 ( .A1(n5902), .A2(n5124), .ZN(n5126) );
  AND2_X1 U6260 ( .A1(n5139), .A2(n5125), .ZN(n5190) );
  INV_X1 U6261 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5650) );
  INV_X1 U6262 ( .A(n6076), .ZN(n5342) );
  INV_X1 U6263 ( .A(n5329), .ZN(n6077) );
  INV_X1 U6264 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6497) );
  NAND3_X1 U6265 ( .A1(REIP_REG_14__SCAN_IN), .A2(REIP_REG_13__SCAN_IN), .A3(
        REIP_REG_12__SCAN_IN), .ZN(n6006) );
  INV_X1 U6266 ( .A(n6006), .ZN(n5290) );
  NAND3_X1 U6267 ( .A1(REIP_REG_15__SCAN_IN), .A2(n5127), .A3(n5290), .ZN(
        n6004) );
  NOR2_X1 U6268 ( .A1(n6497), .A2(n6004), .ZN(n5994) );
  NAND2_X1 U6269 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5994), .ZN(n5132) );
  NOR2_X1 U6270 ( .A1(n6077), .A2(n5132), .ZN(n5210) );
  NOR2_X1 U6271 ( .A1(n5342), .A2(n5210), .ZN(n5997) );
  AOI22_X1 U6272 ( .A1(EBX_REG_18__SCAN_IN), .A2(n3003), .B1(
        REIP_REG_18__SCAN_IN), .B2(n5997), .ZN(n5128) );
  OAI211_X1 U6273 ( .C1(n6078), .C2(n5650), .A(n5128), .B(n6070), .ZN(n5135)
         );
  INV_X1 U6274 ( .A(n5205), .ZN(n5130) );
  MUX2_X1 U6275 ( .A(n5130), .B(n5129), .S(n5204), .Z(n5196) );
  OR2_X1 U6276 ( .A1(n5916), .A2(n5196), .ZN(n5194) );
  NAND2_X1 U6277 ( .A1(n5916), .A2(n5196), .ZN(n5131) );
  AND2_X1 U6278 ( .A1(n5194), .A2(n5131), .ZN(n5907) );
  INV_X1 U6279 ( .A(n5907), .ZN(n5172) );
  NOR2_X1 U6280 ( .A1(n6084), .A2(n5132), .ZN(n5854) );
  INV_X1 U6281 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6500) );
  AOI22_X1 U6282 ( .A1(n5854), .A2(n6500), .B1(n6108), .B2(n5653), .ZN(n5133)
         );
  OAI21_X1 U6283 ( .B1(n5172), .B2(n6100), .A(n5133), .ZN(n5134) );
  NOR2_X1 U6284 ( .A1(n5135), .A2(n5134), .ZN(n5136) );
  OAI21_X1 U6285 ( .B1(n5656), .B2(n6038), .A(n5136), .ZN(U2809) );
  INV_X1 U6286 ( .A(n5175), .ZN(n5177) );
  NAND2_X1 U6287 ( .A1(n5139), .A2(n5138), .ZN(n5900) );
  OAI21_X1 U6288 ( .B1(n5281), .B2(n5140), .A(n5900), .ZN(n5663) );
  INV_X1 U6289 ( .A(EBX_REG_16__SCAN_IN), .ZN(n5144) );
  OR2_X1 U6290 ( .A1(n5932), .A2(n5142), .ZN(n5143) );
  NAND2_X1 U6291 ( .A1(n5141), .A2(n5143), .ZN(n6016) );
  OAI222_X1 U6292 ( .A1(n5663), .A2(n6118), .B1(n6123), .B2(n5144), .C1(n6016), 
        .C2(n5546), .ZN(U2843) );
  INV_X1 U6293 ( .A(n6084), .ZN(n6054) );
  INV_X1 U6294 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6481) );
  AND3_X1 U6295 ( .A1(n6054), .A2(n6481), .A3(n5145), .ZN(n6068) );
  OAI21_X1 U6296 ( .B1(n6068), .B2(n6069), .A(REIP_REG_7__SCAN_IN), .ZN(n5148)
         );
  OR3_X1 U6297 ( .A1(n6084), .A2(REIP_REG_7__SCAN_IN), .A3(n5146), .ZN(n5147)
         );
  OAI211_X1 U6298 ( .C1(n5149), .C2(n6094), .A(n5148), .B(n5147), .ZN(n5153)
         );
  AOI22_X1 U6299 ( .A1(EBX_REG_7__SCAN_IN), .A2(n3003), .B1(n6086), .B2(n6244), 
        .ZN(n5150) );
  OAI211_X1 U6300 ( .C1(n6078), .C2(n5151), .A(n5150), .B(n6070), .ZN(n5152)
         );
  AOI211_X1 U6301 ( .C1(n6073), .C2(n5154), .A(n5153), .B(n5152), .ZN(n5155)
         );
  INV_X1 U6302 ( .A(n5155), .ZN(U2820) );
  NOR2_X2 U6303 ( .A1(n6130), .A2(n5156), .ZN(n6127) );
  AOI22_X1 U6304 ( .A1(n6127), .A2(DATAI_18_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n6130), .ZN(n5159) );
  NAND2_X1 U6305 ( .A1(n6131), .A2(DATAI_2_), .ZN(n5158) );
  OAI211_X1 U6306 ( .C1(n5656), .C2(n5867), .A(n5159), .B(n5158), .ZN(U2873)
         );
  OAI21_X1 U6307 ( .B1(n5160), .B2(INSTADDRPOINTER_REG_11__SCAN_IN), .A(n5891), 
        .ZN(n5162) );
  NAND2_X1 U6308 ( .A1(n5162), .A2(n5161), .ZN(n5274) );
  INV_X1 U6309 ( .A(n5273), .ZN(n5164) );
  NAND2_X1 U6310 ( .A1(n5163), .A2(n6223), .ZN(n5272) );
  NAND2_X1 U6311 ( .A1(n5164), .A2(n5272), .ZN(n5165) );
  XNOR2_X1 U6312 ( .A(n5274), .B(n5165), .ZN(n6220) );
  NAND2_X1 U6313 ( .A1(n6220), .A2(n6204), .ZN(n5170) );
  OAI22_X1 U6314 ( .A1(n5651), .A2(n5166), .B1(n6216), .B2(n6491), .ZN(n5167)
         );
  AOI21_X1 U6315 ( .B1(n6177), .B2(n5168), .A(n5167), .ZN(n5169) );
  OAI211_X1 U6316 ( .C1(n5679), .C2(n5171), .A(n5170), .B(n5169), .ZN(U2974)
         );
  OAI222_X1 U6317 ( .A1(n6118), .A2(n5656), .B1(n5173), .B2(n6123), .C1(n5172), 
        .C2(n5546), .ZN(U2841) );
  INV_X1 U6318 ( .A(n5174), .ZN(n5176) );
  OAI21_X1 U6319 ( .B1(n5177), .B2(n5176), .A(n5288), .ZN(n5280) );
  OR2_X1 U6320 ( .A1(n5179), .A2(n5178), .ZN(n5180) );
  AND2_X1 U6321 ( .A1(n5293), .A2(n5180), .ZN(n5954) );
  NOR2_X1 U6322 ( .A1(n6123), .A2(n6695), .ZN(n5181) );
  AOI21_X1 U6323 ( .B1(n5954), .B2(n6563), .A(n5181), .ZN(n5182) );
  OAI21_X1 U6324 ( .B1(n5280), .B2(n6118), .A(n5182), .ZN(U2846) );
  AOI22_X1 U6325 ( .A1(PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n6097), .B1(n6086), 
        .B2(n5954), .ZN(n5183) );
  OAI211_X1 U6326 ( .C1(n6065), .C2(n6695), .A(n5183), .B(n6070), .ZN(n5186)
         );
  INV_X1 U6327 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6493) );
  NAND2_X1 U6328 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6005), .ZN(n5291) );
  OAI222_X1 U6329 ( .A1(n6493), .A2(n6031), .B1(n6493), .B2(n5184), .C1(
        REIP_REG_13__SCAN_IN), .C2(n5291), .ZN(n5185) );
  AOI211_X1 U6330 ( .C1(n5277), .C2(n6108), .A(n5186), .B(n5185), .ZN(n5187)
         );
  OAI21_X1 U6331 ( .B1(n5280), .B2(n6038), .A(n5187), .ZN(U2814) );
  AOI22_X1 U6332 ( .A1(n5301), .A2(DATAI_13_), .B1(n6130), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n5188) );
  OAI21_X1 U6333 ( .B1(n5280), .B2(n5867), .A(n5188), .ZN(U2878) );
  INV_X1 U6334 ( .A(n5189), .ZN(n5192) );
  INV_X1 U6335 ( .A(n5190), .ZN(n5191) );
  AOI21_X1 U6336 ( .B1(n5192), .B2(n5191), .A(n3008), .ZN(n5887) );
  NAND2_X1 U6337 ( .A1(n5194), .A2(n5193), .ZN(n5195) );
  OAI21_X1 U6338 ( .B1(n5203), .B2(n5196), .A(n5195), .ZN(n5857) );
  OAI22_X1 U6339 ( .A1(n5857), .A2(n5546), .B1(n5197), .B2(n6123), .ZN(n5198)
         );
  AOI21_X1 U6340 ( .B1(n5887), .B2(n3906), .A(n5198), .ZN(n5199) );
  INV_X1 U6341 ( .A(n5199), .ZN(U2840) );
  INV_X1 U6342 ( .A(n5265), .ZN(n5200) );
  OAI21_X1 U6343 ( .B1(n5202), .B2(n3008), .A(n5200), .ZN(n5883) );
  MUX2_X1 U6344 ( .A(n5205), .B(n5204), .S(n5203), .Z(n5206) );
  XOR2_X1 U6345 ( .A(n5207), .B(n5206), .Z(n5765) );
  INV_X1 U6346 ( .A(n5765), .ZN(n5213) );
  INV_X1 U6347 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5271) );
  NOR2_X1 U6348 ( .A1(n5633), .A2(n6078), .ZN(n5208) );
  AOI21_X1 U6349 ( .B1(n6108), .B2(n5636), .A(n5208), .ZN(n5209) );
  OAI21_X1 U6350 ( .B1(n6065), .B2(n5271), .A(n5209), .ZN(n5212) );
  INV_X1 U6351 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6503) );
  NAND3_X1 U6352 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        n5854), .ZN(n5339) );
  NAND4_X1 U6353 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        n5210), .A4(REIP_REG_18__SCAN_IN), .ZN(n5341) );
  NAND2_X1 U6354 ( .A1(n6076), .A2(n5341), .ZN(n5844) );
  AOI21_X1 U6355 ( .B1(n6503), .B2(n5339), .A(n5844), .ZN(n5211) );
  AOI211_X1 U6356 ( .C1(n6086), .C2(n5213), .A(n5212), .B(n5211), .ZN(n5214)
         );
  OAI21_X1 U6357 ( .B1(n5883), .B2(n6038), .A(n5214), .ZN(U2807) );
  INV_X1 U6358 ( .A(n6298), .ZN(n5215) );
  NAND3_X1 U6359 ( .A1(n5215), .A2(n4551), .A3(n5257), .ZN(n5218) );
  AOI21_X1 U6360 ( .B1(n5218), .B2(n5217), .A(n5216), .ZN(n5222) );
  NOR2_X1 U6361 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5219), .ZN(n5255)
         );
  NOR2_X1 U6362 ( .A1(n3149), .A2(n5255), .ZN(n5220) );
  NOR4_X2 U6363 ( .A1(n5222), .A2(n6316), .A3(n5221), .A4(n5220), .ZN(n5262)
         );
  INV_X1 U6364 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5230) );
  NAND2_X1 U6365 ( .A1(n5223), .A2(n4551), .ZN(n6309) );
  OAI22_X1 U6366 ( .A1(n6309), .A2(n5226), .B1(n5225), .B2(n5224), .ZN(n5259)
         );
  AOI22_X1 U6367 ( .A1(n6389), .A2(n5255), .B1(n6351), .B2(n6298), .ZN(n5227)
         );
  OAI21_X1 U6368 ( .B1(n6354), .B2(n5257), .A(n5227), .ZN(n5228) );
  AOI21_X1 U6369 ( .B1(n6391), .B2(n5259), .A(n5228), .ZN(n5229) );
  OAI21_X1 U6370 ( .B1(n5262), .B2(n5230), .A(n5229), .ZN(U3058) );
  INV_X1 U6371 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5234) );
  AOI22_X1 U6372 ( .A1(n6375), .A2(n5255), .B1(n6325), .B2(n6298), .ZN(n5231)
         );
  OAI21_X1 U6373 ( .B1(n6328), .B2(n5257), .A(n5231), .ZN(n5232) );
  AOI21_X1 U6374 ( .B1(n6376), .B2(n5259), .A(n5232), .ZN(n5233) );
  OAI21_X1 U6375 ( .B1(n5262), .B2(n5234), .A(n5233), .ZN(U3053) );
  INV_X1 U6376 ( .A(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5238) );
  AOI22_X1 U6377 ( .A1(n6381), .A2(n5255), .B1(n6335), .B2(n6298), .ZN(n5235)
         );
  OAI21_X1 U6378 ( .B1(n6338), .B2(n5257), .A(n5235), .ZN(n5236) );
  AOI21_X1 U6379 ( .B1(n6382), .B2(n5259), .A(n5236), .ZN(n5237) );
  OAI21_X1 U6380 ( .B1(n5262), .B2(n5238), .A(n5237), .ZN(U3055) );
  INV_X1 U6381 ( .A(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5242) );
  AOI22_X1 U6382 ( .A1(n6339), .A2(n5255), .B1(n6341), .B2(n6298), .ZN(n5239)
         );
  OAI21_X1 U6383 ( .B1(n6344), .B2(n5257), .A(n5239), .ZN(n5240) );
  AOI21_X1 U6384 ( .B1(n6340), .B2(n5259), .A(n5240), .ZN(n5241) );
  OAI21_X1 U6385 ( .B1(n5262), .B2(n5242), .A(n5241), .ZN(U3056) );
  INV_X1 U6386 ( .A(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5246) );
  AOI22_X1 U6387 ( .A1(n6356), .A2(n5255), .B1(n6360), .B2(n6298), .ZN(n5243)
         );
  OAI21_X1 U6388 ( .B1(n6364), .B2(n5257), .A(n5243), .ZN(n5244) );
  AOI21_X1 U6389 ( .B1(n6358), .B2(n5259), .A(n5244), .ZN(n5245) );
  OAI21_X1 U6390 ( .B1(n5262), .B2(n5246), .A(n5245), .ZN(U3059) );
  INV_X1 U6391 ( .A(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5250) );
  AOI22_X1 U6392 ( .A1(n6311), .A2(n5255), .B1(n6321), .B2(n6298), .ZN(n5247)
         );
  OAI21_X1 U6393 ( .B1(n6324), .B2(n5257), .A(n5247), .ZN(n5248) );
  AOI21_X1 U6394 ( .B1(n6312), .B2(n5259), .A(n5248), .ZN(n5249) );
  OAI21_X1 U6395 ( .B1(n5262), .B2(n5250), .A(n5249), .ZN(U3052) );
  INV_X1 U6396 ( .A(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5254) );
  AOI22_X1 U6397 ( .A1(n6329), .A2(n5255), .B1(n6331), .B2(n6298), .ZN(n5251)
         );
  OAI21_X1 U6398 ( .B1(n6334), .B2(n5257), .A(n5251), .ZN(n5252) );
  AOI21_X1 U6399 ( .B1(n6330), .B2(n5259), .A(n5252), .ZN(n5253) );
  OAI21_X1 U6400 ( .B1(n5262), .B2(n5254), .A(n5253), .ZN(U3054) );
  INV_X1 U6401 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5261) );
  AOI22_X1 U6402 ( .A1(n6345), .A2(n5255), .B1(n6347), .B2(n6298), .ZN(n5256)
         );
  OAI21_X1 U6403 ( .B1(n6350), .B2(n5257), .A(n5256), .ZN(n5258) );
  AOI21_X1 U6404 ( .B1(n6346), .B2(n5259), .A(n5258), .ZN(n5260) );
  OAI21_X1 U6405 ( .B1(n5262), .B2(n5261), .A(n5260), .ZN(U3057) );
  OAI21_X1 U6406 ( .B1(n5265), .B2(n5264), .A(n5263), .ZN(n5848) );
  INV_X1 U6407 ( .A(n5266), .ZN(n5269) );
  AOI21_X1 U6408 ( .B1(n5269), .B2(n5268), .A(n5267), .ZN(n5849) );
  AOI22_X1 U6409 ( .A1(n5849), .A2(n6563), .B1(EBX_REG_21__SCAN_IN), .B2(n6562), .ZN(n5270) );
  OAI21_X1 U6410 ( .B1(n5848), .B2(n6118), .A(n5270), .ZN(U2838) );
  OAI222_X1 U6411 ( .A1(n6118), .A2(n5883), .B1(n5271), .B2(n6123), .C1(n5765), 
        .C2(n5546), .ZN(U2839) );
  XNOR2_X1 U6412 ( .A(n5163), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5311)
         );
  XNOR2_X1 U6413 ( .A(n3013), .B(n5311), .ZN(n5955) );
  NAND2_X1 U6414 ( .A1(n5955), .A2(n6204), .ZN(n5279) );
  INV_X1 U6415 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5275) );
  OAI22_X1 U6416 ( .A1(n5651), .A2(n5275), .B1(n6216), .B2(n6493), .ZN(n5276)
         );
  AOI21_X1 U6417 ( .B1(n6177), .B2(n5277), .A(n5276), .ZN(n5278) );
  OAI211_X1 U6418 ( .C1(n5679), .C2(n5280), .A(n5279), .B(n5278), .ZN(U2973)
         );
  INV_X1 U6419 ( .A(n5281), .ZN(n5284) );
  NAND2_X1 U6420 ( .A1(n5286), .A2(n5282), .ZN(n5283) );
  NAND2_X1 U6421 ( .A1(n5284), .A2(n5283), .ZN(n6561) );
  AOI22_X1 U6422 ( .A1(n5301), .A2(DATAI_15_), .B1(n6130), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n5285) );
  OAI21_X1 U6423 ( .B1(n6561), .B2(n5867), .A(n5285), .ZN(U2876) );
  INV_X1 U6424 ( .A(n5286), .ZN(n5287) );
  AOI21_X1 U6425 ( .B1(n5289), .B2(n5288), .A(n5287), .ZN(n5321) );
  INV_X1 U6426 ( .A(n5321), .ZN(n5304) );
  OAI21_X1 U6427 ( .B1(n5342), .B2(n5290), .A(n6031), .ZN(n6017) );
  INV_X1 U6428 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6605) );
  OAI21_X1 U6429 ( .B1(n6493), .B2(n5291), .A(n6605), .ZN(n5299) );
  NAND2_X1 U6430 ( .A1(n5293), .A2(n5292), .ZN(n5294) );
  NAND2_X1 U6431 ( .A1(n5930), .A2(n5294), .ZN(n5948) );
  OAI22_X1 U6432 ( .A1(n5295), .A2(n6078), .B1(n6100), .B2(n5948), .ZN(n5296)
         );
  AOI211_X1 U6433 ( .C1(n3003), .C2(EBX_REG_14__SCAN_IN), .A(n5296), .B(n6081), 
        .ZN(n5297) );
  OAI21_X1 U6434 ( .B1(n5319), .B2(n6094), .A(n5297), .ZN(n5298) );
  AOI21_X1 U6435 ( .B1(n6017), .B2(n5299), .A(n5298), .ZN(n5300) );
  OAI21_X1 U6436 ( .B1(n5304), .B2(n6038), .A(n5300), .ZN(U2813) );
  AOI22_X1 U6437 ( .A1(n5301), .A2(DATAI_14_), .B1(n6130), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n5302) );
  OAI21_X1 U6438 ( .B1(n5304), .B2(n5867), .A(n5302), .ZN(U2877) );
  INV_X1 U6439 ( .A(EBX_REG_14__SCAN_IN), .ZN(n5303) );
  OAI222_X1 U6440 ( .A1(n5304), .A2(n6118), .B1(n6123), .B2(n5303), .C1(n5948), 
        .C2(n5546), .ZN(U2845) );
  NAND2_X1 U6441 ( .A1(n5263), .A2(n5306), .ZN(n5307) );
  NAND2_X1 U6442 ( .A1(n5611), .A2(n5307), .ZN(n5832) );
  INV_X1 U6443 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5310) );
  NOR2_X1 U6444 ( .A1(n5267), .A2(n5308), .ZN(n5309) );
  OR2_X1 U6445 ( .A1(n5730), .A2(n5309), .ZN(n5842) );
  OAI222_X1 U6446 ( .A1(n6118), .A2(n5832), .B1(n6123), .B2(n5310), .C1(n5842), 
        .C2(n5546), .ZN(U2837) );
  NAND2_X1 U6447 ( .A1(n5312), .A2(n5311), .ZN(n5314) );
  INV_X1 U6448 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n6571) );
  NAND2_X1 U6449 ( .A1(n5163), .A2(n6571), .ZN(n5313) );
  NAND2_X1 U6450 ( .A1(n5314), .A2(n5313), .ZN(n5356) );
  INV_X1 U6451 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5952) );
  INV_X1 U6452 ( .A(n5668), .ZN(n5316) );
  AND2_X1 U6453 ( .A1(n5163), .A2(n5952), .ZN(n5647) );
  NOR2_X1 U6454 ( .A1(n5316), .A2(n5647), .ZN(n5317) );
  XNOR2_X1 U6455 ( .A(n5315), .B(n5317), .ZN(n5950) );
  INV_X1 U6456 ( .A(n5950), .ZN(n5323) );
  AOI22_X1 U6457 ( .A1(n6199), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6260), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5318) );
  OAI21_X1 U6458 ( .B1(n6210), .B2(n5319), .A(n5318), .ZN(n5320) );
  AOI21_X1 U6459 ( .B1(n5321), .B2(n6205), .A(n5320), .ZN(n5322) );
  OAI21_X1 U6460 ( .B1(n5323), .B2(n6181), .A(n5322), .ZN(U2972) );
  XNOR2_X1 U6461 ( .A(n3015), .B(n5777), .ZN(n5325) );
  AOI22_X1 U6462 ( .A1(n5325), .A2(n4551), .B1(n5324), .B2(n5328), .ZN(n5327)
         );
  NAND2_X1 U6463 ( .A1(n5782), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n5326) );
  OAI21_X1 U6464 ( .B1(n5782), .B2(n5327), .A(n5326), .ZN(U3463) );
  INV_X1 U6465 ( .A(n5328), .ZN(n5338) );
  INV_X1 U6466 ( .A(n6105), .ZN(n6091) );
  NAND2_X1 U6467 ( .A1(n6206), .A2(n6091), .ZN(n5337) );
  OAI21_X1 U6468 ( .B1(n6084), .B2(REIP_REG_1__SCAN_IN), .A(n5329), .ZN(n6095)
         );
  OAI22_X1 U6469 ( .A1(n6094), .A2(n6209), .B1(n5330), .B2(n6078), .ZN(n5333)
         );
  INV_X1 U6470 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5331) );
  NOR3_X1 U6471 ( .A1(n6084), .A2(REIP_REG_2__SCAN_IN), .A3(n5331), .ZN(n5332)
         );
  AOI211_X1 U6472 ( .C1(EBX_REG_2__SCAN_IN), .C2(n3003), .A(n5333), .B(n5332), 
        .ZN(n5334) );
  OAI21_X1 U6473 ( .B1(n6276), .B2(n6100), .A(n5334), .ZN(n5335) );
  AOI21_X1 U6474 ( .B1(REIP_REG_2__SCAN_IN), .B2(n6095), .A(n5335), .ZN(n5336)
         );
  OAI211_X1 U6475 ( .C1(n5338), .C2(n6088), .A(n5337), .B(n5336), .ZN(U2825)
         );
  NOR2_X1 U6476 ( .A1(n6503), .A2(n5339), .ZN(n5834) );
  NAND3_X1 U6477 ( .A1(REIP_REG_22__SCAN_IN), .A2(REIP_REG_21__SCAN_IN), .A3(
        n5834), .ZN(n5825) );
  INV_X1 U6478 ( .A(REIP_REG_23__SCAN_IN), .ZN(n6506) );
  NOR2_X1 U6479 ( .A1(n5825), .A2(n6506), .ZN(n5808) );
  AND3_X1 U6480 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n5343) );
  NAND2_X1 U6481 ( .A1(n5808), .A2(n5343), .ZN(n5791) );
  NAND2_X1 U6482 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5348) );
  NOR3_X1 U6483 ( .A1(n5791), .A2(REIP_REG_29__SCAN_IN), .A3(n5348), .ZN(n5489) );
  INV_X1 U6484 ( .A(n5348), .ZN(n5345) );
  NAND3_X1 U6485 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5340) );
  OAI21_X1 U6486 ( .B1(n5341), .B2(n5340), .A(n6076), .ZN(n5824) );
  OAI21_X1 U6487 ( .B1(n5343), .B2(n5342), .A(n5824), .ZN(n5797) );
  INV_X1 U6488 ( .A(n5797), .ZN(n5344) );
  OAI21_X1 U6489 ( .B1(n6084), .B2(n5345), .A(n5344), .ZN(n5502) );
  NOR2_X1 U6490 ( .A1(n5489), .A2(n5502), .ZN(n5460) );
  INV_X1 U6491 ( .A(n5460), .ZN(n5354) );
  INV_X1 U6492 ( .A(REIP_REG_29__SCAN_IN), .ZN(n5347) );
  OR3_X1 U6493 ( .A1(n5791), .A2(n5348), .A3(n5347), .ZN(n5462) );
  INV_X1 U6494 ( .A(n5349), .ZN(n5378) );
  OAI22_X1 U6495 ( .A1(n6094), .A2(n5378), .B1(n5350), .B2(n6078), .ZN(n5352)
         );
  NOR2_X1 U6496 ( .A1(n6065), .A2(n4020), .ZN(n5351) );
  NAND3_X1 U6497 ( .A1(n3028), .A2(n3022), .A3(n3033), .ZN(n5353) );
  AOI21_X1 U6498 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5354), .A(n5353), .ZN(n5355) );
  OAI21_X1 U6499 ( .B1(n5550), .B2(n6038), .A(n5355), .ZN(U2797) );
  INV_X1 U6500 ( .A(n5356), .ZN(n5359) );
  INV_X1 U6501 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5938) );
  AND2_X1 U6502 ( .A1(n5163), .A2(n5928), .ZN(n5357) );
  NAND2_X1 U6503 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5396) );
  AND2_X1 U6504 ( .A1(n5163), .A2(n5396), .ZN(n5358) );
  NAND2_X1 U6505 ( .A1(n5359), .A2(n3025), .ZN(n5607) );
  INV_X1 U6506 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n6604) );
  INV_X1 U6507 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5759) );
  AND3_X1 U6508 ( .A1(n6604), .A2(n5759), .A3(n5928), .ZN(n5360) );
  XNOR2_X1 U6509 ( .A(n5163), .B(n5938), .ZN(n5670) );
  INV_X1 U6510 ( .A(n5670), .ZN(n5361) );
  NAND2_X1 U6511 ( .A1(n5607), .A2(n5364), .ZN(n5593) );
  NOR2_X1 U6512 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5365) );
  INV_X1 U6513 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5741) );
  INV_X1 U6514 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5735) );
  INV_X1 U6515 ( .A(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5722) );
  NAND4_X1 U6516 ( .A1(n5365), .A2(n5741), .A3(n5735), .A4(n5722), .ZN(n5366)
         );
  OAI21_X1 U6517 ( .B1(n5593), .B2(n5366), .A(n5891), .ZN(n5370) );
  AND2_X1 U6518 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5742) );
  AND2_X1 U6519 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5390) );
  NAND2_X1 U6520 ( .A1(n5742), .A2(n5390), .ZN(n5395) );
  NAND2_X1 U6521 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5397) );
  NOR2_X1 U6522 ( .A1(n5395), .A2(n5397), .ZN(n5368) );
  NAND2_X1 U6523 ( .A1(n5638), .A2(n5368), .ZN(n5369) );
  NAND2_X1 U6524 ( .A1(n5370), .A2(n5369), .ZN(n5588) );
  INV_X1 U6525 ( .A(n5588), .ZN(n5372) );
  INV_X1 U6526 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5714) );
  XNOR2_X1 U6527 ( .A(n5163), .B(n5714), .ZN(n5589) );
  NAND2_X1 U6528 ( .A1(n5163), .A2(n5714), .ZN(n5373) );
  NAND2_X1 U6529 ( .A1(n5561), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5573) );
  NAND2_X1 U6530 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5690) );
  NOR2_X2 U6531 ( .A1(n5573), .A2(n5690), .ZN(n5439) );
  NOR2_X1 U6532 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5692) );
  NAND2_X1 U6533 ( .A1(n5891), .A2(n5692), .ZN(n5436) );
  NOR3_X1 U6534 ( .A1(n5436), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5418) );
  AND2_X1 U6535 ( .A1(n5582), .A2(n5418), .ZN(n5374) );
  XNOR2_X1 U6536 ( .A(n5376), .B(n5375), .ZN(n5404) );
  NAND2_X1 U6537 ( .A1(n6260), .A2(REIP_REG_30__SCAN_IN), .ZN(n5401) );
  NAND2_X1 U6538 ( .A1(n6199), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5377)
         );
  OAI211_X1 U6539 ( .C1(n6210), .C2(n5378), .A(n5401), .B(n5377), .ZN(n5379)
         );
  AOI21_X1 U6540 ( .B1(n5380), .B2(n6205), .A(n5379), .ZN(n5381) );
  OAI21_X1 U6541 ( .B1(n5404), .B2(n6181), .A(n5381), .ZN(U2956) );
  AND2_X1 U6542 ( .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U6543 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5925) );
  NOR2_X1 U6544 ( .A1(n6223), .A2(n5382), .ZN(n5959) );
  INV_X1 U6545 ( .A(n5959), .ZN(n5941) );
  NOR2_X1 U6546 ( .A1(n6571), .A2(n5941), .ZN(n5945) );
  NAND2_X1 U6547 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5945), .ZN(n5922) );
  NOR2_X1 U6548 ( .A1(n5925), .A2(n5922), .ZN(n5385) );
  OAI221_X1 U6549 ( .B1(n5384), .B2(n5960), .C1(n5384), .C2(n5385), .A(n5383), 
        .ZN(n5757) );
  INV_X1 U6550 ( .A(n5742), .ZN(n5762) );
  OAI21_X1 U6551 ( .B1(n5762), .B2(n5396), .A(n5921), .ZN(n5388) );
  NAND2_X1 U6552 ( .A1(n5386), .A2(n5385), .ZN(n5758) );
  NAND2_X1 U6553 ( .A1(n6280), .A2(n5758), .ZN(n5387) );
  NAND2_X1 U6554 ( .A1(n5388), .A2(n5387), .ZN(n5389) );
  OR2_X1 U6555 ( .A1(n5757), .A2(n5389), .ZN(n5753) );
  INV_X1 U6556 ( .A(n5390), .ZN(n5391) );
  AND2_X1 U6557 ( .A1(n5921), .A2(n5391), .ZN(n5392) );
  NOR2_X1 U6558 ( .A1(n5753), .A2(n5392), .ZN(n5736) );
  OAI21_X1 U6559 ( .B1(n6287), .B2(n6280), .A(n5397), .ZN(n5393) );
  NAND2_X1 U6560 ( .A1(n5736), .A2(n5393), .ZN(n5726) );
  AND2_X1 U6561 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5399) );
  INV_X1 U6562 ( .A(n5399), .ZN(n5708) );
  AND2_X1 U6563 ( .A1(n5921), .A2(n5708), .ZN(n5394) );
  AOI21_X1 U6564 ( .B1(n5690), .B2(n5921), .A(n5703), .ZN(n5447) );
  OAI21_X1 U6565 ( .B1(n5681), .B2(n6228), .A(n5447), .ZN(n5680) );
  INV_X1 U6566 ( .A(n5395), .ZN(n5604) );
  NAND2_X1 U6567 ( .A1(n5945), .A2(n6211), .ZN(n5953) );
  NAND3_X1 U6568 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5934), .ZN(n5920) );
  NOR2_X2 U6569 ( .A1(n5396), .A2(n5920), .ZN(n5770) );
  INV_X1 U6570 ( .A(n5397), .ZN(n5398) );
  NAND2_X1 U6571 ( .A1(n5715), .A2(n5399), .ZN(n5700) );
  NOR2_X1 U6572 ( .A1(n5700), .A2(n5690), .ZN(n5682) );
  NAND3_X1 U6573 ( .A1(n5682), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5375), .ZN(n5400) );
  OAI211_X1 U6574 ( .C1(n5346), .C2(n6217), .A(n5401), .B(n5400), .ZN(n5402)
         );
  AOI21_X1 U6575 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5680), .A(n5402), 
        .ZN(n5403) );
  OAI21_X1 U6576 ( .B1(n5404), .B2(n5906), .A(n5403), .ZN(U2988) );
  AOI21_X1 U6577 ( .B1(n5407), .B2(n5405), .A(n5412), .ZN(n5415) );
  INV_X1 U6578 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n5414) );
  INV_X1 U6579 ( .A(n5406), .ZN(n5409) );
  NAND3_X1 U6580 ( .A1(n4067), .A2(n5407), .A3(n5414), .ZN(n5408) );
  OAI21_X1 U6581 ( .B1(n5410), .B2(n5409), .A(n5408), .ZN(n5411) );
  AOI21_X1 U6582 ( .B1(n6399), .B2(n5967), .A(n5411), .ZN(n5413) );
  OAI22_X1 U6583 ( .A1(n5415), .A2(n5414), .B1(n5413), .B2(n5412), .ZN(U3459)
         );
  INV_X1 U6584 ( .A(n5418), .ZN(n5419) );
  NOR3_X1 U6585 ( .A1(n5417), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5419), 
        .ZN(n5420) );
  AOI21_X1 U6586 ( .B1(n5439), .B2(n5681), .A(n5420), .ZN(n5421) );
  XNOR2_X1 U6587 ( .A(n5421), .B(n5685), .ZN(n5689) );
  NAND2_X1 U6588 ( .A1(n5452), .A2(n5422), .ZN(n5427) );
  AOI22_X1 U6589 ( .A1(n5424), .A2(EAX_REG_31__SCAN_IN), .B1(n5423), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5425) );
  INV_X1 U6590 ( .A(n5425), .ZN(n5426) );
  XNOR2_X2 U6591 ( .A(n5427), .B(n5426), .ZN(n5459) );
  NAND2_X1 U6592 ( .A1(n6260), .A2(REIP_REG_31__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U6593 ( .A1(n6199), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5428)
         );
  OAI211_X1 U6594 ( .C1(n6210), .C2(n5429), .A(n5684), .B(n5428), .ZN(n5430)
         );
  AOI21_X1 U6595 ( .B1(n5459), .B2(n6205), .A(n5430), .ZN(n5431) );
  OAI21_X1 U6596 ( .B1(n5689), .B2(n6181), .A(n5431), .ZN(U2955) );
  NAND3_X1 U6597 ( .A1(n5459), .A2(n5433), .A3(n5432), .ZN(n5435) );
  AOI22_X1 U6598 ( .A1(n6127), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6130), .ZN(n5434) );
  NAND2_X1 U6599 ( .A1(n5435), .A2(n5434), .ZN(U2860) );
  NOR2_X1 U6600 ( .A1(n5436), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5437)
         );
  NOR2_X1 U6601 ( .A1(n5439), .A2(n5438), .ZN(n5441) );
  INV_X1 U6602 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5440) );
  XNOR2_X1 U6603 ( .A(n5441), .B(n5440), .ZN(n5458) );
  MUX2_X1 U6604 ( .A(EBX_REG_29__SCAN_IN), .B(n5442), .S(n3956), .Z(n5443) );
  AOI21_X1 U6605 ( .B1(n5444), .B2(n6724), .A(n5443), .ZN(n5463) );
  XNOR2_X1 U6606 ( .A(n5445), .B(n5463), .ZN(n5517) );
  INV_X1 U6607 ( .A(n5682), .ZN(n5446) );
  NAND2_X1 U6608 ( .A1(n6260), .A2(REIP_REG_29__SCAN_IN), .ZN(n5455) );
  OAI21_X1 U6609 ( .B1(n5446), .B2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5455), 
        .ZN(n5449) );
  NOR2_X1 U6610 ( .A1(n5447), .A2(n5440), .ZN(n5448) );
  AOI211_X1 U6611 ( .C1(n6279), .C2(n5517), .A(n5449), .B(n5448), .ZN(n5450)
         );
  OAI21_X1 U6612 ( .B1(n5458), .B2(n5906), .A(n5450), .ZN(U2989) );
  AOI21_X1 U6613 ( .B1(n5453), .B2(n5493), .A(n5452), .ZN(n5484) );
  NAND2_X1 U6614 ( .A1(n6199), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5454)
         );
  OAI211_X1 U6615 ( .C1(n6210), .C2(n5485), .A(n5455), .B(n5454), .ZN(n5456)
         );
  AOI21_X1 U6616 ( .B1(n5484), .B2(n6205), .A(n5456), .ZN(n5457) );
  OAI21_X1 U6617 ( .B1(n5458), .B2(n6181), .A(n5457), .ZN(U2957) );
  INV_X1 U6618 ( .A(n5459), .ZN(n5483) );
  INV_X1 U6619 ( .A(REIP_REG_31__SCAN_IN), .ZN(n5480) );
  OAI21_X1 U6620 ( .B1(REIP_REG_30__SCAN_IN), .B2(n6084), .A(n5460), .ZN(n5461) );
  INV_X1 U6621 ( .A(n5461), .ZN(n5479) );
  INV_X1 U6622 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6519) );
  NAND3_X1 U6623 ( .A1(n5495), .A2(n5464), .A3(n5463), .ZN(n5465) );
  NAND2_X1 U6624 ( .A1(n5466), .A2(n5465), .ZN(n5471) );
  OAI22_X1 U6625 ( .A1(n5468), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n5467), .B2(EBX_REG_31__SCAN_IN), .ZN(n5469) );
  INV_X1 U6626 ( .A(n5469), .ZN(n5470) );
  XNOR2_X2 U6627 ( .A(n5471), .B(n5470), .ZN(n5514) );
  NAND3_X1 U6628 ( .A1(n5473), .A2(EBX_REG_31__SCAN_IN), .A3(n5472), .ZN(n5474) );
  OAI211_X1 U6629 ( .C1(n5476), .C2(n6078), .A(n5475), .B(n5474), .ZN(n5477)
         );
  INV_X1 U6630 ( .A(n5477), .ZN(n5478) );
  INV_X1 U6631 ( .A(n5481), .ZN(n5482) );
  OAI21_X1 U6632 ( .B1(n5483), .B2(n6038), .A(n5482), .ZN(U2796) );
  INV_X1 U6633 ( .A(n5484), .ZN(n5553) );
  NAND2_X1 U6634 ( .A1(n5517), .A2(n6086), .ZN(n5488) );
  INV_X1 U6635 ( .A(n5485), .ZN(n5486) );
  AOI22_X1 U6636 ( .A1(PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n6097), .B1(n6108), 
        .B2(n5486), .ZN(n5487) );
  OAI211_X1 U6637 ( .C1(n6724), .C2(n6065), .A(n5488), .B(n5487), .ZN(n5490)
         );
  AOI211_X1 U6638 ( .C1(REIP_REG_29__SCAN_IN), .C2(n5502), .A(n5490), .B(n5489), .ZN(n5491) );
  OAI21_X1 U6639 ( .B1(n5553), .B2(n6038), .A(n5491), .ZN(U2798) );
  OAI21_X1 U6640 ( .B1(n5492), .B2(n5494), .A(n5493), .ZN(n5567) );
  INV_X1 U6641 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6513) );
  NOR3_X1 U6642 ( .A1(n5791), .A2(REIP_REG_28__SCAN_IN), .A3(n6513), .ZN(n5501) );
  AOI21_X1 U6643 ( .B1(n5496), .B2(n5524), .A(n5495), .ZN(n5695) );
  INV_X1 U6644 ( .A(n5695), .ZN(n5499) );
  AOI22_X1 U6645 ( .A1(PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n6097), .B1(n6108), 
        .B2(n5566), .ZN(n5498) );
  NAND2_X1 U6646 ( .A1(n3003), .A2(EBX_REG_28__SCAN_IN), .ZN(n5497) );
  OAI211_X1 U6647 ( .C1(n5499), .C2(n6100), .A(n5498), .B(n5497), .ZN(n5500)
         );
  AOI211_X1 U6648 ( .C1(REIP_REG_28__SCAN_IN), .C2(n5502), .A(n5501), .B(n5500), .ZN(n5503) );
  OAI21_X1 U6649 ( .B1(n5567), .B2(n6038), .A(n5503), .ZN(U2799) );
  NAND2_X1 U6650 ( .A1(n5504), .A2(n6091), .ZN(n5513) );
  AOI22_X1 U6651 ( .A1(n6054), .A2(n5331), .B1(n3003), .B2(EBX_REG_1__SCAN_IN), 
        .ZN(n5512) );
  INV_X1 U6652 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5507) );
  NAND2_X1 U6653 ( .A1(n6108), .A2(n5507), .ZN(n5506) );
  NAND2_X1 U6654 ( .A1(n6077), .A2(REIP_REG_1__SCAN_IN), .ZN(n5505) );
  OAI211_X1 U6655 ( .C1(n5507), .C2(n6078), .A(n5506), .B(n5505), .ZN(n5508)
         );
  AOI21_X1 U6656 ( .B1(n6086), .B2(n5509), .A(n5508), .ZN(n5511) );
  NAND2_X1 U6657 ( .A1(n4104), .A2(n6102), .ZN(n5510) );
  NAND4_X1 U6658 ( .A1(n5513), .A2(n5512), .A3(n5511), .A4(n5510), .ZN(U2826)
         );
  INV_X1 U6659 ( .A(n5514), .ZN(n5516) );
  INV_X1 U6660 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5515) );
  OAI22_X1 U6661 ( .A1(n5516), .A2(n5546), .B1(n6123), .B2(n5515), .ZN(U2828)
         );
  INV_X1 U6662 ( .A(n5517), .ZN(n5518) );
  OAI222_X1 U6663 ( .A1(n6118), .A2(n5553), .B1(n6724), .B2(n6123), .C1(n5518), 
        .C2(n5546), .ZN(U2830) );
  AOI22_X1 U6664 ( .A1(n5695), .A2(n6563), .B1(EBX_REG_28__SCAN_IN), .B2(n6562), .ZN(n5519) );
  OAI21_X1 U6665 ( .B1(n5567), .B2(n6118), .A(n5519), .ZN(U2831) );
  AND2_X1 U6666 ( .A1(n5528), .A2(n5520), .ZN(n5521) );
  OR2_X1 U6667 ( .A1(n5521), .A2(n5492), .ZN(n5866) );
  INV_X1 U6668 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5525) );
  OR2_X1 U6669 ( .A1(n5531), .A2(n5522), .ZN(n5523) );
  AND2_X1 U6670 ( .A1(n5524), .A2(n5523), .ZN(n5702) );
  INV_X1 U6671 ( .A(n5702), .ZN(n5787) );
  OAI222_X1 U6672 ( .A1(n6118), .A2(n5866), .B1(n5525), .B2(n6123), .C1(n5787), 
        .C2(n5546), .ZN(U2832) );
  NAND2_X1 U6673 ( .A1(n5534), .A2(n5526), .ZN(n5527) );
  NAND2_X1 U6674 ( .A1(n5528), .A2(n5527), .ZN(n5794) );
  NOR2_X1 U6675 ( .A1(n5537), .A2(n5529), .ZN(n5530) );
  OR2_X1 U6676 ( .A1(n5531), .A2(n5530), .ZN(n5793) );
  INV_X1 U6677 ( .A(n5793), .ZN(n5532) );
  AOI22_X1 U6678 ( .A1(n5532), .A2(n6563), .B1(EBX_REG_26__SCAN_IN), .B2(n6562), .ZN(n5533) );
  OAI21_X1 U6679 ( .B1(n5794), .B2(n6118), .A(n5533), .ZN(U2833) );
  OAI21_X1 U6680 ( .B1(n5540), .B2(n5535), .A(n5534), .ZN(n5800) );
  INV_X1 U6681 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5806) );
  AND2_X1 U6682 ( .A1(n5545), .A2(n5536), .ZN(n5538) );
  OR2_X1 U6683 ( .A1(n5538), .A2(n5537), .ZN(n5812) );
  OAI222_X1 U6684 ( .A1(n6118), .A2(n5800), .B1(n6123), .B2(n5806), .C1(n5812), 
        .C2(n5546), .ZN(U2834) );
  INV_X1 U6685 ( .A(n5539), .ZN(n5542) );
  INV_X1 U6686 ( .A(n5612), .ZN(n5541) );
  AOI21_X1 U6687 ( .B1(n5542), .B2(n5541), .A(n5540), .ZN(n5818) );
  INV_X1 U6688 ( .A(n5818), .ZN(n5560) );
  INV_X1 U6689 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5547) );
  NAND2_X1 U6690 ( .A1(n5731), .A2(n5543), .ZN(n5544) );
  NAND2_X1 U6691 ( .A1(n5545), .A2(n5544), .ZN(n5823) );
  OAI222_X1 U6692 ( .A1(n6118), .A2(n5560), .B1(n6123), .B2(n5547), .C1(n5823), 
        .C2(n5546), .ZN(U2835) );
  AOI22_X1 U6693 ( .A1(n6127), .A2(DATAI_30_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6130), .ZN(n5549) );
  NAND2_X1 U6694 ( .A1(n6131), .A2(DATAI_14_), .ZN(n5548) );
  OAI211_X1 U6695 ( .C1(n5550), .C2(n5867), .A(n5549), .B(n5548), .ZN(U2861)
         );
  AOI22_X1 U6696 ( .A1(n6127), .A2(DATAI_29_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6130), .ZN(n5552) );
  NAND2_X1 U6697 ( .A1(n6131), .A2(DATAI_13_), .ZN(n5551) );
  OAI211_X1 U6698 ( .C1(n5553), .C2(n5867), .A(n5552), .B(n5551), .ZN(U2862)
         );
  AOI22_X1 U6699 ( .A1(n6127), .A2(DATAI_28_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6130), .ZN(n5555) );
  NAND2_X1 U6700 ( .A1(n6131), .A2(DATAI_12_), .ZN(n5554) );
  OAI211_X1 U6701 ( .C1(n5567), .C2(n5867), .A(n5555), .B(n5554), .ZN(U2863)
         );
  AOI22_X1 U6702 ( .A1(n6131), .A2(DATAI_10_), .B1(n6130), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U6703 ( .A1(n6127), .A2(DATAI_26_), .ZN(n5556) );
  OAI211_X1 U6704 ( .C1(n5794), .C2(n5867), .A(n5557), .B(n5556), .ZN(U2865)
         );
  AOI22_X1 U6705 ( .A1(n6131), .A2(DATAI_8_), .B1(n6130), .B2(
        EAX_REG_24__SCAN_IN), .ZN(n5559) );
  NAND2_X1 U6706 ( .A1(n6127), .A2(DATAI_24_), .ZN(n5558) );
  OAI211_X1 U6707 ( .C1(n5560), .C2(n5867), .A(n5559), .B(n5558), .ZN(U2867)
         );
  NAND2_X1 U6708 ( .A1(n5714), .A2(n5580), .ZN(n5707) );
  NOR3_X1 U6709 ( .A1(n5588), .A2(n5163), .A3(n5707), .ZN(n5571) );
  AOI21_X1 U6710 ( .B1(n5561), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5571), 
        .ZN(n5562) );
  AOI21_X1 U6711 ( .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5580), .A(n5562), 
        .ZN(n5563) );
  XNOR2_X1 U6712 ( .A(n5563), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5698)
         );
  AND2_X1 U6713 ( .A1(n6260), .A2(REIP_REG_28__SCAN_IN), .ZN(n5694) );
  NOR2_X1 U6714 ( .A1(n5651), .A2(n5564), .ZN(n5565) );
  AOI211_X1 U6715 ( .C1(n6177), .C2(n5566), .A(n5694), .B(n5565), .ZN(n5570)
         );
  INV_X1 U6716 ( .A(n5567), .ZN(n5568) );
  NAND2_X1 U6717 ( .A1(n5568), .A2(n6205), .ZN(n5569) );
  OAI211_X1 U6718 ( .C1(n5698), .C2(n6181), .A(n5570), .B(n5569), .ZN(U2958)
         );
  INV_X1 U6719 ( .A(n5571), .ZN(n5572) );
  NAND2_X1 U6720 ( .A1(n5573), .A2(n5572), .ZN(n5574) );
  XNOR2_X1 U6721 ( .A(n5574), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5706)
         );
  NAND2_X1 U6722 ( .A1(n6260), .A2(REIP_REG_27__SCAN_IN), .ZN(n5699) );
  OAI21_X1 U6723 ( .B1(n5651), .B2(n5575), .A(n5699), .ZN(n5577) );
  NOR2_X1 U6724 ( .A1(n5866), .A2(n5679), .ZN(n5576) );
  OAI21_X1 U6725 ( .B1(n5706), .B2(n6181), .A(n5579), .ZN(U2959) );
  XNOR2_X1 U6726 ( .A(n5163), .B(n5580), .ZN(n5581) );
  XNOR2_X1 U6727 ( .A(n3006), .B(n5581), .ZN(n5713) );
  NAND2_X1 U6728 ( .A1(n6260), .A2(REIP_REG_26__SCAN_IN), .ZN(n5710) );
  OAI21_X1 U6729 ( .B1(n5651), .B2(n5583), .A(n5710), .ZN(n5585) );
  NOR2_X1 U6730 ( .A1(n5794), .A2(n5679), .ZN(n5584) );
  AOI211_X1 U6731 ( .C1(n6177), .C2(n5792), .A(n5585), .B(n5584), .ZN(n5586)
         );
  OAI21_X1 U6732 ( .B1(n6181), .B2(n5713), .A(n5586), .ZN(U2960) );
  INV_X1 U6733 ( .A(n5417), .ZN(n5587) );
  AOI21_X1 U6734 ( .B1(n5589), .B2(n5588), .A(n5587), .ZN(n5720) );
  NAND2_X1 U6735 ( .A1(n6260), .A2(REIP_REG_25__SCAN_IN), .ZN(n5717) );
  OAI21_X1 U6736 ( .B1(n5651), .B2(n5802), .A(n5717), .ZN(n5591) );
  NOR2_X1 U6737 ( .A1(n5800), .A2(n5679), .ZN(n5590) );
  AOI211_X1 U6738 ( .C1(n6177), .C2(n5804), .A(n5591), .B(n5590), .ZN(n5592)
         );
  OAI21_X1 U6739 ( .B1(n5720), .B2(n6181), .A(n5592), .ZN(U2961) );
  BUF_X1 U6740 ( .A(n5593), .Z(n5639) );
  NAND2_X1 U6741 ( .A1(n5639), .A2(n5891), .ZN(n5595) );
  XNOR2_X1 U6742 ( .A(n5163), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5631)
         );
  INV_X1 U6743 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5596) );
  NOR2_X1 U6744 ( .A1(n5163), .A2(n5596), .ZN(n5597) );
  XNOR2_X1 U6745 ( .A(n5163), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5626)
         );
  NOR2_X1 U6746 ( .A1(n5163), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5618)
         );
  NAND2_X1 U6747 ( .A1(n5598), .A2(n5618), .ZN(n5605) );
  NAND3_X1 U6748 ( .A1(n5163), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5599) );
  XNOR2_X1 U6749 ( .A(n5600), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5728)
         );
  NAND2_X1 U6750 ( .A1(n6260), .A2(REIP_REG_24__SCAN_IN), .ZN(n5723) );
  NAND2_X1 U6751 ( .A1(n6199), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5601)
         );
  OAI211_X1 U6752 ( .C1(n6210), .C2(n5813), .A(n5723), .B(n5601), .ZN(n5602)
         );
  AOI21_X1 U6753 ( .B1(n5818), .B2(n6205), .A(n5602), .ZN(n5603) );
  OAI21_X1 U6754 ( .B1(n5728), .B2(n6181), .A(n5603), .ZN(U2962) );
  NAND2_X1 U6755 ( .A1(n5163), .A2(n5604), .ZN(n5606) );
  OAI21_X1 U6756 ( .B1(n3012), .B2(n5606), .A(n5605), .ZN(n5608) );
  XNOR2_X1 U6757 ( .A(n5608), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5740)
         );
  NAND2_X1 U6758 ( .A1(n6260), .A2(REIP_REG_23__SCAN_IN), .ZN(n5733) );
  OAI21_X1 U6759 ( .B1(n5651), .B2(n5609), .A(n5733), .ZN(n5615) );
  AND2_X1 U6760 ( .A1(n5611), .A2(n5610), .ZN(n5613) );
  OR2_X1 U6761 ( .A1(n5613), .A2(n5612), .ZN(n5829) );
  NOR2_X1 U6762 ( .A1(n5829), .A2(n5679), .ZN(n5614) );
  AOI211_X1 U6763 ( .C1(n6177), .C2(n5616), .A(n5615), .B(n5614), .ZN(n5617)
         );
  OAI21_X1 U6764 ( .B1(n5740), .B2(n6181), .A(n5617), .ZN(U2963) );
  AOI21_X1 U6765 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5163), .A(n5618), 
        .ZN(n5619) );
  XNOR2_X1 U6766 ( .A(n5620), .B(n5619), .ZN(n5749) );
  NAND2_X1 U6767 ( .A1(n6260), .A2(REIP_REG_22__SCAN_IN), .ZN(n5744) );
  OAI21_X1 U6768 ( .B1(n5651), .B2(n5838), .A(n5744), .ZN(n5622) );
  NOR2_X1 U6769 ( .A1(n5832), .A2(n5679), .ZN(n5621) );
  AOI211_X1 U6770 ( .C1(n6177), .C2(n5835), .A(n5622), .B(n5621), .ZN(n5623)
         );
  OAI21_X1 U6771 ( .B1(n5749), .B2(n6181), .A(n5623), .ZN(U2964) );
  OAI21_X1 U6772 ( .B1(n5626), .B2(n5625), .A(n5624), .ZN(n5750) );
  NAND2_X1 U6773 ( .A1(n5750), .A2(n6204), .ZN(n5630) );
  INV_X1 U6774 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5627) );
  NOR2_X1 U6775 ( .A1(n6216), .A2(n5627), .ZN(n5752) );
  NOR2_X1 U6776 ( .A1(n6210), .A2(n5852), .ZN(n5628) );
  AOI211_X1 U6777 ( .C1(n6199), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5752), 
        .B(n5628), .ZN(n5629) );
  OAI211_X1 U6778 ( .C1(n5679), .C2(n5848), .A(n5630), .B(n5629), .ZN(U2965)
         );
  XNOR2_X1 U6779 ( .A(n5632), .B(n5631), .ZN(n5768) );
  NAND2_X1 U6780 ( .A1(n6260), .A2(REIP_REG_20__SCAN_IN), .ZN(n5764) );
  OAI21_X1 U6781 ( .B1(n5651), .B2(n5633), .A(n5764), .ZN(n5635) );
  NOR2_X1 U6782 ( .A1(n5883), .A2(n5679), .ZN(n5634) );
  AOI211_X1 U6783 ( .C1(n6177), .C2(n5636), .A(n5635), .B(n5634), .ZN(n5637)
         );
  OAI21_X1 U6784 ( .B1(n5768), .B2(n6181), .A(n5637), .ZN(U2966) );
  INV_X1 U6785 ( .A(n5638), .ZN(n5640) );
  OAI21_X1 U6786 ( .B1(n5640), .B2(n5769), .A(n5639), .ZN(n5641) );
  XNOR2_X1 U6787 ( .A(n5641), .B(n5163), .ZN(n5776) );
  NAND2_X1 U6788 ( .A1(n6260), .A2(REIP_REG_19__SCAN_IN), .ZN(n5772) );
  NAND2_X1 U6789 ( .A1(n6199), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5642)
         );
  OAI211_X1 U6790 ( .C1(n6210), .C2(n5862), .A(n5772), .B(n5642), .ZN(n5643)
         );
  AOI21_X1 U6791 ( .B1(n5887), .B2(n6205), .A(n5643), .ZN(n5644) );
  OAI21_X1 U6792 ( .B1(n5776), .B2(n6181), .A(n5644), .ZN(U2967) );
  OR2_X1 U6793 ( .A1(n5315), .A2(n5645), .ZN(n5646) );
  AND2_X1 U6794 ( .A1(n5646), .A2(n5658), .ZN(n5890) );
  NOR3_X1 U6795 ( .A1(n5890), .A2(n5891), .A3(n5759), .ZN(n5898) );
  OR2_X1 U6796 ( .A1(n5315), .A2(n5647), .ZN(n5669) );
  NAND2_X1 U6797 ( .A1(n5669), .A2(n5648), .ZN(n5673) );
  OR2_X1 U6798 ( .A1(n5163), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5893)
         );
  NOR3_X1 U6799 ( .A1(n5673), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .A3(n5893), 
        .ZN(n5895) );
  NOR2_X1 U6800 ( .A1(n5898), .A2(n5895), .ZN(n5649) );
  XNOR2_X1 U6801 ( .A(n5649), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5908)
         );
  NAND2_X1 U6802 ( .A1(n5908), .A2(n6204), .ZN(n5655) );
  OAI22_X1 U6803 ( .A1(n5651), .A2(n5650), .B1(n6216), .B2(n6500), .ZN(n5652)
         );
  AOI21_X1 U6804 ( .B1(n6177), .B2(n5653), .A(n5652), .ZN(n5654) );
  OAI211_X1 U6805 ( .C1(n5679), .C2(n5656), .A(n5655), .B(n5654), .ZN(U2968)
         );
  MUX2_X1 U6806 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .B(n5928), .S(n5163), 
        .Z(n5662) );
  INV_X1 U6807 ( .A(n5662), .ZN(n5661) );
  OR2_X1 U6808 ( .A1(n5315), .A2(n5657), .ZN(n5659) );
  AND2_X1 U6809 ( .A1(n5659), .A2(n5658), .ZN(n5660) );
  MUX2_X1 U6810 ( .A(n5662), .B(n5661), .S(n5660), .Z(n5924) );
  INV_X1 U6811 ( .A(n5924), .ZN(n5667) );
  INV_X1 U6812 ( .A(n5663), .ZN(n6129) );
  AOI22_X1 U6813 ( .A1(n6199), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n6260), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5664) );
  OAI21_X1 U6814 ( .B1(n6012), .B2(n6210), .A(n5664), .ZN(n5665) );
  AOI21_X1 U6815 ( .B1(n6129), .B2(n6205), .A(n5665), .ZN(n5666) );
  OAI21_X1 U6816 ( .B1(n5667), .B2(n6181), .A(n5666), .ZN(U2970) );
  NAND2_X1 U6817 ( .A1(n5669), .A2(n5668), .ZN(n5671) );
  NAND2_X1 U6818 ( .A1(n5671), .A2(n5670), .ZN(n5672) );
  NAND2_X1 U6819 ( .A1(n5673), .A2(n5672), .ZN(n5935) );
  NAND2_X1 U6820 ( .A1(n5935), .A2(n6204), .ZN(n5678) );
  INV_X1 U6821 ( .A(REIP_REG_15__SCAN_IN), .ZN(n5674) );
  NOR2_X1 U6822 ( .A1(n6216), .A2(n5674), .ZN(n5933) );
  NOR2_X1 U6823 ( .A1(n5675), .A2(n6210), .ZN(n5676) );
  AOI211_X1 U6824 ( .C1(n6199), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5933), 
        .B(n5676), .ZN(n5677) );
  OAI211_X1 U6825 ( .C1(n5679), .C2(n6561), .A(n5678), .B(n5677), .ZN(U2971)
         );
  INV_X1 U6826 ( .A(n5680), .ZN(n5686) );
  NAND3_X1 U6827 ( .A1(n5682), .A2(n5681), .A3(n5685), .ZN(n5683) );
  OAI211_X1 U6828 ( .C1(n5686), .C2(n5685), .A(n5684), .B(n5683), .ZN(n5687)
         );
  AOI21_X1 U6829 ( .B1(n5514), .B2(n6279), .A(n5687), .ZN(n5688) );
  OAI21_X1 U6830 ( .B1(n5689), .B2(n5906), .A(n5688), .ZN(U2987) );
  INV_X1 U6831 ( .A(n5690), .ZN(n5691) );
  NOR3_X1 U6832 ( .A1(n5700), .A2(n5692), .A3(n5691), .ZN(n5693) );
  AOI211_X1 U6833 ( .C1(n5695), .C2(n6279), .A(n5694), .B(n5693), .ZN(n5697)
         );
  NAND2_X1 U6834 ( .A1(n5703), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5696) );
  OAI211_X1 U6835 ( .C1(n5698), .C2(n5906), .A(n5697), .B(n5696), .ZN(U2990)
         );
  OAI21_X1 U6836 ( .B1(n5700), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5699), 
        .ZN(n5701) );
  AOI21_X1 U6837 ( .B1(n5702), .B2(n6279), .A(n5701), .ZN(n5705) );
  NAND2_X1 U6838 ( .A1(n5703), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5704) );
  OAI211_X1 U6839 ( .C1(n5706), .C2(n5906), .A(n5705), .B(n5704), .ZN(U2991)
         );
  NAND3_X1 U6840 ( .A1(n5715), .A2(n5708), .A3(n5707), .ZN(n5709) );
  OAI211_X1 U6841 ( .C1(n5793), .C2(n6217), .A(n5710), .B(n5709), .ZN(n5711)
         );
  AOI21_X1 U6842 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5726), .A(n5711), 
        .ZN(n5712) );
  OAI21_X1 U6843 ( .B1(n5713), .B2(n5906), .A(n5712), .ZN(U2992) );
  NAND2_X1 U6844 ( .A1(n5715), .A2(n5714), .ZN(n5716) );
  OAI211_X1 U6845 ( .C1(n5812), .C2(n6217), .A(n5717), .B(n5716), .ZN(n5718)
         );
  AOI21_X1 U6846 ( .B1(INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n5726), .A(n5718), 
        .ZN(n5719) );
  OAI21_X1 U6847 ( .B1(n5720), .B2(n5906), .A(n5719), .ZN(U2993) );
  INV_X1 U6848 ( .A(n5721), .ZN(n5734) );
  OAI21_X1 U6849 ( .B1(n5734), .B2(n5735), .A(n5722), .ZN(n5725) );
  OAI21_X1 U6850 ( .B1(n5823), .B2(n6217), .A(n5723), .ZN(n5724) );
  AOI21_X1 U6851 ( .B1(n5726), .B2(n5725), .A(n5724), .ZN(n5727) );
  OAI21_X1 U6852 ( .B1(n5728), .B2(n5906), .A(n5727), .ZN(U2994) );
  OR2_X1 U6853 ( .A1(n5730), .A2(n5729), .ZN(n5732) );
  AND2_X1 U6854 ( .A1(n5732), .A2(n5731), .ZN(n5863) );
  OAI21_X1 U6855 ( .B1(INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n5734), .A(n5733), 
        .ZN(n5738) );
  NOR2_X1 U6856 ( .A1(n5736), .A2(n5735), .ZN(n5737) );
  AOI211_X1 U6857 ( .C1(n6279), .C2(n5863), .A(n5738), .B(n5737), .ZN(n5739)
         );
  OAI21_X1 U6858 ( .B1(n5740), .B2(n5906), .A(n5739), .ZN(U2995) );
  NAND4_X1 U6859 ( .A1(n5770), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n5742), .A4(n5741), .ZN(n5743) );
  OAI211_X1 U6860 ( .C1(n5842), .C2(n6217), .A(n5744), .B(n5743), .ZN(n5745)
         );
  INV_X1 U6861 ( .A(n5745), .ZN(n5748) );
  INV_X1 U6862 ( .A(n5770), .ZN(n5746) );
  NOR3_X1 U6863 ( .A1(n5746), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n5762), 
        .ZN(n5751) );
  OAI21_X1 U6864 ( .B1(n5753), .B2(n5751), .A(INSTADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n5747) );
  OAI211_X1 U6865 ( .C1(n5749), .C2(n5906), .A(n5748), .B(n5747), .ZN(U2996)
         );
  INV_X1 U6866 ( .A(n5750), .ZN(n5756) );
  AOI211_X1 U6867 ( .C1(n5849), .C2(n6279), .A(n5752), .B(n5751), .ZN(n5755)
         );
  NAND2_X1 U6868 ( .A1(n5753), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5754) );
  OAI211_X1 U6869 ( .C1(n5756), .C2(n5906), .A(n5755), .B(n5754), .ZN(U2997)
         );
  INV_X1 U6870 ( .A(n6287), .ZN(n5760) );
  AOI221_X1 U6871 ( .B1(n5759), .B2(n6280), .C1(n5758), .C2(n6280), .A(n5757), 
        .ZN(n5912) );
  OAI21_X1 U6872 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5760), .A(n5912), 
        .ZN(n5905) );
  INV_X1 U6873 ( .A(n5905), .ZN(n5761) );
  OAI21_X1 U6874 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n6228), .A(n5761), 
        .ZN(n5774) );
  OAI211_X1 U6875 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5770), .B(n5762), .ZN(n5763) );
  OAI211_X1 U6876 ( .C1(n5765), .C2(n6217), .A(n5764), .B(n5763), .ZN(n5766)
         );
  AOI21_X1 U6877 ( .B1(n5774), .B2(INSTADDRPOINTER_REG_20__SCAN_IN), .A(n5766), 
        .ZN(n5767) );
  OAI21_X1 U6878 ( .B1(n5768), .B2(n5906), .A(n5767), .ZN(U2998) );
  NAND2_X1 U6879 ( .A1(n5770), .A2(n5769), .ZN(n5771) );
  OAI211_X1 U6880 ( .C1(n5857), .C2(n6217), .A(n5772), .B(n5771), .ZN(n5773)
         );
  AOI21_X1 U6881 ( .B1(n5774), .B2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n5773), 
        .ZN(n5775) );
  OAI21_X1 U6882 ( .B1(n5776), .B2(n5906), .A(n5775), .ZN(U2999) );
  OAI211_X1 U6883 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n5778), .A(n5777), .B(
        n4551), .ZN(n5779) );
  OAI21_X1 U6884 ( .B1(n5781), .B2(n5780), .A(n5779), .ZN(n5783) );
  MUX2_X1 U6885 ( .A(n5783), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(n5782), 
        .Z(U3464) );
  AND2_X1 U6886 ( .A1(n6163), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI22_X1 U6887 ( .A1(EBX_REG_27__SCAN_IN), .A2(n3003), .B1(
        PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n6097), .ZN(n5784) );
  OAI21_X1 U6888 ( .B1(n5785), .B2(n6094), .A(n5784), .ZN(n5786) );
  AOI21_X1 U6889 ( .B1(REIP_REG_27__SCAN_IN), .B2(n5797), .A(n5786), .ZN(n5790) );
  OAI22_X1 U6890 ( .A1(n5866), .A2(n6038), .B1(n5787), .B2(n6100), .ZN(n5788)
         );
  INV_X1 U6891 ( .A(n5788), .ZN(n5789) );
  OAI211_X1 U6892 ( .C1(REIP_REG_27__SCAN_IN), .C2(n5791), .A(n5790), .B(n5789), .ZN(U2800) );
  AOI22_X1 U6893 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6097), .B1(n5792), 
        .B2(n6108), .ZN(n5799) );
  INV_X1 U6894 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6510) );
  NAND2_X1 U6895 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5808), .ZN(n5801) );
  INV_X1 U6896 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6512) );
  OAI21_X1 U6897 ( .B1(n6510), .B2(n5801), .A(n6512), .ZN(n5796) );
  OAI22_X1 U6898 ( .A1(n5794), .A2(n6038), .B1(n5793), .B2(n6100), .ZN(n5795)
         );
  AOI21_X1 U6899 ( .B1(n5797), .B2(n5796), .A(n5795), .ZN(n5798) );
  OAI211_X1 U6900 ( .C1(n6704), .C2(n6065), .A(n5799), .B(n5798), .ZN(U2801)
         );
  INV_X1 U6901 ( .A(n5800), .ZN(n5871) );
  OAI22_X1 U6902 ( .A1(n6078), .A2(n5802), .B1(REIP_REG_25__SCAN_IN), .B2(
        n5801), .ZN(n5803) );
  AOI21_X1 U6903 ( .B1(n5804), .B2(n6108), .A(n5803), .ZN(n5805) );
  OAI21_X1 U6904 ( .B1(n6065), .B2(n5806), .A(n5805), .ZN(n5807) );
  AOI21_X1 U6905 ( .B1(n5871), .B2(n6073), .A(n5807), .ZN(n5811) );
  INV_X1 U6906 ( .A(n5824), .ZN(n5809) );
  INV_X1 U6907 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6508) );
  AND2_X1 U6908 ( .A1(n6508), .A2(n5808), .ZN(n5820) );
  OAI21_X1 U6909 ( .B1(n5809), .B2(n5820), .A(REIP_REG_25__SCAN_IN), .ZN(n5810) );
  OAI211_X1 U6910 ( .C1(n6100), .C2(n5812), .A(n5811), .B(n5810), .ZN(U2802)
         );
  INV_X1 U6911 ( .A(n5813), .ZN(n5814) );
  AOI22_X1 U6912 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n6097), .B1(n6108), 
        .B2(n5814), .ZN(n5816) );
  NAND2_X1 U6913 ( .A1(n3003), .A2(EBX_REG_24__SCAN_IN), .ZN(n5815) );
  OAI211_X1 U6914 ( .C1(n5824), .C2(n6508), .A(n5816), .B(n5815), .ZN(n5817)
         );
  AOI21_X1 U6915 ( .B1(n5818), .B2(n6073), .A(n5817), .ZN(n5819) );
  INV_X1 U6916 ( .A(n5819), .ZN(n5821) );
  NOR2_X1 U6917 ( .A1(n5821), .A2(n5820), .ZN(n5822) );
  OAI21_X1 U6918 ( .B1(n5823), .B2(n6100), .A(n5822), .ZN(U2803) );
  AOI21_X1 U6919 ( .B1(n6506), .B2(n5825), .A(n5824), .ZN(n5828) );
  OAI22_X1 U6920 ( .A1(n5609), .A2(n6078), .B1(n5826), .B2(n6094), .ZN(n5827)
         );
  AOI211_X1 U6921 ( .C1(n3003), .C2(EBX_REG_23__SCAN_IN), .A(n5828), .B(n5827), 
        .ZN(n5831) );
  AOI22_X1 U6922 ( .A1(n5874), .A2(n6073), .B1(n5863), .B2(n6086), .ZN(n5830)
         );
  NAND2_X1 U6923 ( .A1(n5831), .A2(n5830), .ZN(U2804) );
  INV_X1 U6924 ( .A(n5832), .ZN(n5877) );
  NAND2_X1 U6925 ( .A1(n5834), .A2(n5627), .ZN(n5843) );
  INV_X1 U6926 ( .A(REIP_REG_22__SCAN_IN), .ZN(n5833) );
  AOI21_X1 U6927 ( .B1(n5844), .B2(n5843), .A(n5833), .ZN(n5840) );
  NAND3_X1 U6928 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5834), .A3(n5833), .ZN(
        n5837) );
  AOI22_X1 U6929 ( .A1(EBX_REG_22__SCAN_IN), .A2(n3003), .B1(n5835), .B2(n6108), .ZN(n5836) );
  OAI211_X1 U6930 ( .C1(n5838), .C2(n6078), .A(n5837), .B(n5836), .ZN(n5839)
         );
  AOI211_X1 U6931 ( .C1(n5877), .C2(n6073), .A(n5840), .B(n5839), .ZN(n5841)
         );
  OAI21_X1 U6932 ( .B1(n5842), .B2(n6100), .A(n5841), .ZN(U2805) );
  INV_X1 U6933 ( .A(n5843), .ZN(n5847) );
  INV_X1 U6934 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5845) );
  OAI22_X1 U6935 ( .A1(n5845), .A2(n6078), .B1(n5627), .B2(n5844), .ZN(n5846)
         );
  AOI211_X1 U6936 ( .C1(n3003), .C2(EBX_REG_21__SCAN_IN), .A(n5847), .B(n5846), 
        .ZN(n5851) );
  INV_X1 U6937 ( .A(n5848), .ZN(n5880) );
  AOI22_X1 U6938 ( .A1(n5880), .A2(n6073), .B1(n5849), .B2(n6086), .ZN(n5850)
         );
  OAI211_X1 U6939 ( .C1(n5852), .C2(n6094), .A(n5851), .B(n5850), .ZN(U2806)
         );
  INV_X1 U6940 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5856) );
  XOR2_X1 U6941 ( .A(REIP_REG_19__SCAN_IN), .B(REIP_REG_18__SCAN_IN), .Z(n5853) );
  AOI22_X1 U6942 ( .A1(REIP_REG_19__SCAN_IN), .A2(n5997), .B1(n5854), .B2(
        n5853), .ZN(n5855) );
  OAI211_X1 U6943 ( .C1(n6078), .C2(n5856), .A(n5855), .B(n6070), .ZN(n5860)
         );
  INV_X1 U6944 ( .A(n5887), .ZN(n5858) );
  OAI22_X1 U6945 ( .A1(n5858), .A2(n6038), .B1(n5857), .B2(n6100), .ZN(n5859)
         );
  AOI211_X1 U6946 ( .C1(EBX_REG_19__SCAN_IN), .C2(n3003), .A(n5860), .B(n5859), 
        .ZN(n5861) );
  OAI21_X1 U6947 ( .B1(n5862), .B2(n6094), .A(n5861), .ZN(U2808) );
  AOI22_X1 U6948 ( .A1(n5874), .A2(n3906), .B1(n5863), .B2(n6563), .ZN(n5864)
         );
  OAI21_X1 U6949 ( .B1(n6123), .B2(n5865), .A(n5864), .ZN(U2836) );
  INV_X1 U6950 ( .A(n5866), .ZN(n5868) );
  AOI22_X1 U6951 ( .A1(n5868), .A2(n6128), .B1(n6127), .B2(DATAI_27_), .ZN(
        n5870) );
  AOI22_X1 U6952 ( .A1(n6131), .A2(DATAI_11_), .B1(n6130), .B2(
        EAX_REG_27__SCAN_IN), .ZN(n5869) );
  NAND2_X1 U6953 ( .A1(n5870), .A2(n5869), .ZN(U2864) );
  AOI22_X1 U6954 ( .A1(n5871), .A2(n6128), .B1(n6127), .B2(DATAI_25_), .ZN(
        n5873) );
  AOI22_X1 U6955 ( .A1(n6131), .A2(DATAI_9_), .B1(n6130), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n5872) );
  NAND2_X1 U6956 ( .A1(n5873), .A2(n5872), .ZN(U2866) );
  AOI22_X1 U6957 ( .A1(n5874), .A2(n6128), .B1(n6127), .B2(DATAI_23_), .ZN(
        n5876) );
  AOI22_X1 U6958 ( .A1(n6131), .A2(DATAI_7_), .B1(n6130), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n5875) );
  NAND2_X1 U6959 ( .A1(n5876), .A2(n5875), .ZN(U2868) );
  AOI22_X1 U6960 ( .A1(n5877), .A2(n6128), .B1(n6127), .B2(DATAI_22_), .ZN(
        n5879) );
  AOI22_X1 U6961 ( .A1(n6131), .A2(DATAI_6_), .B1(n6130), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5878) );
  NAND2_X1 U6962 ( .A1(n5879), .A2(n5878), .ZN(U2869) );
  AOI22_X1 U6963 ( .A1(n5880), .A2(n6128), .B1(n6127), .B2(DATAI_21_), .ZN(
        n5882) );
  AOI22_X1 U6964 ( .A1(n6131), .A2(DATAI_5_), .B1(n6130), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5881) );
  NAND2_X1 U6965 ( .A1(n5882), .A2(n5881), .ZN(U2870) );
  INV_X1 U6966 ( .A(n5883), .ZN(n5884) );
  AOI22_X1 U6967 ( .A1(n5884), .A2(n6128), .B1(n6127), .B2(DATAI_20_), .ZN(
        n5886) );
  AOI22_X1 U6968 ( .A1(n6131), .A2(DATAI_4_), .B1(n6130), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U6969 ( .A1(n5886), .A2(n5885), .ZN(U2871) );
  AOI22_X1 U6970 ( .A1(n5887), .A2(n6128), .B1(n6127), .B2(DATAI_19_), .ZN(
        n5889) );
  AOI22_X1 U6971 ( .A1(n6131), .A2(DATAI_3_), .B1(n6130), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U6972 ( .A1(n5889), .A2(n5888), .ZN(U2872) );
  AOI22_X1 U6973 ( .A1(n6277), .A2(REIP_REG_17__SCAN_IN), .B1(n6199), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5904) );
  INV_X1 U6974 ( .A(n5890), .ZN(n5894) );
  INV_X1 U6975 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5928) );
  NAND2_X1 U6976 ( .A1(n5891), .A2(n5928), .ZN(n5892) );
  AOI22_X1 U6977 ( .A1(n5894), .A2(n5893), .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5892), .ZN(n5897) );
  INV_X1 U6978 ( .A(n5895), .ZN(n5896) );
  OAI21_X1 U6979 ( .B1(n5898), .B2(n5897), .A(n5896), .ZN(n5917) );
  NAND2_X1 U6980 ( .A1(n5900), .A2(n5899), .ZN(n5901) );
  AOI22_X1 U6981 ( .A1(n5917), .A2(n6204), .B1(n6205), .B2(n6124), .ZN(n5903)
         );
  OAI211_X1 U6982 ( .C1(n6210), .C2(n6003), .A(n5904), .B(n5903), .ZN(U2969)
         );
  NAND2_X1 U6983 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n6604), .ZN(n5911) );
  AOI22_X1 U6984 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5905), .B1(n6277), .B2(REIP_REG_18__SCAN_IN), .ZN(n5910) );
  AOI22_X1 U6985 ( .A1(n5908), .A2(n6284), .B1(n6279), .B2(n5907), .ZN(n5909)
         );
  OAI211_X1 U6986 ( .C1(n5920), .C2(n5911), .A(n5910), .B(n5909), .ZN(U3000)
         );
  INV_X1 U6987 ( .A(n5912), .ZN(n5913) );
  AOI22_X1 U6988 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5913), .B1(n6277), .B2(REIP_REG_17__SCAN_IN), .ZN(n5919) );
  NAND2_X1 U6989 ( .A1(n5141), .A2(n5914), .ZN(n5915) );
  AND2_X1 U6990 ( .A1(n5916), .A2(n5915), .ZN(n6113) );
  AOI22_X1 U6991 ( .A1(n5917), .A2(n6284), .B1(n6279), .B2(n6113), .ZN(n5918)
         );
  OAI211_X1 U6992 ( .C1(INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n5920), .A(n5919), .B(n5918), .ZN(U3001) );
  AOI21_X1 U6993 ( .B1(n5922), .B2(n5921), .A(n6214), .ZN(n5939) );
  OAI22_X1 U6994 ( .A1(n6016), .A2(n6217), .B1(n6497), .B2(n6216), .ZN(n5923)
         );
  AOI21_X1 U6995 ( .B1(n5924), .B2(n6284), .A(n5923), .ZN(n5927) );
  OAI211_X1 U6996 ( .C1(INSTADDRPOINTER_REG_15__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .A(n5934), .B(n5925), .ZN(n5926) );
  OAI211_X1 U6997 ( .C1(n5939), .C2(n5928), .A(n5927), .B(n5926), .ZN(U3002)
         );
  AND2_X1 U6998 ( .A1(n5930), .A2(n5929), .ZN(n5931) );
  NOR2_X1 U6999 ( .A1(n5932), .A2(n5931), .ZN(n6564) );
  AOI21_X1 U7000 ( .B1(n6564), .B2(n6279), .A(n5933), .ZN(n5937) );
  AOI22_X1 U7001 ( .A1(n5935), .A2(n6284), .B1(n5934), .B2(n5938), .ZN(n5936)
         );
  OAI211_X1 U7002 ( .C1(n5939), .C2(n5938), .A(n5937), .B(n5936), .ZN(U3003)
         );
  NAND3_X1 U7003 ( .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n5940), .A3(n5960), 
        .ZN(n5942) );
  AOI211_X1 U7004 ( .C1(n5943), .C2(n5942), .A(INSTADDRPOINTER_REG_13__SCAN_IN), .B(n5941), .ZN(n5958) );
  OAI22_X1 U7005 ( .A1(n5959), .A2(n5946), .B1(n5945), .B2(n5944), .ZN(n5947)
         );
  NOR3_X1 U7006 ( .A1(n5958), .A2(n6214), .A3(n5947), .ZN(n5956) );
  OAI22_X1 U7007 ( .A1(n5948), .A2(n6217), .B1(n6605), .B2(n6216), .ZN(n5949)
         );
  AOI21_X1 U7008 ( .B1(n5950), .B2(n6284), .A(n5949), .ZN(n5951) );
  OAI221_X1 U7009 ( .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5953), .C1(
        n5952), .C2(n5956), .A(n5951), .ZN(U3004) );
  AOI22_X1 U7010 ( .A1(n5955), .A2(n6284), .B1(n6279), .B2(n5954), .ZN(n5965)
         );
  NAND2_X1 U7011 ( .A1(n6277), .A2(REIP_REG_13__SCAN_IN), .ZN(n5964) );
  INV_X1 U7012 ( .A(n5956), .ZN(n5957) );
  OAI21_X1 U7013 ( .B1(INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n5958), .A(n5957), 
        .ZN(n5963) );
  NAND4_X1 U7014 ( .A1(n5961), .A2(n5960), .A3(n5959), .A4(n6571), .ZN(n5962)
         );
  NAND4_X1 U7015 ( .A1(n5965), .A2(n5964), .A3(n5963), .A4(n5962), .ZN(U3005)
         );
  NAND3_X1 U7016 ( .A1(n6082), .A2(n5967), .A3(n5966), .ZN(n5968) );
  OAI22_X1 U7017 ( .A1(n5969), .A2(n5968), .B1(n3851), .B2(n6537), .ZN(U3455)
         );
  INV_X1 U7018 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6455) );
  AOI21_X1 U7019 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6455), .A(n6463), .ZN(n5974) );
  INV_X1 U7020 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5970) );
  AND2_X1 U7021 ( .A1(n6463), .A2(STATE_REG_1__SCAN_IN), .ZN(n6548) );
  AOI21_X1 U7022 ( .B1(n5974), .B2(n5970), .A(n6548), .ZN(U2789) );
  OAI21_X1 U7023 ( .B1(n5971), .B2(n6443), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5972) );
  OAI21_X1 U7024 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6444), .A(n5972), .ZN(
        U2790) );
  INV_X2 U7025 ( .A(n6548), .ZN(n6560) );
  NOR2_X1 U7026 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5975) );
  OAI21_X1 U7027 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5975), .A(n6560), .ZN(n5973)
         );
  OAI21_X1 U7028 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6560), .A(n5973), .ZN(
        U2791) );
  NOR2_X1 U7029 ( .A1(n6548), .A2(n5974), .ZN(n6526) );
  OAI21_X1 U7030 ( .B1(BS16_N), .B2(n5975), .A(n6526), .ZN(n6524) );
  OAI21_X1 U7031 ( .B1(n6526), .B2(n6743), .A(n6524), .ZN(U2792) );
  INV_X1 U7032 ( .A(n5976), .ZN(n5978) );
  OAI21_X1 U7033 ( .B1(n5978), .B2(n5977), .A(n6181), .ZN(U2793) );
  NOR4_X1 U7034 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_20__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n5982) );
  NOR4_X1 U7035 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(
        DATAWIDTH_REG_15__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n5981) );
  NOR4_X1 U7036 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(
        DATAWIDTH_REG_29__SCAN_IN), .A3(DATAWIDTH_REG_30__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5980) );
  NOR4_X1 U7037 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(
        DATAWIDTH_REG_25__SCAN_IN), .A3(DATAWIDTH_REG_26__SCAN_IN), .A4(
        DATAWIDTH_REG_27__SCAN_IN), .ZN(n5979) );
  NAND4_X1 U7038 ( .A1(n5982), .A2(n5981), .A3(n5980), .A4(n5979), .ZN(n5988)
         );
  NOR4_X1 U7039 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), 
        .A3(DATAWIDTH_REG_4__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(
        n5986) );
  AOI211_X1 U7040 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_23__SCAN_IN), .B(
        DATAWIDTH_REG_21__SCAN_IN), .ZN(n5985) );
  NOR4_X1 U7041 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_12__SCAN_IN), .A4(
        DATAWIDTH_REG_13__SCAN_IN), .ZN(n5984) );
  NOR4_X1 U7042 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_7__SCAN_IN), 
        .A3(DATAWIDTH_REG_8__SCAN_IN), .A4(DATAWIDTH_REG_9__SCAN_IN), .ZN(
        n5983) );
  NAND4_X1 U7043 ( .A1(n5986), .A2(n5985), .A3(n5984), .A4(n5983), .ZN(n5987)
         );
  NOR2_X1 U7044 ( .A1(n5988), .A2(n5987), .ZN(n6547) );
  INV_X1 U7045 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5990) );
  NOR3_X1 U7046 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5991) );
  OAI21_X1 U7047 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5991), .A(n6547), .ZN(n5989)
         );
  OAI21_X1 U7048 ( .B1(n6547), .B2(n5990), .A(n5989), .ZN(U2794) );
  INV_X1 U7049 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6525) );
  AOI21_X1 U7050 ( .B1(n5331), .B2(n6525), .A(n5991), .ZN(n5993) );
  INV_X1 U7051 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5992) );
  INV_X1 U7052 ( .A(n6547), .ZN(n6542) );
  AOI22_X1 U7053 ( .A1(n6547), .A2(n5993), .B1(n5992), .B2(n6542), .ZN(U2795)
         );
  INV_X1 U7054 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6115) );
  INV_X1 U7055 ( .A(n5994), .ZN(n5996) );
  INV_X1 U7056 ( .A(REIP_REG_17__SCAN_IN), .ZN(n5995) );
  OAI21_X1 U7057 ( .B1(n6084), .B2(n5996), .A(n5995), .ZN(n5998) );
  AOI22_X1 U7058 ( .A1(n5998), .A2(n5997), .B1(PHYADDRPOINTER_REG_17__SCAN_IN), 
        .B2(n6097), .ZN(n5999) );
  OAI211_X1 U7059 ( .C1(n6065), .C2(n6115), .A(n6070), .B(n5999), .ZN(n6000)
         );
  INV_X1 U7060 ( .A(n6000), .ZN(n6002) );
  AOI22_X1 U7061 ( .A1(n6124), .A2(n6073), .B1(n6086), .B2(n6113), .ZN(n6001)
         );
  OAI211_X1 U7062 ( .C1(n6003), .C2(n6094), .A(n6002), .B(n6001), .ZN(U2810)
         );
  NOR3_X1 U7063 ( .A1(n6084), .A2(REIP_REG_16__SCAN_IN), .A3(n6004), .ZN(n6011) );
  INV_X1 U7064 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n6009) );
  INV_X1 U7065 ( .A(n6005), .ZN(n6007) );
  NOR3_X1 U7066 ( .A1(n6007), .A2(REIP_REG_15__SCAN_IN), .A3(n6006), .ZN(n6021) );
  OAI21_X1 U7067 ( .B1(n6021), .B2(n6017), .A(REIP_REG_16__SCAN_IN), .ZN(n6008) );
  OAI211_X1 U7068 ( .C1(n6078), .C2(n6009), .A(n6070), .B(n6008), .ZN(n6010)
         );
  AOI211_X1 U7069 ( .C1(n3003), .C2(EBX_REG_16__SCAN_IN), .A(n6011), .B(n6010), 
        .ZN(n6015) );
  INV_X1 U7070 ( .A(n6012), .ZN(n6013) );
  AOI22_X1 U7071 ( .A1(n6129), .A2(n6073), .B1(n6013), .B2(n6108), .ZN(n6014)
         );
  OAI211_X1 U7072 ( .C1(n6100), .C2(n6016), .A(n6015), .B(n6014), .ZN(U2811)
         );
  INV_X1 U7073 ( .A(n6561), .ZN(n6022) );
  AOI22_X1 U7074 ( .A1(EBX_REG_15__SCAN_IN), .A2(n3003), .B1(
        REIP_REG_15__SCAN_IN), .B2(n6017), .ZN(n6018) );
  OAI211_X1 U7075 ( .C1(n6078), .C2(n6019), .A(n6018), .B(n6070), .ZN(n6020)
         );
  AOI211_X1 U7076 ( .C1(n6022), .C2(n6073), .A(n6021), .B(n6020), .ZN(n6025)
         );
  AOI22_X1 U7077 ( .A1(n6023), .A2(n6108), .B1(n6086), .B2(n6564), .ZN(n6024)
         );
  NAND2_X1 U7078 ( .A1(n6025), .A2(n6024), .ZN(U2812) );
  INV_X1 U7079 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6486) );
  NOR3_X1 U7080 ( .A1(n6084), .A2(n6486), .A3(n6026), .ZN(n6035) );
  AOI21_X1 U7081 ( .B1(REIP_REG_10__SCAN_IN), .B2(n6035), .A(
        REIP_REG_11__SCAN_IN), .ZN(n6032) );
  AOI22_X1 U7082 ( .A1(EBX_REG_11__SCAN_IN), .A2(n3003), .B1(
        PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n6097), .ZN(n6027) );
  INV_X1 U7083 ( .A(n6027), .ZN(n6028) );
  AOI211_X1 U7084 ( .C1(n6086), .C2(n6116), .A(n6081), .B(n6028), .ZN(n6030)
         );
  INV_X1 U7085 ( .A(n6119), .ZN(n6178) );
  AOI22_X1 U7086 ( .A1(n6178), .A2(n6073), .B1(n6108), .B2(n6176), .ZN(n6029)
         );
  OAI211_X1 U7087 ( .C1(n6032), .C2(n6031), .A(n6030), .B(n6029), .ZN(U2816)
         );
  NAND2_X1 U7088 ( .A1(n6076), .A2(n6033), .ZN(n6063) );
  NAND3_X1 U7089 ( .A1(n6054), .A2(n6486), .A3(n6034), .ZN(n6050) );
  AOI22_X1 U7090 ( .A1(n6086), .A2(n6227), .B1(n6035), .B2(n5046), .ZN(n6036)
         );
  OAI211_X1 U7091 ( .C1(n6078), .C2(n6690), .A(n6036), .B(n6070), .ZN(n6041)
         );
  OAI22_X1 U7092 ( .A1(n6039), .A2(n6038), .B1(n6037), .B2(n6094), .ZN(n6040)
         );
  AOI211_X1 U7093 ( .C1(EBX_REG_10__SCAN_IN), .C2(n3003), .A(n6041), .B(n6040), 
        .ZN(n6042) );
  OAI221_X1 U7094 ( .B1(n5046), .B2(n6063), .C1(n5046), .C2(n6050), .A(n6042), 
        .ZN(U2817) );
  OAI22_X1 U7095 ( .A1(n6043), .A2(n6078), .B1(n6486), .B2(n6063), .ZN(n6044)
         );
  AOI211_X1 U7096 ( .C1(n3003), .C2(EBX_REG_9__SCAN_IN), .A(n6081), .B(n6044), 
        .ZN(n6052) );
  INV_X1 U7097 ( .A(n6045), .ZN(n6047) );
  AOI22_X1 U7098 ( .A1(n6047), .A2(n6073), .B1(n6108), .B2(n6046), .ZN(n6051)
         );
  INV_X1 U7099 ( .A(n6048), .ZN(n6236) );
  NAND2_X1 U7100 ( .A1(n6086), .A2(n6236), .ZN(n6049) );
  NAND4_X1 U7101 ( .A1(n6052), .A2(n6051), .A3(n6050), .A4(n6049), .ZN(U2818)
         );
  AOI21_X1 U7102 ( .B1(n6054), .B2(n6053), .A(REIP_REG_8__SCAN_IN), .ZN(n6064)
         );
  OAI22_X1 U7103 ( .A1(n6056), .A2(n6065), .B1(n6100), .B2(n6055), .ZN(n6057)
         );
  AOI211_X1 U7104 ( .C1(n6097), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n6081), 
        .B(n6057), .ZN(n6062) );
  INV_X1 U7105 ( .A(n6058), .ZN(n6059) );
  AOI22_X1 U7106 ( .A1(n6060), .A2(n6073), .B1(n6059), .B2(n6108), .ZN(n6061)
         );
  OAI211_X1 U7107 ( .C1(n6064), .C2(n6063), .A(n6062), .B(n6061), .ZN(U2819)
         );
  NOR2_X1 U7108 ( .A1(n6066), .A2(n6065), .ZN(n6067) );
  AOI211_X1 U7109 ( .C1(n6069), .C2(REIP_REG_6__SCAN_IN), .A(n6068), .B(n6067), 
        .ZN(n6075) );
  NAND2_X1 U7110 ( .A1(n6253), .A2(n6086), .ZN(n6071) );
  OAI211_X1 U7111 ( .C1(n3396), .C2(n6078), .A(n6071), .B(n6070), .ZN(n6072)
         );
  AOI21_X1 U7112 ( .B1(n6187), .B2(n6073), .A(n6072), .ZN(n6074) );
  OAI211_X1 U7113 ( .C1(n6190), .C2(n6094), .A(n6075), .B(n6074), .ZN(U2821)
         );
  INV_X1 U7114 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6079) );
  OAI21_X1 U7115 ( .B1(n6077), .B2(n6083), .A(n6076), .ZN(n6112) );
  OAI22_X1 U7116 ( .A1(n6079), .A2(n6078), .B1(n6477), .B2(n6112), .ZN(n6080)
         );
  AOI211_X1 U7117 ( .C1(n3003), .C2(EBX_REG_4__SCAN_IN), .A(n6081), .B(n6080), 
        .ZN(n6093) );
  INV_X1 U7118 ( .A(n6082), .ZN(n6089) );
  NOR3_X1 U7119 ( .A1(n6084), .A2(REIP_REG_4__SCAN_IN), .A3(n6083), .ZN(n6085)
         );
  AOI21_X1 U7120 ( .B1(n6259), .B2(n6086), .A(n6085), .ZN(n6087) );
  OAI21_X1 U7121 ( .B1(n6089), .B2(n6088), .A(n6087), .ZN(n6090) );
  AOI21_X1 U7122 ( .B1(n6195), .B2(n6091), .A(n6090), .ZN(n6092) );
  OAI211_X1 U7123 ( .C1(n6198), .C2(n6094), .A(n6093), .B(n6092), .ZN(U2823)
         );
  INV_X1 U7124 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6475) );
  INV_X1 U7125 ( .A(n6095), .ZN(n6096) );
  NAND2_X1 U7126 ( .A1(n6096), .A2(REIP_REG_2__SCAN_IN), .ZN(n6111) );
  AOI22_X1 U7127 ( .A1(n3003), .A2(EBX_REG_3__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n6097), .ZN(n6099) );
  OAI21_X1 U7128 ( .B1(n6100), .B2(n6266), .A(n6099), .ZN(n6101) );
  AOI21_X1 U7129 ( .B1(n6103), .B2(n6102), .A(n6101), .ZN(n6104) );
  OAI21_X1 U7130 ( .B1(n6106), .B2(n6105), .A(n6104), .ZN(n6107) );
  AOI21_X1 U7131 ( .B1(n6109), .B2(n6108), .A(n6107), .ZN(n6110) );
  OAI221_X1 U7132 ( .B1(n6112), .B2(n6475), .C1(n6112), .C2(n6111), .A(n6110), 
        .ZN(U2824) );
  AOI22_X1 U7133 ( .A1(n6124), .A2(n3906), .B1(n6563), .B2(n6113), .ZN(n6114)
         );
  OAI21_X1 U7134 ( .B1(n6123), .B2(n6115), .A(n6114), .ZN(U2842) );
  INV_X1 U7135 ( .A(EBX_REG_11__SCAN_IN), .ZN(n6122) );
  INV_X1 U7136 ( .A(n6116), .ZN(n6117) );
  OAI22_X1 U7137 ( .A1(n6119), .A2(n6118), .B1(n5546), .B2(n6117), .ZN(n6120)
         );
  INV_X1 U7138 ( .A(n6120), .ZN(n6121) );
  OAI21_X1 U7139 ( .B1(n6123), .B2(n6122), .A(n6121), .ZN(U2848) );
  AOI22_X1 U7140 ( .A1(n6124), .A2(n6128), .B1(n6127), .B2(DATAI_17_), .ZN(
        n6126) );
  AOI22_X1 U7141 ( .A1(n6131), .A2(DATAI_1_), .B1(n6130), .B2(
        EAX_REG_17__SCAN_IN), .ZN(n6125) );
  NAND2_X1 U7142 ( .A1(n6126), .A2(n6125), .ZN(U2874) );
  AOI22_X1 U7143 ( .A1(n6129), .A2(n6128), .B1(n6127), .B2(DATAI_16_), .ZN(
        n6133) );
  AOI22_X1 U7144 ( .A1(n6131), .A2(DATAI_0_), .B1(n6130), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n6132) );
  NAND2_X1 U7145 ( .A1(n6133), .A2(n6132), .ZN(U2875) );
  INV_X1 U7146 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n6705) );
  INV_X1 U7147 ( .A(n6134), .ZN(n6136) );
  AOI22_X1 U7148 ( .A1(n6136), .A2(EAX_REG_30__SCAN_IN), .B1(n6552), .B2(
        UWORD_REG_14__SCAN_IN), .ZN(n6135) );
  OAI21_X1 U7149 ( .B1(n6705), .B2(n6145), .A(n6135), .ZN(U2893) );
  INV_X1 U7150 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n6737) );
  AOI22_X1 U7151 ( .A1(n6136), .A2(EAX_REG_22__SCAN_IN), .B1(n6552), .B2(
        UWORD_REG_6__SCAN_IN), .ZN(n6137) );
  OAI21_X1 U7152 ( .B1(n6737), .B2(n6145), .A(n6137), .ZN(U2901) );
  AOI22_X1 U7153 ( .A1(n6552), .A2(LWORD_REG_15__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6138) );
  OAI21_X1 U7154 ( .B1(n6139), .B2(n6166), .A(n6138), .ZN(U2908) );
  INV_X1 U7155 ( .A(LWORD_REG_14__SCAN_IN), .ZN(n6736) );
  AOI22_X1 U7156 ( .A1(EAX_REG_14__SCAN_IN), .A2(n6162), .B1(n6163), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6140) );
  OAI21_X1 U7157 ( .B1(n6736), .B2(n6148), .A(n6140), .ZN(U2909) );
  AOI22_X1 U7158 ( .A1(n6552), .A2(LWORD_REG_13__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6141) );
  OAI21_X1 U7159 ( .B1(n6142), .B2(n6166), .A(n6141), .ZN(U2910) );
  AOI22_X1 U7160 ( .A1(n6552), .A2(LWORD_REG_12__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6143) );
  OAI21_X1 U7161 ( .B1(n5090), .B2(n6166), .A(n6143), .ZN(U2911) );
  INV_X1 U7162 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n6574) );
  AOI22_X1 U7163 ( .A1(EAX_REG_11__SCAN_IN), .A2(n6162), .B1(n6160), .B2(
        LWORD_REG_11__SCAN_IN), .ZN(n6144) );
  OAI21_X1 U7164 ( .B1(n6574), .B2(n6145), .A(n6144), .ZN(U2912) );
  AOI22_X1 U7165 ( .A1(EAX_REG_10__SCAN_IN), .A2(n6162), .B1(n6163), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6146) );
  OAI21_X1 U7166 ( .B1(n6591), .B2(n6148), .A(n6146), .ZN(U2913) );
  AOI22_X1 U7167 ( .A1(EAX_REG_9__SCAN_IN), .A2(n6162), .B1(n6163), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6147) );
  OAI21_X1 U7168 ( .B1(n6725), .B2(n6148), .A(n6147), .ZN(U2914) );
  AOI22_X1 U7169 ( .A1(n6552), .A2(LWORD_REG_8__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6149) );
  OAI21_X1 U7170 ( .B1(n6150), .B2(n6166), .A(n6149), .ZN(U2915) );
  INV_X1 U7171 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6152) );
  AOI22_X1 U7172 ( .A1(n6552), .A2(LWORD_REG_7__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6151) );
  OAI21_X1 U7173 ( .B1(n6152), .B2(n6166), .A(n6151), .ZN(U2916) );
  AOI22_X1 U7174 ( .A1(n6552), .A2(LWORD_REG_6__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6153) );
  OAI21_X1 U7175 ( .B1(n3397), .B2(n6166), .A(n6153), .ZN(U2917) );
  AOI22_X1 U7176 ( .A1(n6552), .A2(LWORD_REG_5__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6154) );
  OAI21_X1 U7177 ( .B1(n6155), .B2(n6166), .A(n6154), .ZN(U2918) );
  AOI22_X1 U7178 ( .A1(n6552), .A2(LWORD_REG_4__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6156) );
  OAI21_X1 U7179 ( .B1(n6157), .B2(n6166), .A(n6156), .ZN(U2919) );
  AOI22_X1 U7180 ( .A1(n6552), .A2(LWORD_REG_3__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6158) );
  OAI21_X1 U7181 ( .B1(n6159), .B2(n6166), .A(n6158), .ZN(U2920) );
  AOI222_X1 U7182 ( .A1(n6163), .A2(DATAO_REG_2__SCAN_IN), .B1(n6162), .B2(
        EAX_REG_2__SCAN_IN), .C1(n6160), .C2(LWORD_REG_2__SCAN_IN), .ZN(n6161)
         );
  INV_X1 U7183 ( .A(n6161), .ZN(U2921) );
  AOI222_X1 U7184 ( .A1(n6163), .A2(DATAO_REG_1__SCAN_IN), .B1(n6162), .B2(
        EAX_REG_1__SCAN_IN), .C1(n6552), .C2(LWORD_REG_1__SCAN_IN), .ZN(n6164)
         );
  INV_X1 U7185 ( .A(n6164), .ZN(U2922) );
  AOI22_X1 U7186 ( .A1(n6552), .A2(LWORD_REG_0__SCAN_IN), .B1(n6163), .B2(
        DATAO_REG_0__SCAN_IN), .ZN(n6165) );
  OAI21_X1 U7187 ( .B1(n6167), .B2(n6166), .A(n6165), .ZN(U2923) );
  AOI22_X1 U7188 ( .A1(n6173), .A2(EAX_REG_30__SCAN_IN), .B1(
        UWORD_REG_14__SCAN_IN), .B2(n6172), .ZN(n6169) );
  NAND2_X1 U7189 ( .A1(n6168), .A2(DATAI_14_), .ZN(n6174) );
  NAND2_X1 U7190 ( .A1(n6169), .A2(n6174), .ZN(U2938) );
  AOI22_X1 U7191 ( .A1(n6173), .A2(EAX_REG_11__SCAN_IN), .B1(
        LWORD_REG_11__SCAN_IN), .B2(n6172), .ZN(n6171) );
  NAND2_X1 U7192 ( .A1(n6171), .A2(n6170), .ZN(U2950) );
  AOI22_X1 U7193 ( .A1(n6173), .A2(EAX_REG_14__SCAN_IN), .B1(
        LWORD_REG_14__SCAN_IN), .B2(n6172), .ZN(n6175) );
  NAND2_X1 U7194 ( .A1(n6175), .A2(n6174), .ZN(U2953) );
  AOI22_X1 U7195 ( .A1(n6277), .A2(REIP_REG_11__SCAN_IN), .B1(n6199), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n6180) );
  AOI22_X1 U7196 ( .A1(n6178), .A2(n6205), .B1(n6177), .B2(n6176), .ZN(n6179)
         );
  OAI211_X1 U7197 ( .C1(n6182), .C2(n6181), .A(n6180), .B(n6179), .ZN(U2975)
         );
  AOI22_X1 U7198 ( .A1(n6277), .A2(REIP_REG_6__SCAN_IN), .B1(n6199), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n6189) );
  OAI21_X1 U7199 ( .B1(n3005), .B2(n6184), .A(n6183), .ZN(n6186) );
  INV_X1 U7200 ( .A(n6186), .ZN(n6252) );
  AOI22_X1 U7201 ( .A1(n6252), .A2(n6204), .B1(n6205), .B2(n6187), .ZN(n6188)
         );
  OAI211_X1 U7202 ( .C1(n6210), .C2(n6190), .A(n6189), .B(n6188), .ZN(U2980)
         );
  AOI22_X1 U7203 ( .A1(n6277), .A2(REIP_REG_4__SCAN_IN), .B1(n6199), .B2(
        PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6197) );
  OAI21_X1 U7204 ( .B1(n6193), .B2(n6192), .A(n6191), .ZN(n6194) );
  INV_X1 U7205 ( .A(n6194), .ZN(n6258) );
  AOI22_X1 U7206 ( .A1(n6258), .A2(n6204), .B1(n6205), .B2(n6195), .ZN(n6196)
         );
  OAI211_X1 U7207 ( .C1(n6210), .C2(n6198), .A(n6197), .B(n6196), .ZN(U2982)
         );
  AOI22_X1 U7208 ( .A1(n6277), .A2(REIP_REG_2__SCAN_IN), .B1(n6199), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6208) );
  CLKBUF_X1 U7209 ( .A(n6200), .Z(n6201) );
  XNOR2_X1 U7210 ( .A(n6201), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6203)
         );
  XNOR2_X1 U7211 ( .A(n6203), .B(n6202), .ZN(n6283) );
  AOI22_X1 U7212 ( .A1(n6206), .A2(n6205), .B1(n6283), .B2(n6204), .ZN(n6207)
         );
  OAI211_X1 U7213 ( .C1(n6210), .C2(n6209), .A(n6208), .B(n6207), .ZN(U2984)
         );
  NAND2_X1 U7214 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n6211), .ZN(n6224) );
  AOI21_X1 U7215 ( .B1(n6213), .B2(n6212), .A(INSTADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n6215) );
  NOR2_X1 U7216 ( .A1(n6215), .A2(n6214), .ZN(n6222) );
  OAI22_X1 U7217 ( .A1(n6218), .A2(n6217), .B1(n6491), .B2(n6216), .ZN(n6219)
         );
  AOI21_X1 U7218 ( .B1(n6220), .B2(n6284), .A(n6219), .ZN(n6221) );
  OAI221_X1 U7219 ( .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n6224), .C1(
        n6223), .C2(n6222), .A(n6221), .ZN(U3006) );
  NAND2_X1 U7220 ( .A1(n6229), .A2(n6247), .ZN(n6241) );
  AOI22_X1 U7221 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n6225), .B1(
        INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n5099), .ZN(n6233) );
  AOI21_X1 U7222 ( .B1(n6227), .B2(n6279), .A(n6226), .ZN(n6232) );
  OAI21_X1 U7223 ( .B1(n6229), .B2(n6228), .A(n6251), .ZN(n6237) );
  AOI22_X1 U7224 ( .A1(n6230), .A2(n6284), .B1(INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n6237), .ZN(n6231) );
  OAI211_X1 U7225 ( .C1(n6241), .C2(n6233), .A(n6232), .B(n6231), .ZN(U3008)
         );
  INV_X1 U7226 ( .A(n6234), .ZN(n6235) );
  AOI21_X1 U7227 ( .B1(n6236), .B2(n6279), .A(n6235), .ZN(n6240) );
  AOI22_X1 U7228 ( .A1(n6238), .A2(n6284), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n6237), .ZN(n6239) );
  OAI211_X1 U7229 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n6241), .A(n6240), 
        .B(n6239), .ZN(U3009) );
  INV_X1 U7230 ( .A(n6242), .ZN(n6243) );
  AOI21_X1 U7231 ( .B1(n6244), .B2(n6279), .A(n6243), .ZN(n6249) );
  INV_X1 U7232 ( .A(n6245), .ZN(n6246) );
  AOI22_X1 U7233 ( .A1(n6247), .A2(n6250), .B1(n6246), .B2(n6284), .ZN(n6248)
         );
  OAI211_X1 U7234 ( .C1(n6251), .C2(n6250), .A(n6249), .B(n6248), .ZN(U3011)
         );
  AOI222_X1 U7235 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6260), .B1(n6279), .B2(
        n6253), .C1(n6284), .C2(n6252), .ZN(n6254) );
  OAI221_X1 U7236 ( .B1(INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n6257), .C1(n6256), .C2(n6255), .A(n6254), .ZN(U3012) );
  AOI21_X1 U7237 ( .B1(n6280), .B2(n6282), .A(n6285), .ZN(n6275) );
  AOI222_X1 U7238 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6260), .B1(n6279), .B2(
        n6259), .C1(n6284), .C2(n6258), .ZN(n6264) );
  NOR2_X1 U7239 ( .A1(n6282), .A2(n6261), .ZN(n6271) );
  OAI211_X1 U7240 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n6271), .B(n6262), .ZN(n6263) );
  OAI211_X1 U7241 ( .C1(n6275), .C2(n6265), .A(n6264), .B(n6263), .ZN(U3014)
         );
  INV_X1 U7242 ( .A(n6266), .ZN(n6268) );
  AOI21_X1 U7243 ( .B1(n6279), .B2(n6268), .A(n6267), .ZN(n6273) );
  INV_X1 U7244 ( .A(n6269), .ZN(n6270) );
  AOI22_X1 U7245 ( .A1(n6271), .A2(n6274), .B1(n6270), .B2(n6284), .ZN(n6272)
         );
  OAI211_X1 U7246 ( .C1(n6275), .C2(n6274), .A(n6273), .B(n6272), .ZN(U3015)
         );
  INV_X1 U7247 ( .A(n6276), .ZN(n6278) );
  AOI22_X1 U7248 ( .A1(n6279), .A2(n6278), .B1(n6277), .B2(REIP_REG_2__SCAN_IN), .ZN(n6291) );
  OAI221_X1 U7249 ( .B1(n6282), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .C1(n6282), .C2(n6281), .A(n6280), .ZN(n6290) );
  AOI22_X1 U7250 ( .A1(n6285), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6284), 
        .B2(n6283), .ZN(n6289) );
  NAND3_X1 U7251 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6287), .A3(n6286), 
        .ZN(n6288) );
  NAND4_X1 U7252 ( .A1(n6291), .A2(n6290), .A3(n6289), .A4(n6288), .ZN(U3016)
         );
  NOR2_X1 U7253 ( .A1(n6293), .A2(n6292), .ZN(U3019) );
  AOI22_X1 U7254 ( .A1(n6375), .A2(n6299), .B1(n6374), .B2(n6298), .ZN(n6295)
         );
  AOI22_X1 U7255 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6301), .B1(n6376), 
        .B2(n6300), .ZN(n6294) );
  OAI211_X1 U7256 ( .C1(n6304), .C2(n6379), .A(n6295), .B(n6294), .ZN(U3045)
         );
  AOI22_X1 U7257 ( .A1(n6381), .A2(n6299), .B1(n6380), .B2(n6298), .ZN(n6297)
         );
  AOI22_X1 U7258 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6301), .B1(n6382), 
        .B2(n6300), .ZN(n6296) );
  OAI211_X1 U7259 ( .C1(n6304), .C2(n6385), .A(n6297), .B(n6296), .ZN(U3047)
         );
  AOI22_X1 U7260 ( .A1(n6389), .A2(n6299), .B1(n6387), .B2(n6298), .ZN(n6303)
         );
  AOI22_X1 U7261 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6301), .B1(n6391), 
        .B2(n6300), .ZN(n6302) );
  OAI211_X1 U7262 ( .C1(n6304), .C2(n6396), .A(n6303), .B(n6302), .ZN(U3050)
         );
  NAND3_X1 U7263 ( .A1(n6306), .A2(n6305), .A3(n6718), .ZN(n6307) );
  OAI21_X1 U7264 ( .B1(n6309), .B2(n6308), .A(n6307), .ZN(n6357) );
  NAND2_X1 U7265 ( .A1(n6406), .A2(n6310), .ZN(n6317) );
  INV_X1 U7266 ( .A(n6317), .ZN(n6355) );
  AOI22_X1 U7267 ( .A1(n6312), .A2(n6357), .B1(n6311), .B2(n6355), .ZN(n6323)
         );
  AOI21_X1 U7268 ( .B1(n6313), .B2(n6373), .A(n6743), .ZN(n6320) );
  NAND2_X1 U7269 ( .A1(n6314), .A2(n4551), .ZN(n6319) );
  AOI211_X1 U7270 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6317), .A(n6316), .B(
        n6315), .ZN(n6318) );
  OAI211_X1 U7271 ( .C1(n6320), .C2(n6319), .A(n6318), .B(n6718), .ZN(n6361)
         );
  AOI22_X1 U7272 ( .A1(n6361), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6321), 
        .B2(n6359), .ZN(n6322) );
  OAI211_X1 U7273 ( .C1(n6324), .C2(n6373), .A(n6323), .B(n6322), .ZN(U3068)
         );
  AOI22_X1 U7274 ( .A1(n6376), .A2(n6357), .B1(n6375), .B2(n6355), .ZN(n6327)
         );
  AOI22_X1 U7275 ( .A1(n6361), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6325), 
        .B2(n6359), .ZN(n6326) );
  OAI211_X1 U7276 ( .C1(n6328), .C2(n6373), .A(n6327), .B(n6326), .ZN(U3069)
         );
  AOI22_X1 U7277 ( .A1(n6330), .A2(n6357), .B1(n6329), .B2(n6355), .ZN(n6333)
         );
  AOI22_X1 U7278 ( .A1(n6361), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6331), 
        .B2(n6359), .ZN(n6332) );
  OAI211_X1 U7279 ( .C1(n6334), .C2(n6373), .A(n6333), .B(n6332), .ZN(U3070)
         );
  AOI22_X1 U7280 ( .A1(n6382), .A2(n6357), .B1(n6381), .B2(n6355), .ZN(n6337)
         );
  AOI22_X1 U7281 ( .A1(n6361), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6335), 
        .B2(n6359), .ZN(n6336) );
  OAI211_X1 U7282 ( .C1(n6338), .C2(n6373), .A(n6337), .B(n6336), .ZN(U3071)
         );
  AOI22_X1 U7283 ( .A1(n6340), .A2(n6357), .B1(n6339), .B2(n6355), .ZN(n6343)
         );
  AOI22_X1 U7284 ( .A1(n6361), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6341), 
        .B2(n6359), .ZN(n6342) );
  OAI211_X1 U7285 ( .C1(n6344), .C2(n6373), .A(n6343), .B(n6342), .ZN(U3072)
         );
  AOI22_X1 U7286 ( .A1(n6346), .A2(n6357), .B1(n6345), .B2(n6355), .ZN(n6349)
         );
  AOI22_X1 U7287 ( .A1(n6361), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6347), 
        .B2(n6359), .ZN(n6348) );
  OAI211_X1 U7288 ( .C1(n6350), .C2(n6373), .A(n6349), .B(n6348), .ZN(U3073)
         );
  AOI22_X1 U7289 ( .A1(n6391), .A2(n6357), .B1(n6389), .B2(n6355), .ZN(n6353)
         );
  AOI22_X1 U7290 ( .A1(n6361), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6351), 
        .B2(n6359), .ZN(n6352) );
  OAI211_X1 U7291 ( .C1(n6354), .C2(n6373), .A(n6353), .B(n6352), .ZN(U3074)
         );
  AOI22_X1 U7292 ( .A1(n6358), .A2(n6357), .B1(n6356), .B2(n6355), .ZN(n6363)
         );
  AOI22_X1 U7293 ( .A1(n6361), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6360), 
        .B2(n6359), .ZN(n6362) );
  OAI211_X1 U7294 ( .C1(n6364), .C2(n6373), .A(n6363), .B(n6362), .ZN(U3075)
         );
  INV_X1 U7295 ( .A(n6365), .ZN(n6368) );
  INV_X1 U7296 ( .A(n6366), .ZN(n6367) );
  AOI22_X1 U7297 ( .A1(n6375), .A2(n6368), .B1(n6374), .B2(n6367), .ZN(n6372)
         );
  AOI22_X1 U7298 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6370), .B1(n6376), 
        .B2(n6369), .ZN(n6371) );
  OAI211_X1 U7299 ( .C1(n6379), .C2(n6373), .A(n6372), .B(n6371), .ZN(U3077)
         );
  AOI22_X1 U7300 ( .A1(n6375), .A2(n6388), .B1(n6374), .B2(n6386), .ZN(n6378)
         );
  AOI22_X1 U7301 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6392), .B1(n6376), 
        .B2(n6390), .ZN(n6377) );
  OAI211_X1 U7302 ( .C1(n6379), .C2(n6395), .A(n6378), .B(n6377), .ZN(U3109)
         );
  AOI22_X1 U7303 ( .A1(n6381), .A2(n6388), .B1(n6380), .B2(n6386), .ZN(n6384)
         );
  AOI22_X1 U7304 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6392), .B1(n6382), 
        .B2(n6390), .ZN(n6383) );
  OAI211_X1 U7305 ( .C1(n6385), .C2(n6395), .A(n6384), .B(n6383), .ZN(U3111)
         );
  AOI22_X1 U7306 ( .A1(n6389), .A2(n6388), .B1(n6387), .B2(n6386), .ZN(n6394)
         );
  AOI22_X1 U7307 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6392), .B1(n6391), 
        .B2(n6390), .ZN(n6393) );
  OAI211_X1 U7308 ( .C1(n6396), .C2(n6395), .A(n6394), .B(n6393), .ZN(U3114)
         );
  AND2_X1 U7309 ( .A1(n6398), .A2(n6397), .ZN(n6417) );
  INV_X1 U7310 ( .A(n6398), .ZN(n6410) );
  NAND2_X1 U7311 ( .A1(n6398), .A2(n6399), .ZN(n6415) );
  INV_X1 U7312 ( .A(n6400), .ZN(n6403) );
  INV_X1 U7313 ( .A(n6401), .ZN(n6402) );
  OAI22_X1 U7314 ( .A1(n6404), .A2(n6403), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6402), .ZN(n6531) );
  NAND2_X1 U7315 ( .A1(n6405), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6540) );
  INV_X1 U7316 ( .A(n6540), .ZN(n6407) );
  NOR3_X1 U7317 ( .A1(n6531), .A2(n6407), .A3(n6406), .ZN(n6411) );
  NAND2_X1 U7318 ( .A1(n6411), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6413) );
  INV_X1 U7319 ( .A(n6408), .ZN(n6409) );
  OAI22_X1 U7320 ( .A1(n6411), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n6410), .B2(n6409), .ZN(n6412) );
  NAND2_X1 U7321 ( .A1(n6413), .A2(n6412), .ZN(n6414) );
  AOI222_X1 U7322 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6415), .B1(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6414), .C1(n6415), .C2(n6414), 
        .ZN(n6416) );
  AOI222_X1 U7323 ( .A1(n6417), .A2(n6416), .B1(n6417), .B2(n6718), .C1(n6416), 
        .C2(n6718), .ZN(n6420) );
  OAI21_X1 U7324 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6418), 
        .ZN(n6419) );
  OAI21_X1 U7325 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n6420), .A(n6419), 
        .ZN(n6426) );
  INV_X1 U7326 ( .A(n6421), .ZN(n6422) );
  NAND3_X1 U7327 ( .A1(n6424), .A2(n6423), .A3(n6422), .ZN(n6425) );
  NOR2_X1 U7328 ( .A1(n6426), .A2(n6425), .ZN(n6442) );
  NOR2_X1 U7329 ( .A1(n6428), .A2(n6427), .ZN(n6432) );
  AOI22_X1 U7330 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), 
        .B1(READY_N), .B2(n6429), .ZN(n6430) );
  AOI21_X1 U7331 ( .B1(n6432), .B2(n6431), .A(n6430), .ZN(n6437) );
  NAND2_X1 U7332 ( .A1(n6437), .A2(n6442), .ZN(n6529) );
  NAND2_X1 U7333 ( .A1(READY_N), .A2(n6433), .ZN(n6450) );
  NAND3_X1 U7334 ( .A1(n6434), .A2(n6529), .A3(n6450), .ZN(n6436) );
  AOI21_X1 U7335 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6436), .A(n6435), .ZN(
        n6441) );
  NOR2_X1 U7336 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6437), .ZN(n6445) );
  OAI21_X1 U7337 ( .B1(n6439), .B2(n6438), .A(n6445), .ZN(n6440) );
  OAI211_X1 U7338 ( .C1(n6442), .C2(n6443), .A(n6441), .B(n6440), .ZN(U3148)
         );
  OAI21_X1 U7339 ( .B1(READY_N), .B2(n6444), .A(n6443), .ZN(n6448) );
  AOI211_X1 U7340 ( .C1(STATE2_REG_0__SCAN_IN), .C2(n6450), .A(n6445), .B(
        n6532), .ZN(n6446) );
  AOI211_X1 U7341 ( .C1(n6529), .C2(n6448), .A(n6447), .B(n6446), .ZN(n6449)
         );
  INV_X1 U7342 ( .A(n6449), .ZN(U3149) );
  INV_X1 U7343 ( .A(n6527), .ZN(n6453) );
  OAI221_X1 U7344 ( .B1(STATE2_REG_2__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(STATE2_REG_2__SCAN_IN), .C2(STATE2_REG_1__SCAN_IN), .A(n6450), 
        .ZN(n6452) );
  OAI21_X1 U7345 ( .B1(n6453), .B2(n6452), .A(n6451), .ZN(U3150) );
  INV_X1 U7346 ( .A(n6526), .ZN(n6454) );
  AND2_X1 U7347 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6454), .ZN(U3151) );
  AND2_X1 U7348 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6454), .ZN(U3152) );
  AND2_X1 U7349 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6454), .ZN(U3153) );
  AND2_X1 U7350 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6454), .ZN(U3154) );
  AND2_X1 U7351 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6454), .ZN(U3155) );
  AND2_X1 U7352 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6454), .ZN(U3156) );
  AND2_X1 U7353 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6454), .ZN(U3157) );
  AND2_X1 U7354 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6454), .ZN(U3158) );
  INV_X1 U7355 ( .A(DATAWIDTH_REG_23__SCAN_IN), .ZN(n6607) );
  NOR2_X1 U7356 ( .A1(n6526), .A2(n6607), .ZN(U3159) );
  AND2_X1 U7357 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6454), .ZN(U3160) );
  INV_X1 U7358 ( .A(DATAWIDTH_REG_21__SCAN_IN), .ZN(n6589) );
  NOR2_X1 U7359 ( .A1(n6526), .A2(n6589), .ZN(U3161) );
  AND2_X1 U7360 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(n6454), .ZN(U3162) );
  AND2_X1 U7361 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6454), .ZN(U3163) );
  AND2_X1 U7362 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6454), .ZN(U3164) );
  AND2_X1 U7363 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6454), .ZN(U3165) );
  AND2_X1 U7364 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6454), .ZN(U3166) );
  AND2_X1 U7365 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6454), .ZN(U3167) );
  AND2_X1 U7366 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6454), .ZN(U3168) );
  AND2_X1 U7367 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6454), .ZN(U3169) );
  AND2_X1 U7368 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6454), .ZN(U3170) );
  AND2_X1 U7369 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6454), .ZN(U3171) );
  AND2_X1 U7370 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6454), .ZN(U3172) );
  AND2_X1 U7371 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6454), .ZN(U3173) );
  AND2_X1 U7372 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6454), .ZN(U3174) );
  AND2_X1 U7373 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6454), .ZN(U3175) );
  AND2_X1 U7374 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6454), .ZN(U3176) );
  AND2_X1 U7375 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6454), .ZN(U3177) );
  AND2_X1 U7376 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6454), .ZN(U3178) );
  AND2_X1 U7377 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6454), .ZN(U3179) );
  AND2_X1 U7378 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6454), .ZN(U3180) );
  NOR2_X1 U7379 ( .A1(n6462), .A2(n6455), .ZN(n6465) );
  AOI22_X1 U7380 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6469) );
  AND2_X1 U7381 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6459) );
  INV_X1 U7382 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6457) );
  INV_X1 U7383 ( .A(NA_N), .ZN(n6466) );
  AOI211_X1 U7384 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6466), .A(
        STATE_REG_0__SCAN_IN), .B(n6465), .ZN(n6471) );
  AOI221_X1 U7385 ( .B1(n6459), .B2(n6560), .C1(n6457), .C2(n6560), .A(n6471), 
        .ZN(n6456) );
  OAI21_X1 U7386 ( .B1(n6465), .B2(n6469), .A(n6456), .ZN(U3181) );
  NOR2_X1 U7387 ( .A1(n6463), .A2(n6457), .ZN(n6467) );
  NAND2_X1 U7388 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6458) );
  OAI21_X1 U7389 ( .B1(n6467), .B2(n6459), .A(n6458), .ZN(n6460) );
  OAI211_X1 U7390 ( .C1(n6462), .C2(n6551), .A(n6461), .B(n6460), .ZN(U3182)
         );
  AOI221_X1 U7391 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6551), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6464) );
  AOI221_X1 U7392 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6464), .C2(HOLD), .A(n6463), .ZN(n6470) );
  AOI21_X1 U7393 ( .B1(n6467), .B2(n6466), .A(n6465), .ZN(n6468) );
  OAI22_X1 U7394 ( .A1(n6471), .A2(n6470), .B1(n6469), .B2(n6468), .ZN(U3183)
         );
  INV_X1 U7395 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6473) );
  INV_X1 U7396 ( .A(n6514), .ZN(n6522) );
  NAND2_X1 U7397 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6548), .ZN(n6516) );
  INV_X1 U7398 ( .A(n6516), .ZN(n6520) );
  AOI22_X1 U7399 ( .A1(REIP_REG_1__SCAN_IN), .A2(n6520), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6560), .ZN(n6472) );
  OAI21_X1 U7400 ( .B1(n6473), .B2(n6522), .A(n6472), .ZN(U3184) );
  AOI22_X1 U7401 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6520), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6560), .ZN(n6474) );
  OAI21_X1 U7402 ( .B1(n6475), .B2(n6522), .A(n6474), .ZN(U3185) );
  AOI22_X1 U7403 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6520), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6560), .ZN(n6476) );
  OAI21_X1 U7404 ( .B1(n6477), .B2(n6522), .A(n6476), .ZN(U3186) );
  AOI22_X1 U7405 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6520), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6560), .ZN(n6478) );
  OAI21_X1 U7406 ( .B1(n6479), .B2(n6522), .A(n6478), .ZN(U3187) );
  AOI22_X1 U7407 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6520), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6560), .ZN(n6480) );
  OAI21_X1 U7408 ( .B1(n6481), .B2(n6522), .A(n6480), .ZN(U3188) );
  AOI22_X1 U7409 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6520), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6560), .ZN(n6482) );
  OAI21_X1 U7410 ( .B1(n6484), .B2(n6522), .A(n6482), .ZN(U3189) );
  AOI22_X1 U7411 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6514), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6560), .ZN(n6483) );
  OAI21_X1 U7412 ( .B1(n6484), .B2(n6516), .A(n6483), .ZN(U3190) );
  AOI22_X1 U7413 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6520), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6560), .ZN(n6485) );
  OAI21_X1 U7414 ( .B1(n6486), .B2(n6522), .A(n6485), .ZN(U3191) );
  AOI22_X1 U7415 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6520), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6560), .ZN(n6487) );
  OAI21_X1 U7416 ( .B1(n5046), .B2(n6522), .A(n6487), .ZN(U3192) );
  AOI22_X1 U7417 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6514), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6560), .ZN(n6488) );
  OAI21_X1 U7418 ( .B1(n5046), .B2(n6516), .A(n6488), .ZN(U3193) );
  AOI22_X1 U7419 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6520), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6560), .ZN(n6489) );
  OAI21_X1 U7420 ( .B1(n6491), .B2(n6522), .A(n6489), .ZN(U3194) );
  AOI22_X1 U7421 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6514), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6560), .ZN(n6490) );
  OAI21_X1 U7422 ( .B1(n6491), .B2(n6516), .A(n6490), .ZN(U3195) );
  AOI22_X1 U7423 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6514), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6560), .ZN(n6492) );
  OAI21_X1 U7424 ( .B1(n6493), .B2(n6516), .A(n6492), .ZN(U3196) );
  AOI22_X1 U7425 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6514), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6560), .ZN(n6494) );
  OAI21_X1 U7426 ( .B1(n6605), .B2(n6516), .A(n6494), .ZN(U3197) );
  AOI22_X1 U7427 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6520), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6560), .ZN(n6495) );
  OAI21_X1 U7428 ( .B1(n6497), .B2(n6522), .A(n6495), .ZN(U3198) );
  AOI22_X1 U7429 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6514), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6560), .ZN(n6496) );
  OAI21_X1 U7430 ( .B1(n6497), .B2(n6516), .A(n6496), .ZN(U3199) );
  AOI22_X1 U7431 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6520), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6560), .ZN(n6498) );
  OAI21_X1 U7432 ( .B1(n6500), .B2(n6522), .A(n6498), .ZN(U3200) );
  AOI22_X1 U7433 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6514), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6560), .ZN(n6499) );
  OAI21_X1 U7434 ( .B1(n6500), .B2(n6516), .A(n6499), .ZN(U3201) );
  AOI22_X1 U7435 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6520), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6560), .ZN(n6501) );
  OAI21_X1 U7436 ( .B1(n6503), .B2(n6522), .A(n6501), .ZN(U3202) );
  AOI22_X1 U7437 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6514), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6560), .ZN(n6502) );
  OAI21_X1 U7438 ( .B1(n6503), .B2(n6516), .A(n6502), .ZN(U3203) );
  AOI22_X1 U7439 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6514), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6560), .ZN(n6504) );
  OAI21_X1 U7440 ( .B1(n5627), .B2(n6516), .A(n6504), .ZN(U3204) );
  AOI22_X1 U7441 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6520), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6560), .ZN(n6505) );
  OAI21_X1 U7442 ( .B1(n6506), .B2(n6522), .A(n6505), .ZN(U3205) );
  INV_X1 U7443 ( .A(ADDRESS_REG_22__SCAN_IN), .ZN(n6689) );
  OAI222_X1 U7444 ( .A1(n6516), .A2(n6506), .B1(n6689), .B2(n6548), .C1(n6508), 
        .C2(n6522), .ZN(U3206) );
  AOI22_X1 U7445 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6514), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6560), .ZN(n6507) );
  OAI21_X1 U7446 ( .B1(n6508), .B2(n6516), .A(n6507), .ZN(U3207) );
  AOI22_X1 U7447 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6514), .B1(
        ADDRESS_REG_24__SCAN_IN), .B2(n6560), .ZN(n6509) );
  OAI21_X1 U7448 ( .B1(n6510), .B2(n6516), .A(n6509), .ZN(U3208) );
  AOI22_X1 U7449 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6514), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6560), .ZN(n6511) );
  OAI21_X1 U7450 ( .B1(n6512), .B2(n6516), .A(n6511), .ZN(U3209) );
  INV_X1 U7451 ( .A(ADDRESS_REG_26__SCAN_IN), .ZN(n6722) );
  INV_X1 U7452 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6517) );
  OAI222_X1 U7453 ( .A1(n6516), .A2(n6513), .B1(n6722), .B2(n6548), .C1(n6517), 
        .C2(n6522), .ZN(U3210) );
  AOI22_X1 U7454 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6514), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6560), .ZN(n6515) );
  OAI21_X1 U7455 ( .B1(n6517), .B2(n6516), .A(n6515), .ZN(U3211) );
  AOI22_X1 U7456 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6520), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6560), .ZN(n6518) );
  OAI21_X1 U7457 ( .B1(n6519), .B2(n6522), .A(n6518), .ZN(U3212) );
  AOI22_X1 U7458 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6520), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6560), .ZN(n6521) );
  OAI21_X1 U7459 ( .B1(n5480), .B2(n6522), .A(n6521), .ZN(U3213) );
  MUX2_X1 U7460 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6560), .Z(U3445) );
  MUX2_X1 U7461 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6560), .Z(U3446) );
  MUX2_X1 U7462 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6560), .Z(U3447) );
  MUX2_X1 U7463 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6560), .Z(U3448) );
  OAI21_X1 U7464 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6526), .A(n6524), .ZN(
        n6523) );
  INV_X1 U7465 ( .A(n6523), .ZN(U3451) );
  OAI21_X1 U7466 ( .B1(n6526), .B2(n6525), .A(n6524), .ZN(U3452) );
  OAI211_X1 U7467 ( .C1(n3149), .C2(n6529), .A(n6528), .B(n6527), .ZN(U3453)
         );
  INV_X1 U7468 ( .A(n6530), .ZN(n6535) );
  NAND2_X1 U7469 ( .A1(n6531), .A2(n3149), .ZN(n6533) );
  MUX2_X1 U7470 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .B(n6533), .S(n6532), 
        .Z(n6534) );
  NAND3_X1 U7471 ( .A1(n6537), .A2(n6535), .A3(n6534), .ZN(n6536) );
  OAI21_X1 U7472 ( .B1(n6537), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n6536), 
        .ZN(n6538) );
  OAI21_X1 U7473 ( .B1(n6540), .B2(n6539), .A(n6538), .ZN(U3461) );
  AOI21_X1 U7474 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6541) );
  AOI22_X1 U7475 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6541), .B2(n5331), .ZN(n6544) );
  INV_X1 U7476 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6543) );
  AOI22_X1 U7477 ( .A1(n6547), .A2(n6544), .B1(n6543), .B2(n6542), .ZN(U3468)
         );
  INV_X1 U7478 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6546) );
  OAI21_X1 U7479 ( .B1(REIP_REG_1__SCAN_IN), .B2(REIP_REG_0__SCAN_IN), .A(
        n6547), .ZN(n6545) );
  OAI21_X1 U7480 ( .B1(n6547), .B2(n6546), .A(n6545), .ZN(U3469) );
  INV_X1 U7481 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6692) );
  AOI22_X1 U7482 ( .A1(n6548), .A2(READREQUEST_REG_SCAN_IN), .B1(n6692), .B2(
        n6560), .ZN(U3470) );
  AOI211_X1 U7483 ( .C1(n6552), .C2(n6551), .A(n6550), .B(n6549), .ZN(n6559)
         );
  OAI211_X1 U7484 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6554), .A(n6553), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6556) );
  AOI21_X1 U7485 ( .B1(n6556), .B2(STATE2_REG_0__SCAN_IN), .A(n6555), .ZN(
        n6558) );
  NAND2_X1 U7486 ( .A1(n6559), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6557) );
  OAI21_X1 U7487 ( .B1(n6559), .B2(n6558), .A(n6557), .ZN(U3472) );
  MUX2_X1 U7488 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6560), .Z(U3473) );
  OR2_X1 U7489 ( .A1(n6561), .A2(n6118), .ZN(n6566) );
  AOI22_X1 U7490 ( .A1(n6564), .A2(n6563), .B1(EBX_REG_15__SCAN_IN), .B2(n6562), .ZN(n6565) );
  INV_X1 U7491 ( .A(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n6739) );
  AOI22_X1 U7492 ( .A1(n6739), .A2(keyinput100), .B1(keyinput72), .B2(n6718), 
        .ZN(n6567) );
  OAI221_X1 U7493 ( .B1(n6739), .B2(keyinput100), .C1(n6718), .C2(keyinput72), 
        .A(n6567), .ZN(n6578) );
  AOI22_X1 U7494 ( .A1(n4492), .A2(keyinput115), .B1(keyinput105), .B2(n6569), 
        .ZN(n6568) );
  OAI221_X1 U7495 ( .B1(n4492), .B2(keyinput115), .C1(n6569), .C2(keyinput105), 
        .A(n6568), .ZN(n6577) );
  AOI22_X1 U7496 ( .A1(n6571), .A2(keyinput110), .B1(keyinput73), .B2(n6690), 
        .ZN(n6570) );
  OAI221_X1 U7497 ( .B1(n6571), .B2(keyinput110), .C1(n6690), .C2(keyinput73), 
        .A(n6570), .ZN(n6576) );
  AOI22_X1 U7498 ( .A1(n6574), .A2(keyinput71), .B1(n6573), .B2(keyinput85), 
        .ZN(n6572) );
  OAI221_X1 U7499 ( .B1(n6574), .B2(keyinput71), .C1(n6573), .C2(keyinput85), 
        .A(n6572), .ZN(n6575) );
  NOR4_X1 U7500 ( .A1(n6578), .A2(n6577), .A3(n6576), .A4(n6575), .ZN(n6615)
         );
  AOI22_X1 U7501 ( .A1(DATAI_4_), .A2(keyinput96), .B1(EBX_REG_26__SCAN_IN), 
        .B2(keyinput99), .ZN(n6579) );
  OAI221_X1 U7502 ( .B1(DATAI_4_), .B2(keyinput96), .C1(EBX_REG_26__SCAN_IN), 
        .C2(keyinput99), .A(n6579), .ZN(n6587) );
  AOI22_X1 U7503 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput76), .B1(
        INSTQUEUE_REG_15__7__SCAN_IN), .B2(keyinput119), .ZN(n6580) );
  OAI221_X1 U7504 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput76), .C1(
        INSTQUEUE_REG_15__7__SCAN_IN), .C2(keyinput119), .A(n6580), .ZN(n6586)
         );
  AOI22_X1 U7505 ( .A1(n5234), .A2(keyinput94), .B1(keyinput89), .B2(n6725), 
        .ZN(n6581) );
  OAI221_X1 U7506 ( .B1(n5234), .B2(keyinput94), .C1(n6725), .C2(keyinput89), 
        .A(n6581), .ZN(n6585) );
  INV_X1 U7507 ( .A(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n6583) );
  AOI22_X1 U7508 ( .A1(EBX_REG_13__SCAN_IN), .A2(keyinput70), .B1(n6583), .B2(
        keyinput91), .ZN(n6582) );
  OAI221_X1 U7509 ( .B1(EBX_REG_13__SCAN_IN), .B2(keyinput70), .C1(n6583), 
        .C2(keyinput91), .A(n6582), .ZN(n6584) );
  NOR4_X1 U7510 ( .A1(n6587), .A2(n6586), .A3(n6585), .A4(n6584), .ZN(n6614)
         );
  AOI22_X1 U7511 ( .A1(n6589), .A2(keyinput66), .B1(n4481), .B2(keyinput116), 
        .ZN(n6588) );
  OAI221_X1 U7512 ( .B1(n6589), .B2(keyinput66), .C1(n4481), .C2(keyinput116), 
        .A(n6588), .ZN(n6599) );
  INV_X1 U7513 ( .A(DATAI_20_), .ZN(n6696) );
  AOI22_X1 U7514 ( .A1(n6591), .A2(keyinput82), .B1(n6696), .B2(keyinput95), 
        .ZN(n6590) );
  OAI221_X1 U7515 ( .B1(n6591), .B2(keyinput82), .C1(n6696), .C2(keyinput95), 
        .A(n6590), .ZN(n6598) );
  INV_X1 U7516 ( .A(BS16_N), .ZN(n6742) );
  AOI22_X1 U7517 ( .A1(n6593), .A2(keyinput122), .B1(keyinput124), .B2(n6742), 
        .ZN(n6592) );
  OAI221_X1 U7518 ( .B1(n6593), .B2(keyinput122), .C1(n6742), .C2(keyinput124), 
        .A(n6592), .ZN(n6597) );
  INV_X1 U7519 ( .A(UWORD_REG_11__SCAN_IN), .ZN(n6595) );
  AOI22_X1 U7520 ( .A1(n6743), .A2(keyinput64), .B1(keyinput125), .B2(n6595), 
        .ZN(n6594) );
  OAI221_X1 U7521 ( .B1(n6743), .B2(keyinput64), .C1(n6595), .C2(keyinput125), 
        .A(n6594), .ZN(n6596) );
  NOR4_X1 U7522 ( .A1(n6599), .A2(n6598), .A3(n6597), .A4(n6596), .ZN(n6613)
         );
  AOI22_X1 U7523 ( .A1(n6692), .A2(keyinput79), .B1(n6719), .B2(keyinput83), 
        .ZN(n6600) );
  OAI221_X1 U7524 ( .B1(n6692), .B2(keyinput79), .C1(n6719), .C2(keyinput83), 
        .A(n6600), .ZN(n6611) );
  INV_X1 U7525 ( .A(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n6602) );
  AOI22_X1 U7526 ( .A1(n6737), .A2(keyinput120), .B1(n6602), .B2(keyinput90), 
        .ZN(n6601) );
  OAI221_X1 U7527 ( .B1(n6737), .B2(keyinput120), .C1(n6602), .C2(keyinput90), 
        .A(n6601), .ZN(n6610) );
  AOI22_X1 U7528 ( .A1(n6605), .A2(keyinput109), .B1(n6604), .B2(keyinput117), 
        .ZN(n6603) );
  OAI221_X1 U7529 ( .B1(n6605), .B2(keyinput109), .C1(n6604), .C2(keyinput117), 
        .A(n6603), .ZN(n6609) );
  AOI22_X1 U7530 ( .A1(n6607), .A2(keyinput77), .B1(keyinput98), .B2(n6736), 
        .ZN(n6606) );
  OAI221_X1 U7531 ( .B1(n6607), .B2(keyinput77), .C1(n6736), .C2(keyinput98), 
        .A(n6606), .ZN(n6608) );
  NOR4_X1 U7532 ( .A1(n6611), .A2(n6610), .A3(n6609), .A4(n6608), .ZN(n6612)
         );
  AND4_X1 U7533 ( .A1(n6615), .A2(n6614), .A3(n6613), .A4(n6612), .ZN(n6755)
         );
  OAI22_X1 U7534 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(keyinput123), .B1(
        keyinput74), .B2(EAX_REG_22__SCAN_IN), .ZN(n6616) );
  AOI221_X1 U7535 ( .B1(INSTQUEUE_REG_12__7__SCAN_IN), .B2(keyinput123), .C1(
        EAX_REG_22__SCAN_IN), .C2(keyinput74), .A(n6616), .ZN(n6623) );
  OAI22_X1 U7536 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(keyinput80), .B1(
        keyinput121), .B2(DATAO_REG_30__SCAN_IN), .ZN(n6617) );
  AOI221_X1 U7537 ( .B1(INSTQUEUE_REG_8__1__SCAN_IN), .B2(keyinput80), .C1(
        DATAO_REG_30__SCAN_IN), .C2(keyinput121), .A(n6617), .ZN(n6622) );
  OAI22_X1 U7538 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(keyinput65), .B1(
        keyinput81), .B2(DATAI_31_), .ZN(n6618) );
  AOI221_X1 U7539 ( .B1(INSTQUEUE_REG_10__4__SCAN_IN), .B2(keyinput65), .C1(
        DATAI_31_), .C2(keyinput81), .A(n6618), .ZN(n6621) );
  OAI22_X1 U7540 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(keyinput103), .B1(
        keyinput114), .B2(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6619) );
  AOI221_X1 U7541 ( .B1(INSTQUEUE_REG_9__3__SCAN_IN), .B2(keyinput103), .C1(
        INSTADDRPOINTER_REG_12__SCAN_IN), .C2(keyinput114), .A(n6619), .ZN(
        n6620) );
  NAND4_X1 U7542 ( .A1(n6623), .A2(n6622), .A3(n6621), .A4(n6620), .ZN(n6651)
         );
  OAI22_X1 U7543 ( .A1(EBX_REG_7__SCAN_IN), .A2(keyinput68), .B1(keyinput108), 
        .B2(REIP_REG_19__SCAN_IN), .ZN(n6624) );
  AOI221_X1 U7544 ( .B1(EBX_REG_7__SCAN_IN), .B2(keyinput68), .C1(
        REIP_REG_19__SCAN_IN), .C2(keyinput108), .A(n6624), .ZN(n6631) );
  OAI22_X1 U7545 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(keyinput97), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(keyinput118), .ZN(n6625) );
  AOI221_X1 U7546 ( .B1(INSTQUEUE_REG_9__0__SCAN_IN), .B2(keyinput97), .C1(
        keyinput118), .C2(ADDRESS_REG_26__SCAN_IN), .A(n6625), .ZN(n6630) );
  OAI22_X1 U7547 ( .A1(EBX_REG_29__SCAN_IN), .A2(keyinput88), .B1(
        DATAO_REG_1__SCAN_IN), .B2(keyinput104), .ZN(n6626) );
  AOI221_X1 U7548 ( .B1(EBX_REG_29__SCAN_IN), .B2(keyinput88), .C1(keyinput104), .C2(DATAO_REG_1__SCAN_IN), .A(n6626), .ZN(n6629) );
  OAI22_X1 U7549 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(keyinput78), .B1(
        DATAI_23_), .B2(keyinput106), .ZN(n6627) );
  AOI221_X1 U7550 ( .B1(INSTQUEUE_REG_7__6__SCAN_IN), .B2(keyinput78), .C1(
        keyinput106), .C2(DATAI_23_), .A(n6627), .ZN(n6628) );
  NAND4_X1 U7551 ( .A1(n6631), .A2(n6630), .A3(n6629), .A4(n6628), .ZN(n6650)
         );
  OAI22_X1 U7552 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(keyinput84), .B1(
        keyinput127), .B2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n6632) );
  AOI221_X1 U7553 ( .B1(INSTQUEUE_REG_7__5__SCAN_IN), .B2(keyinput84), .C1(
        INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(keyinput127), .A(n6632), .ZN(
        n6639) );
  OAI22_X1 U7554 ( .A1(INSTQUEUE_REG_14__3__SCAN_IN), .A2(keyinput86), .B1(
        keyinput126), .B2(EAX_REG_26__SCAN_IN), .ZN(n6633) );
  AOI221_X1 U7555 ( .B1(INSTQUEUE_REG_14__3__SCAN_IN), .B2(keyinput86), .C1(
        EAX_REG_26__SCAN_IN), .C2(keyinput126), .A(n6633), .ZN(n6638) );
  OAI22_X1 U7556 ( .A1(REIP_REG_1__SCAN_IN), .A2(keyinput111), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(keyinput93), .ZN(n6634) );
  AOI221_X1 U7557 ( .B1(REIP_REG_1__SCAN_IN), .B2(keyinput111), .C1(keyinput93), .C2(ADDRESS_REG_22__SCAN_IN), .A(n6634), .ZN(n6637) );
  OAI22_X1 U7558 ( .A1(STATE_REG_1__SCAN_IN), .A2(keyinput92), .B1(keyinput107), .B2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n6635) );
  AOI221_X1 U7559 ( .B1(STATE_REG_1__SCAN_IN), .B2(keyinput92), .C1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .C2(keyinput107), .A(n6635), .ZN(
        n6636) );
  NAND4_X1 U7560 ( .A1(n6639), .A2(n6638), .A3(n6637), .A4(n6636), .ZN(n6649)
         );
  OAI22_X1 U7561 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(keyinput101), .B1(
        INSTQUEUE_REG_1__6__SCAN_IN), .B2(keyinput102), .ZN(n6640) );
  AOI221_X1 U7562 ( .B1(INSTQUEUE_REG_8__0__SCAN_IN), .B2(keyinput101), .C1(
        keyinput102), .C2(INSTQUEUE_REG_1__6__SCAN_IN), .A(n6640), .ZN(n6647)
         );
  OAI22_X1 U7563 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(keyinput69), .B1(
        DATAO_REG_2__SCAN_IN), .B2(keyinput75), .ZN(n6641) );
  AOI221_X1 U7564 ( .B1(INSTQUEUE_REG_0__6__SCAN_IN), .B2(keyinput69), .C1(
        keyinput75), .C2(DATAO_REG_2__SCAN_IN), .A(n6641), .ZN(n6646) );
  OAI22_X1 U7565 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(keyinput112), 
        .B1(keyinput113), .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6642) );
  AOI221_X1 U7566 ( .B1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(keyinput112), 
        .C1(INSTQUEUE_REG_10__6__SCAN_IN), .C2(keyinput113), .A(n6642), .ZN(
        n6645) );
  OAI22_X1 U7567 ( .A1(EBX_REG_6__SCAN_IN), .A2(keyinput87), .B1(DATAI_26_), 
        .B2(keyinput67), .ZN(n6643) );
  AOI221_X1 U7568 ( .B1(EBX_REG_6__SCAN_IN), .B2(keyinput87), .C1(keyinput67), 
        .C2(DATAI_26_), .A(n6643), .ZN(n6644) );
  NAND4_X1 U7569 ( .A1(n6647), .A2(n6646), .A3(n6645), .A4(n6644), .ZN(n6648)
         );
  NOR4_X1 U7570 ( .A1(n6651), .A2(n6650), .A3(n6649), .A4(n6648), .ZN(n6754)
         );
  AOI22_X1 U7571 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(keyinput55), .B1(
        INSTQUEUE_REG_9__4__SCAN_IN), .B2(keyinput27), .ZN(n6652) );
  OAI221_X1 U7572 ( .B1(INSTQUEUE_REG_15__7__SCAN_IN), .B2(keyinput55), .C1(
        INSTQUEUE_REG_9__4__SCAN_IN), .C2(keyinput27), .A(n6652), .ZN(n6659)
         );
  AOI22_X1 U7573 ( .A1(DATAI_31_), .A2(keyinput17), .B1(
        INSTQUEUE_REG_10__4__SCAN_IN), .B2(keyinput1), .ZN(n6653) );
  OAI221_X1 U7574 ( .B1(DATAI_31_), .B2(keyinput17), .C1(
        INSTQUEUE_REG_10__4__SCAN_IN), .C2(keyinput1), .A(n6653), .ZN(n6658)
         );
  AOI22_X1 U7575 ( .A1(PHYADDRPOINTER_REG_17__SCAN_IN), .A2(keyinput43), .B1(
        INSTQUEUE_REG_1__6__SCAN_IN), .B2(keyinput38), .ZN(n6654) );
  OAI221_X1 U7576 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput43), .C1(
        INSTQUEUE_REG_1__6__SCAN_IN), .C2(keyinput38), .A(n6654), .ZN(n6657)
         );
  AOI22_X1 U7577 ( .A1(UWORD_REG_11__SCAN_IN), .A2(keyinput61), .B1(
        INSTADDRPOINTER_REG_13__SCAN_IN), .B2(keyinput46), .ZN(n6655) );
  OAI221_X1 U7578 ( .B1(UWORD_REG_11__SCAN_IN), .B2(keyinput61), .C1(
        INSTADDRPOINTER_REG_13__SCAN_IN), .C2(keyinput46), .A(n6655), .ZN(
        n6656) );
  NOR4_X1 U7579 ( .A1(n6659), .A2(n6658), .A3(n6657), .A4(n6656), .ZN(n6687)
         );
  AOI22_X1 U7580 ( .A1(EBX_REG_7__SCAN_IN), .A2(keyinput4), .B1(
        INSTQUEUE_REG_8__0__SCAN_IN), .B2(keyinput37), .ZN(n6660) );
  OAI221_X1 U7581 ( .B1(EBX_REG_7__SCAN_IN), .B2(keyinput4), .C1(
        INSTQUEUE_REG_8__0__SCAN_IN), .C2(keyinput37), .A(n6660), .ZN(n6667)
         );
  AOI22_X1 U7582 ( .A1(DATAO_REG_11__SCAN_IN), .A2(keyinput7), .B1(
        REIP_REG_1__SCAN_IN), .B2(keyinput47), .ZN(n6661) );
  OAI221_X1 U7583 ( .B1(DATAO_REG_11__SCAN_IN), .B2(keyinput7), .C1(
        REIP_REG_1__SCAN_IN), .C2(keyinput47), .A(n6661), .ZN(n6666) );
  AOI22_X1 U7584 ( .A1(DATAI_6_), .A2(keyinput58), .B1(STATE_REG_1__SCAN_IN), 
        .B2(keyinput28), .ZN(n6662) );
  OAI221_X1 U7585 ( .B1(DATAI_6_), .B2(keyinput58), .C1(STATE_REG_1__SCAN_IN), 
        .C2(keyinput28), .A(n6662), .ZN(n6665) );
  AOI22_X1 U7586 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(keyinput2), .B1(
        EBX_REG_6__SCAN_IN), .B2(keyinput23), .ZN(n6663) );
  OAI221_X1 U7587 ( .B1(DATAWIDTH_REG_21__SCAN_IN), .B2(keyinput2), .C1(
        EBX_REG_6__SCAN_IN), .C2(keyinput23), .A(n6663), .ZN(n6664) );
  NOR4_X1 U7588 ( .A1(n6667), .A2(n6666), .A3(n6665), .A4(n6664), .ZN(n6686)
         );
  AOI22_X1 U7589 ( .A1(REIP_REG_14__SCAN_IN), .A2(keyinput45), .B1(
        INSTQUEUE_REG_9__0__SCAN_IN), .B2(keyinput33), .ZN(n6668) );
  OAI221_X1 U7590 ( .B1(REIP_REG_14__SCAN_IN), .B2(keyinput45), .C1(
        INSTQUEUE_REG_9__0__SCAN_IN), .C2(keyinput33), .A(n6668), .ZN(n6675)
         );
  AOI22_X1 U7591 ( .A1(DATAI_5_), .A2(keyinput41), .B1(
        INSTADDRPOINTER_REG_12__SCAN_IN), .B2(keyinput50), .ZN(n6669) );
  OAI221_X1 U7592 ( .B1(DATAI_5_), .B2(keyinput41), .C1(
        INSTADDRPOINTER_REG_12__SCAN_IN), .C2(keyinput50), .A(n6669), .ZN(
        n6674) );
  AOI22_X1 U7593 ( .A1(INSTQUEUE_REG_12__3__SCAN_IN), .A2(keyinput52), .B1(
        INSTQUEUE_REG_14__3__SCAN_IN), .B2(keyinput22), .ZN(n6670) );
  OAI221_X1 U7594 ( .B1(INSTQUEUE_REG_12__3__SCAN_IN), .B2(keyinput52), .C1(
        INSTQUEUE_REG_14__3__SCAN_IN), .C2(keyinput22), .A(n6670), .ZN(n6673)
         );
  AOI22_X1 U7595 ( .A1(CODEFETCH_REG_SCAN_IN), .A2(keyinput12), .B1(
        INSTQUEUE_REG_8__1__SCAN_IN), .B2(keyinput16), .ZN(n6671) );
  OAI221_X1 U7596 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(keyinput12), .C1(
        INSTQUEUE_REG_8__1__SCAN_IN), .C2(keyinput16), .A(n6671), .ZN(n6672)
         );
  NOR4_X1 U7597 ( .A1(n6675), .A2(n6674), .A3(n6673), .A4(n6672), .ZN(n6685)
         );
  AOI22_X1 U7598 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(keyinput63), .B1(
        INSTQUEUE_REG_12__0__SCAN_IN), .B2(keyinput51), .ZN(n6676) );
  OAI221_X1 U7599 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(keyinput63), 
        .C1(INSTQUEUE_REG_12__0__SCAN_IN), .C2(keyinput51), .A(n6676), .ZN(
        n6683) );
  AOI22_X1 U7600 ( .A1(DATAI_23_), .A2(keyinput42), .B1(
        INSTQUEUE_REG_12__6__SCAN_IN), .B2(keyinput26), .ZN(n6677) );
  OAI221_X1 U7601 ( .B1(DATAI_23_), .B2(keyinput42), .C1(
        INSTQUEUE_REG_12__6__SCAN_IN), .C2(keyinput26), .A(n6677), .ZN(n6682)
         );
  AOI22_X1 U7602 ( .A1(REIP_REG_19__SCAN_IN), .A2(keyinput44), .B1(
        EAX_REG_22__SCAN_IN), .B2(keyinput10), .ZN(n6678) );
  OAI221_X1 U7603 ( .B1(REIP_REG_19__SCAN_IN), .B2(keyinput44), .C1(
        EAX_REG_22__SCAN_IN), .C2(keyinput10), .A(n6678), .ZN(n6681) );
  AOI22_X1 U7604 ( .A1(LWORD_REG_10__SCAN_IN), .A2(keyinput18), .B1(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(keyinput48), .ZN(n6679) );
  OAI221_X1 U7605 ( .B1(LWORD_REG_10__SCAN_IN), .B2(keyinput18), .C1(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(keyinput48), .A(n6679), .ZN(
        n6680) );
  NOR4_X1 U7606 ( .A1(n6683), .A2(n6682), .A3(n6681), .A4(n6680), .ZN(n6684)
         );
  NAND4_X1 U7607 ( .A1(n6687), .A2(n6686), .A3(n6685), .A4(n6684), .ZN(n6753)
         );
  AOI22_X1 U7608 ( .A1(n6690), .A2(keyinput9), .B1(keyinput29), .B2(n6689), 
        .ZN(n6688) );
  OAI221_X1 U7609 ( .B1(n6690), .B2(keyinput9), .C1(n6689), .C2(keyinput29), 
        .A(n6688), .ZN(n6702) );
  AOI22_X1 U7610 ( .A1(n6692), .A2(keyinput15), .B1(n5234), .B2(keyinput30), 
        .ZN(n6691) );
  OAI221_X1 U7611 ( .B1(n6692), .B2(keyinput15), .C1(n5234), .C2(keyinput30), 
        .A(n6691), .ZN(n6701) );
  INV_X1 U7612 ( .A(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n6694) );
  AOI22_X1 U7613 ( .A1(n6695), .A2(keyinput6), .B1(n6694), .B2(keyinput39), 
        .ZN(n6693) );
  OAI221_X1 U7614 ( .B1(n6695), .B2(keyinput6), .C1(n6694), .C2(keyinput39), 
        .A(n6693), .ZN(n6700) );
  XOR2_X1 U7615 ( .A(n6696), .B(keyinput31), .Z(n6698) );
  XNOR2_X1 U7616 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .B(keyinput5), .ZN(n6697)
         );
  NAND2_X1 U7617 ( .A1(n6698), .A2(n6697), .ZN(n6699) );
  NOR4_X1 U7618 ( .A1(n6702), .A2(n6701), .A3(n6700), .A4(n6699), .ZN(n6751)
         );
  AOI22_X1 U7619 ( .A1(n6705), .A2(keyinput57), .B1(n6704), .B2(keyinput35), 
        .ZN(n6703) );
  OAI221_X1 U7620 ( .B1(n6705), .B2(keyinput57), .C1(n6704), .C2(keyinput35), 
        .A(n6703), .ZN(n6716) );
  AOI22_X1 U7621 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(keyinput13), .B1(
        EAX_REG_25__SCAN_IN), .B2(keyinput21), .ZN(n6706) );
  OAI221_X1 U7622 ( .B1(DATAWIDTH_REG_23__SCAN_IN), .B2(keyinput13), .C1(
        EAX_REG_25__SCAN_IN), .C2(keyinput21), .A(n6706), .ZN(n6715) );
  INV_X1 U7623 ( .A(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n6709) );
  INV_X1 U7624 ( .A(DATAO_REG_1__SCAN_IN), .ZN(n6708) );
  AOI22_X1 U7625 ( .A1(n6709), .A2(keyinput14), .B1(keyinput40), .B2(n6708), 
        .ZN(n6707) );
  OAI221_X1 U7626 ( .B1(n6709), .B2(keyinput14), .C1(n6708), .C2(keyinput40), 
        .A(n6707), .ZN(n6714) );
  INV_X1 U7627 ( .A(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n6712) );
  INV_X1 U7628 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n6711) );
  AOI22_X1 U7629 ( .A1(n6712), .A2(keyinput20), .B1(keyinput11), .B2(n6711), 
        .ZN(n6710) );
  OAI221_X1 U7630 ( .B1(n6712), .B2(keyinput20), .C1(n6711), .C2(keyinput11), 
        .A(n6710), .ZN(n6713) );
  NOR4_X1 U7631 ( .A1(n6716), .A2(n6715), .A3(n6714), .A4(n6713), .ZN(n6750)
         );
  AOI22_X1 U7632 ( .A1(n6719), .A2(keyinput19), .B1(n6718), .B2(keyinput8), 
        .ZN(n6717) );
  OAI221_X1 U7633 ( .B1(n6719), .B2(keyinput19), .C1(n6718), .C2(keyinput8), 
        .A(n6717), .ZN(n6731) );
  AOI22_X1 U7634 ( .A1(n6722), .A2(keyinput54), .B1(n6721), .B2(keyinput32), 
        .ZN(n6720) );
  OAI221_X1 U7635 ( .B1(n6722), .B2(keyinput54), .C1(n6721), .C2(keyinput32), 
        .A(n6720), .ZN(n6730) );
  AOI22_X1 U7636 ( .A1(n6725), .A2(keyinput25), .B1(n6724), .B2(keyinput24), 
        .ZN(n6723) );
  OAI221_X1 U7637 ( .B1(n6725), .B2(keyinput25), .C1(n6724), .C2(keyinput24), 
        .A(n6723), .ZN(n6729) );
  XNOR2_X1 U7638 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(keyinput53), .ZN(
        n6727) );
  XNOR2_X1 U7639 ( .A(INSTQUEUE_REG_12__7__SCAN_IN), .B(keyinput59), .ZN(n6726) );
  NAND2_X1 U7640 ( .A1(n6727), .A2(n6726), .ZN(n6728) );
  NOR4_X1 U7641 ( .A1(n6731), .A2(n6730), .A3(n6729), .A4(n6728), .ZN(n6749)
         );
  INV_X1 U7642 ( .A(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n6734) );
  AOI22_X1 U7643 ( .A1(n6734), .A2(keyinput49), .B1(keyinput62), .B2(n6733), 
        .ZN(n6732) );
  OAI221_X1 U7644 ( .B1(n6734), .B2(keyinput49), .C1(n6733), .C2(keyinput62), 
        .A(n6732), .ZN(n6747) );
  AOI22_X1 U7645 ( .A1(n6737), .A2(keyinput56), .B1(keyinput34), .B2(n6736), 
        .ZN(n6735) );
  OAI221_X1 U7646 ( .B1(n6737), .B2(keyinput56), .C1(n6736), .C2(keyinput34), 
        .A(n6735), .ZN(n6746) );
  AOI22_X1 U7647 ( .A1(n6740), .A2(keyinput3), .B1(n6739), .B2(keyinput36), 
        .ZN(n6738) );
  OAI221_X1 U7648 ( .B1(n6740), .B2(keyinput3), .C1(n6739), .C2(keyinput36), 
        .A(n6738), .ZN(n6745) );
  AOI22_X1 U7649 ( .A1(n6743), .A2(keyinput0), .B1(keyinput60), .B2(n6742), 
        .ZN(n6741) );
  OAI221_X1 U7650 ( .B1(n6743), .B2(keyinput0), .C1(n6742), .C2(keyinput60), 
        .A(n6741), .ZN(n6744) );
  NOR4_X1 U7651 ( .A1(n6747), .A2(n6746), .A3(n6745), .A4(n6744), .ZN(n6748)
         );
  NAND4_X1 U7652 ( .A1(n6751), .A2(n6750), .A3(n6749), .A4(n6748), .ZN(n6752)
         );
  AOI211_X1 U7653 ( .C1(n6755), .C2(n6754), .A(n6753), .B(n6752), .ZN(n6756)
         );
  XNOR2_X1 U7654 ( .A(n6757), .B(n6756), .ZN(U2844) );
  CLKBUF_X2 U3457 ( .A(n3017), .Z(n3794) );
  BUF_X2 U3569 ( .A(n3133), .Z(n3279) );
  CLKBUF_X1 U3655 ( .A(n3932), .Z(n4004) );
endmodule

