

module b14_C_SARLock_k_64_4 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386,
         n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396,
         n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406,
         n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
         n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426,
         n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436,
         n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446,
         n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456,
         n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466,
         n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476,
         n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486,
         n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496,
         n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506,
         n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
         n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536,
         n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546,
         n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556,
         n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566,
         n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576,
         n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586,
         n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596,
         n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606,
         n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616,
         n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626,
         n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636,
         n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
         n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
         n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666,
         n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676,
         n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686,
         n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694;

  AOI21_X1 U2259 ( .B1(n4215), .B2(n4533), .A(n2136), .ZN(n2139) );
  CLKBUF_X1 U2260 ( .A(n2330), .Z(n2705) );
  CLKBUF_X2 U2261 ( .A(n2370), .Z(n3622) );
  INV_X2 U2262 ( .A(n2321), .ZN(n2737) );
  INV_X1 U2263 ( .A(n2741), .ZN(n2753) );
  OR2_X1 U2264 ( .A1(n3921), .A2(n3903), .ZN(n3907) );
  CLKBUF_X2 U2265 ( .A(n2370), .Z(n2712) );
  AND2_X1 U2266 ( .A1(n2930), .A2(n2744), .ZN(n2787) );
  OR2_X1 U2267 ( .A1(n2019), .A2(n2064), .ZN(n2063) );
  XNOR2_X1 U2268 ( .A(n2278), .B(IR_REG_30__SCAN_IN), .ZN(n4337) );
  NAND2_X4 U2269 ( .A1(n2304), .A2(n2295), .ZN(n2321) );
  INV_X1 U2270 ( .A(n2442), .ZN(n2016) );
  NOR2_X2 U2271 ( .A1(n3218), .A2(n3204), .ZN(n3249) );
  NAND2_X2 U2272 ( .A1(n2400), .A2(n2399), .ZN(n3288) );
  INV_X2 U2273 ( .A(n4195), .ZN(n2017) );
  OAI21_X1 U2274 ( .B1(n4215), .B2(n2063), .A(n4692), .ZN(n2062) );
  MUX2_X1 U2275 ( .A(n2925), .B(REG0_REG_28__SCAN_IN), .S(n4690), .Z(n2926) );
  AOI21_X1 U2276 ( .B1(n2019), .B2(n4533), .A(n2056), .ZN(n2137) );
  MUX2_X1 U2277 ( .A(REG1_REG_28__SCAN_IN), .B(n2925), .S(n4533), .Z(n2915) );
  OAI21_X1 U2278 ( .B1(n3952), .B2(n3693), .A(n2899), .ZN(n3912) );
  OR2_X1 U2279 ( .A1(n4136), .A2(n3745), .ZN(n4137) );
  NAND2_X1 U2280 ( .A1(n3345), .A2(n2482), .ZN(n3370) );
  NAND2_X1 U2281 ( .A1(n3341), .A2(n2477), .ZN(n3345) );
  OAI21_X1 U2282 ( .B1(n3211), .B2(n2873), .A(n3653), .ZN(n3200) );
  AOI21_X1 U2283 ( .B1(n3392), .B2(n3391), .A(n2240), .ZN(n2239) );
  NAND2_X1 U2284 ( .A1(n4364), .A2(n2170), .ZN(n3831) );
  NAND2_X2 U2285 ( .A1(n3111), .A2(n4193), .ZN(n4195) );
  NAND2_X1 U2286 ( .A1(n2877), .A2(n3658), .ZN(n3240) );
  AND2_X1 U2287 ( .A1(n3647), .A2(n3644), .ZN(n3708) );
  XNOR2_X1 U2288 ( .A(n2163), .B(n2162), .ZN(n3031) );
  NAND2_X1 U2289 ( .A1(n3779), .A2(n3231), .ZN(n3658) );
  INV_X1 U2290 ( .A(n2833), .ZN(n3779) );
  NOR2_X2 U2291 ( .A1(n3004), .A2(n3003), .ZN(n4429) );
  OR2_X1 U2292 ( .A1(n2206), .A2(n2252), .ZN(n3780) );
  INV_X1 U2293 ( .A(n2874), .ZN(n3204) );
  NAND4_X1 U2294 ( .A1(n2260), .A2(n2285), .A3(n2284), .A4(n2283), .ZN(n3784)
         );
  CLKBUF_X1 U2295 ( .A(n2672), .Z(n3606) );
  NAND2_X1 U2296 ( .A1(n2302), .A2(n2301), .ZN(n2370) );
  AND2_X1 U2297 ( .A1(n2791), .A2(n3757), .ZN(n4452) );
  AND2_X1 U2298 ( .A1(n4339), .A2(n2968), .ZN(n2100) );
  XNOR2_X1 U2299 ( .A(n2288), .B(IR_REG_24__SCAN_IN), .ZN(n4340) );
  OR2_X1 U2300 ( .A1(n2989), .A2(n2298), .ZN(n2300) );
  XNOR2_X1 U2301 ( .A(n2306), .B(IR_REG_22__SCAN_IN), .ZN(n4341) );
  XNOR2_X1 U2302 ( .A(n2292), .B(n2291), .ZN(n2795) );
  XNOR2_X1 U2303 ( .A(n2294), .B(IR_REG_21__SCAN_IN), .ZN(n3641) );
  OR2_X1 U2304 ( .A1(n3444), .A2(n2601), .ZN(n2278) );
  XNOR2_X1 U2305 ( .A(n2286), .B(IR_REG_26__SCAN_IN), .ZN(n2968) );
  INV_X1 U2306 ( .A(IR_REG_3__SCAN_IN), .ZN(n2353) );
  INV_X1 U2307 ( .A(IR_REG_27__SCAN_IN), .ZN(n2298) );
  INV_X1 U2308 ( .A(IR_REG_15__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U2309 ( .A1(n2312), .A2(n2311), .ZN(n2314) );
  NOR2_X1 U2310 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2335)
         );
  INV_X1 U2311 ( .A(n2705), .ZN(n2806) );
  CLKBUF_X3 U2312 ( .A(n2347), .Z(n2973) );
  NOR2_X1 U2313 ( .A1(n4337), .A2(n2962), .ZN(n2347) );
  NAND2_X1 U2314 ( .A1(n2122), .A2(n2697), .ZN(n2121) );
  NAND2_X1 U2315 ( .A1(n2123), .A2(n2234), .ZN(n2122) );
  NAND2_X1 U2316 ( .A1(n3812), .A2(n2034), .ZN(n2166) );
  NAND2_X1 U2317 ( .A1(n3012), .A2(n4347), .ZN(n2160) );
  AOI21_X1 U2318 ( .B1(n3849), .B2(REG1_REG_13__SCAN_IN), .A(n4390), .ZN(n3850) );
  NOR2_X1 U2319 ( .A1(n2185), .A2(n2027), .ZN(n2184) );
  NOR2_X1 U2320 ( .A1(n2244), .A2(n2204), .ZN(n2203) );
  INV_X1 U2321 ( .A(n2270), .ZN(n2204) );
  INV_X1 U2322 ( .A(IR_REG_19__SCAN_IN), .ZN(n2311) );
  AND4_X1 U2323 ( .A1(n2264), .A2(n2263), .A3(n2262), .A4(n2502), .ZN(n2265)
         );
  NOR2_X1 U2324 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .ZN(n2263)
         );
  NOR2_X1 U2325 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2262)
         );
  NAND2_X1 U2326 ( .A1(n2118), .A2(n3598), .ZN(n2117) );
  AND2_X1 U2327 ( .A1(n3513), .A2(n3520), .ZN(n2232) );
  INV_X1 U2328 ( .A(n2559), .ZN(n2118) );
  AND2_X1 U2329 ( .A1(n2985), .A2(n2796), .ZN(n2908) );
  NAND2_X1 U2330 ( .A1(n2992), .A2(n2993), .ZN(n3804) );
  AOI21_X1 U2331 ( .B1(n2084), .B2(n2080), .A(n3055), .ZN(n2079) );
  NAND2_X1 U2332 ( .A1(n3038), .A2(n2211), .ZN(n2210) );
  INV_X1 U2333 ( .A(n4360), .ZN(n2211) );
  XNOR2_X1 U2334 ( .A(n3831), .B(n2169), .ZN(n3032) );
  OR2_X1 U2335 ( .A1(n4403), .A2(n4404), .ZN(n2090) );
  NOR2_X1 U2336 ( .A1(n2733), .A2(n4662), .ZN(n2745) );
  OR2_X1 U2337 ( .A1(n4073), .A2(n4094), .ZN(n2853) );
  NAND2_X1 U2338 ( .A1(n2845), .A2(n2181), .ZN(n2176) );
  INV_X1 U2339 ( .A(n2178), .ZN(n2177) );
  NAND2_X1 U2340 ( .A1(n3273), .A2(n3659), .ZN(n2879) );
  NAND2_X1 U2341 ( .A1(n2300), .A2(n2299), .ZN(n2302) );
  AND3_X1 U2342 ( .A1(n2751), .A2(n2750), .A3(n2749), .ZN(n3898) );
  OR2_X1 U2343 ( .A1(n4351), .A2(n2903), .ZN(n4184) );
  NAND2_X1 U2344 ( .A1(n3112), .A2(n4453), .ZN(n3185) );
  AND2_X1 U2345 ( .A1(n2265), .A2(n2266), .ZN(n2205) );
  INV_X1 U2346 ( .A(IR_REG_13__SCAN_IN), .ZN(n2266) );
  AND2_X1 U2347 ( .A1(n4671), .A2(n2226), .ZN(n2224) );
  INV_X1 U2348 ( .A(IR_REG_5__SCAN_IN), .ZN(n2226) );
  NAND2_X1 U2349 ( .A1(n4433), .A2(n2221), .ZN(n2220) );
  NAND2_X1 U2350 ( .A1(n4468), .A2(n4596), .ZN(n2221) );
  XNOR2_X1 U2351 ( .A(n2175), .B(n2174), .ZN(n4214) );
  INV_X1 U2352 ( .A(n3906), .ZN(n2174) );
  NAND2_X1 U2353 ( .A1(n2144), .A2(n2142), .ZN(n2141) );
  AND2_X1 U2354 ( .A1(n2143), .A2(n4502), .ZN(n2142) );
  NAND2_X1 U2355 ( .A1(n2106), .A2(n2108), .ZN(n2103) );
  XNOR2_X1 U2356 ( .A(n2243), .B(n2753), .ZN(n2357) );
  OAI21_X1 U2357 ( .B1(n3178), .B2(n2321), .A(n2356), .ZN(n2243) );
  NOR2_X1 U2358 ( .A1(n3392), .A2(n2131), .ZN(n2130) );
  INV_X1 U2359 ( .A(n2133), .ZN(n2131) );
  AOI21_X1 U2360 ( .B1(n3010), .B2(REG2_REG_3__SCAN_IN), .A(n2039), .ZN(n3011)
         );
  AOI21_X1 U2361 ( .B1(n3017), .B2(REG1_REG_3__SCAN_IN), .A(n2038), .ZN(n3018)
         );
  AOI21_X1 U2362 ( .B1(n4475), .B2(REG1_REG_11__SCAN_IN), .A(n4369), .ZN(n3847) );
  NAND2_X1 U2363 ( .A1(n3861), .A2(n3860), .ZN(n2168) );
  INV_X1 U2364 ( .A(n2860), .ZN(n2193) );
  NAND2_X1 U2365 ( .A1(n4126), .A2(n2065), .ZN(n4046) );
  NOR2_X1 U2366 ( .A1(n3685), .A2(n2066), .ZN(n2065) );
  AND2_X1 U2367 ( .A1(n3773), .A2(n3524), .ZN(n2852) );
  INV_X1 U2368 ( .A(n3710), .ZN(n2843) );
  NOR2_X1 U2369 ( .A1(n3421), .A2(n3407), .ZN(n2152) );
  AND2_X1 U2370 ( .A1(n3248), .A2(n3231), .ZN(n2151) );
  NOR2_X1 U2371 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2270)
         );
  INV_X1 U2372 ( .A(IR_REG_11__SCAN_IN), .ZN(n2502) );
  NAND2_X1 U2373 ( .A1(n2112), .A2(n2111), .ZN(n2110) );
  INV_X1 U2374 ( .A(n3312), .ZN(n2111) );
  INV_X1 U2375 ( .A(n3311), .ZN(n2112) );
  NAND2_X1 U2376 ( .A1(n3311), .A2(n3312), .ZN(n2109) );
  AND2_X1 U2377 ( .A1(n2682), .A2(n2124), .ZN(n2123) );
  NAND2_X1 U2378 ( .A1(n2233), .A2(n2125), .ZN(n2124) );
  INV_X1 U2379 ( .A(n2256), .ZN(n2125) );
  INV_X1 U2380 ( .A(n2109), .ZN(n2108) );
  INV_X1 U2381 ( .A(n2107), .ZN(n2106) );
  OAI21_X1 U2382 ( .B1(n2110), .B2(n2108), .A(n3286), .ZN(n2107) );
  OR2_X1 U2383 ( .A1(n3367), .A2(n3368), .ZN(n2134) );
  INV_X1 U2384 ( .A(n4112), .ZN(n3524) );
  NAND2_X1 U2385 ( .A1(n3595), .A2(n3598), .ZN(n2575) );
  NAND2_X1 U2386 ( .A1(n3130), .A2(n3131), .ZN(n2113) );
  OR2_X1 U2387 ( .A1(n2608), .A2(n2607), .ZN(n2628) );
  NOR2_X1 U2388 ( .A1(n2576), .A2(n2231), .ZN(n2230) );
  INV_X1 U2389 ( .A(n3520), .ZN(n2231) );
  INV_X1 U2390 ( .A(n3519), .ZN(n2228) );
  NAND2_X1 U2391 ( .A1(n2024), .A2(n2051), .ZN(n2115) );
  INV_X1 U2392 ( .A(n3598), .ZN(n2119) );
  OR2_X1 U2393 ( .A1(n2546), .A2(n3588), .ZN(n2579) );
  NAND2_X1 U2394 ( .A1(n2558), .A2(n2559), .ZN(n3595) );
  OR2_X1 U2395 ( .A1(n2558), .A2(n2559), .ZN(n3596) );
  NAND2_X1 U2396 ( .A1(n2973), .A2(REG0_REG_5__SCAN_IN), .ZN(n2207) );
  NAND2_X1 U2397 ( .A1(n2398), .A2(REG1_REG_5__SCAN_IN), .ZN(n2208) );
  AOI21_X1 U2398 ( .B1(n2160), .B2(n2157), .A(n3052), .ZN(n2156) );
  INV_X1 U2399 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2157) );
  INV_X1 U2400 ( .A(n2160), .ZN(n2158) );
  NAND2_X1 U2401 ( .A1(n2077), .A2(n2082), .ZN(n2075) );
  NAND2_X1 U2402 ( .A1(n2212), .A2(n2048), .ZN(n2074) );
  OR2_X1 U2403 ( .A1(n3067), .A2(n2164), .ZN(n2163) );
  AND2_X1 U2404 ( .A1(n4344), .A2(REG2_REG_7__SCAN_IN), .ZN(n2164) );
  OR2_X1 U2405 ( .A1(n4478), .A2(n4604), .ZN(n2170) );
  NAND2_X1 U2406 ( .A1(n3032), .A2(REG2_REG_10__SCAN_IN), .ZN(n3832) );
  XNOR2_X1 U2407 ( .A(n3847), .B(n2167), .ZN(n4381) );
  NAND2_X1 U2408 ( .A1(n4374), .A2(n3834), .ZN(n3835) );
  NAND2_X1 U2409 ( .A1(n2090), .A2(n2031), .ZN(n2089) );
  NAND2_X1 U2410 ( .A1(n2089), .A2(n2088), .ZN(n3869) );
  INV_X1 U2411 ( .A(n3852), .ZN(n2088) );
  XNOR2_X1 U2412 ( .A(n2168), .B(n4470), .ZN(n4420) );
  NAND2_X1 U2413 ( .A1(n4420), .A2(n4419), .ZN(n4418) );
  XNOR2_X1 U2414 ( .A(n3870), .B(n2566), .ZN(n4423) );
  AND2_X1 U2415 ( .A1(n3869), .A2(n3868), .ZN(n3870) );
  NAND2_X1 U2416 ( .A1(n4423), .A2(n4422), .ZN(n4421) );
  NAND2_X1 U2417 ( .A1(n2901), .A2(n2900), .ZN(n3914) );
  INV_X1 U2418 ( .A(n3912), .ZN(n2901) );
  OR2_X1 U2419 ( .A1(n2719), .A2(n2718), .ZN(n2733) );
  OR2_X1 U2420 ( .A1(n2628), .A2(n4583), .ZN(n2658) );
  NAND2_X1 U2421 ( .A1(n2197), .A2(n2196), .ZN(n4008) );
  AOI21_X1 U2422 ( .B1(n2188), .B2(n2186), .A(n2040), .ZN(n2185) );
  INV_X1 U2423 ( .A(n2851), .ZN(n2186) );
  INV_X1 U2424 ( .A(n2188), .ZN(n2187) );
  NOR2_X1 U2425 ( .A1(n2850), .A2(n2189), .ZN(n2188) );
  NAND2_X1 U2426 ( .A1(n4135), .A2(n2851), .ZN(n2190) );
  AOI21_X1 U2427 ( .B1(n4174), .B2(n2848), .A(n2180), .ZN(n4151) );
  AND2_X1 U2428 ( .A1(n4158), .A2(n4181), .ZN(n2180) );
  NAND2_X1 U2429 ( .A1(n2839), .A2(n2199), .ZN(n2198) );
  NOR2_X1 U2430 ( .A1(n2840), .A2(n2200), .ZN(n2199) );
  AND4_X1 U2431 ( .A1(n2488), .A2(n2487), .A3(n2486), .A4(n2485), .ZN(n3402)
         );
  OAI21_X1 U2432 ( .B1(n3226), .B2(n2878), .A(n3658), .ZN(n3273) );
  OAI21_X1 U2433 ( .B1(n3200), .B2(n3198), .A(n3663), .ZN(n3244) );
  NAND2_X1 U2434 ( .A1(n3220), .A2(n3219), .ZN(n3218) );
  NAND2_X1 U2435 ( .A1(n2872), .A2(n3649), .ZN(n3211) );
  NAND2_X1 U2436 ( .A1(n2795), .A2(n3641), .ZN(n3125) );
  NOR2_X2 U2437 ( .A1(n4190), .A2(n2916), .ZN(n4163) );
  NOR2_X1 U2438 ( .A1(n3185), .A2(n3186), .ZN(n3184) );
  AND2_X1 U2439 ( .A1(n2203), .A2(n2276), .ZN(n2202) );
  NOR2_X1 U2440 ( .A1(IR_REG_26__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2276)
         );
  NAND2_X1 U2441 ( .A1(n2272), .A2(n2248), .ZN(n2247) );
  INV_X1 U2442 ( .A(IR_REG_22__SCAN_IN), .ZN(n2272) );
  INV_X1 U2443 ( .A(IR_REG_21__SCAN_IN), .ZN(n2248) );
  OAI21_X1 U2444 ( .B1(n2293), .B2(n2247), .A(IR_REG_31__SCAN_IN), .ZN(n2780)
         );
  INV_X1 U2445 ( .A(IR_REG_23__SCAN_IN), .ZN(n2779) );
  NAND2_X1 U2446 ( .A1(n2314), .A2(n2313), .ZN(n4451) );
  INV_X1 U2447 ( .A(IR_REG_16__SCAN_IN), .ZN(n4670) );
  OR2_X1 U2448 ( .A1(n2404), .A2(n2403), .ZN(n3077) );
  NOR2_X1 U2449 ( .A1(n2335), .A2(n2601), .ZN(n2222) );
  INV_X1 U2450 ( .A(n4349), .ZN(n2148) );
  INV_X1 U2451 ( .A(n3780), .ZN(n2828) );
  OR2_X1 U2452 ( .A1(n2811), .A2(n2805), .ZN(n3581) );
  OR2_X1 U2453 ( .A1(n2811), .A2(n2810), .ZN(n3593) );
  OAI211_X1 U2454 ( .C1(n3924), .C2(n2806), .A(n2736), .B(n2735), .ZN(n3937)
         );
  INV_X1 U2455 ( .A(n4156), .ZN(n3774) );
  NAND2_X1 U2456 ( .A1(n2070), .A2(n2991), .ZN(n3800) );
  XNOR2_X1 U2457 ( .A(n3020), .B(n4345), .ZN(n3075) );
  NOR2_X1 U2458 ( .A1(n3069), .A2(n3068), .ZN(n3067) );
  NAND2_X1 U2459 ( .A1(n2210), .A2(n2025), .ZN(n2086) );
  AND2_X1 U2460 ( .A1(n2085), .A2(n3843), .ZN(n3844) );
  AND2_X1 U2461 ( .A1(n2086), .A2(REG1_REG_10__SCAN_IN), .ZN(n2085) );
  XNOR2_X1 U2462 ( .A(n3835), .B(n2167), .ZN(n4387) );
  NAND2_X1 U2463 ( .A1(n4387), .A2(REG2_REG_12__SCAN_IN), .ZN(n4386) );
  OAI21_X1 U2464 ( .B1(n3878), .B2(n2218), .A(n2217), .ZN(n2216) );
  AOI21_X1 U2465 ( .B1(n4429), .B2(ADDR_REG_18__SCAN_IN), .A(n3874), .ZN(n2217) );
  NOR2_X1 U2466 ( .A1(n2220), .A2(n3873), .ZN(n3878) );
  NAND2_X1 U2467 ( .A1(n2219), .A2(n4437), .ZN(n2218) );
  AND2_X1 U2468 ( .A1(n3044), .A2(n3765), .ZN(n4439) );
  NAND2_X1 U2469 ( .A1(n2220), .A2(n2057), .ZN(n2091) );
  INV_X1 U2470 ( .A(n2095), .ZN(n2092) );
  AND2_X1 U2471 ( .A1(n4096), .A2(n4502), .ZN(n4444) );
  INV_X1 U2473 ( .A(n2141), .ZN(n2064) );
  NAND2_X1 U2474 ( .A1(n3901), .A2(n3900), .ZN(n4215) );
  NAND2_X1 U2475 ( .A1(n3895), .A2(n4281), .ZN(n3901) );
  AND3_X1 U2476 ( .A1(n2205), .A2(n2380), .A3(n2028), .ZN(n2602) );
  INV_X1 U2477 ( .A(n2247), .ZN(n2245) );
  INV_X1 U2478 ( .A(n2274), .ZN(n2246) );
  INV_X1 U2479 ( .A(n3112), .ZN(n3117) );
  INV_X1 U2480 ( .A(n2079), .ZN(n2077) );
  NAND2_X1 U2481 ( .A1(n3970), .A2(n2897), .ZN(n3952) );
  OAI21_X1 U2482 ( .B1(n2843), .B2(n2179), .A(n2847), .ZN(n2178) );
  NAND2_X1 U2483 ( .A1(n3175), .A2(n3644), .ZN(n3141) );
  AND2_X1 U2484 ( .A1(n4341), .A2(n3641), .ZN(n2985) );
  INV_X1 U2485 ( .A(n3708), .ZN(n2871) );
  OR2_X1 U2486 ( .A1(n3524), .A2(n4122), .ZN(n2154) );
  INV_X1 U2487 ( .A(n2965), .ZN(n2911) );
  INV_X1 U2488 ( .A(IR_REG_6__SCAN_IN), .ZN(n2402) );
  AND2_X1 U2489 ( .A1(n2236), .A2(n2103), .ZN(n2102) );
  AND2_X1 U2490 ( .A1(n2042), .A2(n2423), .ZN(n2236) );
  AND2_X1 U2491 ( .A1(n2799), .A2(n3125), .ZN(n2741) );
  NAND2_X1 U2492 ( .A1(n3367), .A2(n3368), .ZN(n2133) );
  NAND2_X1 U2493 ( .A1(n3468), .A2(n2698), .ZN(n3532) );
  AOI21_X1 U2494 ( .B1(n2651), .B2(n2123), .A(n2121), .ZN(n2120) );
  NAND2_X1 U2495 ( .A1(n3084), .A2(n3083), .ZN(n3082) );
  AOI21_X1 U2496 ( .B1(n2130), .B2(n2128), .A(n2127), .ZN(n2126) );
  INV_X1 U2497 ( .A(n2130), .ZN(n2129) );
  INV_X1 U2498 ( .A(n2134), .ZN(n2128) );
  NAND2_X1 U2499 ( .A1(n2235), .A2(n2233), .ZN(n3566) );
  NAND2_X1 U2500 ( .A1(n2651), .A2(n2256), .ZN(n2235) );
  NAND2_X1 U2501 ( .A1(n3622), .A2(DATAI_22_), .ZN(n4020) );
  OR2_X1 U2502 ( .A1(n2483), .A2(n3371), .ZN(n2496) );
  XNOR2_X1 U2503 ( .A(n2337), .B(n2753), .ZN(n2342) );
  OAI21_X1 U2504 ( .B1(n2822), .B2(n2321), .A(n2336), .ZN(n2337) );
  OR2_X1 U2505 ( .A1(n3102), .A2(n2752), .ZN(n2336) );
  INV_X1 U2506 ( .A(n3593), .ZN(n3579) );
  INV_X1 U2507 ( .A(n3641), .ZN(n3757) );
  NAND2_X1 U2508 ( .A1(n2362), .A2(n2361), .ZN(n2365) );
  NAND2_X1 U2509 ( .A1(n3804), .A2(n2033), .ZN(n2099) );
  XNOR2_X1 U2510 ( .A(n2166), .B(n2165), .ZN(n3010) );
  INV_X1 U2511 ( .A(n2352), .ZN(n2225) );
  OAI22_X1 U2512 ( .A1(n2155), .A2(n2158), .B1(n2156), .B2(n2029), .ZN(n3013)
         );
  OR2_X1 U2513 ( .A1(n3818), .A2(n2029), .ZN(n2155) );
  NAND2_X1 U2514 ( .A1(n3036), .A2(n2072), .ZN(n3038) );
  NAND2_X1 U2515 ( .A1(n2073), .A2(n2162), .ZN(n2072) );
  INV_X1 U2516 ( .A(n2074), .ZN(n2073) );
  OAI21_X1 U2517 ( .B1(n2214), .B2(n4381), .A(n2213), .ZN(n4390) );
  NAND2_X1 U2518 ( .A1(n2215), .A2(REG1_REG_12__SCAN_IN), .ZN(n2214) );
  NAND2_X1 U2519 ( .A1(n3848), .A2(n2215), .ZN(n2213) );
  NOR2_X1 U2520 ( .A1(n4381), .A2(n4382), .ZN(n4380) );
  NAND2_X1 U2521 ( .A1(n4418), .A2(n3863), .ZN(n4431) );
  INV_X1 U2522 ( .A(n2168), .ZN(n3862) );
  NAND2_X1 U2523 ( .A1(n2220), .A2(n3873), .ZN(n2219) );
  NOR2_X1 U2524 ( .A1(n3879), .A2(n2058), .ZN(n2095) );
  AND2_X1 U2525 ( .A1(n3003), .A2(n3002), .ZN(n3044) );
  INV_X1 U2526 ( .A(n2867), .ZN(n2172) );
  NAND2_X1 U2527 ( .A1(n3622), .A2(DATAI_27_), .ZN(n3922) );
  INV_X1 U2528 ( .A(n2195), .ZN(n2194) );
  AOI21_X1 U2529 ( .B1(n2195), .B2(n2193), .A(n2037), .ZN(n2192) );
  AOI21_X1 U2530 ( .B1(n4011), .B2(n2860), .A(n2035), .ZN(n2195) );
  AND2_X1 U2531 ( .A1(n2711), .A2(n2710), .ZN(n3973) );
  INV_X1 U2532 ( .A(n3957), .ZN(n3994) );
  INV_X1 U2533 ( .A(n4020), .ZN(n4012) );
  AND4_X1 U2534 ( .A1(n2676), .A2(n2675), .A3(n2674), .A4(n2673), .ZN(n4016)
         );
  NOR2_X1 U2535 ( .A1(n2658), .A2(n2657), .ZN(n2669) );
  NAND2_X1 U2536 ( .A1(n3622), .A2(DATAI_21_), .ZN(n4028) );
  NAND2_X1 U2537 ( .A1(n4046), .A2(n3615), .ZN(n2892) );
  OR2_X1 U2538 ( .A1(n3733), .A2(n3732), .ZN(n4070) );
  INV_X1 U2539 ( .A(n2182), .ZN(n4086) );
  NOR2_X1 U2540 ( .A1(n2184), .A2(n2852), .ZN(n2183) );
  NAND2_X1 U2541 ( .A1(n4126), .A2(n3683), .ZN(n4104) );
  AND4_X1 U2542 ( .A1(n2535), .A2(n2534), .A3(n2533), .A4(n2532), .ZN(n4143)
         );
  OAI21_X1 U2543 ( .B1(n2887), .B2(n4152), .A(n2059), .ZN(n4136) );
  AND2_X1 U2544 ( .A1(n2060), .A2(n3610), .ZN(n2059) );
  OR2_X1 U2545 ( .A1(n3676), .A2(n4152), .ZN(n2060) );
  NAND2_X1 U2546 ( .A1(n2887), .A2(n3676), .ZN(n4153) );
  AND2_X1 U2547 ( .A1(n2513), .A2(REG3_REG_13__SCAN_IN), .ZN(n2530) );
  OR2_X1 U2548 ( .A1(n3736), .A2(n3735), .ZN(n4180) );
  AND4_X1 U2549 ( .A1(n2519), .A2(n2518), .A3(n2517), .A4(n2516), .ZN(n3461)
         );
  AND2_X1 U2550 ( .A1(n3399), .A2(n3401), .ZN(n3710) );
  INV_X1 U2551 ( .A(n4184), .ZN(n4159) );
  OAI21_X1 U2552 ( .B1(n3321), .B2(n3320), .A(n3660), .ZN(n3377) );
  NOR2_X1 U2553 ( .A1(n2440), .A2(n3359), .ZN(n2466) );
  OR2_X1 U2554 ( .A1(n2411), .A2(n2410), .ZN(n2425) );
  INV_X1 U2555 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2424) );
  INV_X1 U2556 ( .A(n3292), .ZN(n3231) );
  NAND2_X1 U2557 ( .A1(n2876), .A2(n3655), .ZN(n3226) );
  INV_X1 U2558 ( .A(n4450), .ZN(n4154) );
  NOR2_X1 U2559 ( .A1(n2988), .A2(n2908), .ZN(n3109) );
  INV_X1 U2560 ( .A(n3196), .ZN(n3709) );
  OAI21_X1 U2561 ( .B1(n3113), .B2(n3730), .A(n3643), .ZN(n3176) );
  NAND2_X1 U2562 ( .A1(n3176), .A2(n3708), .ZN(n3175) );
  AND4_X1 U2563 ( .A1(n2351), .A2(n2350), .A3(n2349), .A4(n2348), .ZN(n3178)
         );
  NAND2_X1 U2564 ( .A1(n3907), .A2(n3908), .ZN(n2143) );
  AND2_X1 U2565 ( .A1(n4452), .A2(n3759), .ZN(n4450) );
  AOI21_X1 U2566 ( .B1(n3893), .B2(n3892), .A(n3891), .ZN(n3894) );
  NAND2_X1 U2567 ( .A1(n2902), .A2(n3635), .ZN(n4281) );
  NAND2_X1 U2568 ( .A1(n3942), .A2(n3922), .ZN(n3921) );
  NOR2_X1 U2569 ( .A1(n3960), .A2(n3936), .ZN(n3942) );
  NAND2_X1 U2570 ( .A1(n2153), .A2(n3961), .ZN(n3960) );
  NAND2_X1 U2571 ( .A1(n3622), .A2(DATAI_24_), .ZN(n3979) );
  INV_X1 U2572 ( .A(n3473), .ZN(n4000) );
  AND2_X1 U2573 ( .A1(n4035), .A2(n4020), .ZN(n4237) );
  NOR2_X1 U2574 ( .A1(n4056), .A2(n4034), .ZN(n4035) );
  AND2_X1 U2575 ( .A1(n3622), .A2(DATAI_20_), .ZN(n4054) );
  OR2_X1 U2576 ( .A1(n4079), .A2(n4054), .ZN(n4056) );
  NOR3_X1 U2577 ( .A1(n4121), .A2(n4094), .A3(n2154), .ZN(n4077) );
  NAND2_X1 U2578 ( .A1(n4077), .A2(n4076), .ZN(n4079) );
  NOR2_X1 U2579 ( .A1(n4121), .A2(n2154), .ZN(n4110) );
  NOR2_X1 U2580 ( .A1(n4121), .A2(n4122), .ZN(n2918) );
  NAND2_X1 U2581 ( .A1(n3430), .A2(n2050), .ZN(n4190) );
  NAND2_X1 U2582 ( .A1(n3430), .A2(n2152), .ZN(n4189) );
  NAND2_X1 U2583 ( .A1(n3430), .A2(n3429), .ZN(n3428) );
  AND2_X1 U2584 ( .A1(n3249), .A2(n2022), .ZN(n3383) );
  AND2_X1 U2585 ( .A1(n3383), .A2(n3382), .ZN(n3430) );
  INV_X1 U2586 ( .A(n3350), .ZN(n3382) );
  NAND2_X1 U2587 ( .A1(n3249), .A2(n2151), .ZN(n3280) );
  NAND2_X1 U2588 ( .A1(n3249), .A2(n2018), .ZN(n3327) );
  NAND2_X1 U2589 ( .A1(n4455), .A2(n4480), .ZN(n4513) );
  INV_X1 U2590 ( .A(n3308), .ZN(n3248) );
  AND2_X1 U2591 ( .A1(n3249), .A2(n3248), .ZN(n3251) );
  INV_X1 U2592 ( .A(n3108), .ZN(n2923) );
  INV_X1 U2593 ( .A(n4453), .ZN(n4282) );
  INV_X1 U2594 ( .A(n4513), .ZN(n4496) );
  NAND2_X1 U2595 ( .A1(n2149), .A2(IR_REG_31__SCAN_IN), .ZN(n2989) );
  INV_X1 U2596 ( .A(IR_REG_20__SCAN_IN), .ZN(n2291) );
  NAND2_X1 U2597 ( .A1(n2314), .A2(IR_REG_31__SCAN_IN), .ZN(n2292) );
  INV_X1 U2598 ( .A(IR_REG_17__SCAN_IN), .ZN(n2268) );
  INV_X1 U2599 ( .A(n2242), .ZN(n2241) );
  NOR2_X1 U2600 ( .A1(n2536), .A2(n2242), .ZN(n2585) );
  AND2_X1 U2601 ( .A1(n2380), .A2(n2265), .ZN(n2520) );
  AND4_X1 U2602 ( .A1(n2430), .A2(n2429), .A3(n2428), .A4(n2427), .ZN(n3360)
         );
  NAND2_X1 U2603 ( .A1(n3314), .A2(n2110), .ZN(n2105) );
  AND2_X1 U2604 ( .A1(n3622), .A2(DATAI_23_), .ZN(n3473) );
  OAI21_X1 U2605 ( .B1(n3314), .B2(n2108), .A(n2106), .ZN(n2237) );
  INV_X1 U2606 ( .A(n4028), .ZN(n4034) );
  INV_X1 U2607 ( .A(n4122), .ZN(n4128) );
  NAND2_X1 U2608 ( .A1(n2229), .A2(n2576), .ZN(n3521) );
  INV_X1 U2609 ( .A(n3979), .ZN(n3539) );
  NAND2_X1 U2610 ( .A1(n2113), .A2(n2360), .ZN(n3156) );
  AND4_X1 U2611 ( .A1(n2501), .A2(n2500), .A3(n2499), .A4(n2498), .ZN(n4185)
         );
  NOR2_X2 U2612 ( .A1(n2792), .A2(n2793), .ZN(n3563) );
  NAND2_X1 U2613 ( .A1(n2235), .A2(n3490), .ZN(n3568) );
  AND2_X1 U2614 ( .A1(n2115), .A2(n2227), .ZN(n2114) );
  NOR2_X1 U2615 ( .A1(n2230), .A2(n2228), .ZN(n2227) );
  AND4_X1 U2616 ( .A1(n2563), .A2(n2562), .A3(n2561), .A4(n2560), .ZN(n3594)
         );
  NOR2_X1 U2617 ( .A1(n2321), .A2(n2801), .ZN(n3766) );
  INV_X1 U2618 ( .A(n3973), .ZN(n3535) );
  INV_X1 U2619 ( .A(n4016), .ZN(n3975) );
  INV_X1 U2620 ( .A(n4106), .ZN(n4073) );
  INV_X1 U2621 ( .A(n3594), .ZN(n4140) );
  INV_X1 U2622 ( .A(n4143), .ZN(n4182) );
  INV_X1 U2623 ( .A(n3461), .ZN(n4158) );
  INV_X1 U2624 ( .A(n4185), .ZN(n3775) );
  NAND2_X1 U2625 ( .A1(n2330), .A2(n3206), .ZN(n2209) );
  INV_X1 U2626 ( .A(n3178), .ZN(n3213) );
  OR2_X1 U2627 ( .A1(n2304), .A2(n2967), .ZN(n3783) );
  NAND2_X1 U2628 ( .A1(n2996), .A2(n2997), .ZN(n3812) );
  XNOR2_X1 U2629 ( .A(n2099), .B(n2165), .ZN(n3017) );
  OAI21_X1 U2630 ( .B1(n3818), .B2(n2158), .A(n2156), .ZN(n2159) );
  AOI21_X1 U2631 ( .B1(n3818), .B2(REG2_REG_4__SCAN_IN), .A(n2158), .ZN(n3053)
         );
  AOI21_X1 U2632 ( .B1(n3817), .B2(REG1_REG_4__SCAN_IN), .A(n2081), .ZN(n3056)
         );
  XNOR2_X1 U2633 ( .A(n3013), .B(n4345), .ZN(n3074) );
  AOI22_X1 U2634 ( .A1(n3075), .A2(REG1_REG_6__SCAN_IN), .B1(n4345), .B2(n3021), .ZN(n3064) );
  XNOR2_X1 U2635 ( .A(n2074), .B(n2162), .ZN(n3022) );
  NAND2_X1 U2636 ( .A1(n3022), .A2(REG1_REG_8__SCAN_IN), .ZN(n3036) );
  OAI22_X1 U2637 ( .A1(n3031), .A2(n3030), .B1(n3037), .B2(n2161), .ZN(n4365)
         );
  INV_X1 U2638 ( .A(n2163), .ZN(n2161) );
  INV_X1 U2639 ( .A(n2210), .ZN(n4359) );
  INV_X1 U2640 ( .A(n3038), .ZN(n4361) );
  NAND2_X1 U2641 ( .A1(n3832), .A2(n3833), .ZN(n4375) );
  NOR2_X1 U2642 ( .A1(n3844), .A2(n3845), .ZN(n4371) );
  NAND2_X1 U2643 ( .A1(n4386), .A2(n3836), .ZN(n4397) );
  INV_X1 U2644 ( .A(n2090), .ZN(n4402) );
  INV_X1 U2645 ( .A(n2089), .ZN(n3853) );
  NAND2_X1 U2646 ( .A1(n4421), .A2(n3871), .ZN(n4434) );
  AOI21_X1 U2647 ( .B1(n2095), .B2(n3873), .A(n2026), .ZN(n2094) );
  NAND2_X1 U2648 ( .A1(n2097), .A2(n3879), .ZN(n2096) );
  INV_X1 U2649 ( .A(n3873), .ZN(n2097) );
  NOR2_X1 U2650 ( .A1(n2140), .A2(n4208), .ZN(n4216) );
  INV_X1 U2651 ( .A(n2143), .ZN(n2140) );
  OR2_X1 U2652 ( .A1(n2734), .A2(n2745), .ZN(n3924) );
  NAND2_X1 U2653 ( .A1(n4008), .A2(n2860), .ZN(n3987) );
  OAI21_X1 U2654 ( .B1(n4135), .B2(n2187), .A(n2185), .ZN(n4103) );
  AND2_X1 U2655 ( .A1(n2190), .A2(n2191), .ZN(n4120) );
  NAND2_X1 U2656 ( .A1(n2190), .A2(n2188), .ZN(n4118) );
  NAND2_X1 U2657 ( .A1(n3418), .A2(n2845), .ZN(n3414) );
  NAND2_X1 U2658 ( .A1(n2198), .A2(n2201), .ZN(n3381) );
  OR2_X1 U2659 ( .A1(n2988), .A2(n2912), .ZN(n4193) );
  NAND2_X1 U2660 ( .A1(n2135), .A2(n3150), .ZN(n4485) );
  INV_X1 U2661 ( .A(n3220), .ZN(n2135) );
  AND2_X1 U2662 ( .A1(n3730), .A2(n3729), .ZN(n4456) );
  INV_X1 U2663 ( .A(n4193), .ZN(n4459) );
  INV_X2 U2664 ( .A(n4690), .ZN(n4692) );
  NAND2_X1 U2665 ( .A1(n2966), .A2(n2965), .ZN(n4464) );
  NAND2_X1 U2666 ( .A1(n2277), .A2(n2069), .ZN(n2068) );
  XNOR2_X1 U2667 ( .A(n2804), .B(n2277), .ZN(n4351) );
  OR2_X1 U2668 ( .A1(n2297), .A2(n2601), .ZN(n2286) );
  XNOR2_X1 U2669 ( .A(n2289), .B(IR_REG_25__SCAN_IN), .ZN(n4339) );
  NAND2_X1 U2670 ( .A1(n2287), .A2(IR_REG_31__SCAN_IN), .ZN(n2288) );
  NAND2_X1 U2671 ( .A1(n2780), .A2(n2779), .ZN(n2287) );
  AND2_X1 U2672 ( .A1(n2987), .A2(STATE_REG_SCAN_IN), .ZN(n4466) );
  INV_X1 U2673 ( .A(n2795), .ZN(n3759) );
  INV_X1 U2674 ( .A(n4451), .ZN(n4342) );
  INV_X1 U2675 ( .A(n3849), .ZN(n4473) );
  XNOR2_X1 U2676 ( .A(n2369), .B(IR_REG_4__SCAN_IN), .ZN(n4347) );
  NAND2_X1 U2677 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2071)
         );
  NAND2_X1 U2678 ( .A1(n3843), .A2(n2086), .ZN(n3040) );
  INV_X1 U2679 ( .A(n2216), .ZN(n3875) );
  OAI211_X1 U2680 ( .C1(n2220), .C2(n2093), .A(n4437), .B(n2091), .ZN(n2098)
         );
  NAND2_X1 U2681 ( .A1(n2094), .A2(n2096), .ZN(n2093) );
  AOI22_X1 U2682 ( .A1(n4356), .A2(n4444), .B1(REG2_REG_30__SCAN_IN), .B2(
        n2017), .ZN(n4357) );
  INV_X1 U2683 ( .A(n2137), .ZN(n2136) );
  OR2_X1 U2684 ( .A1(n3447), .A2(n4278), .ZN(n2921) );
  NAND2_X1 U2685 ( .A1(n2062), .A2(n2055), .ZN(U3515) );
  INV_X1 U2686 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2061) );
  INV_X1 U2687 ( .A(IR_REG_31__SCAN_IN), .ZN(n2601) );
  AND2_X1 U2688 ( .A1(n2151), .A2(n3302), .ZN(n2018) );
  AND2_X1 U2689 ( .A1(n4214), .A2(n4513), .ZN(n2019) );
  INV_X2 U2690 ( .A(n2755), .ZN(n2307) );
  NAND2_X1 U2691 ( .A1(n2225), .A2(n2250), .ZN(n2381) );
  OR2_X1 U2692 ( .A1(n2536), .A2(IR_REG_14__SCAN_IN), .ZN(n2020) );
  NOR2_X1 U2693 ( .A1(n2834), .A2(n3240), .ZN(n2021) );
  INV_X1 U2694 ( .A(n2846), .ZN(n2181) );
  AND2_X1 U2695 ( .A1(n2018), .A2(n2150), .ZN(n2022) );
  INV_X1 U2696 ( .A(n3555), .ZN(n2240) );
  OR2_X1 U2697 ( .A1(n4478), .A2(n4528), .ZN(n2023) );
  AND2_X1 U2698 ( .A1(n2232), .A2(n2117), .ZN(n2024) );
  AND2_X1 U2699 ( .A1(n2169), .A2(n2023), .ZN(n2025) );
  AND2_X1 U2700 ( .A1(n3879), .A2(n2058), .ZN(n2026) );
  AND3_X1 U2701 ( .A1(n2250), .A2(n2335), .A3(n2224), .ZN(n2380) );
  AND2_X1 U2702 ( .A1(n2962), .A2(n4337), .ZN(n2330) );
  AND2_X1 U2703 ( .A1(n4129), .A2(n4112), .ZN(n2027) );
  AND2_X1 U2704 ( .A1(n2241), .A2(n2268), .ZN(n2028) );
  XNOR2_X1 U2705 ( .A(n2280), .B(IR_REG_29__SCAN_IN), .ZN(n2962) );
  AND4_X1 U2706 ( .A1(n2416), .A2(n2415), .A3(n2414), .A4(n2413), .ZN(n2833)
         );
  AND2_X1 U2707 ( .A1(n4346), .A2(REG2_REG_5__SCAN_IN), .ZN(n2029) );
  AND4_X1 U2708 ( .A1(n2334), .A2(n2333), .A3(n2332), .A4(n2331), .ZN(n2822)
         );
  NAND2_X1 U2709 ( .A1(n2116), .A2(n2114), .ZN(n3476) );
  INV_X1 U2710 ( .A(IR_REG_2__SCAN_IN), .ZN(n4671) );
  NAND2_X1 U2711 ( .A1(n4337), .A2(n2282), .ZN(n2442) );
  INV_X2 U2712 ( .A(n2442), .ZN(n2672) );
  OR2_X1 U2713 ( .A1(n2293), .A2(IR_REG_21__SCAN_IN), .ZN(n2030) );
  INV_X1 U2714 ( .A(n3904), .ZN(n2173) );
  INV_X1 U2715 ( .A(n3302), .ZN(n3279) );
  OR2_X1 U2716 ( .A1(n3850), .A2(n4472), .ZN(n2031) );
  NAND2_X1 U2717 ( .A1(n3288), .A2(n3308), .ZN(n2032) );
  OR2_X1 U2718 ( .A1(n2998), .A2(n2994), .ZN(n2033) );
  OR2_X1 U2719 ( .A1(n2998), .A2(n2999), .ZN(n2034) );
  NOR2_X1 U2720 ( .A1(n3975), .A2(n3473), .ZN(n2035) );
  NAND2_X1 U2721 ( .A1(n2335), .A2(n4671), .ZN(n2352) );
  NAND2_X1 U2722 ( .A1(n4346), .A2(REG1_REG_5__SCAN_IN), .ZN(n2082) );
  INV_X1 U2723 ( .A(n4208), .ZN(n2144) );
  NOR2_X1 U2724 ( .A1(n3907), .A2(n3908), .ZN(n4208) );
  OR3_X1 U2725 ( .A1(n2293), .A2(n2247), .A3(n2274), .ZN(n2036) );
  AND2_X1 U2726 ( .A1(n3975), .A2(n3473), .ZN(n2037) );
  AND2_X1 U2727 ( .A1(n2099), .A2(n4348), .ZN(n2038) );
  AND2_X1 U2728 ( .A1(n2166), .A2(n4348), .ZN(n2039) );
  INV_X1 U2729 ( .A(n2845), .ZN(n2179) );
  NOR2_X1 U2730 ( .A1(n3594), .A2(n4128), .ZN(n2040) );
  OR2_X1 U2731 ( .A1(n3776), .A2(n3350), .ZN(n2041) );
  NOR2_X1 U2732 ( .A1(n3354), .A2(n2465), .ZN(n2042) );
  AND2_X1 U2733 ( .A1(n2360), .A2(n2374), .ZN(n2043) );
  AND2_X1 U2734 ( .A1(n2041), .A2(n2201), .ZN(n2044) );
  NAND2_X1 U2735 ( .A1(n4282), .A2(n2738), .ZN(n2045) );
  INV_X1 U2736 ( .A(n2084), .ZN(n2081) );
  NAND2_X1 U2737 ( .A1(n3019), .A2(n4347), .ZN(n2084) );
  OR2_X1 U2738 ( .A1(n2187), .A2(n2027), .ZN(n2046) );
  INV_X1 U2739 ( .A(n3037), .ZN(n2162) );
  INV_X1 U2740 ( .A(n4119), .ZN(n2189) );
  NAND2_X1 U2741 ( .A1(n2237), .A2(n2423), .ZN(n3296) );
  INV_X1 U2742 ( .A(n4094), .ZN(n3582) );
  AND2_X1 U2743 ( .A1(n3772), .A2(n3936), .ZN(n2047) );
  INV_X1 U2744 ( .A(n3322), .ZN(n2150) );
  OAI21_X1 U2745 ( .B1(n3370), .B2(n2129), .A(n2126), .ZN(n3553) );
  INV_X1 U2746 ( .A(n2234), .ZN(n2233) );
  NAND2_X1 U2747 ( .A1(n2668), .A2(n3490), .ZN(n2234) );
  OR2_X1 U2748 ( .A1(n4344), .A2(REG1_REG_7__SCAN_IN), .ZN(n2048) );
  NAND2_X1 U2749 ( .A1(n2132), .A2(n2133), .ZN(n3390) );
  NAND2_X1 U2750 ( .A1(n2529), .A2(n2528), .ZN(n3456) );
  NAND2_X1 U2751 ( .A1(n2205), .A2(n2380), .ZN(n2536) );
  NOR2_X1 U2752 ( .A1(n4380), .A2(n3848), .ZN(n2049) );
  AND2_X1 U2753 ( .A1(n2152), .A2(n4191), .ZN(n2050) );
  INV_X1 U2754 ( .A(n2153), .ZN(n3978) );
  NOR2_X1 U2755 ( .A1(n3999), .A2(n3539), .ZN(n2153) );
  AND2_X1 U2756 ( .A1(n2559), .A2(n2119), .ZN(n2051) );
  AND2_X1 U2757 ( .A1(n3991), .A2(n2893), .ZN(n4011) );
  INV_X1 U2758 ( .A(n4011), .ZN(n2196) );
  INV_X1 U2759 ( .A(IR_REG_14__SCAN_IN), .ZN(n2267) );
  AND2_X1 U2760 ( .A1(n3917), .A2(n3903), .ZN(n2052) );
  OR2_X1 U2761 ( .A1(n3066), .A2(n4598), .ZN(n2053) );
  OR2_X1 U2762 ( .A1(n2257), .A2(n2047), .ZN(n2054) );
  INV_X1 U2763 ( .A(n3846), .ZN(n2167) );
  NAND2_X1 U2764 ( .A1(n2087), .A2(n3830), .ZN(n3843) );
  INV_X2 U2765 ( .A(n4530), .ZN(n4533) );
  OR2_X1 U2766 ( .A1(n2924), .A2(n3108), .ZN(n4530) );
  NAND2_X1 U2767 ( .A1(n2105), .A2(n2109), .ZN(n3285) );
  INV_X1 U2768 ( .A(n3683), .ZN(n2066) );
  INV_X1 U2769 ( .A(n3391), .ZN(n2127) );
  NAND2_X1 U2770 ( .A1(n2104), .A2(n2102), .ZN(n3341) );
  NAND2_X1 U2771 ( .A1(n2844), .A2(n2843), .ZN(n3418) );
  OR2_X1 U2772 ( .A1(n4692), .A2(n2061), .ZN(n2055) );
  NOR2_X1 U2773 ( .A1(n4533), .A2(n4557), .ZN(n2056) );
  INV_X1 U2774 ( .A(n2850), .ZN(n2191) );
  INV_X1 U2775 ( .A(n4502), .ZN(n2101) );
  AND4_X1 U2776 ( .A1(n2320), .A2(n2319), .A3(n2318), .A4(n2317), .ZN(n3087)
         );
  INV_X1 U2777 ( .A(n4437), .ZN(n4401) );
  AND2_X1 U2778 ( .A1(n3044), .A2(n3794), .ZN(n4437) );
  AND2_X1 U2779 ( .A1(n2094), .A2(n2092), .ZN(n2057) );
  AND2_X1 U2780 ( .A1(n2712), .A2(DATAI_25_), .ZN(n3508) );
  INV_X1 U2781 ( .A(n3830), .ZN(n2169) );
  INV_X1 U2782 ( .A(n3872), .ZN(n4468) );
  AND2_X1 U2783 ( .A1(n3881), .A2(REG1_REG_18__SCAN_IN), .ZN(n2058) );
  INV_X1 U2784 ( .A(DATAI_0_), .ZN(n2145) );
  INV_X1 U2785 ( .A(DATAI_1_), .ZN(n2147) );
  INV_X1 U2786 ( .A(IR_REG_29__SCAN_IN), .ZN(n2069) );
  INV_X1 U2787 ( .A(IR_REG_0__SCAN_IN), .ZN(n2146) );
  AND2_X1 U2788 ( .A1(n2368), .A2(n2355), .ZN(n4348) );
  INV_X1 U2789 ( .A(n4348), .ZN(n2165) );
  INV_X1 U2790 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2080) );
  INV_X1 U2791 ( .A(n2803), .ZN(n2067) );
  NAND2_X1 U2792 ( .A1(n2067), .A2(n2277), .ZN(n2279) );
  NOR2_X1 U2793 ( .A1(n2803), .A2(n2068), .ZN(n3444) );
  NAND3_X1 U2794 ( .A1(n4670), .A2(n2552), .A3(n2267), .ZN(n2242) );
  MUX2_X1 U2795 ( .A(REG1_REG_1__SCAN_IN), .B(n2990), .S(n4349), .Z(n2070) );
  XNOR2_X2 U2796 ( .A(n2071), .B(IR_REG_1__SCAN_IN), .ZN(n4349) );
  NAND2_X1 U2797 ( .A1(n2076), .A2(n2075), .ZN(n3020) );
  NAND3_X1 U2798 ( .A1(n2078), .A2(n2082), .A3(n2084), .ZN(n2076) );
  OAI21_X1 U2799 ( .B1(n3817), .B2(n2081), .A(n2079), .ZN(n2083) );
  INV_X1 U2800 ( .A(n3817), .ZN(n2078) );
  INV_X1 U2801 ( .A(n2083), .ZN(n3054) );
  NAND2_X1 U2802 ( .A1(n2210), .A2(n2023), .ZN(n2087) );
  NAND2_X1 U2803 ( .A1(n2098), .A2(n3889), .ZN(U3259) );
  NAND2_X4 U2804 ( .A1(n2101), .A2(n2738), .ZN(n2755) );
  NAND2_X2 U2805 ( .A1(n2304), .A2(n3125), .ZN(n2752) );
  NAND2_X2 U2806 ( .A1(n4340), .A2(n2100), .ZN(n2304) );
  NAND2_X1 U2807 ( .A1(n3314), .A2(n2106), .ZN(n2104) );
  NAND2_X1 U2808 ( .A1(n2113), .A2(n2043), .ZN(n3157) );
  NAND2_X1 U2809 ( .A1(n2558), .A2(n2024), .ZN(n2116) );
  OAI21_X1 U2810 ( .B1(n2651), .B2(n2234), .A(n2123), .ZN(n3468) );
  INV_X1 U2811 ( .A(n2120), .ZN(n2695) );
  NAND2_X1 U2812 ( .A1(n3370), .A2(n2134), .ZN(n2132) );
  INV_X1 U2813 ( .A(n3553), .ZN(n2527) );
  AND2_X2 U2814 ( .A1(n3184), .A2(n3149), .ZN(n3220) );
  OAI21_X1 U2815 ( .B1(n2141), .B2(n4530), .A(n2139), .ZN(U3547) );
  MUX2_X1 U2816 ( .A(n2146), .B(n2145), .S(n2370), .Z(n4453) );
  MUX2_X1 U2817 ( .A(n2148), .B(n2147), .S(n2370), .Z(n3112) );
  NAND2_X1 U2818 ( .A1(n2297), .A2(n2296), .ZN(n2149) );
  AND2_X1 U2819 ( .A1(n2271), .A2(n2203), .ZN(n2297) );
  NAND2_X1 U2820 ( .A1(n2695), .A2(n2694), .ZN(n3531) );
  NAND2_X1 U2821 ( .A1(n3163), .A2(n2392), .ZN(n3314) );
  NAND2_X1 U2822 ( .A1(n3531), .A2(n2702), .ZN(n3504) );
  AOI21_X1 U2823 ( .B1(n2943), .B2(n2940), .A(n2939), .ZN(n2930) );
  NAND2_X1 U2824 ( .A1(n3064), .A2(n2053), .ZN(n2212) );
  NAND2_X1 U2825 ( .A1(n2223), .A2(n3457), .ZN(n2558) );
  NAND2_X1 U2826 ( .A1(n2341), .A2(n2340), .ZN(n3100) );
  OAI21_X1 U2827 ( .B1(n3087), .B2(n2321), .A(n2322), .ZN(n2323) );
  INV_X1 U2828 ( .A(n2159), .ZN(n3051) );
  NAND2_X1 U2829 ( .A1(n2868), .A2(n2867), .ZN(n3905) );
  OAI21_X1 U2830 ( .B1(n2868), .B2(n2173), .A(n2171), .ZN(n2175) );
  AOI21_X1 U2831 ( .B1(n3904), .B2(n2172), .A(n2052), .ZN(n2171) );
  OAI22_X2 U2832 ( .A1(n2844), .A2(n2176), .B1(n2177), .B2(n2846), .ZN(n4174)
         );
  OAI21_X1 U2833 ( .B1(n4135), .B2(n2046), .A(n2183), .ZN(n2182) );
  OAI21_X1 U2834 ( .B1(n4007), .B2(n2194), .A(n2192), .ZN(n3968) );
  INV_X1 U2835 ( .A(n4007), .ZN(n2197) );
  NAND2_X1 U2836 ( .A1(n2198), .A2(n2044), .ZN(n2842) );
  NAND2_X1 U2837 ( .A1(n2839), .A2(n2838), .ZN(n3326) );
  INV_X1 U2838 ( .A(n2838), .ZN(n2200) );
  OR2_X1 U2839 ( .A1(n3777), .A2(n3322), .ZN(n2201) );
  OAI21_X1 U2840 ( .B1(n2864), .B2(n2054), .A(n2865), .ZN(n3918) );
  NOR2_X1 U2841 ( .A1(n2864), .A2(n2257), .ZN(n3929) );
  INV_X1 U2842 ( .A(n3918), .ZN(n2866) );
  NAND2_X1 U2843 ( .A1(n2271), .A2(n2202), .ZN(n2803) );
  NAND2_X1 U2844 ( .A1(n2271), .A2(n2270), .ZN(n2293) );
  NAND4_X1 U2845 ( .A1(n2028), .A2(n2205), .A3(n2380), .A4(n2269), .ZN(n2290)
         );
  NAND3_X1 U2846 ( .A1(n2209), .A2(n2208), .A3(n2207), .ZN(n2206) );
  INV_X1 U2847 ( .A(n4391), .ZN(n2215) );
  XNOR2_X2 U2848 ( .A(n2222), .B(n4671), .ZN(n3807) );
  NAND3_X1 U2849 ( .A1(n2529), .A2(n2528), .A3(n2541), .ZN(n2223) );
  NAND3_X1 U2850 ( .A1(n2575), .A2(n3596), .A3(n3513), .ZN(n2229) );
  NAND2_X1 U2851 ( .A1(n2238), .A2(n2239), .ZN(n2526) );
  NAND2_X1 U2852 ( .A1(n3390), .A2(n3391), .ZN(n2238) );
  NAND3_X1 U2853 ( .A1(n2246), .A2(n2275), .A3(n2245), .ZN(n2244) );
  NAND2_X1 U2854 ( .A1(n4237), .A2(n4000), .ZN(n3999) );
  NAND2_X1 U2855 ( .A1(n3117), .A2(n2738), .ZN(n2322) );
  NAND2_X1 U2856 ( .A1(n3087), .A2(n3117), .ZN(n3643) );
  CLKBUF_X1 U2857 ( .A(n2870), .Z(n3113) );
  NAND2_X1 U2858 ( .A1(n3784), .A2(n2307), .ZN(n2310) );
  AND2_X1 U2859 ( .A1(n3784), .A2(n4282), .ZN(n3114) );
  XNOR2_X1 U2860 ( .A(n2780), .B(n2779), .ZN(n2987) );
  NAND2_X1 U2861 ( .A1(n2347), .A2(REG0_REG_1__SCAN_IN), .ZN(n2318) );
  NAND2_X1 U2862 ( .A1(n2279), .A2(IR_REG_31__SCAN_IN), .ZN(n2280) );
  OR2_X1 U2863 ( .A1(n3557), .A2(n3940), .ZN(n2249) );
  AND2_X1 U2864 ( .A1(n2353), .A2(n2261), .ZN(n2250) );
  NAND2_X1 U2865 ( .A1(n3590), .A2(n3936), .ZN(n2251) );
  AND2_X1 U2866 ( .A1(n2672), .A2(REG2_REG_5__SCAN_IN), .ZN(n2252) );
  AND2_X1 U2867 ( .A1(n2672), .A2(REG2_REG_6__SCAN_IN), .ZN(n2253) );
  OR2_X1 U2868 ( .A1(n3937), .A2(n3638), .ZN(n2254) );
  OR2_X1 U2869 ( .A1(n2944), .A2(n3599), .ZN(n2255) );
  NAND2_X1 U2870 ( .A1(n2652), .A2(n2653), .ZN(n2256) );
  AND2_X1 U2871 ( .A1(n3535), .A2(n3508), .ZN(n2257) );
  AND2_X1 U2872 ( .A1(n2816), .A2(n2815), .ZN(n2258) );
  NAND2_X1 U2873 ( .A1(n2828), .A2(n2874), .ZN(n2259) );
  AND4_X1 U2874 ( .A1(n2551), .A2(n2550), .A3(n2549), .A4(n2548), .ZN(n4156)
         );
  OR2_X1 U2875 ( .A1(n2442), .A2(n2281), .ZN(n2260) );
  INV_X1 U2876 ( .A(IR_REG_4__SCAN_IN), .ZN(n2261) );
  INV_X1 U2877 ( .A(IR_REG_18__SCAN_IN), .ZN(n2269) );
  INV_X1 U2878 ( .A(IR_REG_24__SCAN_IN), .ZN(n2273) );
  NAND2_X1 U2879 ( .A1(n2989), .A2(n2277), .ZN(n2299) );
  OR2_X1 U2880 ( .A1(n4031), .A2(n4054), .ZN(n2856) );
  NAND2_X1 U2881 ( .A1(n3178), .A2(n3149), .ZN(n3194) );
  INV_X1 U2882 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2410) );
  INV_X1 U2883 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2495) );
  INV_X1 U2884 ( .A(n3569), .ZN(n2668) );
  NOR2_X1 U2885 ( .A1(n2579), .A2(n2578), .ZN(n2595) );
  OAI21_X1 U2886 ( .B1(n3898), .B2(n4184), .A(n3897), .ZN(n3899) );
  INV_X1 U2887 ( .A(n3919), .ZN(n2900) );
  AND2_X1 U2888 ( .A1(n2686), .A2(REG3_REG_24__SCAN_IN), .ZN(n2703) );
  INV_X1 U2889 ( .A(n4144), .ZN(n2917) );
  OR2_X1 U2890 ( .A1(n4182), .A2(n2916), .ZN(n2849) );
  AND2_X1 U2891 ( .A1(n3649), .A2(n3646), .ZN(n3746) );
  AND2_X1 U2892 ( .A1(n3622), .A2(DATAI_28_), .ZN(n3903) );
  NAND2_X1 U2893 ( .A1(n2870), .A2(n3114), .ZN(n3116) );
  INV_X1 U2894 ( .A(n4340), .ZN(n2775) );
  OR3_X1 U2895 ( .A1(n2447), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2449) );
  INV_X1 U2896 ( .A(n3922), .ZN(n3638) );
  AND2_X1 U2897 ( .A1(n2788), .A2(n3563), .ZN(n2783) );
  OR2_X1 U2898 ( .A1(n2425), .A2(n2424), .ZN(n2440) );
  NOR2_X1 U2899 ( .A1(n2496), .A2(n2495), .ZN(n2513) );
  INV_X1 U2900 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4583) );
  INV_X1 U2901 ( .A(n3421), .ZN(n3429) );
  OR2_X1 U2902 ( .A1(n2782), .A2(n4450), .ZN(n2793) );
  INV_X1 U2903 ( .A(n3944), .ZN(n3936) );
  OR2_X1 U2904 ( .A1(n3449), .A2(n2806), .ZN(n2751) );
  INV_X1 U2905 ( .A(REG3_REG_5__SCAN_IN), .ZN(n3059) );
  INV_X1 U2906 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3359) );
  INV_X1 U2907 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3371) );
  INV_X1 U2908 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3588) );
  AND2_X1 U2909 ( .A1(n3622), .A2(n2986), .ZN(n3003) );
  INV_X1 U2910 ( .A(n3899), .ZN(n3900) );
  OAI22_X1 U2911 ( .A1(n4025), .A2(n2859), .B1(n4034), .B2(n4013), .ZN(n4007)
         );
  NOR2_X1 U2912 ( .A1(n3774), .A2(n4144), .ZN(n2850) );
  AND2_X1 U2913 ( .A1(n2882), .A2(n4185), .ZN(n2846) );
  AND2_X1 U2914 ( .A1(n3671), .A2(n3672), .ZN(n3750) );
  NAND2_X1 U2915 ( .A1(n4351), .A2(n2985), .ZN(n4155) );
  INV_X1 U2916 ( .A(n3714), .ZN(n3908) );
  INV_X1 U2917 ( .A(n2888), .ZN(n4076) );
  INV_X1 U2918 ( .A(n4191), .ZN(n4181) );
  INV_X1 U2919 ( .A(n4281), .ZN(n4161) );
  NAND2_X1 U2920 ( .A1(n2869), .A2(n4451), .ZN(n4455) );
  NAND2_X1 U2921 ( .A1(n2304), .A2(n4466), .ZN(n2988) );
  NOR2_X1 U2922 ( .A1(n2449), .A2(IR_REG_9__SCAN_IN), .ZN(n2490) );
  NAND2_X1 U2923 ( .A1(n2934), .A2(n3603), .ZN(n2935) );
  AND2_X1 U2924 ( .A1(n2669), .A2(REG3_REG_23__SCAN_IN), .ZN(n2686) );
  INV_X1 U2925 ( .A(n3581), .ZN(n3589) );
  INV_X1 U2926 ( .A(n3557), .ZN(n3603) );
  AND4_X1 U2927 ( .A1(n2600), .A2(n2599), .A3(n2598), .A4(n2597), .ZN(n4106)
         );
  AND4_X1 U2928 ( .A1(n2584), .A2(n2583), .A3(n2582), .A4(n2581), .ZN(n4129)
         );
  INV_X1 U2929 ( .A(n4155), .ZN(n4280) );
  AND2_X1 U2930 ( .A1(n4195), .A2(n4451), .ZN(n4096) );
  AND2_X1 U2931 ( .A1(n4195), .A2(n3193), .ZN(n3920) );
  NAND2_X1 U2932 ( .A1(n2778), .A2(n2777), .ZN(n3108) );
  NAND2_X1 U2933 ( .A1(n3622), .A2(DATAI_26_), .ZN(n3944) );
  AND2_X1 U2934 ( .A1(n4452), .A2(n2795), .ZN(n4502) );
  AND3_X1 U2935 ( .A1(n2791), .A2(n4342), .A3(n2795), .ZN(n4520) );
  NAND2_X1 U2936 ( .A1(n2761), .A2(n2968), .ZN(n2965) );
  INV_X1 U2937 ( .A(n3590), .ZN(n3583) );
  AND2_X1 U2938 ( .A1(n2802), .A2(n3086), .ZN(n3557) );
  INV_X1 U2939 ( .A(n3563), .ZN(n3599) );
  INV_X1 U2940 ( .A(n4129), .ZN(n3773) );
  INV_X1 U2941 ( .A(n2822), .ZN(n3782) );
  INV_X1 U2942 ( .A(n4439), .ZN(n4405) );
  INV_X1 U2943 ( .A(n4412), .ZN(n4442) );
  XNOR2_X1 U2944 ( .A(n3905), .B(n3904), .ZN(n3455) );
  INV_X1 U2945 ( .A(n3920), .ZN(n4172) );
  INV_X1 U2946 ( .A(n4444), .ZN(n4169) );
  NAND2_X1 U2947 ( .A1(n4533), .A2(n4502), .ZN(n4278) );
  OR2_X1 U2948 ( .A1(n3447), .A2(n4335), .ZN(n2927) );
  OR2_X1 U2949 ( .A1(n3430), .A2(n3384), .ZN(n3443) );
  NAND2_X1 U2950 ( .A1(n4692), .A2(n4502), .ZN(n4335) );
  OR2_X1 U2951 ( .A1(n2924), .A2(n2923), .ZN(n4690) );
  INV_X1 U2952 ( .A(n4464), .ZN(n4465) );
  AND2_X1 U2953 ( .A1(n2554), .A2(n2564), .ZN(n4343) );
  INV_X1 U2954 ( .A(n3077), .ZN(n4345) );
  INV_X2 U2955 ( .A(n3783), .ZN(U4043) );
  INV_X2 U2956 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NOR2_X1 U2957 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2264)
         );
  INV_X1 U2958 ( .A(n2290), .ZN(n2271) );
  NAND2_X1 U2959 ( .A1(n2779), .A2(n2273), .ZN(n2274) );
  INV_X1 U2960 ( .A(IR_REG_25__SCAN_IN), .ZN(n2275) );
  INV_X1 U2961 ( .A(IR_REG_28__SCAN_IN), .ZN(n2277) );
  INV_X1 U2962 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2281) );
  NAND2_X1 U2963 ( .A1(n2330), .A2(REG3_REG_0__SCAN_IN), .ZN(n2285) );
  NAND2_X1 U2964 ( .A1(n2347), .A2(REG0_REG_0__SCAN_IN), .ZN(n2284) );
  INV_X1 U2965 ( .A(n2962), .ZN(n2282) );
  NOR2_X2 U2966 ( .A1(n4337), .A2(n2282), .ZN(n2398) );
  NAND2_X1 U2967 ( .A1(n2398), .A2(REG1_REG_0__SCAN_IN), .ZN(n2283) );
  NAND2_X1 U2968 ( .A1(n2036), .A2(IR_REG_31__SCAN_IN), .ZN(n2289) );
  NAND2_X1 U2969 ( .A1(n2290), .A2(IR_REG_31__SCAN_IN), .ZN(n2312) );
  NAND2_X1 U2970 ( .A1(n2293), .A2(IR_REG_31__SCAN_IN), .ZN(n2294) );
  INV_X1 U2971 ( .A(n3125), .ZN(n2295) );
  NAND2_X1 U2972 ( .A1(n3784), .A2(n2737), .ZN(n2303) );
  INV_X1 U2973 ( .A(IR_REG_26__SCAN_IN), .ZN(n2296) );
  NAND2_X1 U2974 ( .A1(n2277), .A2(IR_REG_27__SCAN_IN), .ZN(n2301) );
  INV_X2 U2975 ( .A(n2752), .ZN(n2738) );
  AND2_X1 U2976 ( .A1(n2303), .A2(n2045), .ZN(n2315) );
  INV_X1 U2977 ( .A(REG1_REG_0__SCAN_IN), .ZN(n3787) );
  OR2_X1 U2978 ( .A1(n2304), .A2(n3787), .ZN(n2305) );
  NAND2_X1 U2979 ( .A1(n2315), .A2(n2305), .ZN(n3084) );
  NAND2_X1 U2980 ( .A1(n2030), .A2(IR_REG_31__SCAN_IN), .ZN(n2306) );
  INV_X1 U2981 ( .A(n4341), .ZN(n2791) );
  INV_X1 U2982 ( .A(n2304), .ZN(n2308) );
  AOI22_X1 U2983 ( .A1(n4282), .A2(n2737), .B1(IR_REG_0__SCAN_IN), .B2(n2308), 
        .ZN(n2309) );
  NAND2_X1 U2984 ( .A1(n2310), .A2(n2309), .ZN(n3083) );
  OR2_X1 U2985 ( .A1(n2312), .A2(n2311), .ZN(n2313) );
  NAND2_X1 U2986 ( .A1(n4341), .A2(n4451), .ZN(n2799) );
  NAND2_X1 U2987 ( .A1(n2315), .A2(n2741), .ZN(n2316) );
  NAND2_X1 U2988 ( .A1(n3082), .A2(n2316), .ZN(n3093) );
  NAND2_X1 U2989 ( .A1(n2672), .A2(REG2_REG_1__SCAN_IN), .ZN(n2320) );
  NAND2_X1 U2990 ( .A1(n2398), .A2(REG1_REG_1__SCAN_IN), .ZN(n2319) );
  NAND2_X1 U2991 ( .A1(n2330), .A2(REG3_REG_1__SCAN_IN), .ZN(n2317) );
  XNOR2_X1 U2992 ( .A(n2323), .B(n2741), .ZN(n2326) );
  OR2_X1 U2993 ( .A1(n3087), .A2(n2755), .ZN(n2325) );
  NAND2_X1 U2994 ( .A1(n3117), .A2(n2737), .ZN(n2324) );
  NAND2_X1 U2995 ( .A1(n2325), .A2(n2324), .ZN(n2327) );
  XNOR2_X1 U2996 ( .A(n2326), .B(n2327), .ZN(n3091) );
  NAND2_X1 U2997 ( .A1(n3093), .A2(n3091), .ZN(n3092) );
  INV_X1 U2998 ( .A(n2326), .ZN(n2328) );
  NAND2_X1 U2999 ( .A1(n2328), .A2(n2327), .ZN(n2329) );
  NAND2_X1 U3000 ( .A1(n3092), .A2(n2329), .ZN(n3099) );
  INV_X1 U3001 ( .A(n3099), .ZN(n2341) );
  NAND2_X1 U3002 ( .A1(n2330), .A2(REG3_REG_2__SCAN_IN), .ZN(n2334) );
  NAND2_X1 U3003 ( .A1(n2398), .A2(REG1_REG_2__SCAN_IN), .ZN(n2333) );
  NAND2_X1 U3004 ( .A1(n2016), .A2(REG2_REG_2__SCAN_IN), .ZN(n2332) );
  NAND2_X1 U3005 ( .A1(n2347), .A2(REG0_REG_2__SCAN_IN), .ZN(n2331) );
  MUX2_X1 U3006 ( .A(n3807), .B(DATAI_2_), .S(n2370), .Z(n3186) );
  INV_X1 U3007 ( .A(n3186), .ZN(n3102) );
  OR2_X1 U3008 ( .A1(n2822), .A2(n2755), .ZN(n2339) );
  NAND2_X1 U3009 ( .A1(n3186), .A2(n2737), .ZN(n2338) );
  NAND2_X1 U3010 ( .A1(n2339), .A2(n2338), .ZN(n2343) );
  XNOR2_X1 U3011 ( .A(n2342), .B(n2343), .ZN(n3098) );
  INV_X1 U3012 ( .A(n3098), .ZN(n2340) );
  INV_X1 U3013 ( .A(n2342), .ZN(n2345) );
  INV_X1 U3014 ( .A(n2343), .ZN(n2344) );
  NAND2_X1 U3015 ( .A1(n2345), .A2(n2344), .ZN(n2346) );
  NAND2_X1 U3016 ( .A1(n3100), .A2(n2346), .ZN(n3130) );
  NAND2_X1 U3017 ( .A1(n2330), .A2(n3151), .ZN(n2351) );
  NAND2_X1 U3018 ( .A1(n2973), .A2(REG0_REG_3__SCAN_IN), .ZN(n2350) );
  NAND2_X1 U3019 ( .A1(n2672), .A2(REG2_REG_3__SCAN_IN), .ZN(n2349) );
  NAND2_X1 U3020 ( .A1(n2398), .A2(REG1_REG_3__SCAN_IN), .ZN(n2348) );
  NAND2_X1 U3021 ( .A1(n2352), .A2(IR_REG_31__SCAN_IN), .ZN(n2354) );
  NAND2_X1 U3022 ( .A1(n2354), .A2(n2353), .ZN(n2368) );
  OR2_X1 U3023 ( .A1(n2354), .A2(n2353), .ZN(n2355) );
  MUX2_X1 U3024 ( .A(n4348), .B(DATAI_3_), .S(n2712), .Z(n3142) );
  NAND2_X1 U3025 ( .A1(n3142), .A2(n2738), .ZN(n2356) );
  AOI22_X1 U3026 ( .A1(n3213), .A2(n2307), .B1(n3142), .B2(n2737), .ZN(n2358)
         );
  XNOR2_X1 U3027 ( .A(n2357), .B(n2358), .ZN(n3131) );
  INV_X1 U3028 ( .A(n2357), .ZN(n2359) );
  NAND2_X1 U3029 ( .A1(n2359), .A2(n2358), .ZN(n2360) );
  NAND2_X1 U3030 ( .A1(n2973), .A2(REG0_REG_4__SCAN_IN), .ZN(n2367) );
  NAND2_X1 U3031 ( .A1(n2672), .A2(REG2_REG_4__SCAN_IN), .ZN(n2362) );
  NAND2_X1 U3032 ( .A1(n2398), .A2(REG1_REG_4__SCAN_IN), .ZN(n2361) );
  NAND2_X1 U3033 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2378) );
  OAI21_X1 U3034 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        n2378), .ZN(n3221) );
  INV_X1 U3035 ( .A(n3221), .ZN(n2363) );
  AND2_X1 U3036 ( .A1(n2330), .A2(n2363), .ZN(n2364) );
  NOR2_X1 U3037 ( .A1(n2365), .A2(n2364), .ZN(n2366) );
  NAND2_X1 U3038 ( .A1(n2367), .A2(n2366), .ZN(n3781) );
  INV_X1 U3039 ( .A(n3781), .ZN(n2825) );
  NAND2_X1 U3040 ( .A1(n2368), .A2(IR_REG_31__SCAN_IN), .ZN(n2369) );
  MUX2_X1 U3041 ( .A(n4347), .B(DATAI_4_), .S(n3622), .Z(n3212) );
  INV_X1 U3042 ( .A(n3212), .ZN(n3219) );
  OAI22_X1 U3043 ( .A1(n2825), .A2(n2321), .B1(n2752), .B2(n3219), .ZN(n2371)
         );
  XNOR2_X1 U3044 ( .A(n2371), .B(n2753), .ZN(n2376) );
  OR2_X1 U3045 ( .A1(n2825), .A2(n2755), .ZN(n2373) );
  NAND2_X1 U3046 ( .A1(n3212), .A2(n2737), .ZN(n2372) );
  NAND2_X1 U3047 ( .A1(n2373), .A2(n2372), .ZN(n2375) );
  XNOR2_X1 U3048 ( .A(n2376), .B(n2375), .ZN(n3155) );
  INV_X1 U3049 ( .A(n3155), .ZN(n2374) );
  NAND2_X1 U3050 ( .A1(n2376), .A2(n2375), .ZN(n2377) );
  NAND2_X1 U3051 ( .A1(n3157), .A2(n2377), .ZN(n3165) );
  NOR2_X1 U3052 ( .A1(n2378), .A2(n3059), .ZN(n2393) );
  AND2_X1 U3053 ( .A1(n2378), .A2(n3059), .ZN(n2379) );
  NOR2_X1 U3054 ( .A1(n2393), .A2(n2379), .ZN(n3206) );
  INV_X1 U3055 ( .A(n2380), .ZN(n2384) );
  NAND2_X1 U3056 ( .A1(n2381), .A2(IR_REG_31__SCAN_IN), .ZN(n2382) );
  MUX2_X1 U3057 ( .A(IR_REG_31__SCAN_IN), .B(n2382), .S(IR_REG_5__SCAN_IN), 
        .Z(n2383) );
  NAND2_X1 U3058 ( .A1(n2384), .A2(n2383), .ZN(n3062) );
  INV_X1 U3059 ( .A(DATAI_5_), .ZN(n2385) );
  MUX2_X1 U3060 ( .A(n3062), .B(n2385), .S(n3622), .Z(n2874) );
  OAI22_X1 U3061 ( .A1(n2828), .A2(n2321), .B1(n2752), .B2(n2874), .ZN(n2386)
         );
  XNOR2_X1 U3062 ( .A(n2386), .B(n2741), .ZN(n2389) );
  OR2_X1 U3063 ( .A1(n2828), .A2(n2755), .ZN(n2388) );
  NAND2_X1 U3064 ( .A1(n3204), .A2(n2737), .ZN(n2387) );
  NAND2_X1 U3065 ( .A1(n2388), .A2(n2387), .ZN(n2390) );
  XNOR2_X1 U3066 ( .A(n2389), .B(n2390), .ZN(n3164) );
  NAND2_X1 U3067 ( .A1(n3165), .A2(n3164), .ZN(n3163) );
  INV_X1 U3068 ( .A(n2389), .ZN(n2391) );
  NAND2_X1 U3069 ( .A1(n2391), .A2(n2390), .ZN(n2392) );
  NAND2_X1 U3070 ( .A1(n2393), .A2(REG3_REG_6__SCAN_IN), .ZN(n2411) );
  OR2_X1 U3071 ( .A1(n2393), .A2(REG3_REG_6__SCAN_IN), .ZN(n2394) );
  AND2_X1 U3072 ( .A1(n2411), .A2(n2394), .ZN(n3318) );
  NAND2_X1 U3073 ( .A1(n2330), .A2(n3318), .ZN(n2396) );
  NAND2_X1 U3074 ( .A1(n2973), .A2(REG0_REG_6__SCAN_IN), .ZN(n2395) );
  NAND2_X1 U3075 ( .A1(n2396), .A2(n2395), .ZN(n2397) );
  NOR2_X1 U3076 ( .A1(n2397), .A2(n2253), .ZN(n2400) );
  CLKBUF_X3 U3077 ( .A(n2398), .Z(n3605) );
  NAND2_X1 U3078 ( .A1(n3605), .A2(REG1_REG_6__SCAN_IN), .ZN(n2399) );
  NAND2_X1 U3079 ( .A1(n3288), .A2(n2307), .ZN(n2406) );
  NOR2_X1 U3080 ( .A1(n2380), .A2(n2601), .ZN(n2401) );
  MUX2_X1 U3081 ( .A(n2601), .B(n2401), .S(IR_REG_6__SCAN_IN), .Z(n2404) );
  NAND2_X1 U3082 ( .A1(n2380), .A2(n2402), .ZN(n2447) );
  INV_X1 U3083 ( .A(n2447), .ZN(n2403) );
  MUX2_X1 U3084 ( .A(n4345), .B(DATAI_6_), .S(n2712), .Z(n3308) );
  NAND2_X1 U3085 ( .A1(n3308), .A2(n2737), .ZN(n2405) );
  NAND2_X1 U3086 ( .A1(n2406), .A2(n2405), .ZN(n3312) );
  NAND2_X1 U3087 ( .A1(n3288), .A2(n2737), .ZN(n2408) );
  NAND2_X1 U3088 ( .A1(n3308), .A2(n2738), .ZN(n2407) );
  NAND2_X1 U3089 ( .A1(n2408), .A2(n2407), .ZN(n2409) );
  XNOR2_X1 U3090 ( .A(n2409), .B(n2753), .ZN(n3311) );
  NAND2_X1 U3091 ( .A1(n2411), .A2(n2410), .ZN(n2412) );
  AND2_X1 U3092 ( .A1(n2425), .A2(n2412), .ZN(n3232) );
  NAND2_X1 U3093 ( .A1(n2330), .A2(n3232), .ZN(n2416) );
  NAND2_X1 U3094 ( .A1(n2973), .A2(REG0_REG_7__SCAN_IN), .ZN(n2415) );
  NAND2_X1 U3095 ( .A1(n3605), .A2(REG1_REG_7__SCAN_IN), .ZN(n2414) );
  NAND2_X1 U3096 ( .A1(n2672), .A2(REG2_REG_7__SCAN_IN), .ZN(n2413) );
  NAND2_X1 U3097 ( .A1(n2447), .A2(IR_REG_31__SCAN_IN), .ZN(n2432) );
  XNOR2_X1 U3098 ( .A(n2432), .B(IR_REG_7__SCAN_IN), .ZN(n4344) );
  MUX2_X1 U3099 ( .A(n4344), .B(DATAI_7_), .S(n2712), .Z(n3292) );
  OAI22_X1 U3100 ( .A1(n2833), .A2(n2321), .B1(n2752), .B2(n3231), .ZN(n2417)
         );
  XNOR2_X1 U3101 ( .A(n2417), .B(n2741), .ZN(n2420) );
  OR2_X1 U3102 ( .A1(n2833), .A2(n2755), .ZN(n2419) );
  NAND2_X1 U3103 ( .A1(n3292), .A2(n2737), .ZN(n2418) );
  NAND2_X1 U3104 ( .A1(n2419), .A2(n2418), .ZN(n2421) );
  XNOR2_X1 U3105 ( .A(n2420), .B(n2421), .ZN(n3286) );
  INV_X1 U3106 ( .A(n2420), .ZN(n2422) );
  NAND2_X1 U3107 ( .A1(n2422), .A2(n2421), .ZN(n2423) );
  NAND2_X1 U3108 ( .A1(n2425), .A2(n2424), .ZN(n2426) );
  AND2_X1 U3109 ( .A1(n2440), .A2(n2426), .ZN(n3304) );
  NAND2_X1 U3110 ( .A1(n2705), .A2(n3304), .ZN(n2430) );
  NAND2_X1 U3111 ( .A1(n2973), .A2(REG0_REG_8__SCAN_IN), .ZN(n2429) );
  NAND2_X1 U3112 ( .A1(n3605), .A2(REG1_REG_8__SCAN_IN), .ZN(n2428) );
  NAND2_X1 U3113 ( .A1(n2672), .A2(REG2_REG_8__SCAN_IN), .ZN(n2427) );
  INV_X1 U3114 ( .A(IR_REG_7__SCAN_IN), .ZN(n2431) );
  NAND2_X1 U3115 ( .A1(n2432), .A2(n2431), .ZN(n2433) );
  NAND2_X1 U3116 ( .A1(n2433), .A2(IR_REG_31__SCAN_IN), .ZN(n2435) );
  INV_X1 U3117 ( .A(IR_REG_8__SCAN_IN), .ZN(n2434) );
  XNOR2_X1 U3118 ( .A(n2435), .B(n2434), .ZN(n3037) );
  INV_X1 U3119 ( .A(DATAI_8_), .ZN(n2436) );
  MUX2_X1 U3120 ( .A(n3037), .B(n2436), .S(n2712), .Z(n3302) );
  OAI22_X1 U3121 ( .A1(n3360), .A2(n2321), .B1(n2752), .B2(n3302), .ZN(n2437)
         );
  XNOR2_X1 U3122 ( .A(n2437), .B(n2753), .ZN(n2459) );
  OR2_X1 U3123 ( .A1(n3360), .A2(n2755), .ZN(n2439) );
  NAND2_X1 U3124 ( .A1(n3279), .A2(n2737), .ZN(n2438) );
  NAND2_X1 U3125 ( .A1(n2439), .A2(n2438), .ZN(n2460) );
  AND2_X1 U3126 ( .A1(n2459), .A2(n2460), .ZN(n3354) );
  AND2_X1 U3127 ( .A1(n2440), .A2(n3359), .ZN(n2441) );
  NOR2_X1 U3128 ( .A1(n2466), .A2(n2441), .ZN(n3364) );
  NAND2_X1 U3129 ( .A1(n2705), .A2(n3364), .ZN(n2446) );
  NAND2_X1 U3130 ( .A1(n2973), .A2(REG0_REG_9__SCAN_IN), .ZN(n2445) );
  NAND2_X1 U3131 ( .A1(n3605), .A2(REG1_REG_9__SCAN_IN), .ZN(n2444) );
  NAND2_X1 U3132 ( .A1(n2672), .A2(REG2_REG_9__SCAN_IN), .ZN(n2443) );
  NAND4_X1 U3133 ( .A1(n2446), .A2(n2445), .A3(n2444), .A4(n2443), .ZN(n3777)
         );
  NAND2_X1 U3134 ( .A1(n3777), .A2(n2737), .ZN(n2453) );
  NAND2_X1 U3135 ( .A1(n2449), .A2(IR_REG_31__SCAN_IN), .ZN(n2448) );
  MUX2_X1 U3136 ( .A(IR_REG_31__SCAN_IN), .B(n2448), .S(IR_REG_9__SCAN_IN), 
        .Z(n2451) );
  INV_X1 U3137 ( .A(n2490), .ZN(n2450) );
  NAND2_X1 U3138 ( .A1(n2451), .A2(n2450), .ZN(n4478) );
  INV_X1 U3139 ( .A(n4478), .ZN(n3039) );
  MUX2_X1 U3140 ( .A(n3039), .B(DATAI_9_), .S(n2712), .Z(n3322) );
  NAND2_X1 U3141 ( .A1(n3322), .A2(n2738), .ZN(n2452) );
  NAND2_X1 U3142 ( .A1(n2453), .A2(n2452), .ZN(n2454) );
  XNOR2_X1 U3143 ( .A(n2454), .B(n2753), .ZN(n2457) );
  INV_X1 U3144 ( .A(n2457), .ZN(n2455) );
  AOI22_X1 U3145 ( .A1(n3777), .A2(n2307), .B1(n3322), .B2(n2737), .ZN(n2456)
         );
  NAND2_X1 U3146 ( .A1(n2455), .A2(n2456), .ZN(n2463) );
  INV_X1 U3147 ( .A(n2463), .ZN(n2458) );
  XNOR2_X1 U31480 ( .A(n2457), .B(n2456), .ZN(n3358) );
  NOR2_X1 U31490 ( .A1(n2458), .A2(n3358), .ZN(n2465) );
  INV_X1 U3150 ( .A(n2459), .ZN(n2462) );
  INV_X1 U3151 ( .A(n2460), .ZN(n2461) );
  NAND2_X1 U3152 ( .A1(n2462), .A2(n2461), .ZN(n3355) );
  AND2_X1 U3153 ( .A1(n3355), .A2(n2463), .ZN(n2464) );
  OR2_X1 U3154 ( .A1(n2465), .A2(n2464), .ZN(n3342) );
  OR2_X1 U3155 ( .A1(n2466), .A2(REG3_REG_10__SCAN_IN), .ZN(n2467) );
  NAND2_X1 U3156 ( .A1(n2466), .A2(REG3_REG_10__SCAN_IN), .ZN(n2483) );
  AND2_X1 U3157 ( .A1(n2467), .A2(n2483), .ZN(n3385) );
  NAND2_X1 U3158 ( .A1(n2705), .A2(n3385), .ZN(n2471) );
  NAND2_X1 U3159 ( .A1(n2973), .A2(REG0_REG_10__SCAN_IN), .ZN(n2470) );
  NAND2_X1 U3160 ( .A1(n3605), .A2(REG1_REG_10__SCAN_IN), .ZN(n2469) );
  NAND2_X1 U3161 ( .A1(n2672), .A2(REG2_REG_10__SCAN_IN), .ZN(n2468) );
  NAND4_X1 U3162 ( .A1(n2471), .A2(n2470), .A3(n2469), .A4(n2468), .ZN(n3776)
         );
  NAND2_X1 U3163 ( .A1(n3776), .A2(n2737), .ZN(n2474) );
  OR2_X1 U3164 ( .A1(n2490), .A2(n2601), .ZN(n2472) );
  XNOR2_X1 U3165 ( .A(n2472), .B(IR_REG_10__SCAN_IN), .ZN(n3830) );
  MUX2_X1 U3166 ( .A(n3830), .B(DATAI_10_), .S(n2712), .Z(n3350) );
  NAND2_X1 U3167 ( .A1(n3350), .A2(n2738), .ZN(n2473) );
  NAND2_X1 U3168 ( .A1(n2474), .A2(n2473), .ZN(n2475) );
  XNOR2_X1 U3169 ( .A(n2475), .B(n2741), .ZN(n2478) );
  AOI22_X1 U3170 ( .A1(n3776), .A2(n2307), .B1(n2737), .B2(n3350), .ZN(n2479)
         );
  XNOR2_X1 U3171 ( .A(n2478), .B(n2479), .ZN(n3343) );
  INV_X1 U3172 ( .A(n3343), .ZN(n2476) );
  AND2_X1 U3173 ( .A1(n3342), .A2(n2476), .ZN(n2477) );
  INV_X1 U3174 ( .A(n2478), .ZN(n2481) );
  INV_X1 U3175 ( .A(n2479), .ZN(n2480) );
  NAND2_X1 U3176 ( .A1(n2481), .A2(n2480), .ZN(n2482) );
  NAND2_X1 U3177 ( .A1(n2483), .A2(n3371), .ZN(n2484) );
  AND2_X1 U3178 ( .A1(n2496), .A2(n2484), .ZN(n3431) );
  NAND2_X1 U3179 ( .A1(n2705), .A2(n3431), .ZN(n2488) );
  NAND2_X1 U3180 ( .A1(n2973), .A2(REG0_REG_11__SCAN_IN), .ZN(n2487) );
  NAND2_X1 U3181 ( .A1(n3605), .A2(REG1_REG_11__SCAN_IN), .ZN(n2486) );
  NAND2_X1 U3182 ( .A1(n2672), .A2(REG2_REG_11__SCAN_IN), .ZN(n2485) );
  OR2_X1 U3183 ( .A1(n3402), .A2(n2755), .ZN(n2493) );
  INV_X1 U3184 ( .A(IR_REG_10__SCAN_IN), .ZN(n2489) );
  NAND2_X1 U3185 ( .A1(n2490), .A2(n2489), .ZN(n2491) );
  NAND2_X1 U3186 ( .A1(n2491), .A2(IR_REG_31__SCAN_IN), .ZN(n2503) );
  XNOR2_X1 U3187 ( .A(n2503), .B(IR_REG_11__SCAN_IN), .ZN(n4475) );
  MUX2_X1 U3188 ( .A(n4475), .B(DATAI_11_), .S(n2712), .Z(n3421) );
  NAND2_X1 U3189 ( .A1(n3421), .A2(n2737), .ZN(n2492) );
  NAND2_X1 U3190 ( .A1(n2493), .A2(n2492), .ZN(n3368) );
  OAI22_X1 U3191 ( .A1(n3402), .A2(n2321), .B1(n2752), .B2(n3429), .ZN(n2494)
         );
  XNOR2_X1 U3192 ( .A(n2494), .B(n2753), .ZN(n3367) );
  AND2_X1 U3193 ( .A1(n2496), .A2(n2495), .ZN(n2497) );
  NOR2_X1 U3194 ( .A1(n2513), .A2(n2497), .ZN(n3409) );
  NAND2_X1 U3195 ( .A1(n2705), .A2(n3409), .ZN(n2501) );
  NAND2_X1 U3196 ( .A1(n2973), .A2(REG0_REG_12__SCAN_IN), .ZN(n2500) );
  NAND2_X1 U3197 ( .A1(n3605), .A2(REG1_REG_12__SCAN_IN), .ZN(n2499) );
  NAND2_X1 U3198 ( .A1(n3606), .A2(REG2_REG_12__SCAN_IN), .ZN(n2498) );
  NAND2_X1 U3199 ( .A1(n2503), .A2(n2502), .ZN(n2504) );
  NAND2_X1 U3200 ( .A1(n2504), .A2(IR_REG_31__SCAN_IN), .ZN(n2505) );
  XNOR2_X1 U3201 ( .A(n2505), .B(IR_REG_12__SCAN_IN), .ZN(n3846) );
  MUX2_X1 U3202 ( .A(n3846), .B(DATAI_12_), .S(n2712), .Z(n3407) );
  INV_X1 U3203 ( .A(n3407), .ZN(n2882) );
  OAI22_X1 U3204 ( .A1(n4185), .A2(n2321), .B1(n2752), .B2(n2882), .ZN(n2506)
         );
  XNOR2_X1 U3205 ( .A(n2506), .B(n2753), .ZN(n2509) );
  OR2_X1 U3206 ( .A1(n4185), .A2(n2755), .ZN(n2508) );
  NAND2_X1 U3207 ( .A1(n3407), .A2(n2737), .ZN(n2507) );
  NAND2_X1 U3208 ( .A1(n2508), .A2(n2507), .ZN(n2510) );
  AND2_X1 U3209 ( .A1(n2509), .A2(n2510), .ZN(n3392) );
  INV_X1 U32100 ( .A(n2509), .ZN(n2512) );
  INV_X1 U32110 ( .A(n2510), .ZN(n2511) );
  NAND2_X1 U32120 ( .A1(n2512), .A2(n2511), .ZN(n3391) );
  NOR2_X1 U32130 ( .A1(n2513), .A2(REG3_REG_13__SCAN_IN), .ZN(n2514) );
  OR2_X1 U32140 ( .A1(n2530), .A2(n2514), .ZN(n4194) );
  INV_X1 U32150 ( .A(n4194), .ZN(n2515) );
  NAND2_X1 U32160 ( .A1(n2705), .A2(n2515), .ZN(n2519) );
  NAND2_X1 U32170 ( .A1(n2973), .A2(REG0_REG_13__SCAN_IN), .ZN(n2518) );
  NAND2_X1 U32180 ( .A1(n3605), .A2(REG1_REG_13__SCAN_IN), .ZN(n2517) );
  NAND2_X1 U32190 ( .A1(n3606), .A2(REG2_REG_13__SCAN_IN), .ZN(n2516) );
  OR2_X1 U32200 ( .A1(n2520), .A2(n2601), .ZN(n2521) );
  XNOR2_X1 U32210 ( .A(n2521), .B(IR_REG_13__SCAN_IN), .ZN(n3849) );
  INV_X1 U32220 ( .A(DATAI_13_), .ZN(n2522) );
  MUX2_X1 U32230 ( .A(n4473), .B(n2522), .S(n3622), .Z(n4191) );
  OAI22_X1 U32240 ( .A1(n3461), .A2(n2321), .B1(n2752), .B2(n4191), .ZN(n2523)
         );
  XNOR2_X1 U32250 ( .A(n2523), .B(n2741), .ZN(n3555) );
  OR2_X1 U32260 ( .A1(n3461), .A2(n2755), .ZN(n2525) );
  NAND2_X1 U32270 ( .A1(n4181), .A2(n2737), .ZN(n2524) );
  NAND2_X1 U32280 ( .A1(n2525), .A2(n2524), .ZN(n3554) );
  NAND2_X1 U32290 ( .A1(n2526), .A2(n3554), .ZN(n2529) );
  NAND2_X1 U32300 ( .A1(n2527), .A2(n2240), .ZN(n2528) );
  NAND2_X1 U32310 ( .A1(n2530), .A2(REG3_REG_14__SCAN_IN), .ZN(n2546) );
  OR2_X1 U32320 ( .A1(n2530), .A2(REG3_REG_14__SCAN_IN), .ZN(n2531) );
  AND2_X1 U32330 ( .A1(n2546), .A2(n2531), .ZN(n4167) );
  NAND2_X1 U32340 ( .A1(n2705), .A2(n4167), .ZN(n2535) );
  NAND2_X1 U32350 ( .A1(n2973), .A2(REG0_REG_14__SCAN_IN), .ZN(n2534) );
  NAND2_X1 U32360 ( .A1(n3605), .A2(REG1_REG_14__SCAN_IN), .ZN(n2533) );
  NAND2_X1 U32370 ( .A1(n3606), .A2(REG2_REG_14__SCAN_IN), .ZN(n2532) );
  NAND2_X1 U32380 ( .A1(n2536), .A2(IR_REG_31__SCAN_IN), .ZN(n2537) );
  XNOR2_X1 U32390 ( .A(n2537), .B(IR_REG_14__SCAN_IN), .ZN(n4411) );
  MUX2_X1 U32400 ( .A(n4411), .B(DATAI_14_), .S(n2712), .Z(n2916) );
  INV_X1 U32410 ( .A(n2916), .ZN(n4165) );
  OAI22_X1 U32420 ( .A1(n4143), .A2(n2321), .B1(n4165), .B2(n2752), .ZN(n2538)
         );
  XNOR2_X1 U32430 ( .A(n2538), .B(n2753), .ZN(n2542) );
  OR2_X1 U32440 ( .A1(n4143), .A2(n2755), .ZN(n2540) );
  NAND2_X1 U32450 ( .A1(n2916), .A2(n2737), .ZN(n2539) );
  NAND2_X1 U32460 ( .A1(n2540), .A2(n2539), .ZN(n2543) );
  AND2_X1 U32470 ( .A1(n2542), .A2(n2543), .ZN(n3458) );
  INV_X1 U32480 ( .A(n3458), .ZN(n2541) );
  INV_X1 U32490 ( .A(n2542), .ZN(n2545) );
  INV_X1 U32500 ( .A(n2543), .ZN(n2544) );
  NAND2_X1 U32510 ( .A1(n2545), .A2(n2544), .ZN(n3457) );
  NAND2_X1 U32520 ( .A1(n2546), .A2(n3588), .ZN(n2547) );
  AND2_X1 U32530 ( .A1(n2579), .A2(n2547), .ZN(n4145) );
  NAND2_X1 U32540 ( .A1(n2705), .A2(n4145), .ZN(n2551) );
  NAND2_X1 U32550 ( .A1(n2973), .A2(REG0_REG_15__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U32560 ( .A1(n3605), .A2(REG1_REG_15__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U32570 ( .A1(n3606), .A2(REG2_REG_15__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U32580 ( .A1(n2020), .A2(IR_REG_31__SCAN_IN), .ZN(n2553) );
  OR2_X1 U32590 ( .A1(n2553), .A2(n2552), .ZN(n2554) );
  NAND2_X1 U32600 ( .A1(n2553), .A2(n2552), .ZN(n2564) );
  MUX2_X1 U32610 ( .A(n4343), .B(DATAI_15_), .S(n2712), .Z(n4144) );
  OAI22_X1 U32620 ( .A1(n4156), .A2(n2321), .B1(n2752), .B2(n2917), .ZN(n2555)
         );
  XNOR2_X1 U32630 ( .A(n2555), .B(n2741), .ZN(n2559) );
  OR2_X1 U32640 ( .A1(n4156), .A2(n2755), .ZN(n2557) );
  NAND2_X1 U32650 ( .A1(n4144), .A2(n2737), .ZN(n2556) );
  NAND2_X1 U32660 ( .A1(n2557), .A2(n2556), .ZN(n3598) );
  XNOR2_X1 U32670 ( .A(n2579), .B(REG3_REG_16__SCAN_IN), .ZN(n4123) );
  NAND2_X1 U32680 ( .A1(n2705), .A2(n4123), .ZN(n2563) );
  NAND2_X1 U32690 ( .A1(n2973), .A2(REG0_REG_16__SCAN_IN), .ZN(n2562) );
  NAND2_X1 U32700 ( .A1(n3605), .A2(REG1_REG_16__SCAN_IN), .ZN(n2561) );
  NAND2_X1 U32710 ( .A1(n2672), .A2(REG2_REG_16__SCAN_IN), .ZN(n2560) );
  NAND2_X1 U32720 ( .A1(n2564), .A2(IR_REG_31__SCAN_IN), .ZN(n2565) );
  XNOR2_X1 U32730 ( .A(n2565), .B(n4670), .ZN(n4470) );
  INV_X1 U32740 ( .A(n4470), .ZN(n2566) );
  MUX2_X1 U32750 ( .A(n2566), .B(DATAI_16_), .S(n2712), .Z(n4122) );
  OAI22_X1 U32760 ( .A1(n3594), .A2(n2321), .B1(n4128), .B2(n2752), .ZN(n2567)
         );
  XNOR2_X1 U32770 ( .A(n2567), .B(n2741), .ZN(n2570) );
  OR2_X1 U32780 ( .A1(n3594), .A2(n2755), .ZN(n2569) );
  NAND2_X1 U32790 ( .A1(n4122), .A2(n2737), .ZN(n2568) );
  AND2_X1 U32800 ( .A1(n2569), .A2(n2568), .ZN(n2571) );
  NAND2_X1 U32810 ( .A1(n2570), .A2(n2571), .ZN(n2576) );
  INV_X1 U32820 ( .A(n2570), .ZN(n2573) );
  INV_X1 U32830 ( .A(n2571), .ZN(n2572) );
  NAND2_X1 U32840 ( .A1(n2573), .A2(n2572), .ZN(n2574) );
  AND2_X1 U32850 ( .A1(n2576), .A2(n2574), .ZN(n3513) );
  INV_X1 U32860 ( .A(n2579), .ZN(n2577) );
  AOI21_X1 U32870 ( .B1(n2577), .B2(REG3_REG_16__SCAN_IN), .A(
        REG3_REG_17__SCAN_IN), .ZN(n2580) );
  NAND2_X1 U32880 ( .A1(REG3_REG_16__SCAN_IN), .A2(REG3_REG_17__SCAN_IN), .ZN(
        n2578) );
  OR2_X1 U32890 ( .A1(n2580), .A2(n2595), .ZN(n3523) );
  INV_X1 U32900 ( .A(n3523), .ZN(n4113) );
  NAND2_X1 U32910 ( .A1(n2705), .A2(n4113), .ZN(n2584) );
  NAND2_X1 U32920 ( .A1(n2973), .A2(REG0_REG_17__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U32930 ( .A1(n3605), .A2(REG1_REG_17__SCAN_IN), .ZN(n2582) );
  NAND2_X1 U32940 ( .A1(n3606), .A2(REG2_REG_17__SCAN_IN), .ZN(n2581) );
  OR2_X1 U32950 ( .A1(n2585), .A2(n2601), .ZN(n2586) );
  XNOR2_X1 U32960 ( .A(n2586), .B(IR_REG_17__SCAN_IN), .ZN(n3872) );
  INV_X1 U32970 ( .A(DATAI_17_), .ZN(n2587) );
  MUX2_X1 U32980 ( .A(n4468), .B(n2587), .S(n2712), .Z(n4112) );
  OAI22_X1 U32990 ( .A1(n4129), .A2(n2321), .B1(n2752), .B2(n4112), .ZN(n2588)
         );
  XNOR2_X1 U33000 ( .A(n2588), .B(n2753), .ZN(n2591) );
  OR2_X1 U33010 ( .A1(n4129), .A2(n2755), .ZN(n2590) );
  NAND2_X1 U33020 ( .A1(n3524), .A2(n2737), .ZN(n2589) );
  NAND2_X1 U33030 ( .A1(n2590), .A2(n2589), .ZN(n2592) );
  NAND2_X1 U33040 ( .A1(n2591), .A2(n2592), .ZN(n3520) );
  INV_X1 U33050 ( .A(n2591), .ZN(n2594) );
  INV_X1 U33060 ( .A(n2592), .ZN(n2593) );
  NAND2_X1 U33070 ( .A1(n2594), .A2(n2593), .ZN(n3519) );
  NAND2_X1 U33080 ( .A1(n2595), .A2(REG3_REG_18__SCAN_IN), .ZN(n2608) );
  OR2_X1 U33090 ( .A1(n2595), .A2(REG3_REG_18__SCAN_IN), .ZN(n2596) );
  AND2_X1 U33100 ( .A1(n2608), .A2(n2596), .ZN(n4097) );
  NAND2_X1 U33110 ( .A1(n2705), .A2(n4097), .ZN(n2600) );
  NAND2_X1 U33120 ( .A1(n2973), .A2(REG0_REG_18__SCAN_IN), .ZN(n2599) );
  NAND2_X1 U33130 ( .A1(n3605), .A2(REG1_REG_18__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U33140 ( .A1(n3606), .A2(REG2_REG_18__SCAN_IN), .ZN(n2597) );
  OR2_X1 U33150 ( .A1(n4106), .A2(n2755), .ZN(n2605) );
  OR2_X1 U33160 ( .A1(n2602), .A2(n2601), .ZN(n2603) );
  XNOR2_X1 U33170 ( .A(n2603), .B(IR_REG_18__SCAN_IN), .ZN(n3881) );
  MUX2_X1 U33180 ( .A(n3881), .B(DATAI_18_), .S(n3622), .Z(n4094) );
  NAND2_X1 U33190 ( .A1(n4094), .A2(n2737), .ZN(n2604) );
  NAND2_X1 U33200 ( .A1(n2605), .A2(n2604), .ZN(n3576) );
  OAI22_X1 U33210 ( .A1(n4106), .A2(n2321), .B1(n2752), .B2(n3582), .ZN(n2606)
         );
  XNOR2_X1 U33220 ( .A(n2606), .B(n2753), .ZN(n3577) );
  INV_X1 U33230 ( .A(REG3_REG_19__SCAN_IN), .ZN(n2607) );
  NAND2_X1 U33240 ( .A1(n2608), .A2(n2607), .ZN(n2609) );
  AND2_X1 U33250 ( .A1(n2628), .A2(n2609), .ZN(n4080) );
  NAND2_X1 U33260 ( .A1(n2705), .A2(n4080), .ZN(n2613) );
  NAND2_X1 U33270 ( .A1(n2973), .A2(REG0_REG_19__SCAN_IN), .ZN(n2612) );
  NAND2_X1 U33280 ( .A1(n3605), .A2(REG1_REG_19__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U33290 ( .A1(n3606), .A2(REG2_REG_19__SCAN_IN), .ZN(n2610) );
  NAND4_X1 U33300 ( .A1(n2613), .A2(n2612), .A3(n2611), .A4(n2610), .ZN(n4090)
         );
  NAND2_X1 U33310 ( .A1(n4090), .A2(n2737), .ZN(n2615) );
  MUX2_X1 U33320 ( .A(n4342), .B(DATAI_19_), .S(n2712), .Z(n2888) );
  NAND2_X1 U33330 ( .A1(n2888), .A2(n2738), .ZN(n2614) );
  NAND2_X1 U33340 ( .A1(n2615), .A2(n2614), .ZN(n2616) );
  XNOR2_X1 U33350 ( .A(n2616), .B(n2753), .ZN(n2621) );
  NAND2_X1 U33360 ( .A1(n4090), .A2(n2307), .ZN(n2618) );
  NAND2_X1 U33370 ( .A1(n2888), .A2(n2737), .ZN(n2617) );
  NAND2_X1 U33380 ( .A1(n2618), .A2(n2617), .ZN(n2622) );
  AND2_X1 U33390 ( .A1(n2621), .A2(n2622), .ZN(n2620) );
  AOI21_X1 U33400 ( .B1(n3576), .B2(n3577), .A(n2620), .ZN(n2619) );
  NAND2_X1 U33410 ( .A1(n3476), .A2(n2619), .ZN(n2627) );
  INV_X1 U33420 ( .A(n3577), .ZN(n3477) );
  INV_X1 U33430 ( .A(n3576), .ZN(n3478) );
  INV_X1 U33440 ( .A(n2620), .ZN(n3482) );
  NAND3_X1 U33450 ( .A1(n3477), .A2(n3478), .A3(n3482), .ZN(n2625) );
  INV_X1 U33460 ( .A(n2621), .ZN(n2624) );
  INV_X1 U33470 ( .A(n2622), .ZN(n2623) );
  NAND2_X1 U33480 ( .A1(n2624), .A2(n2623), .ZN(n3481) );
  AND2_X1 U33490 ( .A1(n2625), .A2(n3481), .ZN(n2626) );
  NAND2_X1 U33500 ( .A1(n2627), .A2(n2626), .ZN(n3491) );
  NAND2_X1 U33510 ( .A1(n2628), .A2(n4583), .ZN(n2629) );
  NAND2_X1 U33520 ( .A1(n2658), .A2(n2629), .ZN(n3552) );
  INV_X1 U3353 ( .A(n3552), .ZN(n4057) );
  NAND2_X1 U33540 ( .A1(n2705), .A2(n4057), .ZN(n2633) );
  NAND2_X1 U3355 ( .A1(n2973), .A2(REG0_REG_20__SCAN_IN), .ZN(n2632) );
  NAND2_X1 U3356 ( .A1(n3605), .A2(REG1_REG_20__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U3357 ( .A1(n3606), .A2(REG2_REG_20__SCAN_IN), .ZN(n2630) );
  NAND4_X1 U3358 ( .A1(n2633), .A2(n2632), .A3(n2631), .A4(n2630), .ZN(n4031)
         );
  NAND2_X1 U3359 ( .A1(n4031), .A2(n2737), .ZN(n2635) );
  NAND2_X1 U3360 ( .A1(n4054), .A2(n2738), .ZN(n2634) );
  NAND2_X1 U3361 ( .A1(n2635), .A2(n2634), .ZN(n2636) );
  XNOR2_X1 U3362 ( .A(n2636), .B(n2753), .ZN(n2639) );
  NAND2_X1 U3363 ( .A1(n4031), .A2(n2307), .ZN(n2638) );
  NAND2_X1 U3364 ( .A1(n4054), .A2(n2737), .ZN(n2637) );
  NAND2_X1 U3365 ( .A1(n2638), .A2(n2637), .ZN(n2640) );
  NAND2_X1 U3366 ( .A1(n2639), .A2(n2640), .ZN(n3545) );
  NAND2_X1 U3367 ( .A1(n3491), .A2(n3545), .ZN(n3543) );
  INV_X1 U3368 ( .A(n2639), .ZN(n2642) );
  INV_X1 U3369 ( .A(n2640), .ZN(n2641) );
  NAND2_X1 U3370 ( .A1(n2642), .A2(n2641), .ZN(n3544) );
  NAND2_X1 U3371 ( .A1(n3543), .A2(n3544), .ZN(n3494) );
  INV_X1 U3372 ( .A(n3494), .ZN(n2651) );
  XNOR2_X1 U3373 ( .A(n2658), .B(REG3_REG_21__SCAN_IN), .ZN(n4037) );
  NAND2_X1 U3374 ( .A1(n2705), .A2(n4037), .ZN(n2646) );
  NAND2_X1 U3375 ( .A1(n2973), .A2(REG0_REG_21__SCAN_IN), .ZN(n2645) );
  NAND2_X1 U3376 ( .A1(n2398), .A2(REG1_REG_21__SCAN_IN), .ZN(n2644) );
  NAND2_X1 U3377 ( .A1(n3606), .A2(REG2_REG_21__SCAN_IN), .ZN(n2643) );
  NAND4_X1 U3378 ( .A1(n2646), .A2(n2645), .A3(n2644), .A4(n2643), .ZN(n4013)
         );
  NAND2_X1 U3379 ( .A1(n4013), .A2(n2737), .ZN(n2648) );
  NAND2_X1 U3380 ( .A1(n4034), .A2(n2738), .ZN(n2647) );
  NAND2_X1 U3381 ( .A1(n2648), .A2(n2647), .ZN(n2649) );
  XNOR2_X1 U3382 ( .A(n2649), .B(n2741), .ZN(n2652) );
  NOR2_X1 U3383 ( .A1(n4028), .A2(n2321), .ZN(n2650) );
  AOI21_X1 U3384 ( .B1(n4013), .B2(n2307), .A(n2650), .ZN(n2653) );
  INV_X1 U3385 ( .A(n2652), .ZN(n2655) );
  INV_X1 U3386 ( .A(n2653), .ZN(n2654) );
  NAND2_X1 U3387 ( .A1(n2655), .A2(n2654), .ZN(n3490) );
  INV_X1 U3388 ( .A(n2658), .ZN(n2656) );
  AOI21_X1 U3389 ( .B1(n2656), .B2(REG3_REG_21__SCAN_IN), .A(
        REG3_REG_22__SCAN_IN), .ZN(n2659) );
  NAND2_X1 U3390 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2657) );
  NOR2_X1 U3391 ( .A1(n2659), .A2(n2669), .ZN(n4019) );
  NAND2_X1 U3392 ( .A1(n2705), .A2(n4019), .ZN(n2663) );
  NAND2_X1 U3393 ( .A1(n3605), .A2(REG1_REG_22__SCAN_IN), .ZN(n2662) );
  NAND2_X1 U3394 ( .A1(n3606), .A2(REG2_REG_22__SCAN_IN), .ZN(n2661) );
  NAND2_X1 U3395 ( .A1(n2973), .A2(REG0_REG_22__SCAN_IN), .ZN(n2660) );
  NAND4_X1 U3396 ( .A1(n2663), .A2(n2662), .A3(n2661), .A4(n2660), .ZN(n3996)
         );
  NAND2_X1 U3397 ( .A1(n3996), .A2(n2737), .ZN(n2665) );
  NAND2_X1 U3398 ( .A1(n4012), .A2(n2738), .ZN(n2664) );
  NAND2_X1 U3399 ( .A1(n2665), .A2(n2664), .ZN(n2666) );
  XNOR2_X1 U3400 ( .A(n2666), .B(n2741), .ZN(n2681) );
  NOR2_X1 U3401 ( .A1(n4020), .A2(n2321), .ZN(n2667) );
  AOI21_X1 U3402 ( .B1(n3996), .B2(n2307), .A(n2667), .ZN(n2680) );
  XNOR2_X1 U3403 ( .A(n2681), .B(n2680), .ZN(n3569) );
  NOR2_X1 U3404 ( .A1(n2669), .A2(REG3_REG_23__SCAN_IN), .ZN(n2670) );
  OR2_X1 U3405 ( .A1(n2686), .A2(n2670), .ZN(n4001) );
  INV_X1 U3406 ( .A(n4001), .ZN(n2671) );
  NAND2_X1 U3407 ( .A1(n2705), .A2(n2671), .ZN(n2676) );
  NAND2_X1 U3408 ( .A1(n2973), .A2(REG0_REG_23__SCAN_IN), .ZN(n2675) );
  NAND2_X1 U3409 ( .A1(n3605), .A2(REG1_REG_23__SCAN_IN), .ZN(n2674) );
  NAND2_X1 U3410 ( .A1(n3606), .A2(REG2_REG_23__SCAN_IN), .ZN(n2673) );
  OAI22_X1 U3411 ( .A1(n4016), .A2(n2321), .B1(n2752), .B2(n4000), .ZN(n2677)
         );
  XNOR2_X1 U3412 ( .A(n2677), .B(n2741), .ZN(n2683) );
  OR2_X1 U3413 ( .A1(n4016), .A2(n2755), .ZN(n2679) );
  NAND2_X1 U3414 ( .A1(n3473), .A2(n2737), .ZN(n2678) );
  NAND2_X1 U3415 ( .A1(n2679), .A2(n2678), .ZN(n2684) );
  XNOR2_X1 U3416 ( .A(n2683), .B(n2684), .ZN(n3469) );
  NAND2_X1 U3417 ( .A1(n2681), .A2(n2680), .ZN(n3467) );
  AND2_X1 U3418 ( .A1(n3469), .A2(n3467), .ZN(n2682) );
  INV_X1 U3419 ( .A(n2683), .ZN(n2685) );
  NAND2_X1 U3420 ( .A1(n2685), .A2(n2684), .ZN(n2697) );
  NOR2_X1 U3421 ( .A1(n2686), .A2(REG3_REG_24__SCAN_IN), .ZN(n2687) );
  OR2_X1 U3422 ( .A1(n2703), .A2(n2687), .ZN(n3981) );
  INV_X1 U3423 ( .A(n3981), .ZN(n2688) );
  NAND2_X1 U3424 ( .A1(n2705), .A2(n2688), .ZN(n2692) );
  NAND2_X1 U3425 ( .A1(n2973), .A2(REG0_REG_24__SCAN_IN), .ZN(n2691) );
  NAND2_X1 U3426 ( .A1(n3605), .A2(REG1_REG_24__SCAN_IN), .ZN(n2690) );
  NAND2_X1 U3427 ( .A1(n3606), .A2(REG2_REG_24__SCAN_IN), .ZN(n2689) );
  NAND4_X1 U3428 ( .A1(n2692), .A2(n2691), .A3(n2690), .A4(n2689), .ZN(n3957)
         );
  NOR2_X1 U3429 ( .A1(n3979), .A2(n2321), .ZN(n2693) );
  AOI21_X1 U3430 ( .B1(n3957), .B2(n2307), .A(n2693), .ZN(n2696) );
  INV_X1 U3431 ( .A(n2696), .ZN(n2694) );
  AND2_X1 U3432 ( .A1(n2697), .A2(n2696), .ZN(n2698) );
  NAND2_X1 U3433 ( .A1(n3957), .A2(n2737), .ZN(n2700) );
  NAND2_X1 U3434 ( .A1(n3539), .A2(n2738), .ZN(n2699) );
  NAND2_X1 U3435 ( .A1(n2700), .A2(n2699), .ZN(n2701) );
  XNOR2_X1 U3436 ( .A(n2701), .B(n2753), .ZN(n3534) );
  NAND2_X1 U3437 ( .A1(n3532), .A2(n3534), .ZN(n2702) );
  NAND2_X1 U3438 ( .A1(n2703), .A2(REG3_REG_25__SCAN_IN), .ZN(n2719) );
  OR2_X1 U3439 ( .A1(n2703), .A2(REG3_REG_25__SCAN_IN), .ZN(n2704) );
  NAND2_X1 U3440 ( .A1(n2719), .A2(n2704), .ZN(n3962) );
  NAND2_X1 U3441 ( .A1(n3606), .A2(REG2_REG_25__SCAN_IN), .ZN(n2706) );
  OAI21_X1 U3442 ( .B1(n3962), .B2(n2806), .A(n2706), .ZN(n2707) );
  INV_X1 U3443 ( .A(n2707), .ZN(n2711) );
  NAND2_X1 U3444 ( .A1(n2973), .A2(REG0_REG_25__SCAN_IN), .ZN(n2709) );
  NAND2_X1 U3445 ( .A1(n3605), .A2(REG1_REG_25__SCAN_IN), .ZN(n2708) );
  AND2_X1 U3446 ( .A1(n2709), .A2(n2708), .ZN(n2710) );
  INV_X1 U3447 ( .A(n3508), .ZN(n3961) );
  OAI22_X1 U3448 ( .A1(n3973), .A2(n2321), .B1(n2752), .B2(n3961), .ZN(n2713)
         );
  XNOR2_X1 U3449 ( .A(n2713), .B(n2753), .ZN(n2717) );
  INV_X1 U3450 ( .A(n2717), .ZN(n2715) );
  OAI22_X1 U3451 ( .A1(n3973), .A2(n2755), .B1(n2321), .B2(n3961), .ZN(n2716)
         );
  INV_X1 U3452 ( .A(n2716), .ZN(n2714) );
  NAND2_X1 U3453 ( .A1(n2715), .A2(n2714), .ZN(n3500) );
  AND2_X1 U3454 ( .A1(n2717), .A2(n2716), .ZN(n3501) );
  AOI21_X2 U3455 ( .B1(n3504), .B2(n3500), .A(n3501), .ZN(n2943) );
  INV_X1 U3456 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2718) );
  NAND2_X1 U3457 ( .A1(n2719), .A2(n2718), .ZN(n2720) );
  NAND2_X1 U34580 ( .A1(n2733), .A2(n2720), .ZN(n3940) );
  NAND2_X1 U34590 ( .A1(n2973), .A2(REG0_REG_26__SCAN_IN), .ZN(n2722) );
  NAND2_X1 U3460 ( .A1(n3605), .A2(REG1_REG_26__SCAN_IN), .ZN(n2721) );
  AND2_X1 U3461 ( .A1(n2722), .A2(n2721), .ZN(n2724) );
  NAND2_X1 U3462 ( .A1(n3606), .A2(REG2_REG_26__SCAN_IN), .ZN(n2723) );
  OAI211_X1 U3463 ( .C1(n3940), .C2(n2806), .A(n2724), .B(n2723), .ZN(n3772)
         );
  NAND2_X1 U3464 ( .A1(n3772), .A2(n2737), .ZN(n2726) );
  NAND2_X1 U3465 ( .A1(n3936), .A2(n2738), .ZN(n2725) );
  NAND2_X1 U3466 ( .A1(n2726), .A2(n2725), .ZN(n2727) );
  XNOR2_X1 U34670 ( .A(n2727), .B(n2741), .ZN(n2732) );
  INV_X1 U3468 ( .A(n2732), .ZN(n2730) );
  NOR2_X1 U34690 ( .A1(n3944), .A2(n2321), .ZN(n2728) );
  AOI21_X1 U3470 ( .B1(n3772), .B2(n2307), .A(n2728), .ZN(n2731) );
  INV_X1 U34710 ( .A(n2731), .ZN(n2729) );
  NAND2_X1 U3472 ( .A1(n2730), .A2(n2729), .ZN(n2940) );
  AND2_X1 U34730 ( .A1(n2732), .A2(n2731), .ZN(n2939) );
  INV_X1 U3474 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4662) );
  AND2_X1 U34750 ( .A1(n2733), .A2(n4662), .ZN(n2734) );
  AOI22_X1 U3476 ( .A1(n3605), .A2(REG1_REG_27__SCAN_IN), .B1(n2973), .B2(
        REG0_REG_27__SCAN_IN), .ZN(n2736) );
  NAND2_X1 U34770 ( .A1(n3606), .A2(REG2_REG_27__SCAN_IN), .ZN(n2735) );
  NAND2_X1 U3478 ( .A1(n3937), .A2(n2737), .ZN(n2740) );
  NAND2_X1 U34790 ( .A1(n3638), .A2(n2738), .ZN(n2739) );
  NAND2_X1 U3480 ( .A1(n2740), .A2(n2739), .ZN(n2742) );
  XNOR2_X1 U34810 ( .A(n2742), .B(n2741), .ZN(n2759) );
  NOR2_X1 U3482 ( .A1(n3922), .A2(n2321), .ZN(n2743) );
  AOI21_X1 U34830 ( .B1(n3937), .B2(n2307), .A(n2743), .ZN(n2758) );
  XNOR2_X1 U3484 ( .A(n2759), .B(n2758), .ZN(n2929) );
  INV_X1 U34850 ( .A(n2929), .ZN(n2744) );
  INV_X1 U3486 ( .A(n2787), .ZN(n2786) );
  NAND2_X1 U34870 ( .A1(n2745), .A2(REG3_REG_28__SCAN_IN), .ZN(n3890) );
  INV_X1 U3488 ( .A(n2745), .ZN(n2747) );
  INV_X1 U34890 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2746) );
  NAND2_X1 U3490 ( .A1(n2747), .A2(n2746), .ZN(n2748) );
  NAND2_X1 U34910 ( .A1(n3890), .A2(n2748), .ZN(n3449) );
  AOI22_X1 U3492 ( .A1(n3605), .A2(REG1_REG_28__SCAN_IN), .B1(n2973), .B2(
        REG0_REG_28__SCAN_IN), .ZN(n2750) );
  NAND2_X1 U34930 ( .A1(n3606), .A2(REG2_REG_28__SCAN_IN), .ZN(n2749) );
  INV_X1 U3494 ( .A(n3903), .ZN(n2919) );
  OAI22_X1 U34950 ( .A1(n3898), .A2(n2321), .B1(n2919), .B2(n2752), .ZN(n2754)
         );
  XNOR2_X1 U3496 ( .A(n2754), .B(n2753), .ZN(n2757) );
  OAI22_X1 U34970 ( .A1(n3898), .A2(n2755), .B1(n2919), .B2(n2321), .ZN(n2756)
         );
  XNOR2_X1 U3498 ( .A(n2757), .B(n2756), .ZN(n2790) );
  INV_X1 U34990 ( .A(n2790), .ZN(n2784) );
  OR2_X1 U3500 ( .A1(n2759), .A2(n2758), .ZN(n2788) );
  INV_X1 U35010 ( .A(n4339), .ZN(n2773) );
  NAND2_X1 U3502 ( .A1(n2775), .A2(n2773), .ZN(n2760) );
  MUX2_X1 U35030 ( .A(n2775), .B(n2760), .S(B_REG_SCAN_IN), .Z(n2761) );
  NOR4_X1 U3504 ( .A1(D_REG_14__SCAN_IN), .A2(D_REG_15__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n2765) );
  NOR4_X1 U35050 ( .A1(D_REG_12__SCAN_IN), .A2(D_REG_10__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2764) );
  NOR4_X1 U35060 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2763) );
  NOR4_X1 U35070 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_24__SCAN_IN), .ZN(n2762) );
  AND4_X1 U35080 ( .A1(n2765), .A2(n2764), .A3(n2763), .A4(n2762), .ZN(n2771)
         );
  NOR2_X1 U35090 ( .A1(D_REG_25__SCAN_IN), .A2(D_REG_4__SCAN_IN), .ZN(n2769)
         );
  NOR4_X1 U35100 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2768) );
  NOR4_X1 U35110 ( .A1(D_REG_5__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2767) );
  NOR4_X1 U35120 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n2766) );
  AND4_X1 U35130 ( .A1(n2769), .A2(n2768), .A3(n2767), .A4(n2766), .ZN(n2770)
         );
  NAND2_X1 U35140 ( .A1(n2771), .A2(n2770), .ZN(n2910) );
  INV_X1 U35150 ( .A(n2910), .ZN(n2772) );
  NAND2_X1 U35160 ( .A1(n2772), .A2(D_REG_1__SCAN_IN), .ZN(n2774) );
  INV_X1 U35170 ( .A(n2968), .ZN(n2776) );
  NAND2_X1 U35180 ( .A1(n2776), .A2(n2773), .ZN(n2909) );
  INV_X1 U35190 ( .A(n2909), .ZN(n2971) );
  AOI21_X1 U35200 ( .B1(n2911), .B2(n2774), .A(n2971), .ZN(n3110) );
  INV_X1 U35210 ( .A(D_REG_0__SCAN_IN), .ZN(n2970) );
  NAND2_X1 U35220 ( .A1(n2911), .A2(n2970), .ZN(n2778) );
  NAND2_X1 U35230 ( .A1(n2776), .A2(n2775), .ZN(n2777) );
  NAND2_X1 U35240 ( .A1(n3110), .A2(n2923), .ZN(n2811) );
  OR2_X1 U35250 ( .A1(n2811), .A2(n2988), .ZN(n2792) );
  INV_X1 U35260 ( .A(n2985), .ZN(n2903) );
  NAND2_X1 U35270 ( .A1(n4452), .A2(n4342), .ZN(n2781) );
  NAND2_X1 U35280 ( .A1(n2903), .A2(n2781), .ZN(n2782) );
  AND2_X1 U35290 ( .A1(n2784), .A2(n2783), .ZN(n2785) );
  NAND2_X1 U35300 ( .A1(n2786), .A2(n2785), .ZN(n2818) );
  NAND3_X1 U35310 ( .A1(n2787), .A2(n3563), .A3(n2790), .ZN(n2817) );
  INV_X1 U35320 ( .A(n2788), .ZN(n2789) );
  NAND3_X1 U35330 ( .A1(n2790), .A2(n3563), .A3(n2789), .ZN(n2816) );
  NAND2_X1 U35340 ( .A1(n4520), .A2(n3757), .ZN(n2912) );
  OAI21_X2 U35350 ( .B1(n2792), .B2(n4154), .A(n4193), .ZN(n3590) );
  NAND2_X1 U35360 ( .A1(n2793), .A2(n4154), .ZN(n2794) );
  NAND2_X1 U35370 ( .A1(n2811), .A2(n2794), .ZN(n3085) );
  NAND2_X1 U35380 ( .A1(n2795), .A2(n4451), .ZN(n2796) );
  INV_X1 U35390 ( .A(n2908), .ZN(n2797) );
  NAND4_X1 U35400 ( .A1(n3085), .A2(n2797), .A3(n2987), .A4(n2304), .ZN(n2798)
         );
  NAND2_X1 U35410 ( .A1(n2798), .A2(STATE_REG_SCAN_IN), .ZN(n2802) );
  INV_X1 U35420 ( .A(n2799), .ZN(n2800) );
  NAND2_X1 U35430 ( .A1(n4466), .A2(n2800), .ZN(n2801) );
  NAND2_X1 U35440 ( .A1(n2811), .A2(n3766), .ZN(n3086) );
  NOR2_X1 U35450 ( .A1(n3557), .A2(n3449), .ZN(n2814) );
  INV_X1 U35460 ( .A(n3937), .ZN(n3639) );
  NAND2_X1 U35470 ( .A1(n2803), .A2(IR_REG_31__SCAN_IN), .ZN(n2804) );
  INV_X1 U35480 ( .A(n4351), .ZN(n3796) );
  NAND2_X1 U35490 ( .A1(n3766), .A2(n3796), .ZN(n2805) );
  INV_X1 U35500 ( .A(REG2_REG_29__SCAN_IN), .ZN(n2809) );
  OR2_X1 U35510 ( .A1(n3890), .A2(n2806), .ZN(n2808) );
  AOI22_X1 U35520 ( .A1(REG1_REG_29__SCAN_IN), .A2(n3605), .B1(n2973), .B2(
        REG0_REG_29__SCAN_IN), .ZN(n2807) );
  OAI211_X1 U35530 ( .C1(n2442), .C2(n2809), .A(n2808), .B(n2807), .ZN(n3771)
         );
  NAND2_X1 U35540 ( .A1(n3766), .A2(n4351), .ZN(n2810) );
  AOI22_X1 U35550 ( .A1(n3771), .A2(n3579), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n2812) );
  OAI21_X1 U35560 ( .B1(n3639), .B2(n3581), .A(n2812), .ZN(n2813) );
  AOI211_X1 U35570 ( .C1(n3903), .C2(n3590), .A(n2814), .B(n2813), .ZN(n2815)
         );
  NAND3_X1 U35580 ( .A1(n2818), .A2(n2817), .A3(n2258), .ZN(U3217) );
  INV_X1 U35590 ( .A(n3087), .ZN(n2819) );
  NAND2_X1 U35600 ( .A1(n2819), .A2(n3112), .ZN(n3640) );
  NAND2_X1 U35610 ( .A1(n3640), .A2(n3643), .ZN(n2870) );
  CLKBUF_X1 U35620 ( .A(n2819), .Z(n4279) );
  NAND2_X1 U35630 ( .A1(n4279), .A2(n3117), .ZN(n2820) );
  NAND2_X1 U35640 ( .A1(n3116), .A2(n2820), .ZN(n3174) );
  INV_X1 U35650 ( .A(n3174), .ZN(n2821) );
  NAND2_X1 U35660 ( .A1(n3782), .A2(n3102), .ZN(n3647) );
  NAND2_X1 U35670 ( .A1(n2822), .A2(n3186), .ZN(n3644) );
  NAND2_X1 U35680 ( .A1(n2821), .A2(n2871), .ZN(n3172) );
  NAND2_X1 U35690 ( .A1(n2822), .A2(n3102), .ZN(n2823) );
  NAND2_X1 U35700 ( .A1(n3172), .A2(n2823), .ZN(n3139) );
  NAND2_X1 U35710 ( .A1(n3213), .A2(n3142), .ZN(n2824) );
  NAND2_X1 U35720 ( .A1(n3139), .A2(n2824), .ZN(n3195) );
  NAND2_X1 U35730 ( .A1(n3781), .A2(n3219), .ZN(n3653) );
  NAND2_X1 U35740 ( .A1(n2825), .A2(n3212), .ZN(n3650) );
  NAND2_X1 U35750 ( .A1(n3653), .A2(n3650), .ZN(n3196) );
  NAND2_X1 U35760 ( .A1(n3196), .A2(n2259), .ZN(n3254) );
  INV_X2 U35770 ( .A(n3142), .ZN(n3149) );
  INV_X1 U35780 ( .A(n3288), .ZN(n2875) );
  NAND2_X1 U35790 ( .A1(n2875), .A2(n3248), .ZN(n3235) );
  NAND2_X1 U35800 ( .A1(n3194), .A2(n3235), .ZN(n2826) );
  NOR2_X1 U35810 ( .A1(n3254), .A2(n2826), .ZN(n2827) );
  NAND2_X1 U3582 ( .A1(n3195), .A2(n2827), .ZN(n2836) );
  NAND2_X1 U3583 ( .A1(n3781), .A2(n3212), .ZN(n3197) );
  NAND2_X1 U3584 ( .A1(n3780), .A2(n3204), .ZN(n2829) );
  NAND2_X1 U3585 ( .A1(n3197), .A2(n2829), .ZN(n2830) );
  NAND2_X1 U3586 ( .A1(n2830), .A2(n2259), .ZN(n3256) );
  NAND2_X1 U3587 ( .A1(n3256), .A2(n2032), .ZN(n2831) );
  NAND2_X1 U3588 ( .A1(n2831), .A2(n3235), .ZN(n3238) );
  NAND2_X1 U3589 ( .A1(n3779), .A2(n3292), .ZN(n2832) );
  AND2_X1 U3590 ( .A1(n3238), .A2(n2832), .ZN(n2835) );
  INV_X1 U3591 ( .A(n2832), .ZN(n2834) );
  NAND2_X1 U3592 ( .A1(n2833), .A2(n3292), .ZN(n2877) );
  AOI21_X1 U3593 ( .B1(n2836), .B2(n2835), .A(n2021), .ZN(n3277) );
  NAND2_X1 U3594 ( .A1(n3360), .A2(n3302), .ZN(n2837) );
  NAND2_X1 U3595 ( .A1(n3277), .A2(n2837), .ZN(n2839) );
  INV_X1 U3596 ( .A(n3360), .ZN(n3778) );
  NAND2_X1 U3597 ( .A1(n3778), .A2(n3279), .ZN(n2838) );
  AND2_X1 U3598 ( .A1(n3777), .A2(n3322), .ZN(n2840) );
  NAND2_X1 U3599 ( .A1(n3776), .A2(n3350), .ZN(n2841) );
  NAND2_X1 U3600 ( .A1(n2842), .A2(n2841), .ZN(n3419) );
  INV_X1 U3601 ( .A(n3419), .ZN(n2844) );
  NAND2_X1 U3602 ( .A1(n3402), .A2(n3421), .ZN(n3399) );
  INV_X1 U3603 ( .A(n3402), .ZN(n3007) );
  NAND2_X1 U3604 ( .A1(n3007), .A2(n3429), .ZN(n3401) );
  NAND2_X1 U3605 ( .A1(n3402), .A2(n3429), .ZN(n2845) );
  NAND2_X1 U3606 ( .A1(n3775), .A2(n3407), .ZN(n2847) );
  NAND2_X1 U3607 ( .A1(n3461), .A2(n4191), .ZN(n2848) );
  NAND2_X1 U3608 ( .A1(n4143), .A2(n2916), .ZN(n3610) );
  NAND2_X1 U3609 ( .A1(n4182), .A2(n4165), .ZN(n3611) );
  NAND2_X1 U3610 ( .A1(n3610), .A2(n3611), .ZN(n4152) );
  NAND2_X1 U3611 ( .A1(n4151), .A2(n4152), .ZN(n4150) );
  NAND2_X1 U3612 ( .A1(n4150), .A2(n2849), .ZN(n4135) );
  NAND2_X1 U3613 ( .A1(n3774), .A2(n4144), .ZN(n2851) );
  NAND2_X1 U3614 ( .A1(n3594), .A2(n4122), .ZN(n3686) );
  NAND2_X1 U3615 ( .A1(n4140), .A2(n4128), .ZN(n3683) );
  NAND2_X1 U3616 ( .A1(n3686), .A2(n3683), .ZN(n4119) );
  NAND2_X1 U3617 ( .A1(n4106), .A2(n4094), .ZN(n4066) );
  NAND2_X1 U3618 ( .A1(n4073), .A2(n3582), .ZN(n4067) );
  NAND2_X1 U3619 ( .A1(n4066), .A2(n4067), .ZN(n4089) );
  NAND2_X1 U3620 ( .A1(n4086), .A2(n4089), .ZN(n4085) );
  NAND2_X1 U3621 ( .A1(n4085), .A2(n2853), .ZN(n4062) );
  NAND2_X1 U3622 ( .A1(n4090), .A2(n2888), .ZN(n2855) );
  NOR2_X1 U3623 ( .A1(n4090), .A2(n2888), .ZN(n2854) );
  AOI21_X1 U3624 ( .B1(n4062), .B2(n2855), .A(n2854), .ZN(n4042) );
  NAND2_X1 U3625 ( .A1(n4042), .A2(n2856), .ZN(n2858) );
  NAND2_X1 U3626 ( .A1(n4031), .A2(n4054), .ZN(n2857) );
  NAND2_X1 U3627 ( .A1(n2858), .A2(n2857), .ZN(n4025) );
  INV_X1 U3628 ( .A(n4013), .ZN(n4044) );
  NOR2_X1 U3629 ( .A1(n4044), .A2(n4028), .ZN(n2859) );
  INV_X1 U3630 ( .A(n3996), .ZN(n4029) );
  NAND2_X1 U3631 ( .A1(n4029), .A2(n4012), .ZN(n3991) );
  NAND2_X1 U3632 ( .A1(n3996), .A2(n4020), .ZN(n2893) );
  NAND2_X1 U3633 ( .A1(n3996), .A2(n4012), .ZN(n2860) );
  NOR2_X1 U3634 ( .A1(n3994), .A2(n3979), .ZN(n2862) );
  NAND2_X1 U3635 ( .A1(n3994), .A2(n3979), .ZN(n2861) );
  OAI21_X1 U3636 ( .B1(n3968), .B2(n2862), .A(n2861), .ZN(n3950) );
  NOR2_X1 U3637 ( .A1(n3535), .A2(n3508), .ZN(n2863) );
  NOR2_X1 U3638 ( .A1(n3950), .A2(n2863), .ZN(n2864) );
  INV_X1 U3639 ( .A(n3772), .ZN(n3955) );
  NAND2_X1 U3640 ( .A1(n3955), .A2(n3944), .ZN(n2865) );
  NAND2_X1 U3641 ( .A1(n2866), .A2(n2254), .ZN(n2868) );
  NAND2_X1 U3642 ( .A1(n3937), .A2(n3638), .ZN(n2867) );
  OR2_X1 U3643 ( .A1(n3898), .A2(n3903), .ZN(n3892) );
  NAND2_X1 U3644 ( .A1(n3898), .A2(n3903), .ZN(n3623) );
  NAND2_X1 U3645 ( .A1(n3892), .A2(n3623), .ZN(n3904) );
  XNOR2_X1 U3646 ( .A(n4341), .B(n3125), .ZN(n2869) );
  INV_X1 U3647 ( .A(n4520), .ZN(n4480) );
  INV_X1 U3648 ( .A(n3784), .ZN(n3094) );
  NAND2_X1 U3649 ( .A1(n3094), .A2(n4282), .ZN(n3730) );
  NAND2_X1 U3650 ( .A1(n3178), .A2(n3142), .ZN(n3649) );
  NAND2_X1 U3651 ( .A1(n3213), .A2(n3149), .ZN(n3646) );
  NAND2_X1 U3652 ( .A1(n3141), .A2(n3746), .ZN(n2872) );
  INV_X1 U3653 ( .A(n3650), .ZN(n2873) );
  AND2_X1 U3654 ( .A1(n3780), .A2(n2874), .ZN(n3198) );
  NAND2_X1 U3655 ( .A1(n2828), .A2(n3204), .ZN(n3663) );
  NAND2_X1 U3656 ( .A1(n3288), .A2(n3248), .ZN(n3664) );
  NAND2_X1 U3657 ( .A1(n3244), .A2(n3664), .ZN(n2876) );
  NAND2_X1 U3658 ( .A1(n2875), .A2(n3308), .ZN(n3655) );
  INV_X1 U3659 ( .A(n2877), .ZN(n2878) );
  NAND2_X1 U3660 ( .A1(n3360), .A2(n3279), .ZN(n3659) );
  NAND2_X1 U3661 ( .A1(n3778), .A2(n3302), .ZN(n3657) );
  NAND2_X1 U3662 ( .A1(n2879), .A2(n3657), .ZN(n3321) );
  AND2_X1 U3663 ( .A1(n3777), .A2(n2150), .ZN(n3320) );
  INV_X1 U3664 ( .A(n3777), .ZN(n2880) );
  NAND2_X1 U3665 ( .A1(n2880), .A2(n3322), .ZN(n3660) );
  NAND2_X1 U3666 ( .A1(n3776), .A2(n3382), .ZN(n3672) );
  NAND2_X1 U3667 ( .A1(n3377), .A2(n3672), .ZN(n2881) );
  INV_X1 U3668 ( .A(n3776), .ZN(n3423) );
  NAND2_X1 U3669 ( .A1(n3423), .A2(n3350), .ZN(n3671) );
  NAND2_X1 U3670 ( .A1(n2881), .A2(n3671), .ZN(n3417) );
  NAND2_X1 U3671 ( .A1(n3775), .A2(n2882), .ZN(n4175) );
  NAND2_X1 U3672 ( .A1(n4158), .A2(n4191), .ZN(n3734) );
  NAND2_X1 U3673 ( .A1(n4175), .A2(n3734), .ZN(n2884) );
  INV_X1 U3674 ( .A(n3401), .ZN(n2883) );
  NOR2_X1 U3675 ( .A1(n2884), .A2(n2883), .ZN(n3673) );
  NAND2_X1 U3676 ( .A1(n3417), .A2(n3673), .ZN(n2887) );
  NAND2_X1 U3677 ( .A1(n4185), .A2(n3407), .ZN(n4177) );
  NAND2_X1 U3678 ( .A1(n3399), .A2(n4177), .ZN(n2886) );
  INV_X1 U3679 ( .A(n2884), .ZN(n2885) );
  NOR2_X1 U3680 ( .A1(n4158), .A2(n4191), .ZN(n3735) );
  AOI21_X1 U3681 ( .B1(n2886), .B2(n2885), .A(n3735), .ZN(n3676) );
  NAND2_X1 U3682 ( .A1(n4156), .A2(n4144), .ZN(n3613) );
  NAND2_X1 U3683 ( .A1(n3774), .A2(n2917), .ZN(n3612) );
  NAND2_X1 U3684 ( .A1(n3613), .A2(n3612), .ZN(n3745) );
  NAND2_X1 U3685 ( .A1(n4137), .A2(n3612), .ZN(n4127) );
  NAND2_X1 U3686 ( .A1(n4127), .A2(n2189), .ZN(n4126) );
  NAND2_X1 U3687 ( .A1(n4090), .A2(n4076), .ZN(n3731) );
  AND2_X1 U3688 ( .A1(n4067), .A2(n3731), .ZN(n2889) );
  NAND2_X1 U3689 ( .A1(n3773), .A2(n4112), .ZN(n4063) );
  NAND2_X1 U3690 ( .A1(n2889), .A2(n4063), .ZN(n3685) );
  NAND2_X1 U3691 ( .A1(n4129), .A2(n3524), .ZN(n4064) );
  NAND2_X1 U3692 ( .A1(n4066), .A2(n4064), .ZN(n2890) );
  NOR2_X1 U3693 ( .A1(n4090), .A2(n4076), .ZN(n3732) );
  AOI21_X1 U3694 ( .B1(n2890), .B2(n2889), .A(n3732), .ZN(n4045) );
  INV_X1 U3695 ( .A(n4031), .ZN(n4071) );
  NAND2_X1 U3696 ( .A1(n4071), .A2(n4054), .ZN(n2891) );
  AND2_X1 U3697 ( .A1(n4045), .A2(n2891), .ZN(n3615) );
  INV_X1 U3698 ( .A(n4054), .ZN(n4043) );
  NAND2_X1 U3699 ( .A1(n4031), .A2(n4043), .ZN(n3688) );
  NAND2_X1 U3700 ( .A1(n2892), .A2(n3688), .ZN(n4026) );
  NAND2_X1 U3701 ( .A1(n4044), .A2(n4034), .ZN(n3989) );
  AND2_X1 U3702 ( .A1(n3991), .A2(n3989), .ZN(n3692) );
  NAND2_X1 U3703 ( .A1(n4026), .A2(n3692), .ZN(n2896) );
  OR2_X1 U3704 ( .A1(n4016), .A2(n3473), .ZN(n3718) );
  AND2_X1 U3705 ( .A1(n3718), .A2(n2893), .ZN(n3696) );
  AND2_X1 U3706 ( .A1(n4013), .A2(n4028), .ZN(n3988) );
  NAND2_X1 U3707 ( .A1(n3991), .A2(n3988), .ZN(n2894) );
  NAND2_X1 U3708 ( .A1(n3696), .A2(n2894), .ZN(n3617) );
  INV_X1 U3709 ( .A(n3617), .ZN(n2895) );
  NAND2_X1 U3710 ( .A1(n2896), .A2(n2895), .ZN(n3970) );
  NAND2_X1 U3711 ( .A1(n4016), .A2(n3473), .ZN(n3969) );
  NAND2_X1 U3712 ( .A1(n3994), .A2(n3539), .ZN(n3717) );
  NAND2_X1 U3713 ( .A1(n3969), .A2(n3717), .ZN(n3694) );
  INV_X1 U3714 ( .A(n3694), .ZN(n2897) );
  NAND2_X1 U3715 ( .A1(n3955), .A2(n3936), .ZN(n3727) );
  NAND2_X1 U3716 ( .A1(n3973), .A2(n3508), .ZN(n3930) );
  AND2_X1 U3717 ( .A1(n3727), .A2(n3930), .ZN(n3621) );
  INV_X1 U3718 ( .A(n3621), .ZN(n3693) );
  NAND2_X1 U3719 ( .A1(n3535), .A2(n3961), .ZN(n3716) );
  NAND2_X1 U3720 ( .A1(n3957), .A2(n3979), .ZN(n3951) );
  AND2_X1 U3721 ( .A1(n3716), .A2(n3951), .ZN(n3932) );
  OR2_X1 U3722 ( .A1(n3693), .A2(n3932), .ZN(n2898) );
  AND2_X1 U3723 ( .A1(n3772), .A2(n3944), .ZN(n3629) );
  INV_X1 U3724 ( .A(n3629), .ZN(n3728) );
  NAND2_X1 U3725 ( .A1(n2898), .A2(n3728), .ZN(n3698) );
  INV_X1 U3726 ( .A(n3698), .ZN(n2899) );
  XNOR2_X1 U3727 ( .A(n3937), .B(n3922), .ZN(n3919) );
  OR2_X1 U3728 ( .A1(n3937), .A2(n3922), .ZN(n3624) );
  NAND2_X1 U3729 ( .A1(n3914), .A2(n3624), .ZN(n3893) );
  XNOR2_X1 U3730 ( .A(n3893), .B(n2173), .ZN(n2907) );
  NAND2_X1 U3731 ( .A1(n4341), .A2(n4342), .ZN(n2902) );
  NAND2_X1 U3732 ( .A1(n3759), .A2(n3641), .ZN(n3635) );
  NAND2_X1 U3733 ( .A1(n3937), .A2(n4159), .ZN(n2905) );
  NAND2_X1 U3734 ( .A1(n3771), .A2(n4280), .ZN(n2904) );
  OAI211_X1 U3735 ( .C1(n4154), .C2(n2919), .A(n2905), .B(n2904), .ZN(n2906)
         );
  AOI21_X1 U3736 ( .B1(n2907), .B2(n4281), .A(n2906), .ZN(n3450) );
  OAI21_X1 U3737 ( .B1(n3455), .B2(n4496), .A(n3450), .ZN(n2925) );
  OAI21_X1 U3738 ( .B1(n2965), .B2(D_REG_1__SCAN_IN), .A(n2909), .ZN(n2914) );
  NAND2_X1 U3739 ( .A1(n2911), .A2(n2910), .ZN(n2913) );
  NAND4_X1 U3740 ( .A1(n3109), .A2(n2914), .A3(n2913), .A4(n2912), .ZN(n2924)
         );
  INV_X1 U3741 ( .A(n2915), .ZN(n2922) );
  NAND2_X1 U3742 ( .A1(n4163), .A2(n2917), .ZN(n4121) );
  INV_X1 U3743 ( .A(n3921), .ZN(n2920) );
  OAI21_X1 U3744 ( .B1(n2920), .B2(n2919), .A(n3907), .ZN(n3447) );
  NAND2_X1 U3745 ( .A1(n2922), .A2(n2921), .ZN(U3546) );
  INV_X1 U3746 ( .A(n2926), .ZN(n2928) );
  NAND2_X1 U3747 ( .A1(n2928), .A2(n2927), .ZN(U3514) );
  XNOR2_X1 U3748 ( .A(n2930), .B(n2929), .ZN(n2931) );
  NAND2_X1 U3749 ( .A1(n2931), .A2(n3563), .ZN(n2938) );
  NOR2_X1 U3750 ( .A1(n3955), .A2(n3581), .ZN(n2933) );
  OAI22_X1 U3751 ( .A1(n3898), .A2(n3593), .B1(STATE_REG_SCAN_IN), .B2(n4662), 
        .ZN(n2932) );
  AOI211_X1 U3752 ( .C1(n3638), .C2(n3590), .A(n2933), .B(n2932), .ZN(n2936)
         );
  INV_X1 U3753 ( .A(n3924), .ZN(n2934) );
  AND2_X1 U3754 ( .A1(n2936), .A2(n2935), .ZN(n2937) );
  NAND2_X1 U3755 ( .A1(n2938), .A2(n2937), .ZN(U3211) );
  INV_X1 U3756 ( .A(n2939), .ZN(n2941) );
  NAND2_X1 U3757 ( .A1(n2941), .A2(n2940), .ZN(n2942) );
  XNOR2_X1 U3758 ( .A(n2943), .B(n2942), .ZN(n2944) );
  NAND2_X1 U3759 ( .A1(n3937), .A2(n3579), .ZN(n2946) );
  NAND2_X1 U3760 ( .A1(U3149), .A2(REG3_REG_26__SCAN_IN), .ZN(n2945) );
  OAI211_X1 U3761 ( .C1(n3973), .C2(n3581), .A(n2946), .B(n2945), .ZN(n2947)
         );
  INV_X1 U3762 ( .A(n2947), .ZN(n2948) );
  NAND4_X1 U3763 ( .A1(n2255), .A2(n2249), .A3(n2251), .A4(n2948), .ZN(U3237)
         );
  INV_X1 U3764 ( .A(n4466), .ZN(n2967) );
  INV_X1 U3765 ( .A(n3807), .ZN(n2998) );
  INV_X1 U3766 ( .A(DATAI_2_), .ZN(n2949) );
  MUX2_X1 U3767 ( .A(n2998), .B(n2949), .S(U3149), .Z(n2950) );
  INV_X1 U3768 ( .A(n2950), .ZN(U3350) );
  MUX2_X1 U3769 ( .A(n2436), .B(n3037), .S(STATE_REG_SCAN_IN), .Z(n2951) );
  INV_X1 U3770 ( .A(n2951), .ZN(U3344) );
  INV_X1 U3771 ( .A(DATAI_18_), .ZN(n2953) );
  NAND2_X1 U3772 ( .A1(n3881), .A2(STATE_REG_SCAN_IN), .ZN(n2952) );
  OAI21_X1 U3773 ( .B1(STATE_REG_SCAN_IN), .B2(n2953), .A(n2952), .ZN(U3334)
         );
  INV_X1 U3774 ( .A(DATAI_10_), .ZN(n2954) );
  MUX2_X1 U3775 ( .A(n2169), .B(n2954), .S(U3149), .Z(n2955) );
  INV_X1 U3776 ( .A(n2955), .ZN(U3342) );
  INV_X1 U3777 ( .A(DATAI_20_), .ZN(n2957) );
  NAND2_X1 U3778 ( .A1(n3759), .A2(STATE_REG_SCAN_IN), .ZN(n2956) );
  OAI21_X1 U3779 ( .B1(STATE_REG_SCAN_IN), .B2(n2957), .A(n2956), .ZN(U3332)
         );
  INV_X1 U3780 ( .A(DATAI_21_), .ZN(n2959) );
  NAND2_X1 U3781 ( .A1(n3641), .A2(STATE_REG_SCAN_IN), .ZN(n2958) );
  OAI21_X1 U3782 ( .B1(STATE_REG_SCAN_IN), .B2(n2959), .A(n2958), .ZN(U3331)
         );
  INV_X1 U3783 ( .A(DATAI_26_), .ZN(n2961) );
  NAND2_X1 U3784 ( .A1(n2968), .A2(STATE_REG_SCAN_IN), .ZN(n2960) );
  OAI21_X1 U3785 ( .B1(STATE_REG_SCAN_IN), .B2(n2961), .A(n2960), .ZN(U3326)
         );
  INV_X1 U3786 ( .A(DATAI_29_), .ZN(n2964) );
  NAND2_X1 U3787 ( .A1(n2962), .A2(STATE_REG_SCAN_IN), .ZN(n2963) );
  OAI21_X1 U3788 ( .B1(STATE_REG_SCAN_IN), .B2(n2964), .A(n2963), .ZN(U3323)
         );
  INV_X1 U3789 ( .A(n2988), .ZN(n2966) );
  NOR3_X1 U3790 ( .A1(n2968), .A2(n2967), .A3(n4340), .ZN(n2969) );
  AOI21_X1 U3791 ( .B1(n4464), .B2(n2970), .A(n2969), .ZN(U3458) );
  INV_X1 U3792 ( .A(D_REG_1__SCAN_IN), .ZN(n2972) );
  AOI22_X1 U3793 ( .A1(n4464), .A2(n2972), .B1(n2971), .B2(n4466), .ZN(U3459)
         );
  INV_X1 U3794 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n2978) );
  NAND2_X1 U3795 ( .A1(n3605), .A2(REG1_REG_30__SCAN_IN), .ZN(n2976) );
  NAND2_X1 U3796 ( .A1(n3606), .A2(REG2_REG_30__SCAN_IN), .ZN(n2975) );
  NAND2_X1 U3797 ( .A1(n2973), .A2(REG0_REG_30__SCAN_IN), .ZN(n2974) );
  NAND3_X1 U3798 ( .A1(n2976), .A2(n2975), .A3(n2974), .ZN(n3896) );
  NAND2_X1 U3799 ( .A1(n3896), .A2(U4043), .ZN(n2977) );
  OAI21_X1 U3800 ( .B1(U4043), .B2(n2978), .A(n2977), .ZN(U3580) );
  INV_X1 U3801 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n2980) );
  NAND2_X1 U3802 ( .A1(n3288), .A2(U4043), .ZN(n2979) );
  OAI21_X1 U3803 ( .B1(U4043), .B2(n2980), .A(n2979), .ZN(U3556) );
  INV_X1 U3804 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n2982) );
  NAND2_X1 U3805 ( .A1(n3213), .A2(U4043), .ZN(n2981) );
  OAI21_X1 U3806 ( .B1(U4043), .B2(n2982), .A(n2981), .ZN(U3553) );
  INV_X1 U3807 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n2984) );
  NAND2_X1 U3808 ( .A1(n4031), .A2(U4043), .ZN(n2983) );
  OAI21_X1 U3809 ( .B1(U4043), .B2(n2984), .A(n2983), .ZN(U3570) );
  NAND2_X1 U3810 ( .A1(n2987), .A2(n2985), .ZN(n2986) );
  OR2_X1 U3811 ( .A1(n2987), .A2(U3149), .ZN(n3769) );
  NAND2_X1 U3812 ( .A1(n2988), .A2(n3769), .ZN(n3002) );
  AND2_X1 U3813 ( .A1(n3044), .A2(n4351), .ZN(n4412) );
  XNOR2_X1 U3814 ( .A(n2989), .B(IR_REG_27__SCAN_IN), .ZN(n4338) );
  INV_X1 U3815 ( .A(n4338), .ZN(n3794) );
  INV_X1 U3816 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2994) );
  MUX2_X1 U3817 ( .A(REG1_REG_2__SCAN_IN), .B(n2994), .S(n3807), .Z(n2993) );
  INV_X1 U3818 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2990) );
  AND2_X1 U3819 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n2991)
         );
  NAND2_X1 U3820 ( .A1(n4349), .A2(REG1_REG_1__SCAN_IN), .ZN(n3801) );
  NAND2_X1 U3821 ( .A1(n3800), .A2(n3801), .ZN(n2992) );
  XOR2_X1 U3822 ( .A(REG1_REG_3__SCAN_IN), .B(n3017), .Z(n3001) );
  NOR2_X1 U3823 ( .A1(n3794), .A2(n4351), .ZN(n3765) );
  INV_X1 U3824 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2999) );
  MUX2_X1 U3825 ( .A(REG2_REG_2__SCAN_IN), .B(n2999), .S(n3807), .Z(n2997) );
  INV_X1 U3826 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2995) );
  MUX2_X1 U3827 ( .A(REG2_REG_1__SCAN_IN), .B(n2995), .S(n4349), .Z(n3785) );
  AND2_X1 U3828 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3793)
         );
  NAND2_X1 U3829 ( .A1(n3785), .A2(n3793), .ZN(n3808) );
  NAND2_X1 U3830 ( .A1(n4349), .A2(REG2_REG_1__SCAN_IN), .ZN(n3809) );
  NAND2_X1 U3831 ( .A1(n3808), .A2(n3809), .ZN(n2996) );
  XOR2_X1 U3832 ( .A(REG2_REG_3__SCAN_IN), .B(n3010), .Z(n3000) );
  AOI22_X1 U3833 ( .A1(n4437), .A2(n3001), .B1(n4439), .B2(n3000), .ZN(n3006)
         );
  INV_X1 U3834 ( .A(n3002), .ZN(n3004) );
  INV_X1 U3835 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3151) );
  NOR2_X1 U3836 ( .A1(STATE_REG_SCAN_IN), .A2(n3151), .ZN(n3132) );
  AOI21_X1 U3837 ( .B1(n4429), .B2(ADDR_REG_3__SCAN_IN), .A(n3132), .ZN(n3005)
         );
  OAI211_X1 U3838 ( .C1(n2165), .C2(n4442), .A(n3006), .B(n3005), .ZN(U3243)
         );
  INV_X1 U3839 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n3009) );
  NAND2_X1 U3840 ( .A1(n3007), .A2(U4043), .ZN(n3008) );
  OAI21_X1 U3841 ( .B1(U4043), .B2(n3009), .A(n3008), .ZN(U3561) );
  INV_X1 U3842 ( .A(n3062), .ZN(n4346) );
  XNOR2_X1 U3843 ( .A(n3011), .B(n4347), .ZN(n3818) );
  INV_X1 U3844 ( .A(n3011), .ZN(n3012) );
  INV_X1 U3845 ( .A(REG2_REG_5__SCAN_IN), .ZN(n4601) );
  MUX2_X1 U3846 ( .A(REG2_REG_5__SCAN_IN), .B(n4601), .S(n3062), .Z(n3052) );
  INV_X1 U3847 ( .A(n3013), .ZN(n3014) );
  AOI22_X1 U3848 ( .A1(n3074), .A2(REG2_REG_6__SCAN_IN), .B1(n4345), .B2(n3014), .ZN(n3069) );
  INV_X1 U3849 ( .A(REG2_REG_7__SCAN_IN), .ZN(n4600) );
  MUX2_X1 U3850 ( .A(n4600), .B(REG2_REG_7__SCAN_IN), .S(n4344), .Z(n3068) );
  XOR2_X1 U3851 ( .A(REG2_REG_8__SCAN_IN), .B(n3031), .Z(n3025) );
  NAND2_X1 U3852 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3299) );
  INV_X1 U3853 ( .A(n3299), .ZN(n3016) );
  NOR2_X1 U3854 ( .A1(n4442), .A2(n3037), .ZN(n3015) );
  AOI211_X1 U3855 ( .C1(n4429), .C2(ADDR_REG_8__SCAN_IN), .A(n3016), .B(n3015), 
        .ZN(n3024) );
  INV_X1 U3856 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4598) );
  INV_X1 U3857 ( .A(n4344), .ZN(n3066) );
  XNOR2_X1 U3858 ( .A(n3018), .B(n4347), .ZN(n3817) );
  INV_X1 U3859 ( .A(n3018), .ZN(n3019) );
  INV_X1 U3860 ( .A(REG1_REG_5__SCAN_IN), .ZN(n4525) );
  MUX2_X1 U3861 ( .A(REG1_REG_5__SCAN_IN), .B(n4525), .S(n3062), .Z(n3055) );
  INV_X1 U3862 ( .A(n3020), .ZN(n3021) );
  OAI211_X1 U3863 ( .C1(n3022), .C2(REG1_REG_8__SCAN_IN), .A(n3036), .B(n4437), 
        .ZN(n3023) );
  OAI211_X1 U3864 ( .C1(n3025), .C2(n4405), .A(n3024), .B(n3023), .ZN(U3248)
         );
  INV_X1 U3865 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n3027) );
  NAND2_X1 U3866 ( .A1(n3937), .A2(U4043), .ZN(n3026) );
  OAI21_X1 U3867 ( .B1(U4043), .B2(n3027), .A(n3026), .ZN(U3577) );
  NOR2_X1 U3868 ( .A1(n4429), .A2(U4043), .ZN(U3148) );
  INV_X1 U3869 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n3029) );
  NAND2_X1 U3870 ( .A1(n3535), .A2(U4043), .ZN(n3028) );
  OAI21_X1 U3871 ( .B1(U4043), .B2(n3029), .A(n3028), .ZN(U3575) );
  INV_X1 U3872 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4604) );
  AOI22_X1 U3873 ( .A1(n3039), .A2(REG2_REG_9__SCAN_IN), .B1(n4604), .B2(n4478), .ZN(n4366) );
  INV_X1 U3874 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3030) );
  NAND2_X1 U3875 ( .A1(n4366), .A2(n4365), .ZN(n4364) );
  OAI211_X1 U3876 ( .C1(n3032), .C2(REG2_REG_10__SCAN_IN), .A(n4439), .B(n3832), .ZN(n3035) );
  NAND2_X1 U3877 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n3348) );
  INV_X1 U3878 ( .A(n3348), .ZN(n3033) );
  AOI21_X1 U3879 ( .B1(n4429), .B2(ADDR_REG_10__SCAN_IN), .A(n3033), .ZN(n3034) );
  OAI211_X1 U3880 ( .C1(n4442), .C2(n2169), .A(n3035), .B(n3034), .ZN(n3042)
         );
  INV_X1 U3881 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3441) );
  INV_X1 U3882 ( .A(REG1_REG_9__SCAN_IN), .ZN(n4528) );
  AOI22_X1 U3883 ( .A1(n3039), .A2(n4528), .B1(REG1_REG_9__SCAN_IN), .B2(n4478), .ZN(n4360) );
  AOI211_X1 U3884 ( .C1(n3441), .C2(n3040), .A(n3844), .B(n4401), .ZN(n3041)
         );
  OR2_X1 U3885 ( .A1(n3042), .A2(n3041), .ZN(U3250) );
  INV_X1 U3886 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3047) );
  AOI21_X1 U3887 ( .B1(n4338), .B2(n2281), .A(n4351), .ZN(n3799) );
  NOR2_X1 U3888 ( .A1(n4338), .A2(REG1_REG_0__SCAN_IN), .ZN(n3043) );
  OAI21_X1 U3889 ( .B1(IR_REG_0__SCAN_IN), .B2(n3043), .A(n3799), .ZN(n3045)
         );
  OAI211_X1 U3890 ( .C1(n3799), .C2(IR_REG_0__SCAN_IN), .A(n3045), .B(n3044), 
        .ZN(n3046) );
  OAI21_X1 U3891 ( .B1(STATE_REG_SCAN_IN), .B2(n3047), .A(n3046), .ZN(n3049)
         );
  NOR3_X1 U3892 ( .A1(n4401), .A2(REG1_REG_0__SCAN_IN), .A3(n2146), .ZN(n3048)
         );
  AOI211_X1 U3893 ( .C1(n4429), .C2(ADDR_REG_0__SCAN_IN), .A(n3049), .B(n3048), 
        .ZN(n3050) );
  INV_X1 U3894 ( .A(n3050), .ZN(U3240) );
  AOI211_X1 U3895 ( .C1(n3053), .C2(n3052), .A(n3051), .B(n4405), .ZN(n3058)
         );
  AOI211_X1 U3896 ( .C1(n3056), .C2(n3055), .A(n3054), .B(n4401), .ZN(n3057)
         );
  NOR2_X1 U3897 ( .A1(n3058), .A2(n3057), .ZN(n3061) );
  NOR2_X1 U3898 ( .A1(n3059), .A2(STATE_REG_SCAN_IN), .ZN(n3166) );
  AOI21_X1 U3899 ( .B1(n4429), .B2(ADDR_REG_5__SCAN_IN), .A(n3166), .ZN(n3060)
         );
  OAI211_X1 U3900 ( .C1(n3062), .C2(n4442), .A(n3061), .B(n3060), .ZN(U3245)
         );
  XNOR2_X1 U3901 ( .A(n4344), .B(n4598), .ZN(n3063) );
  XNOR2_X1 U3902 ( .A(n3064), .B(n3063), .ZN(n3072) );
  NAND2_X1 U3903 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3290) );
  NAND2_X1 U3904 ( .A1(n4429), .A2(ADDR_REG_7__SCAN_IN), .ZN(n3065) );
  OAI211_X1 U3905 ( .C1(n4442), .C2(n3066), .A(n3290), .B(n3065), .ZN(n3071)
         );
  AOI211_X1 U3906 ( .C1(n3069), .C2(n3068), .A(n4405), .B(n3067), .ZN(n3070)
         );
  AOI211_X1 U3907 ( .C1(n3072), .C2(n4437), .A(n3071), .B(n3070), .ZN(n3073)
         );
  INV_X1 U3908 ( .A(n3073), .ZN(U3247) );
  XNOR2_X1 U3909 ( .A(n3074), .B(REG2_REG_6__SCAN_IN), .ZN(n3081) );
  XOR2_X1 U3910 ( .A(REG1_REG_6__SCAN_IN), .B(n3075), .Z(n3079) );
  INV_X1 U3911 ( .A(REG3_REG_6__SCAN_IN), .ZN(n4659) );
  NOR2_X1 U3912 ( .A1(STATE_REG_SCAN_IN), .A2(n4659), .ZN(n3307) );
  AOI21_X1 U3913 ( .B1(n4429), .B2(ADDR_REG_6__SCAN_IN), .A(n3307), .ZN(n3076)
         );
  OAI21_X1 U3914 ( .B1(n4442), .B2(n3077), .A(n3076), .ZN(n3078) );
  AOI21_X1 U3915 ( .B1(n4437), .B2(n3079), .A(n3078), .ZN(n3080) );
  OAI21_X1 U3916 ( .B1(n3081), .B2(n4405), .A(n3080), .ZN(U3246) );
  OAI21_X1 U3917 ( .B1(n3084), .B2(n3083), .A(n3082), .ZN(n3797) );
  OAI22_X1 U3918 ( .A1(n3797), .A2(n3599), .B1(n3583), .B2(n4453), .ZN(n3090)
         );
  NAND3_X1 U3919 ( .A1(n3086), .A2(n3085), .A3(n3109), .ZN(n3105) );
  INV_X1 U3920 ( .A(n3105), .ZN(n3088) );
  OAI22_X1 U3921 ( .A1(n3088), .A2(n3047), .B1(n3087), .B2(n3593), .ZN(n3089)
         );
  OR2_X1 U3922 ( .A1(n3090), .A2(n3089), .ZN(U3229) );
  OAI211_X1 U3923 ( .C1(n3091), .C2(n3093), .A(n3092), .B(n3563), .ZN(n3097)
         );
  OAI22_X1 U3924 ( .A1(n3094), .A2(n3581), .B1(n2822), .B2(n3593), .ZN(n3095)
         );
  AOI21_X1 U3925 ( .B1(REG3_REG_1__SCAN_IN), .B2(n3105), .A(n3095), .ZN(n3096)
         );
  OAI211_X1 U3926 ( .C1(n3583), .C2(n3112), .A(n3097), .B(n3096), .ZN(U3219)
         );
  INV_X1 U3927 ( .A(n3100), .ZN(n3101) );
  AOI21_X1 U3928 ( .B1(n3098), .B2(n3099), .A(n3101), .ZN(n3107) );
  OAI22_X1 U3929 ( .A1(n3178), .A2(n3593), .B1(n3087), .B2(n3581), .ZN(n3104)
         );
  NOR2_X1 U3930 ( .A1(n3583), .A2(n3102), .ZN(n3103) );
  AOI211_X1 U3931 ( .C1(REG3_REG_2__SCAN_IN), .C2(n3105), .A(n3104), .B(n3103), 
        .ZN(n3106) );
  OAI21_X1 U3932 ( .B1(n3107), .B2(n3599), .A(n3106), .ZN(U3234) );
  NAND3_X1 U3933 ( .A1(n3110), .A2(n3109), .A3(n3108), .ZN(n3111) );
  OAI21_X1 U3934 ( .B1(n4453), .B2(n3112), .A(n3185), .ZN(n4479) );
  OR2_X1 U3935 ( .A1(n3113), .A2(n3114), .ZN(n3115) );
  NAND2_X1 U3936 ( .A1(n3116), .A2(n3115), .ZN(n4481) );
  NAND2_X1 U3937 ( .A1(n3117), .A2(n4450), .ZN(n3119) );
  NAND2_X1 U3938 ( .A1(n3784), .A2(n4159), .ZN(n3118) );
  OAI211_X1 U3939 ( .C1(n2822), .C2(n4155), .A(n3119), .B(n3118), .ZN(n3120)
         );
  INV_X1 U3940 ( .A(n3120), .ZN(n3123) );
  XNOR2_X1 U3941 ( .A(n3113), .B(n3730), .ZN(n3121) );
  NAND2_X1 U3942 ( .A1(n3121), .A2(n4281), .ZN(n3122) );
  OAI211_X1 U3943 ( .C1(n4481), .C2(n4455), .A(n3123), .B(n3122), .ZN(n4483)
         );
  MUX2_X1 U3944 ( .A(n4483), .B(REG2_REG_1__SCAN_IN), .S(n2017), .Z(n3124) );
  INV_X1 U3945 ( .A(n3124), .ZN(n3129) );
  INV_X1 U3946 ( .A(n4481), .ZN(n3127) );
  OR2_X1 U3947 ( .A1(n3125), .A2(n4451), .ZN(n3192) );
  INV_X1 U3948 ( .A(n3192), .ZN(n3126) );
  AND2_X1 U3949 ( .A1(n4195), .A2(n3126), .ZN(n4460) );
  AOI22_X1 U3950 ( .A1(n3127), .A2(n4460), .B1(REG3_REG_1__SCAN_IN), .B2(n4459), .ZN(n3128) );
  OAI211_X1 U3951 ( .C1(n4169), .C2(n4479), .A(n3129), .B(n3128), .ZN(U3289)
         );
  XNOR2_X1 U3952 ( .A(n3131), .B(n3130), .ZN(n3137) );
  NOR2_X1 U3953 ( .A1(n3557), .A2(REG3_REG_3__SCAN_IN), .ZN(n3136) );
  AOI21_X1 U3954 ( .B1(n3782), .B2(n3589), .A(n3132), .ZN(n3134) );
  NAND2_X1 U3955 ( .A1(n3590), .A2(n3142), .ZN(n3133) );
  OAI211_X1 U3956 ( .C1(n2825), .C2(n3593), .A(n3134), .B(n3133), .ZN(n3135)
         );
  AOI211_X1 U3957 ( .C1(n3137), .C2(n3563), .A(n3136), .B(n3135), .ZN(n3138)
         );
  INV_X1 U3958 ( .A(n3138), .ZN(U3215) );
  INV_X1 U3959 ( .A(n3746), .ZN(n3140) );
  XNOR2_X1 U3960 ( .A(n3139), .B(n3140), .ZN(n4487) );
  INV_X1 U3961 ( .A(n4455), .ZN(n3425) );
  NAND2_X1 U3962 ( .A1(n4487), .A2(n3425), .ZN(n3148) );
  XNOR2_X1 U3963 ( .A(n3141), .B(n3746), .ZN(n3146) );
  OR2_X1 U3964 ( .A1(n2822), .A2(n4184), .ZN(n3144) );
  NAND2_X1 U3965 ( .A1(n3142), .A2(n4450), .ZN(n3143) );
  OAI211_X1 U3966 ( .C1(n2825), .C2(n4155), .A(n3144), .B(n3143), .ZN(n3145)
         );
  AOI21_X1 U3967 ( .B1(n3146), .B2(n4281), .A(n3145), .ZN(n3147) );
  AND2_X1 U3968 ( .A1(n3148), .A2(n3147), .ZN(n4489) );
  OR2_X1 U3969 ( .A1(n3184), .A2(n3149), .ZN(n3150) );
  AOI22_X1 U3970 ( .A1(n2017), .A2(REG2_REG_3__SCAN_IN), .B1(n4459), .B2(n3151), .ZN(n3152) );
  OAI21_X1 U3971 ( .B1(n4169), .B2(n4485), .A(n3152), .ZN(n3153) );
  AOI21_X1 U3972 ( .B1(n4487), .B2(n4460), .A(n3153), .ZN(n3154) );
  OAI21_X1 U3973 ( .B1(n4489), .B2(n2017), .A(n3154), .ZN(U3287) );
  AOI21_X1 U3974 ( .B1(n3156), .B2(n3155), .A(n3599), .ZN(n3158) );
  NAND2_X1 U3975 ( .A1(n3158), .A2(n3157), .ZN(n3162) );
  NAND2_X1 U3976 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3816) );
  NAND2_X1 U3977 ( .A1(n3589), .A2(n3213), .ZN(n3159) );
  OAI211_X1 U3978 ( .C1(n2828), .C2(n3593), .A(n3816), .B(n3159), .ZN(n3160)
         );
  AOI21_X1 U3979 ( .B1(n3212), .B2(n3590), .A(n3160), .ZN(n3161) );
  OAI211_X1 U3980 ( .C1(n3557), .C2(n3221), .A(n3162), .B(n3161), .ZN(U3227)
         );
  INV_X1 U3981 ( .A(n3206), .ZN(n3171) );
  OAI211_X1 U3982 ( .C1(n3165), .C2(n3164), .A(n3163), .B(n3563), .ZN(n3170)
         );
  AOI21_X1 U3983 ( .B1(n3579), .B2(n3288), .A(n3166), .ZN(n3167) );
  OAI21_X1 U3984 ( .B1(n2825), .B2(n3581), .A(n3167), .ZN(n3168) );
  AOI21_X1 U3985 ( .B1(n3204), .B2(n3590), .A(n3168), .ZN(n3169) );
  OAI211_X1 U3986 ( .C1(n3557), .C2(n3171), .A(n3170), .B(n3169), .ZN(U3224)
         );
  INV_X1 U3987 ( .A(n3172), .ZN(n3173) );
  AOI21_X1 U3988 ( .B1(n3708), .B2(n3174), .A(n3173), .ZN(n3179) );
  INV_X1 U3989 ( .A(n3179), .ZN(n4445) );
  OAI21_X1 U3990 ( .B1(n3708), .B2(n3176), .A(n3175), .ZN(n3182) );
  AOI22_X1 U3991 ( .A1(n4279), .A2(n4159), .B1(n3186), .B2(n4450), .ZN(n3177)
         );
  OAI21_X1 U3992 ( .B1(n3178), .B2(n4155), .A(n3177), .ZN(n3181) );
  NOR2_X1 U3993 ( .A1(n3179), .A2(n4455), .ZN(n3180) );
  AOI211_X1 U3994 ( .C1(n4281), .C2(n3182), .A(n3181), .B(n3180), .ZN(n4448)
         );
  INV_X1 U3995 ( .A(n4448), .ZN(n3183) );
  AOI21_X1 U3996 ( .B1(n4520), .B2(n4445), .A(n3183), .ZN(n3191) );
  AOI21_X1 U3997 ( .B1(n3186), .B2(n3185), .A(n3184), .ZN(n4443) );
  INV_X1 U3998 ( .A(n4335), .ZN(n3187) );
  AOI22_X1 U3999 ( .A1(n4443), .A2(n3187), .B1(n4690), .B2(REG0_REG_2__SCAN_IN), .ZN(n3188) );
  OAI21_X1 U4000 ( .B1(n3191), .B2(n4690), .A(n3188), .ZN(U3471) );
  INV_X1 U4001 ( .A(n4278), .ZN(n3189) );
  AOI22_X1 U4002 ( .A1(n4443), .A2(n3189), .B1(n4530), .B2(REG1_REG_2__SCAN_IN), .ZN(n3190) );
  OAI21_X1 U4003 ( .B1(n3191), .B2(n4530), .A(n3190), .ZN(U3520) );
  NAND2_X1 U4004 ( .A1(n4455), .A2(n3192), .ZN(n3193) );
  NAND2_X1 U4005 ( .A1(n3195), .A2(n3194), .ZN(n3255) );
  OR2_X1 U4006 ( .A1(n3255), .A2(n3709), .ZN(n3210) );
  NAND2_X1 U4007 ( .A1(n3210), .A2(n3197), .ZN(n3199) );
  INV_X1 U4008 ( .A(n3198), .ZN(n3652) );
  NAND2_X1 U4009 ( .A1(n3652), .A2(n3663), .ZN(n3722) );
  XNOR2_X1 U4010 ( .A(n3199), .B(n3722), .ZN(n4497) );
  XNOR2_X1 U4011 ( .A(n3200), .B(n3722), .ZN(n3203) );
  AOI22_X1 U4012 ( .A1(n3288), .A2(n4280), .B1(n4450), .B2(n3204), .ZN(n3201)
         );
  OAI21_X1 U4013 ( .B1(n2825), .B2(n4184), .A(n3201), .ZN(n3202) );
  AOI21_X1 U4014 ( .B1(n3203), .B2(n4281), .A(n3202), .ZN(n4498) );
  MUX2_X1 U4015 ( .A(n4498), .B(n4601), .S(n2017), .Z(n3208) );
  AND2_X1 U4016 ( .A1(n3218), .A2(n3204), .ZN(n3205) );
  NOR2_X1 U4017 ( .A1(n3249), .A2(n3205), .ZN(n4501) );
  AOI22_X1 U4018 ( .A1(n4501), .A2(n4444), .B1(n3206), .B2(n4459), .ZN(n3207)
         );
  OAI211_X1 U4019 ( .C1(n4172), .C2(n4497), .A(n3208), .B(n3207), .ZN(U3285)
         );
  NAND2_X1 U4020 ( .A1(n3255), .A2(n3709), .ZN(n3209) );
  AND2_X1 U4021 ( .A1(n3210), .A2(n3209), .ZN(n4494) );
  INV_X1 U4022 ( .A(n4494), .ZN(n3225) );
  INV_X1 U4023 ( .A(n4460), .ZN(n4200) );
  XOR2_X1 U4024 ( .A(n3211), .B(n3709), .Z(n3217) );
  AOI22_X1 U4025 ( .A1(n3213), .A2(n4159), .B1(n3212), .B2(n4450), .ZN(n3214)
         );
  OAI21_X1 U4026 ( .B1(n2828), .B2(n4155), .A(n3214), .ZN(n3215) );
  AOI21_X1 U4027 ( .B1(n4494), .B2(n3425), .A(n3215), .ZN(n3216) );
  OAI21_X1 U4028 ( .B1(n4161), .B2(n3217), .A(n3216), .ZN(n4492) );
  OAI211_X1 U4029 ( .C1(n3220), .C2(n3219), .A(n4502), .B(n3218), .ZN(n4491)
         );
  OAI22_X1 U4030 ( .A1(n4491), .A2(n4342), .B1(n4193), .B2(n3221), .ZN(n3222)
         );
  OAI21_X1 U4031 ( .B1(n4492), .B2(n3222), .A(n4195), .ZN(n3224) );
  NAND2_X1 U4032 ( .A1(n2017), .A2(REG2_REG_4__SCAN_IN), .ZN(n3223) );
  OAI211_X1 U4033 ( .C1(n3225), .C2(n4200), .A(n3224), .B(n3223), .ZN(U3286)
         );
  INV_X1 U4034 ( .A(n3240), .ZN(n3711) );
  XNOR2_X1 U4035 ( .A(n3226), .B(n3711), .ZN(n3230) );
  NAND2_X1 U4036 ( .A1(n3292), .A2(n4450), .ZN(n3228) );
  NAND2_X1 U4037 ( .A1(n3288), .A2(n4159), .ZN(n3227) );
  OAI211_X1 U4038 ( .C1(n3360), .C2(n4155), .A(n3228), .B(n3227), .ZN(n3229)
         );
  AOI21_X1 U4039 ( .B1(n3230), .B2(n4281), .A(n3229), .ZN(n4508) );
  OAI211_X1 U4040 ( .C1(n3251), .C2(n3231), .A(n4502), .B(n3280), .ZN(n4506)
         );
  INV_X1 U4041 ( .A(n4506), .ZN(n3234) );
  INV_X1 U4042 ( .A(n3232), .ZN(n3295) );
  OAI22_X1 U40430 ( .A1(n4195), .A2(n4600), .B1(n3295), .B2(n4193), .ZN(n3233)
         );
  AOI21_X1 U4044 ( .B1(n3234), .B2(n4096), .A(n3233), .ZN(n3243) );
  INV_X1 U4045 ( .A(n3235), .ZN(n3236) );
  OR2_X1 U4046 ( .A1(n3254), .A2(n3236), .ZN(n3237) );
  OR2_X1 U4047 ( .A1(n3255), .A2(n3237), .ZN(n3239) );
  NAND2_X1 U4048 ( .A1(n3239), .A2(n3238), .ZN(n3241) );
  OR2_X1 U4049 ( .A1(n3241), .A2(n3240), .ZN(n4505) );
  NAND2_X1 U4050 ( .A1(n3241), .A2(n3240), .ZN(n4504) );
  NAND3_X1 U4051 ( .A1(n4505), .A2(n3920), .A3(n4504), .ZN(n3242) );
  OAI211_X1 U4052 ( .C1(n4508), .C2(n2017), .A(n3243), .B(n3242), .ZN(U3283)
         );
  AND2_X1 U4053 ( .A1(n3655), .A2(n3664), .ZN(n3749) );
  XNOR2_X1 U4054 ( .A(n3244), .B(n3749), .ZN(n3247) );
  NOR2_X1 U4055 ( .A1(n2828), .A2(n4184), .ZN(n3246) );
  OAI22_X1 U4056 ( .A1(n2833), .A2(n4155), .B1(n4154), .B2(n3248), .ZN(n3245)
         );
  AOI211_X1 U4057 ( .C1(n3247), .C2(n4281), .A(n3246), .B(n3245), .ZN(n3263)
         );
  NOR2_X1 U4058 ( .A1(n3249), .A2(n3248), .ZN(n3250) );
  OR2_X1 U4059 ( .A1(n3251), .A2(n3250), .ZN(n3269) );
  INV_X1 U4060 ( .A(n3269), .ZN(n3261) );
  INV_X1 U4061 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3253) );
  INV_X1 U4062 ( .A(n3318), .ZN(n3252) );
  OAI22_X1 U4063 ( .A1(n4195), .A2(n3253), .B1(n3252), .B2(n4193), .ZN(n3260)
         );
  OR2_X1 U4064 ( .A1(n3255), .A2(n3254), .ZN(n3257) );
  NAND2_X1 U4065 ( .A1(n3257), .A2(n3256), .ZN(n3258) );
  XOR2_X1 U4066 ( .A(n3749), .B(n3258), .Z(n3264) );
  NOR2_X1 U4067 ( .A1(n3264), .A2(n4172), .ZN(n3259) );
  AOI211_X1 U4068 ( .C1(n3261), .C2(n4444), .A(n3260), .B(n3259), .ZN(n3262)
         );
  OAI21_X1 U4069 ( .B1(n2017), .B2(n3263), .A(n3262), .ZN(U3284) );
  OAI21_X1 U4070 ( .B1(n3264), .B2(n4496), .A(n3263), .ZN(n3271) );
  INV_X1 U4071 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3265) );
  OAI22_X1 U4072 ( .A1(n3269), .A2(n4278), .B1(n4533), .B2(n3265), .ZN(n3266)
         );
  AOI21_X1 U4073 ( .B1(n3271), .B2(n4533), .A(n3266), .ZN(n3267) );
  INV_X1 U4074 ( .A(n3267), .ZN(U3524) );
  INV_X1 U4075 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3268) );
  OAI22_X1 U4076 ( .A1(n3269), .A2(n4335), .B1(n4692), .B2(n3268), .ZN(n3270)
         );
  AOI21_X1 U4077 ( .B1(n3271), .B2(n4692), .A(n3270), .ZN(n3272) );
  INV_X1 U4078 ( .A(n3272), .ZN(U3479) );
  NAND2_X1 U4079 ( .A1(n3659), .A2(n3657), .ZN(n3721) );
  XNOR2_X1 U4080 ( .A(n3273), .B(n3721), .ZN(n3276) );
  AOI22_X1 U4081 ( .A1(n3777), .A2(n4280), .B1(n4450), .B2(n3279), .ZN(n3274)
         );
  OAI21_X1 U4082 ( .B1(n2833), .B2(n4184), .A(n3274), .ZN(n3275) );
  AOI21_X1 U4083 ( .B1(n3276), .B2(n4281), .A(n3275), .ZN(n3335) );
  INV_X1 U4084 ( .A(n3721), .ZN(n3278) );
  XNOR2_X1 U4085 ( .A(n3277), .B(n3278), .ZN(n3333) );
  NAND2_X1 U4086 ( .A1(n3280), .A2(n3279), .ZN(n3281) );
  NAND2_X1 U4087 ( .A1(n3327), .A2(n3281), .ZN(n3340) );
  AOI22_X1 U4088 ( .A1(n2017), .A2(REG2_REG_8__SCAN_IN), .B1(n3304), .B2(n4459), .ZN(n3282) );
  OAI21_X1 U4089 ( .B1(n3340), .B2(n4169), .A(n3282), .ZN(n3283) );
  AOI21_X1 U4090 ( .B1(n3333), .B2(n3920), .A(n3283), .ZN(n3284) );
  OAI21_X1 U4091 ( .B1(n3335), .B2(n2017), .A(n3284), .ZN(U3282) );
  XOR2_X1 U4092 ( .A(n3285), .B(n3286), .Z(n3287) );
  NAND2_X1 U4093 ( .A1(n3287), .A2(n3563), .ZN(n3294) );
  NAND2_X1 U4094 ( .A1(n3589), .A2(n3288), .ZN(n3289) );
  OAI211_X1 U4095 ( .C1(n3360), .C2(n3593), .A(n3290), .B(n3289), .ZN(n3291)
         );
  AOI21_X1 U4096 ( .B1(n3292), .B2(n3590), .A(n3291), .ZN(n3293) );
  OAI211_X1 U4097 ( .C1(n3557), .C2(n3295), .A(n3294), .B(n3293), .ZN(U3210)
         );
  INV_X1 U4098 ( .A(n3355), .ZN(n3297) );
  NOR2_X1 U4099 ( .A1(n3297), .A2(n3354), .ZN(n3298) );
  XNOR2_X1 U4100 ( .A(n3296), .B(n3298), .ZN(n3306) );
  OAI21_X1 U4101 ( .B1(n2833), .B2(n3581), .A(n3299), .ZN(n3300) );
  AOI21_X1 U4102 ( .B1(n3579), .B2(n3777), .A(n3300), .ZN(n3301) );
  OAI21_X1 U4103 ( .B1(n3583), .B2(n3302), .A(n3301), .ZN(n3303) );
  AOI21_X1 U4104 ( .B1(n3304), .B2(n3603), .A(n3303), .ZN(n3305) );
  OAI21_X1 U4105 ( .B1(n3306), .B2(n3599), .A(n3305), .ZN(U3218) );
  AOI21_X1 U4106 ( .B1(n3780), .B2(n3589), .A(n3307), .ZN(n3310) );
  NAND2_X1 U4107 ( .A1(n3590), .A2(n3308), .ZN(n3309) );
  OAI211_X1 U4108 ( .C1(n2833), .C2(n3593), .A(n3310), .B(n3309), .ZN(n3317)
         );
  XOR2_X1 U4109 ( .A(n3312), .B(n3311), .Z(n3313) );
  XNOR2_X1 U4110 ( .A(n3314), .B(n3313), .ZN(n3315) );
  NOR2_X1 U4111 ( .A1(n3315), .A2(n3599), .ZN(n3316) );
  AOI211_X1 U4112 ( .C1(n3318), .C2(n3603), .A(n3317), .B(n3316), .ZN(n3319)
         );
  INV_X1 U4113 ( .A(n3319), .ZN(U3236) );
  INV_X1 U4114 ( .A(n3320), .ZN(n3674) );
  NAND2_X1 U4115 ( .A1(n3674), .A2(n3660), .ZN(n3720) );
  XNOR2_X1 U4116 ( .A(n3321), .B(n3720), .ZN(n3325) );
  AOI22_X1 U4117 ( .A1(n3776), .A2(n4280), .B1(n4450), .B2(n3322), .ZN(n3323)
         );
  OAI21_X1 U4118 ( .B1(n3360), .B2(n4184), .A(n3323), .ZN(n3324) );
  AOI21_X1 U4119 ( .B1(n3325), .B2(n4281), .A(n3324), .ZN(n4510) );
  XOR2_X1 U4120 ( .A(n3326), .B(n3720), .Z(n4514) );
  INV_X1 U4121 ( .A(n3327), .ZN(n3329) );
  INV_X1 U4122 ( .A(n3383), .ZN(n3328) );
  OAI21_X1 U4123 ( .B1(n3329), .B2(n2150), .A(n3328), .ZN(n4511) );
  AOI22_X1 U4124 ( .A1(n2017), .A2(REG2_REG_9__SCAN_IN), .B1(n3364), .B2(n4459), .ZN(n3330) );
  OAI21_X1 U4125 ( .B1(n4511), .B2(n4169), .A(n3330), .ZN(n3331) );
  AOI21_X1 U4126 ( .B1(n4514), .B2(n3920), .A(n3331), .ZN(n3332) );
  OAI21_X1 U4127 ( .B1(n2017), .B2(n4510), .A(n3332), .ZN(U3281) );
  NAND2_X1 U4128 ( .A1(n3333), .A2(n4513), .ZN(n3334) );
  AND2_X1 U4129 ( .A1(n3335), .A2(n3334), .ZN(n3338) );
  INV_X1 U4130 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3336) );
  MUX2_X1 U4131 ( .A(n3338), .B(n3336), .S(n4690), .Z(n3337) );
  OAI21_X1 U4132 ( .B1(n3340), .B2(n4335), .A(n3337), .ZN(U3483) );
  INV_X1 U4133 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4614) );
  MUX2_X1 U4134 ( .A(n4614), .B(n3338), .S(n4533), .Z(n3339) );
  OAI21_X1 U4135 ( .B1(n3340), .B2(n4278), .A(n3339), .ZN(U3526) );
  INV_X1 U4136 ( .A(n3385), .ZN(n3353) );
  NAND2_X1 U4137 ( .A1(n3341), .A2(n3342), .ZN(n3344) );
  AOI21_X1 U4138 ( .B1(n3344), .B2(n3343), .A(n3599), .ZN(n3346) );
  NAND2_X1 U4139 ( .A1(n3346), .A2(n3345), .ZN(n3352) );
  NAND2_X1 U4140 ( .A1(n3589), .A2(n3777), .ZN(n3347) );
  OAI211_X1 U4141 ( .C1(n3402), .C2(n3593), .A(n3348), .B(n3347), .ZN(n3349)
         );
  AOI21_X1 U4142 ( .B1(n3350), .B2(n3590), .A(n3349), .ZN(n3351) );
  OAI211_X1 U4143 ( .C1(n3557), .C2(n3353), .A(n3352), .B(n3351), .ZN(U3214)
         );
  OR2_X1 U4144 ( .A1(n3296), .A2(n3354), .ZN(n3356) );
  NAND2_X1 U4145 ( .A1(n3356), .A2(n3355), .ZN(n3357) );
  XOR2_X1 U4146 ( .A(n3358), .B(n3357), .Z(n3366) );
  NOR2_X1 U4147 ( .A1(STATE_REG_SCAN_IN), .A2(n3359), .ZN(n4362) );
  NOR2_X1 U4148 ( .A1(n3360), .A2(n3581), .ZN(n3361) );
  AOI211_X1 U4149 ( .C1(n3579), .C2(n3776), .A(n4362), .B(n3361), .ZN(n3362)
         );
  OAI21_X1 U4150 ( .B1(n3583), .B2(n2150), .A(n3362), .ZN(n3363) );
  AOI21_X1 U4151 ( .B1(n3364), .B2(n3603), .A(n3363), .ZN(n3365) );
  OAI21_X1 U4152 ( .B1(n3366), .B2(n3599), .A(n3365), .ZN(U3228) );
  XOR2_X1 U4153 ( .A(n3368), .B(n3367), .Z(n3369) );
  XNOR2_X1 U4154 ( .A(n3370), .B(n3369), .ZN(n3376) );
  NOR2_X1 U4155 ( .A1(STATE_REG_SCAN_IN), .A2(n3371), .ZN(n4372) );
  NOR2_X1 U4156 ( .A1(n4185), .A2(n3593), .ZN(n3372) );
  AOI211_X1 U4157 ( .C1(n3589), .C2(n3776), .A(n4372), .B(n3372), .ZN(n3373)
         );
  OAI21_X1 U4158 ( .B1(n3583), .B2(n3429), .A(n3373), .ZN(n3374) );
  AOI21_X1 U4159 ( .B1(n3431), .B2(n3603), .A(n3374), .ZN(n3375) );
  OAI21_X1 U4160 ( .B1(n3376), .B2(n3599), .A(n3375), .ZN(U3233) );
  XOR2_X1 U4161 ( .A(n3377), .B(n3750), .Z(n3380) );
  OAI22_X1 U4162 ( .A1(n3402), .A2(n4155), .B1(n4154), .B2(n3382), .ZN(n3378)
         );
  AOI21_X1 U4163 ( .B1(n4159), .B2(n3777), .A(n3378), .ZN(n3379) );
  OAI21_X1 U4164 ( .B1(n3380), .B2(n4161), .A(n3379), .ZN(n3436) );
  INV_X1 U4165 ( .A(n3436), .ZN(n3389) );
  XOR2_X1 U4166 ( .A(n3381), .B(n3750), .Z(n3437) );
  NOR2_X1 U4167 ( .A1(n3383), .A2(n3382), .ZN(n3384) );
  AOI22_X1 U4168 ( .A1(n2017), .A2(REG2_REG_10__SCAN_IN), .B1(n3385), .B2(
        n4459), .ZN(n3386) );
  OAI21_X1 U4169 ( .B1(n3443), .B2(n4169), .A(n3386), .ZN(n3387) );
  AOI21_X1 U4170 ( .B1(n3437), .B2(n3920), .A(n3387), .ZN(n3388) );
  OAI21_X1 U4171 ( .B1(n3389), .B2(n2017), .A(n3388), .ZN(U3280) );
  NOR2_X1 U4172 ( .A1(n2127), .A2(n3392), .ZN(n3393) );
  XNOR2_X1 U4173 ( .A(n3390), .B(n3393), .ZN(n3398) );
  NOR2_X1 U4174 ( .A1(n3461), .A2(n3593), .ZN(n3395) );
  NAND2_X1 U4175 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4383) );
  OAI21_X1 U4176 ( .B1(n3402), .B2(n3581), .A(n4383), .ZN(n3394) );
  AOI211_X1 U4177 ( .C1(n3407), .C2(n3590), .A(n3395), .B(n3394), .ZN(n3397)
         );
  NAND2_X1 U4178 ( .A1(n3603), .A2(n3409), .ZN(n3396) );
  OAI211_X1 U4179 ( .C1(n3398), .C2(n3599), .A(n3397), .B(n3396), .ZN(U3221)
         );
  INV_X1 U4180 ( .A(n3399), .ZN(n3400) );
  AOI21_X1 U4181 ( .B1(n3417), .B2(n3401), .A(n3400), .ZN(n4178) );
  NAND2_X1 U4182 ( .A1(n4177), .A2(n4175), .ZN(n3719) );
  XNOR2_X1 U4183 ( .A(n4178), .B(n3719), .ZN(n3406) );
  OR2_X1 U4184 ( .A1(n3402), .A2(n4184), .ZN(n3404) );
  NAND2_X1 U4185 ( .A1(n3407), .A2(n4450), .ZN(n3403) );
  OAI211_X1 U4186 ( .C1(n3461), .C2(n4155), .A(n3404), .B(n3403), .ZN(n3405)
         );
  AOI21_X1 U4187 ( .B1(n3406), .B2(n4281), .A(n3405), .ZN(n4274) );
  NAND2_X1 U4188 ( .A1(n3428), .A2(n3407), .ZN(n3408) );
  NAND2_X1 U4189 ( .A1(n4189), .A2(n3408), .ZN(n4336) );
  INV_X1 U4190 ( .A(n4336), .ZN(n3413) );
  INV_X1 U4191 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3411) );
  INV_X1 U4192 ( .A(n3409), .ZN(n3410) );
  OAI22_X1 U4193 ( .A1(n4195), .A2(n3411), .B1(n3410), .B2(n4193), .ZN(n3412)
         );
  AOI21_X1 U4194 ( .B1(n3413), .B2(n4444), .A(n3412), .ZN(n3416) );
  XNOR2_X1 U4195 ( .A(n3414), .B(n3719), .ZN(n4273) );
  NAND2_X1 U4196 ( .A1(n4273), .A2(n3920), .ZN(n3415) );
  OAI211_X1 U4197 ( .C1(n4274), .C2(n2017), .A(n3416), .B(n3415), .ZN(U3278)
         );
  XOR2_X1 U4198 ( .A(n3710), .B(n3417), .Z(n3427) );
  NAND2_X1 U4199 ( .A1(n3419), .A2(n3710), .ZN(n3420) );
  NAND2_X1 U4200 ( .A1(n3418), .A2(n3420), .ZN(n4519) );
  AOI22_X1 U4201 ( .A1(n3775), .A2(n4280), .B1(n3421), .B2(n4450), .ZN(n3422)
         );
  OAI21_X1 U4202 ( .B1(n3423), .B2(n4184), .A(n3422), .ZN(n3424) );
  AOI21_X1 U4203 ( .B1(n4519), .B2(n3425), .A(n3424), .ZN(n3426) );
  OAI21_X1 U4204 ( .B1(n4161), .B2(n3427), .A(n3426), .ZN(n4517) );
  INV_X1 U4205 ( .A(n4517), .ZN(n3435) );
  OAI21_X1 U4206 ( .B1(n3430), .B2(n3429), .A(n3428), .ZN(n4516) );
  AOI22_X1 U4207 ( .A1(n2017), .A2(REG2_REG_11__SCAN_IN), .B1(n3431), .B2(
        n4459), .ZN(n3432) );
  OAI21_X1 U4208 ( .B1(n4516), .B2(n4169), .A(n3432), .ZN(n3433) );
  AOI21_X1 U4209 ( .B1(n4519), .B2(n4460), .A(n3433), .ZN(n3434) );
  OAI21_X1 U4210 ( .B1(n3435), .B2(n2017), .A(n3434), .ZN(U3279) );
  INV_X1 U4211 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3438) );
  AOI21_X1 U4212 ( .B1(n4513), .B2(n3437), .A(n3436), .ZN(n3440) );
  MUX2_X1 U4213 ( .A(n3438), .B(n3440), .S(n4692), .Z(n3439) );
  OAI21_X1 U4214 ( .B1(n3443), .B2(n4335), .A(n3439), .ZN(U3487) );
  MUX2_X1 U4215 ( .A(n3441), .B(n3440), .S(n4533), .Z(n3442) );
  OAI21_X1 U4216 ( .B1(n3443), .B2(n4278), .A(n3442), .ZN(U3528) );
  INV_X1 U4217 ( .A(n3444), .ZN(n3446) );
  INV_X1 U4218 ( .A(IR_REG_30__SCAN_IN), .ZN(n4663) );
  NAND3_X1 U4219 ( .A1(IR_REG_31__SCAN_IN), .A2(STATE_REG_SCAN_IN), .A3(n4663), 
        .ZN(n3445) );
  INV_X1 U4220 ( .A(DATAI_31_), .ZN(n4680) );
  OAI22_X1 U4221 ( .A1(n3446), .A2(n3445), .B1(STATE_REG_SCAN_IN), .B2(n4680), 
        .ZN(U3321) );
  INV_X1 U4222 ( .A(n3447), .ZN(n3453) );
  INV_X1 U4223 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3448) );
  OAI22_X1 U4224 ( .A1(n3449), .A2(n4193), .B1(n3448), .B2(n4195), .ZN(n3452)
         );
  NOR2_X1 U4225 ( .A1(n3450), .A2(n2017), .ZN(n3451) );
  AOI211_X1 U4226 ( .C1(n4444), .C2(n3453), .A(n3452), .B(n3451), .ZN(n3454)
         );
  OAI21_X1 U4227 ( .B1(n3455), .B2(n4172), .A(n3454), .ZN(U3262) );
  INV_X1 U4228 ( .A(n3457), .ZN(n3459) );
  NOR2_X1 U4229 ( .A1(n3459), .A2(n3458), .ZN(n3460) );
  XNOR2_X1 U4230 ( .A(n3456), .B(n3460), .ZN(n3466) );
  NAND2_X1 U4231 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4413) );
  OAI21_X1 U4232 ( .B1(n3461), .B2(n3581), .A(n4413), .ZN(n3462) );
  AOI21_X1 U4233 ( .B1(n3579), .B2(n3774), .A(n3462), .ZN(n3463) );
  OAI21_X1 U4234 ( .B1(n3583), .B2(n4165), .A(n3463), .ZN(n3464) );
  AOI21_X1 U4235 ( .B1(n4167), .B2(n3603), .A(n3464), .ZN(n3465) );
  OAI21_X1 U4236 ( .B1(n3466), .B2(n3599), .A(n3465), .ZN(U3212) );
  AND2_X1 U4237 ( .A1(n3566), .A2(n3467), .ZN(n3470) );
  OAI211_X1 U4238 ( .C1(n3470), .C2(n3469), .A(n3563), .B(n3468), .ZN(n3475)
         );
  AOI22_X1 U4239 ( .A1(n3579), .A2(n3957), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3471) );
  OAI21_X1 U4240 ( .B1(n4029), .B2(n3581), .A(n3471), .ZN(n3472) );
  AOI21_X1 U4241 ( .B1(n3473), .B2(n3590), .A(n3472), .ZN(n3474) );
  OAI211_X1 U4242 ( .C1(n3557), .C2(n4001), .A(n3475), .B(n3474), .ZN(U3213)
         );
  INV_X1 U4243 ( .A(n3476), .ZN(n3480) );
  AOI21_X1 U4244 ( .B1(n3476), .B2(n3478), .A(n3477), .ZN(n3479) );
  AOI21_X1 U4245 ( .B1(n3480), .B2(n3576), .A(n3479), .ZN(n3484) );
  NAND2_X1 U4246 ( .A1(n3482), .A2(n3481), .ZN(n3483) );
  XNOR2_X1 U4247 ( .A(n3484), .B(n3483), .ZN(n3489) );
  NAND2_X1 U4248 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3886) );
  OAI21_X1 U4249 ( .B1(n4071), .B2(n3593), .A(n3886), .ZN(n3485) );
  AOI21_X1 U4250 ( .B1(n3589), .B2(n4073), .A(n3485), .ZN(n3486) );
  OAI21_X1 U4251 ( .B1(n3583), .B2(n4076), .A(n3486), .ZN(n3487) );
  AOI21_X1 U4252 ( .B1(n4080), .B2(n3603), .A(n3487), .ZN(n3488) );
  OAI21_X1 U4253 ( .B1(n3489), .B2(n3599), .A(n3488), .ZN(U3216) );
  INV_X1 U4254 ( .A(n4037), .ZN(n3499) );
  NAND2_X1 U4255 ( .A1(n2256), .A2(n3490), .ZN(n3493) );
  INV_X1 U4256 ( .A(n3544), .ZN(n3542) );
  OAI211_X1 U4257 ( .C1(n3491), .C2(n3542), .A(n3545), .B(n3493), .ZN(n3492)
         );
  OAI211_X1 U4258 ( .C1(n3494), .C2(n3493), .A(n3563), .B(n3492), .ZN(n3498)
         );
  AOI22_X1 U4259 ( .A1(n3579), .A2(n3996), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3495) );
  OAI21_X1 U4260 ( .B1(n4071), .B2(n3581), .A(n3495), .ZN(n3496) );
  AOI21_X1 U4261 ( .B1(n4034), .B2(n3590), .A(n3496), .ZN(n3497) );
  OAI211_X1 U4262 ( .C1(n3557), .C2(n3499), .A(n3498), .B(n3497), .ZN(U3220)
         );
  INV_X1 U4263 ( .A(n3500), .ZN(n3502) );
  NOR2_X1 U4264 ( .A1(n3502), .A2(n3501), .ZN(n3503) );
  XNOR2_X1 U4265 ( .A(n3504), .B(n3503), .ZN(n3510) );
  AOI22_X1 U4266 ( .A1(n3579), .A2(n3772), .B1(REG3_REG_25__SCAN_IN), .B2(
        U3149), .ZN(n3505) );
  OAI21_X1 U4267 ( .B1(n3994), .B2(n3581), .A(n3505), .ZN(n3507) );
  NOR2_X1 U4268 ( .A1(n3557), .A2(n3962), .ZN(n3506) );
  AOI211_X1 U4269 ( .C1(n3508), .C2(n3590), .A(n3507), .B(n3506), .ZN(n3509)
         );
  OAI21_X1 U4270 ( .B1(n3510), .B2(n3599), .A(n3509), .ZN(U3222) );
  INV_X1 U4271 ( .A(n3596), .ZN(n3511) );
  OAI21_X1 U4272 ( .B1(n3511), .B2(n3598), .A(n3595), .ZN(n3512) );
  XOR2_X1 U4273 ( .A(n3513), .B(n3512), .Z(n3518) );
  NAND2_X1 U4274 ( .A1(REG3_REG_16__SCAN_IN), .A2(U3149), .ZN(n4416) );
  OAI21_X1 U4275 ( .B1(n4156), .B2(n3581), .A(n4416), .ZN(n3514) );
  AOI21_X1 U4276 ( .B1(n3579), .B2(n3773), .A(n3514), .ZN(n3515) );
  OAI21_X1 U4277 ( .B1(n3583), .B2(n4128), .A(n3515), .ZN(n3516) );
  AOI21_X1 U4278 ( .B1(n4123), .B2(n3603), .A(n3516), .ZN(n3517) );
  OAI21_X1 U4279 ( .B1(n3518), .B2(n3599), .A(n3517), .ZN(U3223) );
  NAND2_X1 U4280 ( .A1(n3520), .A2(n3519), .ZN(n3522) );
  XOR2_X1 U4281 ( .A(n3522), .B(n3521), .Z(n3529) );
  NOR2_X1 U4282 ( .A1(n3557), .A2(n3523), .ZN(n3528) );
  AND2_X1 U4283 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4428) );
  AOI21_X1 U4284 ( .B1(n4073), .B2(n3579), .A(n4428), .ZN(n3526) );
  NAND2_X1 U4285 ( .A1(n3590), .A2(n3524), .ZN(n3525) );
  OAI211_X1 U4286 ( .C1(n3594), .C2(n3581), .A(n3526), .B(n3525), .ZN(n3527)
         );
  AOI211_X1 U4287 ( .C1(n3529), .C2(n3563), .A(n3528), .B(n3527), .ZN(n3530)
         );
  INV_X1 U4288 ( .A(n3530), .ZN(U3225) );
  NAND2_X1 U4289 ( .A1(n3531), .A2(n3532), .ZN(n3533) );
  XOR2_X1 U4290 ( .A(n3534), .B(n3533), .Z(n3541) );
  NOR2_X1 U4291 ( .A1(n3557), .A2(n3981), .ZN(n3538) );
  AOI22_X1 U4292 ( .A1(n3535), .A2(n3579), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3536) );
  OAI21_X1 U4293 ( .B1(n4016), .B2(n3581), .A(n3536), .ZN(n3537) );
  AOI211_X1 U4294 ( .C1(n3539), .C2(n3590), .A(n3538), .B(n3537), .ZN(n3540)
         );
  OAI21_X1 U4295 ( .B1(n3541), .B2(n3599), .A(n3540), .ZN(U3226) );
  NOR2_X1 U4296 ( .A1(n3543), .A2(n3542), .ZN(n3547) );
  AOI21_X1 U4297 ( .B1(n3545), .B2(n3544), .A(n3491), .ZN(n3546) );
  OAI21_X1 U4298 ( .B1(n3547), .B2(n3546), .A(n3563), .ZN(n3551) );
  OAI22_X1 U4299 ( .A1(n4044), .A2(n3593), .B1(STATE_REG_SCAN_IN), .B2(n4583), 
        .ZN(n3549) );
  NOR2_X1 U4300 ( .A1(n3583), .A2(n4043), .ZN(n3548) );
  AOI211_X1 U4301 ( .C1(n3589), .C2(n4090), .A(n3549), .B(n3548), .ZN(n3550)
         );
  OAI211_X1 U4302 ( .C1(n3557), .C2(n3552), .A(n3551), .B(n3550), .ZN(U3230)
         );
  XNOR2_X1 U4303 ( .A(n3555), .B(n3554), .ZN(n3556) );
  XNOR2_X1 U4304 ( .A(n3553), .B(n3556), .ZN(n3564) );
  NOR2_X1 U4305 ( .A1(n3557), .A2(n4194), .ZN(n3562) );
  INV_X1 U4306 ( .A(REG3_REG_13__SCAN_IN), .ZN(n3558) );
  NOR2_X1 U4307 ( .A1(STATE_REG_SCAN_IN), .A2(n3558), .ZN(n4393) );
  AOI21_X1 U4308 ( .B1(n4182), .B2(n3579), .A(n4393), .ZN(n3560) );
  NAND2_X1 U4309 ( .A1(n3590), .A2(n4181), .ZN(n3559) );
  OAI211_X1 U4310 ( .C1(n4185), .C2(n3581), .A(n3560), .B(n3559), .ZN(n3561)
         );
  AOI211_X1 U4311 ( .C1(n3564), .C2(n3563), .A(n3562), .B(n3561), .ZN(n3565)
         );
  INV_X1 U4312 ( .A(n3565), .ZN(U3231) );
  INV_X1 U4313 ( .A(n3566), .ZN(n3567) );
  AOI21_X1 U4314 ( .B1(n3569), .B2(n3568), .A(n3567), .ZN(n3575) );
  INV_X1 U4315 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3570) );
  OAI22_X1 U4316 ( .A1(n4016), .A2(n3593), .B1(STATE_REG_SCAN_IN), .B2(n3570), 
        .ZN(n3572) );
  NOR2_X1 U4317 ( .A1(n3583), .A2(n4020), .ZN(n3571) );
  AOI211_X1 U4318 ( .C1(n3589), .C2(n4013), .A(n3572), .B(n3571), .ZN(n3574)
         );
  NAND2_X1 U4319 ( .A1(n3603), .A2(n4019), .ZN(n3573) );
  OAI211_X1 U4320 ( .C1(n3575), .C2(n3599), .A(n3574), .B(n3573), .ZN(U3232)
         );
  XNOR2_X1 U4321 ( .A(n3577), .B(n3576), .ZN(n3578) );
  XNOR2_X1 U4322 ( .A(n3476), .B(n3578), .ZN(n3587) );
  NAND2_X1 U4323 ( .A1(n3579), .A2(n4090), .ZN(n3580) );
  NAND2_X1 U4324 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n3867) );
  OAI211_X1 U4325 ( .C1(n4129), .C2(n3581), .A(n3580), .B(n3867), .ZN(n3585)
         );
  NOR2_X1 U4326 ( .A1(n3583), .A2(n3582), .ZN(n3584) );
  AOI211_X1 U4327 ( .C1(n4097), .C2(n3603), .A(n3585), .B(n3584), .ZN(n3586)
         );
  OAI21_X1 U4328 ( .B1(n3587), .B2(n3599), .A(n3586), .ZN(U3235) );
  NOR2_X1 U4329 ( .A1(STATE_REG_SCAN_IN), .A2(n3588), .ZN(n3855) );
  AOI21_X1 U4330 ( .B1(n4182), .B2(n3589), .A(n3855), .ZN(n3592) );
  NAND2_X1 U4331 ( .A1(n3590), .A2(n4144), .ZN(n3591) );
  OAI211_X1 U4332 ( .C1(n3594), .C2(n3593), .A(n3592), .B(n3591), .ZN(n3602)
         );
  NAND2_X1 U4333 ( .A1(n3596), .A2(n3595), .ZN(n3597) );
  XOR2_X1 U4334 ( .A(n3598), .B(n3597), .Z(n3600) );
  NOR2_X1 U4335 ( .A1(n3600), .A2(n3599), .ZN(n3601) );
  AOI211_X1 U4336 ( .C1(n4145), .C2(n3603), .A(n3602), .B(n3601), .ZN(n3604)
         );
  INV_X1 U4337 ( .A(n3604), .ZN(U3238) );
  NAND2_X1 U4338 ( .A1(n3622), .A2(DATAI_30_), .ZN(n4209) );
  NAND2_X1 U4339 ( .A1(n3605), .A2(REG1_REG_31__SCAN_IN), .ZN(n3609) );
  NAND2_X1 U4340 ( .A1(n3606), .A2(REG2_REG_31__SCAN_IN), .ZN(n3608) );
  NAND2_X1 U4341 ( .A1(n2973), .A2(REG0_REG_31__SCAN_IN), .ZN(n3607) );
  NAND3_X1 U4342 ( .A1(n3609), .A2(n3608), .A3(n3607), .ZN(n4203) );
  NAND2_X1 U4343 ( .A1(n3610), .A2(n3613), .ZN(n3678) );
  NAND2_X1 U4344 ( .A1(n3612), .A2(n3611), .ZN(n3662) );
  NAND2_X1 U4345 ( .A1(n3662), .A2(n3613), .ZN(n3677) );
  OAI21_X1 U4346 ( .B1(n4153), .B2(n3678), .A(n3677), .ZN(n3614) );
  AOI211_X1 U4347 ( .C1(n3614), .C2(n3686), .A(n2066), .B(n3685), .ZN(n3616)
         );
  INV_X1 U4348 ( .A(n3615), .ZN(n3689) );
  OAI21_X1 U4349 ( .B1(n3616), .B2(n3689), .A(n3688), .ZN(n3618) );
  AOI21_X1 U4350 ( .B1(n3692), .B2(n3618), .A(n3617), .ZN(n3619) );
  OAI21_X1 U4351 ( .B1(n3619), .B2(n3694), .A(n3932), .ZN(n3620) );
  NAND4_X1 U4352 ( .A1(n3621), .A2(n3623), .A3(n3624), .A4(n3620), .ZN(n3632)
         );
  INV_X1 U4353 ( .A(n3771), .ZN(n3626) );
  NAND2_X1 U4354 ( .A1(n3622), .A2(DATAI_29_), .ZN(n3714) );
  NAND2_X1 U4355 ( .A1(n3622), .A2(DATAI_31_), .ZN(n4201) );
  NAND2_X1 U4356 ( .A1(n4203), .A2(n4201), .ZN(n3705) );
  OAI21_X1 U4357 ( .B1(n3896), .B2(n4209), .A(n3705), .ZN(n3738) );
  AOI21_X1 U4358 ( .B1(n3626), .B2(n3908), .A(n3738), .ZN(n3627) );
  INV_X1 U4359 ( .A(n3627), .ZN(n3631) );
  INV_X1 U4360 ( .A(n3623), .ZN(n3891) );
  INV_X1 U4361 ( .A(n3624), .ZN(n3625) );
  NOR2_X1 U4362 ( .A1(n3891), .A2(n3625), .ZN(n3628) );
  OAI21_X1 U4363 ( .B1(n3626), .B2(n3908), .A(n3892), .ZN(n3697) );
  OAI21_X1 U4364 ( .B1(n3628), .B2(n3697), .A(n3627), .ZN(n3701) );
  NOR3_X1 U4365 ( .A1(n3629), .A2(n3919), .A3(n3697), .ZN(n3630) );
  OAI22_X1 U4366 ( .A1(n3632), .A2(n3631), .B1(n3701), .B2(n3630), .ZN(n3633)
         );
  OAI21_X1 U4367 ( .B1(n4209), .B2(n4203), .A(n3633), .ZN(n3637) );
  AND2_X1 U4368 ( .A1(n3896), .A2(n4209), .ZN(n3703) );
  INV_X1 U4369 ( .A(n4203), .ZN(n3634) );
  INV_X1 U4370 ( .A(n4201), .ZN(n4204) );
  OAI21_X1 U4371 ( .B1(n3703), .B2(n3634), .A(n4204), .ZN(n3636) );
  AOI21_X1 U4372 ( .B1(n3637), .B2(n3636), .A(n3635), .ZN(n3763) );
  NOR2_X1 U4373 ( .A1(n3639), .A2(n3638), .ZN(n3700) );
  INV_X1 U4374 ( .A(n3730), .ZN(n3642) );
  NAND2_X1 U4375 ( .A1(n3784), .A2(n4453), .ZN(n3729) );
  OAI211_X1 U4376 ( .C1(n3642), .C2(n3641), .A(n3729), .B(n3640), .ZN(n3645)
         );
  NAND3_X1 U4377 ( .A1(n3645), .A2(n3644), .A3(n3643), .ZN(n3648) );
  NAND3_X1 U4378 ( .A1(n3648), .A2(n3647), .A3(n3646), .ZN(n3651) );
  NAND3_X1 U4379 ( .A1(n3651), .A2(n3650), .A3(n3649), .ZN(n3654) );
  NAND4_X1 U4380 ( .A1(n3654), .A2(n3653), .A3(n3652), .A4(n3664), .ZN(n3656)
         );
  AND3_X1 U4381 ( .A1(n3656), .A2(n3711), .A3(n3655), .ZN(n3661) );
  NAND2_X1 U4382 ( .A1(n3658), .A2(n3657), .ZN(n3666) );
  OAI211_X1 U4383 ( .C1(n3661), .C2(n3666), .A(n3660), .B(n3659), .ZN(n3670)
         );
  INV_X1 U4384 ( .A(n3662), .ZN(n3669) );
  INV_X1 U4385 ( .A(n3663), .ZN(n3665) );
  NAND2_X1 U4386 ( .A1(n3665), .A2(n3664), .ZN(n3667) );
  OAI21_X1 U4387 ( .B1(n3667), .B2(n3666), .A(n3671), .ZN(n3668) );
  AOI22_X1 U4388 ( .A1(n3670), .A2(n3669), .B1(n3677), .B2(n3668), .ZN(n3682)
         );
  INV_X1 U4389 ( .A(n3671), .ZN(n3675) );
  OAI211_X1 U4390 ( .C1(n3675), .C2(n3674), .A(n3673), .B(n3672), .ZN(n3681)
         );
  INV_X1 U4391 ( .A(n3676), .ZN(n3679) );
  OAI21_X1 U4392 ( .B1(n3679), .B2(n3678), .A(n3677), .ZN(n3680) );
  OAI21_X1 U4393 ( .B1(n3682), .B2(n3681), .A(n3680), .ZN(n3684) );
  NAND2_X1 U4394 ( .A1(n3684), .A2(n3683), .ZN(n3687) );
  AOI21_X1 U4395 ( .B1(n3687), .B2(n3686), .A(n3685), .ZN(n3690) );
  INV_X1 U4396 ( .A(n3988), .ZN(n3744) );
  OAI211_X1 U4397 ( .C1(n3690), .C2(n3689), .A(n3744), .B(n3688), .ZN(n3691)
         );
  NAND2_X1 U4398 ( .A1(n3692), .A2(n3691), .ZN(n3695) );
  AOI211_X1 U4399 ( .C1(n3696), .C2(n3695), .A(n3694), .B(n3693), .ZN(n3699)
         );
  NOR4_X1 U4400 ( .A1(n3700), .A2(n3699), .A3(n3698), .A4(n3697), .ZN(n3702)
         );
  OR2_X1 U4401 ( .A1(n3702), .A2(n3701), .ZN(n3707) );
  INV_X1 U4402 ( .A(n3703), .ZN(n3704) );
  OAI21_X1 U4403 ( .B1(n4203), .B2(n4201), .A(n3704), .ZN(n3737) );
  NAND2_X1 U4404 ( .A1(n3737), .A2(n3705), .ZN(n3706) );
  NAND2_X1 U4405 ( .A1(n3707), .A2(n3706), .ZN(n3761) );
  OR2_X1 U4406 ( .A1(n4089), .A2(n4152), .ZN(n3713) );
  NAND4_X1 U4407 ( .A1(n3711), .A2(n3710), .A3(n3709), .A4(n3708), .ZN(n3712)
         );
  NOR3_X1 U4408 ( .A1(n3904), .A2(n3713), .A3(n3712), .ZN(n3756) );
  XNOR2_X1 U4409 ( .A(n3771), .B(n3714), .ZN(n3906) );
  XNOR2_X1 U4410 ( .A(n4031), .B(n4043), .ZN(n4047) );
  OR2_X1 U4411 ( .A1(n3906), .A2(n4047), .ZN(n3715) );
  NOR2_X1 U4412 ( .A1(n3919), .A2(n3715), .ZN(n3755) );
  NAND2_X1 U4413 ( .A1(n3716), .A2(n3930), .ZN(n3954) );
  NAND2_X1 U4414 ( .A1(n3717), .A2(n3951), .ZN(n3971) );
  NOR2_X1 U4415 ( .A1(n3954), .A2(n3971), .ZN(n3726) );
  NAND2_X1 U4416 ( .A1(n3718), .A2(n3969), .ZN(n3992) );
  NAND2_X1 U4417 ( .A1(n4064), .A2(n4063), .ZN(n4105) );
  NOR2_X1 U4418 ( .A1(n3992), .A2(n4105), .ZN(n3725) );
  NOR2_X1 U4419 ( .A1(n3720), .A2(n3719), .ZN(n3724) );
  NOR2_X1 U4420 ( .A1(n3722), .A2(n3721), .ZN(n3723) );
  NAND4_X1 U4421 ( .A1(n3726), .A2(n3725), .A3(n3724), .A4(n3723), .ZN(n3743)
         );
  NAND2_X1 U4422 ( .A1(n3728), .A2(n3727), .ZN(n3933) );
  INV_X1 U4423 ( .A(n3933), .ZN(n3741) );
  INV_X1 U4424 ( .A(n3731), .ZN(n3733) );
  INV_X1 U4425 ( .A(n3734), .ZN(n3736) );
  NOR2_X1 U4426 ( .A1(n4070), .A2(n4180), .ZN(n3740) );
  NOR2_X1 U4427 ( .A1(n3738), .A2(n3737), .ZN(n3739) );
  NAND4_X1 U4428 ( .A1(n3741), .A2(n4456), .A3(n3740), .A4(n3739), .ZN(n3742)
         );
  NOR2_X1 U4429 ( .A1(n3743), .A2(n3742), .ZN(n3754) );
  NAND2_X1 U4430 ( .A1(n3744), .A2(n3989), .ZN(n4027) );
  INV_X1 U4431 ( .A(n4027), .ZN(n3748) );
  INV_X1 U4432 ( .A(n3113), .ZN(n3747) );
  INV_X1 U4433 ( .A(n3745), .ZN(n4138) );
  NAND4_X1 U4434 ( .A1(n3748), .A2(n3747), .A3(n3746), .A4(n4138), .ZN(n3752)
         );
  NAND4_X1 U4435 ( .A1(n2189), .A2(n4011), .A3(n3750), .A4(n3749), .ZN(n3751)
         );
  NOR2_X1 U4436 ( .A1(n3752), .A2(n3751), .ZN(n3753) );
  NAND4_X1 U4437 ( .A1(n3756), .A2(n3755), .A3(n3754), .A4(n3753), .ZN(n3758)
         );
  AND2_X1 U4438 ( .A1(n3758), .A2(n3757), .ZN(n3760) );
  MUX2_X1 U4439 ( .A(n3761), .B(n3760), .S(n3759), .Z(n3762) );
  NOR2_X1 U4440 ( .A1(n3763), .A2(n3762), .ZN(n3764) );
  XNOR2_X1 U4441 ( .A(n3764), .B(n4342), .ZN(n3770) );
  NAND2_X1 U4442 ( .A1(n3766), .A2(n3765), .ZN(n3767) );
  OAI211_X1 U4443 ( .C1(n4341), .C2(n3769), .A(n3767), .B(B_REG_SCAN_IN), .ZN(
        n3768) );
  OAI21_X1 U4444 ( .B1(n3770), .B2(n3769), .A(n3768), .ZN(U3239) );
  MUX2_X1 U4445 ( .A(n4203), .B(DATAO_REG_31__SCAN_IN), .S(n3783), .Z(U3581)
         );
  MUX2_X1 U4446 ( .A(n3771), .B(DATAO_REG_29__SCAN_IN), .S(n3783), .Z(U3579)
         );
  INV_X1 U4447 ( .A(n3898), .ZN(n3917) );
  MUX2_X1 U4448 ( .A(DATAO_REG_28__SCAN_IN), .B(n3917), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4449 ( .A(n3772), .B(DATAO_REG_26__SCAN_IN), .S(n3783), .Z(U3576)
         );
  MUX2_X1 U4450 ( .A(n3957), .B(DATAO_REG_24__SCAN_IN), .S(n3783), .Z(U3574)
         );
  MUX2_X1 U4451 ( .A(DATAO_REG_23__SCAN_IN), .B(n3975), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4452 ( .A(n3996), .B(DATAO_REG_22__SCAN_IN), .S(n3783), .Z(U3572)
         );
  MUX2_X1 U4453 ( .A(n4013), .B(DATAO_REG_21__SCAN_IN), .S(n3783), .Z(U3571)
         );
  MUX2_X1 U4454 ( .A(n4090), .B(DATAO_REG_19__SCAN_IN), .S(n3783), .Z(U3569)
         );
  MUX2_X1 U4455 ( .A(DATAO_REG_18__SCAN_IN), .B(n4073), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4456 ( .A(DATAO_REG_17__SCAN_IN), .B(n3773), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4457 ( .A(DATAO_REG_16__SCAN_IN), .B(n4140), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4458 ( .A(DATAO_REG_15__SCAN_IN), .B(n3774), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4459 ( .A(DATAO_REG_14__SCAN_IN), .B(n4182), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4460 ( .A(DATAO_REG_13__SCAN_IN), .B(n4158), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4461 ( .A(DATAO_REG_12__SCAN_IN), .B(n3775), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4462 ( .A(n3776), .B(DATAO_REG_10__SCAN_IN), .S(n3783), .Z(U3560)
         );
  MUX2_X1 U4463 ( .A(n3777), .B(DATAO_REG_9__SCAN_IN), .S(n3783), .Z(U3559) );
  MUX2_X1 U4464 ( .A(DATAO_REG_8__SCAN_IN), .B(n3778), .S(U4043), .Z(U3558) );
  MUX2_X1 U4465 ( .A(DATAO_REG_7__SCAN_IN), .B(n3779), .S(U4043), .Z(U3557) );
  MUX2_X1 U4466 ( .A(DATAO_REG_5__SCAN_IN), .B(n3780), .S(U4043), .Z(U3555) );
  MUX2_X1 U4467 ( .A(DATAO_REG_4__SCAN_IN), .B(n3781), .S(U4043), .Z(U3554) );
  MUX2_X1 U4468 ( .A(DATAO_REG_2__SCAN_IN), .B(n3782), .S(U4043), .Z(U3552) );
  MUX2_X1 U4469 ( .A(DATAO_REG_1__SCAN_IN), .B(n4279), .S(U4043), .Z(U3551) );
  MUX2_X1 U4470 ( .A(n3784), .B(DATAO_REG_0__SCAN_IN), .S(n3783), .Z(U3550) );
  AOI22_X1 U4471 ( .A1(n4429), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3792) );
  NAND2_X1 U4472 ( .A1(n4412), .A2(n4349), .ZN(n3791) );
  OAI211_X1 U4473 ( .C1(n3793), .C2(n3785), .A(n4439), .B(n3808), .ZN(n3790)
         );
  MUX2_X1 U4474 ( .A(n2990), .B(REG1_REG_1__SCAN_IN), .S(n4349), .Z(n3786) );
  OAI21_X1 U4475 ( .B1(n2146), .B2(n3787), .A(n3786), .ZN(n3788) );
  NAND3_X1 U4476 ( .A1(n4437), .A2(n3800), .A3(n3788), .ZN(n3789) );
  NAND4_X1 U4477 ( .A1(n3792), .A2(n3791), .A3(n3790), .A4(n3789), .ZN(U3241)
         );
  OR2_X1 U4478 ( .A1(n3794), .A2(n3793), .ZN(n3795) );
  OAI211_X1 U4479 ( .C1(n3797), .C2(n4338), .A(n3796), .B(n3795), .ZN(n3798)
         );
  OAI211_X1 U4480 ( .C1(IR_REG_0__SCAN_IN), .C2(n3799), .A(n3798), .B(U4043), 
        .ZN(n3825) );
  AOI22_X1 U4481 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4429), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3815) );
  MUX2_X1 U4482 ( .A(n2994), .B(REG1_REG_2__SCAN_IN), .S(n3807), .Z(n3802) );
  NAND3_X1 U4483 ( .A1(n3802), .A2(n3801), .A3(n3800), .ZN(n3803) );
  NAND3_X1 U4484 ( .A1(n4437), .A2(n3804), .A3(n3803), .ZN(n3806) );
  NAND2_X1 U4485 ( .A1(n4412), .A2(n3807), .ZN(n3805) );
  AND2_X1 U4486 ( .A1(n3806), .A2(n3805), .ZN(n3814) );
  MUX2_X1 U4487 ( .A(n2999), .B(REG2_REG_2__SCAN_IN), .S(n3807), .Z(n3810) );
  NAND3_X1 U4488 ( .A1(n3810), .A2(n3809), .A3(n3808), .ZN(n3811) );
  NAND3_X1 U4489 ( .A1(n4439), .A2(n3812), .A3(n3811), .ZN(n3813) );
  NAND4_X1 U4490 ( .A1(n3825), .A2(n3815), .A3(n3814), .A4(n3813), .ZN(U3242)
         );
  NAND2_X1 U4491 ( .A1(n4429), .A2(ADDR_REG_4__SCAN_IN), .ZN(n3824) );
  INV_X1 U4492 ( .A(n3816), .ZN(n3822) );
  XNOR2_X1 U4493 ( .A(n3817), .B(REG1_REG_4__SCAN_IN), .ZN(n3820) );
  XNOR2_X1 U4494 ( .A(n3818), .B(REG2_REG_4__SCAN_IN), .ZN(n3819) );
  OAI22_X1 U4495 ( .A1(n3820), .A2(n4401), .B1(n4405), .B2(n3819), .ZN(n3821)
         );
  AOI211_X1 U4496 ( .C1(n4347), .C2(n4412), .A(n3822), .B(n3821), .ZN(n3823)
         );
  NAND3_X1 U4497 ( .A1(n3825), .A2(n3824), .A3(n3823), .ZN(U3244) );
  INV_X1 U4498 ( .A(n4343), .ZN(n3858) );
  NAND2_X1 U4499 ( .A1(n3858), .A2(REG2_REG_15__SCAN_IN), .ZN(n3828) );
  INV_X1 U4500 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3826) );
  NAND2_X1 U4501 ( .A1(n4343), .A2(n3826), .ZN(n3827) );
  AND2_X1 U4502 ( .A1(n3828), .A2(n3827), .ZN(n3841) );
  INV_X1 U4503 ( .A(n4411), .ZN(n4472) );
  INV_X1 U4504 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4395) );
  NOR2_X1 U4505 ( .A1(n4395), .A2(n4473), .ZN(n4394) );
  NAND2_X1 U4506 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4475), .ZN(n3834) );
  INV_X1 U4507 ( .A(n4475), .ZN(n4379) );
  INV_X1 U4508 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4509 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4475), .B1(n4379), .B2(
        n3829), .ZN(n4376) );
  NAND2_X1 U4510 ( .A1(n3831), .A2(n3830), .ZN(n3833) );
  NAND2_X1 U4511 ( .A1(n4376), .A2(n4375), .ZN(n4374) );
  NAND2_X1 U4512 ( .A1(n3846), .A2(n3835), .ZN(n3836) );
  OAI22_X1 U4513 ( .A1(n4394), .A2(n4397), .B1(REG2_REG_13__SCAN_IN), .B2(
        n3849), .ZN(n3837) );
  NOR2_X1 U4514 ( .A1(n4472), .A2(n3837), .ZN(n3838) );
  INV_X1 U4515 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4408) );
  XOR2_X1 U4516 ( .A(n4411), .B(n3837), .Z(n4407) );
  NOR2_X1 U4517 ( .A1(n4408), .A2(n4407), .ZN(n4406) );
  NOR2_X1 U4518 ( .A1(n3838), .A2(n4406), .ZN(n3840) );
  OR2_X1 U4519 ( .A1(n3840), .A2(n3841), .ZN(n3861) );
  INV_X1 U4520 ( .A(n3861), .ZN(n3839) );
  AOI21_X1 U4521 ( .B1(n3841), .B2(n3840), .A(n3839), .ZN(n3842) );
  NAND2_X1 U4522 ( .A1(n4439), .A2(n3842), .ZN(n3857) );
  INV_X1 U4523 ( .A(n3843), .ZN(n3845) );
  INV_X1 U4524 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4531) );
  AOI22_X1 U4525 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4379), .B1(n4475), .B2(
        n4531), .ZN(n4370) );
  NOR2_X1 U4526 ( .A1(n4371), .A2(n4370), .ZN(n4369) );
  NOR2_X1 U4527 ( .A1(n3847), .A2(n2167), .ZN(n3848) );
  INV_X1 U4528 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4382) );
  INV_X1 U4529 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4271) );
  AOI22_X1 U4530 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4473), .B1(n3849), .B2(
        n4271), .ZN(n4391) );
  INV_X1 U4531 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4404) );
  XOR2_X1 U4532 ( .A(n4411), .B(n3850), .Z(n4403) );
  NAND2_X1 U4533 ( .A1(n4343), .A2(REG1_REG_15__SCAN_IN), .ZN(n3868) );
  OAI21_X1 U4534 ( .B1(n4343), .B2(REG1_REG_15__SCAN_IN), .A(n3868), .ZN(n3852) );
  INV_X1 U4535 ( .A(n3869), .ZN(n3851) );
  AOI211_X1 U4536 ( .C1(n3853), .C2(n3852), .A(n3851), .B(n4401), .ZN(n3854)
         );
  AOI211_X1 U4537 ( .C1(n4429), .C2(ADDR_REG_15__SCAN_IN), .A(n3855), .B(n3854), .ZN(n3856) );
  OAI211_X1 U4538 ( .C1(n3858), .C2(n4442), .A(n3857), .B(n3856), .ZN(U3255)
         );
  INV_X1 U4539 ( .A(n3881), .ZN(n3877) );
  XNOR2_X1 U4540 ( .A(n3881), .B(REG2_REG_18__SCAN_IN), .ZN(n3865) );
  NOR2_X1 U4541 ( .A1(n3872), .A2(REG2_REG_17__SCAN_IN), .ZN(n3859) );
  AOI21_X1 U4542 ( .B1(REG2_REG_17__SCAN_IN), .B2(n3872), .A(n3859), .ZN(n4432) );
  NAND2_X1 U4543 ( .A1(n4343), .A2(REG2_REG_15__SCAN_IN), .ZN(n3860) );
  NAND2_X1 U4544 ( .A1(n3862), .A2(n4470), .ZN(n3863) );
  INV_X1 U4545 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4419) );
  NAND2_X1 U4546 ( .A1(n4432), .A2(n4431), .ZN(n4430) );
  OAI21_X1 U4547 ( .B1(n3872), .B2(REG2_REG_17__SCAN_IN), .A(n4430), .ZN(n3864) );
  NOR2_X1 U4548 ( .A1(n3864), .A2(n3865), .ZN(n3880) );
  AOI21_X1 U4549 ( .B1(n3865), .B2(n3864), .A(n3880), .ZN(n3866) );
  NAND2_X1 U4550 ( .A1(n4439), .A2(n3866), .ZN(n3876) );
  INV_X1 U4551 ( .A(n3867), .ZN(n3874) );
  XNOR2_X1 U4552 ( .A(n3881), .B(REG1_REG_18__SCAN_IN), .ZN(n3873) );
  INV_X1 U4553 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4596) );
  AOI22_X1 U4554 ( .A1(n3872), .A2(REG1_REG_17__SCAN_IN), .B1(n4596), .B2(
        n4468), .ZN(n4435) );
  NAND2_X1 U4555 ( .A1(n3870), .A2(n4470), .ZN(n3871) );
  INV_X1 U4556 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4422) );
  NAND2_X1 U4557 ( .A1(n4435), .A2(n4434), .ZN(n4433) );
  OAI211_X1 U4558 ( .C1(n3877), .C2(n4442), .A(n3876), .B(n3875), .ZN(U3258)
         );
  XNOR2_X1 U4559 ( .A(n4342), .B(REG1_REG_19__SCAN_IN), .ZN(n3879) );
  AOI21_X1 U4560 ( .B1(n3881), .B2(REG2_REG_18__SCAN_IN), .A(n3880), .ZN(n3884) );
  INV_X1 U4561 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3882) );
  MUX2_X1 U4562 ( .A(n3882), .B(REG2_REG_19__SCAN_IN), .S(n4451), .Z(n3883) );
  XNOR2_X1 U4563 ( .A(n3884), .B(n3883), .ZN(n3888) );
  NAND2_X1 U4564 ( .A1(n4429), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3885) );
  OAI211_X1 U4565 ( .C1(n4442), .C2(n4451), .A(n3886), .B(n3885), .ZN(n3887)
         );
  AOI21_X1 U4566 ( .B1(n3888), .B2(n4439), .A(n3887), .ZN(n3889) );
  INV_X1 U4567 ( .A(n3890), .ZN(n3902) );
  XNOR2_X1 U4568 ( .A(n3894), .B(n3906), .ZN(n3895) );
  AOI21_X1 U4569 ( .B1(n4338), .B2(B_REG_SCAN_IN), .A(n4155), .ZN(n4202) );
  AOI22_X1 U4570 ( .A1(n3896), .A2(n4202), .B1(n3908), .B2(n4450), .ZN(n3897)
         );
  AOI21_X1 U4571 ( .B1(n3902), .B2(n4459), .A(n4215), .ZN(n3911) );
  NAND2_X1 U4572 ( .A1(n4214), .A2(n3920), .ZN(n3910) );
  AOI22_X1 U4573 ( .A1(n4216), .A2(n4444), .B1(REG2_REG_29__SCAN_IN), .B2(
        n2017), .ZN(n3909) );
  OAI211_X1 U4574 ( .C1(n2017), .C2(n3911), .A(n3910), .B(n3909), .ZN(U3354)
         );
  OAI22_X1 U4575 ( .A1(n3955), .A2(n4184), .B1(n3922), .B2(n4154), .ZN(n3916)
         );
  NAND2_X1 U4576 ( .A1(n3912), .A2(n3919), .ZN(n3913) );
  AOI21_X1 U4577 ( .B1(n3914), .B2(n3913), .A(n4161), .ZN(n3915) );
  AOI211_X1 U4578 ( .C1(n4280), .C2(n3917), .A(n3916), .B(n3915), .ZN(n4218)
         );
  XNOR2_X1 U4579 ( .A(n3918), .B(n3919), .ZN(n4217) );
  NAND2_X1 U4580 ( .A1(n4217), .A2(n3920), .ZN(n3928) );
  OAI21_X1 U4581 ( .B1(n3942), .B2(n3922), .A(n3921), .ZN(n4220) );
  INV_X1 U4582 ( .A(n4220), .ZN(n3926) );
  INV_X1 U4583 ( .A(REG2_REG_27__SCAN_IN), .ZN(n3923) );
  OAI22_X1 U4584 ( .A1(n3924), .A2(n4193), .B1(n4195), .B2(n3923), .ZN(n3925)
         );
  AOI21_X1 U4585 ( .B1(n3926), .B2(n4444), .A(n3925), .ZN(n3927) );
  OAI211_X1 U4586 ( .C1(n4218), .C2(n2017), .A(n3928), .B(n3927), .ZN(U3263)
         );
  XNOR2_X1 U4587 ( .A(n3929), .B(n3933), .ZN(n4222) );
  INV_X1 U4588 ( .A(n4222), .ZN(n3949) );
  INV_X1 U4589 ( .A(n3930), .ZN(n3931) );
  AOI21_X1 U4590 ( .B1(n3952), .B2(n3932), .A(n3931), .ZN(n3934) );
  XNOR2_X1 U4591 ( .A(n3934), .B(n3933), .ZN(n3935) );
  NAND2_X1 U4592 ( .A1(n3935), .A2(n4281), .ZN(n3939) );
  AOI22_X1 U4593 ( .A1(n3937), .A2(n4280), .B1(n4450), .B2(n3936), .ZN(n3938)
         );
  OAI211_X1 U4594 ( .C1(n3973), .C2(n4184), .A(n3939), .B(n3938), .ZN(n4221)
         );
  INV_X1 U4595 ( .A(REG2_REG_26__SCAN_IN), .ZN(n3941) );
  OAI22_X1 U4596 ( .A1(n4195), .A2(n3941), .B1(n3940), .B2(n4193), .ZN(n3947)
         );
  INV_X1 U4597 ( .A(n3960), .ZN(n3945) );
  INV_X1 U4598 ( .A(n3942), .ZN(n3943) );
  OAI21_X1 U4599 ( .B1(n3945), .B2(n3944), .A(n3943), .ZN(n4293) );
  NOR2_X1 U4600 ( .A1(n4293), .A2(n4169), .ZN(n3946) );
  AOI211_X1 U4601 ( .C1(n4221), .C2(n4195), .A(n3947), .B(n3946), .ZN(n3948)
         );
  OAI21_X1 U4602 ( .B1(n3949), .B2(n4172), .A(n3948), .ZN(U3264) );
  XNOR2_X1 U4603 ( .A(n3950), .B(n3954), .ZN(n4226) );
  INV_X1 U4604 ( .A(n4226), .ZN(n3967) );
  NAND2_X1 U4605 ( .A1(n3952), .A2(n3951), .ZN(n3953) );
  XOR2_X1 U4606 ( .A(n3954), .B(n3953), .Z(n3959) );
  OAI22_X1 U4607 ( .A1(n3955), .A2(n4155), .B1(n4154), .B2(n3961), .ZN(n3956)
         );
  AOI21_X1 U4608 ( .B1(n4159), .B2(n3957), .A(n3956), .ZN(n3958) );
  OAI21_X1 U4609 ( .B1(n3959), .B2(n4161), .A(n3958), .ZN(n4225) );
  OAI21_X1 U4610 ( .B1(n2153), .B2(n3961), .A(n3960), .ZN(n4297) );
  NOR2_X1 U4611 ( .A1(n4297), .A2(n4169), .ZN(n3965) );
  INV_X1 U4612 ( .A(REG2_REG_25__SCAN_IN), .ZN(n3963) );
  OAI22_X1 U4613 ( .A1(n4195), .A2(n3963), .B1(n3962), .B2(n4193), .ZN(n3964)
         );
  AOI211_X1 U4614 ( .C1(n4225), .C2(n4195), .A(n3965), .B(n3964), .ZN(n3966)
         );
  OAI21_X1 U4615 ( .B1(n3967), .B2(n4172), .A(n3966), .ZN(U3265) );
  XOR2_X1 U4616 ( .A(n3971), .B(n3968), .Z(n4230) );
  INV_X1 U4617 ( .A(n4230), .ZN(n3986) );
  NAND2_X1 U4618 ( .A1(n3970), .A2(n3969), .ZN(n3972) );
  XNOR2_X1 U4619 ( .A(n3972), .B(n3971), .ZN(n3977) );
  OAI22_X1 U4620 ( .A1(n3973), .A2(n4155), .B1(n4154), .B2(n3979), .ZN(n3974)
         );
  AOI21_X1 U4621 ( .B1(n4159), .B2(n3975), .A(n3974), .ZN(n3976) );
  OAI21_X1 U4622 ( .B1(n3977), .B2(n4161), .A(n3976), .ZN(n4229) );
  INV_X1 U4623 ( .A(n3999), .ZN(n3980) );
  OAI21_X1 U4624 ( .B1(n3980), .B2(n3979), .A(n3978), .ZN(n4300) );
  NOR2_X1 U4625 ( .A1(n4300), .A2(n4169), .ZN(n3984) );
  INV_X1 U4626 ( .A(REG2_REG_24__SCAN_IN), .ZN(n3982) );
  OAI22_X1 U4627 ( .A1(n4195), .A2(n3982), .B1(n3981), .B2(n4193), .ZN(n3983)
         );
  AOI211_X1 U4628 ( .C1(n4229), .C2(n4195), .A(n3984), .B(n3983), .ZN(n3985)
         );
  OAI21_X1 U4629 ( .B1(n3986), .B2(n4172), .A(n3985), .ZN(U3266) );
  XOR2_X1 U4630 ( .A(n3992), .B(n3987), .Z(n4233) );
  INV_X1 U4631 ( .A(n4233), .ZN(n4006) );
  OR2_X1 U4632 ( .A1(n4026), .A2(n3988), .ZN(n3990) );
  NAND2_X1 U4633 ( .A1(n3990), .A2(n3989), .ZN(n4010) );
  NAND2_X1 U4634 ( .A1(n4010), .A2(n4011), .ZN(n4009) );
  NAND2_X1 U4635 ( .A1(n4009), .A2(n3991), .ZN(n3993) );
  XNOR2_X1 U4636 ( .A(n3993), .B(n3992), .ZN(n3998) );
  OAI22_X1 U4637 ( .A1(n3994), .A2(n4155), .B1(n4154), .B2(n4000), .ZN(n3995)
         );
  AOI21_X1 U4638 ( .B1(n4159), .B2(n3996), .A(n3995), .ZN(n3997) );
  OAI21_X1 U4639 ( .B1(n3998), .B2(n4161), .A(n3997), .ZN(n4232) );
  OAI21_X1 U4640 ( .B1(n4237), .B2(n4000), .A(n3999), .ZN(n4304) );
  NOR2_X1 U4641 ( .A1(n4304), .A2(n4169), .ZN(n4004) );
  INV_X1 U4642 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4002) );
  OAI22_X1 U4643 ( .A1(n4195), .A2(n4002), .B1(n4001), .B2(n4193), .ZN(n4003)
         );
  AOI211_X1 U4644 ( .C1(n4232), .C2(n4195), .A(n4004), .B(n4003), .ZN(n4005)
         );
  OAI21_X1 U4645 ( .B1(n4006), .B2(n4172), .A(n4005), .ZN(U3267) );
  OAI21_X1 U4646 ( .B1(n2197), .B2(n2196), .A(n4008), .ZN(n4240) );
  OAI21_X1 U4647 ( .B1(n4011), .B2(n4010), .A(n4009), .ZN(n4018) );
  NAND2_X1 U4648 ( .A1(n4012), .A2(n4450), .ZN(n4015) );
  NAND2_X1 U4649 ( .A1(n4013), .A2(n4159), .ZN(n4014) );
  OAI211_X1 U4650 ( .C1(n4016), .C2(n4155), .A(n4015), .B(n4014), .ZN(n4017)
         );
  AOI21_X1 U4651 ( .B1(n4018), .B2(n4281), .A(n4017), .ZN(n4239) );
  AOI22_X1 U4652 ( .A1(n2017), .A2(REG2_REG_22__SCAN_IN), .B1(n4019), .B2(
        n4459), .ZN(n4022) );
  NOR2_X1 U4653 ( .A1(n4035), .A2(n4020), .ZN(n4236) );
  OR3_X1 U4654 ( .A1(n4237), .A2(n4236), .A3(n4169), .ZN(n4021) );
  OAI211_X1 U4655 ( .C1(n4239), .C2(n2017), .A(n4022), .B(n4021), .ZN(n4023)
         );
  INV_X1 U4656 ( .A(n4023), .ZN(n4024) );
  OAI21_X1 U4657 ( .B1(n4240), .B2(n4172), .A(n4024), .ZN(U3268) );
  XOR2_X1 U4658 ( .A(n4027), .B(n4025), .Z(n4242) );
  INV_X1 U4659 ( .A(n4242), .ZN(n4041) );
  XOR2_X1 U4660 ( .A(n4027), .B(n4026), .Z(n4033) );
  OAI22_X1 U4661 ( .A1(n4029), .A2(n4155), .B1(n4154), .B2(n4028), .ZN(n4030)
         );
  AOI21_X1 U4662 ( .B1(n4159), .B2(n4031), .A(n4030), .ZN(n4032) );
  OAI21_X1 U4663 ( .B1(n4033), .B2(n4161), .A(n4032), .ZN(n4241) );
  AND2_X1 U4664 ( .A1(n4056), .A2(n4034), .ZN(n4036) );
  OR2_X1 U4665 ( .A1(n4036), .A2(n4035), .ZN(n4308) );
  AOI22_X1 U4666 ( .A1(n2017), .A2(REG2_REG_21__SCAN_IN), .B1(n4037), .B2(
        n4459), .ZN(n4038) );
  OAI21_X1 U4667 ( .B1(n4308), .B2(n4169), .A(n4038), .ZN(n4039) );
  AOI21_X1 U4668 ( .B1(n4241), .B2(n4195), .A(n4039), .ZN(n4040) );
  OAI21_X1 U4669 ( .B1(n4041), .B2(n4172), .A(n4040), .ZN(U3269) );
  XNOR2_X1 U4670 ( .A(n4042), .B(n4047), .ZN(n4053) );
  OAI22_X1 U4671 ( .A1(n4044), .A2(n4155), .B1(n4154), .B2(n4043), .ZN(n4051)
         );
  NAND2_X1 U4672 ( .A1(n4046), .A2(n4045), .ZN(n4048) );
  XNOR2_X1 U4673 ( .A(n4048), .B(n4047), .ZN(n4049) );
  NOR2_X1 U4674 ( .A1(n4049), .A2(n4161), .ZN(n4050) );
  AOI211_X1 U4675 ( .C1(n4159), .C2(n4090), .A(n4051), .B(n4050), .ZN(n4052)
         );
  OAI21_X1 U4676 ( .B1(n4053), .B2(n4455), .A(n4052), .ZN(n4244) );
  INV_X1 U4677 ( .A(n4244), .ZN(n4061) );
  INV_X1 U4678 ( .A(n4053), .ZN(n4245) );
  NAND2_X1 U4679 ( .A1(n4079), .A2(n4054), .ZN(n4055) );
  NAND2_X1 U4680 ( .A1(n4056), .A2(n4055), .ZN(n4312) );
  AOI22_X1 U4681 ( .A1(n2017), .A2(REG2_REG_20__SCAN_IN), .B1(n4057), .B2(
        n4459), .ZN(n4058) );
  OAI21_X1 U4682 ( .B1(n4312), .B2(n4169), .A(n4058), .ZN(n4059) );
  AOI21_X1 U4683 ( .B1(n4245), .B2(n4460), .A(n4059), .ZN(n4060) );
  OAI21_X1 U4684 ( .B1(n4061), .B2(n2017), .A(n4060), .ZN(U3270) );
  XNOR2_X1 U4685 ( .A(n4062), .B(n4070), .ZN(n4248) );
  INV_X1 U4686 ( .A(n4248), .ZN(n4084) );
  INV_X1 U4687 ( .A(n4063), .ZN(n4065) );
  OAI21_X1 U4688 ( .B1(n4104), .B2(n4065), .A(n4064), .ZN(n4088) );
  INV_X1 U4689 ( .A(n4066), .ZN(n4068) );
  OAI21_X1 U4690 ( .B1(n4088), .B2(n4068), .A(n4067), .ZN(n4069) );
  XOR2_X1 U4691 ( .A(n4070), .B(n4069), .Z(n4075) );
  OAI22_X1 U4692 ( .A1(n4071), .A2(n4155), .B1(n4154), .B2(n4076), .ZN(n4072)
         );
  AOI21_X1 U4693 ( .B1(n4159), .B2(n4073), .A(n4072), .ZN(n4074) );
  OAI21_X1 U4694 ( .B1(n4075), .B2(n4161), .A(n4074), .ZN(n4247) );
  OR2_X1 U4695 ( .A1(n4077), .A2(n4076), .ZN(n4078) );
  NAND2_X1 U4696 ( .A1(n4079), .A2(n4078), .ZN(n4316) );
  AOI22_X1 U4697 ( .A1(n2017), .A2(REG2_REG_19__SCAN_IN), .B1(n4080), .B2(
        n4459), .ZN(n4081) );
  OAI21_X1 U4698 ( .B1(n4316), .B2(n4169), .A(n4081), .ZN(n4082) );
  AOI21_X1 U4699 ( .B1(n4247), .B2(n4195), .A(n4082), .ZN(n4083) );
  OAI21_X1 U4700 ( .B1(n4084), .B2(n4172), .A(n4083), .ZN(U3271) );
  OAI21_X1 U4701 ( .B1(n4086), .B2(n4089), .A(n4085), .ZN(n4087) );
  INV_X1 U4702 ( .A(n4087), .ZN(n4253) );
  XOR2_X1 U4703 ( .A(n4089), .B(n4088), .Z(n4093) );
  AOI22_X1 U4704 ( .A1(n4090), .A2(n4280), .B1(n4094), .B2(n4450), .ZN(n4091)
         );
  OAI21_X1 U4705 ( .B1(n4129), .B2(n4184), .A(n4091), .ZN(n4092) );
  AOI21_X1 U4706 ( .B1(n4093), .B2(n4281), .A(n4092), .ZN(n4252) );
  INV_X1 U4707 ( .A(n4252), .ZN(n4101) );
  XNOR2_X1 U4708 ( .A(n4110), .B(n4094), .ZN(n4095) );
  NAND2_X1 U4709 ( .A1(n4095), .A2(n4502), .ZN(n4251) );
  INV_X1 U4710 ( .A(n4096), .ZN(n4099) );
  AOI22_X1 U4711 ( .A1(n2017), .A2(REG2_REG_18__SCAN_IN), .B1(n4097), .B2(
        n4459), .ZN(n4098) );
  OAI21_X1 U4712 ( .B1(n4251), .B2(n4099), .A(n4098), .ZN(n4100) );
  AOI21_X1 U4713 ( .B1(n4101), .B2(n4195), .A(n4100), .ZN(n4102) );
  OAI21_X1 U4714 ( .B1(n4253), .B2(n4172), .A(n4102), .ZN(U3272) );
  XOR2_X1 U4715 ( .A(n4105), .B(n4103), .Z(n4255) );
  INV_X1 U4716 ( .A(n4255), .ZN(n4117) );
  XOR2_X1 U4717 ( .A(n4105), .B(n4104), .Z(n4109) );
  OAI22_X1 U4718 ( .A1(n4106), .A2(n4155), .B1(n4154), .B2(n4112), .ZN(n4107)
         );
  AOI21_X1 U4719 ( .B1(n4159), .B2(n4140), .A(n4107), .ZN(n4108) );
  OAI21_X1 U4720 ( .B1(n4109), .B2(n4161), .A(n4108), .ZN(n4254) );
  INV_X1 U4721 ( .A(n4110), .ZN(n4111) );
  OAI21_X1 U4722 ( .B1(n2918), .B2(n4112), .A(n4111), .ZN(n4321) );
  AOI22_X1 U4723 ( .A1(n2017), .A2(REG2_REG_17__SCAN_IN), .B1(n4113), .B2(
        n4459), .ZN(n4114) );
  OAI21_X1 U4724 ( .B1(n4321), .B2(n4169), .A(n4114), .ZN(n4115) );
  AOI21_X1 U4725 ( .B1(n4254), .B2(n4195), .A(n4115), .ZN(n4116) );
  OAI21_X1 U4726 ( .B1(n4117), .B2(n4172), .A(n4116), .ZN(U3273) );
  OAI21_X1 U4727 ( .B1(n4120), .B2(n4119), .A(n4118), .ZN(n4260) );
  AOI21_X1 U4728 ( .B1(n4122), .B2(n4121), .A(n2918), .ZN(n4258) );
  INV_X1 U4729 ( .A(n4123), .ZN(n4124) );
  OAI22_X1 U4730 ( .A1(n4195), .A2(n4419), .B1(n4124), .B2(n4193), .ZN(n4125)
         );
  AOI21_X1 U4731 ( .B1(n4258), .B2(n4444), .A(n4125), .ZN(n4134) );
  OAI211_X1 U4732 ( .C1(n4127), .C2(n2189), .A(n4126), .B(n4281), .ZN(n4132)
         );
  OAI22_X1 U4733 ( .A1(n4129), .A2(n4155), .B1(n4128), .B2(n4154), .ZN(n4130)
         );
  INV_X1 U4734 ( .A(n4130), .ZN(n4131) );
  OAI211_X1 U4735 ( .C1(n4156), .C2(n4184), .A(n4132), .B(n4131), .ZN(n4257)
         );
  NAND2_X1 U4736 ( .A1(n4257), .A2(n4195), .ZN(n4133) );
  OAI211_X1 U4737 ( .C1(n4260), .C2(n4172), .A(n4134), .B(n4133), .ZN(U3274)
         );
  XNOR2_X1 U4738 ( .A(n4135), .B(n4138), .ZN(n4264) );
  INV_X1 U4739 ( .A(n4136), .ZN(n4139) );
  OAI211_X1 U4740 ( .C1(n4139), .C2(n4138), .A(n4281), .B(n4137), .ZN(n4142)
         );
  AOI22_X1 U4741 ( .A1(n4140), .A2(n4280), .B1(n4450), .B2(n4144), .ZN(n4141)
         );
  OAI211_X1 U4742 ( .C1(n4143), .C2(n4184), .A(n4142), .B(n4141), .ZN(n4261)
         );
  XNOR2_X1 U4743 ( .A(n4163), .B(n4144), .ZN(n4262) );
  INV_X1 U4744 ( .A(n4262), .ZN(n4147) );
  AOI22_X1 U4745 ( .A1(n2017), .A2(REG2_REG_15__SCAN_IN), .B1(n4145), .B2(
        n4459), .ZN(n4146) );
  OAI21_X1 U4746 ( .B1(n4147), .B2(n4169), .A(n4146), .ZN(n4148) );
  AOI21_X1 U4747 ( .B1(n4261), .B2(n4195), .A(n4148), .ZN(n4149) );
  OAI21_X1 U4748 ( .B1(n4264), .B2(n4172), .A(n4149), .ZN(U3275) );
  OAI21_X1 U4749 ( .B1(n4151), .B2(n4152), .A(n4150), .ZN(n4266) );
  INV_X1 U4750 ( .A(n4266), .ZN(n4173) );
  XNOR2_X1 U4751 ( .A(n4153), .B(n4152), .ZN(n4162) );
  OAI22_X1 U4752 ( .A1(n4156), .A2(n4155), .B1(n4165), .B2(n4154), .ZN(n4157)
         );
  AOI21_X1 U4753 ( .B1(n4159), .B2(n4158), .A(n4157), .ZN(n4160) );
  OAI21_X1 U4754 ( .B1(n4162), .B2(n4161), .A(n4160), .ZN(n4265) );
  INV_X1 U4755 ( .A(n4190), .ZN(n4166) );
  INV_X1 U4756 ( .A(n4163), .ZN(n4164) );
  OAI21_X1 U4757 ( .B1(n4166), .B2(n4165), .A(n4164), .ZN(n4327) );
  AOI22_X1 U4758 ( .A1(n2017), .A2(REG2_REG_14__SCAN_IN), .B1(n4167), .B2(
        n4459), .ZN(n4168) );
  OAI21_X1 U4759 ( .B1(n4327), .B2(n4169), .A(n4168), .ZN(n4170) );
  AOI21_X1 U4760 ( .B1(n4265), .B2(n4195), .A(n4170), .ZN(n4171) );
  OAI21_X1 U4761 ( .B1(n4173), .B2(n4172), .A(n4171), .ZN(U3276) );
  XNOR2_X1 U4762 ( .A(n4174), .B(n4180), .ZN(n4268) );
  INV_X1 U4763 ( .A(n4175), .ZN(n4176) );
  AOI21_X1 U4764 ( .B1(n4178), .B2(n4177), .A(n4176), .ZN(n4179) );
  XOR2_X1 U4765 ( .A(n4180), .B(n4179), .Z(n4187) );
  AOI22_X1 U4766 ( .A1(n4182), .A2(n4280), .B1(n4450), .B2(n4181), .ZN(n4183)
         );
  OAI21_X1 U4767 ( .B1(n4185), .B2(n4184), .A(n4183), .ZN(n4186) );
  AOI21_X1 U4768 ( .B1(n4187), .B2(n4281), .A(n4186), .ZN(n4188) );
  OAI21_X1 U4769 ( .B1(n4268), .B2(n4455), .A(n4188), .ZN(n4269) );
  NAND2_X1 U4770 ( .A1(n4269), .A2(n4195), .ZN(n4199) );
  INV_X1 U4771 ( .A(n4189), .ZN(n4192) );
  OAI21_X1 U4772 ( .B1(n4192), .B2(n4191), .A(n4190), .ZN(n4331) );
  INV_X1 U4773 ( .A(n4331), .ZN(n4197) );
  OAI22_X1 U4774 ( .A1(n4195), .A2(n4395), .B1(n4194), .B2(n4193), .ZN(n4196)
         );
  AOI21_X1 U4775 ( .B1(n4197), .B2(n4444), .A(n4196), .ZN(n4198) );
  OAI211_X1 U4776 ( .C1(n4268), .C2(n4200), .A(n4199), .B(n4198), .ZN(U3277)
         );
  NAND2_X1 U4777 ( .A1(n4208), .A2(n4209), .ZN(n4207) );
  XNOR2_X1 U4778 ( .A(n4207), .B(n4201), .ZN(n4352) );
  INV_X1 U4779 ( .A(n4352), .ZN(n4286) );
  INV_X1 U4780 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4205) );
  AND2_X1 U4781 ( .A1(n4203), .A2(n4202), .ZN(n4210) );
  AOI21_X1 U4782 ( .B1(n4204), .B2(n4450), .A(n4210), .ZN(n4354) );
  MUX2_X1 U4783 ( .A(n4205), .B(n4354), .S(n4533), .Z(n4206) );
  OAI21_X1 U4784 ( .B1(n4286), .B2(n4278), .A(n4206), .ZN(U3549) );
  OAI21_X1 U4785 ( .B1(n4208), .B2(n4209), .A(n4207), .ZN(n4355) );
  INV_X1 U4786 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4212) );
  INV_X1 U4787 ( .A(n4209), .ZN(n4211) );
  AOI21_X1 U4788 ( .B1(n4211), .B2(n4450), .A(n4210), .ZN(n4358) );
  MUX2_X1 U4789 ( .A(n4212), .B(n4358), .S(n4533), .Z(n4213) );
  OAI21_X1 U4790 ( .B1(n4355), .B2(n4278), .A(n4213), .ZN(U3548) );
  NAND2_X1 U4791 ( .A1(n4217), .A2(n4513), .ZN(n4219) );
  OAI211_X1 U4792 ( .C1(n2101), .C2(n4220), .A(n4219), .B(n4218), .ZN(n4289)
         );
  MUX2_X1 U4793 ( .A(REG1_REG_27__SCAN_IN), .B(n4289), .S(n4533), .Z(U3545) );
  INV_X1 U4794 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4223) );
  AOI21_X1 U4795 ( .B1(n4222), .B2(n4513), .A(n4221), .ZN(n4290) );
  MUX2_X1 U4796 ( .A(n4223), .B(n4290), .S(n4533), .Z(n4224) );
  OAI21_X1 U4797 ( .B1(n4278), .B2(n4293), .A(n4224), .ZN(U3544) );
  INV_X1 U4798 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4227) );
  AOI21_X1 U4799 ( .B1(n4226), .B2(n4513), .A(n4225), .ZN(n4294) );
  MUX2_X1 U4800 ( .A(n4227), .B(n4294), .S(n4533), .Z(n4228) );
  OAI21_X1 U4801 ( .B1(n4278), .B2(n4297), .A(n4228), .ZN(U3543) );
  INV_X1 U4802 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4550) );
  AOI21_X1 U4803 ( .B1(n4230), .B2(n4513), .A(n4229), .ZN(n4298) );
  MUX2_X1 U4804 ( .A(n4550), .B(n4298), .S(n4533), .Z(n4231) );
  OAI21_X1 U4805 ( .B1(n4278), .B2(n4300), .A(n4231), .ZN(U3542) );
  INV_X1 U4806 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4234) );
  AOI21_X1 U4807 ( .B1(n4233), .B2(n4513), .A(n4232), .ZN(n4301) );
  MUX2_X1 U4808 ( .A(n4234), .B(n4301), .S(n4533), .Z(n4235) );
  OAI21_X1 U4809 ( .B1(n4278), .B2(n4304), .A(n4235), .ZN(U3541) );
  OR3_X1 U4810 ( .A1(n4237), .A2(n4236), .A3(n2101), .ZN(n4238) );
  OAI211_X1 U4811 ( .C1(n4240), .C2(n4496), .A(n4239), .B(n4238), .ZN(n4305)
         );
  MUX2_X1 U4812 ( .A(REG1_REG_22__SCAN_IN), .B(n4305), .S(n4533), .Z(U3540) );
  INV_X1 U4813 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4551) );
  AOI21_X1 U4814 ( .B1(n4242), .B2(n4513), .A(n4241), .ZN(n4306) );
  MUX2_X1 U4815 ( .A(n4551), .B(n4306), .S(n4533), .Z(n4243) );
  OAI21_X1 U4816 ( .B1(n4278), .B2(n4308), .A(n4243), .ZN(U3539) );
  INV_X1 U4817 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4611) );
  AOI21_X1 U4818 ( .B1(n4520), .B2(n4245), .A(n4244), .ZN(n4309) );
  MUX2_X1 U4819 ( .A(n4611), .B(n4309), .S(n4533), .Z(n4246) );
  OAI21_X1 U4820 ( .B1(n4278), .B2(n4312), .A(n4246), .ZN(U3538) );
  INV_X1 U4821 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4249) );
  AOI21_X1 U4822 ( .B1(n4248), .B2(n4513), .A(n4247), .ZN(n4313) );
  MUX2_X1 U4823 ( .A(n4249), .B(n4313), .S(n4533), .Z(n4250) );
  OAI21_X1 U4824 ( .B1(n4278), .B2(n4316), .A(n4250), .ZN(U3537) );
  OAI211_X1 U4825 ( .C1(n4253), .C2(n4496), .A(n4252), .B(n4251), .ZN(n4317)
         );
  MUX2_X1 U4826 ( .A(REG1_REG_18__SCAN_IN), .B(n4317), .S(n4533), .Z(U3536) );
  AOI21_X1 U4827 ( .B1(n4255), .B2(n4513), .A(n4254), .ZN(n4318) );
  MUX2_X1 U4828 ( .A(n4596), .B(n4318), .S(n4533), .Z(n4256) );
  OAI21_X1 U4829 ( .B1(n4278), .B2(n4321), .A(n4256), .ZN(U3535) );
  AOI21_X1 U4830 ( .B1(n4502), .B2(n4258), .A(n4257), .ZN(n4259) );
  OAI21_X1 U4831 ( .B1(n4260), .B2(n4496), .A(n4259), .ZN(n4322) );
  MUX2_X1 U4832 ( .A(REG1_REG_16__SCAN_IN), .B(n4322), .S(n4533), .Z(U3534) );
  AOI21_X1 U4833 ( .B1(n4502), .B2(n4262), .A(n4261), .ZN(n4263) );
  OAI21_X1 U4834 ( .B1(n4264), .B2(n4496), .A(n4263), .ZN(n4323) );
  MUX2_X1 U4835 ( .A(REG1_REG_15__SCAN_IN), .B(n4323), .S(n4533), .Z(U3533) );
  AOI21_X1 U4836 ( .B1(n4266), .B2(n4513), .A(n4265), .ZN(n4324) );
  MUX2_X1 U4837 ( .A(n4404), .B(n4324), .S(n4533), .Z(n4267) );
  OAI21_X1 U4838 ( .B1(n4278), .B2(n4327), .A(n4267), .ZN(U3532) );
  INV_X1 U4839 ( .A(n4268), .ZN(n4270) );
  AOI21_X1 U4840 ( .B1(n4520), .B2(n4270), .A(n4269), .ZN(n4328) );
  MUX2_X1 U4841 ( .A(n4271), .B(n4328), .S(n4533), .Z(n4272) );
  OAI21_X1 U4842 ( .B1(n4278), .B2(n4331), .A(n4272), .ZN(U3531) );
  NAND2_X1 U4843 ( .A1(n4273), .A2(n4513), .ZN(n4275) );
  NAND2_X1 U4844 ( .A1(n4275), .A2(n4274), .ZN(n4332) );
  MUX2_X1 U4845 ( .A(n4332), .B(REG1_REG_12__SCAN_IN), .S(n4530), .Z(n4276) );
  INV_X1 U4846 ( .A(n4276), .ZN(n4277) );
  OAI21_X1 U4847 ( .B1(n4278), .B2(n4336), .A(n4277), .ZN(U3530) );
  INV_X1 U4848 ( .A(n4456), .ZN(n4461) );
  AOI22_X1 U4849 ( .A1(n4461), .A2(n4281), .B1(n4280), .B2(n4279), .ZN(n4449)
         );
  NAND2_X1 U4850 ( .A1(n4282), .A2(n4452), .ZN(n4283) );
  OAI211_X1 U4851 ( .C1(n4496), .C2(n4456), .A(n4449), .B(n4283), .ZN(n4691)
         );
  MUX2_X1 U4852 ( .A(REG1_REG_0__SCAN_IN), .B(n4691), .S(n4533), .Z(U3518) );
  INV_X1 U4853 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4284) );
  MUX2_X1 U4854 ( .A(n4284), .B(n4354), .S(n4692), .Z(n4285) );
  OAI21_X1 U4855 ( .B1(n4286), .B2(n4335), .A(n4285), .ZN(U3517) );
  INV_X1 U4856 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4287) );
  MUX2_X1 U4857 ( .A(n4287), .B(n4358), .S(n4692), .Z(n4288) );
  OAI21_X1 U4858 ( .B1(n4355), .B2(n4335), .A(n4288), .ZN(U3516) );
  MUX2_X1 U4859 ( .A(REG0_REG_27__SCAN_IN), .B(n4289), .S(n4692), .Z(U3513) );
  INV_X1 U4860 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4291) );
  MUX2_X1 U4861 ( .A(n4291), .B(n4290), .S(n4692), .Z(n4292) );
  OAI21_X1 U4862 ( .B1(n4293), .B2(n4335), .A(n4292), .ZN(U3512) );
  INV_X1 U4863 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4295) );
  MUX2_X1 U4864 ( .A(n4295), .B(n4294), .S(n4692), .Z(n4296) );
  OAI21_X1 U4865 ( .B1(n4297), .B2(n4335), .A(n4296), .ZN(U3511) );
  INV_X1 U4866 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4553) );
  MUX2_X1 U4867 ( .A(n4553), .B(n4298), .S(n4692), .Z(n4299) );
  OAI21_X1 U4868 ( .B1(n4300), .B2(n4335), .A(n4299), .ZN(U3510) );
  INV_X1 U4869 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4302) );
  MUX2_X1 U4870 ( .A(n4302), .B(n4301), .S(n4692), .Z(n4303) );
  OAI21_X1 U4871 ( .B1(n4304), .B2(n4335), .A(n4303), .ZN(U3509) );
  MUX2_X1 U4872 ( .A(REG0_REG_22__SCAN_IN), .B(n4305), .S(n4692), .Z(U3508) );
  INV_X1 U4873 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4554) );
  MUX2_X1 U4874 ( .A(n4554), .B(n4306), .S(n4692), .Z(n4307) );
  OAI21_X1 U4875 ( .B1(n4308), .B2(n4335), .A(n4307), .ZN(U3507) );
  INV_X1 U4876 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4310) );
  MUX2_X1 U4877 ( .A(n4310), .B(n4309), .S(n4692), .Z(n4311) );
  OAI21_X1 U4878 ( .B1(n4312), .B2(n4335), .A(n4311), .ZN(U3506) );
  INV_X1 U4879 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4314) );
  MUX2_X1 U4880 ( .A(n4314), .B(n4313), .S(n4692), .Z(n4315) );
  OAI21_X1 U4881 ( .B1(n4316), .B2(n4335), .A(n4315), .ZN(U3505) );
  MUX2_X1 U4882 ( .A(REG0_REG_18__SCAN_IN), .B(n4317), .S(n4692), .Z(U3503) );
  INV_X1 U4883 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4319) );
  MUX2_X1 U4884 ( .A(n4319), .B(n4318), .S(n4692), .Z(n4320) );
  OAI21_X1 U4885 ( .B1(n4321), .B2(n4335), .A(n4320), .ZN(U3501) );
  MUX2_X1 U4886 ( .A(REG0_REG_16__SCAN_IN), .B(n4322), .S(n4692), .Z(U3499) );
  MUX2_X1 U4887 ( .A(REG0_REG_15__SCAN_IN), .B(n4323), .S(n4692), .Z(U3497) );
  INV_X1 U4888 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4325) );
  MUX2_X1 U4889 ( .A(n4325), .B(n4324), .S(n4692), .Z(n4326) );
  OAI21_X1 U4890 ( .B1(n4327), .B2(n4335), .A(n4326), .ZN(U3495) );
  INV_X1 U4891 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4329) );
  MUX2_X1 U4892 ( .A(n4329), .B(n4328), .S(n4692), .Z(n4330) );
  OAI21_X1 U4893 ( .B1(n4331), .B2(n4335), .A(n4330), .ZN(U3493) );
  MUX2_X1 U4894 ( .A(n4332), .B(REG0_REG_12__SCAN_IN), .S(n4690), .Z(n4333) );
  INV_X1 U4895 ( .A(n4333), .ZN(n4334) );
  OAI21_X1 U4896 ( .B1(n4336), .B2(n4335), .A(n4334), .ZN(U3491) );
  MUX2_X1 U4897 ( .A(n4337), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U4898 ( .A(n4338), .B(DATAI_27_), .S(U3149), .Z(U3325) );
  MUX2_X1 U4899 ( .A(n4339), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U4900 ( .A(DATAI_24_), .B(n4340), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U4901 ( .A(DATAI_22_), .B(n4341), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4902 ( .A(DATAI_19_), .B(n4342), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U4903 ( .A(n4343), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U4904 ( .A(DATAI_7_), .B(n4344), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U4905 ( .A(n4345), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4906 ( .A(n4346), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4907 ( .A(DATAI_4_), .B(n4347), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4908 ( .A(n4348), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4909 ( .A(n4349), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U4910 ( .A(DATAI_28_), .ZN(n4350) );
  AOI22_X1 U4911 ( .A1(STATE_REG_SCAN_IN), .A2(n4351), .B1(n4350), .B2(U3149), 
        .ZN(U3324) );
  AOI22_X1 U4912 ( .A1(n4352), .A2(n4444), .B1(n2017), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n4353) );
  OAI21_X1 U4913 ( .B1(n2017), .B2(n4354), .A(n4353), .ZN(U3260) );
  INV_X1 U4914 ( .A(n4355), .ZN(n4356) );
  OAI21_X1 U4915 ( .B1(n2017), .B2(n4358), .A(n4357), .ZN(U3261) );
  AOI211_X1 U4916 ( .C1(n4361), .C2(n4360), .A(n4359), .B(n4401), .ZN(n4363)
         );
  AOI211_X1 U4917 ( .C1(n4429), .C2(ADDR_REG_9__SCAN_IN), .A(n4363), .B(n4362), 
        .ZN(n4368) );
  OAI211_X1 U4918 ( .C1(n4366), .C2(n4365), .A(n4439), .B(n4364), .ZN(n4367)
         );
  OAI211_X1 U4919 ( .C1(n4442), .C2(n4478), .A(n4368), .B(n4367), .ZN(U3249)
         );
  AOI211_X1 U4920 ( .C1(n4371), .C2(n4370), .A(n4369), .B(n4401), .ZN(n4373)
         );
  AOI211_X1 U4921 ( .C1(n4429), .C2(ADDR_REG_11__SCAN_IN), .A(n4373), .B(n4372), .ZN(n4378) );
  OAI211_X1 U4922 ( .C1(n4376), .C2(n4375), .A(n4439), .B(n4374), .ZN(n4377)
         );
  OAI211_X1 U4923 ( .C1(n4442), .C2(n4379), .A(n4378), .B(n4377), .ZN(U3251)
         );
  AOI211_X1 U4924 ( .C1(n4382), .C2(n4381), .A(n4380), .B(n4401), .ZN(n4385)
         );
  INV_X1 U4925 ( .A(n4383), .ZN(n4384) );
  AOI211_X1 U4926 ( .C1(n4429), .C2(ADDR_REG_12__SCAN_IN), .A(n4385), .B(n4384), .ZN(n4389) );
  OAI211_X1 U4927 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4387), .A(n4439), .B(n4386), .ZN(n4388) );
  OAI211_X1 U4928 ( .C1(n4442), .C2(n2167), .A(n4389), .B(n4388), .ZN(U3252)
         );
  AOI211_X1 U4929 ( .C1(n2049), .C2(n4391), .A(n4390), .B(n4401), .ZN(n4392)
         );
  AOI211_X1 U4930 ( .C1(n4429), .C2(ADDR_REG_13__SCAN_IN), .A(n4393), .B(n4392), .ZN(n4400) );
  AOI21_X1 U4931 ( .B1(n4395), .B2(n4473), .A(n4394), .ZN(n4398) );
  AOI21_X1 U4932 ( .B1(n4398), .B2(n4397), .A(n4405), .ZN(n4396) );
  OAI21_X1 U4933 ( .B1(n4398), .B2(n4397), .A(n4396), .ZN(n4399) );
  OAI211_X1 U4934 ( .C1(n4442), .C2(n4473), .A(n4400), .B(n4399), .ZN(U3253)
         );
  NAND2_X1 U4935 ( .A1(ADDR_REG_14__SCAN_IN), .A2(n4429), .ZN(n4415) );
  AOI211_X1 U4936 ( .C1(n4404), .C2(n4403), .A(n4402), .B(n4401), .ZN(n4410)
         );
  AOI211_X1 U4937 ( .C1(n4408), .C2(n4407), .A(n4406), .B(n4405), .ZN(n4409)
         );
  AOI211_X1 U4938 ( .C1(n4412), .C2(n4411), .A(n4410), .B(n4409), .ZN(n4414)
         );
  NAND3_X1 U4939 ( .A1(n4415), .A2(n4414), .A3(n4413), .ZN(U3254) );
  INV_X1 U4940 ( .A(n4416), .ZN(n4417) );
  AOI21_X1 U4941 ( .B1(n4429), .B2(ADDR_REG_16__SCAN_IN), .A(n4417), .ZN(n4427) );
  OAI21_X1 U4942 ( .B1(n4420), .B2(n4419), .A(n4418), .ZN(n4425) );
  OAI21_X1 U4943 ( .B1(n4423), .B2(n4422), .A(n4421), .ZN(n4424) );
  AOI22_X1 U4944 ( .A1(n4439), .A2(n4425), .B1(n4437), .B2(n4424), .ZN(n4426)
         );
  OAI211_X1 U4945 ( .C1(n4470), .C2(n4442), .A(n4427), .B(n4426), .ZN(U3256)
         );
  AOI21_X1 U4946 ( .B1(n4429), .B2(ADDR_REG_17__SCAN_IN), .A(n4428), .ZN(n4441) );
  OAI21_X1 U4947 ( .B1(n4432), .B2(n4431), .A(n4430), .ZN(n4438) );
  OAI21_X1 U4948 ( .B1(n4435), .B2(n4434), .A(n4433), .ZN(n4436) );
  AOI22_X1 U4949 ( .A1(n4439), .A2(n4438), .B1(n4437), .B2(n4436), .ZN(n4440)
         );
  OAI211_X1 U4950 ( .C1(n4468), .C2(n4442), .A(n4441), .B(n4440), .ZN(U3257)
         );
  AOI22_X1 U4951 ( .A1(REG3_REG_2__SCAN_IN), .A2(n4459), .B1(
        REG2_REG_2__SCAN_IN), .B2(n2017), .ZN(n4447) );
  AOI22_X1 U4952 ( .A1(n4445), .A2(n4460), .B1(n4444), .B2(n4443), .ZN(n4446)
         );
  OAI211_X1 U4953 ( .C1(n2017), .C2(n4448), .A(n4447), .B(n4446), .ZN(U3288)
         );
  INV_X1 U4954 ( .A(n4449), .ZN(n4458) );
  AOI21_X1 U4955 ( .B1(n4452), .B2(n4451), .A(n4450), .ZN(n4454) );
  OAI22_X1 U4956 ( .A1(n4456), .A2(n4455), .B1(n4454), .B2(n4453), .ZN(n4457)
         );
  NOR2_X1 U4957 ( .A1(n4458), .A2(n4457), .ZN(n4463) );
  AOI22_X1 U4958 ( .A1(n4461), .A2(n4460), .B1(REG3_REG_0__SCAN_IN), .B2(n4459), .ZN(n4462) );
  OAI221_X1 U4959 ( .B1(n2017), .B2(n4463), .C1(n4195), .C2(n2281), .A(n4462), 
        .ZN(U3290) );
  AND2_X1 U4960 ( .A1(D_REG_31__SCAN_IN), .A2(n4464), .ZN(U3291) );
  AND2_X1 U4961 ( .A1(D_REG_30__SCAN_IN), .A2(n4464), .ZN(U3292) );
  AND2_X1 U4962 ( .A1(D_REG_29__SCAN_IN), .A2(n4464), .ZN(U3293) );
  AND2_X1 U4963 ( .A1(D_REG_28__SCAN_IN), .A2(n4464), .ZN(U3294) );
  AND2_X1 U4964 ( .A1(D_REG_27__SCAN_IN), .A2(n4464), .ZN(U3295) );
  AND2_X1 U4965 ( .A1(D_REG_26__SCAN_IN), .A2(n4464), .ZN(U3296) );
  INV_X1 U4966 ( .A(D_REG_25__SCAN_IN), .ZN(n4539) );
  NOR2_X1 U4967 ( .A1(n4465), .A2(n4539), .ZN(U3297) );
  AND2_X1 U4968 ( .A1(D_REG_24__SCAN_IN), .A2(n4464), .ZN(U3298) );
  INV_X1 U4969 ( .A(D_REG_23__SCAN_IN), .ZN(n4543) );
  NOR2_X1 U4970 ( .A1(n4465), .A2(n4543), .ZN(U3299) );
  AND2_X1 U4971 ( .A1(D_REG_22__SCAN_IN), .A2(n4464), .ZN(U3300) );
  AND2_X1 U4972 ( .A1(D_REG_21__SCAN_IN), .A2(n4464), .ZN(U3301) );
  AND2_X1 U4973 ( .A1(D_REG_20__SCAN_IN), .A2(n4464), .ZN(U3302) );
  AND2_X1 U4974 ( .A1(D_REG_19__SCAN_IN), .A2(n4464), .ZN(U3303) );
  INV_X1 U4975 ( .A(D_REG_18__SCAN_IN), .ZN(n4536) );
  NOR2_X1 U4976 ( .A1(n4465), .A2(n4536), .ZN(U3304) );
  AND2_X1 U4977 ( .A1(D_REG_17__SCAN_IN), .A2(n4464), .ZN(U3305) );
  INV_X1 U4978 ( .A(D_REG_16__SCAN_IN), .ZN(n4535) );
  NOR2_X1 U4979 ( .A1(n4465), .A2(n4535), .ZN(U3306) );
  AND2_X1 U4980 ( .A1(D_REG_15__SCAN_IN), .A2(n4464), .ZN(U3307) );
  AND2_X1 U4981 ( .A1(D_REG_14__SCAN_IN), .A2(n4464), .ZN(U3308) );
  AND2_X1 U4982 ( .A1(D_REG_13__SCAN_IN), .A2(n4464), .ZN(U3309) );
  AND2_X1 U4983 ( .A1(D_REG_12__SCAN_IN), .A2(n4464), .ZN(U3310) );
  AND2_X1 U4984 ( .A1(D_REG_11__SCAN_IN), .A2(n4464), .ZN(U3311) );
  AND2_X1 U4985 ( .A1(D_REG_10__SCAN_IN), .A2(n4464), .ZN(U3312) );
  AND2_X1 U4986 ( .A1(D_REG_9__SCAN_IN), .A2(n4464), .ZN(U3313) );
  AND2_X1 U4987 ( .A1(D_REG_8__SCAN_IN), .A2(n4464), .ZN(U3314) );
  AND2_X1 U4988 ( .A1(D_REG_7__SCAN_IN), .A2(n4464), .ZN(U3315) );
  INV_X1 U4989 ( .A(D_REG_6__SCAN_IN), .ZN(n4544) );
  NOR2_X1 U4990 ( .A1(n4465), .A2(n4544), .ZN(U3316) );
  AND2_X1 U4991 ( .A1(D_REG_5__SCAN_IN), .A2(n4464), .ZN(U3317) );
  INV_X1 U4992 ( .A(D_REG_4__SCAN_IN), .ZN(n4538) );
  NOR2_X1 U4993 ( .A1(n4465), .A2(n4538), .ZN(U3318) );
  AND2_X1 U4994 ( .A1(D_REG_3__SCAN_IN), .A2(n4464), .ZN(U3319) );
  INV_X1 U4995 ( .A(D_REG_2__SCAN_IN), .ZN(n4541) );
  NOR2_X1 U4996 ( .A1(n4465), .A2(n4541), .ZN(U3320) );
  INV_X1 U4997 ( .A(DATAI_23_), .ZN(n4467) );
  AOI21_X1 U4998 ( .B1(U3149), .B2(n4467), .A(n4466), .ZN(U3329) );
  AOI22_X1 U4999 ( .A1(STATE_REG_SCAN_IN), .A2(n4468), .B1(n2587), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5000 ( .A(DATAI_16_), .ZN(n4469) );
  AOI22_X1 U5001 ( .A1(STATE_REG_SCAN_IN), .A2(n4470), .B1(n4469), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5002 ( .A(DATAI_14_), .ZN(n4471) );
  AOI22_X1 U5003 ( .A1(STATE_REG_SCAN_IN), .A2(n4472), .B1(n4471), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5004 ( .A1(STATE_REG_SCAN_IN), .A2(n4473), .B1(n2522), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5005 ( .A(DATAI_12_), .ZN(n4474) );
  AOI22_X1 U5006 ( .A1(STATE_REG_SCAN_IN), .A2(n2167), .B1(n4474), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5007 ( .A1(U3149), .A2(n4475), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4476) );
  INV_X1 U5008 ( .A(n4476), .ZN(U3341) );
  INV_X1 U5009 ( .A(DATAI_9_), .ZN(n4477) );
  AOI22_X1 U5010 ( .A1(STATE_REG_SCAN_IN), .A2(n4478), .B1(n4477), .B2(U3149), 
        .ZN(U3343) );
  AOI22_X1 U5011 ( .A1(STATE_REG_SCAN_IN), .A2(n2146), .B1(n2145), .B2(U3149), 
        .ZN(U3352) );
  OAI22_X1 U5012 ( .A1(n4481), .A2(n4480), .B1(n2101), .B2(n4479), .ZN(n4482)
         );
  NOR2_X1 U5013 ( .A1(n4483), .A2(n4482), .ZN(n4521) );
  INV_X1 U5014 ( .A(REG0_REG_1__SCAN_IN), .ZN(n4484) );
  AOI22_X1 U5015 ( .A1(n4692), .A2(n4521), .B1(n4484), .B2(n4690), .ZN(U3469)
         );
  NOR2_X1 U5016 ( .A1(n4485), .A2(n2101), .ZN(n4486) );
  AOI21_X1 U5017 ( .B1(n4487), .B2(n4520), .A(n4486), .ZN(n4488) );
  AND2_X1 U5018 ( .A1(n4489), .A2(n4488), .ZN(n4523) );
  INV_X1 U5019 ( .A(REG0_REG_3__SCAN_IN), .ZN(n4490) );
  AOI22_X1 U5020 ( .A1(n4692), .A2(n4523), .B1(n4490), .B2(n4690), .ZN(U3473)
         );
  INV_X1 U5021 ( .A(n4491), .ZN(n4493) );
  AOI211_X1 U5022 ( .C1(n4494), .C2(n4520), .A(n4493), .B(n4492), .ZN(n4524)
         );
  INV_X1 U5023 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4495) );
  AOI22_X1 U5024 ( .A1(n4692), .A2(n4524), .B1(n4495), .B2(n4690), .ZN(U3475)
         );
  NOR2_X1 U5025 ( .A1(n4497), .A2(n4496), .ZN(n4500) );
  INV_X1 U5026 ( .A(n4498), .ZN(n4499) );
  AOI211_X1 U5027 ( .C1(n4502), .C2(n4501), .A(n4500), .B(n4499), .ZN(n4526)
         );
  INV_X1 U5028 ( .A(REG0_REG_5__SCAN_IN), .ZN(n4503) );
  AOI22_X1 U5029 ( .A1(n4692), .A2(n4526), .B1(n4503), .B2(n4690), .ZN(U3477)
         );
  NAND3_X1 U5030 ( .A1(n4505), .A2(n4513), .A3(n4504), .ZN(n4507) );
  AND3_X1 U5031 ( .A1(n4508), .A2(n4507), .A3(n4506), .ZN(n4527) );
  INV_X1 U5032 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4509) );
  AOI22_X1 U5033 ( .A1(n4692), .A2(n4527), .B1(n4509), .B2(n4690), .ZN(U3481)
         );
  OAI21_X1 U5034 ( .B1(n2101), .B2(n4511), .A(n4510), .ZN(n4512) );
  AOI21_X1 U5035 ( .B1(n4514), .B2(n4513), .A(n4512), .ZN(n4529) );
  INV_X1 U5036 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4515) );
  AOI22_X1 U5037 ( .A1(n4692), .A2(n4529), .B1(n4515), .B2(n4690), .ZN(U3485)
         );
  NOR2_X1 U5038 ( .A1(n4516), .A2(n2101), .ZN(n4518) );
  AOI211_X1 U5039 ( .C1(n4520), .C2(n4519), .A(n4518), .B(n4517), .ZN(n4532)
         );
  INV_X1 U5040 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4613) );
  AOI22_X1 U5041 ( .A1(n4692), .A2(n4532), .B1(n4613), .B2(n4690), .ZN(U3489)
         );
  AOI22_X1 U5042 ( .A1(n4533), .A2(n4521), .B1(n2990), .B2(n4530), .ZN(U3519)
         );
  INV_X1 U5043 ( .A(REG1_REG_3__SCAN_IN), .ZN(n4522) );
  AOI22_X1 U5044 ( .A1(n4533), .A2(n4523), .B1(n4522), .B2(n4530), .ZN(U3521)
         );
  AOI22_X1 U5045 ( .A1(n4533), .A2(n4524), .B1(n2080), .B2(n4530), .ZN(U3522)
         );
  AOI22_X1 U5046 ( .A1(n4533), .A2(n4526), .B1(n4525), .B2(n4530), .ZN(U3523)
         );
  AOI22_X1 U5047 ( .A1(n4533), .A2(n4527), .B1(n4598), .B2(n4530), .ZN(U3525)
         );
  AOI22_X1 U5048 ( .A1(n4533), .A2(n4529), .B1(n4528), .B2(n4530), .ZN(U3527)
         );
  AOI22_X1 U5049 ( .A1(n4533), .A2(n4532), .B1(n4531), .B2(n4530), .ZN(U3529)
         );
  OAI22_X1 U5050 ( .A1(n4536), .A2(keyinput2), .B1(n4535), .B2(keyinput35), 
        .ZN(n4534) );
  AOI221_X1 U5051 ( .B1(n4536), .B2(keyinput2), .C1(keyinput35), .C2(n4535), 
        .A(n4534), .ZN(n4548) );
  OAI22_X1 U5052 ( .A1(n4539), .A2(keyinput61), .B1(n4538), .B2(keyinput33), 
        .ZN(n4537) );
  AOI221_X1 U5053 ( .B1(n4539), .B2(keyinput61), .C1(keyinput33), .C2(n4538), 
        .A(n4537), .ZN(n4547) );
  OAI22_X1 U5054 ( .A1(n4541), .A2(keyinput25), .B1(n2147), .B2(keyinput18), 
        .ZN(n4540) );
  AOI221_X1 U5055 ( .B1(n4541), .B2(keyinput25), .C1(keyinput18), .C2(n2147), 
        .A(n4540), .ZN(n4546) );
  OAI22_X1 U5056 ( .A1(n4544), .A2(keyinput47), .B1(n4543), .B2(keyinput8), 
        .ZN(n4542) );
  AOI221_X1 U5057 ( .B1(n4544), .B2(keyinput47), .C1(keyinput8), .C2(n4543), 
        .A(n4542), .ZN(n4545) );
  NAND4_X1 U5058 ( .A1(n4548), .A2(n4547), .A3(n4546), .A4(n4545), .ZN(n4689)
         );
  OAI22_X1 U5059 ( .A1(n4551), .A2(keyinput10), .B1(n4550), .B2(keyinput38), 
        .ZN(n4549) );
  AOI221_X1 U5060 ( .B1(n4551), .B2(keyinput10), .C1(keyinput38), .C2(n4550), 
        .A(n4549), .ZN(n4564) );
  OAI22_X1 U5061 ( .A1(n4554), .A2(keyinput62), .B1(n4553), .B2(keyinput59), 
        .ZN(n4552) );
  AOI221_X1 U5062 ( .B1(n4554), .B2(keyinput62), .C1(keyinput59), .C2(n4553), 
        .A(n4552), .ZN(n4563) );
  INV_X1 U5063 ( .A(REG1_REG_29__SCAN_IN), .ZN(n4557) );
  INV_X1 U5064 ( .A(keyinput32), .ZN(n4556) );
  OAI22_X1 U5065 ( .A1(n4557), .A2(keyinput54), .B1(n4556), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4555) );
  AOI221_X1 U5066 ( .B1(n4557), .B2(keyinput54), .C1(DATAO_REG_30__SCAN_IN), 
        .C2(n4556), .A(n4555), .ZN(n4562) );
  INV_X1 U5067 ( .A(keyinput16), .ZN(n4560) );
  INV_X1 U5068 ( .A(keyinput19), .ZN(n4559) );
  OAI22_X1 U5069 ( .A1(n4560), .A2(DATAO_REG_25__SCAN_IN), .B1(n4559), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4558) );
  AOI221_X1 U5070 ( .B1(n4560), .B2(DATAO_REG_25__SCAN_IN), .C1(
        DATAO_REG_27__SCAN_IN), .C2(n4559), .A(n4558), .ZN(n4561) );
  NAND4_X1 U5071 ( .A1(n4564), .A2(n4563), .A3(n4562), .A4(n4561), .ZN(n4688)
         );
  INV_X1 U5072 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n4566) );
  NAND2_X1 U5073 ( .A1(U3149), .A2(keyinput6), .ZN(n4565) );
  OAI221_X1 U5074 ( .B1(n4566), .B2(keyinput9), .C1(U3149), .C2(keyinput6), 
        .A(n4565), .ZN(n4578) );
  INV_X1 U5075 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4569) );
  INV_X1 U5076 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4568) );
  AOI22_X1 U5077 ( .A1(n4569), .A2(keyinput3), .B1(n4568), .B2(keyinput30), 
        .ZN(n4567) );
  OAI221_X1 U5078 ( .B1(n4569), .B2(keyinput3), .C1(n4568), .C2(keyinput30), 
        .A(n4567), .ZN(n4577) );
  INV_X1 U5079 ( .A(keyinput50), .ZN(n4572) );
  INV_X1 U5080 ( .A(keyinput48), .ZN(n4571) );
  AOI22_X1 U5081 ( .A1(n4572), .A2(DATAO_REG_6__SCAN_IN), .B1(
        DATAO_REG_3__SCAN_IN), .B2(n4571), .ZN(n4570) );
  OAI221_X1 U5082 ( .B1(n4572), .B2(DATAO_REG_6__SCAN_IN), .C1(n4571), .C2(
        DATAO_REG_3__SCAN_IN), .A(n4570), .ZN(n4576) );
  INV_X1 U5083 ( .A(keyinput41), .ZN(n4574) );
  AOI22_X1 U5084 ( .A1(n2809), .A2(keyinput23), .B1(DATAO_REG_11__SCAN_IN), 
        .B2(n4574), .ZN(n4573) );
  OAI221_X1 U5085 ( .B1(n2809), .B2(keyinput23), .C1(n4574), .C2(
        DATAO_REG_11__SCAN_IN), .A(n4573), .ZN(n4575) );
  NOR4_X1 U5086 ( .A1(n4578), .A2(n4577), .A3(n4576), .A4(n4575), .ZN(n4625)
         );
  INV_X1 U5087 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4580) );
  INV_X1 U5088 ( .A(keyinput56), .ZN(n4626) );
  AOI22_X1 U5089 ( .A1(n4580), .A2(keyinput55), .B1(ADDR_REG_8__SCAN_IN), .B2(
        n4626), .ZN(n4579) );
  OAI221_X1 U5090 ( .B1(n4580), .B2(keyinput55), .C1(n4626), .C2(
        ADDR_REG_8__SCAN_IN), .A(n4579), .ZN(n4593) );
  INV_X1 U5091 ( .A(DATAI_30_), .ZN(n4582) );
  AOI22_X1 U5092 ( .A1(n4583), .A2(keyinput11), .B1(keyinput46), .B2(n4582), 
        .ZN(n4581) );
  OAI221_X1 U5093 ( .B1(n4583), .B2(keyinput11), .C1(n4582), .C2(keyinput46), 
        .A(n4581), .ZN(n4592) );
  INV_X1 U5094 ( .A(REG2_REG_10__SCAN_IN), .ZN(n4586) );
  INV_X1 U5095 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n4585) );
  AOI22_X1 U5096 ( .A1(n4586), .A2(keyinput4), .B1(keyinput21), .B2(n4585), 
        .ZN(n4584) );
  OAI221_X1 U5097 ( .B1(n4586), .B2(keyinput4), .C1(n4585), .C2(keyinput21), 
        .A(n4584), .ZN(n4591) );
  INV_X1 U5098 ( .A(keyinput29), .ZN(n4587) );
  XOR2_X1 U5099 ( .A(ADDR_REG_1__SCAN_IN), .B(n4587), .Z(n4589) );
  XNOR2_X1 U5100 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput63), .ZN(n4588) );
  NAND2_X1 U5101 ( .A1(n4589), .A2(n4588), .ZN(n4590) );
  NOR4_X1 U5102 ( .A1(n4593), .A2(n4592), .A3(n4591), .A4(n4590), .ZN(n4624)
         );
  INV_X1 U5103 ( .A(keyinput5), .ZN(n4595) );
  AOI22_X1 U5104 ( .A1(n4596), .A2(keyinput22), .B1(ADDR_REG_17__SCAN_IN), 
        .B2(n4595), .ZN(n4594) );
  OAI221_X1 U5105 ( .B1(n4596), .B2(keyinput22), .C1(n4595), .C2(
        ADDR_REG_17__SCAN_IN), .A(n4594), .ZN(n4608) );
  AOI22_X1 U5106 ( .A1(n4598), .A2(keyinput0), .B1(keyinput31), .B2(n2990), 
        .ZN(n4597) );
  OAI221_X1 U5107 ( .B1(n4598), .B2(keyinput0), .C1(n2990), .C2(keyinput31), 
        .A(n4597), .ZN(n4607) );
  AOI22_X1 U5108 ( .A1(n4601), .A2(keyinput45), .B1(n4600), .B2(keyinput57), 
        .ZN(n4599) );
  OAI221_X1 U5109 ( .B1(n4601), .B2(keyinput45), .C1(n4600), .C2(keyinput57), 
        .A(n4599), .ZN(n4606) );
  INV_X1 U5110 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4603) );
  AOI22_X1 U5111 ( .A1(n4604), .A2(keyinput44), .B1(n4603), .B2(keyinput42), 
        .ZN(n4602) );
  OAI221_X1 U5112 ( .B1(n4604), .B2(keyinput44), .C1(n4603), .C2(keyinput42), 
        .A(n4602), .ZN(n4605) );
  NOR4_X1 U5113 ( .A1(n4608), .A2(n4607), .A3(n4606), .A4(n4605), .ZN(n4623)
         );
  INV_X1 U5114 ( .A(keyinput43), .ZN(n4610) );
  AOI22_X1 U5115 ( .A1(n4611), .A2(keyinput37), .B1(DATAO_REG_20__SCAN_IN), 
        .B2(n4610), .ZN(n4609) );
  OAI221_X1 U5116 ( .B1(n4611), .B2(keyinput37), .C1(n4610), .C2(
        DATAO_REG_20__SCAN_IN), .A(n4609), .ZN(n4621) );
  AOI22_X1 U5117 ( .A1(n4614), .A2(keyinput34), .B1(n4613), .B2(keyinput17), 
        .ZN(n4612) );
  OAI221_X1 U5118 ( .B1(n4614), .B2(keyinput34), .C1(n4613), .C2(keyinput17), 
        .A(n4612), .ZN(n4620) );
  XNOR2_X1 U5119 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput36), .ZN(n4618) );
  XNOR2_X1 U5120 ( .A(DATAI_9_), .B(keyinput39), .ZN(n4617) );
  XNOR2_X1 U5121 ( .A(IR_REG_7__SCAN_IN), .B(keyinput58), .ZN(n4616) );
  XNOR2_X1 U5122 ( .A(keyinput13), .B(REG0_REG_2__SCAN_IN), .ZN(n4615) );
  NAND4_X1 U5123 ( .A1(n4618), .A2(n4617), .A3(n4616), .A4(n4615), .ZN(n4619)
         );
  NOR3_X1 U5124 ( .A1(n4621), .A2(n4620), .A3(n4619), .ZN(n4622) );
  NAND4_X1 U5125 ( .A1(n4625), .A2(n4624), .A3(n4623), .A4(n4622), .ZN(n4687)
         );
  NAND2_X1 U5126 ( .A1(keyinput3), .A2(keyinput1), .ZN(n4631) );
  NAND4_X1 U5127 ( .A1(keyinput55), .A2(keyinput29), .A3(keyinput4), .A4(n4626), .ZN(n4630) );
  NOR3_X1 U5128 ( .A1(keyinput30), .A2(keyinput50), .A3(keyinput41), .ZN(n4628) );
  NOR3_X1 U5129 ( .A1(keyinput11), .A2(keyinput46), .A3(keyinput63), .ZN(n4627) );
  NAND4_X1 U5130 ( .A1(keyinput48), .A2(n4628), .A3(keyinput23), .A4(n4627), 
        .ZN(n4629) );
  NOR4_X1 U5131 ( .A1(keyinput6), .A2(n4631), .A3(n4630), .A4(n4629), .ZN(
        n4656) );
  NOR2_X1 U5132 ( .A1(keyinput21), .A2(keyinput22), .ZN(n4632) );
  NAND3_X1 U5133 ( .A1(keyinput5), .A2(keyinput0), .A3(n4632), .ZN(n4654) );
  NOR2_X1 U5134 ( .A1(keyinput31), .A2(keyinput44), .ZN(n4637) );
  NAND2_X1 U5135 ( .A1(keyinput36), .A2(keyinput34), .ZN(n4635) );
  NOR2_X1 U5136 ( .A1(keyinput17), .A2(keyinput43), .ZN(n4633) );
  NAND3_X1 U5137 ( .A1(keyinput58), .A2(keyinput39), .A3(n4633), .ZN(n4634) );
  NOR4_X1 U5138 ( .A1(keyinput42), .A2(keyinput13), .A3(n4635), .A4(n4634), 
        .ZN(n4636) );
  NAND4_X1 U5139 ( .A1(keyinput45), .A2(keyinput57), .A3(n4637), .A4(n4636), 
        .ZN(n4653) );
  NOR2_X1 U5140 ( .A1(keyinput37), .A2(keyinput62), .ZN(n4644) );
  NAND2_X1 U5141 ( .A1(keyinput19), .A2(keyinput54), .ZN(n4642) );
  NOR3_X1 U5142 ( .A1(keyinput32), .A2(keyinput61), .A3(keyinput33), .ZN(n4640) );
  INV_X1 U5143 ( .A(keyinput8), .ZN(n4638) );
  NOR3_X1 U5144 ( .A1(keyinput35), .A2(keyinput25), .A3(n4638), .ZN(n4639) );
  NAND4_X1 U5145 ( .A1(keyinput2), .A2(n4640), .A3(keyinput47), .A4(n4639), 
        .ZN(n4641) );
  NOR4_X1 U5146 ( .A1(keyinput38), .A2(keyinput16), .A3(n4642), .A4(n4641), 
        .ZN(n4643) );
  NAND4_X1 U5147 ( .A1(keyinput10), .A2(keyinput59), .A3(n4644), .A4(n4643), 
        .ZN(n4652) );
  NOR3_X1 U5148 ( .A1(keyinput15), .A2(keyinput14), .A3(keyinput51), .ZN(n4650) );
  NAND2_X1 U5149 ( .A1(keyinput28), .A2(keyinput60), .ZN(n4645) );
  NOR3_X1 U5150 ( .A1(keyinput40), .A2(keyinput24), .A3(n4645), .ZN(n4649) );
  NAND4_X1 U5151 ( .A1(keyinput18), .A2(keyinput26), .A3(keyinput27), .A4(
        keyinput7), .ZN(n4647) );
  NAND2_X1 U5152 ( .A1(keyinput12), .A2(keyinput49), .ZN(n4646) );
  NOR4_X1 U5153 ( .A1(keyinput53), .A2(keyinput20), .A3(n4647), .A4(n4646), 
        .ZN(n4648) );
  NAND4_X1 U5154 ( .A1(keyinput52), .A2(n4650), .A3(n4649), .A4(n4648), .ZN(
        n4651) );
  NOR4_X1 U5155 ( .A1(n4654), .A2(n4653), .A3(n4652), .A4(n4651), .ZN(n4655)
         );
  AOI21_X1 U5156 ( .B1(n4656), .B2(n4655), .A(keyinput9), .ZN(n4685) );
  INV_X1 U5157 ( .A(DATAI_22_), .ZN(n4658) );
  AOI22_X1 U5158 ( .A1(n4659), .A2(keyinput40), .B1(keyinput28), .B2(n4658), 
        .ZN(n4657) );
  OAI221_X1 U5159 ( .B1(n4659), .B2(keyinput40), .C1(n4658), .C2(keyinput28), 
        .A(n4657), .ZN(n4669) );
  AOI22_X1 U5160 ( .A1(n2385), .A2(keyinput24), .B1(n2436), .B2(keyinput20), 
        .ZN(n4660) );
  OAI221_X1 U5161 ( .B1(n2385), .B2(keyinput24), .C1(n2436), .C2(keyinput20), 
        .A(n4660), .ZN(n4668) );
  AOI22_X1 U5162 ( .A1(n2069), .A2(keyinput1), .B1(keyinput53), .B2(n4662), 
        .ZN(n4661) );
  OAI221_X1 U5163 ( .B1(n2069), .B2(keyinput1), .C1(n4662), .C2(keyinput53), 
        .A(n4661), .ZN(n4667) );
  XOR2_X1 U5164 ( .A(n4663), .B(keyinput49), .Z(n4665) );
  XNOR2_X1 U5165 ( .A(DATAI_4_), .B(keyinput12), .ZN(n4664) );
  NAND2_X1 U5166 ( .A1(n4665), .A2(n4664), .ZN(n4666) );
  NOR4_X1 U5167 ( .A1(n4669), .A2(n4668), .A3(n4667), .A4(n4666), .ZN(n4684)
         );
  XOR2_X1 U5168 ( .A(IR_REG_21__SCAN_IN), .B(keyinput60), .Z(n4675) );
  XOR2_X1 U5169 ( .A(REG3_REG_18__SCAN_IN), .B(keyinput51), .Z(n4674) );
  XNOR2_X1 U5170 ( .A(n4670), .B(keyinput14), .ZN(n4673) );
  XNOR2_X1 U5171 ( .A(keyinput15), .B(n4671), .ZN(n4672) );
  NOR4_X1 U5172 ( .A1(n4675), .A2(n4674), .A3(n4673), .A4(n4672), .ZN(n4679)
         );
  XOR2_X1 U5173 ( .A(n2145), .B(keyinput26), .Z(n4678) );
  XNOR2_X1 U5174 ( .A(IR_REG_8__SCAN_IN), .B(keyinput7), .ZN(n4677) );
  XNOR2_X1 U5175 ( .A(IR_REG_13__SCAN_IN), .B(keyinput27), .ZN(n4676) );
  NAND4_X1 U5176 ( .A1(n4679), .A2(n4678), .A3(n4677), .A4(n4676), .ZN(n4682)
         );
  XNOR2_X1 U5177 ( .A(n4680), .B(keyinput52), .ZN(n4681) );
  NOR2_X1 U5178 ( .A1(n4682), .A2(n4681), .ZN(n4683) );
  OAI211_X1 U5179 ( .C1(ADDR_REG_3__SCAN_IN), .C2(n4685), .A(n4684), .B(n4683), 
        .ZN(n4686) );
  NOR4_X1 U5180 ( .A1(n4689), .A2(n4688), .A3(n4687), .A4(n4686), .ZN(n4694)
         );
  AOI22_X1 U5181 ( .A1(n4692), .A2(n4691), .B1(REG0_REG_0__SCAN_IN), .B2(n4690), .ZN(n4693) );
  XNOR2_X1 U5182 ( .A(n4694), .B(n4693), .ZN(U3467) );
endmodule

