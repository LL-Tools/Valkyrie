

module b22_C_gen_AntiSAT_k_256_3 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, 
        keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, 
        keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, 
        keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, 
        keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, 
        keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, 
        keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, 
        keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, 
        keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104, 
        keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108, 
        keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112, 
        keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116, 
        keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120, 
        keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124, 
        keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, 
        keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, 
        keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, 
        keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, 
        keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, 
        keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, 
        keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, 
        keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65,
         keyinput_f66, keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70,
         keyinput_f71, keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75,
         keyinput_f76, keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80,
         keyinput_f81, keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85,
         keyinput_f86, keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90,
         keyinput_f91, keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95,
         keyinput_f96, keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100,
         keyinput_f101, keyinput_f102, keyinput_f103, keyinput_f104,
         keyinput_f105, keyinput_f106, keyinput_f107, keyinput_f108,
         keyinput_f109, keyinput_f110, keyinput_f111, keyinput_f112,
         keyinput_f113, keyinput_f114, keyinput_f115, keyinput_f116,
         keyinput_f117, keyinput_f118, keyinput_f119, keyinput_f120,
         keyinput_f121, keyinput_f122, keyinput_f123, keyinput_f124,
         keyinput_f125, keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66,
         keyinput_g67, keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71,
         keyinput_g72, keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76,
         keyinput_g77, keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81,
         keyinput_g82, keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86,
         keyinput_g87, keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91,
         keyinput_g92, keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96,
         keyinput_g97, keyinput_g98, keyinput_g99, keyinput_g100,
         keyinput_g101, keyinput_g102, keyinput_g103, keyinput_g104,
         keyinput_g105, keyinput_g106, keyinput_g107, keyinput_g108,
         keyinput_g109, keyinput_g110, keyinput_g111, keyinput_g112,
         keyinput_g113, keyinput_g114, keyinput_g115, keyinput_g116,
         keyinput_g117, keyinput_g118, keyinput_g119, keyinput_g120,
         keyinput_g121, keyinput_g122, keyinput_g123, keyinput_g124,
         keyinput_g125, keyinput_g126, keyinput_g127;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164,
         n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         n10357, n10358, n10359, n10360, n10361, n10362, n10363, n10364,
         n10365, n10366, n10367, n10368, n10369, n10370, n10371, n10372,
         n10373, n10374, n10375, n10376, n10377, n10378, n10379, n10380,
         n10381, n10382, n10383, n10384, n10385, n10386, n10387, n10388,
         n10389, n10390, n10391, n10392, n10393, n10394, n10395, n10396,
         n10397, n10398, n10399, n10400, n10401, n10402, n10403, n10404,
         n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
         n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
         n10421, n10422, n10423, n10424, n10425, n10426, n10427, n10428,
         n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436,
         n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444,
         n10445, n10446, n10447, n10448, n10449, n10450, n10451, n10452,
         n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
         n10461, n10462, n10463, n10464, n10465, n10466, n10467, n10468,
         n10469, n10470, n10471, n10472, n10473, n10474, n10475, n10476,
         n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
         n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492,
         n10493, n10494, n10495, n10496, n10497, n10498, n10499, n10500,
         n10501, n10502, n10503, n10504, n10505, n10506, n10507, n10508,
         n10509, n10510, n10511, n10512, n10513, n10514, n10515, n10516,
         n10517, n10518, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10529, n10530, n10531, n10532,
         n10533, n10534, n10535, n10536, n10537, n10538, n10539, n10540,
         n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
         n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
         n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
         n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572,
         n10573, n10574, n10575, n10576, n10577, n10578, n10579, n10580,
         n10581, n10582, n10583, n10584, n10585, n10586, n10587, n10588,
         n10589, n10590, n10591, n10592, n10593, n10594, n10595, n10596,
         n10597, n10598, n10599, n10600, n10601, n10602, n10603, n10604,
         n10605, n10606, n10607, n10608, n10609, n10610, n10611, n10612,
         n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
         n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644,
         n10645, n10646, n10647, n10648, n10649, n10650, n10651, n10652,
         n10653, n10654, n10655, n10656, n10657, n10658, n10659, n10660,
         n10661, n10662, n10663, n10664, n10665, n10666, n10667, n10668,
         n10669, n10670, n10671, n10672, n10673, n10674, n10675, n10676,
         n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
         n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
         n10693, n10694, n10695, n10696, n10697, n10698, n10699, n10700,
         n10701, n10702, n10703, n10704, n10705, n10706, n10707, n10708,
         n10709, n10710, n10711, n10712, n10713, n10714, n10715, n10716,
         n10717, n10718, n10719, n10720, n10721, n10722, n10723, n10724,
         n10725, n10726, n10727, n10728, n10729, n10730, n10731, n10732,
         n10733, n10734, n10735, n10736, n10737, n10738, n10739, n10740,
         n10741, n10742, n10743, n10744, n10745, n10746, n10747, n10748,
         n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756,
         n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
         n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10777, n10778, n10779, n10780,
         n10781, n10782, n10783, n10784, n10785, n10786, n10787, n10788,
         n10789, n10790, n10791, n10792, n10793, n10794, n10795, n10796,
         n10797, n10798, n10799, n10800, n10801, n10802, n10803, n10804,
         n10805, n10806, n10807, n10808, n10809, n10810, n10811, n10812,
         n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
         n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844,
         n10845, n10846, n10847, n10848, n10849, n10850, n10851, n10852,
         n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
         n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868,
         n10869, n10870, n10871, n10872, n10873, n10874, n10875, n10876,
         n10877, n10878, n10879, n10880, n10881, n10882, n10883, n10884,
         n10885, n10886, n10887, n10888, n10889, n10890, n10891, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268,
         n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
         n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284,
         n12285, n12286, n12287, n12288, n12289, n12290, n12291, n12292,
         n12293, n12294, n12295, n12296, n12297, n12298, n12299, n12300,
         n12301, n12302, n12303, n12304, n12305, n12306, n12307, n12308,
         n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316,
         n12317, n12318, n12319, n12320, n12321, n12322, n12323, n12324,
         n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
         n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340,
         n12341, n12342, n12343, n12344, n12345, n12346, n12347, n12348,
         n12349, n12350, n12351, n12352, n12353, n12354, n12355, n12356,
         n12357, n12358, n12359, n12360, n12361, n12362, n12363, n12364,
         n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
         n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380,
         n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
         n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396,
         n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
         n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412,
         n12413, n12414, n12415, n12416, n12417, n12418, n12419, n12420,
         n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
         n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436,
         n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
         n12445, n12446, n12447, n12448, n12449, n12450, n12451, n12452,
         n12453, n12454, n12455, n12456, n12457, n12458, n12459, n12460,
         n12461, n12462, n12463, n12464, n12465, n12466, n12467, n12468,
         n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
         n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484,
         n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
         n12493, n12494, n12495, n12496, n12497, n12498, n12499, n12500,
         n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
         n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516,
         n12517, n12518, n12519, n12520, n12521, n12522, n12523, n12524,
         n12525, n12526, n12527, n12528, n12529, n12530, n12531, n12532,
         n12533, n12534, n12535, n12536, n12537, n12538, n12539, n12540,
         n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
         n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556,
         n12557, n12558, n12559, n12560, n12561, n12562, n12563, n12564,
         n12565, n12566, n12567, n12568, n12569, n12570, n12571, n12572,
         n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
         n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
         n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596,
         n12597, n12598, n12599, n12600, n12601, n12602, n12603, n12604,
         n12605, n12606, n12607, n12608, n12609, n12610, n12611, n12612,
         n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
         n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
         n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636,
         n12637, n12638, n12639, n12640, n12641, n12642, n12643, n12644,
         n12645, n12646, n12647, n12648, n12649, n12650, n12651, n12652,
         n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
         n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668,
         n12669, n12670, n12671, n12672, n12673, n12674, n12675, n12676,
         n12677, n12678, n12679, n12680, n12681, n12682, n12683, n12684,
         n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
         n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700,
         n12701, n12702, n12703, n12704, n12705, n12706, n12707, n12708,
         n12709, n12710, n12711, n12712, n12713, n12714, n12715, n12716,
         n12717, n12718, n12719, n12720, n12721, n12722, n12723, n12724,
         n12725, n12726, n12727, n12728, n12729, n12730, n12731, n12732,
         n12733, n12734, n12735, n12736, n12737, n12738, n12739, n12740,
         n12741, n12742, n12743, n12744, n12745, n12746, n12747, n12748,
         n12749, n12750, n12751, n12752, n12753, n12754, n12755, n12756,
         n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764,
         n12765, n12766, n12767, n12768, n12769, n12770, n12771, n12772,
         n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
         n12781, n12782, n12783, n12784, n12785, n12786, n12787, n12788,
         n12789, n12790, n12791, n12792, n12793, n12794, n12795, n12796,
         n12797, n12798, n12799, n12800, n12801, n12802, n12803, n12804,
         n12805, n12806, n12807, n12808, n12809, n12810, n12811, n12812,
         n12813, n12814, n12815, n12816, n12817, n12818, n12819, n12820,
         n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
         n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836,
         n12837, n12838, n12839, n12840, n12841, n12842, n12843, n12844,
         n12845, n12846, n12847, n12848, n12849, n12850, n12851, n12852,
         n12853, n12854, n12855, n12856, n12857, n12858, n12859, n12860,
         n12861, n12862, n12863, n12864, n12865, n12866, n12867, n12868,
         n12869, n12870, n12871, n12872, n12873, n12874, n12875, n12876,
         n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884,
         n12885, n12886, n12887, n12888, n12889, n12890, n12891, n12892,
         n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
         n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908,
         n12909, n12910, n12911, n12912, n12913, n12914, n12915, n12916,
         n12917, n12918, n12919, n12920, n12921, n12922, n12923, n12924,
         n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
         n12933, n12934, n12935, n12936, n12937, n12938, n12939, n12940,
         n12941, n12942, n12943, n12944, n12945, n12946, n12947, n12948,
         n12949, n12950, n12951, n12952, n12953, n12954, n12955, n12956,
         n12957, n12958, n12959, n12960, n12961, n12962, n12963, n12964,
         n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
         n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980,
         n12981, n12982, n12983, n12984, n12985, n12986, n12987, n12988,
         n12989, n12990, n12991, n12992, n12993, n12994, n12995, n12996,
         n12997, n12998, n12999, n13000, n13001, n13002, n13003, n13004,
         n13005, n13006, n13007, n13008, n13009, n13010, n13011, n13012,
         n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020,
         n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
         n13029, n13030, n13031, n13032, n13033, n13034, n13035, n13036,
         n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
         n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052,
         n13053, n13054, n13055, n13056, n13057, n13058, n13059, n13060,
         n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
         n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076,
         n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
         n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092,
         n13093, n13094, n13095, n13096, n13097, n13098, n13099, n13100,
         n13101, n13102, n13103, n13104, n13105, n13106, n13107, n13108,
         n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
         n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124,
         n13125, n13126, n13127, n13128, n13129, n13130, n13131, n13132,
         n13133, n13134, n13135, n13136, n13137, n13138, n13139, n13140,
         n13141, n13142, n13143, n13144, n13145, n13146, n13147, n13148,
         n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
         n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164,
         n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172,
         n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
         n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
         n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196,
         n13197, n13198, n13199, n13200, n13201, n13202, n13203, n13204,
         n13205, n13206, n13207, n13208, n13209, n13210, n13211, n13212,
         n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220,
         n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
         n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236,
         n13237, n13238, n13239, n13240, n13241, n13242, n13243, n13244,
         n13245, n13246, n13247, n13248, n13249, n13250, n13251, n13252,
         n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
         n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268,
         n13269, n13270, n13271, n13272, n13273, n13274, n13275, n13276,
         n13277, n13278, n13279, n13280, n13281, n13282, n13283, n13284,
         n13285, n13286, n13287, n13288, n13289, n13290, n13291, n13292,
         n13293, n13294, n13295, n13296, n13297, n13298, n13299, n13300,
         n13301, n13302, n13303, n13304, n13305, n13306, n13307, n13308,
         n13309, n13310, n13311, n13312, n13313, n13314, n13315, n13316,
         n13317, n13318, n13319, n13320, n13321, n13322, n13323, n13324,
         n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
         n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340,
         n13341, n13342, n13343, n13344, n13345, n13346, n13347, n13348,
         n13349, n13350, n13351, n13352, n13353, n13354, n13355, n13356,
         n13357, n13358, n13359, n13360, n13361, n13362, n13363, n13364,
         n13365, n13366, n13367, n13368, n13369, n13370, n13371, n13372,
         n13373, n13374, n13375, n13376, n13377, n13378, n13379, n13380,
         n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388,
         n13389, n13390, n13391, n13392, n13393, n13394, n13395, n13396,
         n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
         n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
         n13413, n13414, n13415, n13416, n13417, n13418, n13419, n13420,
         n13421, n13422, n13423, n13424, n13425, n13426, n13427, n13428,
         n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
         n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444,
         n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
         n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460,
         n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
         n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476,
         n13477, n13478, n13479, n13480, n13481, n13482, n13483, n13484,
         n13485, n13486, n13487, n13488, n13489, n13490, n13491, n13492,
         n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
         n13501, n13502, n13503, n13504, n13505, n13506, n13507, n13508,
         n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
         n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
         n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
         n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540,
         n13541, n13542, n13543, n13544, n13545, n13546, n13547, n13548,
         n13549, n13550, n13551, n13552, n13553, n13554, n13555, n13556,
         n13557, n13558, n13559, n13560, n13561, n13562, n13563, n13564,
         n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
         n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
         n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588,
         n13589, n13590, n13591, n13592, n13593, n13594, n13595, n13596,
         n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
         n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612,
         n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
         n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628,
         n13629, n13630, n13631, n13632, n13633, n13634, n13635, n13636,
         n13637, n13638, n13639, n13640, n13641, n13642, n13643, n13644,
         n13645, n13646, n13647, n13648, n13649, n13650, n13651, n13652,
         n13653, n13654, n13655, n13656, n13657, n13658, n13659, n13660,
         n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
         n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
         n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684,
         n13685, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624;

  INV_X1 U7414 ( .A(n10727), .ZN(n13729) );
  INV_X2 U7415 ( .A(n9341), .ZN(n9616) );
  INV_X1 U7416 ( .A(n9523), .ZN(n7251) );
  INV_X1 U7417 ( .A(n15300), .ZN(n10725) );
  CLKBUF_X2 U7420 ( .A(n8764), .Z(n8752) );
  AND4_X1 U7421 ( .A1(n8416), .A2(n8415), .A3(n8414), .A4(n8413), .ZN(n8952)
         );
  CLKBUF_X2 U7422 ( .A(n9420), .Z(n6666) );
  NOR2_X2 U7423 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n8447) );
  XNOR2_X1 U7424 ( .A(n7168), .B(n6849), .ZN(n10160) );
  NAND2_X2 U7425 ( .A1(n7761), .A2(n12947), .ZN(n8361) );
  NAND2_X1 U7426 ( .A1(n8382), .A2(n13679), .ZN(n13685) );
  AND2_X1 U7427 ( .A1(n10135), .A2(n10030), .ZN(n7377) );
  INV_X1 U7428 ( .A(n10005), .ZN(n9908) );
  NOR4_X1 U7429 ( .A1(n12875), .A2(n12861), .A3(n13114), .A4(n12860), .ZN(
        n12862) );
  INV_X1 U7430 ( .A(n9015), .ZN(n9026) );
  XNOR2_X1 U7431 ( .A(n7728), .B(n10153), .ZN(n11045) );
  INV_X1 U7432 ( .A(n10727), .ZN(n13734) );
  NOR2_X1 U7433 ( .A1(n15480), .A2(n6811), .ZN(n7780) );
  AND2_X1 U7434 ( .A1(n8916), .A2(n13422), .ZN(n13435) );
  INV_X1 U7435 ( .A(n8361), .ZN(n8636) );
  OR2_X1 U7436 ( .A1(n8324), .A2(n10287), .ZN(n8325) );
  CLKBUF_X2 U7437 ( .A(n9599), .Z(n9924) );
  OR2_X1 U7438 ( .A1(n13699), .A2(n14981), .ZN(n14092) );
  AND2_X1 U7439 ( .A1(n11139), .A2(n11130), .ZN(n11024) );
  INV_X1 U7440 ( .A(n10886), .ZN(n13057) );
  INV_X2 U7441 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n7593) );
  NAND2_X1 U7442 ( .A1(n15060), .A2(n12412), .ZN(n15063) );
  INV_X1 U7443 ( .A(n15131), .ZN(n11582) );
  INV_X1 U7444 ( .A(n12530), .ZN(n11632) );
  OAI211_X1 U7445 ( .C1(n8663), .C2(n10158), .A(n7120), .B(n7119), .ZN(n10719)
         );
  INV_X1 U7446 ( .A(n12390), .ZN(n12398) );
  NAND2_X1 U7447 ( .A1(n8684), .A2(n8683), .ZN(n13494) );
  NAND2_X1 U7448 ( .A1(n8834), .A2(n8835), .ZN(n11940) );
  NAND2_X1 U7449 ( .A1(n8378), .A2(n8377), .ZN(n13679) );
  NAND2_X1 U7450 ( .A1(n8380), .A2(n7751), .ZN(n12947) );
  INV_X1 U7451 ( .A(n13957), .ZN(n14122) );
  NAND2_X1 U7452 ( .A1(n9629), .A2(n9628), .ZN(n14110) );
  NAND2_X1 U7453 ( .A1(n9685), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9081) );
  INV_X2 U7454 ( .A(n12475), .ZN(n14483) );
  NAND2_X2 U7455 ( .A1(n14872), .A2(n10247), .ZN(n12738) );
  AND2_X1 U7456 ( .A1(n7117), .A2(n7118), .ZN(n7115) );
  XNOR2_X1 U7457 ( .A(n7671), .B(n7670), .ZN(n10768) );
  INV_X1 U7458 ( .A(n9722), .ZN(n13890) );
  AOI21_X1 U7459 ( .B1(n12913), .B2(n14618), .A(n12912), .ZN(n14736) );
  INV_X2 U7460 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n9093) );
  NOR2_X2 U7461 ( .A1(n10568), .A2(n7714), .ZN(n7718) );
  AND2_X2 U7462 ( .A1(n6700), .A2(n9109), .ZN(n9233) );
  AND2_X1 U7463 ( .A1(n11568), .A2(n15341), .ZN(n11642) );
  NOR2_X2 U7464 ( .A1(n11170), .A2(n11272), .ZN(n11568) );
  AOI21_X2 U7465 ( .B1(n14016), .B2(n14015), .A(n7272), .ZN(n13999) );
  NAND4_X4 U7466 ( .A1(n10837), .A2(n10836), .A3(n10835), .A4(n10834), .ZN(
        n14376) );
  NAND2_X2 U7467 ( .A1(n7925), .A2(n15615), .ZN(n14896) );
  OAI21_X1 U7468 ( .B1(n14109), .B2(n15000), .A(n6714), .ZN(n14173) );
  XNOR2_X2 U7469 ( .A(n14375), .B(n11797), .ZN(n11479) );
  OAI222_X1 U7470 ( .A1(n14874), .A2(n14195), .B1(P1_U3086), .B2(n12951), .C1(
        n12950), .C2(n14876), .ZN(P1_U3326) );
  OAI21_X2 U7471 ( .B1(n9039), .B2(n8924), .A(n8922), .ZN(n8951) );
  AOI21_X2 U7472 ( .B1(n13423), .B2(n13422), .A(n13421), .ZN(n9039) );
  OAI22_X2 U7473 ( .A1(n13939), .A2(n13944), .B1(n13943), .B2(n9907), .ZN(
        n13924) );
  NOR4_X2 U7474 ( .A1(n8934), .A2(n8795), .A3(n8930), .A4(n8793), .ZN(n8794)
         );
  OAI21_X1 U7475 ( .B1(n10160), .B2(n10954), .A(n7708), .ZN(n10598) );
  AOI21_X2 U7476 ( .B1(n13283), .B2(n13197), .A(n13196), .ZN(n13263) );
  OAI22_X2 U7477 ( .A1(n9608), .A2(n7328), .B1(n7327), .B2(n12139), .ZN(n9626)
         );
  OAI21_X2 U7478 ( .B1(n9675), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9657) );
  OAI22_X2 U7479 ( .A1(n13235), .A2(n13236), .B1(n13173), .B2(n13302), .ZN(
        n13300) );
  AOI21_X2 U7480 ( .B1(n13195), .B2(n13171), .A(n13170), .ZN(n13235) );
  NOR2_X2 U7481 ( .A1(n15512), .A2(n15511), .ZN(n15510) );
  NOR2_X2 U7482 ( .A1(n7735), .A2(n13331), .ZN(n15512) );
  INV_X1 U7483 ( .A(n7761), .ZN(n7844) );
  XNOR2_X2 U7484 ( .A(n7753), .B(n7752), .ZN(n7761) );
  NOR2_X2 U7485 ( .A1(n9741), .A2(n6721), .ZN(n7641) );
  NOR2_X2 U7486 ( .A1(n14992), .A2(n14993), .ZN(n9741) );
  AND3_X4 U7487 ( .A1(n6725), .A2(n7052), .A3(n7051), .ZN(n15300) );
  XOR2_X2 U7488 ( .A(n7866), .B(P3_ADDR_REG_4__SCAN_IN), .Z(n6694) );
  NAND2_X2 U7489 ( .A1(n7864), .A2(n7865), .ZN(n7866) );
  NOR2_X2 U7490 ( .A1(n13367), .A2(n13366), .ZN(n13365) );
  NOR2_X2 U7491 ( .A1(n7737), .A2(n13349), .ZN(n13367) );
  XNOR2_X1 U7492 ( .A(n10945), .B(n7021), .ZN(n10942) );
  INV_X1 U7493 ( .A(n13886), .ZN(n7021) );
  AOI21_X2 U7494 ( .B1(P3_REG2_REG_14__SCAN_IN), .B2(n15519), .A(n15510), .ZN(
        n7736) );
  NAND2_X1 U7495 ( .A1(n9922), .A2(n9921), .ZN(n13910) );
  NAND2_X1 U7496 ( .A1(n8922), .A2(n8777), .ZN(n13216) );
  XNOR2_X1 U7497 ( .A(n9644), .B(n9643), .ZN(n14869) );
  AND2_X1 U7498 ( .A1(n9595), .A2(n9594), .ZN(n13957) );
  NAND2_X1 U7499 ( .A1(n9752), .A2(n9751), .ZN(n14014) );
  AOI21_X1 U7500 ( .B1(n6922), .B2(n6925), .A(n6921), .ZN(n13780) );
  XNOR2_X1 U7501 ( .A(n14126), .B(n13866), .ZN(n13971) );
  INV_X1 U7502 ( .A(n13975), .ZN(n14126) );
  NAND2_X1 U7503 ( .A1(n12749), .A2(n12748), .ZN(n14757) );
  NAND2_X1 U7504 ( .A1(n12774), .A2(n12773), .ZN(n14751) );
  CLKBUF_X1 U7505 ( .A(n14224), .Z(n14311) );
  AND2_X1 U7506 ( .A1(n9458), .A2(n9457), .ZN(n14072) );
  OR2_X1 U7507 ( .A1(n9810), .A2(n7424), .ZN(n7423) );
  INV_X2 U7508 ( .A(n12555), .ZN(n11797) );
  NAND2_X1 U7509 ( .A1(n11091), .A2(n15539), .ZN(n8817) );
  INV_X2 U7510 ( .A(n11755), .ZN(n11543) );
  INV_X1 U7511 ( .A(n11713), .ZN(n6816) );
  INV_X1 U7512 ( .A(n13888), .ZN(n9786) );
  CLKBUF_X3 U7513 ( .A(n11713), .Z(n12432) );
  OR2_X1 U7514 ( .A1(n8601), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8613) );
  CLKBUF_X1 U7515 ( .A(n8995), .Z(n10242) );
  CLKBUF_X2 U7516 ( .A(n8752), .Z(n8737) );
  INV_X2 U7517 ( .A(n10734), .ZN(n10697) );
  NAND2_X2 U7518 ( .A1(n10768), .A2(n11039), .ZN(n10706) );
  XNOR2_X1 U7519 ( .A(n9121), .B(n9142), .ZN(n9106) );
  INV_X1 U7520 ( .A(n11474), .ZN(n10691) );
  CLKBUF_X2 U7522 ( .A(n12753), .Z(n12786) );
  INV_X1 U7523 ( .A(n9928), .ZN(n9097) );
  NAND2_X1 U7524 ( .A1(n9070), .A2(n9072), .ZN(n9131) );
  NAND2_X1 U7526 ( .A1(n6857), .A2(n6854), .ZN(n14194) );
  NAND2_X1 U7527 ( .A1(n6864), .A2(n6861), .ZN(n14872) );
  NAND2_X1 U7528 ( .A1(n7377), .A2(n10029), .ZN(n10489) );
  INV_X1 U7529 ( .A(n9181), .ZN(n10170) );
  AND2_X1 U7530 ( .A1(n8487), .A2(n8486), .ZN(n8500) );
  NAND2_X1 U7531 ( .A1(n10026), .A2(n10025), .ZN(n10495) );
  NAND2_X1 U7532 ( .A1(n8360), .A2(n8359), .ZN(n6670) );
  NAND2_X1 U7533 ( .A1(n7437), .A2(n7433), .ZN(n9970) );
  NOR2_X1 U7534 ( .A1(n9955), .A2(n7434), .ZN(n7433) );
  NAND2_X1 U7535 ( .A1(n9904), .A2(n7432), .ZN(n7437) );
  NAND2_X1 U7536 ( .A1(n12936), .A2(n12935), .ZN(n14507) );
  INV_X1 U7537 ( .A(n14497), .ZN(n14824) );
  NAND2_X1 U7538 ( .A1(n12473), .A2(n12472), .ZN(n14488) );
  OAI21_X1 U7539 ( .B1(n7534), .B2(n6907), .A(n6748), .ZN(n6906) );
  NAND2_X1 U7540 ( .A1(n12495), .A2(n12494), .ZN(n14497) );
  NAND2_X1 U7541 ( .A1(n14532), .A2(n12907), .ZN(n14521) );
  NAND2_X1 U7542 ( .A1(n14547), .A2(n7223), .ZN(n14532) );
  OAI211_X1 U7543 ( .C1(n9947), .C2(n9946), .A(n9945), .B(n9944), .ZN(n14186)
         );
  XNOR2_X1 U7544 ( .A(n14106), .B(n13862), .ZN(n9995) );
  NAND2_X1 U7545 ( .A1(n12518), .A2(n12517), .ZN(n13101) );
  XNOR2_X1 U7546 ( .A(n9920), .B(n9919), .ZN(n12885) );
  NAND2_X1 U7547 ( .A1(n9642), .A2(n9641), .ZN(n13923) );
  NAND2_X1 U7548 ( .A1(n7331), .A2(n9649), .ZN(n14106) );
  OR2_X1 U7549 ( .A1(n14110), .A2(n13769), .ZN(n9642) );
  AOI21_X1 U7550 ( .B1(n7293), .B2(n7291), .A(n7290), .ZN(n7289) );
  NAND2_X1 U7551 ( .A1(n14578), .A2(n12903), .ZN(n14563) );
  NAND2_X1 U7552 ( .A1(n9914), .A2(n9913), .ZN(n9943) );
  XNOR2_X1 U7553 ( .A(n9914), .B(n9913), .ZN(n12949) );
  NAND2_X2 U7554 ( .A1(n12822), .A2(n12821), .ZN(n14734) );
  NAND2_X1 U7555 ( .A1(n9648), .A2(n9647), .ZN(n9914) );
  NAND2_X1 U7556 ( .A1(n14579), .A2(n12902), .ZN(n14578) );
  AND2_X1 U7557 ( .A1(n9972), .A2(n9971), .ZN(n13959) );
  NAND2_X1 U7558 ( .A1(n9644), .A2(n9643), .ZN(n9648) );
  AND2_X1 U7559 ( .A1(n6970), .A2(n7625), .ZN(n6969) );
  NAND2_X1 U7560 ( .A1(n12806), .A2(n12805), .ZN(n14508) );
  NAND2_X1 U7561 ( .A1(n9627), .A2(n6806), .ZN(n9644) );
  NAND2_X1 U7562 ( .A1(n14014), .A2(n7412), .ZN(n7411) );
  NOR2_X1 U7563 ( .A1(n14533), .A2(n7626), .ZN(n7625) );
  NAND2_X1 U7564 ( .A1(n9611), .A2(n9610), .ZN(n14116) );
  OR2_X1 U7565 ( .A1(n7628), .A2(n14562), .ZN(n6970) );
  OAI21_X1 U7566 ( .B1(n12713), .B2(n12712), .A(n12711), .ZN(n12715) );
  CLKBUF_X1 U7567 ( .A(n14641), .Z(n6860) );
  NAND2_X1 U7568 ( .A1(n7266), .A2(n7269), .ZN(n14016) );
  XNOR2_X1 U7569 ( .A(n14757), .B(n6822), .ZN(n14550) );
  AND2_X1 U7570 ( .A1(n12907), .A2(n12837), .ZN(n14533) );
  AOI21_X1 U7571 ( .B1(n6925), .B2(n6924), .A(n13713), .ZN(n6923) );
  XNOR2_X1 U7572 ( .A(n9608), .B(n9593), .ZN(n12792) );
  NAND2_X1 U7573 ( .A1(n9592), .A2(n9591), .ZN(n9608) );
  AND2_X1 U7574 ( .A1(n9572), .A2(n9562), .ZN(n12746) );
  NAND2_X1 U7575 ( .A1(n7259), .A2(n6736), .ZN(n14063) );
  XNOR2_X1 U7576 ( .A(n9585), .B(n9586), .ZN(n12771) );
  NAND2_X1 U7577 ( .A1(n7336), .A2(n9571), .ZN(n9585) );
  AND2_X1 U7578 ( .A1(n6971), .A2(n12928), .ZN(n6696) );
  NAND2_X1 U7579 ( .A1(n6829), .A2(SI_24_), .ZN(n9571) );
  NOR2_X1 U7580 ( .A1(n13837), .A2(n13702), .ZN(n7533) );
  NAND2_X1 U7581 ( .A1(n14877), .A2(n12738), .ZN(n14843) );
  NAND2_X1 U7582 ( .A1(n8676), .A2(n8675), .ZN(n13288) );
  AOI21_X1 U7583 ( .B1(n13694), .B2(n13693), .A(n6912), .ZN(n13795) );
  NAND2_X1 U7584 ( .A1(n12663), .A2(n12662), .ZN(n14794) );
  XNOR2_X1 U7585 ( .A(n6914), .B(n13692), .ZN(n13694) );
  NAND2_X1 U7586 ( .A1(n9441), .A2(n9440), .ZN(n14161) );
  NAND2_X1 U7587 ( .A1(n8653), .A2(n8652), .ZN(n13274) );
  NAND2_X1 U7588 ( .A1(n9509), .A2(n9508), .ZN(n14146) );
  NAND2_X1 U7589 ( .A1(n12725), .A2(n12724), .ZN(n14601) );
  NAND2_X1 U7590 ( .A1(n12651), .A2(n12650), .ZN(n14650) );
  NAND2_X1 U7591 ( .A1(n12357), .A2(n12356), .ZN(n6914) );
  AND2_X1 U7592 ( .A1(n9483), .A2(n9482), .ZN(n14052) );
  NAND2_X1 U7593 ( .A1(n12710), .A2(n12709), .ZN(n14633) );
  NAND2_X1 U7594 ( .A1(n15371), .A2(n12226), .ZN(n12228) );
  NAND2_X1 U7595 ( .A1(n9499), .A2(n9481), .ZN(n12707) );
  XNOR2_X1 U7596 ( .A(n6933), .B(n13361), .ZN(n13348) );
  NOR2_X1 U7597 ( .A1(n15513), .A2(n6798), .ZN(n6933) );
  NAND2_X1 U7598 ( .A1(n9397), .A2(n9396), .ZN(n14975) );
  NAND2_X1 U7599 ( .A1(n12630), .A2(n12629), .ZN(n14807) );
  OR2_X1 U7600 ( .A1(n9475), .A2(n10541), .ZN(n9453) );
  OAI21_X1 U7601 ( .B1(n9433), .B2(n6676), .A(n7314), .ZN(n9501) );
  NAND2_X1 U7602 ( .A1(n12446), .A2(n12445), .ZN(n14810) );
  NAND2_X1 U7603 ( .A1(n9429), .A2(n9428), .ZN(n9433) );
  OAI21_X1 U7604 ( .B1(n11895), .B2(n7155), .A(n7154), .ZN(n15494) );
  AND2_X1 U7605 ( .A1(n9296), .A2(n9295), .ZN(n11680) );
  NOR2_X1 U7606 ( .A1(n11154), .A2(n6873), .ZN(n7731) );
  OR2_X1 U7607 ( .A1(n9354), .A2(SI_14_), .ZN(n9369) );
  OAI21_X1 U7608 ( .B1(n9353), .B2(n9352), .A(n9351), .ZN(n9354) );
  NAND2_X1 U7609 ( .A1(n9291), .A2(n9290), .ZN(n9293) );
  NAND2_X1 U7610 ( .A1(n11340), .A2(n11339), .ZN(n15158) );
  AND2_X1 U7611 ( .A1(n9218), .A2(n9217), .ZN(n11265) );
  CLKBUF_X1 U7612 ( .A(n10988), .Z(n15139) );
  AOI21_X1 U7613 ( .B1(n14380), .B2(n13038), .A(n10494), .ZN(n10627) );
  NAND2_X1 U7614 ( .A1(n8821), .A2(n8824), .ZN(n11742) );
  INV_X1 U7615 ( .A(n12974), .ZN(n13087) );
  AND2_X1 U7616 ( .A1(n9170), .A2(n9169), .ZN(n15332) );
  NAND2_X1 U7617 ( .A1(n9129), .A2(n9130), .ZN(n15314) );
  NAND2_X1 U7618 ( .A1(n10617), .A2(n12465), .ZN(n12974) );
  INV_X1 U7619 ( .A(n10616), .ZN(n13026) );
  NAND2_X1 U7620 ( .A1(n9194), .A2(n9193), .ZN(n9212) );
  AND4_X1 U7621 ( .A1(n8438), .A2(n8437), .A3(n8436), .A4(n8435), .ZN(n11755)
         );
  BUF_X2 U7622 ( .A(n11689), .Z(n12812) );
  NOR2_X1 U7623 ( .A1(n15608), .A2(n7912), .ZN(n7914) );
  CLKBUF_X3 U7624 ( .A(n8449), .Z(n8757) );
  INV_X2 U7625 ( .A(n13329), .ZN(n6667) );
  CLKBUF_X1 U7626 ( .A(n10734), .Z(n13735) );
  NAND2_X2 U7627 ( .A1(n10884), .A2(n10620), .ZN(n10886) );
  XNOR2_X1 U7628 ( .A(n10031), .B(n10035), .ZN(n12324) );
  AND2_X2 U7629 ( .A1(n10888), .A2(n12478), .ZN(n14811) );
  NAND2_X2 U7631 ( .A1(n8361), .A2(n10170), .ZN(n8663) );
  INV_X2 U7632 ( .A(n12721), .ZN(n12819) );
  OR2_X1 U7633 ( .A1(n9928), .A2(n10079), .ZN(n9116) );
  INV_X1 U7634 ( .A(n12474), .ZN(n14878) );
  OR2_X1 U7635 ( .A1(n9192), .A2(n9191), .ZN(n9193) );
  CLKBUF_X1 U7636 ( .A(n12947), .Z(n6812) );
  OAI21_X1 U7637 ( .B1(n10032), .B2(P1_IR_REG_24__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n10031) );
  INV_X2 U7638 ( .A(n9096), .ZN(n10062) );
  XNOR2_X1 U7639 ( .A(n10213), .B(n10212), .ZN(n12474) );
  NAND2_X1 U7640 ( .A1(n9096), .A2(n10170), .ZN(n9150) );
  NAND2_X1 U7641 ( .A1(n9070), .A2(n14194), .ZN(n9420) );
  MUX2_X1 U7642 ( .A(P3_IR_REG_31__SCAN_IN), .B(n8381), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n8382) );
  OR2_X1 U7643 ( .A1(n9190), .A2(n9197), .ZN(n9188) );
  NOR2_X1 U7644 ( .A1(n7739), .A2(P3_IR_REG_17__SCAN_IN), .ZN(n6874) );
  NAND2_X4 U7645 ( .A1(n9668), .A2(n10070), .ZN(n9096) );
  XNOR2_X1 U7646 ( .A(n7697), .B(n7696), .ZN(n15483) );
  NAND2_X1 U7647 ( .A1(n14862), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10477) );
  NAND2_X2 U7648 ( .A1(n10170), .A2(P2_U3088), .ZN(n14201) );
  XNOR2_X1 U7649 ( .A(n7699), .B(P3_IR_REG_7__SCAN_IN), .ZN(n15464) );
  OR2_X1 U7650 ( .A1(n7139), .A2(n7715), .ZN(n7659) );
  CLKBUF_X1 U7651 ( .A(n9710), .Z(n11287) );
  NAND2_X1 U7652 ( .A1(n7376), .A2(n7375), .ZN(n10215) );
  OR2_X1 U7653 ( .A1(n10478), .A2(n14864), .ZN(n10480) );
  INV_X1 U7654 ( .A(n10489), .ZN(n7376) );
  NAND2_X1 U7655 ( .A1(n14190), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n7523) );
  AND2_X1 U7656 ( .A1(n7676), .A2(n7668), .ZN(n7674) );
  AND2_X1 U7657 ( .A1(n7749), .A2(n6770), .ZN(n7139) );
  NAND2_X1 U7658 ( .A1(n9082), .A2(n6737), .ZN(n14190) );
  AND2_X1 U7659 ( .A1(n7667), .A2(n7678), .ZN(n7676) );
  NAND2_X1 U7660 ( .A1(n7748), .A2(n7103), .ZN(n7102) );
  NAND2_X2 U7661 ( .A1(n8360), .A2(n8359), .ZN(n9181) );
  AND2_X1 U7662 ( .A1(n7624), .A2(n7237), .ZN(n7243) );
  XNOR2_X1 U7663 ( .A(n7712), .B(n7711), .ZN(n7766) );
  NOR2_X1 U7664 ( .A1(n10037), .A2(P1_IR_REG_20__SCAN_IN), .ZN(n7624) );
  AND2_X1 U7665 ( .A1(n7014), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n7907) );
  AND3_X1 U7666 ( .A1(n7107), .A2(n7106), .A3(n7105), .ZN(n7645) );
  NAND4_X1 U7667 ( .A1(n9066), .A2(n9065), .A3(n6825), .A4(n9064), .ZN(n9077)
         );
  AND4_X1 U7668 ( .A1(n10758), .A2(n10757), .A3(n10023), .A4(n10022), .ZN(
        n10026) );
  NOR2_X1 U7669 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), .ZN(
        n6825) );
  INV_X4 U7670 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NOR2_X1 U7671 ( .A1(P2_IR_REG_20__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), .ZN(
        n9065) );
  NOR2_X1 U7672 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_21__SCAN_IN), .ZN(
        n9066) );
  NOR2_X1 U7673 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .ZN(
        n9055) );
  NOR2_X1 U7674 ( .A1(P2_IR_REG_16__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n9056) );
  INV_X1 U7675 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n9080) );
  NOR2_X1 U7676 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n10234) );
  INV_X1 U7677 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n10133) );
  INV_X1 U7678 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n9254) );
  INV_X1 U7679 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n9064) );
  INV_X1 U7680 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n8355) );
  INV_X1 U7681 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n9313) );
  INV_X4 U7682 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X2 U7683 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n7709) );
  INV_X1 U7684 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n10212) );
  INV_X4 U7685 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7686 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10476) );
  NOR2_X1 U7687 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n10022) );
  NOR2_X1 U7688 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n10024) );
  INV_X1 U7689 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n10035) );
  OAI21_X2 U7690 ( .B1(n11866), .B2(n11865), .A(n14318), .ZN(n11871) );
  NOR2_X2 U7691 ( .A1(n13954), .A2(n14116), .ZN(n7058) );
  INV_X1 U7692 ( .A(n12702), .ZN(n6668) );
  OAI21_X2 U7693 ( .B1(n11558), .B2(n7393), .A(n7391), .ZN(n11593) );
  NAND2_X2 U7694 ( .A1(n7029), .A2(n9734), .ZN(n11558) );
  OAI21_X2 U7695 ( .B1(n11138), .B2(n7399), .A(n7019), .ZN(n11023) );
  NAND2_X2 U7696 ( .A1(n9728), .A2(n9727), .ZN(n11138) );
  INV_X1 U7697 ( .A(n9948), .ZN(n6669) );
  BUF_X4 U7698 ( .A(n9150), .Z(n9948) );
  OAI21_X2 U7699 ( .B1(n14046), .B2(n9746), .A(n9747), .ZN(n14042) );
  INV_X4 U7700 ( .A(n10170), .ZN(n9213) );
  NOR2_X2 U7701 ( .A1(n13969), .A2(n6723), .ZN(n13952) );
  NOR2_X2 U7702 ( .A1(n13970), .A2(n13971), .ZN(n13969) );
  INV_X1 U7703 ( .A(n15265), .ZN(n15272) );
  XNOR2_X2 U7704 ( .A(n13890), .B(n15271), .ZN(n15265) );
  NAND2_X1 U7705 ( .A1(n10691), .A2(n9763), .ZN(n11466) );
  NAND4_X2 U7706 ( .A1(n9101), .A2(n9100), .A3(n9099), .A4(n9098), .ZN(n9763)
         );
  AOI21_X2 U7707 ( .B1(n13952), .B2(n9754), .A(n6884), .ZN(n13939) );
  AOI21_X1 U7708 ( .B1(n7489), .B2(n7492), .A(n7487), .ZN(n7486) );
  INV_X1 U7709 ( .A(n9876), .ZN(n7487) );
  NOR2_X1 U7710 ( .A1(n9350), .A2(SI_13_), .ZN(n9352) );
  INV_X1 U7711 ( .A(n9349), .ZN(n9350) );
  OR2_X1 U7712 ( .A1(n14933), .A2(n13140), .ZN(n8873) );
  INV_X1 U7713 ( .A(n14194), .ZN(n9072) );
  NOR2_X1 U7714 ( .A1(n9655), .A2(P2_IR_REG_19__SCAN_IN), .ZN(n9659) );
  NAND2_X1 U7715 ( .A1(n13275), .A2(n6726), .ZN(n13226) );
  INV_X1 U7716 ( .A(n13229), .ZN(n13160) );
  AND2_X1 U7717 ( .A1(n8743), .A2(n8742), .ZN(n13218) );
  AOI21_X1 U7718 ( .B1(n13461), .B2(n8757), .A(n8706), .ZN(n13265) );
  NOR2_X1 U7719 ( .A1(n7543), .A2(n13786), .ZN(n7542) );
  NOR2_X1 U7720 ( .A1(n13813), .A2(n6677), .ZN(n7543) );
  NAND2_X1 U7721 ( .A1(n12738), .A2(n10170), .ZN(n12721) );
  NAND2_X1 U7722 ( .A1(n9763), .A2(n9767), .ZN(n7419) );
  OR2_X1 U7723 ( .A1(n9811), .A2(n7425), .ZN(n7422) );
  AND2_X1 U7724 ( .A1(n7425), .A2(n9811), .ZN(n7424) );
  NAND2_X1 U7725 ( .A1(n7481), .A2(n7480), .ZN(n7479) );
  NAND2_X1 U7726 ( .A1(n7453), .A2(n9885), .ZN(n7452) );
  NAND2_X1 U7727 ( .A1(n7456), .A2(n7454), .ZN(n7453) );
  NAND2_X1 U7728 ( .A1(n7578), .A2(n7577), .ZN(n7576) );
  INV_X1 U7729 ( .A(n12739), .ZN(n7577) );
  INV_X1 U7730 ( .A(n12740), .ZN(n7578) );
  AND2_X1 U7731 ( .A1(n6947), .A2(n12807), .ZN(n6946) );
  NAND2_X1 U7732 ( .A1(n6690), .A2(n12808), .ZN(n6947) );
  NAND2_X1 U7733 ( .A1(n7771), .A2(n8429), .ZN(n7772) );
  NAND2_X1 U7734 ( .A1(n9389), .A2(n10442), .ZN(n9408) );
  OR2_X1 U7735 ( .A1(n10704), .A2(n11039), .ZN(n10702) );
  NAND2_X1 U7736 ( .A1(n8395), .A2(n7220), .ZN(n8772) );
  AND2_X1 U7737 ( .A1(n7221), .A2(n8394), .ZN(n7220) );
  INV_X1 U7738 ( .A(n13685), .ZN(n8384) );
  NOR2_X1 U7739 ( .A1(n15496), .A2(n6789), .ZN(n7786) );
  NAND2_X1 U7740 ( .A1(n7066), .A2(n7068), .ZN(n7065) );
  OR2_X1 U7741 ( .A1(n13274), .A2(n13519), .ZN(n8898) );
  OR2_X1 U7742 ( .A1(n13128), .A2(n13219), .ZN(n8931) );
  NAND2_X1 U7743 ( .A1(n7748), .A2(n7504), .ZN(n7503) );
  NOR2_X1 U7744 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_27__SCAN_IN), .ZN(
        n7504) );
  AOI21_X1 U7745 ( .B1(n7235), .B2(n7233), .A(n6795), .ZN(n7232) );
  INV_X1 U7746 ( .A(n7235), .ZN(n7234) );
  NAND2_X1 U7747 ( .A1(n8549), .A2(n8323), .ZN(n8324) );
  INV_X1 U7748 ( .A(P3_IR_REG_13__SCAN_IN), .ZN(n7497) );
  NAND2_X1 U7749 ( .A1(n10188), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n8308) );
  NAND2_X1 U7750 ( .A1(n7687), .A2(n7716), .ZN(n7705) );
  NAND2_X1 U7751 ( .A1(n10186), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n8303) );
  INV_X1 U7752 ( .A(P3_IR_REG_3__SCAN_IN), .ZN(n7716) );
  NAND2_X1 U7753 ( .A1(n14126), .A2(n9895), .ZN(n7298) );
  AND2_X1 U7754 ( .A1(n6763), .A2(n9745), .ZN(n7404) );
  NOR2_X1 U7755 ( .A1(n14029), .A2(n7273), .ZN(n7272) );
  INV_X1 U7756 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n9660) );
  NOR2_X1 U7757 ( .A1(P2_IR_REG_18__SCAN_IN), .A2(n9060), .ZN(n6929) );
  INV_X1 U7758 ( .A(n14274), .ZN(n7348) );
  AOI21_X1 U7759 ( .B1(n14274), .B2(n7347), .A(n7346), .ZN(n7345) );
  NOR2_X1 U7760 ( .A1(n14609), .A2(n7617), .ZN(n7616) );
  INV_X1 U7761 ( .A(n12926), .ZN(n7617) );
  NAND2_X1 U7762 ( .A1(n6989), .A2(n14697), .ZN(n6988) );
  NAND2_X1 U7763 ( .A1(n12915), .A2(n12917), .ZN(n6989) );
  AND2_X1 U7764 ( .A1(n9388), .A2(n9374), .ZN(n9386) );
  INV_X1 U7765 ( .A(n9370), .ZN(n7326) );
  XNOR2_X1 U7766 ( .A(n9308), .B(SI_11_), .ZN(n9311) );
  INV_X1 U7767 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n10140) );
  AOI21_X1 U7768 ( .B1(n7123), .B2(n7125), .A(n11715), .ZN(n7122) );
  INV_X1 U7769 ( .A(n13494), .ZN(n13197) );
  AND2_X1 U7770 ( .A1(n11095), .A2(n11093), .ZN(n7147) );
  NAND2_X1 U7771 ( .A1(n8365), .A2(n8364), .ZN(n8559) );
  INV_X1 U7772 ( .A(n8540), .ZN(n8365) );
  NAND2_X1 U7773 ( .A1(n13226), .A2(n13162), .ZN(n13195) );
  CLKBUF_X1 U7774 ( .A(n8668), .Z(n6813) );
  AND2_X2 U7775 ( .A1(n13685), .A2(n8383), .ZN(n8668) );
  NAND2_X1 U7776 ( .A1(n7153), .A2(n7152), .ZN(n7151) );
  INV_X1 U7777 ( .A(n15445), .ZN(n7152) );
  OR2_X1 U7778 ( .A1(n13341), .A2(n14947), .ZN(n6941) );
  NOR2_X1 U7779 ( .A1(n8597), .A2(n7738), .ZN(n6869) );
  NOR2_X1 U7780 ( .A1(n13383), .A2(n7789), .ZN(n14920) );
  OR2_X1 U7781 ( .A1(n14920), .A2(n14919), .ZN(n6940) );
  AND2_X1 U7782 ( .A1(n7086), .A2(n7085), .ZN(n9044) );
  AND2_X1 U7783 ( .A1(n9040), .A2(n8744), .ZN(n13417) );
  OAI21_X1 U7784 ( .B1(n13498), .B2(n13284), .A(n13491), .ZN(n13481) );
  NOR2_X1 U7785 ( .A1(n13544), .A2(n13150), .ZN(n7071) );
  OR2_X1 U7786 ( .A1(n13544), .A2(n13517), .ZN(n8885) );
  AOI21_X1 U7787 ( .B1(n7428), .B2(n7431), .A(n8880), .ZN(n7426) );
  AND2_X1 U7788 ( .A1(n7429), .A2(n13556), .ZN(n7428) );
  NAND2_X1 U7789 ( .A1(n8977), .A2(n6691), .ZN(n7088) );
  NAND2_X1 U7790 ( .A1(n11756), .A2(n8960), .ZN(n11540) );
  INV_X1 U7791 ( .A(n8663), .ZN(n8760) );
  INV_X1 U7792 ( .A(n8761), .ZN(n8637) );
  NAND2_X1 U7793 ( .A1(n8350), .A2(n8349), .ZN(n8731) );
  OR2_X1 U7794 ( .A1(n8719), .A2(n8348), .ZN(n8350) );
  AND2_X1 U7795 ( .A1(n8323), .A2(n8322), .ZN(n8546) );
  AOI21_X1 U7796 ( .B1(n8534), .B2(n7189), .A(n7188), .ZN(n7187) );
  INV_X1 U7797 ( .A(n8321), .ZN(n7188) );
  INV_X1 U7798 ( .A(n8319), .ZN(n7189) );
  INV_X1 U7799 ( .A(n8534), .ZN(n7190) );
  NAND2_X1 U7800 ( .A1(n8466), .A2(n8309), .ZN(n8311) );
  NAND2_X1 U7801 ( .A1(n10182), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n8306) );
  OAI21_X1 U7802 ( .B1(n6905), .B2(n13772), .A(n6901), .ZN(n6900) );
  NAND2_X1 U7803 ( .A1(n6905), .A2(n6902), .ZN(n6901) );
  NAND2_X1 U7804 ( .A1(n6903), .A2(n6907), .ZN(n6902) );
  NAND2_X1 U7805 ( .A1(n9575), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n9597) );
  XNOR2_X1 U7806 ( .A(n10726), .B(n15306), .ZN(n10737) );
  NAND2_X1 U7807 ( .A1(n7541), .A2(n7539), .ZN(n6817) );
  INV_X1 U7808 ( .A(n13849), .ZN(n7539) );
  AND2_X1 U7809 ( .A1(n9605), .A2(n9604), .ZN(n13789) );
  AND2_X1 U7810 ( .A1(n9493), .A2(n9492), .ZN(n13759) );
  AND4_X1 U7811 ( .A1(n9178), .A2(n9177), .A3(n9176), .A4(n9175), .ZN(n9794)
         );
  NOR2_X1 U7812 ( .A1(n7409), .A2(n7408), .ZN(n7407) );
  INV_X1 U7813 ( .A(n7410), .ZN(n7409) );
  NOR2_X1 U7814 ( .A1(n14036), .A2(n14029), .ZN(n14025) );
  AND2_X1 U7815 ( .A1(n14969), .A2(n9742), .ZN(n7401) );
  INV_X1 U7816 ( .A(n9348), .ZN(n7282) );
  NAND2_X1 U7817 ( .A1(n7284), .A2(n6701), .ZN(n7283) );
  INV_X1 U7818 ( .A(n11879), .ZN(n7284) );
  NAND2_X1 U7819 ( .A1(n10947), .A2(n10946), .ZN(n7256) );
  AND2_X1 U7820 ( .A1(n9687), .A2(n9704), .ZN(n15283) );
  NAND2_X1 U7821 ( .A1(n12738), .A2(n9213), .ZN(n10978) );
  INV_X1 U7822 ( .A(n10622), .ZN(n10625) );
  NAND2_X1 U7823 ( .A1(n14507), .A2(n7618), .ZN(n13098) );
  NOR2_X1 U7824 ( .A1(n12939), .A2(n7619), .ZN(n7618) );
  INV_X1 U7825 ( .A(n12937), .ZN(n7619) );
  NAND2_X1 U7826 ( .A1(n14567), .A2(n7627), .ZN(n14543) );
  NAND2_X1 U7827 ( .A1(n14678), .A2(n12896), .ZN(n7204) );
  NOR2_X1 U7828 ( .A1(n12854), .A2(n7615), .ZN(n7614) );
  INV_X1 U7829 ( .A(n12295), .ZN(n7615) );
  NOR2_X1 U7830 ( .A1(n6982), .A2(n6981), .ZN(n6980) );
  INV_X1 U7831 ( .A(n7608), .ZN(n6981) );
  NOR2_X1 U7832 ( .A1(n6671), .A2(n11832), .ZN(n6982) );
  AOI21_X1 U7833 ( .B1(n12087), .B2(n7609), .A(n6739), .ZN(n7608) );
  OR2_X1 U7834 ( .A1(n7610), .A2(n7607), .ZN(n6671) );
  OR2_X1 U7835 ( .A1(n12659), .A2(n12721), .ZN(n12663) );
  INV_X1 U7836 ( .A(n12738), .ZN(n12660) );
  OR2_X1 U7837 ( .A1(n9480), .A2(n9500), .ZN(n9499) );
  NAND2_X1 U7838 ( .A1(n10141), .A2(n10140), .ZN(n10761) );
  AND2_X1 U7839 ( .A1(n10135), .A2(n10137), .ZN(n10141) );
  INV_X1 U7840 ( .A(n13267), .ZN(n7130) );
  NOR2_X1 U7841 ( .A1(n7537), .A2(n13733), .ZN(n7536) );
  INV_X1 U7842 ( .A(n7542), .ZN(n7537) );
  NAND2_X1 U7843 ( .A1(n12273), .A2(n12272), .ZN(n15060) );
  NAND2_X1 U7844 ( .A1(n12552), .A2(n11578), .ZN(n7565) );
  NAND2_X1 U7845 ( .A1(n12551), .A2(n15139), .ZN(n7566) );
  INV_X1 U7846 ( .A(n9801), .ZN(n7444) );
  NAND2_X1 U7847 ( .A1(n7423), .A2(n6735), .ZN(n9817) );
  NAND2_X1 U7848 ( .A1(n12591), .A2(n7560), .ZN(n7559) );
  INV_X1 U7849 ( .A(n12590), .ZN(n7560) );
  INV_X1 U7850 ( .A(n9824), .ZN(n7502) );
  INV_X1 U7851 ( .A(n7479), .ZN(n7478) );
  AND2_X1 U7852 ( .A1(n7633), .A2(n7476), .ZN(n7475) );
  NAND2_X1 U7853 ( .A1(n7479), .A2(n7477), .ZN(n7476) );
  NOR2_X1 U7854 ( .A1(n14642), .A2(n7632), .ZN(n12689) );
  NAND2_X1 U7855 ( .A1(n7484), .A2(n7483), .ZN(n7482) );
  OR2_X1 U7856 ( .A1(n7486), .A2(n7491), .ZN(n7485) );
  AND2_X1 U7857 ( .A1(n9882), .A2(n9884), .ZN(n7456) );
  INV_X1 U7858 ( .A(n7451), .ZN(n7450) );
  OAI21_X1 U7859 ( .B1(n7452), .B2(n7454), .A(n9886), .ZN(n7451) );
  NOR2_X1 U7860 ( .A1(n9885), .A2(n7449), .ZN(n7448) );
  INV_X1 U7861 ( .A(n7454), .ZN(n7449) );
  INV_X1 U7862 ( .A(n12760), .ZN(n7557) );
  AND2_X1 U7863 ( .A1(n7555), .A2(n12778), .ZN(n7553) );
  NAND2_X1 U7864 ( .A1(n6678), .A2(n7556), .ZN(n7555) );
  OAI21_X1 U7865 ( .B1(n12741), .B2(n7575), .A(n7572), .ZN(n12743) );
  NAND2_X1 U7866 ( .A1(n7580), .A2(n12745), .ZN(n7575) );
  OR2_X1 U7867 ( .A1(n7557), .A2(n12762), .ZN(n7556) );
  NAND2_X1 U7868 ( .A1(n9909), .A2(n6710), .ZN(n7436) );
  NAND2_X1 U7869 ( .A1(n12825), .A2(n7583), .ZN(n7582) );
  INV_X1 U7870 ( .A(n12824), .ZN(n7583) );
  NAND2_X1 U7871 ( .A1(n6757), .A2(n6944), .ZN(n6943) );
  NAND2_X1 U7872 ( .A1(n12797), .A2(n7591), .ZN(n7590) );
  NAND2_X1 U7873 ( .A1(n6946), .A2(n12809), .ZN(n6945) );
  INV_X1 U7874 ( .A(n9585), .ZN(n9588) );
  OAI21_X1 U7875 ( .B1(n9557), .B2(n9556), .A(n9555), .ZN(n9558) );
  INV_X1 U7876 ( .A(n7315), .ZN(n7314) );
  OAI21_X1 U7877 ( .B1(n7316), .B2(n6676), .A(n9478), .ZN(n7315) );
  NOR2_X1 U7878 ( .A1(n9474), .A2(n7317), .ZN(n7316) );
  AND2_X1 U7879 ( .A1(n7323), .A2(n9329), .ZN(n7319) );
  INV_X1 U7880 ( .A(n9310), .ZN(n7321) );
  INV_X1 U7881 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n8364) );
  NAND2_X1 U7882 ( .A1(n10770), .A2(n8804), .ZN(n10712) );
  NAND2_X1 U7883 ( .A1(P3_REG2_REG_2__SCAN_IN), .A2(n7766), .ZN(n7713) );
  INV_X1 U7884 ( .A(n7713), .ZN(n7714) );
  AOI21_X1 U7885 ( .B1(P3_REG1_REG_6__SCAN_IN), .B2(n15442), .A(n15439), .ZN(
        n7777) );
  AND2_X1 U7886 ( .A1(n7151), .A2(n7150), .ZN(n7725) );
  NAND2_X1 U7887 ( .A1(n15442), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7150) );
  NOR2_X1 U7888 ( .A1(n11152), .A2(n6810), .ZN(n7783) );
  AND2_X1 U7889 ( .A1(n10163), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n6810) );
  INV_X1 U7890 ( .A(n8751), .ZN(n13123) );
  INV_X1 U7891 ( .A(n6702), .ZN(n7093) );
  OR2_X1 U7892 ( .A1(n13454), .A2(n13455), .ZN(n8800) );
  NAND2_X1 U7893 ( .A1(n13274), .A2(n13493), .ZN(n7074) );
  AOI21_X1 U7894 ( .B1(n7080), .B2(n8971), .A(n6740), .ZN(n7079) );
  INV_X1 U7895 ( .A(n8970), .ZN(n7080) );
  INV_X1 U7896 ( .A(n8971), .ZN(n7081) );
  NOR2_X1 U7897 ( .A1(n11778), .A2(n7114), .ZN(n7113) );
  INV_X1 U7898 ( .A(n8967), .ZN(n7114) );
  NAND2_X1 U7899 ( .A1(n8961), .A2(n8445), .ZN(n11539) );
  INV_X1 U7900 ( .A(P3_IR_REG_23__SCAN_IN), .ZN(n7664) );
  INV_X1 U7901 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7653) );
  INV_X1 U7902 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7647) );
  INV_X1 U7903 ( .A(n8476), .ZN(n7208) );
  NOR2_X1 U7904 ( .A1(n7527), .A2(n13709), .ZN(n7526) );
  INV_X1 U7905 ( .A(n7533), .ZN(n7527) );
  NAND2_X1 U7906 ( .A1(n7293), .A2(n9972), .ZN(n7292) );
  XNOR2_X1 U7907 ( .A(n14131), .B(n13867), .ZN(n7408) );
  NOR2_X1 U7908 ( .A1(n9516), .A2(n7268), .ZN(n7267) );
  INV_X1 U7909 ( .A(n9495), .ZN(n7268) );
  INV_X1 U7910 ( .A(n7271), .ZN(n7270) );
  AOI21_X1 U7911 ( .B1(n14054), .B2(n9495), .A(n6742), .ZN(n7271) );
  INV_X1 U7912 ( .A(n9735), .ZN(n7395) );
  INV_X1 U7913 ( .A(n11562), .ZN(n7392) );
  NAND2_X1 U7914 ( .A1(n9757), .A2(n9710), .ZN(n10723) );
  NOR2_X1 U7915 ( .A1(n11022), .A2(n10942), .ZN(n7253) );
  INV_X1 U7916 ( .A(n9210), .ZN(n7255) );
  AND2_X1 U7917 ( .A1(n10942), .A2(n7398), .ZN(n7020) );
  INV_X1 U7918 ( .A(n12282), .ZN(n7265) );
  NOR2_X1 U7919 ( .A1(n9077), .A2(n9068), .ZN(n7257) );
  OR2_X1 U7920 ( .A1(n13008), .A2(n14283), .ZN(n13016) );
  NAND2_X1 U7921 ( .A1(n14258), .A2(n12983), .ZN(n7387) );
  INV_X1 U7922 ( .A(n14265), .ZN(n7383) );
  INV_X1 U7923 ( .A(n12983), .ZN(n7384) );
  INV_X1 U7924 ( .A(n14291), .ZN(n7339) );
  OR2_X1 U7925 ( .A1(n13101), .A2(n14734), .ZN(n7039) );
  NOR2_X1 U7926 ( .A1(n7605), .A2(n7601), .ZN(n7600) );
  NAND2_X1 U7927 ( .A1(n6986), .A2(n6988), .ZN(n6984) );
  INV_X1 U7928 ( .A(n12919), .ZN(n7601) );
  NAND2_X1 U7929 ( .A1(n12921), .A2(n7604), .ZN(n7603) );
  INV_X1 U7930 ( .A(n12920), .ZN(n7604) );
  OR2_X1 U7931 ( .A1(n15050), .A2(n14295), .ZN(n12613) );
  NAND2_X1 U7932 ( .A1(n6868), .A2(n12530), .ZN(n11356) );
  OAI21_X1 U7933 ( .B1(n12951), .B2(n11629), .A(n7620), .ZN(n7621) );
  NAND2_X1 U7934 ( .A1(n12951), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n7620) );
  AND2_X1 U7935 ( .A1(n14599), .A2(n14843), .ZN(n14589) );
  NAND2_X1 U7936 ( .A1(n7239), .A2(n7243), .ZN(n10211) );
  NOR2_X1 U7937 ( .A1(n10495), .A2(n7240), .ZN(n7239) );
  NAND2_X1 U7938 ( .A1(n7241), .A2(n7242), .ZN(n7240) );
  NOR2_X1 U7939 ( .A1(n9607), .A2(SI_26_), .ZN(n7328) );
  INV_X1 U7940 ( .A(n9607), .ZN(n7327) );
  NAND2_X1 U7941 ( .A1(n9559), .A2(n9571), .ZN(n9561) );
  INV_X1 U7942 ( .A(n9500), .ZN(n9502) );
  INV_X1 U7943 ( .A(n9473), .ZN(n6957) );
  INV_X1 U7944 ( .A(n9453), .ZN(n6959) );
  NAND2_X1 U7945 ( .A1(n9434), .A2(n9470), .ZN(n6960) );
  NAND2_X1 U7946 ( .A1(n9433), .A2(n9432), .ZN(n9475) );
  AOI21_X1 U7947 ( .B1(n6952), .B2(n6954), .A(n6950), .ZN(n6949) );
  INV_X1 U7948 ( .A(n9408), .ZN(n6950) );
  AND2_X1 U7949 ( .A1(n9408), .A2(n9391), .ZN(n9406) );
  NAND2_X1 U7950 ( .A1(n9372), .A2(n10316), .ZN(n9388) );
  NAND2_X1 U7951 ( .A1(n9275), .A2(SI_10_), .ZN(n9292) );
  INV_X1 U7952 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n10137) );
  XNOR2_X1 U7953 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n7906) );
  NAND2_X1 U7954 ( .A1(n6994), .A2(n6992), .ZN(n7863) );
  NAND2_X1 U7955 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6993), .ZN(n6992) );
  INV_X1 U7956 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6993) );
  NAND2_X1 U7957 ( .A1(n6999), .A2(n7867), .ZN(n7869) );
  NAND2_X1 U7958 ( .A1(n6694), .A2(n10669), .ZN(n6999) );
  XNOR2_X1 U7959 ( .A(n7869), .B(n7868), .ZN(n7913) );
  OAI21_X1 U7960 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n15453), .A(n7872), .ZN(
        n7873) );
  OAI21_X1 U7961 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n15493), .A(n7876), .ZN(
        n7899) );
  OAI21_X1 U7962 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n7882), .A(n7881), .ZN(
        n7895) );
  AOI21_X1 U7963 ( .B1(n7126), .B2(n7124), .A(n6717), .ZN(n7123) );
  INV_X1 U7964 ( .A(n11710), .ZN(n7124) );
  INV_X1 U7965 ( .A(n7126), .ZN(n7125) );
  INV_X1 U7966 ( .A(n15374), .ZN(n6876) );
  XNOR2_X1 U7967 ( .A(n12432), .B(n11759), .ZN(n11090) );
  INV_X1 U7968 ( .A(n13174), .ZN(n13215) );
  INV_X1 U7969 ( .A(n8712), .ZN(n8375) );
  AND3_X1 U7970 ( .A1(n8421), .A2(n8420), .A3(n8419), .ZN(n11309) );
  OR2_X1 U7971 ( .A1(n8761), .A2(SI_2_), .ZN(n8421) );
  AND2_X1 U7972 ( .A1(n6708), .A2(n15392), .ZN(n7126) );
  XNOR2_X1 U7973 ( .A(n7458), .B(n9014), .ZN(n6835) );
  NOR2_X1 U7974 ( .A1(n8934), .A2(n6712), .ZN(n7459) );
  INV_X1 U7975 ( .A(n6813), .ZN(n8767) );
  AND4_X1 U7976 ( .A1(n8464), .A2(n8463), .A3(n8462), .A4(n8461), .ZN(n11942)
         );
  AND4_X1 U7977 ( .A1(n8453), .A2(n8452), .A3(n8451), .A4(n8450), .ZN(n11767)
         );
  NOR2_X1 U7978 ( .A1(n15425), .A2(n7775), .ZN(n15441) );
  OR2_X1 U7979 ( .A1(n15422), .A2(n7723), .ZN(n7153) );
  XNOR2_X1 U7980 ( .A(n7777), .B(n15464), .ZN(n15462) );
  XNOR2_X1 U7981 ( .A(n7725), .B(n15464), .ZN(n15455) );
  NOR2_X1 U7982 ( .A1(n15456), .A2(n15455), .ZN(n15454) );
  NAND2_X1 U7983 ( .A1(n6935), .A2(n6934), .ZN(n15480) );
  NAND2_X1 U7984 ( .A1(n7778), .A2(n6939), .ZN(n6934) );
  OR2_X1 U7985 ( .A1(n15462), .A2(n6936), .ZN(n6935) );
  NAND2_X1 U7986 ( .A1(n6939), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n6936) );
  OR2_X1 U7987 ( .A1(n15462), .A2(n15600), .ZN(n6938) );
  AND2_X1 U7988 ( .A1(n15483), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n6811) );
  AND2_X1 U7989 ( .A1(n10163), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n6873) );
  AND2_X1 U7990 ( .A1(n6941), .A2(n6758), .ZN(n15515) );
  NOR2_X1 U7991 ( .A1(n15515), .A2(n15514), .ZN(n15513) );
  NAND2_X1 U7992 ( .A1(n6872), .A2(n6871), .ZN(n6858) );
  NAND2_X1 U7993 ( .A1(n15500), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n6871) );
  INV_X1 U7994 ( .A(n15494), .ZN(n6872) );
  NOR2_X1 U7995 ( .A1(n13351), .A2(n13350), .ZN(n13349) );
  NAND2_X1 U7996 ( .A1(n13444), .A2(n7636), .ZN(n13432) );
  OR2_X1 U7997 ( .A1(n13641), .A2(n13268), .ZN(n7636) );
  NAND2_X1 U7998 ( .A1(n7091), .A2(n7470), .ZN(n7469) );
  INV_X1 U7999 ( .A(n8800), .ZN(n7470) );
  INV_X1 U8000 ( .A(n7468), .ZN(n7467) );
  OAI21_X1 U8001 ( .B1(n13447), .B2(n8798), .A(n8797), .ZN(n7468) );
  OR2_X1 U8002 ( .A1(n7099), .A2(n7098), .ZN(n7097) );
  INV_X1 U8003 ( .A(n7101), .ZN(n7098) );
  AND2_X1 U8004 ( .A1(n6715), .A2(n13466), .ZN(n7099) );
  NAND2_X1 U8005 ( .A1(n13481), .A2(n6702), .ZN(n7096) );
  NAND2_X1 U8006 ( .A1(n13492), .A2(n13496), .ZN(n13491) );
  AND3_X1 U8007 ( .A1(n8671), .A2(n8670), .A3(n8669), .ZN(n13506) );
  NAND2_X1 U8008 ( .A1(n13153), .A2(n13534), .ZN(n7075) );
  NAND2_X1 U8009 ( .A1(n7073), .A2(n13546), .ZN(n7072) );
  INV_X1 U8010 ( .A(n13529), .ZN(n7073) );
  NAND2_X1 U8011 ( .A1(n7088), .A2(n6727), .ZN(n13551) );
  AND2_X1 U8012 ( .A1(n8879), .A2(n8882), .ZN(n13556) );
  NAND2_X1 U8013 ( .A1(n8592), .A2(n8873), .ZN(n12371) );
  NAND2_X1 U8014 ( .A1(n12371), .A2(n12370), .ZN(n12369) );
  AND4_X1 U8015 ( .A1(n8545), .A2(n8544), .A3(n8543), .A4(n8542), .ZN(n12388)
         );
  NAND2_X1 U8016 ( .A1(n6847), .A2(n6846), .ZN(n7498) );
  INV_X1 U8017 ( .A(n8847), .ZN(n6846) );
  OR2_X1 U8018 ( .A1(n11941), .A2(n7112), .ZN(n7109) );
  INV_X1 U8019 ( .A(n7113), .ZN(n7112) );
  AOI21_X1 U8020 ( .B1(n7113), .B2(n8781), .A(n7111), .ZN(n7110) );
  NOR2_X1 U8021 ( .A1(n12004), .A2(n11721), .ZN(n7111) );
  AND4_X1 U8022 ( .A1(n8475), .A2(n8474), .A3(n8473), .A4(n8472), .ZN(n11780)
         );
  AND2_X1 U8023 ( .A1(n8839), .A2(n8846), .ZN(n11778) );
  AND3_X1 U8024 ( .A1(n8482), .A2(n8481), .A3(n8480), .ZN(n8966) );
  NAND2_X1 U8025 ( .A1(n11941), .A2(n11940), .ZN(n11939) );
  AND2_X1 U8026 ( .A1(n8830), .A2(n11937), .ZN(n11765) );
  AND3_X1 U8027 ( .A1(n8458), .A2(n8457), .A3(n8456), .ZN(n11550) );
  OR2_X1 U8028 ( .A1(n8663), .A2(n10127), .ZN(n8457) );
  NOR2_X1 U8029 ( .A1(n11753), .A2(n8954), .ZN(n8958) );
  INV_X1 U8030 ( .A(n13552), .ZN(n13515) );
  NAND2_X1 U8031 ( .A1(n8599), .A2(n8598), .ZN(n13143) );
  NAND2_X1 U8032 ( .A1(n9013), .A2(n11313), .ZN(n15582) );
  NAND2_X1 U8033 ( .A1(n8987), .A2(n9015), .ZN(n13520) );
  OAI22_X1 U8034 ( .A1(n8759), .A2(n8354), .B1(P2_DATAO_REG_29__SCAN_IN), .B2(
        n14193), .ZN(n8391) );
  XNOR2_X1 U8035 ( .A(n7661), .B(P3_IR_REG_26__SCAN_IN), .ZN(n8993) );
  OAI21_X1 U8036 ( .B1(n8698), .B2(n7247), .A(n7244), .ZN(n8719) );
  NAND2_X1 U8037 ( .A1(n8346), .A2(n12747), .ZN(n7247) );
  OAI21_X1 U8038 ( .B1(n8345), .B2(n7246), .A(n8347), .ZN(n7245) );
  OR2_X1 U8039 ( .A1(n8343), .A2(n12142), .ZN(n8345) );
  NOR2_X1 U8040 ( .A1(n7757), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n7754) );
  XNOR2_X1 U8041 ( .A(n7758), .B(P3_IR_REG_21__SCAN_IN), .ZN(n10704) );
  AND4_X1 U8042 ( .A1(n7650), .A2(n7649), .A3(n7648), .A4(n7678), .ZN(n7651)
         );
  INV_X1 U8043 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n7648) );
  INV_X1 U8044 ( .A(n7182), .ZN(n7181) );
  OAI21_X1 U8045 ( .B1(n8580), .B2(n7183), .A(n8593), .ZN(n7182) );
  INV_X1 U8046 ( .A(n8330), .ZN(n7183) );
  NAND2_X1 U8047 ( .A1(n8569), .A2(n8328), .ZN(n8581) );
  NAND2_X1 U8048 ( .A1(n8581), .A2(n8580), .ZN(n8583) );
  AND2_X1 U8049 ( .A1(n8326), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n7211) );
  NAND2_X1 U8050 ( .A1(n8324), .A2(n10287), .ZN(n8326) );
  INV_X1 U8051 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7107) );
  INV_X1 U8052 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7106) );
  INV_X1 U8053 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7105) );
  AND2_X1 U8054 ( .A1(n7643), .A2(n7642), .ZN(n7644) );
  NAND2_X1 U8055 ( .A1(n7186), .A2(n7184), .ZN(n8549) );
  AOI21_X1 U8056 ( .B1(n7187), .B2(n7190), .A(n7185), .ZN(n7184) );
  INV_X1 U8057 ( .A(n8546), .ZN(n7185) );
  AND2_X1 U8058 ( .A1(n8321), .A2(n8320), .ZN(n8534) );
  NAND2_X1 U8059 ( .A1(n8509), .A2(n8317), .ZN(n8521) );
  AND2_X1 U8060 ( .A1(n8319), .A2(n8318), .ZN(n8520) );
  OR2_X1 U8061 ( .A1(n7693), .A2(P3_IR_REG_9__SCAN_IN), .ZN(n7690) );
  AND2_X1 U8062 ( .A1(n7698), .A2(n7688), .ZN(n7695) );
  NAND2_X1 U8063 ( .A1(n10166), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n8313) );
  AND2_X1 U8064 ( .A1(n8315), .A2(n8314), .ZN(n8493) );
  OAI21_X1 U8065 ( .B1(n8311), .B2(n7207), .A(n7205), .ZN(n8496) );
  INV_X1 U8066 ( .A(n7206), .ZN(n7205) );
  OAI21_X1 U8067 ( .B1(n6703), .B2(n7207), .A(n8493), .ZN(n7206) );
  INV_X1 U8068 ( .A(n8313), .ZN(n7207) );
  NAND2_X1 U8069 ( .A1(n8311), .A2(n6703), .ZN(n8479) );
  AND2_X1 U8070 ( .A1(n7700), .A2(n7701), .ZN(n7698) );
  NAND2_X1 U8071 ( .A1(n7212), .A2(n7213), .ZN(n8466) );
  AOI21_X1 U8072 ( .B1(n7216), .B2(n7218), .A(n7214), .ZN(n7213) );
  INV_X1 U8073 ( .A(n8308), .ZN(n7214) );
  NOR2_X1 U8074 ( .A1(n7703), .A2(P3_IR_REG_5__SCAN_IN), .ZN(n7700) );
  INV_X1 U8075 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7701) );
  AND2_X1 U8076 ( .A1(n8308), .A2(n8307), .ZN(n8454) );
  OR2_X1 U8077 ( .A1(n7705), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n7703) );
  XNOR2_X1 U8078 ( .A(n7707), .B(n7706), .ZN(n15417) );
  INV_X1 U8079 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7706) );
  AND2_X1 U8080 ( .A1(n8306), .A2(n8305), .ZN(n8439) );
  NAND2_X1 U8081 ( .A1(n8301), .A2(n8300), .ZN(n8428) );
  OR2_X1 U8082 ( .A1(n7687), .A2(n7715), .ZN(n7717) );
  INV_X1 U8083 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7711) );
  NAND2_X1 U8084 ( .A1(n6817), .A2(n13732), .ZN(n7534) );
  NAND2_X1 U8085 ( .A1(n7551), .A2(n7550), .ZN(n12357) );
  AND2_X1 U8086 ( .A1(n12156), .A2(n12155), .ZN(n7550) );
  NAND2_X1 U8087 ( .A1(n12151), .A2(n12150), .ZN(n7551) );
  INV_X1 U8088 ( .A(n7526), .ZN(n6924) );
  INV_X1 U8089 ( .A(n9543), .ZN(n9541) );
  NAND2_X1 U8090 ( .A1(n11206), .A2(n11208), .ZN(n11203) );
  INV_X1 U8091 ( .A(n13821), .ZN(n6926) );
  NAND2_X1 U8092 ( .A1(n7525), .A2(n13708), .ZN(n7524) );
  INV_X1 U8093 ( .A(n7528), .ZN(n7525) );
  INV_X1 U8094 ( .A(n6919), .ZN(n6918) );
  OAI21_X1 U8095 ( .B1(n11672), .B2(n6920), .A(n11961), .ZN(n6919) );
  INV_X1 U8096 ( .A(n11922), .ZN(n6920) );
  NAND2_X1 U8097 ( .A1(n13803), .A2(n13804), .ZN(n13802) );
  AND2_X1 U8098 ( .A1(n10931), .A2(n10922), .ZN(n7546) );
  AOI21_X1 U8099 ( .B1(n7542), .B2(n6677), .A(n6753), .ZN(n7541) );
  INV_X1 U8100 ( .A(n13727), .ZN(n7544) );
  INV_X1 U8101 ( .A(n13728), .ZN(n7545) );
  AND2_X1 U8102 ( .A1(n9584), .A2(n9583), .ZN(n9895) );
  AND2_X1 U8103 ( .A1(n9467), .A2(n9466), .ZN(n13842) );
  AND3_X1 U8104 ( .A1(n9385), .A2(n9384), .A3(n9383), .ZN(n12358) );
  AND4_X1 U8105 ( .A1(n9305), .A2(n9304), .A3(n9303), .A4(n9302), .ZN(n11587)
         );
  AND4_X1 U8106 ( .A1(n9226), .A2(n9225), .A3(n9224), .A4(n9223), .ZN(n11075)
         );
  AND2_X1 U8107 ( .A1(n9630), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n9714) );
  INV_X1 U8108 ( .A(n9971), .ZN(n7290) );
  NOR2_X1 U8109 ( .A1(n9606), .A2(n7294), .ZN(n7291) );
  OR2_X1 U8110 ( .A1(n13982), .A2(n7292), .ZN(n7285) );
  AND2_X1 U8111 ( .A1(n14122), .A2(n13865), .ZN(n6884) );
  NAND2_X1 U8112 ( .A1(n7296), .A2(n7298), .ZN(n7293) );
  NAND2_X1 U8113 ( .A1(n7297), .A2(n13971), .ZN(n7296) );
  NAND2_X1 U8114 ( .A1(n13992), .A2(n6695), .ZN(n7297) );
  AND2_X1 U8115 ( .A1(n7298), .A2(n6695), .ZN(n7294) );
  INV_X1 U8116 ( .A(n7408), .ZN(n13992) );
  OR2_X1 U8117 ( .A1(n14053), .A2(n14054), .ZN(n14055) );
  OR2_X1 U8118 ( .A1(n14081), .A2(n14082), .ZN(n14079) );
  AOI21_X1 U8119 ( .B1(n7281), .B2(n7279), .A(n6755), .ZN(n7278) );
  INV_X1 U8120 ( .A(n6701), .ZN(n7279) );
  NAND2_X1 U8121 ( .A1(n9328), .A2(n9327), .ZN(n11879) );
  NAND2_X1 U8122 ( .A1(n9203), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9221) );
  NAND2_X1 U8123 ( .A1(n9180), .A2(n9179), .ZN(n10947) );
  NOR2_X1 U8124 ( .A1(n15332), .A2(n9794), .ZN(n7398) );
  INV_X1 U8125 ( .A(n11296), .ZN(n7050) );
  AND2_X1 U8126 ( .A1(n15300), .A2(n11474), .ZN(n15275) );
  AND2_X1 U8127 ( .A1(n9378), .A2(n9377), .ZN(n15008) );
  OR2_X1 U8128 ( .A1(n11062), .A2(n10693), .ZN(n15340) );
  AND2_X1 U8129 ( .A1(n10021), .A2(n10063), .ZN(n9708) );
  INV_X1 U8130 ( .A(n7258), .ZN(n9082) );
  INV_X1 U8131 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n9069) );
  INV_X1 U8132 ( .A(n14190), .ZN(n6856) );
  NOR2_X1 U8133 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), .ZN(
        n6855) );
  OR2_X1 U8134 ( .A1(n9675), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n9676) );
  CLKBUF_X1 U8135 ( .A(n9233), .Z(n9234) );
  AND2_X1 U8136 ( .A1(n15042), .A2(n15043), .ZN(n12967) );
  INV_X1 U8137 ( .A(n10615), .ZN(n6866) );
  INV_X1 U8138 ( .A(n12721), .ZN(n6867) );
  NAND2_X1 U8139 ( .A1(n7365), .A2(n7364), .ZN(n10622) );
  NAND2_X1 U8140 ( .A1(n13059), .A2(n14378), .ZN(n7365) );
  NAND2_X1 U8141 ( .A1(n13070), .A2(n12530), .ZN(n7364) );
  AND2_X1 U8142 ( .A1(n13066), .A2(n13065), .ZN(n14245) );
  AND2_X1 U8143 ( .A1(n14244), .A2(n13054), .ZN(n14274) );
  NAND2_X1 U8144 ( .A1(n7351), .A2(n7349), .ZN(n14214) );
  AOI21_X1 U8145 ( .B1(n7352), .B2(n7355), .A(n7350), .ZN(n7349) );
  INV_X1 U8146 ( .A(n14302), .ZN(n7350) );
  NOR2_X1 U8147 ( .A1(n12875), .A2(n12874), .ZN(n7598) );
  AOI21_X1 U8148 ( .B1(n12240), .B2(P1_REG1_REG_13__SCAN_IN), .A(n11732), .ZN(
        n14446) );
  NAND2_X1 U8149 ( .A1(n14824), .A2(n7038), .ZN(n7037) );
  INV_X1 U8150 ( .A(n7039), .ZN(n7038) );
  OR2_X1 U8151 ( .A1(n14508), .A2(n14517), .ZN(n14509) );
  NAND2_X1 U8152 ( .A1(n12905), .A2(n7225), .ZN(n14547) );
  NOR2_X1 U8153 ( .A1(n14550), .A2(n7226), .ZN(n7225) );
  INV_X1 U8154 ( .A(n12904), .ZN(n7226) );
  INV_X1 U8155 ( .A(n14533), .ZN(n14531) );
  NAND2_X1 U8156 ( .A1(n14563), .A2(n14569), .ZN(n12905) );
  AND2_X1 U8157 ( .A1(n14567), .A2(n12930), .ZN(n14544) );
  OR2_X1 U8158 ( .A1(n14566), .A2(n14569), .ZN(n14567) );
  AOI21_X1 U8159 ( .B1(n12925), .B2(n6696), .A(n6973), .ZN(n6972) );
  NAND2_X1 U8160 ( .A1(n6974), .A2(n14587), .ZN(n6973) );
  NAND2_X1 U8161 ( .A1(n6696), .A2(n6975), .ZN(n6974) );
  NAND2_X1 U8162 ( .A1(n12900), .A2(n12697), .ZN(n14639) );
  INV_X1 U8163 ( .A(n6860), .ZN(n12900) );
  NAND2_X1 U8164 ( .A1(n14694), .A2(n12895), .ZN(n14678) );
  OR2_X1 U8165 ( .A1(n12452), .A2(n12451), .ZN(n12632) );
  NAND2_X1 U8166 ( .A1(n12894), .A2(n7209), .ZN(n14694) );
  NOR2_X1 U8167 ( .A1(n14697), .A2(n7210), .ZN(n7209) );
  INV_X1 U8168 ( .A(n12893), .ZN(n7210) );
  OR2_X1 U8169 ( .A1(n14810), .A2(n15040), .ZN(n12893) );
  AOI21_X1 U8170 ( .B1(n12914), .B2(n12917), .A(n6988), .ZN(n6985) );
  OR2_X1 U8171 ( .A1(n12245), .A2(n12244), .ZN(n12309) );
  AOI21_X1 U8172 ( .B1(n6980), .B2(n6671), .A(n12849), .ZN(n6978) );
  INV_X1 U8173 ( .A(n6980), .ZN(n6979) );
  INV_X1 U8174 ( .A(n14370), .ZN(n12082) );
  INV_X1 U8175 ( .A(n14371), .ZN(n12123) );
  NAND2_X1 U8176 ( .A1(n11421), .A2(n11319), .ZN(n7613) );
  MUX2_X1 U8177 ( .A(n7593), .B(n14879), .S(n12738), .Z(n11786) );
  OR2_X1 U8178 ( .A1(n14734), .A2(n13111), .ZN(n6883) );
  NAND2_X1 U8179 ( .A1(n12242), .A2(n12241), .ZN(n12957) );
  AOI21_X1 U8180 ( .B1(n10977), .B2(n12819), .A(n7177), .ZN(n7176) );
  OAI22_X1 U8181 ( .A1(n9106), .A2(n12721), .B1(n12738), .B2(n10825), .ZN(
        n6991) );
  INV_X1 U8182 ( .A(n14811), .ZN(n14781) );
  AND2_X1 U8183 ( .A1(n10500), .A2(n10499), .ZN(n11514) );
  AND2_X1 U8184 ( .A1(n10248), .A2(n12484), .ZN(n14771) );
  INV_X1 U8185 ( .A(n14618), .ZN(n14699) );
  XNOR2_X1 U8186 ( .A(n10208), .B(n10207), .ZN(n10247) );
  INV_X1 U8187 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n10207) );
  NAND2_X1 U8188 ( .A1(n10211), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10208) );
  INV_X1 U8189 ( .A(n10211), .ZN(n6863) );
  INV_X1 U8190 ( .A(n6960), .ZN(n6955) );
  NAND2_X1 U8191 ( .A1(n9355), .A2(n9369), .ZN(n9371) );
  OR2_X1 U8192 ( .A1(n10256), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n10257) );
  NAND2_X1 U8193 ( .A1(n7322), .A2(n9310), .ZN(n9330) );
  NAND2_X1 U8194 ( .A1(n9293), .A2(n7323), .ZN(n7322) );
  INV_X1 U8195 ( .A(n9197), .ZN(n7028) );
  NAND4_X1 U8196 ( .A1(n10133), .A2(n10146), .A3(n10117), .A4(n7593), .ZN(
        n10119) );
  NAND2_X1 U8197 ( .A1(n9181), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n6848) );
  XNOR2_X1 U8198 ( .A(n7907), .B(n7310), .ZN(n7909) );
  INV_X1 U8199 ( .A(n7906), .ZN(n7310) );
  XNOR2_X1 U8200 ( .A(n7863), .B(n8246), .ZN(n7903) );
  INV_X1 U8201 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14393) );
  XNOR2_X1 U8202 ( .A(n7913), .B(P1_ADDR_REG_5__SCAN_IN), .ZN(n7915) );
  NOR2_X1 U8203 ( .A1(n14892), .A2(n7920), .ZN(n7922) );
  NOR2_X1 U8204 ( .A1(n7011), .A2(P2_ADDR_REG_9__SCAN_IN), .ZN(n7008) );
  AOI22_X1 U8205 ( .A1(n13300), .A2(n13301), .B1(n13419), .B2(n13176), .ZN(
        n13214) );
  NAND2_X1 U8206 ( .A1(n8733), .A2(n8732), .ZN(n13180) );
  NAND2_X1 U8207 ( .A1(n8689), .A2(n8688), .ZN(n13470) );
  AND3_X1 U8208 ( .A1(n8526), .A2(n8525), .A3(n8524), .ZN(n15378) );
  NAND2_X1 U8209 ( .A1(n11718), .A2(n11717), .ZN(n12007) );
  OR2_X1 U8210 ( .A1(n8761), .A2(n10159), .ZN(n7120) );
  AND3_X1 U8211 ( .A1(n8658), .A2(n8657), .A3(n8656), .ZN(n13519) );
  NAND2_X1 U8212 ( .A1(n8665), .A2(n8664), .ZN(n13498) );
  OR2_X1 U8213 ( .A1(n11136), .A2(n8663), .ZN(n8665) );
  NAND2_X1 U8214 ( .A1(n11184), .A2(n11183), .ZN(n11711) );
  NAND2_X1 U8215 ( .A1(n7134), .A2(n7132), .ZN(n7131) );
  OR2_X1 U8216 ( .A1(n13267), .A2(n7136), .ZN(n7134) );
  NAND2_X1 U8217 ( .A1(n13267), .A2(n7133), .ZN(n7132) );
  NAND2_X1 U8218 ( .A1(n13267), .A2(n13163), .ZN(n7135) );
  NAND2_X1 U8219 ( .A1(n8700), .A2(n8699), .ZN(n13272) );
  NAND2_X1 U8220 ( .A1(n13277), .A2(n13276), .ZN(n13275) );
  XNOR2_X1 U8221 ( .A(n13195), .B(n13193), .ZN(n13283) );
  NAND2_X1 U8222 ( .A1(n10554), .A2(n13538), .ZN(n15377) );
  INV_X1 U8223 ( .A(n11780), .ZN(n11714) );
  XNOR2_X1 U8224 ( .A(n7731), .B(n11906), .ZN(n11895) );
  XNOR2_X1 U8225 ( .A(n6858), .B(n10253), .ZN(n13332) );
  NOR2_X1 U8226 ( .A1(n13385), .A2(n7741), .ZN(n13388) );
  OAI211_X1 U8227 ( .C1(n14930), .C2(n15516), .A(n14929), .B(n7171), .ZN(n7170) );
  NOR2_X1 U8228 ( .A1(n7173), .A2(n7172), .ZN(n7171) );
  OAI21_X1 U8229 ( .B1(n13385), .B2(n7163), .A(n7162), .ZN(n14921) );
  NAND2_X1 U8230 ( .A1(n7164), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7163) );
  INV_X1 U8231 ( .A(n14922), .ZN(n7164) );
  OR2_X1 U8232 ( .A1(n7850), .A2(n8986), .ZN(n15530) );
  INV_X1 U8233 ( .A(n8989), .ZN(n7118) );
  NAND2_X1 U8234 ( .A1(n8763), .A2(n8762), .ZN(n13128) );
  OR2_X1 U8235 ( .A1(n13126), .A2(n13125), .ZN(n6839) );
  NOR2_X1 U8236 ( .A1(n7634), .A2(n9045), .ZN(n9046) );
  CLKBUF_X1 U8237 ( .A(n13545), .Z(n13610) );
  NAND2_X1 U8238 ( .A1(n8624), .A2(n8623), .ZN(n13544) );
  OR2_X1 U8239 ( .A1(n10542), .A2(n8663), .ZN(n8624) );
  NAND2_X1 U8240 ( .A1(n10553), .A2(n11310), .ZN(n13538) );
  INV_X1 U8241 ( .A(n13562), .ZN(n13543) );
  NAND2_X1 U8242 ( .A1(n8990), .A2(n13552), .ZN(n7116) );
  OR2_X1 U8243 ( .A1(n13420), .A2(n13410), .ZN(n7635) );
  NAND2_X1 U8244 ( .A1(n15607), .A2(n15561), .ZN(n13623) );
  INV_X1 U8245 ( .A(n13222), .ZN(n13410) );
  INV_X1 U8246 ( .A(n13180), .ZN(n13633) );
  NAND2_X1 U8247 ( .A1(n7549), .A2(n7547), .ZN(n11671) );
  AND2_X1 U8248 ( .A1(n11456), .A2(n6685), .ZN(n7547) );
  NOR2_X1 U8249 ( .A1(n13749), .A2(n6894), .ZN(n6893) );
  INV_X1 U8250 ( .A(n10738), .ZN(n6894) );
  AND2_X1 U8251 ( .A1(n6898), .A2(n6908), .ZN(n6896) );
  NAND2_X1 U8252 ( .A1(n6900), .A2(n6904), .ZN(n6899) );
  NAND2_X1 U8253 ( .A1(n13772), .A2(n13767), .ZN(n6904) );
  INV_X1 U8254 ( .A(n11247), .ZN(n11215) );
  AND2_X1 U8255 ( .A1(n10729), .A2(n10728), .ZN(n10915) );
  OR2_X1 U8256 ( .A1(n13722), .A2(n13721), .ZN(n13723) );
  INV_X1 U8257 ( .A(n14052), .ZN(n14151) );
  NAND2_X1 U8258 ( .A1(n10905), .A2(n10906), .ZN(n10904) );
  OR2_X1 U8259 ( .A1(n12659), .A2(n9523), .ZN(n9441) );
  INV_X1 U8260 ( .A(n15008), .ZN(n12363) );
  NAND2_X1 U8261 ( .A1(n10685), .A2(n14086), .ZN(n13857) );
  NAND2_X1 U8262 ( .A1(n9622), .A2(n9621), .ZN(n13864) );
  INV_X1 U8263 ( .A(n9895), .ZN(n13866) );
  INV_X1 U8264 ( .A(n11589), .ZN(n13878) );
  INV_X1 U8265 ( .A(n11587), .ZN(n13880) );
  OR2_X1 U8266 ( .A1(n6666), .A2(n9071), .ZN(n9074) );
  OR2_X1 U8267 ( .A1(n9928), .A2(n10075), .ZN(n9073) );
  NAND2_X1 U8268 ( .A1(n9599), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n9098) );
  AOI21_X1 U8269 ( .B1(n7248), .B2(n14065), .A(n9674), .ZN(n14108) );
  INV_X1 U8270 ( .A(n9673), .ZN(n9674) );
  AOI22_X1 U8271 ( .A1(n13863), .A2(n13851), .B1(n13913), .B2(n13861), .ZN(
        n9673) );
  OR2_X1 U8272 ( .A1(n11555), .A2(n9523), .ZN(n9525) );
  INV_X1 U8273 ( .A(n15280), .ZN(n14099) );
  NAND2_X1 U8274 ( .A1(n9706), .A2(n9705), .ZN(n15287) );
  INV_X1 U8275 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n11113) );
  NAND2_X1 U8276 ( .A1(n11381), .A2(n11380), .ZN(n12577) );
  INV_X1 U8277 ( .A(n7379), .ZN(n7378) );
  OAI21_X1 U8278 ( .B1(n6672), .B2(n6680), .A(n6785), .ZN(n7379) );
  NOR2_X1 U8279 ( .A1(n7369), .A2(n15062), .ZN(n7367) );
  NOR2_X1 U8280 ( .A1(n7372), .A2(n7370), .ZN(n7369) );
  INV_X1 U8281 ( .A(n7373), .ZN(n7370) );
  NAND2_X1 U8282 ( .A1(n7373), .A2(n7374), .ZN(n7371) );
  INV_X1 U8283 ( .A(n13091), .ZN(n7374) );
  INV_X1 U8284 ( .A(n14372), .ZN(n12080) );
  INV_X1 U8285 ( .A(n14368), .ZN(n12424) );
  NOR2_X1 U8286 ( .A1(n12422), .A2(n7363), .ZN(n7362) );
  INV_X1 U8287 ( .A(n12416), .ZN(n7363) );
  NAND2_X1 U8288 ( .A1(n15063), .A2(n12416), .ZN(n12421) );
  INV_X1 U8289 ( .A(n14364), .ZN(n15040) );
  OR2_X1 U8290 ( .A1(n12707), .A2(n12721), .ZN(n12710) );
  OR2_X1 U8291 ( .A1(n10822), .A2(n10821), .ZN(n7361) );
  AND2_X1 U8292 ( .A1(n10641), .A2(n12484), .ZN(n14620) );
  OR2_X1 U8293 ( .A1(n14479), .A2(n15124), .ZN(n6820) );
  AOI21_X1 U8294 ( .B1(n14481), .B2(n14482), .A(n14480), .ZN(n6819) );
  NAND2_X1 U8295 ( .A1(n6976), .A2(n13098), .ZN(n14737) );
  NAND2_X1 U8296 ( .A1(n12938), .A2(n12939), .ZN(n6976) );
  NAND2_X1 U8297 ( .A1(n14676), .A2(n12919), .ZN(n7606) );
  NAND2_X1 U8298 ( .A1(n12880), .A2(n11513), .ZN(n14706) );
  INV_X1 U8299 ( .A(n14508), .ZN(n14830) );
  NAND2_X1 U8300 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), 
        .ZN(n7596) );
  NOR2_X1 U8301 ( .A1(n10487), .A2(n7595), .ZN(n7594) );
  NOR2_X1 U8302 ( .A1(n10761), .A2(n10495), .ZN(n7597) );
  INV_X1 U8303 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n11112) );
  XNOR2_X1 U8304 ( .A(n7909), .B(n7309), .ZN(n15623) );
  NAND2_X1 U8305 ( .A1(n14888), .A2(n7303), .ZN(n15620) );
  OAI21_X1 U8306 ( .B1(n14889), .B2(n14890), .A(n7304), .ZN(n7303) );
  INV_X1 U8307 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n7304) );
  NOR2_X1 U8308 ( .A1(n14893), .A2(n14894), .ZN(n14892) );
  OR2_X1 U8309 ( .A1(n14901), .A2(n14900), .ZN(n7006) );
  NAND2_X1 U8310 ( .A1(n7004), .A2(n7001), .ZN(n7003) );
  NOR2_X1 U8311 ( .A1(n14915), .A2(n7953), .ZN(n7001) );
  AND2_X1 U8312 ( .A1(n7952), .A2(n7953), .ZN(n14882) );
  AND2_X1 U8313 ( .A1(n7003), .A2(n7002), .ZN(n7308) );
  INV_X1 U8314 ( .A(P2_ADDR_REG_18__SCAN_IN), .ZN(n7002) );
  INV_X1 U8315 ( .A(n7419), .ZN(n7416) );
  AND3_X1 U8316 ( .A1(n7565), .A2(n7566), .A3(n12554), .ZN(n7564) );
  OR2_X1 U8317 ( .A1(n7444), .A2(n7445), .ZN(n6774) );
  INV_X1 U8318 ( .A(n9803), .ZN(n9806) );
  INV_X1 U8319 ( .A(n9813), .ZN(n7421) );
  NAND2_X1 U8320 ( .A1(n7588), .A2(n12578), .ZN(n7587) );
  OR2_X1 U8321 ( .A1(n12578), .A2(n7588), .ZN(n7586) );
  NAND2_X1 U8322 ( .A1(n12590), .A2(n7562), .ZN(n7561) );
  NAND2_X1 U8323 ( .A1(n7502), .A2(n7501), .ZN(n7500) );
  INV_X1 U8324 ( .A(n9825), .ZN(n7501) );
  INV_X1 U8325 ( .A(n9837), .ZN(n7481) );
  NOR2_X1 U8326 ( .A1(n7481), .A2(n7480), .ZN(n7477) );
  NAND2_X1 U8327 ( .A1(n12612), .A2(n7571), .ZN(n7568) );
  NOR2_X1 U8328 ( .A1(n6730), .A2(n7570), .ZN(n7569) );
  NOR2_X1 U8329 ( .A1(n7571), .A2(n12612), .ZN(n7570) );
  AND2_X1 U8330 ( .A1(n7474), .A2(n9864), .ZN(n7473) );
  NAND2_X1 U8331 ( .A1(n7475), .A2(n7478), .ZN(n7474) );
  AND2_X1 U8332 ( .A1(n7490), .A2(n9875), .ZN(n7489) );
  NAND2_X1 U8333 ( .A1(n7494), .A2(n7493), .ZN(n7490) );
  AND2_X1 U8334 ( .A1(n9872), .A2(n7495), .ZN(n7494) );
  INV_X1 U8335 ( .A(n9874), .ZN(n7495) );
  NOR2_X1 U8336 ( .A1(n7492), .A2(n9875), .ZN(n7491) );
  NAND2_X1 U8337 ( .A1(n7486), .A2(n7488), .ZN(n7484) );
  INV_X1 U8338 ( .A(n7489), .ZN(n7488) );
  NAND2_X1 U8339 ( .A1(n7491), .A2(n7494), .ZN(n7483) );
  CLKBUF_X1 U8340 ( .A(n9764), .Z(n9826) );
  NAND2_X1 U8341 ( .A1(n9883), .A2(n7455), .ZN(n7454) );
  INV_X1 U8342 ( .A(n9884), .ZN(n7455) );
  AOI21_X1 U8343 ( .B1(n12696), .B2(n12697), .A(n12695), .ZN(n12698) );
  NOR2_X1 U8344 ( .A1(n7450), .A2(n7448), .ZN(n7447) );
  AOI22_X1 U8345 ( .A1(n7450), .A2(n7452), .B1(n7448), .B2(n7456), .ZN(n7446)
         );
  INV_X1 U8346 ( .A(n7573), .ZN(n7572) );
  OAI21_X1 U8347 ( .B1(n7576), .B2(n7574), .A(n12742), .ZN(n7573) );
  INV_X1 U8348 ( .A(n12745), .ZN(n7574) );
  OAI22_X1 U8349 ( .A1(n13990), .A2(n9908), .B1(n13788), .B2(n10005), .ZN(
        n9890) );
  OAI21_X1 U8350 ( .B1(n8914), .B2(n6837), .A(n6750), .ZN(n8918) );
  NAND2_X1 U8351 ( .A1(n6754), .A2(n7091), .ZN(n6837) );
  INV_X1 U8352 ( .A(n12796), .ZN(n7591) );
  INV_X1 U8353 ( .A(n7556), .ZN(n7554) );
  INV_X1 U8354 ( .A(n9432), .ZN(n7317) );
  NOR2_X1 U8355 ( .A1(n9470), .A2(SI_18_), .ZN(n9474) );
  AOI21_X1 U8356 ( .B1(n7772), .B2(n7519), .A(n15408), .ZN(n7517) );
  NOR2_X1 U8357 ( .A1(n7747), .A2(P3_IR_REG_26__SCAN_IN), .ZN(n7748) );
  AOI21_X1 U8358 ( .B1(n8673), .B2(n8342), .A(n7236), .ZN(n7235) );
  INV_X1 U8359 ( .A(n8686), .ZN(n7236) );
  INV_X1 U8360 ( .A(n8342), .ZN(n7233) );
  AND2_X1 U8361 ( .A1(n9762), .A2(n11556), .ZN(n9764) );
  NAND2_X1 U8362 ( .A1(n9953), .A2(n10006), .ZN(n9959) );
  INV_X1 U8363 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n9238) );
  INV_X1 U8364 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n9059) );
  INV_X1 U8365 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n9061) );
  NOR2_X1 U8366 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_4__SCAN_IN), .ZN(
        n9062) );
  INV_X1 U8367 ( .A(n12921), .ZN(n7605) );
  NOR2_X1 U8368 ( .A1(n14751), .A2(n7046), .ZN(n7045) );
  INV_X1 U8369 ( .A(n7047), .ZN(n7046) );
  NAND2_X1 U8370 ( .A1(n9558), .A2(n12890), .ZN(n9559) );
  INV_X1 U8371 ( .A(n6953), .ZN(n6952) );
  OAI21_X1 U8372 ( .B1(n9386), .B2(n6954), .A(n9406), .ZN(n6953) );
  INV_X1 U8373 ( .A(n9388), .ZN(n6954) );
  NAND2_X1 U8374 ( .A1(n9253), .A2(SI_9_), .ZN(n9273) );
  NAND2_X1 U8375 ( .A1(n7390), .A2(n7388), .ZN(n7016) );
  NAND2_X1 U8376 ( .A1(n9143), .A2(SI_2_), .ZN(n7017) );
  NAND2_X1 U8377 ( .A1(n9181), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n6830) );
  NOR2_X1 U8378 ( .A1(n8795), .A2(n8774), .ZN(n7461) );
  INV_X1 U8379 ( .A(n8931), .ZN(n7462) );
  NOR2_X1 U8380 ( .A1(n13626), .A2(n7221), .ZN(n8934) );
  OR2_X1 U8381 ( .A1(n10572), .A2(n7770), .ZN(n7771) );
  OAI21_X1 U8382 ( .B1(n10584), .B2(n7159), .A(n7157), .ZN(n7161) );
  AOI21_X1 U8383 ( .B1(n7720), .B2(n7158), .A(n15405), .ZN(n7157) );
  AND2_X1 U8384 ( .A1(n10583), .A2(n7720), .ZN(n15404) );
  AND2_X1 U8385 ( .A1(n7521), .A2(n7520), .ZN(n7774) );
  NAND2_X1 U8386 ( .A1(n15417), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7520) );
  AND2_X1 U8387 ( .A1(n7161), .A2(n7160), .ZN(n7722) );
  NAND2_X1 U8388 ( .A1(n15417), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7160) );
  INV_X1 U8389 ( .A(n15481), .ZN(n6939) );
  XNOR2_X1 U8390 ( .A(n7841), .B(n10540), .ZN(n14927) );
  NOR2_X1 U8391 ( .A1(n13392), .A2(n7839), .ZN(n7841) );
  OR2_X1 U8392 ( .A1(n13222), .A2(n13420), .ZN(n8922) );
  OR2_X1 U8393 ( .A1(n8722), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8734) );
  NAND2_X1 U8394 ( .A1(n13322), .A2(n13470), .ZN(n7101) );
  OR2_X1 U8395 ( .A1(n13288), .A2(n13197), .ZN(n8907) );
  OR2_X1 U8396 ( .A1(n13498), .A2(n13506), .ZN(n8903) );
  NAND2_X1 U8397 ( .A1(n7430), .A2(n8874), .ZN(n7429) );
  INV_X1 U8398 ( .A(n12370), .ZN(n7430) );
  INV_X1 U8399 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n8486) );
  NOR2_X1 U8400 ( .A1(n8959), .A2(n11544), .ZN(n8961) );
  AND2_X1 U8401 ( .A1(n8809), .A2(n8812), .ZN(n8806) );
  NAND2_X1 U8402 ( .A1(n13633), .A2(n13218), .ZN(n7085) );
  INV_X1 U8403 ( .A(n8352), .ZN(n7230) );
  INV_X1 U8404 ( .A(n8346), .ZN(n7246) );
  INV_X1 U8405 ( .A(n7217), .ZN(n7216) );
  OAI21_X1 U8406 ( .B1(n8439), .B2(n7218), .A(n8454), .ZN(n7217) );
  INV_X1 U8407 ( .A(n8306), .ZN(n7218) );
  OR2_X1 U8408 ( .A1(n9239), .A2(n9238), .ZN(n9261) );
  NOR2_X1 U8409 ( .A1(n6720), .A2(n7438), .ZN(n7432) );
  NOR2_X1 U8410 ( .A1(n7439), .A2(n9905), .ZN(n7438) );
  NAND2_X1 U8411 ( .A1(n7436), .A2(n7435), .ZN(n7434) );
  NAND2_X1 U8412 ( .A1(n9956), .A2(n6682), .ZN(n7435) );
  NAND2_X1 U8413 ( .A1(n13990), .A2(n7054), .ZN(n7053) );
  INV_X1 U8414 ( .A(n7055), .ZN(n7054) );
  NAND2_X1 U8415 ( .A1(n14008), .A2(n7056), .ZN(n7055) );
  INV_X1 U8416 ( .A(n9427), .ZN(n7262) );
  NAND2_X1 U8417 ( .A1(n7261), .A2(n9426), .ZN(n7260) );
  NAND2_X1 U8418 ( .A1(n6749), .A2(n15014), .ZN(n7060) );
  OR2_X1 U8419 ( .A1(n9261), .A2(n11275), .ZN(n9282) );
  AND2_X1 U8420 ( .A1(n11556), .A2(n9664), .ZN(n9713) );
  NAND2_X1 U8421 ( .A1(n7058), .A2(n7057), .ZN(n13932) );
  INV_X1 U8422 ( .A(n14110), .ZN(n7057) );
  INV_X1 U8423 ( .A(n12540), .ZN(n10620) );
  AOI21_X1 U8424 ( .B1(n13025), .B2(n7354), .A(n7353), .ZN(n7352) );
  INV_X1 U8425 ( .A(n13009), .ZN(n7354) );
  INV_X1 U8426 ( .A(n13025), .ZN(n7355) );
  NAND2_X1 U8427 ( .A1(n12826), .A2(n12824), .ZN(n7584) );
  NAND2_X1 U8428 ( .A1(n7622), .A2(n12951), .ZN(n10989) );
  INV_X1 U8429 ( .A(n10989), .ZN(n11689) );
  NOR2_X1 U8430 ( .A1(n14757), .A2(n13039), .ZN(n7047) );
  INV_X1 U8431 ( .A(n12700), .ZN(n12506) );
  OR2_X1 U8432 ( .A1(n12668), .A2(n12652), .ZN(n12700) );
  NOR2_X1 U8433 ( .A1(n14807), .A2(n14810), .ZN(n7034) );
  INV_X1 U8434 ( .A(n11971), .ZN(n7609) );
  AND2_X1 U8435 ( .A1(n6673), .A2(n7041), .ZN(n7040) );
  NOR2_X1 U8436 ( .A1(n12589), .A2(n12580), .ZN(n7043) );
  NOR2_X1 U8437 ( .A1(n11386), .A2(n11385), .ZN(n11690) );
  AND2_X1 U8438 ( .A1(n12500), .A2(n12478), .ZN(n12540) );
  XNOR2_X1 U8439 ( .A(n14376), .B(n10988), .ZN(n7175) );
  INV_X1 U8440 ( .A(n12486), .ZN(n12500) );
  AOI21_X1 U8441 ( .B1(n6675), .B2(n14642), .A(n6741), .ZN(n7219) );
  AND2_X1 U8442 ( .A1(n12318), .A2(n15074), .ZN(n12462) );
  INV_X1 U8443 ( .A(n11435), .ZN(n7033) );
  NAND2_X1 U8444 ( .A1(n6878), .A2(n6799), .ZN(n9945) );
  INV_X1 U8445 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n10027) );
  NOR2_X1 U8446 ( .A1(n10119), .A2(n7238), .ZN(n7237) );
  NAND2_X1 U8447 ( .A1(n10039), .A2(n10121), .ZN(n7238) );
  INV_X1 U8448 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n10039) );
  NAND2_X1 U8449 ( .A1(n9559), .A2(n7337), .ZN(n7336) );
  INV_X1 U8450 ( .A(n9560), .ZN(n7337) );
  INV_X1 U8451 ( .A(n9558), .ZN(n6829) );
  INV_X1 U8452 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n10044) );
  AOI21_X1 U8453 ( .B1(n7314), .B2(n6676), .A(n6784), .ZN(n7313) );
  AOI21_X1 U8454 ( .B1(n7321), .B2(n9329), .A(n6744), .ZN(n7320) );
  NOR2_X1 U8455 ( .A1(n9311), .A2(n7324), .ZN(n7323) );
  INV_X1 U8456 ( .A(n9292), .ZN(n7324) );
  OAI21_X1 U8457 ( .B1(n9275), .B2(SI_10_), .A(n9292), .ZN(n9289) );
  OAI21_X1 U8458 ( .B1(n9253), .B2(SI_9_), .A(n9273), .ZN(n9270) );
  NAND2_X1 U8459 ( .A1(n6670), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n6852) );
  INV_X1 U8460 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n8246) );
  OAI21_X1 U8461 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n7878), .A(n7877), .ZN(
        n7879) );
  NAND2_X1 U8462 ( .A1(n12391), .A2(n12390), .ZN(n7146) );
  NAND2_X1 U8463 ( .A1(n13163), .A2(n7138), .ZN(n7133) );
  INV_X1 U8464 ( .A(n8640), .ZN(n8372) );
  INV_X1 U8465 ( .A(n7144), .ZN(n7143) );
  OAI21_X1 U8466 ( .B1(n12227), .B2(n12398), .A(n12393), .ZN(n7144) );
  NAND2_X1 U8467 ( .A1(n8367), .A2(n8366), .ZN(n8572) );
  INV_X1 U8468 ( .A(n8559), .ZN(n8367) );
  NAND2_X1 U8469 ( .A1(n12228), .A2(n12227), .ZN(n12391) );
  OR2_X1 U8470 ( .A1(n12228), .A2(n12227), .ZN(n12392) );
  OR2_X1 U8471 ( .A1(n8528), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8540) );
  NAND2_X1 U8472 ( .A1(n11713), .A2(n10708), .ZN(n6814) );
  INV_X1 U8473 ( .A(n8613), .ZN(n8371) );
  NAND2_X1 U8474 ( .A1(n8447), .A2(n8092), .ZN(n8459) );
  AND4_X1 U8475 ( .A1(n8519), .A2(n8518), .A3(n8517), .A4(n8516), .ZN(n12223)
         );
  AND4_X1 U8476 ( .A1(n8492), .A2(n8491), .A3(n8490), .A4(n8489), .ZN(n12013)
         );
  OR2_X1 U8477 ( .A1(n12033), .A2(n7663), .ZN(n7745) );
  AND2_X1 U8478 ( .A1(n10602), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10605) );
  NOR2_X1 U8479 ( .A1(n10598), .A2(n11665), .ZN(n10597) );
  NAND2_X1 U8480 ( .A1(n7505), .A2(n7769), .ZN(n10573) );
  NAND2_X1 U8481 ( .A1(n7768), .A2(n7767), .ZN(n7505) );
  XNOR2_X1 U8482 ( .A(n7771), .B(n10594), .ZN(n10587) );
  NAND2_X1 U8483 ( .A1(n10587), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n10586) );
  NAND2_X1 U8484 ( .A1(n10584), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n10583) );
  NOR2_X1 U8485 ( .A1(n15426), .A2(n15596), .ZN(n15425) );
  NOR2_X1 U8486 ( .A1(n7726), .A2(n15454), .ZN(n15475) );
  NOR2_X1 U8487 ( .A1(n15475), .A2(n15474), .ZN(n15473) );
  AOI21_X1 U8488 ( .B1(n15459), .B2(n15458), .A(n7819), .ZN(n15478) );
  NAND2_X1 U8489 ( .A1(n7167), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7166) );
  INV_X1 U8490 ( .A(n11155), .ZN(n7167) );
  NOR2_X1 U8491 ( .A1(n11045), .A2(n11533), .ZN(n11044) );
  NAND2_X1 U8492 ( .A1(n7511), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7510) );
  NAND2_X1 U8493 ( .A1(n7784), .A2(n7511), .ZN(n7509) );
  INV_X1 U8494 ( .A(n15497), .ZN(n7511) );
  NOR2_X1 U8495 ( .A1(n11902), .A2(n14958), .ZN(n11901) );
  NOR2_X1 U8496 ( .A1(n15525), .A2(n15526), .ZN(n15524) );
  NOR2_X1 U8497 ( .A1(n13356), .A2(n13357), .ZN(n13355) );
  NOR2_X1 U8498 ( .A1(n6933), .A2(n13361), .ZN(n7787) );
  OAI21_X1 U8499 ( .B1(n13348), .B2(n7515), .A(n6932), .ZN(n13375) );
  NAND2_X1 U8500 ( .A1(n7516), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7515) );
  NAND2_X1 U8501 ( .A1(n7787), .A2(n7516), .ZN(n6932) );
  INV_X1 U8502 ( .A(n13376), .ZN(n7516) );
  NOR2_X1 U8503 ( .A1(n13375), .A2(n6931), .ZN(n7788) );
  NOR2_X1 U8504 ( .A1(n8597), .A2(n13621), .ZN(n6931) );
  INV_X1 U8505 ( .A(n14931), .ZN(n7173) );
  NOR2_X1 U8506 ( .A1(n14932), .A2(P3_STATE_REG_SCAN_IN), .ZN(n7172) );
  NOR2_X1 U8507 ( .A1(n13417), .A2(n7084), .ZN(n7083) );
  INV_X1 U8508 ( .A(n7087), .ZN(n7084) );
  NAND2_X1 U8509 ( .A1(n13306), .A2(n13238), .ZN(n7087) );
  AOI21_X1 U8510 ( .B1(n7467), .B2(n7469), .A(n7466), .ZN(n7465) );
  INV_X1 U8511 ( .A(n8916), .ZN(n7466) );
  INV_X1 U8512 ( .A(n13417), .ZN(n13421) );
  AOI21_X1 U8513 ( .B1(n7092), .B2(n7095), .A(n7091), .ZN(n7090) );
  AOI21_X1 U8514 ( .B1(n7094), .B2(n7093), .A(n13442), .ZN(n7092) );
  INV_X1 U8515 ( .A(n8701), .ZN(n8374) );
  OR2_X1 U8516 ( .A1(n8690), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8701) );
  OR2_X1 U8517 ( .A1(n8654), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8666) );
  NAND2_X1 U8518 ( .A1(n8373), .A2(n8049), .ZN(n8677) );
  INV_X1 U8519 ( .A(n8666), .ZN(n8373) );
  OAI22_X1 U8520 ( .A1(n13529), .A2(n7063), .B1(n6738), .B2(n7062), .ZN(n13492) );
  INV_X1 U8521 ( .A(n7074), .ZN(n7062) );
  NAND2_X1 U8522 ( .A1(n7066), .A2(n7074), .ZN(n7063) );
  NAND2_X1 U8523 ( .A1(n7077), .A2(n7076), .ZN(n12130) );
  AOI21_X1 U8524 ( .B1(n7079), .B2(n7081), .A(n6777), .ZN(n7076) );
  NAND2_X1 U8525 ( .A1(n7078), .A2(n8971), .ZN(n12035) );
  NAND2_X1 U8526 ( .A1(n12046), .A2(n8970), .ZN(n7078) );
  INV_X1 U8527 ( .A(n14953), .ZN(n12054) );
  AND3_X1 U8528 ( .A1(n8512), .A2(n8511), .A3(n8510), .ZN(n11531) );
  NAND2_X1 U8529 ( .A1(n7109), .A2(n6716), .ZN(n11527) );
  OR2_X1 U8530 ( .A1(n8459), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8469) );
  AND2_X1 U8531 ( .A1(n11763), .A2(n8822), .ZN(n11544) );
  INV_X1 U8532 ( .A(n13520), .ZN(n13533) );
  AND2_X1 U8533 ( .A1(n8813), .A2(n8817), .ZN(n11753) );
  INV_X1 U8534 ( .A(n8806), .ZN(n11303) );
  AND4_X1 U8535 ( .A1(n8426), .A2(n8425), .A3(n8424), .A4(n8423), .ZN(n11304)
         );
  NAND2_X1 U8536 ( .A1(n8804), .A2(n10708), .ZN(n10772) );
  NAND2_X1 U8537 ( .A1(n7086), .A2(n7082), .ZN(n9043) );
  AND2_X1 U8538 ( .A1(n13216), .A2(n7085), .ZN(n7082) );
  NAND2_X1 U8539 ( .A1(n8395), .A2(n8394), .ZN(n7222) );
  NAND2_X1 U8540 ( .A1(n8363), .A2(n8362), .ZN(n8773) );
  OR2_X1 U8541 ( .A1(n11037), .A2(n8663), .ZN(n8653) );
  NAND2_X1 U8542 ( .A1(n7227), .A2(n7228), .ZN(n8759) );
  AOI21_X1 U8543 ( .B1(n7229), .B2(n8351), .A(n6800), .ZN(n7228) );
  NAND2_X1 U8544 ( .A1(n6891), .A2(n6889), .ZN(n7751) );
  NAND2_X1 U8545 ( .A1(n6890), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n6889) );
  AND2_X1 U8546 ( .A1(n7653), .A2(n7664), .ZN(n7141) );
  NAND2_X1 U8547 ( .A1(n8345), .A2(n8344), .ZN(n8698) );
  NAND2_X1 U8548 ( .A1(n8651), .A2(n8339), .ZN(n8660) );
  NAND2_X1 U8549 ( .A1(n7199), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n8339) );
  NAND2_X1 U8550 ( .A1(n8635), .A2(n8338), .ZN(n7199) );
  NAND2_X1 U8551 ( .A1(n8660), .A2(n8659), .ZN(n8662) );
  NAND2_X1 U8552 ( .A1(n7201), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7200) );
  INV_X1 U8553 ( .A(n8338), .ZN(n7201) );
  NAND2_X1 U8554 ( .A1(n8635), .A2(n6790), .ZN(n7202) );
  NAND3_X1 U8555 ( .A1(n7198), .A2(n7197), .A3(n7202), .ZN(n8651) );
  AND2_X1 U8556 ( .A1(n7200), .A2(n12708), .ZN(n7197) );
  NAND2_X1 U8557 ( .A1(n8622), .A2(n8336), .ZN(n8633) );
  NAND2_X1 U8558 ( .A1(n7180), .A2(n7178), .ZN(n8608) );
  AOI21_X1 U8559 ( .B1(n7181), .B2(n7183), .A(n7179), .ZN(n7178) );
  INV_X1 U8560 ( .A(n8332), .ZN(n7179) );
  INV_X1 U8561 ( .A(P3_IR_REG_14__SCAN_IN), .ZN(n7678) );
  AND2_X1 U8562 ( .A1(n8328), .A2(n8327), .ZN(n8566) );
  AND2_X1 U8563 ( .A1(n7647), .A2(n7646), .ZN(n7496) );
  NAND2_X1 U8564 ( .A1(n8496), .A2(n8315), .ZN(n8507) );
  NAND2_X1 U8565 ( .A1(n8507), .A2(n8506), .ZN(n8509) );
  XNOR2_X1 U8566 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n8412) );
  NAND2_X1 U8567 ( .A1(n9093), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8411) );
  INV_X1 U8568 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9220) );
  OR2_X1 U8569 ( .A1(n9221), .A2(n9220), .ZN(n9239) );
  NOR2_X1 U8570 ( .A1(n13756), .A2(n7529), .ZN(n7528) );
  INV_X1 U8571 ( .A(n7531), .ZN(n7529) );
  NAND2_X1 U8572 ( .A1(n13704), .A2(n7532), .ZN(n7531) );
  INV_X1 U8573 ( .A(n13705), .ZN(n7532) );
  NAND2_X1 U8574 ( .A1(n13802), .A2(n7533), .ZN(n7530) );
  INV_X1 U8575 ( .A(n13772), .ZN(n6903) );
  INV_X1 U8576 ( .A(n6906), .ZN(n6905) );
  NOR2_X1 U8577 ( .A1(n6914), .A2(n6913), .ZN(n6912) );
  INV_X1 U8578 ( .A(n13692), .ZN(n6913) );
  OR2_X1 U8579 ( .A1(n9565), .A2(n13815), .ZN(n9577) );
  INV_X1 U8580 ( .A(n11204), .ZN(n7548) );
  NAND2_X1 U8581 ( .A1(n13802), .A2(n7526), .ZN(n6927) );
  NAND2_X1 U8582 ( .A1(n9318), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n9339) );
  INV_X1 U8583 ( .A(n9320), .ZN(n9318) );
  INV_X1 U8584 ( .A(n9443), .ZN(n9442) );
  INV_X1 U8585 ( .A(n13841), .ZN(n13852) );
  AND2_X1 U8586 ( .A1(n10018), .A2(n9757), .ZN(n10692) );
  AND4_X1 U8587 ( .A1(n9347), .A2(n9346), .A3(n9345), .A4(n9344), .ZN(n11589)
         );
  AND4_X1 U8588 ( .A1(n9326), .A2(n9325), .A3(n9324), .A4(n9323), .ZN(n11914)
         );
  AND4_X1 U8589 ( .A1(n9245), .A2(n9244), .A3(n9243), .A4(n9242), .ZN(n11198)
         );
  OR2_X1 U8590 ( .A1(n9131), .A2(n11472), .ZN(n9075) );
  NAND2_X1 U8591 ( .A1(n13918), .A2(n14104), .ZN(n13917) );
  INV_X1 U8592 ( .A(n9995), .ZN(n9654) );
  INV_X1 U8593 ( .A(n14106), .ZN(n9934) );
  AND2_X1 U8594 ( .A1(n9634), .A2(n9633), .ZN(n13934) );
  AND2_X1 U8595 ( .A1(n9614), .A2(n9598), .ZN(n13955) );
  NAND2_X1 U8596 ( .A1(n14008), .A2(n13832), .ZN(n7410) );
  NOR2_X1 U8597 ( .A1(n14036), .A2(n7053), .ZN(n13986) );
  NOR2_X1 U8598 ( .A1(n14036), .A2(n7055), .ZN(n14005) );
  NOR2_X1 U8599 ( .A1(n14000), .A2(n7413), .ZN(n7412) );
  NAND2_X1 U8600 ( .A1(n9527), .A2(n9526), .ZN(n9543) );
  INV_X1 U8601 ( .A(n9529), .ZN(n9527) );
  OR2_X1 U8602 ( .A1(n9485), .A2(n9484), .ZN(n9529) );
  NAND2_X1 U8603 ( .A1(n7270), .A2(n7274), .ZN(n7269) );
  AOI21_X1 U8604 ( .B1(n14082), .B2(n7404), .A(n7403), .ZN(n7402) );
  NOR2_X1 U8605 ( .A1(n14072), .A2(n13842), .ZN(n7403) );
  AND2_X1 U8606 ( .A1(n14072), .A2(n14090), .ZN(n14067) );
  INV_X1 U8607 ( .A(n9984), .ZN(n12281) );
  AOI21_X1 U8608 ( .B1(n6752), .B2(n7278), .A(n6687), .ZN(n7276) );
  NAND2_X1 U8609 ( .A1(n7278), .A2(n6699), .ZN(n7277) );
  NAND2_X1 U8610 ( .A1(n9379), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n9418) );
  INV_X1 U8611 ( .A(n9381), .ZN(n9379) );
  NOR3_X1 U8612 ( .A1(n11885), .A2(n14991), .A3(n11888), .ZN(n14994) );
  OR2_X1 U8613 ( .A1(n9361), .A2(n12160), .ZN(n9381) );
  NOR2_X1 U8614 ( .A1(n11885), .A2(n11888), .ZN(n14996) );
  INV_X1 U8615 ( .A(n7394), .ZN(n7393) );
  AOI21_X1 U8616 ( .B1(n7392), .B2(n7394), .A(n6733), .ZN(n7391) );
  NOR2_X1 U8617 ( .A1(n9736), .A2(n7395), .ZN(n7394) );
  OR2_X1 U8618 ( .A1(n9299), .A2(n9298), .ZN(n9320) );
  XNOR2_X1 U8619 ( .A(n10723), .B(n11556), .ZN(n11641) );
  AOI21_X1 U8620 ( .B1(n11028), .B2(n7255), .A(n6743), .ZN(n7254) );
  NAND2_X1 U8621 ( .A1(n11024), .A2(n11265), .ZN(n11072) );
  NAND2_X1 U8622 ( .A1(n10942), .A2(n7400), .ZN(n7399) );
  NOR2_X1 U8623 ( .A1(n6709), .A2(n7020), .ZN(n7019) );
  INV_X1 U8624 ( .A(n9729), .ZN(n7400) );
  NAND2_X1 U8625 ( .A1(n9171), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9204) );
  NAND2_X1 U8626 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9173) );
  NAND2_X1 U8627 ( .A1(n9138), .A2(n9137), .ZN(n11120) );
  AND2_X1 U8628 ( .A1(n9699), .A2(n15283), .ZN(n10686) );
  AND2_X1 U8629 ( .A1(n9757), .A2(n11063), .ZN(n9762) );
  NAND2_X1 U8630 ( .A1(n7263), .A2(n9427), .ZN(n14083) );
  NAND2_X1 U8631 ( .A1(n7265), .A2(n7264), .ZN(n7263) );
  AND2_X1 U8632 ( .A1(n9317), .A2(n9316), .ZN(n15026) );
  CLKBUF_X1 U8633 ( .A(n10724), .Z(n15335) );
  INV_X1 U8634 ( .A(n15340), .ZN(n15313) );
  INV_X1 U8635 ( .A(n9077), .ZN(n7406) );
  INV_X1 U8636 ( .A(n9521), .ZN(n7332) );
  XNOR2_X1 U8637 ( .A(n9663), .B(n9662), .ZN(n9667) );
  OR2_X1 U8638 ( .A1(n9163), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n9166) );
  INV_X1 U8639 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n9063) );
  INV_X1 U8640 ( .A(n12113), .ZN(n7380) );
  INV_X1 U8641 ( .A(n12078), .ZN(n7381) );
  OR2_X1 U8642 ( .A1(n13023), .A2(n13022), .ZN(n14234) );
  NAND2_X1 U8643 ( .A1(n14311), .A2(n13009), .ZN(n14235) );
  AND2_X1 U8644 ( .A1(n7342), .A2(n14245), .ZN(n7341) );
  NAND2_X1 U8645 ( .A1(n7345), .A2(n7348), .ZN(n7342) );
  OR2_X1 U8646 ( .A1(n12763), .A2(n14250), .ZN(n12784) );
  OR2_X1 U8647 ( .A1(n14257), .A2(n14258), .ZN(n14255) );
  NAND2_X1 U8648 ( .A1(n12075), .A2(n6672), .ZN(n12114) );
  AND2_X1 U8649 ( .A1(n14215), .A2(n13033), .ZN(n14302) );
  OR2_X1 U8650 ( .A1(n12729), .A2(n14305), .ZN(n12751) );
  NAND2_X1 U8651 ( .A1(n11690), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n11982) );
  INV_X1 U8652 ( .A(n7386), .ZN(n7385) );
  AOI21_X1 U8653 ( .B1(n7386), .B2(n7384), .A(n7383), .ZN(n7382) );
  AND2_X1 U8654 ( .A1(n7387), .A2(n14264), .ZN(n7386) );
  AOI21_X1 U8655 ( .B1(n12967), .B2(n7339), .A(n6746), .ZN(n7338) );
  INV_X1 U8656 ( .A(n12967), .ZN(n7340) );
  AND2_X1 U8657 ( .A1(n14878), .A2(n12500), .ZN(n12484) );
  NAND2_X1 U8658 ( .A1(n14382), .A2(n14383), .ZN(n14381) );
  NAND2_X1 U8659 ( .A1(n10178), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10236) );
  NOR2_X1 U8660 ( .A1(n15107), .A2(n6821), .ZN(n11734) );
  NAND2_X1 U8661 ( .A1(n11734), .A2(n11735), .ZN(n12021) );
  XNOR2_X1 U8662 ( .A(n14464), .B(n6818), .ZN(n15117) );
  NAND2_X1 U8663 ( .A1(n15117), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n15116) );
  OR2_X1 U8664 ( .A1(n14509), .A2(n14734), .ZN(n13100) );
  AOI21_X1 U8665 ( .B1(n6969), .B2(n7628), .A(n6732), .ZN(n6967) );
  INV_X1 U8666 ( .A(n12932), .ZN(n14520) );
  NOR2_X1 U8667 ( .A1(n14531), .A2(n7224), .ZN(n7223) );
  INV_X1 U8668 ( .A(n12906), .ZN(n7224) );
  NAND2_X1 U8669 ( .A1(n14589), .A2(n14839), .ZN(n14571) );
  NAND2_X1 U8670 ( .A1(n7616), .A2(n14627), .ZN(n6971) );
  INV_X1 U8671 ( .A(n7616), .ZN(n6975) );
  AND2_X1 U8672 ( .A1(n14628), .A2(n14847), .ZN(n14599) );
  AND2_X1 U8673 ( .A1(n12922), .A2(n7603), .ZN(n7602) );
  OR2_X1 U8674 ( .A1(n14666), .A2(n14650), .ZN(n14651) );
  NAND2_X1 U8675 ( .A1(n12505), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n12666) );
  OR2_X1 U8676 ( .A1(n12666), .A2(n12665), .ZN(n12668) );
  OR2_X1 U8677 ( .A1(n7035), .A2(n14794), .ZN(n14666) );
  OAI21_X1 U8678 ( .B1(n12914), .B2(n6988), .A(n6986), .ZN(n14676) );
  NAND2_X1 U8679 ( .A1(n12462), .A2(n14353), .ZN(n14703) );
  NAND2_X1 U8680 ( .A1(n12462), .A2(n7034), .ZN(n14704) );
  INV_X1 U8681 ( .A(n12309), .ZN(n12307) );
  CLKBUF_X1 U8682 ( .A(n12447), .Z(n12304) );
  AND2_X1 U8683 ( .A1(n12257), .A2(n14300), .ZN(n12318) );
  NAND2_X1 U8684 ( .A1(n11702), .A2(n6673), .ZN(n12105) );
  NAND2_X1 U8685 ( .A1(n11833), .A2(n11832), .ZN(n11838) );
  NAND2_X1 U8686 ( .A1(n11838), .A2(n12847), .ZN(n11972) );
  NOR2_X1 U8687 ( .A1(n11400), .A2(n12577), .ZN(n11702) );
  OR2_X1 U8688 ( .A1(n11506), .A2(n15158), .ZN(n11400) );
  NAND2_X1 U8689 ( .A1(n11331), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n11386) );
  NOR2_X1 U8690 ( .A1(n11496), .A2(n12555), .ZN(n11507) );
  NAND2_X1 U8691 ( .A1(n11578), .A2(n7032), .ZN(n11496) );
  NAND2_X1 U8692 ( .A1(n7613), .A2(n12528), .ZN(n11433) );
  NAND2_X1 U8693 ( .A1(n11632), .A2(n11786), .ZN(n11435) );
  NAND2_X1 U8694 ( .A1(n7622), .A2(n7621), .ZN(n7623) );
  AND2_X1 U8695 ( .A1(n14510), .A2(n14509), .ZN(n14738) );
  AND2_X1 U8696 ( .A1(n12474), .A2(n12486), .ZN(n10888) );
  NAND2_X1 U8697 ( .A1(n10225), .A2(n10224), .ZN(n10512) );
  NAND2_X1 U8698 ( .A1(n9943), .A2(n9935), .ZN(n9920) );
  INV_X1 U8699 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n10479) );
  NAND2_X1 U8700 ( .A1(n6807), .A2(n12215), .ZN(n6806) );
  XNOR2_X1 U8701 ( .A(n9626), .B(n9609), .ZN(n12887) );
  NOR2_X1 U8702 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n7595) );
  NAND2_X1 U8703 ( .A1(n6958), .A2(n6956), .ZN(n12649) );
  AOI22_X1 U8704 ( .A1(n6959), .A2(n9473), .B1(n6776), .B2(n9434), .ZN(n6958)
         );
  NAND2_X1 U8705 ( .A1(n6951), .A2(n9388), .ZN(n9407) );
  NAND2_X1 U8706 ( .A1(n9387), .A2(n9386), .ZN(n6951) );
  AND2_X1 U8707 ( .A1(n10534), .A2(n10285), .ZN(n12240) );
  NAND2_X1 U8708 ( .A1(n9293), .A2(n9292), .ZN(n9312) );
  NOR2_X1 U8709 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .ZN(
        n10132) );
  NAND2_X1 U8710 ( .A1(n7861), .A2(n6995), .ZN(n7905) );
  NAND2_X1 U8711 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n6996), .ZN(n6995) );
  INV_X1 U8712 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6996) );
  NAND2_X1 U8713 ( .A1(n15611), .A2(n7916), .ZN(n7919) );
  NAND2_X1 U8714 ( .A1(n7871), .A2(n7870), .ZN(n7918) );
  AND2_X1 U8715 ( .A1(n7879), .A2(n14415), .ZN(n7929) );
  NOR2_X1 U8716 ( .A1(n7879), .A2(n14415), .ZN(n7930) );
  NOR2_X1 U8717 ( .A1(n7930), .A2(n7880), .ZN(n7897) );
  NOR2_X1 U8718 ( .A1(P3_ADDR_REG_10__SCAN_IN), .A2(n7929), .ZN(n7880) );
  OAI21_X1 U8719 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n7884), .A(n7883), .ZN(
        n7893) );
  OAI21_X1 U8720 ( .B1(n15102), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7299), .ZN(
        n7946) );
  NOR2_X1 U8721 ( .A1(n14914), .A2(P2_ADDR_REG_17__SCAN_IN), .ZN(n7000) );
  OAI21_X1 U8722 ( .B1(n11711), .B2(n7125), .A(n7123), .ZN(n15360) );
  OR2_X1 U8723 ( .A1(n13212), .A2(n13303), .ZN(n6844) );
  NAND2_X1 U8724 ( .A1(n15358), .A2(n11716), .ZN(n11718) );
  NAND2_X1 U8725 ( .A1(n13275), .A2(n13159), .ZN(n13228) );
  NAND2_X1 U8726 ( .A1(n8711), .A2(n8710), .ZN(n13240) );
  AND2_X1 U8727 ( .A1(n15387), .A2(n11093), .ZN(n11094) );
  INV_X1 U8728 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n12012) );
  NAND2_X1 U8729 ( .A1(n12007), .A2(n12006), .ZN(n12010) );
  NAND2_X1 U8730 ( .A1(n13204), .A2(n13156), .ZN(n13277) );
  CLKBUF_X1 U8731 ( .A(n8955), .Z(n11305) );
  NAND2_X1 U8732 ( .A1(n7127), .A2(n7126), .ZN(n15391) );
  NAND2_X1 U8733 ( .A1(n11711), .A2(n11710), .ZN(n7127) );
  INV_X1 U8734 ( .A(n8985), .ZN(n6834) );
  AND2_X1 U8735 ( .A1(n8770), .A2(n8769), .ZN(n13219) );
  INV_X1 U8736 ( .A(n12223), .ZN(n13324) );
  INV_X1 U8737 ( .A(n12013), .ZN(n12004) );
  INV_X1 U8738 ( .A(n11767), .ZN(n11181) );
  INV_X1 U8739 ( .A(n11304), .ZN(n11091) );
  INV_X1 U8740 ( .A(n8952), .ZN(n13327) );
  NAND4_X2 U8741 ( .A1(n8401), .A2(n8403), .A3(n8402), .A4(n8400), .ZN(n13330)
         );
  OR2_X1 U8742 ( .A1(n7745), .A2(n10218), .ZN(n13329) );
  INV_X1 U8743 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n10957) );
  AND2_X1 U8744 ( .A1(n10963), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n10962) );
  INV_X1 U8745 ( .A(n7153), .ZN(n15446) );
  INV_X1 U8746 ( .A(n7151), .ZN(n15444) );
  INV_X1 U8747 ( .A(n6938), .ZN(n15461) );
  INV_X1 U8748 ( .A(n7778), .ZN(n6937) );
  XNOR2_X1 U8749 ( .A(n7780), .B(n10153), .ZN(n11043) );
  NOR2_X1 U8750 ( .A1(n11043), .A2(n15604), .ZN(n11042) );
  OAI21_X1 U8751 ( .B1(n11043), .B2(n7513), .A(n7512), .ZN(n11152) );
  NAND2_X1 U8752 ( .A1(n7514), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7513) );
  NAND2_X1 U8753 ( .A1(n7781), .A2(n7514), .ZN(n7512) );
  INV_X1 U8754 ( .A(n11153), .ZN(n7514) );
  NOR2_X1 U8755 ( .A1(n11895), .A2(n12056), .ZN(n11894) );
  NAND2_X1 U8756 ( .A1(n7156), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7155) );
  INV_X1 U8757 ( .A(n15495), .ZN(n7156) );
  AND2_X1 U8758 ( .A1(n7826), .A2(n11906), .ZN(n6888) );
  INV_X1 U8759 ( .A(n6941), .ZN(n13340) );
  INV_X1 U8760 ( .A(n6858), .ZN(n7734) );
  NOR2_X1 U8761 ( .A1(n13348), .A2(n14937), .ZN(n13347) );
  NOR2_X1 U8762 ( .A1(n13384), .A2(n13617), .ZN(n13383) );
  NAND2_X1 U8763 ( .A1(n10540), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n7508) );
  OR2_X1 U8764 ( .A1(n14921), .A2(n6828), .ZN(n6827) );
  NOR2_X1 U8765 ( .A1(n14917), .A2(n13540), .ZN(n6828) );
  NAND2_X1 U8766 ( .A1(n7464), .A2(n7467), .ZN(n13436) );
  OR2_X1 U8767 ( .A1(n13474), .A2(n7469), .ZN(n7464) );
  AND2_X1 U8768 ( .A1(n7471), .A2(n8798), .ZN(n13448) );
  NAND2_X1 U8769 ( .A1(n7096), .A2(n7097), .ZN(n13457) );
  AND2_X1 U8770 ( .A1(n7100), .A2(n6715), .ZN(n13467) );
  NAND2_X1 U8771 ( .A1(n13481), .A2(n8981), .ZN(n7100) );
  NAND2_X1 U8772 ( .A1(n7064), .A2(n7066), .ZN(n13503) );
  NAND2_X1 U8773 ( .A1(n13529), .A2(n7070), .ZN(n7064) );
  NAND2_X1 U8774 ( .A1(n7072), .A2(n7069), .ZN(n13514) );
  INV_X1 U8775 ( .A(n7071), .ZN(n7069) );
  NAND2_X1 U8776 ( .A1(n13610), .A2(n8885), .ZN(n13522) );
  AND2_X1 U8777 ( .A1(n7088), .A2(n6707), .ZN(n13553) );
  NAND2_X1 U8778 ( .A1(n12369), .A2(n8874), .ZN(n13557) );
  NAND2_X1 U8779 ( .A1(n8977), .A2(n8976), .ZN(n12367) );
  NAND2_X1 U8780 ( .A1(n8585), .A2(n8584), .ZN(n14933) );
  NAND2_X1 U8781 ( .A1(n7498), .A2(n8840), .ZN(n11822) );
  NAND2_X1 U8782 ( .A1(n11939), .A2(n8967), .ZN(n11777) );
  NAND2_X1 U8783 ( .A1(n11540), .A2(n8963), .ZN(n11766) );
  AND3_X1 U8784 ( .A1(n8443), .A2(n8442), .A3(n8441), .ZN(n15545) );
  AND3_X1 U8785 ( .A1(n8432), .A2(n8431), .A3(n8430), .ZN(n11759) );
  INV_X1 U8786 ( .A(n13538), .ZN(n13559) );
  INV_X1 U8787 ( .A(n7222), .ZN(n13626) );
  INV_X1 U8788 ( .A(n8773), .ZN(n13629) );
  INV_X1 U8789 ( .A(n13240), .ZN(n13641) );
  OR2_X1 U8790 ( .A1(n13614), .A2(n13613), .ZN(n13666) );
  NAND2_X1 U8791 ( .A1(n8612), .A2(n8611), .ZN(n13670) );
  AND2_X1 U8792 ( .A1(n8997), .A2(n8996), .ZN(n11006) );
  NAND2_X1 U8793 ( .A1(n13679), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8379) );
  XNOR2_X1 U8794 ( .A(n8759), .B(n8758), .ZN(n13684) );
  NAND2_X1 U8795 ( .A1(n7231), .A2(n8352), .ZN(n8746) );
  OR2_X1 U8796 ( .A1(n8731), .A2(n8351), .ZN(n7231) );
  XNOR2_X1 U8797 ( .A(n7756), .B(P3_IR_REG_22__SCAN_IN), .ZN(n11190) );
  INV_X1 U8798 ( .A(n10704), .ZN(n11313) );
  XNOR2_X1 U8799 ( .A(n8776), .B(n7103), .ZN(n11039) );
  INV_X1 U8800 ( .A(SI_19_), .ZN(n10767) );
  INV_X1 U8801 ( .A(SI_16_), .ZN(n10442) );
  OAI21_X1 U8802 ( .B1(n8581), .B2(n7183), .A(n7181), .ZN(n8596) );
  NAND2_X1 U8803 ( .A1(n8583), .A2(n8330), .ZN(n8594) );
  INV_X1 U8804 ( .A(SI_15_), .ZN(n10316) );
  NAND2_X1 U8805 ( .A1(n8325), .A2(n8326), .ZN(n8554) );
  OAI21_X1 U8806 ( .B1(n8523), .B2(n7190), .A(n7187), .ZN(n8547) );
  INV_X1 U8807 ( .A(SI_11_), .ZN(n10167) );
  NAND2_X1 U8808 ( .A1(n8535), .A2(n8534), .ZN(n8537) );
  NAND2_X1 U8809 ( .A1(n8523), .A2(n8319), .ZN(n8535) );
  XNOR2_X1 U8810 ( .A(n7692), .B(n7691), .ZN(n10163) );
  OR2_X1 U8811 ( .A1(n7695), .A2(n7715), .ZN(n7697) );
  NAND2_X1 U8812 ( .A1(n8479), .A2(n8313), .ZN(n8494) );
  NAND2_X1 U8813 ( .A1(n8311), .A2(n8310), .ZN(n8477) );
  XNOR2_X1 U8814 ( .A(n7702), .B(n7701), .ZN(n15442) );
  NAND2_X1 U8815 ( .A1(n7215), .A2(n8306), .ZN(n8455) );
  NAND2_X1 U8816 ( .A1(n8440), .A2(n8439), .ZN(n7215) );
  XNOR2_X1 U8817 ( .A(n7704), .B(P3_IR_REG_5__SCAN_IN), .ZN(n15434) );
  NAND2_X1 U8818 ( .A1(n7710), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7712) );
  NAND2_X1 U8819 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(P3_IR_REG_0__SCAN_IN), .ZN(
        n7168) );
  INV_X1 U8820 ( .A(P3_IR_REG_1__SCAN_IN), .ZN(n6849) );
  OAI211_X1 U8821 ( .C1(n10923), .C2(n6911), .A(n6909), .B(n11017), .ZN(n11197) );
  INV_X1 U8822 ( .A(n11015), .ZN(n6911) );
  NAND2_X1 U8823 ( .A1(n11016), .A2(n11015), .ZN(n11018) );
  NAND2_X1 U8824 ( .A1(n7551), .A2(n12155), .ZN(n12158) );
  AND2_X1 U8825 ( .A1(n7549), .A2(n6685), .ZN(n11457) );
  NAND2_X1 U8826 ( .A1(n10904), .A2(n10738), .ZN(n13750) );
  NAND2_X1 U8827 ( .A1(n7530), .A2(n7531), .ZN(n13757) );
  INV_X1 U8828 ( .A(n6923), .ZN(n6921) );
  NAND2_X1 U8829 ( .A1(n11923), .A2(n11922), .ZN(n11962) );
  AOI21_X1 U8830 ( .B1(n13814), .B2(n13813), .A(n6677), .ZN(n13787) );
  INV_X1 U8831 ( .A(n15332), .ZN(n11141) );
  NAND2_X1 U8832 ( .A1(n13751), .A2(n10744), .ZN(n10747) );
  NAND2_X1 U8833 ( .A1(n10118), .A2(n7251), .ZN(n9152) );
  INV_X1 U8834 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n11275) );
  AND2_X1 U8835 ( .A1(n6927), .A2(n6925), .ZN(n13820) );
  NAND2_X1 U8836 ( .A1(n6927), .A2(n7524), .ZN(n13822) );
  AOI21_X1 U8837 ( .B1(n6918), .B2(n6920), .A(n6916), .ZN(n6915) );
  INV_X1 U8838 ( .A(n11963), .ZN(n6916) );
  NAND2_X1 U8839 ( .A1(n11673), .A2(n11672), .ZN(n11923) );
  NAND2_X1 U8840 ( .A1(n10913), .A2(n10733), .ZN(n10905) );
  XNOR2_X1 U8841 ( .A(n10737), .B(n10735), .ZN(n10906) );
  INV_X1 U8842 ( .A(n13855), .ZN(n13843) );
  NAND2_X1 U8843 ( .A1(n13802), .A2(n13703), .ZN(n13838) );
  NAND2_X1 U8844 ( .A1(n10923), .A2(n7546), .ZN(n11016) );
  NAND2_X1 U8845 ( .A1(n10923), .A2(n10922), .ZN(n10929) );
  INV_X1 U8846 ( .A(n6817), .ZN(n7538) );
  NAND2_X1 U8847 ( .A1(n7540), .A2(n7541), .ZN(n13850) );
  AND2_X1 U8848 ( .A1(n10752), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13853) );
  INV_X1 U8849 ( .A(n11816), .ZN(n7329) );
  NOR2_X1 U8850 ( .A1(n10011), .A2(n6684), .ZN(n7330) );
  INV_X1 U8851 ( .A(n10010), .ZN(n10014) );
  OAI21_X1 U8852 ( .B1(n10004), .B2(n11063), .A(n10009), .ZN(n10010) );
  INV_X1 U8853 ( .A(n13789), .ZN(n13865) );
  INV_X1 U8854 ( .A(n9794), .ZN(n13887) );
  AND2_X1 U8855 ( .A1(n9257), .A2(n9411), .ZN(n10455) );
  INV_X1 U8856 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n8356) );
  INV_X1 U8857 ( .A(n9952), .ZN(n14101) );
  INV_X1 U8858 ( .A(n13910), .ZN(n14104) );
  AND2_X1 U8859 ( .A1(n13931), .A2(n13930), .ZN(n14113) );
  NAND2_X1 U8860 ( .A1(n7285), .A2(n7289), .ZN(n13945) );
  NAND2_X1 U8861 ( .A1(n7288), .A2(n7293), .ZN(n13960) );
  NAND2_X1 U8862 ( .A1(n7295), .A2(n6695), .ZN(n13966) );
  OR2_X1 U8863 ( .A1(n13982), .A2(n13992), .ZN(n7295) );
  NAND2_X1 U8864 ( .A1(n14055), .A2(n9495), .ZN(n14032) );
  OR2_X1 U8865 ( .A1(n12707), .A2(n9523), .ZN(n9483) );
  NAND2_X1 U8866 ( .A1(n14079), .A2(n9745), .ZN(n14074) );
  NAND2_X1 U8867 ( .A1(n9414), .A2(n9413), .ZN(n13699) );
  NAND2_X1 U8868 ( .A1(n12062), .A2(n9742), .ZN(n14978) );
  NAND2_X1 U8869 ( .A1(n7275), .A2(n7278), .ZN(n12060) );
  NAND2_X1 U8870 ( .A1(n11879), .A2(n7281), .ZN(n7275) );
  NAND2_X1 U8871 ( .A1(n7283), .A2(n9348), .ZN(n14986) );
  INV_X1 U8872 ( .A(n15026), .ZN(n11930) );
  NAND2_X1 U8873 ( .A1(n7396), .A2(n9735), .ZN(n11640) );
  NAND2_X1 U8874 ( .A1(n11558), .A2(n11562), .ZN(n7396) );
  AND2_X1 U8875 ( .A1(n9237), .A2(n9236), .ZN(n11247) );
  NAND2_X1 U8876 ( .A1(n7256), .A2(n9210), .ZN(n11029) );
  OAI21_X1 U8877 ( .B1(n11138), .B2(n9729), .A(n7397), .ZN(n10943) );
  INV_X1 U8878 ( .A(n7398), .ZN(n7397) );
  OAI211_X2 U8879 ( .C1(n9523), .C2(n9106), .A(n9113), .B(n9112), .ZN(n15271)
         );
  OR2_X1 U8880 ( .A1(n14078), .A2(n10684), .ZN(n14094) );
  OR2_X1 U8881 ( .A1(n9150), .A2(n10171), .ZN(n7052) );
  OR3_X1 U8882 ( .A1(n14144), .A2(n14143), .A3(n14142), .ZN(n14180) );
  AND2_X2 U8883 ( .A1(n10968), .A2(n15287), .ZN(n15347) );
  AND2_X1 U8884 ( .A1(n9708), .A2(P2_STATE_REG_SCAN_IN), .ZN(n15289) );
  INV_X1 U8885 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n14187) );
  NAND2_X1 U8886 ( .A1(n9084), .A2(n6804), .ZN(n6857) );
  NOR2_X1 U8887 ( .A1(n7522), .A2(n9658), .ZN(n6804) );
  XNOR2_X1 U8888 ( .A(n9678), .B(P2_IR_REG_24__SCAN_IN), .ZN(n12141) );
  CLKBUF_X1 U8889 ( .A(n9667), .Z(n9664) );
  INV_X1 U8890 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n10871) );
  INV_X1 U8891 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n10766) );
  INV_X1 U8892 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n10192) );
  INV_X1 U8893 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n10195) );
  INV_X1 U8894 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n10198) );
  INV_X1 U8895 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n10189) );
  INV_X1 U8896 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n10188) );
  INV_X1 U8897 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n10182) );
  INV_X1 U8898 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n10186) );
  INV_X1 U8899 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n10183) );
  INV_X1 U8900 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n10171) );
  NAND2_X1 U8901 ( .A1(n15044), .A2(n12967), .ZN(n15046) );
  OAI21_X1 U8902 ( .B1(n10822), .B2(n7359), .A(n7358), .ZN(n10986) );
  NAND2_X1 U8903 ( .A1(n7360), .A2(n10820), .ZN(n7359) );
  NAND2_X1 U8904 ( .A1(n7356), .A2(n10976), .ZN(n7360) );
  NAND2_X1 U8905 ( .A1(n10986), .A2(n10985), .ZN(n11228) );
  NAND2_X1 U8906 ( .A1(n12075), .A2(n12074), .ZN(n12077) );
  NAND2_X1 U8907 ( .A1(n6867), .A2(n6866), .ZN(n6865) );
  NAND2_X1 U8908 ( .A1(n14255), .A2(n12983), .ZN(n14267) );
  NAND2_X1 U8909 ( .A1(n14218), .A2(n14273), .ZN(n7344) );
  NAND2_X1 U8910 ( .A1(n12114), .A2(n12113), .ZN(n12269) );
  NAND2_X1 U8911 ( .A1(n14292), .A2(n14291), .ZN(n15044) );
  AND2_X1 U8912 ( .A1(n15058), .A2(n15059), .ZN(n12412) );
  INV_X1 U8913 ( .A(n14369), .ZN(n15057) );
  INV_X1 U8914 ( .A(n14367), .ZN(n15054) );
  INV_X1 U8915 ( .A(n10829), .ZN(n7357) );
  NAND2_X1 U8916 ( .A1(n14344), .A2(n14343), .ZN(n14342) );
  XNOR2_X1 U8917 ( .A(n12978), .B(n12976), .ZN(n14344) );
  AND2_X1 U8918 ( .A1(n10527), .A2(n12879), .ZN(n14349) );
  NAND2_X1 U8919 ( .A1(n6963), .A2(n7598), .ZN(n6962) );
  NAND2_X1 U8920 ( .A1(n12804), .A2(n12803), .ZN(n14357) );
  NAND2_X1 U8921 ( .A1(n12791), .A2(n12790), .ZN(n14358) );
  OAI21_X1 U8922 ( .B1(n10322), .B2(n14396), .A(n10321), .ZN(n14401) );
  AOI21_X1 U8923 ( .B1(n10672), .B2(P1_REG1_REG_4__SCAN_IN), .A(n10661), .ZN(
        n10323) );
  OAI21_X1 U8924 ( .B1(n10472), .B2(n10467), .A(n10401), .ZN(n10470) );
  NOR2_X1 U8925 ( .A1(n10413), .A2(n10414), .ZN(n10412) );
  NOR2_X1 U8926 ( .A1(n10429), .A2(n10430), .ZN(n14430) );
  NOR2_X1 U8927 ( .A1(n14489), .A2(n14781), .ZN(n14717) );
  NAND2_X1 U8928 ( .A1(n6713), .A2(n7036), .ZN(n14489) );
  OAI21_X1 U8929 ( .B1(n14509), .B2(n7037), .A(n14488), .ZN(n7036) );
  AND2_X1 U8930 ( .A1(n6851), .A2(n6850), .ZN(n14721) );
  OR2_X1 U8931 ( .A1(n7037), .A2(n14509), .ZN(n6851) );
  XNOR2_X1 U8932 ( .A(n13099), .B(n13114), .ZN(n14731) );
  NAND2_X1 U8933 ( .A1(n13098), .A2(n6734), .ZN(n13099) );
  NAND2_X1 U8934 ( .A1(n6966), .A2(n6969), .ZN(n14530) );
  NAND2_X1 U8935 ( .A1(n14566), .A2(n7627), .ZN(n6966) );
  NAND2_X1 U8936 ( .A1(n12905), .A2(n12904), .ZN(n14549) );
  NAND2_X1 U8937 ( .A1(n14639), .A2(n6675), .ZN(n14617) );
  NAND2_X1 U8938 ( .A1(n7204), .A2(n12897), .ZN(n14661) );
  NAND2_X1 U8939 ( .A1(n12894), .A2(n12893), .ZN(n14696) );
  OAI21_X1 U8940 ( .B1(n12914), .B2(n12915), .A(n12917), .ZN(n14692) );
  INV_X1 U8941 ( .A(n6985), .ZN(n14691) );
  NAND2_X1 U8942 ( .A1(n12294), .A2(n12293), .ZN(n15050) );
  NAND2_X1 U8943 ( .A1(n12296), .A2(n12295), .ZN(n12298) );
  NAND2_X1 U8944 ( .A1(n12169), .A2(n12168), .ZN(n12608) );
  CLKBUF_X1 U8945 ( .A(n12253), .Z(n12174) );
  OAI21_X1 U8946 ( .B1(n11833), .B2(n6671), .A(n6980), .ZN(n12093) );
  NAND2_X1 U8947 ( .A1(n11397), .A2(n11681), .ZN(n11687) );
  INV_X1 U8948 ( .A(n14709), .ZN(n15140) );
  CLKBUF_X1 U8949 ( .A(n11481), .Z(n11482) );
  NAND2_X1 U8950 ( .A1(n7612), .A2(n12528), .ZN(n11420) );
  INV_X1 U8951 ( .A(n7613), .ZN(n7612) );
  CLKBUF_X1 U8952 ( .A(n11355), .Z(n14378) );
  NOR2_X1 U8953 ( .A1(n11516), .A2(n10893), .ZN(n14801) );
  INV_X1 U8954 ( .A(n14801), .ZN(n15181) );
  INV_X1 U8955 ( .A(n12957), .ZN(n14300) );
  CLKBUF_X1 U8956 ( .A(n10247), .Z(n10248) );
  NOR2_X1 U8957 ( .A1(n6863), .A2(n6862), .ZN(n6861) );
  OR2_X1 U8958 ( .A1(n10210), .A2(n7242), .ZN(n6864) );
  NOR2_X1 U8959 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_31__SCAN_IN), .ZN(
        n6862) );
  NAND2_X1 U8960 ( .A1(n9454), .A2(n9436), .ZN(n12659) );
  INV_X1 U8961 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10879) );
  INV_X1 U8962 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n10763) );
  INV_X1 U8963 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n10259) );
  INV_X1 U8964 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n10240) );
  INV_X1 U8965 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n10205) );
  INV_X1 U8966 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n10175) );
  INV_X1 U8967 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n10166) );
  INV_X1 U8968 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n10144) );
  NAND2_X1 U8969 ( .A1(n9212), .A2(n7026), .ZN(n11338) );
  NAND2_X1 U8970 ( .A1(n9198), .A2(n7027), .ZN(n7026) );
  NOR2_X1 U8971 ( .A1(n9199), .A2(n7028), .ZN(n7027) );
  OR2_X1 U8972 ( .A1(n10143), .A2(n10142), .ZN(n10400) );
  INV_X1 U8973 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n11326) );
  NOR2_X1 U8974 ( .A1(n10135), .A2(n14864), .ZN(n10136) );
  INV_X1 U8975 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n11220) );
  CLKBUF_X1 U8976 ( .A(n10119), .Z(n10120) );
  NOR2_X1 U8977 ( .A1(n15622), .A2(n7910), .ZN(n14889) );
  NOR2_X1 U8978 ( .A1(n15620), .A2(n15619), .ZN(n7911) );
  XNOR2_X1 U8979 ( .A(n7914), .B(n7302), .ZN(n15613) );
  INV_X1 U8980 ( .A(n7915), .ZN(n7302) );
  NAND2_X1 U8981 ( .A1(n15613), .A2(n15612), .ZN(n15611) );
  XNOR2_X1 U8982 ( .A(n7919), .B(n7005), .ZN(n14893) );
  NAND2_X1 U8983 ( .A1(n14903), .A2(n7305), .ZN(n7010) );
  NAND2_X1 U8984 ( .A1(n6681), .A2(n7008), .ZN(n7007) );
  NOR2_X1 U8985 ( .A1(n7934), .A2(n7935), .ZN(n15085) );
  NAND2_X1 U8986 ( .A1(n15087), .A2(n15088), .ZN(n15084) );
  NAND2_X1 U8987 ( .A1(n15086), .A2(n15084), .ZN(n15090) );
  NAND2_X1 U8988 ( .A1(n15089), .A2(n7300), .ZN(n15094) );
  OAI21_X1 U8989 ( .B1(n15090), .B2(n15091), .A(n7301), .ZN(n7300) );
  INV_X1 U8990 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n7301) );
  NAND2_X1 U8991 ( .A1(n15094), .A2(n15095), .ZN(n15093) );
  NAND2_X1 U8992 ( .A1(n6997), .A2(n15093), .ZN(n15098) );
  OAI21_X1 U8993 ( .B1(n15094), .B2(n15095), .A(n6998), .ZN(n6997) );
  INV_X1 U8994 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n6998) );
  NOR2_X1 U8995 ( .A1(n7940), .A2(n7941), .ZN(n15101) );
  AND2_X1 U8996 ( .A1(n7940), .A2(n7941), .ZN(n15102) );
  NOR2_X1 U8997 ( .A1(n7946), .A2(n7947), .ZN(n14914) );
  AND2_X1 U8998 ( .A1(n7946), .A2(n7947), .ZN(n14915) );
  NAND2_X1 U8999 ( .A1(n6683), .A2(n7135), .ZN(n7129) );
  NOR2_X1 U9000 ( .A1(n13388), .A2(n7743), .ZN(n14923) );
  OAI21_X1 U9001 ( .B1(n7860), .B2(n15530), .A(n6845), .ZN(P3_U3201) );
  AOI21_X1 U9002 ( .B1(n7506), .B2(n10603), .A(n7859), .ZN(n6845) );
  XNOR2_X1 U9003 ( .A(n6827), .B(n7845), .ZN(n7860) );
  XNOR2_X1 U9004 ( .A(n7507), .B(n7843), .ZN(n7506) );
  AOI21_X1 U9005 ( .B1(n13128), .B2(n13543), .A(n13127), .ZN(n6838) );
  OAI21_X1 U9006 ( .B1(n7115), .B2(n9022), .A(n6880), .ZN(P3_U3488) );
  INV_X1 U9007 ( .A(n6881), .ZN(n6880) );
  OAI21_X1 U9008 ( .B1(n7116), .B2(n9022), .A(n9025), .ZN(n6881) );
  AND2_X1 U9009 ( .A1(n9024), .A2(n9023), .ZN(n9025) );
  MUX2_X1 U9010 ( .A(n13573), .B(n13630), .S(n15607), .Z(n13574) );
  OAI21_X1 U9011 ( .B1(n9035), .B2(n13674), .A(n9034), .ZN(n9036) );
  OAI22_X1 U9012 ( .A1(n13410), .A2(n13674), .B1(n15591), .B2(n9048), .ZN(
        n9049) );
  MUX2_X1 U9013 ( .A(n13631), .B(n13630), .S(n15591), .Z(n13632) );
  NAND2_X1 U9014 ( .A1(n6899), .A2(n6908), .ZN(n6897) );
  INV_X1 U9015 ( .A(n9718), .ZN(n9761) );
  OAI21_X1 U9016 ( .B1(n14108), .B2(n15269), .A(n9717), .ZN(n9718) );
  NAND2_X1 U9017 ( .A1(n15355), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6802) );
  INV_X1 U9018 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n7023) );
  CLKBUF_X1 U9019 ( .A(n14379), .Z(P1_U4016) );
  INV_X1 U9020 ( .A(n6841), .ZN(n6840) );
  OAI21_X1 U9021 ( .B1(n14830), .B2(n14352), .A(n14213), .ZN(n6841) );
  NAND2_X1 U9022 ( .A1(n7371), .A2(n14341), .ZN(n7368) );
  AND2_X1 U9023 ( .A1(n6820), .A2(n6819), .ZN(n14484) );
  INV_X1 U9024 ( .A(n14737), .ZN(n14732) );
  INV_X1 U9025 ( .A(n7006), .ZN(n14899) );
  NAND2_X1 U9026 ( .A1(n6796), .A2(n14903), .ZN(n14902) );
  XNOR2_X1 U9027 ( .A(n8295), .B(n8288), .ZN(n7306) );
  NOR2_X1 U9028 ( .A1(n14882), .A2(n7308), .ZN(n7307) );
  AND2_X1 U9029 ( .A1(n7381), .A2(n12074), .ZN(n6672) );
  AND2_X1 U9030 ( .A1(n7043), .A2(n7042), .ZN(n6673) );
  AND2_X1 U9031 ( .A1(n7600), .A2(n6984), .ZN(n6674) );
  NOR2_X1 U9032 ( .A1(n13262), .A2(n13483), .ZN(n7136) );
  MUX2_X2 U9033 ( .A(n12500), .B(n12478), .S(n12499), .Z(n12496) );
  XNOR2_X1 U9034 ( .A(n9455), .B(P2_IR_REG_19__SCAN_IN), .ZN(n9709) );
  INV_X2 U9035 ( .A(n13026), .ZN(n13085) );
  INV_X2 U9036 ( .A(n13026), .ZN(n13070) );
  AND2_X1 U9037 ( .A1(n12901), .A2(n14627), .ZN(n6675) );
  INV_X1 U9038 ( .A(n11116), .ZN(n7049) );
  INV_X2 U9039 ( .A(n9764), .ZN(n9870) );
  CLKBUF_X3 U9040 ( .A(n9764), .Z(n10005) );
  AND2_X1 U9041 ( .A1(n10029), .A2(n10135), .ZN(n10487) );
  OR2_X1 U9042 ( .A1(n9473), .A2(n9472), .ZN(n6676) );
  INV_X1 U9043 ( .A(n12847), .ZN(n7607) );
  AND2_X1 U9044 ( .A1(n13725), .A2(n13726), .ZN(n6677) );
  AND2_X1 U9045 ( .A1(n12762), .A2(n7557), .ZN(n6678) );
  XNOR2_X1 U9046 ( .A(n14650), .B(n14619), .ZN(n12697) );
  INV_X1 U9047 ( .A(n12697), .ZN(n14642) );
  AND2_X1 U9048 ( .A1(n14589), .A2(n7045), .ZN(n6679) );
  INV_X1 U9049 ( .A(n13447), .ZN(n7091) );
  INV_X1 U9050 ( .A(n7175), .ZN(n11490) );
  OR2_X1 U9051 ( .A1(n12268), .A2(n7380), .ZN(n6680) );
  INV_X1 U9052 ( .A(n11355), .ZN(n6868) );
  INV_X1 U9053 ( .A(n14903), .ZN(n7013) );
  OR2_X1 U9054 ( .A1(n7928), .A2(n7927), .ZN(n6681) );
  INV_X1 U9055 ( .A(n8874), .ZN(n7431) );
  AND2_X1 U9056 ( .A1(n9905), .A2(n7439), .ZN(n6682) );
  NAND2_X1 U9057 ( .A1(n9874), .A2(n9873), .ZN(n7493) );
  INV_X1 U9058 ( .A(n7493), .ZN(n7492) );
  AND2_X1 U9059 ( .A1(n7131), .A2(n15390), .ZN(n6683) );
  NAND2_X1 U9060 ( .A1(n9525), .A2(n9524), .ZN(n14029) );
  INV_X1 U9061 ( .A(n14029), .ZN(n7056) );
  AND3_X1 U9062 ( .A1(n14101), .A2(n10005), .A3(n13912), .ZN(n6684) );
  NAND2_X1 U9063 ( .A1(n11449), .A2(n11448), .ZN(n6685) );
  NAND2_X1 U9064 ( .A1(n11837), .A2(n11836), .ZN(n12589) );
  INV_X1 U9065 ( .A(n13238), .ZN(n13419) );
  NAND2_X1 U9066 ( .A1(n8729), .A2(n8728), .ZN(n13238) );
  INV_X1 U9067 ( .A(n7628), .ZN(n7627) );
  NAND2_X1 U9068 ( .A1(n14550), .A2(n12930), .ZN(n7628) );
  AND2_X1 U9069 ( .A1(n12728), .A2(n6961), .ZN(n6686) );
  AND2_X1 U9070 ( .A1(n15008), .A2(n13876), .ZN(n6687) );
  INV_X1 U9071 ( .A(n12609), .ZN(n7571) );
  NOR2_X1 U9072 ( .A1(n11274), .A2(n7548), .ZN(n6688) );
  INV_X1 U9073 ( .A(n6987), .ZN(n6986) );
  OAI21_X1 U9074 ( .B1(n6988), .B2(n12917), .A(n12918), .ZN(n6987) );
  NAND2_X1 U9075 ( .A1(n12227), .A2(n12398), .ZN(n6689) );
  AND2_X1 U9076 ( .A1(n7592), .A2(n12796), .ZN(n6690) );
  INV_X1 U9077 ( .A(n14273), .ZN(n7347) );
  AND2_X1 U9078 ( .A1(n6786), .A2(n8976), .ZN(n6691) );
  INV_X1 U9079 ( .A(n11525), .ZN(n7108) );
  NAND2_X1 U9080 ( .A1(n11975), .A2(n11974), .ZN(n12592) );
  INV_X1 U9081 ( .A(n12592), .ZN(n7042) );
  NAND2_X1 U9082 ( .A1(n11702), .A2(n15166), .ZN(n6692) );
  INV_X1 U9083 ( .A(n8600), .ZN(n8646) );
  AND3_X1 U9084 ( .A1(n10992), .A2(n10993), .A3(n10994), .ZN(n6693) );
  INV_X1 U9085 ( .A(n12087), .ZN(n7610) );
  OR2_X1 U9086 ( .A1(n13990), .A2(n13867), .ZN(n6695) );
  INV_X1 U9087 ( .A(n9838), .ZN(n7480) );
  AND2_X1 U9088 ( .A1(n14235), .A2(n13025), .ZN(n6697) );
  AND2_X1 U9089 ( .A1(n7344), .A2(n14274), .ZN(n6698) );
  INV_X1 U9090 ( .A(n10617), .ZN(n11858) );
  OR2_X1 U9091 ( .A1(n15008), .A2(n13876), .ZN(n6699) );
  AND4_X1 U9092 ( .A1(n9062), .A2(n9061), .A3(n9127), .A4(n9164), .ZN(n6700)
         );
  AND2_X1 U9093 ( .A1(n9360), .A2(n9359), .ZN(n15014) );
  OR2_X1 U9094 ( .A1(n15021), .A2(n13878), .ZN(n6701) );
  AND2_X1 U9095 ( .A1(n7101), .A2(n8981), .ZN(n6702) );
  AND2_X1 U9096 ( .A1(n7208), .A2(n8310), .ZN(n6703) );
  INV_X1 U9097 ( .A(n14131), .ZN(n13990) );
  NAND2_X1 U9098 ( .A1(n9564), .A2(n9563), .ZN(n14131) );
  AND2_X1 U9099 ( .A1(n12893), .A2(n12624), .ZN(n12915) );
  NAND2_X1 U9100 ( .A1(n14507), .A2(n12937), .ZN(n12938) );
  AND2_X1 U9101 ( .A1(n9881), .A2(n9880), .ZN(n6704) );
  AND2_X1 U9102 ( .A1(n7096), .A2(n7094), .ZN(n6705) );
  AND2_X1 U9103 ( .A1(n9574), .A2(n9573), .ZN(n13975) );
  AND2_X1 U9104 ( .A1(n9075), .A2(n9076), .ZN(n6706) );
  NAND2_X1 U9105 ( .A1(n12527), .A2(n12526), .ZN(n13039) );
  OR2_X1 U9106 ( .A1(n13143), .A2(n13256), .ZN(n6707) );
  NAND2_X1 U9107 ( .A1(n11709), .A2(n11767), .ZN(n6708) );
  XNOR2_X1 U9108 ( .A(n13722), .B(n13721), .ZN(n13742) );
  NAND2_X1 U9109 ( .A1(n14624), .A2(n12926), .ZN(n14598) );
  NAND2_X1 U9110 ( .A1(n7606), .A2(n12920), .ZN(n14657) );
  NAND2_X1 U9111 ( .A1(n12640), .A2(n12639), .ZN(n14683) );
  INV_X1 U9112 ( .A(n14619), .ZN(n14658) );
  INV_X1 U9113 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n7862) );
  AND2_X1 U9114 ( .A1(n10945), .A2(n13886), .ZN(n6709) );
  NAND2_X1 U9115 ( .A1(n12795), .A2(n12794), .ZN(n14329) );
  INV_X1 U9116 ( .A(n14329), .ZN(n7044) );
  OR2_X1 U9117 ( .A1(n9956), .A2(n6682), .ZN(n6710) );
  OR2_X1 U9118 ( .A1(n13990), .A2(n13788), .ZN(n6711) );
  AND2_X1 U9119 ( .A1(n8930), .A2(n7222), .ZN(n6712) );
  INV_X1 U9120 ( .A(n13767), .ZN(n6907) );
  INV_X1 U9121 ( .A(n10942), .ZN(n10946) );
  OR3_X1 U9122 ( .A1(n14509), .A2(n14488), .A3(n7037), .ZN(n6713) );
  AND2_X1 U9123 ( .A1(n14108), .A2(n14107), .ZN(n6714) );
  NAND2_X1 U9124 ( .A1(n13653), .A2(n13197), .ZN(n6715) );
  INV_X1 U9125 ( .A(n15021), .ZN(n11888) );
  AND2_X1 U9126 ( .A1(n9338), .A2(n9337), .ZN(n15021) );
  AND2_X1 U9127 ( .A1(n7110), .A2(n7108), .ZN(n6716) );
  NAND2_X1 U9128 ( .A1(n10132), .A2(n10133), .ZN(n10145) );
  AND2_X1 U9129 ( .A1(n11712), .A2(n13326), .ZN(n6717) );
  OR2_X1 U9130 ( .A1(n9835), .A2(n9834), .ZN(n6718) );
  NOR2_X1 U9131 ( .A1(n13347), .A2(n7787), .ZN(n6719) );
  NAND2_X1 U9132 ( .A1(n11686), .A2(n11685), .ZN(n12580) );
  NAND2_X1 U9133 ( .A1(n8639), .A2(n8638), .ZN(n13153) );
  INV_X1 U9134 ( .A(n7058), .ZN(n13940) );
  INV_X1 U9135 ( .A(n9426), .ZN(n7264) );
  NOR2_X1 U9136 ( .A1(n9956), .A2(n9909), .ZN(n6720) );
  NOR2_X1 U9137 ( .A1(n15014), .A2(n12144), .ZN(n6721) );
  AND2_X1 U9138 ( .A1(n14547), .A2(n12906), .ZN(n6722) );
  INV_X1 U9139 ( .A(n13528), .ZN(n13546) );
  AND2_X1 U9140 ( .A1(n8885), .A2(n8884), .ZN(n13528) );
  AND2_X1 U9141 ( .A1(n13975), .A2(n9895), .ZN(n6723) );
  NAND2_X1 U9142 ( .A1(n14589), .A2(n7047), .ZN(n7048) );
  AND2_X1 U9143 ( .A1(n14543), .A2(n12931), .ZN(n6724) );
  INV_X1 U9144 ( .A(n7095), .ZN(n7094) );
  NAND2_X1 U9145 ( .A1(n13454), .A2(n7097), .ZN(n7095) );
  OR2_X1 U9146 ( .A1(n9096), .A2(n15185), .ZN(n6725) );
  AND2_X1 U9147 ( .A1(n7524), .A2(n6926), .ZN(n6925) );
  AND2_X1 U9148 ( .A1(n12613), .A2(n12615), .ZN(n12854) );
  AND2_X1 U9149 ( .A1(n13160), .A2(n13159), .ZN(n6726) );
  INV_X1 U9150 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n7309) );
  AND2_X1 U9151 ( .A1(n8978), .A2(n6707), .ZN(n6727) );
  AND2_X1 U9152 ( .A1(n7540), .A2(n7538), .ZN(n6728) );
  AND2_X1 U9153 ( .A1(n7191), .A2(n7194), .ZN(n6729) );
  NAND2_X1 U9154 ( .A1(n12854), .A2(n12611), .ZN(n6730) );
  AND2_X1 U9155 ( .A1(n8647), .A2(n8885), .ZN(n6731) );
  AND2_X1 U9156 ( .A1(n14751), .A2(n14524), .ZN(n6732) );
  AND2_X1 U9157 ( .A1(n11680), .A2(n11587), .ZN(n6733) );
  NAND2_X1 U9158 ( .A1(n14734), .A2(n14356), .ZN(n6734) );
  AND2_X1 U9159 ( .A1(n7422), .A2(n7421), .ZN(n6735) );
  AND2_X1 U9160 ( .A1(n7260), .A2(n9452), .ZN(n6736) );
  AND2_X1 U9161 ( .A1(n9069), .A2(n7522), .ZN(n6737) );
  AND2_X1 U9162 ( .A1(n7065), .A2(n13508), .ZN(n6738) );
  INV_X1 U9163 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n7522) );
  NOR2_X1 U9164 ( .A1(n12592), .A2(n14369), .ZN(n6739) );
  AND2_X1 U9165 ( .A1(n8856), .A2(n8855), .ZN(n6740) );
  NOR2_X1 U9166 ( .A1(n14633), .A2(n14239), .ZN(n6741) );
  NOR2_X1 U9167 ( .A1(n14146), .A2(n13831), .ZN(n6742) );
  NOR2_X1 U9168 ( .A1(n11265), .A2(n13885), .ZN(n6743) );
  OR2_X1 U9169 ( .A1(n13670), .A2(n13532), .ZN(n8879) );
  INV_X1 U9170 ( .A(n9516), .ZN(n7274) );
  INV_X1 U9171 ( .A(n9972), .ZN(n9606) );
  OR2_X1 U9172 ( .A1(n14122), .A2(n13789), .ZN(n9972) );
  NAND2_X1 U9173 ( .A1(n12925), .A2(n12856), .ZN(n14624) );
  AND2_X1 U9174 ( .A1(n9332), .A2(n10180), .ZN(n6744) );
  NAND2_X1 U9175 ( .A1(n7130), .A2(n7137), .ZN(n6745) );
  INV_X1 U9176 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9658) );
  INV_X1 U9177 ( .A(n12591), .ZN(n7562) );
  NOR2_X1 U9178 ( .A1(n12970), .A2(n12969), .ZN(n6746) );
  NAND2_X1 U9179 ( .A1(n12504), .A2(n12503), .ZN(n6747) );
  NAND2_X1 U9180 ( .A1(n13766), .A2(n13765), .ZN(n6748) );
  INV_X1 U9181 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7140) );
  AND2_X1 U9182 ( .A1(n15008), .A2(n15021), .ZN(n6749) );
  AND2_X1 U9183 ( .A1(n8915), .A2(n13435), .ZN(n6750) );
  INV_X1 U9184 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n10030) );
  AND2_X1 U9185 ( .A1(n12602), .A2(n12601), .ZN(n6751) );
  OR2_X1 U9186 ( .A1(n13474), .A2(n8800), .ZN(n7471) );
  AND2_X1 U9187 ( .A1(n7280), .A2(n6699), .ZN(n6752) );
  INV_X1 U9188 ( .A(n13306), .ZN(n13637) );
  NAND2_X1 U9189 ( .A1(n8721), .A2(n8720), .ZN(n13306) );
  AND2_X1 U9190 ( .A1(n9540), .A2(n9539), .ZN(n14008) );
  INV_X1 U9191 ( .A(n14008), .ZN(n14136) );
  AND2_X1 U9192 ( .A1(n7545), .A2(n7544), .ZN(n6753) );
  NAND2_X1 U9193 ( .A1(n13458), .A2(n8913), .ZN(n6754) );
  NOR2_X1 U9194 ( .A1(n15014), .A2(n13877), .ZN(n6755) );
  INV_X1 U9195 ( .A(n13454), .ZN(n13458) );
  NAND2_X1 U9196 ( .A1(n8707), .A2(n8798), .ZN(n13454) );
  AND2_X1 U9197 ( .A1(n8931), .A2(n8928), .ZN(n6756) );
  INV_X1 U9198 ( .A(n7067), .ZN(n7066) );
  OAI21_X1 U9199 ( .B1(n7068), .B2(n13546), .A(n7075), .ZN(n7067) );
  INV_X1 U9200 ( .A(P3_ADDR_REG_1__SCAN_IN), .ZN(n8245) );
  INV_X1 U9201 ( .A(n7580), .ZN(n7579) );
  NAND2_X1 U9202 ( .A1(n12740), .A2(n12739), .ZN(n7580) );
  INV_X1 U9203 ( .A(n12797), .ZN(n7592) );
  OR2_X1 U9204 ( .A1(n12808), .A2(n6690), .ZN(n6757) );
  OR2_X1 U9205 ( .A1(n6870), .A2(n7786), .ZN(n6758) );
  INV_X1 U9206 ( .A(n9991), .ZN(n13944) );
  OR2_X1 U9207 ( .A1(n13720), .A2(n13719), .ZN(n6759) );
  AND2_X1 U9208 ( .A1(n8840), .A2(n8842), .ZN(n6760) );
  XNOR2_X1 U9209 ( .A(n9331), .B(n10180), .ZN(n9329) );
  MUX2_X1 U9210 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n9181), .Z(n9143) );
  INV_X1 U9211 ( .A(n9143), .ZN(n9142) );
  AND2_X1 U9212 ( .A1(n7034), .A2(n14859), .ZN(n6761) );
  AND2_X1 U9213 ( .A1(n7045), .A2(n7044), .ZN(n6762) );
  INV_X1 U9214 ( .A(n13402), .ZN(n7221) );
  NOR2_X1 U9215 ( .A1(n9451), .A2(n7262), .ZN(n7261) );
  NAND2_X1 U9216 ( .A1(n14072), .A2(n13842), .ZN(n6763) );
  AND2_X1 U9217 ( .A1(n7411), .A2(n7410), .ZN(n6764) );
  AND2_X1 U9218 ( .A1(n6839), .A2(n6838), .ZN(n6765) );
  AND2_X1 U9219 ( .A1(n12898), .A2(n12897), .ZN(n6766) );
  AND2_X1 U9220 ( .A1(n11688), .A2(n11681), .ZN(n6767) );
  AND2_X1 U9221 ( .A1(n12008), .A2(n12006), .ZN(n6768) );
  AND2_X1 U9222 ( .A1(n14639), .A2(n12901), .ZN(n6769) );
  AND2_X1 U9223 ( .A1(n7141), .A2(n7140), .ZN(n6770) );
  AND2_X1 U9224 ( .A1(n7566), .A2(n7565), .ZN(n6771) );
  INV_X1 U9225 ( .A(n9802), .ZN(n7445) );
  AND2_X1 U9226 ( .A1(n6683), .A2(n6745), .ZN(n6772) );
  NAND3_X1 U9227 ( .A1(n10029), .A2(n10135), .A3(n7624), .ZN(n6773) );
  INV_X1 U9228 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n6890) );
  INV_X1 U9229 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n7242) );
  INV_X1 U9230 ( .A(n12579), .ZN(n7588) );
  INV_X1 U9231 ( .A(n7012), .ZN(n7011) );
  NAND2_X1 U9232 ( .A1(n7013), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n7012) );
  INV_X1 U9233 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n9078) );
  NAND2_X1 U9234 ( .A1(n6905), .A2(n6903), .ZN(n6775) );
  INV_X1 U9235 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n7375) );
  INV_X1 U9236 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n10979) );
  AND2_X1 U9237 ( .A1(n12528), .A2(n11319), .ZN(n11419) );
  INV_X1 U9238 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7103) );
  OR2_X1 U9239 ( .A1(n11561), .A2(n11562), .ZN(n11559) );
  INV_X1 U9240 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6853) );
  AND4_X1 U9241 ( .A1(n8533), .A2(n8532), .A3(n8531), .A4(n8530), .ZN(n12390)
         );
  INV_X1 U9242 ( .A(n14359), .ZN(n6822) );
  NAND2_X1 U9243 ( .A1(n11972), .A2(n11971), .ZN(n12088) );
  INV_X1 U9244 ( .A(n14244), .ZN(n7346) );
  INV_X1 U9245 ( .A(n14301), .ZN(n7353) );
  NAND2_X1 U9246 ( .A1(n12243), .A2(n12852), .ZN(n12296) );
  AND2_X1 U9247 ( .A1(n9470), .A2(n9473), .ZN(n6776) );
  NOR2_X2 U9248 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_12__SCAN_IN), .ZN(
        n10757) );
  AND2_X1 U9249 ( .A1(n14948), .A2(n13323), .ZN(n6777) );
  OR2_X1 U9250 ( .A1(n12954), .A2(n12953), .ZN(n6778) );
  NOR2_X1 U9251 ( .A1(n11901), .A2(n7784), .ZN(n6779) );
  NOR2_X1 U9252 ( .A1(n11894), .A2(n7732), .ZN(n6780) );
  INV_X1 U9253 ( .A(n7281), .ZN(n7280) );
  NOR2_X1 U9254 ( .A1(n9368), .A2(n7282), .ZN(n7281) );
  INV_X1 U9255 ( .A(n7070), .ZN(n7068) );
  NOR2_X1 U9256 ( .A1(n8980), .A2(n7071), .ZN(n7070) );
  INV_X1 U9257 ( .A(n7138), .ZN(n7137) );
  NOR2_X1 U9258 ( .A1(n13198), .A2(n13322), .ZN(n7138) );
  AND2_X1 U9259 ( .A1(n7530), .A2(n7528), .ZN(n6781) );
  NAND3_X1 U9260 ( .A1(n6928), .A2(n9234), .A3(n7406), .ZN(n6782) );
  INV_X1 U9261 ( .A(n7145), .ZN(n12394) );
  NAND2_X1 U9262 ( .A1(n7146), .A2(n12392), .ZN(n7145) );
  NAND2_X1 U9263 ( .A1(n7754), .A2(n7653), .ZN(n6783) );
  AND2_X1 U9264 ( .A1(n9502), .A2(SI_20_), .ZN(n6784) );
  OR2_X1 U9265 ( .A1(n12266), .A2(n12267), .ZN(n6785) );
  NAND2_X1 U9266 ( .A1(n13143), .A2(n13256), .ZN(n6786) );
  INV_X1 U9267 ( .A(n7059), .ZN(n14980) );
  NOR2_X1 U9268 ( .A1(n11885), .A2(n7060), .ZN(n7059) );
  NAND2_X1 U9269 ( .A1(n9824), .A2(n9825), .ZN(n6787) );
  INV_X1 U9270 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n10278) );
  INV_X1 U9271 ( .A(n13566), .ZN(n13541) );
  INV_X2 U9272 ( .A(n15355), .ZN(n15357) );
  NAND2_X1 U9273 ( .A1(n11203), .A2(n11204), .ZN(n11273) );
  AND2_X1 U9274 ( .A1(n11702), .A2(n7043), .ZN(n6788) );
  AND2_X2 U9275 ( .A1(n9031), .A2(n10562), .ZN(n15591) );
  INV_X1 U9276 ( .A(n13869), .ZN(n7273) );
  AND2_X1 U9277 ( .A1(n15500), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n6789) );
  INV_X1 U9278 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n12708) );
  AND2_X1 U9279 ( .A1(n8338), .A2(n7203), .ZN(n6790) );
  NOR2_X1 U9280 ( .A1(n11042), .A2(n7781), .ZN(n6791) );
  NOR2_X1 U9281 ( .A1(n11044), .A2(n7729), .ZN(n6792) );
  INV_X1 U9282 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n7005) );
  AND2_X1 U9283 ( .A1(n6938), .A2(n6937), .ZN(n6793) );
  AND2_X1 U9284 ( .A1(n7109), .A2(n7110), .ZN(n6794) );
  AND2_X1 U9285 ( .A1(n11818), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n6795) );
  AND2_X1 U9286 ( .A1(n7006), .A2(n6681), .ZN(n6796) );
  AND2_X1 U9287 ( .A1(n7127), .A2(n6708), .ZN(n6797) );
  INV_X1 U9288 ( .A(n13859), .ZN(n6908) );
  OR2_X1 U9289 ( .A1(n10696), .A2(n10695), .ZN(n13859) );
  INV_X1 U9290 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7203) );
  INV_X1 U9291 ( .A(n14474), .ZN(n6818) );
  INV_X1 U9292 ( .A(n10253), .ZN(n6870) );
  INV_X1 U9293 ( .A(SI_22_), .ZN(n6885) );
  AND2_X1 U9294 ( .A1(n10527), .A2(n10516), .ZN(n14341) );
  INV_X1 U9295 ( .A(n14341), .ZN(n15062) );
  NAND2_X1 U9296 ( .A1(n10550), .A2(n10562), .ZN(n15381) );
  INV_X1 U9297 ( .A(n15381), .ZN(n15390) );
  AND2_X1 U9298 ( .A1(n15519), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n6798) );
  NAND2_X1 U9299 ( .A1(n12092), .A2(n12091), .ZN(n15068) );
  INV_X1 U9300 ( .A(n15068), .ZN(n7041) );
  INV_X1 U9301 ( .A(n9014), .ZN(n7457) );
  INV_X1 U9302 ( .A(n10768), .ZN(n9014) );
  AND2_X1 U9303 ( .A1(n9940), .A2(n9939), .ZN(n6799) );
  NAND2_X1 U9304 ( .A1(n6859), .A2(n11433), .ZN(n11432) );
  AND2_X1 U9305 ( .A1(n10586), .A2(n7772), .ZN(n15406) );
  AND2_X1 U9306 ( .A1(n14200), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n6800) );
  NAND2_X1 U9307 ( .A1(n7033), .A2(n12533), .ZN(n11495) );
  INV_X1 U9308 ( .A(n11495), .ZN(n7032) );
  INV_X1 U9309 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n7305) );
  AND2_X1 U9310 ( .A1(n15557), .A2(n15583), .ZN(n15570) );
  NOR2_X1 U9311 ( .A1(n8353), .A2(n7230), .ZN(n7229) );
  AND2_X1 U9312 ( .A1(n7361), .A2(n7357), .ZN(n6801) );
  INV_X1 U9313 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n7014) );
  INV_X1 U9314 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n7519) );
  INV_X1 U9315 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n7158) );
  INV_X1 U9316 ( .A(n15279), .ZN(n14026) );
  AOI21_X1 U9317 ( .B1(n14105), .B2(n15279), .A(n9716), .ZN(n9717) );
  NOR2_X2 U9318 ( .A1(n10523), .A2(n10046), .ZN(n14379) );
  INV_X1 U9319 ( .A(n9681), .ZN(n9079) );
  NAND3_X1 U9320 ( .A1(n7405), .A2(n9233), .A3(n7414), .ZN(n9681) );
  NAND2_X1 U9321 ( .A1(n12280), .A2(n9744), .ZN(n14081) );
  NOR2_X1 U9322 ( .A1(n6856), .A2(n6855), .ZN(n6854) );
  XNOR2_X1 U9323 ( .A(n13891), .B(n10725), .ZN(n11468) );
  NAND2_X1 U9324 ( .A1(n14173), .A2(n15357), .ZN(n6803) );
  NAND2_X1 U9325 ( .A1(n6803), .A2(n6802), .ZN(P2_U3528) );
  NAND2_X1 U9326 ( .A1(n11169), .A2(n11168), .ZN(n7029) );
  NAND2_X1 U9327 ( .A1(n12053), .A2(n12052), .ZN(n12051) );
  OAI21_X1 U9328 ( .B1(n12128), .B2(n8565), .A(n8861), .ZN(n12204) );
  NAND2_X1 U9329 ( .A1(n11545), .A2(n11544), .ZN(n11936) );
  NAND2_X1 U9330 ( .A1(n6805), .A2(n14957), .ZN(n7117) );
  INV_X1 U9331 ( .A(n13126), .ZN(n6805) );
  OAI21_X1 U9332 ( .B1(n13507), .B2(n13508), .A(n8898), .ZN(n13497) );
  NAND2_X1 U9333 ( .A1(n11301), .A2(n8806), .ZN(n8422) );
  NAND2_X1 U9334 ( .A1(n7641), .A2(n12063), .ZN(n12062) );
  NAND2_X1 U9335 ( .A1(n13991), .A2(n6711), .ZN(n13970) );
  NOR2_X1 U9336 ( .A1(n15610), .A2(n15609), .ZN(n15608) );
  XNOR2_X1 U9337 ( .A(n7902), .B(P2_ADDR_REG_4__SCAN_IN), .ZN(n15610) );
  INV_X1 U9338 ( .A(n7003), .ZN(n14881) );
  INV_X1 U9339 ( .A(n15101), .ZN(n7299) );
  NOR2_X1 U9340 ( .A1(n15098), .A2(n15099), .ZN(n15097) );
  NOR2_X1 U9341 ( .A1(n15082), .A2(n15081), .ZN(n7932) );
  NAND2_X1 U9342 ( .A1(n7905), .A2(n7904), .ZN(n6994) );
  INV_X1 U9343 ( .A(n10930), .ZN(n10931) );
  NAND2_X1 U9344 ( .A1(n13827), .A2(n6759), .ZN(n13722) );
  NAND2_X1 U9345 ( .A1(n6910), .A2(n11015), .ZN(n6909) );
  NAND2_X1 U9346 ( .A1(n6917), .A2(n6915), .ZN(n12151) );
  NAND2_X1 U9347 ( .A1(n9759), .A2(n9758), .ZN(n10724) );
  NAND2_X1 U9348 ( .A1(n6877), .A2(n6876), .ZN(n15371) );
  INV_X1 U9349 ( .A(n8646), .ZN(n8736) );
  NAND2_X1 U9350 ( .A1(n13185), .A2(n13184), .ZN(n13183) );
  NAND2_X1 U9351 ( .A1(n13293), .A2(n13292), .ZN(n13291) );
  NAND2_X1 U9352 ( .A1(n7142), .A2(n7143), .ZN(n12431) );
  NAND2_X1 U9353 ( .A1(n10716), .A2(n10713), .ZN(n10896) );
  AND2_X1 U9354 ( .A1(n10895), .A2(n10710), .ZN(n10716) );
  NAND2_X1 U9355 ( .A1(n15387), .A2(n7147), .ZN(n11184) );
  INV_X1 U9356 ( .A(n7139), .ZN(n7657) );
  NAND2_X1 U9357 ( .A1(n10709), .A2(n6816), .ZN(n6815) );
  INV_X1 U9358 ( .A(n9190), .ZN(n9199) );
  NAND2_X1 U9359 ( .A1(n9184), .A2(n9211), .ZN(n9190) );
  INV_X1 U9360 ( .A(n9626), .ZN(n6807) );
  NAND3_X1 U9361 ( .A1(n7333), .A2(n7332), .A3(n7334), .ZN(n9537) );
  NAND2_X1 U9362 ( .A1(n6808), .A2(n10019), .ZN(P2_U3328) );
  NAND3_X1 U9363 ( .A1(n10016), .A2(n6832), .A3(n6831), .ZN(n6808) );
  NAND2_X1 U9364 ( .A1(n10004), .A2(n10003), .ZN(n10012) );
  NAND2_X1 U9365 ( .A1(n6814), .A2(n6815), .ZN(n10895) );
  OAI21_X1 U9366 ( .B1(n9181), .B2(n10979), .A(n6830), .ZN(n9124) );
  AOI21_X1 U9367 ( .B1(n7289), .B2(n7292), .A(n9991), .ZN(n7286) );
  XNOR2_X1 U9368 ( .A(n7249), .B(n9654), .ZN(n7248) );
  OR2_X1 U9369 ( .A1(n6668), .A2(n10991), .ZN(n10992) );
  NAND2_X2 U9370 ( .A1(n6693), .A2(n10995), .ZN(n14375) );
  NAND2_X1 U9371 ( .A1(n8433), .A2(n8813), .ZN(n11740) );
  AND2_X4 U9372 ( .A1(n13133), .A2(n13685), .ZN(n8764) );
  NAND2_X1 U9373 ( .A1(n10482), .A2(n10481), .ZN(n10832) );
  NAND2_X1 U9374 ( .A1(n12448), .A2(n12613), .ZN(n12450) );
  OAI21_X1 U9375 ( .B1(n11502), .B2(n11361), .A(n11360), .ZN(n11362) );
  NAND2_X1 U9376 ( .A1(n11491), .A2(n7175), .ZN(n6809) );
  NAND2_X1 U9377 ( .A1(n6809), .A2(n11357), .ZN(n11481) );
  AND2_X2 U9378 ( .A1(n13472), .A2(n13471), .ZN(n13474) );
  NAND2_X1 U9379 ( .A1(n8685), .A2(n8907), .ZN(n13472) );
  XNOR2_X1 U9380 ( .A(n7786), .B(n6870), .ZN(n13341) );
  NAND2_X1 U9381 ( .A1(n10712), .A2(n10708), .ZN(n11301) );
  NAND2_X1 U9382 ( .A1(n8485), .A2(n8834), .ZN(n11776) );
  XNOR2_X1 U9383 ( .A(n9125), .B(n9145), .ZN(n10977) );
  NAND2_X1 U9384 ( .A1(n8992), .A2(n8993), .ZN(n8995) );
  NOR2_X2 U9385 ( .A1(n8775), .A2(P3_IR_REG_20__SCAN_IN), .ZN(n7749) );
  OAI22_X2 U9386 ( .A1(n14501), .A2(n12935), .B1(n14830), .B2(n14357), .ZN(
        n13113) );
  NAND2_X1 U9387 ( .A1(n11978), .A2(n7610), .ZN(n12101) );
  NAND2_X1 U9388 ( .A1(n9369), .A2(n7325), .ZN(n9387) );
  NAND2_X1 U9389 ( .A1(n6948), .A2(n6949), .ZN(n9429) );
  NAND2_X1 U9390 ( .A1(n6775), .A2(n6900), .ZN(n6898) );
  NAND2_X1 U9391 ( .A1(n9571), .A2(n7335), .ZN(n9572) );
  INV_X1 U9392 ( .A(n7336), .ZN(n7335) );
  NAND2_X1 U9393 ( .A1(n9274), .A2(n9273), .ZN(n9291) );
  NAND2_X1 U9394 ( .A1(n6886), .A2(n6885), .ZN(n7333) );
  INV_X1 U9395 ( .A(n6969), .ZN(n6968) );
  AND2_X1 U9396 ( .A1(n11733), .A2(n15111), .ZN(n6821) );
  NOR2_X1 U9397 ( .A1(n9145), .A2(n9144), .ZN(n9146) );
  NAND2_X1 U9398 ( .A1(n7115), .A2(n7116), .ZN(n9032) );
  NAND2_X1 U9399 ( .A1(n8579), .A2(n8867), .ZN(n12328) );
  NAND2_X1 U9400 ( .A1(n12051), .A2(n8843), .ZN(n12042) );
  NAND2_X1 U9401 ( .A1(n11936), .A2(n11935), .ZN(n8484) );
  NAND2_X1 U9402 ( .A1(n8631), .A2(n13528), .ZN(n13545) );
  XNOR2_X1 U9403 ( .A(n8951), .B(n6756), .ZN(n13126) );
  NAND2_X2 U9404 ( .A1(n11689), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10635) );
  NAND2_X1 U9405 ( .A1(n6882), .A2(n7219), .ZN(n14608) );
  NAND2_X1 U9406 ( .A1(n14659), .A2(n12899), .ZN(n14641) );
  NAND2_X1 U9407 ( .A1(n12255), .A2(n12254), .ZN(n12300) );
  NAND2_X1 U9408 ( .A1(n11840), .A2(n11839), .ZN(n11841) );
  NAND2_X1 U9409 ( .A1(n6823), .A2(n7607), .ZN(n11977) );
  INV_X1 U9410 ( .A(n11841), .ZN(n6823) );
  NAND2_X1 U9411 ( .A1(n7204), .A2(n6766), .ZN(n14659) );
  NAND2_X1 U9412 ( .A1(n6824), .A2(n8938), .ZN(n8943) );
  NAND2_X1 U9413 ( .A1(n6833), .A2(n6729), .ZN(n6824) );
  NAND2_X1 U9414 ( .A1(n14641), .A2(n6675), .ZN(n6882) );
  OAI22_X1 U9415 ( .A1(n11437), .A2(n12839), .B1(n12533), .B2(n14377), .ZN(
        n11491) );
  AOI22_X1 U9416 ( .A1(n6669), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n10062), .B2(
        n10184), .ZN(n9129) );
  NAND2_X1 U9417 ( .A1(n9733), .A2(n9732), .ZN(n11169) );
  BUF_X1 U9418 ( .A(n11468), .Z(n6826) );
  NAND2_X1 U9419 ( .A1(n13927), .A2(n9642), .ZN(n7249) );
  NAND2_X1 U9420 ( .A1(n7287), .A2(n7286), .ZN(n13925) );
  NAND2_X1 U9421 ( .A1(n10014), .A2(n10015), .ZN(n6831) );
  INV_X1 U9422 ( .A(n10013), .ZN(n6832) );
  NAND2_X1 U9423 ( .A1(n9355), .A2(n7326), .ZN(n7325) );
  NAND2_X1 U9424 ( .A1(n9252), .A2(n9251), .ZN(n9272) );
  NAND2_X1 U9425 ( .A1(n9537), .A2(n7334), .ZN(n9557) );
  NOR2_X1 U9426 ( .A1(n13336), .A2(n13335), .ZN(n13334) );
  OAI21_X1 U9427 ( .B1(n14924), .B2(n15530), .A(n7169), .ZN(P3_U3200) );
  NOR2_X1 U9428 ( .A1(n11159), .A2(n11160), .ZN(n11158) );
  NAND2_X2 U9429 ( .A1(n7666), .A2(n7651), .ZN(n8775) );
  NAND2_X1 U9430 ( .A1(n8567), .A2(n8566), .ZN(n8569) );
  NAND2_X1 U9431 ( .A1(n8925), .A2(n8926), .ZN(n8923) );
  NAND2_X1 U9432 ( .A1(n8921), .A2(n8920), .ZN(n8925) );
  NAND2_X1 U9433 ( .A1(n8620), .A2(n8619), .ZN(n8622) );
  NAND2_X1 U9434 ( .A1(n8608), .A2(n8607), .ZN(n8610) );
  NAND2_X1 U9435 ( .A1(n7211), .A2(n8325), .ZN(n8556) );
  NAND2_X1 U9436 ( .A1(n6835), .A2(n6834), .ZN(n6833) );
  AOI21_X2 U9437 ( .B1(n6836), .B2(n8935), .A(n8934), .ZN(n8936) );
  NAND3_X1 U9438 ( .A1(n8933), .A2(n8931), .A3(n8932), .ZN(n6836) );
  OR2_X1 U9439 ( .A1(n7750), .A2(n7715), .ZN(n6892) );
  NAND2_X1 U9440 ( .A1(n8553), .A2(n8855), .ZN(n12128) );
  NAND2_X1 U9441 ( .A1(n8499), .A2(n8839), .ZN(n11526) );
  NAND2_X1 U9442 ( .A1(n7427), .A2(n7426), .ZN(n13547) );
  NAND2_X2 U9443 ( .A1(n11871), .A2(n11870), .ZN(n12075) );
  NAND2_X1 U9444 ( .A1(n6842), .A2(n6840), .ZN(P1_U3214) );
  NAND2_X1 U9445 ( .A1(n14207), .A2(n14341), .ZN(n6842) );
  AOI22_X2 U9446 ( .A1(n11864), .A2(n11863), .B1(n11862), .B2(n11861), .ZN(
        n14320) );
  OAI21_X1 U9447 ( .B1(n14292), .B2(n7340), .A(n7338), .ZN(n12978) );
  NAND2_X1 U9448 ( .A1(n7343), .A2(n7341), .ZN(n14246) );
  INV_X1 U9449 ( .A(n12204), .ZN(n8578) );
  INV_X1 U9450 ( .A(n11526), .ZN(n6847) );
  NAND2_X1 U9451 ( .A1(n12431), .A2(n12430), .ZN(n12435) );
  NAND2_X1 U9452 ( .A1(n13244), .A2(n13146), .ZN(n13255) );
  NAND2_X1 U9453 ( .A1(n13183), .A2(n13139), .ZN(n13311) );
  NAND2_X1 U9454 ( .A1(n13253), .A2(n13148), .ZN(n13293) );
  NAND2_X1 U9455 ( .A1(n13246), .A2(n13245), .ZN(n13244) );
  OAI21_X4 U9456 ( .B1(n10703), .B2(n10702), .A(n10707), .ZN(n11713) );
  XNOR2_X1 U9457 ( .A(n6843), .B(n13217), .ZN(n13225) );
  OAI21_X1 U9458 ( .B1(n13214), .B2(n13213), .A(n6844), .ZN(n6843) );
  NAND2_X1 U9459 ( .A1(n12222), .A2(n12221), .ZN(n15373) );
  NOR2_X1 U9460 ( .A1(n11896), .A2(n6888), .ZN(n15506) );
  OAI21_X1 U9462 ( .B1(n7637), .B2(n7858), .A(n7857), .ZN(n7859) );
  NOR2_X1 U9463 ( .A1(n11897), .A2(n11898), .ZN(n11896) );
  NAND2_X1 U9464 ( .A1(n9354), .A2(SI_14_), .ZN(n9355) );
  NAND2_X1 U9465 ( .A1(n9950), .A2(n9949), .ZN(n9952) );
  INV_X1 U9466 ( .A(n9943), .ZN(n6878) );
  INV_X1 U9467 ( .A(n9959), .ZN(n9997) );
  OAI21_X1 U9468 ( .B1(n10012), .B2(n7330), .A(n7329), .ZN(n10013) );
  INV_X1 U9469 ( .A(n9103), .ZN(n7388) );
  NAND2_X1 U9470 ( .A1(n9588), .A2(n9587), .ZN(n9592) );
  OAI21_X1 U9471 ( .B1(n9181), .B2(n8404), .A(n6848), .ZN(n9092) );
  AOI21_X2 U9472 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n15483), .A(n15473), .ZN(
        n7728) );
  NOR2_X2 U9473 ( .A1(n13365), .A2(n6869), .ZN(n7742) );
  NAND2_X1 U9474 ( .A1(n9518), .A2(n9517), .ZN(n9519) );
  NOR2_X1 U9475 ( .A1(n15423), .A2(n15424), .ZN(n15422) );
  NAND2_X1 U9476 ( .A1(n7460), .A2(n7459), .ZN(n7458) );
  AOI21_X1 U9477 ( .B1(n14496), .B2(n14497), .A(n14781), .ZN(n6850) );
  XNOR2_X1 U9478 ( .A(n7783), .B(n11906), .ZN(n11902) );
  INV_X1 U9479 ( .A(n6940), .ZN(n14918) );
  NOR2_X1 U9480 ( .A1(n10573), .A2(n10574), .ZN(n10572) );
  INV_X1 U9481 ( .A(n7170), .ZN(n7169) );
  NAND2_X1 U9482 ( .A1(n11023), .A2(n11022), .ZN(n9731) );
  OR2_X1 U9483 ( .A1(n9105), .A2(n10615), .ZN(n7051) );
  OAI21_X1 U9484 ( .B1(n6670), .B2(n6853), .A(n6852), .ZN(n9091) );
  NAND2_X1 U9485 ( .A1(n7390), .A2(n7389), .ZN(n9104) );
  NAND3_X2 U9486 ( .A1(n6706), .A2(n9074), .A3(n9073), .ZN(n13891) );
  NAND2_X1 U9487 ( .A1(n7729), .A2(n7167), .ZN(n7165) );
  NAND2_X1 U9488 ( .A1(n7732), .A2(n7156), .ZN(n7154) );
  INV_X1 U9489 ( .A(n9519), .ZN(n6886) );
  OAI211_X1 U9490 ( .C1(n12877), .C2(n6963), .A(n12876), .B(n6962), .ZN(n12878) );
  NAND4_X4 U9491 ( .A1(n10636), .A2(n10635), .A3(n10634), .A4(n10633), .ZN(
        n14377) );
  CLKBUF_X1 U9492 ( .A(n12839), .Z(n6859) );
  INV_X1 U9493 ( .A(n10028), .ZN(n7241) );
  OAI21_X1 U9494 ( .B1(n13113), .B2(n13112), .A(n6883), .ZN(n13115) );
  INV_X1 U9495 ( .A(n12951), .ZN(n10482) );
  NAND2_X1 U9496 ( .A1(n11393), .A2(n11392), .ZN(n11682) );
  NOR2_X2 U9497 ( .A1(n10211), .A2(P1_IR_REG_28__SCAN_IN), .ZN(n10478) );
  OAI211_X2 U9498 ( .C1(n12738), .C2(n11224), .A(n11223), .B(n11222), .ZN(
        n12555) );
  NAND2_X2 U9500 ( .A1(n7030), .A2(n6865), .ZN(n12530) );
  NAND2_X1 U9501 ( .A1(n11288), .A2(n11289), .ZN(n9726) );
  NAND2_X1 U9502 ( .A1(n9724), .A2(n9723), .ZN(n11288) );
  NAND2_X1 U9503 ( .A1(n9082), .A2(n9069), .ZN(n9084) );
  NAND2_X1 U9504 ( .A1(n14173), .A2(n15347), .ZN(n7024) );
  NAND2_X1 U9505 ( .A1(n7025), .A2(n7402), .ZN(n14046) );
  BUF_X2 U9506 ( .A(n7666), .Z(n7667) );
  INV_X1 U9507 ( .A(n6874), .ZN(n7672) );
  INV_X1 U9508 ( .A(n15373), .ZN(n6877) );
  INV_X1 U9509 ( .A(n15382), .ZN(n7148) );
  NAND2_X1 U9510 ( .A1(n6887), .A2(n6689), .ZN(n7142) );
  NAND2_X1 U9511 ( .A1(n6875), .A2(n11089), .ZN(n15383) );
  NAND2_X1 U9512 ( .A1(n11086), .A2(n11087), .ZN(n6875) );
  NAND2_X1 U9513 ( .A1(n7149), .A2(n7148), .ZN(n15387) );
  INV_X1 U9514 ( .A(n12228), .ZN(n6887) );
  OR2_X2 U9515 ( .A1(n10015), .A2(n10012), .ZN(n10016) );
  NAND2_X1 U9516 ( .A1(n9506), .A2(n9505), .ZN(n9518) );
  AND4_X2 U9517 ( .A1(n7645), .A2(n7646), .A3(n7497), .A4(n7647), .ZN(n7104)
         );
  NAND2_X1 U9518 ( .A1(n6892), .A2(P3_IR_REG_28__SCAN_IN), .ZN(n6891) );
  NAND2_X1 U9519 ( .A1(n8422), .A2(n8812), .ZN(n11750) );
  INV_X1 U9520 ( .A(n10760), .ZN(n10025) );
  AND2_X4 U9521 ( .A1(n10481), .A2(n12951), .ZN(n12702) );
  NAND2_X1 U9522 ( .A1(n9231), .A2(n9230), .ZN(n9250) );
  NAND2_X1 U9523 ( .A1(n9146), .A2(n7015), .ZN(n7018) );
  INV_X1 U9524 ( .A(n7031), .ZN(n7030) );
  NAND2_X1 U9525 ( .A1(n7243), .A2(n10029), .ZN(n10209) );
  NAND2_X1 U9526 ( .A1(n10209), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10210) );
  INV_X2 U9527 ( .A(n11713), .ZN(n13174) );
  NAND2_X1 U9528 ( .A1(n12007), .A2(n6768), .ZN(n12222) );
  INV_X1 U9529 ( .A(n15383), .ZN(n7149) );
  XNOR2_X1 U9530 ( .A(n12892), .B(P3_B_REG_SCAN_IN), .ZN(n8991) );
  XNOR2_X2 U9531 ( .A(n15314), .B(n13889), .ZN(n11290) );
  NAND2_X1 U9532 ( .A1(n14081), .A2(n7404), .ZN(n7025) );
  NAND2_X1 U9533 ( .A1(n6893), .A2(n10904), .ZN(n13751) );
  NAND2_X1 U9534 ( .A1(n10743), .A2(n10744), .ZN(n13749) );
  NAND2_X1 U9535 ( .A1(n6896), .A2(n7535), .ZN(n6895) );
  OAI211_X1 U9536 ( .C1(n7535), .C2(n6897), .A(n6895), .B(n13778), .ZN(
        P2_U3192) );
  NAND2_X1 U9537 ( .A1(n7535), .A2(n7534), .ZN(n13768) );
  INV_X1 U9538 ( .A(n7546), .ZN(n6910) );
  NAND2_X1 U9539 ( .A1(n11197), .A2(n11196), .ZN(n11206) );
  NAND2_X1 U9540 ( .A1(n11673), .A2(n6918), .ZN(n6917) );
  INV_X1 U9541 ( .A(n13802), .ZN(n6922) );
  INV_X1 U9542 ( .A(n9410), .ZN(n6930) );
  CLKBUF_X1 U9543 ( .A(n7414), .Z(n6928) );
  NAND4_X1 U9544 ( .A1(n6700), .A2(n9109), .A3(n6930), .A4(n6929), .ZN(n9655)
         );
  NAND2_X1 U9545 ( .A1(n9234), .A2(n6928), .ZN(n9437) );
  NOR2_X2 U9546 ( .A1(n9410), .A2(n9060), .ZN(n7414) );
  NAND2_X1 U9547 ( .A1(n6940), .A2(n7508), .ZN(n7507) );
  NAND2_X1 U9548 ( .A1(n7318), .A2(n7320), .ZN(n9353) );
  NAND2_X1 U9549 ( .A1(n7589), .A2(n6943), .ZN(n6942) );
  NAND3_X1 U9550 ( .A1(n6942), .A2(n6945), .A3(n7582), .ZN(n7581) );
  INV_X1 U9551 ( .A(n6946), .ZN(n6944) );
  NAND2_X1 U9552 ( .A1(n9387), .A2(n6952), .ZN(n6948) );
  NAND2_X1 U9553 ( .A1(n6955), .A2(n9453), .ZN(n9454) );
  NAND2_X1 U9554 ( .A1(n9453), .A2(n9434), .ZN(n9435) );
  NAND3_X1 U9555 ( .A1(n9453), .A2(n6957), .A3(n6960), .ZN(n6956) );
  OAI21_X1 U9556 ( .B1(n12741), .B2(n7579), .A(n7576), .ZN(n12744) );
  OAI22_X1 U9557 ( .A1(n12727), .A2(n6686), .B1(n12728), .B2(n6961), .ZN(
        n12741) );
  INV_X1 U9558 ( .A(n12726), .ZN(n6961) );
  OAI21_X2 U9559 ( .B1(n12836), .B2(n7639), .A(n6747), .ZN(n6963) );
  NAND2_X1 U9560 ( .A1(n9147), .A2(SI_2_), .ZN(n9122) );
  NAND2_X1 U9561 ( .A1(n6964), .A2(n7389), .ZN(n9147) );
  NAND3_X1 U9562 ( .A1(n7388), .A2(n7389), .A3(n7390), .ZN(n6964) );
  NAND2_X1 U9563 ( .A1(n9090), .A2(n10159), .ZN(n7390) );
  NAND2_X1 U9564 ( .A1(n9091), .A2(SI_1_), .ZN(n7389) );
  OR2_X1 U9565 ( .A1(n14566), .A2(n6968), .ZN(n6965) );
  NAND2_X1 U9566 ( .A1(n6965), .A2(n6967), .ZN(n14516) );
  INV_X1 U9567 ( .A(n6972), .ZN(n14586) );
  OAI21_X1 U9568 ( .B1(n12925), .B2(n6975), .A(n6696), .ZN(n14588) );
  INV_X1 U9569 ( .A(n11833), .ZN(n6977) );
  OAI21_X1 U9570 ( .B1(n6977), .B2(n6979), .A(n6978), .ZN(n12166) );
  INV_X1 U9571 ( .A(n12914), .ZN(n6983) );
  OAI21_X1 U9572 ( .B1(n6983), .B2(n6987), .A(n6674), .ZN(n7599) );
  NAND2_X2 U9573 ( .A1(n6990), .A2(n10824), .ZN(n11434) );
  INV_X1 U9574 ( .A(n6991), .ZN(n6990) );
  XNOR2_X1 U9575 ( .A(n7307), .B(n7306), .ZN(SUB_1596_U4) );
  INV_X1 U9576 ( .A(n7000), .ZN(n7004) );
  OR2_X1 U9577 ( .A1(n7000), .A2(n14915), .ZN(n7952) );
  NAND3_X1 U9578 ( .A1(n7009), .A2(n7007), .A3(n7010), .ZN(n15082) );
  NAND3_X1 U9579 ( .A1(n6681), .A2(n14901), .A3(n7012), .ZN(n7009) );
  NAND3_X1 U9580 ( .A1(n7017), .A2(n7389), .A3(n7016), .ZN(n7015) );
  NAND2_X1 U9581 ( .A1(n7018), .A2(n9148), .ZN(n9161) );
  NAND2_X1 U9582 ( .A1(n7024), .A2(n7022), .ZN(P2_U3496) );
  OR2_X1 U9583 ( .A1(n15347), .A2(n7023), .ZN(n7022) );
  XNOR2_X1 U9584 ( .A(n9755), .B(n9995), .ZN(n14109) );
  OR2_X1 U9585 ( .A1(n11338), .A2(n9523), .ZN(n9202) );
  OAI22_X1 U9586 ( .A1(n10978), .A2(n6853), .B1(n14387), .B2(n12738), .ZN(
        n7031) );
  NAND2_X1 U9587 ( .A1(n12462), .A2(n6761), .ZN(n7035) );
  INV_X1 U9588 ( .A(n7035), .ZN(n14682) );
  NOR2_X1 U9589 ( .A1(n14509), .A2(n7039), .ZN(n14495) );
  NAND2_X1 U9590 ( .A1(n11702), .A2(n7040), .ZN(n12187) );
  NAND2_X1 U9591 ( .A1(n14589), .A2(n6762), .ZN(n14517) );
  INV_X1 U9592 ( .A(n7048), .ZN(n14553) );
  NOR2_X2 U9593 ( .A1(n11140), .A2(n11141), .ZN(n11139) );
  NAND2_X1 U9594 ( .A1(n7050), .A2(n7049), .ZN(n11140) );
  NOR3_X4 U9595 ( .A1(n14036), .A2(n7053), .A3(n14126), .ZN(n13976) );
  NOR2_X2 U9596 ( .A1(n13932), .A2(n14106), .ZN(n13918) );
  NOR3_X2 U9597 ( .A1(n11885), .A2(n14975), .A3(n7060), .ZN(n7061) );
  INV_X1 U9598 ( .A(n7061), .ZN(n14981) );
  NAND2_X1 U9599 ( .A1(n12046), .A2(n7079), .ZN(n7077) );
  NAND2_X1 U9600 ( .A1(n8983), .A2(n7083), .ZN(n7086) );
  NAND2_X1 U9601 ( .A1(n8983), .A2(n7087), .ZN(n13416) );
  INV_X1 U9602 ( .A(n7086), .ZN(n13415) );
  NAND2_X1 U9603 ( .A1(n13481), .A2(n7092), .ZN(n7089) );
  NAND2_X1 U9604 ( .A1(n7089), .A2(n7090), .ZN(n13444) );
  NAND4_X1 U9605 ( .A1(n7654), .A2(n7140), .A3(n7653), .A4(n7664), .ZN(n7747)
         );
  AND3_X2 U9606 ( .A1(n7104), .A2(n7644), .A3(n7687), .ZN(n7666) );
  AND2_X2 U9607 ( .A1(n7709), .A2(n7711), .ZN(n7687) );
  AND2_X1 U9608 ( .A1(n7116), .A2(n7118), .ZN(n13129) );
  OR2_X1 U9609 ( .A1(n6879), .A2(n10160), .ZN(n7119) );
  NAND2_X4 U9610 ( .A1(n8361), .A2(n9213), .ZN(n8761) );
  NAND3_X1 U9611 ( .A1(n11540), .A2(n8964), .A3(n8963), .ZN(n11770) );
  NAND2_X1 U9612 ( .A1(n11711), .A2(n7123), .ZN(n7121) );
  NAND2_X1 U9613 ( .A1(n7121), .A2(n7122), .ZN(n15358) );
  NAND2_X1 U9614 ( .A1(n13263), .A2(n6772), .ZN(n7128) );
  OAI211_X1 U9615 ( .C1(n13263), .C2(n7129), .A(n7128), .B(n13273), .ZN(
        P3_U3169) );
  XNOR2_X1 U9616 ( .A(n13263), .B(n13198), .ZN(n13264) );
  OAI21_X2 U9617 ( .B1(n8995), .B2(P3_D_REG_0__SCAN_IN), .A(n8994), .ZN(n10703) );
  INV_X1 U9618 ( .A(n7720), .ZN(n7159) );
  INV_X1 U9619 ( .A(n7161), .ZN(n15403) );
  NAND2_X1 U9620 ( .A1(n7743), .A2(n7164), .ZN(n7162) );
  XNOR2_X2 U9621 ( .A(n7742), .B(n13397), .ZN(n13385) );
  OAI21_X1 U9622 ( .B1(n11045), .B2(n7166), .A(n7165), .ZN(n11154) );
  CLKBUF_X1 U9623 ( .A(n7175), .Z(n7174) );
  NAND3_X1 U9624 ( .A1(n12549), .A2(n12550), .A3(n7174), .ZN(n12553) );
  NAND3_X1 U9625 ( .A1(n12842), .A2(n12841), .A3(n7174), .ZN(n12846) );
  NAND2_X1 U9626 ( .A1(n10980), .A2(n7176), .ZN(n10988) );
  NOR2_X1 U9627 ( .A1(n12738), .A2(n14402), .ZN(n7177) );
  NAND2_X1 U9628 ( .A1(n8581), .A2(n7181), .ZN(n7180) );
  NAND2_X1 U9629 ( .A1(n8523), .A2(n7187), .ZN(n7186) );
  INV_X1 U9630 ( .A(n7192), .ZN(n7191) );
  OAI21_X1 U9631 ( .B1(n8936), .B2(n11314), .A(n7193), .ZN(n7192) );
  NAND2_X1 U9632 ( .A1(n8936), .A2(n8939), .ZN(n7193) );
  NAND2_X1 U9633 ( .A1(n7195), .A2(n8937), .ZN(n7194) );
  XNOR2_X1 U9634 ( .A(n8794), .B(n7457), .ZN(n7195) );
  INV_X1 U9635 ( .A(n8635), .ZN(n7196) );
  NAND2_X1 U9636 ( .A1(n7196), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n7198) );
  NAND3_X1 U9637 ( .A1(n7202), .A2(n7200), .A3(n7198), .ZN(n8649) );
  NAND2_X2 U9638 ( .A1(n12450), .A2(n12915), .ZN(n12894) );
  NAND2_X1 U9639 ( .A1(n8556), .A2(n8326), .ZN(n8567) );
  NAND2_X1 U9640 ( .A1(n11682), .A2(n6767), .ZN(n11840) );
  NAND2_X1 U9641 ( .A1(n8440), .A2(n7216), .ZN(n7212) );
  NAND2_X1 U9642 ( .A1(n8731), .A2(n7229), .ZN(n7227) );
  OAI21_X1 U9643 ( .B1(n8674), .B2(n7234), .A(n7232), .ZN(n8343) );
  OAI21_X1 U9644 ( .B1(n8674), .B2(n8673), .A(n8342), .ZN(n8687) );
  NOR2_X2 U9645 ( .A1(n10119), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n10135) );
  INV_X1 U9646 ( .A(n7245), .ZN(n7244) );
  OAI21_X1 U9647 ( .B1(n8698), .B2(P2_DATAO_REG_24__SCAN_IN), .A(n8345), .ZN(
        n8709) );
  NAND2_X2 U9648 ( .A1(n14608), .A2(n14609), .ZN(n14579) );
  NOR2_X1 U9649 ( .A1(n13333), .A2(n13332), .ZN(n13331) );
  NOR2_X1 U9650 ( .A1(n10570), .A2(n10569), .ZN(n10568) );
  AOI21_X1 U9651 ( .B1(P3_REG2_REG_0__SCAN_IN), .B2(n7709), .A(n10597), .ZN(
        n10570) );
  CLKBUF_X1 U9652 ( .A(n7251), .Z(n7250) );
  NAND2_X1 U9653 ( .A1(n10977), .A2(n7251), .ZN(n9130) );
  NAND2_X1 U9654 ( .A1(n11325), .A2(n7251), .ZN(n9170) );
  NAND2_X1 U9655 ( .A1(n11378), .A2(n7251), .ZN(n9218) );
  NAND2_X1 U9656 ( .A1(n11683), .A2(n7251), .ZN(n9237) );
  NAND2_X1 U9657 ( .A1(n11834), .A2(n7250), .ZN(n9259) );
  NAND2_X1 U9658 ( .A1(n11973), .A2(n7250), .ZN(n9278) );
  NAND2_X1 U9659 ( .A1(n12089), .A2(n7250), .ZN(n9296) );
  NAND2_X1 U9660 ( .A1(n12167), .A2(n7250), .ZN(n9317) );
  NAND2_X1 U9661 ( .A1(n12239), .A2(n7250), .ZN(n9338) );
  NAND2_X1 U9662 ( .A1(n12292), .A2(n7250), .ZN(n9360) );
  NAND2_X1 U9663 ( .A1(n12443), .A2(n7250), .ZN(n9378) );
  NAND2_X1 U9664 ( .A1(n12627), .A2(n7250), .ZN(n9397) );
  NAND2_X1 U9665 ( .A1(n12638), .A2(n7250), .ZN(n9414) );
  NAND2_X1 U9666 ( .A1(n12649), .A2(n7250), .ZN(n9458) );
  NAND2_X1 U9667 ( .A1(n12524), .A2(n7250), .ZN(n9540) );
  NAND2_X1 U9668 ( .A1(n12746), .A2(n7250), .ZN(n9564) );
  NAND2_X1 U9669 ( .A1(n12771), .A2(n7250), .ZN(n9574) );
  NAND2_X1 U9670 ( .A1(n12792), .A2(n7250), .ZN(n9595) );
  NAND2_X1 U9671 ( .A1(n12887), .A2(n7250), .ZN(n9611) );
  NAND2_X1 U9672 ( .A1(n14869), .A2(n7250), .ZN(n9629) );
  NAND2_X1 U9673 ( .A1(n12949), .A2(n7250), .ZN(n7331) );
  NAND2_X1 U9674 ( .A1(n12885), .A2(n7250), .ZN(n9922) );
  NAND2_X1 U9675 ( .A1(n14186), .A2(n7250), .ZN(n9950) );
  NAND2_X1 U9676 ( .A1(n10947), .A2(n7253), .ZN(n7252) );
  NAND2_X1 U9677 ( .A1(n7252), .A2(n7254), .ZN(n11074) );
  NAND2_X1 U9678 ( .A1(n7258), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9083) );
  NAND3_X1 U9679 ( .A1(n7414), .A2(n9233), .A3(n7257), .ZN(n7258) );
  NAND2_X1 U9680 ( .A1(n12282), .A2(n7261), .ZN(n7259) );
  NAND2_X1 U9681 ( .A1(n14053), .A2(n7267), .ZN(n7266) );
  OAI21_X2 U9682 ( .B1(n11879), .B2(n7277), .A(n7276), .ZN(n14970) );
  NAND2_X1 U9683 ( .A1(n13982), .A2(n7289), .ZN(n7287) );
  NAND2_X1 U9684 ( .A1(n13982), .A2(n7294), .ZN(n7288) );
  NAND2_X1 U9685 ( .A1(n7311), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n8360) );
  NAND3_X1 U9686 ( .A1(n8356), .A2(n8355), .A3(n14886), .ZN(n7311) );
  NAND2_X1 U9687 ( .A1(n9433), .A2(n7314), .ZN(n7312) );
  NAND2_X1 U9688 ( .A1(n7312), .A2(n7313), .ZN(n9506) );
  NAND2_X1 U9689 ( .A1(n9293), .A2(n7319), .ZN(n7318) );
  NAND2_X1 U9690 ( .A1(n9626), .A2(SI_27_), .ZN(n9625) );
  NAND2_X1 U9691 ( .A1(n9519), .A2(SI_22_), .ZN(n7334) );
  NAND2_X1 U9692 ( .A1(n7333), .A2(n7334), .ZN(n12736) );
  NAND2_X1 U9693 ( .A1(n14218), .A2(n7345), .ZN(n7343) );
  NAND2_X1 U9694 ( .A1(n14224), .A2(n7352), .ZN(n7351) );
  XNOR2_X1 U9695 ( .A(n7356), .B(n10976), .ZN(n10829) );
  INV_X1 U9696 ( .A(n10975), .ZN(n7356) );
  NAND2_X1 U9697 ( .A1(n7360), .A2(n10829), .ZN(n7358) );
  INV_X1 U9698 ( .A(n7361), .ZN(n10830) );
  NAND2_X1 U9699 ( .A1(n15063), .A2(n7362), .ZN(n12955) );
  INV_X2 U9700 ( .A(n12974), .ZN(n13059) );
  NAND2_X1 U9701 ( .A1(n14204), .A2(n7367), .ZN(n7366) );
  OAI211_X1 U9702 ( .C1(n14204), .C2(n7368), .A(n7366), .B(n13097), .ZN(
        P1_U3220) );
  NOR2_X1 U9703 ( .A1(n13091), .A2(n13084), .ZN(n7372) );
  NAND2_X1 U9704 ( .A1(n13091), .A2(n13084), .ZN(n7373) );
  OAI21_X2 U9705 ( .B1(n12075), .B2(n6680), .A(n7378), .ZN(n12273) );
  OAI21_X1 U9706 ( .B1(n14257), .B2(n7385), .A(n7382), .ZN(n14310) );
  NAND2_X1 U9707 ( .A1(n12062), .A2(n7401), .ZN(n14976) );
  NOR2_X1 U9708 ( .A1(n9077), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n7405) );
  INV_X2 U9709 ( .A(n15271), .ZN(n15306) );
  NAND2_X1 U9710 ( .A1(n7411), .A2(n7407), .ZN(n13991) );
  NAND2_X1 U9711 ( .A1(n14014), .A2(n9753), .ZN(n13997) );
  INV_X1 U9712 ( .A(n7411), .ZN(n13996) );
  INV_X1 U9713 ( .A(n9753), .ZN(n7413) );
  NAND2_X1 U9714 ( .A1(n7417), .A2(n7415), .ZN(n9769) );
  NAND2_X1 U9715 ( .A1(n7416), .A2(n11474), .ZN(n7415) );
  NAND2_X1 U9716 ( .A1(n7418), .A2(n9766), .ZN(n7417) );
  OAI211_X1 U9717 ( .C1(n9763), .C2(n10691), .A(n7420), .B(n7419), .ZN(n7418)
         );
  NAND2_X1 U9718 ( .A1(n9764), .A2(n10691), .ZN(n7420) );
  NAND2_X1 U9719 ( .A1(n7423), .A2(n7422), .ZN(n9814) );
  INV_X1 U9720 ( .A(n9809), .ZN(n7425) );
  NAND2_X1 U9721 ( .A1(n12371), .A2(n7428), .ZN(n7427) );
  INV_X1 U9722 ( .A(n9906), .ZN(n7439) );
  NAND2_X1 U9723 ( .A1(n7440), .A2(n6774), .ZN(n9803) );
  NAND3_X1 U9724 ( .A1(n7443), .A2(n7442), .A3(n7441), .ZN(n7440) );
  OR2_X1 U9725 ( .A1(n9801), .A2(n9802), .ZN(n7441) );
  NAND2_X1 U9726 ( .A1(n9798), .A2(n9797), .ZN(n7442) );
  NAND2_X1 U9727 ( .A1(n9800), .A2(n9799), .ZN(n7443) );
  OAI21_X2 U9728 ( .B1(n6704), .B2(n7447), .A(n7446), .ZN(n9889) );
  AND2_X2 U9729 ( .A1(n14194), .A2(n13121), .ZN(n9599) );
  OAI21_X1 U9730 ( .B1(n8951), .B2(n7462), .A(n7461), .ZN(n7460) );
  NAND2_X1 U9731 ( .A1(n13474), .A2(n7467), .ZN(n7463) );
  NAND2_X1 U9732 ( .A1(n7463), .A2(n7465), .ZN(n13423) );
  NAND2_X1 U9733 ( .A1(n13545), .A2(n6731), .ZN(n8648) );
  NAND2_X1 U9734 ( .A1(n7472), .A2(n7473), .ZN(n9867) );
  NAND3_X1 U9735 ( .A1(n9836), .A2(n6718), .A3(n7475), .ZN(n7472) );
  AOI21_X1 U9736 ( .B1(n9871), .B2(n7485), .A(n7482), .ZN(n9879) );
  NAND4_X1 U9737 ( .A1(n7645), .A2(n7644), .A3(n7687), .A4(n7496), .ZN(n7680)
         );
  NAND4_X1 U9738 ( .A1(n7645), .A2(n7644), .A3(n7687), .A4(n7646), .ZN(n7684)
         );
  NAND2_X1 U9739 ( .A1(n7498), .A2(n6760), .ZN(n8527) );
  NAND3_X1 U9740 ( .A1(n9823), .A2(n9822), .A3(n6787), .ZN(n7499) );
  NAND2_X1 U9741 ( .A1(n7499), .A2(n7500), .ZN(n9830) );
  NOR2_X2 U9742 ( .A1(n8775), .A2(n7503), .ZN(n7750) );
  OAI21_X1 U9743 ( .B1(n11902), .B2(n7510), .A(n7509), .ZN(n15496) );
  OAI21_X1 U9744 ( .B1(n10587), .B2(n7518), .A(n7517), .ZN(n7521) );
  INV_X1 U9745 ( .A(n7772), .ZN(n7518) );
  INV_X1 U9746 ( .A(n7521), .ZN(n15407) );
  XNOR2_X2 U9747 ( .A(n7523), .B(n14187), .ZN(n13121) );
  NAND2_X1 U9748 ( .A1(n13814), .A2(n7536), .ZN(n7535) );
  NAND2_X1 U9749 ( .A1(n13814), .A2(n7542), .ZN(n7540) );
  NAND2_X1 U9750 ( .A1(n11203), .A2(n6688), .ZN(n7549) );
  INV_X1 U9751 ( .A(n7549), .ZN(n11450) );
  INV_X1 U9752 ( .A(n12761), .ZN(n7552) );
  OAI21_X1 U9753 ( .B1(n7552), .B2(n7554), .A(n7553), .ZN(n12776) );
  OAI21_X1 U9754 ( .B1(n12761), .B2(n6678), .A(n7556), .ZN(n12777) );
  NAND2_X1 U9755 ( .A1(n7558), .A2(n7561), .ZN(n12595) );
  NAND3_X1 U9756 ( .A1(n12588), .A2(n7559), .A3(n12587), .ZN(n7558) );
  NAND2_X1 U9757 ( .A1(n12553), .A2(n6771), .ZN(n12558) );
  NAND2_X1 U9758 ( .A1(n7563), .A2(n12556), .ZN(n12560) );
  NAND2_X1 U9759 ( .A1(n7564), .A2(n12553), .ZN(n7563) );
  NAND2_X1 U9760 ( .A1(n12607), .A2(n7568), .ZN(n7567) );
  OAI21_X1 U9761 ( .B1(n7567), .B2(n6751), .A(n7569), .ZN(n12623) );
  NAND2_X1 U9762 ( .A1(n7581), .A2(n7584), .ZN(n12830) );
  NAND2_X1 U9763 ( .A1(n7585), .A2(n7587), .ZN(n12583) );
  NAND3_X1 U9764 ( .A1(n12576), .A2(n7586), .A3(n12575), .ZN(n7585) );
  NAND3_X1 U9765 ( .A1(n12782), .A2(n7590), .A3(n12781), .ZN(n7589) );
  OAI21_X2 U9766 ( .B1(n7597), .B2(n7596), .A(n7594), .ZN(n12475) );
  NAND2_X1 U9767 ( .A1(n7599), .A2(n7602), .ZN(n14648) );
  INV_X1 U9768 ( .A(n14377), .ZN(n7611) );
  AND2_X1 U9769 ( .A1(n11322), .A2(n11321), .ZN(n12839) );
  NAND2_X1 U9770 ( .A1(n7611), .A2(n12532), .ZN(n11322) );
  NAND2_X1 U9771 ( .A1(n12296), .A2(n7614), .ZN(n12442) );
  INV_X1 U9772 ( .A(n10481), .ZN(n7622) );
  OR2_X2 U9773 ( .A1(n10481), .A2(n12951), .ZN(n12753) );
  NAND3_X1 U9774 ( .A1(n10519), .A2(n10520), .A3(n7623), .ZN(n11355) );
  INV_X1 U9775 ( .A(n12931), .ZN(n7626) );
  NAND2_X1 U9776 ( .A1(n9032), .A2(n15591), .ZN(n9038) );
  AND2_X1 U9777 ( .A1(n13195), .A2(n13194), .ZN(n13196) );
  BUF_X4 U9778 ( .A(n10978), .Z(n12820) );
  NAND2_X1 U9779 ( .A1(n13116), .A2(n14618), .ZN(n14730) );
  XNOR2_X1 U9780 ( .A(n13113), .B(n12939), .ZN(n12913) );
  NAND2_X1 U9781 ( .A1(n8578), .A2(n8866), .ZN(n8579) );
  AND2_X4 U9782 ( .A1(n13133), .A2(n8384), .ZN(n8600) );
  INV_X1 U9783 ( .A(n13133), .ZN(n8383) );
  INV_X1 U9784 ( .A(n10820), .ZN(n10821) );
  NAND2_X1 U9785 ( .A1(n10032), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10034) );
  AOI22_X1 U9786 ( .A1(n10725), .A2(n9767), .B1(n13891), .B2(n9764), .ZN(n9768) );
  INV_X1 U9787 ( .A(n7766), .ZN(n7768) );
  OR2_X4 U9788 ( .A1(n12324), .A2(n10041), .ZN(n10523) );
  INV_X1 U9789 ( .A(n9713), .ZN(n11062) );
  NAND2_X1 U9790 ( .A1(n12539), .A2(n11356), .ZN(n12542) );
  AND2_X1 U9791 ( .A1(n13890), .A2(n10734), .ZN(n10735) );
  OAI21_X2 U9792 ( .B1(n9096), .B2(P2_IR_REG_0__SCAN_IN), .A(n9095), .ZN(
        n11474) );
  NAND2_X1 U9793 ( .A1(n9096), .A2(n14202), .ZN(n9095) );
  NAND2_X1 U9794 ( .A1(n9096), .A2(n9213), .ZN(n9105) );
  OAI211_X1 U9795 ( .C1(n13216), .C2(n9044), .A(n9043), .B(n13552), .ZN(n9047)
         );
  NAND2_X1 U9796 ( .A1(n9097), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n9100) );
  OAI22_X2 U9797 ( .A1(n9773), .A2(n9772), .B1(n9771), .B2(n9770), .ZN(n9774)
         );
  NOR2_X1 U9798 ( .A1(n9769), .A2(n9768), .ZN(n9773) );
  INV_X1 U9799 ( .A(n11641), .ZN(n9759) );
  NAND2_X1 U9800 ( .A1(n6868), .A2(n11632), .ZN(n12528) );
  OR2_X1 U9801 ( .A1(n9659), .A2(n9658), .ZN(n9661) );
  NAND2_X1 U9802 ( .A1(n9675), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9663) );
  NAND2_X4 U9803 ( .A1(n13121), .A2(n9072), .ZN(n9928) );
  NAND2_X1 U9804 ( .A1(n10724), .A2(n10723), .ZN(n10726) );
  NAND2_X1 U9805 ( .A1(n13829), .A2(n13828), .ZN(n13827) );
  INV_X1 U9806 ( .A(n13121), .ZN(n9070) );
  OR2_X1 U9807 ( .A1(n14109), .A2(n14099), .ZN(n7629) );
  XNOR2_X1 U9808 ( .A(n14508), .B(n14357), .ZN(n14504) );
  OR2_X1 U9809 ( .A1(n13410), .A2(n13623), .ZN(n7630) );
  AND2_X2 U9810 ( .A1(n11008), .A2(n9020), .ZN(n15607) );
  OR2_X1 U9811 ( .A1(n9830), .A2(n9829), .ZN(n7631) );
  OR2_X1 U9812 ( .A1(n14662), .A2(n12688), .ZN(n7632) );
  AND2_X1 U9813 ( .A1(n9850), .A2(n9847), .ZN(n7633) );
  AND2_X1 U9814 ( .A1(n13303), .A2(n13531), .ZN(n7634) );
  INV_X1 U9815 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n11981) );
  INV_X1 U9816 ( .A(n13262), .ZN(n13198) );
  INV_X1 U9817 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n7868) );
  INV_X1 U9818 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7715) );
  AND2_X2 U9819 ( .A1(n13103), .A2(n14706), .ZN(n15143) );
  XNOR2_X1 U9820 ( .A(n7848), .B(n7847), .ZN(n7637) );
  INV_X1 U9821 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n8357) );
  AND3_X1 U9822 ( .A1(n12622), .A2(n12621), .A3(n12620), .ZN(n7638) );
  AND2_X1 U9823 ( .A1(n12835), .A2(n12834), .ZN(n7639) );
  AND3_X1 U9824 ( .A1(n9996), .A2(n9995), .A3(n9994), .ZN(n7640) );
  INV_X1 U9825 ( .A(n14015), .ZN(n9751) );
  AND2_X1 U9826 ( .A1(n9712), .A2(n14086), .ZN(n14078) );
  INV_X1 U9827 ( .A(n14078), .ZN(n14088) );
  INV_X1 U9828 ( .A(n9765), .ZN(n9766) );
  AOI22_X1 U9829 ( .A1(n10725), .A2(n9826), .B1(n13891), .B2(n9767), .ZN(n9772) );
  OAI22_X1 U9830 ( .A1(n15306), .A2(n9870), .B1(n9722), .B2(n10005), .ZN(n9775) );
  OAI22_X1 U9831 ( .A1(n15306), .A2(n10005), .B1(n9722), .B2(n9870), .ZN(n9778) );
  OAI21_X1 U9832 ( .B1(n9782), .B2(n9781), .A(n9780), .ZN(n9784) );
  NAND2_X1 U9833 ( .A1(n9793), .A2(n9792), .ZN(n9795) );
  OAI22_X1 U9834 ( .A1(n11247), .A2(n9870), .B1(n11198), .B2(n10005), .ZN(
        n9809) );
  AOI22_X1 U9835 ( .A1(n9808), .A2(n9807), .B1(n9806), .B2(n9805), .ZN(n9810)
         );
  AOI21_X1 U9836 ( .B1(n9817), .B2(n9816), .A(n9815), .ZN(n9821) );
  INV_X1 U9837 ( .A(n9848), .ZN(n9845) );
  AND2_X1 U9838 ( .A1(n9863), .A2(n9862), .ZN(n9864) );
  NAND2_X1 U9839 ( .A1(n9894), .A2(n9893), .ZN(n9898) );
  INV_X1 U9840 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9058) );
  INV_X1 U9841 ( .A(n9553), .ZN(n9554) );
  INV_X1 U9842 ( .A(P3_REG1_REG_2__SCAN_IN), .ZN(n7767) );
  OR2_X1 U9843 ( .A1(n13306), .A2(n13238), .ZN(n8982) );
  INV_X1 U9844 ( .A(n8734), .ZN(n8376) );
  NAND2_X1 U9845 ( .A1(n13432), .A2(n8982), .ZN(n8983) );
  INV_X1 U9846 ( .A(n13556), .ZN(n8978) );
  INV_X1 U9847 ( .A(n9577), .ZN(n9575) );
  OR2_X1 U9848 ( .A1(n9597), .A2(n9596), .ZN(n9614) );
  INV_X1 U9849 ( .A(n9282), .ZN(n9280) );
  INV_X1 U9850 ( .A(n9709), .ZN(n9758) );
  INV_X1 U9851 ( .A(n12716), .ZN(n12507) );
  OR2_X1 U9852 ( .A1(n14508), .A2(n14357), .ZN(n12937) );
  INV_X1 U9853 ( .A(n12632), .ZN(n12505) );
  NAND2_X1 U9854 ( .A1(n12101), .A2(n12100), .ZN(n12171) );
  INV_X1 U9855 ( .A(n11434), .ZN(n12532) );
  OR2_X1 U9856 ( .A1(n8677), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8690) );
  NAND2_X1 U9857 ( .A1(n8376), .A2(n8126), .ZN(n8749) );
  NAND2_X1 U9858 ( .A1(n8374), .A2(n8230), .ZN(n8712) );
  INV_X1 U9859 ( .A(n12011), .ZN(n12008) );
  INV_X1 U9860 ( .A(n8586), .ZN(n8369) );
  NOR2_X1 U9861 ( .A1(n13219), .A2(n13520), .ZN(n9045) );
  OR2_X1 U9862 ( .A1(n13306), .A2(n13419), .ZN(n8916) );
  INV_X1 U9863 ( .A(n11765), .ZN(n8964) );
  INV_X1 U9864 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n9033) );
  AND2_X1 U9865 ( .A1(n8317), .A2(n8316), .ZN(n8506) );
  INV_X1 U9866 ( .A(n12159), .ZN(n12156) );
  XNOR2_X1 U9867 ( .A(n10725), .B(n10726), .ZN(n10730) );
  OR2_X1 U9868 ( .A1(n9460), .A2(n9459), .ZN(n9485) );
  INV_X1 U9869 ( .A(n13863), .ZN(n13769) );
  NAND2_X1 U9870 ( .A1(n9541), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n9565) );
  NAND2_X1 U9871 ( .A1(n9442), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9460) );
  NAND2_X1 U9872 ( .A1(n9280), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9299) );
  OR2_X1 U9873 ( .A1(n11062), .A2(n9711), .ZN(n10688) );
  INV_X1 U9874 ( .A(n9667), .ZN(n9757) );
  OAI21_X1 U9875 ( .B1(n9676), .B2(P2_IR_REG_22__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9702) );
  INV_X1 U9876 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n9127) );
  NOR2_X1 U9877 ( .A1(n12094), .A2(n14433), .ZN(n12175) );
  OR2_X1 U9878 ( .A1(n12415), .A2(n12414), .ZN(n12416) );
  OR2_X1 U9879 ( .A1(n12798), .A2(n14210), .ZN(n13105) );
  NAND2_X1 U9880 ( .A1(n12507), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n12729) );
  INV_X1 U9881 ( .A(n14504), .ZN(n12935) );
  NAND2_X1 U9882 ( .A1(n12307), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n12452) );
  OR2_X1 U9883 ( .A1(n8572), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8586) );
  NAND2_X1 U9884 ( .A1(n8372), .A2(n13207), .ZN(n8654) );
  OR2_X1 U9885 ( .A1(n8749), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8751) );
  NAND2_X1 U9886 ( .A1(n8375), .A2(n8086), .ZN(n8722) );
  NAND2_X1 U9887 ( .A1(n8371), .A2(n8370), .ZN(n8625) );
  NAND2_X1 U9888 ( .A1(n8500), .A2(n12012), .ZN(n8513) );
  OR2_X1 U9889 ( .A1(n8625), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8640) );
  NAND2_X1 U9890 ( .A1(n8369), .A2(n8368), .ZN(n8601) );
  AND2_X1 U9891 ( .A1(n8770), .A2(n8399), .ZN(n13402) );
  INV_X1 U9892 ( .A(n13534), .ZN(n13505) );
  AND4_X1 U9893 ( .A1(n8630), .A2(n8629), .A3(n8628), .A4(n8627), .ZN(n13517)
         );
  AND2_X1 U9894 ( .A1(n8875), .A2(n8874), .ZN(n12370) );
  AND2_X1 U9895 ( .A1(n10562), .A2(n15561), .ZN(n10553) );
  INV_X1 U9896 ( .A(n15607), .ZN(n9022) );
  OR2_X1 U9897 ( .A1(n13402), .A2(n13401), .ZN(n13624) );
  INV_X1 U9898 ( .A(n11531), .ZN(n15575) );
  INV_X1 U9899 ( .A(n11550), .ZN(n15550) );
  AND2_X1 U9900 ( .A1(n7745), .A2(n7759), .ZN(n11083) );
  NAND2_X1 U9901 ( .A1(n8662), .A2(n8341), .ZN(n8674) );
  NAND2_X1 U9902 ( .A1(n8610), .A2(n8334), .ZN(n8620) );
  AND2_X1 U9903 ( .A1(n8303), .A2(n8302), .ZN(n8427) );
  OR2_X1 U9904 ( .A1(n9418), .A2(n9417), .ZN(n9443) );
  OR2_X1 U9905 ( .A1(n9339), .A2(n11964), .ZN(n9361) );
  AND2_X1 U9906 ( .A1(n10692), .A2(n10066), .ZN(n13851) );
  INV_X1 U9907 ( .A(n13864), .ZN(n9907) );
  NAND2_X1 U9908 ( .A1(n11647), .A2(n9307), .ZN(n11586) );
  INV_X1 U9909 ( .A(n15274), .ZN(n14091) );
  INV_X1 U9910 ( .A(n13851), .ZN(n13839) );
  INV_X1 U9911 ( .A(n14969), .ZN(n14979) );
  AND2_X1 U9912 ( .A1(n9666), .A2(n9665), .ZN(n13962) );
  INV_X1 U9913 ( .A(n10686), .ZN(n10941) );
  OR2_X1 U9914 ( .A1(n9256), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n9411) );
  AND2_X1 U9915 ( .A1(n14273), .A2(n13044), .ZN(n14216) );
  NAND2_X1 U9916 ( .A1(n12071), .A2(n12073), .ZN(n12074) );
  INV_X1 U9917 ( .A(n14366), .ZN(n15041) );
  AND3_X1 U9918 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n11331) );
  AND3_X1 U9919 ( .A1(n11345), .A2(n11514), .A3(n10513), .ZN(n10527) );
  AND2_X1 U9920 ( .A1(n13105), .A2(n12799), .ZN(n14511) );
  NAND2_X1 U9921 ( .A1(n12506), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n12716) );
  INV_X1 U9922 ( .A(n12753), .ZN(n12810) );
  INV_X1 U9923 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n14433) );
  INV_X1 U9924 ( .A(n14524), .ZN(n14546) );
  AND2_X1 U9925 ( .A1(n10498), .A2(n10497), .ZN(n11345) );
  INV_X1 U9926 ( .A(n14363), .ZN(n14681) );
  INV_X1 U9927 ( .A(n14771), .ZN(n14702) );
  INV_X1 U9928 ( .A(n7937), .ZN(n7940) );
  NOR2_X1 U9929 ( .A1(n8469), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8487) );
  OR2_X1 U9930 ( .A1(n8513), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8528) );
  NOR2_X1 U9931 ( .A1(n10559), .A2(n10551), .ZN(n15393) );
  INV_X1 U9932 ( .A(n15401), .ZN(n13319) );
  INV_X1 U9933 ( .A(n13218), .ZN(n13303) );
  AND2_X1 U9934 ( .A1(n8697), .A2(n8696), .ZN(n13483) );
  NAND2_X1 U9935 ( .A1(n9047), .A2(n9046), .ZN(n13407) );
  INV_X1 U9936 ( .A(n13518), .ZN(n13531) );
  NAND2_X1 U9937 ( .A1(n9027), .A2(n8985), .ZN(n13552) );
  INV_X1 U9938 ( .A(n13125), .ZN(n13564) );
  NAND2_X1 U9939 ( .A1(n9022), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n9023) );
  AND2_X1 U9940 ( .A1(n9010), .A2(n9009), .ZN(n11008) );
  INV_X1 U9941 ( .A(n15570), .ZN(n14957) );
  AND2_X1 U9942 ( .A1(n11083), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10562) );
  INV_X1 U9943 ( .A(n15582), .ZN(n15561) );
  INV_X1 U9944 ( .A(n14072), .ZN(n14156) );
  AND2_X1 U9945 ( .A1(n9550), .A2(n9549), .ZN(n13832) );
  AND3_X1 U9946 ( .A1(n9367), .A2(n9366), .A3(n9365), .ZN(n12144) );
  INV_X1 U9947 ( .A(n13901), .ZN(n15255) );
  AND2_X1 U9948 ( .A1(n10068), .A2(n10071), .ZN(n15252) );
  INV_X1 U9949 ( .A(n9989), .ZN(n14000) );
  INV_X1 U9950 ( .A(n11680), .ZN(n11910) );
  INV_X1 U9951 ( .A(n13962), .ZN(n14065) );
  NAND2_X1 U9952 ( .A1(n15289), .A2(n10937), .ZN(n14086) );
  INV_X1 U9953 ( .A(n14094), .ZN(n15270) );
  AND2_X1 U9954 ( .A1(n15335), .A2(n15334), .ZN(n15000) );
  AND3_X1 U9955 ( .A1(n10941), .A2(n10940), .A3(n10939), .ZN(n10968) );
  OR3_X1 U9956 ( .A1(n11982), .A2(n11981), .A3(n11980), .ZN(n12094) );
  NAND2_X1 U9957 ( .A1(n10528), .A2(n14706), .ZN(n15067) );
  AND2_X1 U9958 ( .A1(n12735), .A2(n12734), .ZN(n14607) );
  NAND2_X1 U9959 ( .A1(n12702), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n10634) );
  INV_X1 U9960 ( .A(n15124), .ZN(n14477) );
  OR3_X1 U9961 ( .A1(n11730), .A2(n15105), .A3(n11729), .ZN(n12019) );
  NAND2_X1 U9962 ( .A1(n12911), .A2(n12910), .ZN(n12912) );
  INV_X1 U9963 ( .A(n15146), .ZN(n14713) );
  INV_X1 U9964 ( .A(n14716), .ZN(n14649) );
  AND2_X1 U9965 ( .A1(n11347), .A2(n15161), .ZN(n14815) );
  INV_X1 U9966 ( .A(n14815), .ZN(n15175) );
  AND2_X1 U9967 ( .A1(n10523), .A2(n10228), .ZN(n12880) );
  XNOR2_X1 U9968 ( .A(n10535), .B(P1_IR_REG_14__SCAN_IN), .ZN(n14451) );
  AND2_X1 U9969 ( .A1(n7853), .A2(n7852), .ZN(n15523) );
  NAND2_X1 U9970 ( .A1(n11085), .A2(P3_STATE_REG_SCAN_IN), .ZN(n15401) );
  AND2_X1 U9971 ( .A1(n8770), .A2(n8389), .ZN(n11375) );
  INV_X1 U9972 ( .A(n13519), .ZN(n13493) );
  INV_X1 U9973 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n15453) );
  OR2_X1 U9974 ( .A1(n7850), .A2(n7844), .ZN(n15516) );
  OR2_X1 U9975 ( .A1(n11010), .A2(n11663), .ZN(n13562) );
  INV_X1 U9976 ( .A(n13541), .ZN(n13560) );
  AND2_X1 U9977 ( .A1(n11010), .A2(n13538), .ZN(n13566) );
  OR2_X1 U9978 ( .A1(n13560), .A2(n11661), .ZN(n13125) );
  INV_X1 U9979 ( .A(n13153), .ZN(n13665) );
  INV_X1 U9980 ( .A(n15591), .ZN(n15589) );
  NAND2_X1 U9981 ( .A1(n15591), .A2(n15561), .ZN(n13674) );
  NAND2_X1 U9982 ( .A1(n10242), .A2(n10241), .ZN(n10243) );
  INV_X1 U9983 ( .A(SI_17_), .ZN(n10532) );
  INV_X1 U9984 ( .A(SI_12_), .ZN(n10180) );
  INV_X1 U9985 ( .A(n13681), .ZN(n13688) );
  OR2_X1 U9986 ( .A1(n10696), .A2(n10683), .ZN(n13855) );
  INV_X1 U9987 ( .A(n13853), .ZN(n13845) );
  NAND2_X1 U9988 ( .A1(n9640), .A2(n9639), .ZN(n13863) );
  INV_X1 U9989 ( .A(n13842), .ZN(n13872) );
  INV_X1 U9990 ( .A(n12358), .ZN(n13876) );
  OR2_X1 U9991 ( .A1(n10072), .A2(n10071), .ZN(n13901) );
  INV_X1 U9992 ( .A(n15252), .ZN(n12354) );
  OR2_X1 U9993 ( .A1(n10110), .A2(P2_U3088), .ZN(n15228) );
  NAND2_X1 U9994 ( .A1(n10968), .A2(n10967), .ZN(n15355) );
  OR3_X1 U9995 ( .A1(n14170), .A2(n14169), .A3(n14168), .ZN(n14185) );
  INV_X1 U9996 ( .A(n15347), .ZN(n15346) );
  OR2_X1 U9997 ( .A1(n15285), .A2(n15283), .ZN(n15284) );
  INV_X1 U9998 ( .A(n15289), .ZN(n15285) );
  INV_X1 U9999 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n10200) );
  AND2_X1 U10000 ( .A1(n10246), .A2(n10244), .ZN(n14435) );
  NAND2_X1 U10001 ( .A1(n10987), .A2(P1_STATE_REG_SCAN_IN), .ZN(n15072) );
  INV_X1 U10002 ( .A(n14794), .ZN(n14668) );
  NAND2_X1 U10003 ( .A1(n12818), .A2(n12817), .ZN(n14356) );
  INV_X1 U10004 ( .A(n14607), .ZN(n14772) );
  OR2_X1 U10005 ( .A1(n10318), .A2(n13102), .ZN(n15124) );
  INV_X1 U10006 ( .A(n14480), .ZN(n15122) );
  OR2_X1 U10007 ( .A1(n15143), .A2(n11369), .ZN(n14709) );
  OR2_X1 U10008 ( .A1(n15143), .A2(n11605), .ZN(n14716) );
  NAND2_X1 U10009 ( .A1(n15184), .A2(n15157), .ZN(n14804) );
  INV_X2 U10010 ( .A(n15181), .ZN(n15184) );
  INV_X1 U10011 ( .A(n14488), .ZN(n14820) );
  INV_X1 U10012 ( .A(n13039), .ZN(n14839) );
  NAND2_X1 U10013 ( .A1(n14854), .A2(n15157), .ZN(n14858) );
  INV_X1 U10014 ( .A(n14854), .ZN(n15177) );
  AND2_X1 U10015 ( .A1(n10522), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10228) );
  INV_X1 U10016 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n10287) );
  INV_X1 U10017 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n10179) );
  XNOR2_X1 U10018 ( .A(n8294), .B(n8293), .ZN(n8295) );
  INV_X1 U10019 ( .A(n13329), .ZN(P3_U3897) );
  AND2_X1 U10020 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10065), .ZN(P2_U3947) );
  NAND2_X1 U10021 ( .A1(n9761), .A2(n7629), .ZN(P2_U3236) );
  NOR2_X2 U10022 ( .A1(P3_IR_REG_9__SCAN_IN), .A2(P3_IR_REG_8__SCAN_IN), .ZN(
        n7646) );
  NOR2_X1 U10023 ( .A1(P3_IR_REG_3__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n7643) );
  NOR2_X1 U10024 ( .A1(P3_IR_REG_6__SCAN_IN), .A2(P3_IR_REG_11__SCAN_IN), .ZN(
        n7642) );
  NOR2_X1 U10025 ( .A1(P3_IR_REG_16__SCAN_IN), .A2(P3_IR_REG_17__SCAN_IN), 
        .ZN(n7650) );
  NOR2_X1 U10026 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), 
        .ZN(n7649) );
  INV_X1 U10027 ( .A(n7749), .ZN(n7757) );
  OAI21_X1 U10028 ( .B1(n7657), .B2(P3_IR_REG_24__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7652) );
  MUX2_X1 U10029 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7652), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n7656) );
  NOR2_X1 U10030 ( .A1(P3_IR_REG_24__SCAN_IN), .A2(P3_IR_REG_25__SCAN_IN), 
        .ZN(n7654) );
  INV_X1 U10031 ( .A(n7747), .ZN(n7655) );
  NAND2_X1 U10032 ( .A1(n7749), .A2(n7655), .ZN(n7660) );
  NAND2_X1 U10033 ( .A1(n7656), .A2(n7660), .ZN(n12033) );
  INV_X1 U10034 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7658) );
  XNOR2_X2 U10035 ( .A(n7659), .B(n7658), .ZN(n12892) );
  INV_X1 U10036 ( .A(n12892), .ZN(n7662) );
  NAND2_X1 U10037 ( .A1(n7660), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7661) );
  NAND2_X1 U10038 ( .A1(n7662), .A2(n8993), .ZN(n7663) );
  NAND2_X1 U10039 ( .A1(n6783), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7665) );
  XNOR2_X1 U10040 ( .A(n7665), .B(n7664), .ZN(n7759) );
  NAND2_X1 U10041 ( .A1(n7759), .A2(P3_STATE_REG_SCAN_IN), .ZN(n10218) );
  INV_X1 U10042 ( .A(P3_IR_REG_15__SCAN_IN), .ZN(n7668) );
  INV_X1 U10043 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7669) );
  NAND2_X1 U10044 ( .A1(n7674), .A2(n7669), .ZN(n7739) );
  OAI21_X2 U10045 ( .B1(n7672), .B2(P3_IR_REG_18__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7671) );
  INV_X1 U10046 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7670) );
  XNOR2_X1 U10047 ( .A(n7457), .B(P3_REG2_REG_19__SCAN_IN), .ZN(n7845) );
  NAND2_X1 U10048 ( .A1(n7672), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7673) );
  XNOR2_X1 U10049 ( .A(n7673), .B(P3_IR_REG_18__SCAN_IN), .ZN(n14917) );
  INV_X1 U10050 ( .A(n14917), .ZN(n10540) );
  INV_X1 U10051 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n7741) );
  OR2_X1 U10052 ( .A1(n7674), .A2(n7715), .ZN(n7675) );
  XNOR2_X1 U10053 ( .A(n7675), .B(P3_IR_REG_16__SCAN_IN), .ZN(n8597) );
  INV_X1 U10054 ( .A(n8597), .ZN(n13374) );
  OR2_X1 U10055 ( .A1(n7676), .A2(n7715), .ZN(n7677) );
  XNOR2_X1 U10056 ( .A(n7677), .B(P3_IR_REG_15__SCAN_IN), .ZN(n13361) );
  OR2_X1 U10057 ( .A1(n7667), .A2(n7715), .ZN(n7679) );
  XNOR2_X1 U10058 ( .A(n7679), .B(n7678), .ZN(n15519) );
  NAND2_X1 U10059 ( .A1(n7680), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7681) );
  MUX2_X1 U10060 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7681), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n7683) );
  INV_X1 U10061 ( .A(n7667), .ZN(n7682) );
  NAND2_X1 U10062 ( .A1(n7683), .A2(n7682), .ZN(n10253) );
  NAND2_X1 U10063 ( .A1(n7684), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7685) );
  MUX2_X1 U10064 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7685), .S(
        P3_IR_REG_12__SCAN_IN), .Z(n7686) );
  NAND2_X1 U10065 ( .A1(n7686), .A2(n7680), .ZN(n15500) );
  INV_X1 U10066 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7688) );
  INV_X1 U10067 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7696) );
  NAND2_X1 U10068 ( .A1(n7695), .A2(n7696), .ZN(n7693) );
  OAI21_X1 U10069 ( .B1(n7690), .B2(P3_IR_REG_10__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7689) );
  XNOR2_X1 U10070 ( .A(n7689), .B(P3_IR_REG_11__SCAN_IN), .ZN(n11906) );
  NAND2_X1 U10071 ( .A1(n7690), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7692) );
  INV_X1 U10072 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7691) );
  NAND2_X1 U10073 ( .A1(n7693), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7694) );
  XNOR2_X1 U10074 ( .A(n7694), .B(P3_IR_REG_9__SCAN_IN), .ZN(n10153) );
  OR2_X1 U10075 ( .A1(n7698), .A2(n7715), .ZN(n7699) );
  OR2_X1 U10076 ( .A1(n7700), .A2(n7715), .ZN(n7702) );
  NAND2_X1 U10077 ( .A1(n7703), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7704) );
  NAND2_X1 U10078 ( .A1(n7705), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7707) );
  INV_X1 U10079 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n11014) );
  NOR2_X1 U10080 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(n11014), .ZN(n10954) );
  NAND2_X1 U10081 ( .A1(n7709), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7708) );
  INV_X1 U10082 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n11665) );
  INV_X1 U10083 ( .A(n7709), .ZN(n7710) );
  OAI21_X1 U10084 ( .B1(P3_REG2_REG_2__SCAN_IN), .B2(n7766), .A(n7713), .ZN(
        n10569) );
  XNOR2_X1 U10085 ( .A(n7717), .B(n7716), .ZN(n8429) );
  XNOR2_X1 U10086 ( .A(n7718), .B(n8429), .ZN(n10584) );
  INV_X1 U10087 ( .A(n7718), .ZN(n7719) );
  NAND2_X1 U10088 ( .A1(n7719), .A2(n8429), .ZN(n7720) );
  NAND2_X1 U10089 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n15417), .ZN(n7721) );
  OAI21_X1 U10090 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n15417), .A(n7721), .ZN(
        n15405) );
  NOR2_X1 U10091 ( .A1(n15434), .A2(n7722), .ZN(n7723) );
  INV_X1 U10092 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n15424) );
  XNOR2_X1 U10093 ( .A(n7722), .B(n15434), .ZN(n15423) );
  NAND2_X1 U10094 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n15442), .ZN(n7724) );
  OAI21_X1 U10095 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n15442), .A(n7724), .ZN(
        n15445) );
  NOR2_X1 U10096 ( .A1(n15464), .A2(n7725), .ZN(n7726) );
  INV_X1 U10097 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n15456) );
  NAND2_X1 U10098 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n15483), .ZN(n7727) );
  OAI21_X1 U10099 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n15483), .A(n7727), .ZN(
        n15474) );
  NOR2_X1 U10100 ( .A1(n10153), .A2(n7728), .ZN(n7729) );
  INV_X1 U10101 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n11533) );
  NAND2_X1 U10102 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n10163), .ZN(n7730) );
  OAI21_X1 U10103 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n10163), .A(n7730), .ZN(
        n11155) );
  NOR2_X1 U10104 ( .A1(n11906), .A2(n7731), .ZN(n7732) );
  INV_X1 U10105 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n12056) );
  NAND2_X1 U10106 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n15500), .ZN(n7733) );
  OAI21_X1 U10107 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n15500), .A(n7733), .ZN(
        n15495) );
  NOR2_X1 U10108 ( .A1(n6870), .A2(n7734), .ZN(n7735) );
  INV_X1 U10109 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n13333) );
  XNOR2_X1 U10110 ( .A(n15519), .B(P3_REG2_REG_14__SCAN_IN), .ZN(n15511) );
  NOR2_X1 U10111 ( .A1(n13361), .A2(n7736), .ZN(n7737) );
  INV_X1 U10112 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n13351) );
  XNOR2_X1 U10113 ( .A(n7736), .B(n13361), .ZN(n13350) );
  INV_X1 U10114 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n7738) );
  AOI22_X1 U10115 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n8597), .B1(n13374), 
        .B2(n7738), .ZN(n13366) );
  NAND2_X1 U10116 ( .A1(n7739), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7740) );
  XNOR2_X1 U10117 ( .A(n7740), .B(P3_IR_REG_17__SCAN_IN), .ZN(n13397) );
  NOR2_X1 U10118 ( .A1(n13397), .A2(n7742), .ZN(n7743) );
  NAND2_X1 U10119 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n10540), .ZN(n7744) );
  OAI21_X1 U10120 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n10540), .A(n7744), .ZN(
        n14922) );
  INV_X1 U10121 ( .A(n10562), .ZN(n7746) );
  OR2_X1 U10122 ( .A1(n7759), .A2(P3_U3151), .ZN(n11445) );
  NAND2_X1 U10123 ( .A1(n7746), .A2(n11445), .ZN(n7853) );
  AND2_X2 U10124 ( .A1(n7750), .A2(n6890), .ZN(n8378) );
  INV_X1 U10125 ( .A(n8378), .ZN(n8380) );
  INV_X1 U10126 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7752) );
  INV_X1 U10127 ( .A(n7754), .ZN(n7755) );
  NAND2_X1 U10128 ( .A1(n7755), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7756) );
  NAND2_X1 U10129 ( .A1(n7757), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7758) );
  AND2_X2 U10130 ( .A1(n11190), .A2(n10704), .ZN(n9015) );
  NAND2_X1 U10131 ( .A1(n9015), .A2(n7759), .ZN(n7760) );
  AND2_X1 U10132 ( .A1(n6879), .A2(n7760), .ZN(n7851) );
  NAND2_X1 U10133 ( .A1(n7853), .A2(n7851), .ZN(n7850) );
  INV_X1 U10134 ( .A(n6812), .ZN(n7849) );
  NAND2_X1 U10135 ( .A1(n7849), .A2(n7844), .ZN(n8986) );
  INV_X1 U10136 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n10545) );
  NOR2_X1 U10137 ( .A1(n10545), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n7762) );
  INV_X1 U10138 ( .A(n7762), .ZN(n10955) );
  NOR2_X1 U10139 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n10955), .ZN(n7765) );
  NAND2_X1 U10140 ( .A1(n10160), .A2(n10955), .ZN(n7764) );
  NAND2_X1 U10141 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n7762), .ZN(n7763) );
  NAND2_X1 U10142 ( .A1(n7764), .A2(n7763), .ZN(n10602) );
  NOR2_X1 U10143 ( .A1(n7765), .A2(n10605), .ZN(n10574) );
  NAND2_X1 U10144 ( .A1(P3_REG1_REG_2__SCAN_IN), .A2(n7766), .ZN(n7769) );
  INV_X1 U10145 ( .A(n7769), .ZN(n7770) );
  INV_X1 U10146 ( .A(n8429), .ZN(n10594) );
  NAND2_X1 U10147 ( .A1(P3_REG1_REG_4__SCAN_IN), .A2(n15417), .ZN(n7773) );
  OAI21_X1 U10148 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n15417), .A(n7773), .ZN(
        n15408) );
  NOR2_X1 U10149 ( .A1(n15434), .A2(n7774), .ZN(n7775) );
  INV_X1 U10150 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n15596) );
  XNOR2_X1 U10151 ( .A(n7774), .B(n15434), .ZN(n15426) );
  NAND2_X1 U10152 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n15442), .ZN(n7776) );
  OAI21_X1 U10153 ( .B1(P3_REG1_REG_6__SCAN_IN), .B2(n15442), .A(n7776), .ZN(
        n15440) );
  NOR2_X1 U10154 ( .A1(n15441), .A2(n15440), .ZN(n15439) );
  NOR2_X1 U10155 ( .A1(n15464), .A2(n7777), .ZN(n7778) );
  INV_X1 U10156 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15600) );
  NAND2_X1 U10157 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n15483), .ZN(n7779) );
  OAI21_X1 U10158 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n15483), .A(n7779), .ZN(
        n15481) );
  NOR2_X1 U10159 ( .A1(n10153), .A2(n7780), .ZN(n7781) );
  INV_X1 U10160 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15604) );
  NAND2_X1 U10161 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n10163), .ZN(n7782) );
  OAI21_X1 U10162 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n10163), .A(n7782), .ZN(
        n11153) );
  NOR2_X1 U10163 ( .A1(n11906), .A2(n7783), .ZN(n7784) );
  INV_X1 U10164 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14958) );
  NAND2_X1 U10165 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n15500), .ZN(n7785) );
  OAI21_X1 U10166 ( .B1(P3_REG1_REG_12__SCAN_IN), .B2(n15500), .A(n7785), .ZN(
        n15497) );
  INV_X1 U10167 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14947) );
  XNOR2_X1 U10168 ( .A(n15519), .B(P3_REG1_REG_14__SCAN_IN), .ZN(n15514) );
  INV_X1 U10169 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n14937) );
  INV_X1 U10170 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n13621) );
  AOI22_X1 U10171 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n8597), .B1(n13374), 
        .B2(n13621), .ZN(n13376) );
  XNOR2_X1 U10172 ( .A(n7788), .B(n13397), .ZN(n13384) );
  INV_X1 U10173 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n13617) );
  NOR2_X1 U10174 ( .A1(n13397), .A2(n7788), .ZN(n7789) );
  INV_X1 U10175 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n7840) );
  AOI22_X1 U10176 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n14917), .B1(n10540), 
        .B2(n7840), .ZN(n14919) );
  INV_X1 U10177 ( .A(P3_REG1_REG_19__SCAN_IN), .ZN(n13607) );
  XNOR2_X1 U10178 ( .A(n7457), .B(n13607), .ZN(n7843) );
  INV_X4 U10179 ( .A(n7844), .ZN(n12217) );
  MUX2_X1 U10180 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12217), .Z(n7838) );
  INV_X1 U10181 ( .A(n13397), .ZN(n10531) );
  AND2_X1 U10182 ( .A1(n7838), .A2(n10531), .ZN(n7839) );
  MUX2_X1 U10183 ( .A(n7738), .B(n13621), .S(n12217), .Z(n7835) );
  NOR2_X1 U10184 ( .A1(n7835), .A2(n8597), .ZN(n13368) );
  MUX2_X1 U10185 ( .A(P3_REG2_REG_14__SCAN_IN), .B(P3_REG1_REG_14__SCAN_IN), 
        .S(n12217), .Z(n7831) );
  MUX2_X1 U10186 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12217), .Z(n7830) );
  XNOR2_X1 U10187 ( .A(n7830), .B(n10253), .ZN(n13336) );
  MUX2_X1 U10188 ( .A(P3_REG2_REG_12__SCAN_IN), .B(P3_REG1_REG_12__SCAN_IN), 
        .S(n12217), .Z(n7827) );
  NAND2_X1 U10189 ( .A1(n7827), .A2(n15500), .ZN(n7828) );
  MUX2_X1 U10190 ( .A(P3_REG2_REG_11__SCAN_IN), .B(P3_REG1_REG_11__SCAN_IN), 
        .S(n12217), .Z(n7825) );
  INV_X1 U10191 ( .A(n7825), .ZN(n7826) );
  INV_X1 U10192 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n7791) );
  INV_X1 U10193 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n7790) );
  MUX2_X1 U10194 ( .A(n7791), .B(n7790), .S(n12217), .Z(n7823) );
  INV_X1 U10195 ( .A(n10163), .ZN(n11164) );
  AND2_X1 U10196 ( .A1(n7823), .A2(n11164), .ZN(n7824) );
  MUX2_X1 U10197 ( .A(n11533), .B(n15604), .S(n12217), .Z(n7821) );
  OR2_X1 U10198 ( .A1(n7821), .A2(n10153), .ZN(n11048) );
  MUX2_X1 U10199 ( .A(P3_REG2_REG_1__SCAN_IN), .B(P3_REG1_REG_1__SCAN_IN), .S(
        n7761), .Z(n7792) );
  INV_X1 U10200 ( .A(n10160), .ZN(n10613) );
  XNOR2_X1 U10201 ( .A(n7792), .B(n10613), .ZN(n10606) );
  MUX2_X1 U10202 ( .A(n11014), .B(n10545), .S(n7761), .Z(n10963) );
  NAND2_X1 U10203 ( .A1(n10606), .A2(n10962), .ZN(n7795) );
  INV_X1 U10204 ( .A(n7792), .ZN(n7793) );
  NAND2_X1 U10205 ( .A1(n7793), .A2(n10613), .ZN(n7794) );
  NAND2_X1 U10206 ( .A1(n7795), .A2(n7794), .ZN(n10566) );
  MUX2_X1 U10207 ( .A(P3_REG2_REG_2__SCAN_IN), .B(P3_REG1_REG_2__SCAN_IN), .S(
        n12217), .Z(n7796) );
  XNOR2_X1 U10208 ( .A(n7796), .B(n7768), .ZN(n10567) );
  NAND2_X1 U10209 ( .A1(n10566), .A2(n10567), .ZN(n7799) );
  INV_X1 U10210 ( .A(n7796), .ZN(n7797) );
  NAND2_X1 U10211 ( .A1(n7797), .A2(n7768), .ZN(n7798) );
  NAND2_X1 U10212 ( .A1(n7799), .A2(n7798), .ZN(n10581) );
  MUX2_X1 U10213 ( .A(P3_REG2_REG_3__SCAN_IN), .B(P3_REG1_REG_3__SCAN_IN), .S(
        n12217), .Z(n7800) );
  XNOR2_X1 U10214 ( .A(n7800), .B(n10594), .ZN(n10582) );
  NAND2_X1 U10215 ( .A1(n10581), .A2(n10582), .ZN(n7803) );
  INV_X1 U10216 ( .A(n7800), .ZN(n7801) );
  NAND2_X1 U10217 ( .A1(n7801), .A2(n10594), .ZN(n7802) );
  NAND2_X1 U10218 ( .A1(n7803), .A2(n7802), .ZN(n15413) );
  MUX2_X1 U10219 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12217), .Z(n7804) );
  INV_X1 U10220 ( .A(n15417), .ZN(n10129) );
  XNOR2_X1 U10221 ( .A(n7804), .B(n10129), .ZN(n15412) );
  NAND2_X1 U10222 ( .A1(n15413), .A2(n15412), .ZN(n7807) );
  INV_X1 U10223 ( .A(n7804), .ZN(n7805) );
  NAND2_X1 U10224 ( .A1(n7805), .A2(n10129), .ZN(n7806) );
  NAND2_X1 U10225 ( .A1(n7807), .A2(n7806), .ZN(n15429) );
  MUX2_X1 U10226 ( .A(P3_REG2_REG_5__SCAN_IN), .B(P3_REG1_REG_5__SCAN_IN), .S(
        n12217), .Z(n7808) );
  XNOR2_X1 U10227 ( .A(n7808), .B(n15434), .ZN(n15430) );
  NAND2_X1 U10228 ( .A1(n15429), .A2(n15430), .ZN(n7811) );
  INV_X1 U10229 ( .A(n7808), .ZN(n7809) );
  NAND2_X1 U10230 ( .A1(n7809), .A2(n15434), .ZN(n7810) );
  NAND2_X1 U10231 ( .A1(n7811), .A2(n7810), .ZN(n15438) );
  MUX2_X1 U10232 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12217), .Z(n7812) );
  INV_X1 U10233 ( .A(n15442), .ZN(n7813) );
  XNOR2_X1 U10234 ( .A(n7812), .B(n7813), .ZN(n15437) );
  NAND2_X1 U10235 ( .A1(n15438), .A2(n15437), .ZN(n7816) );
  INV_X1 U10236 ( .A(n7812), .ZN(n7814) );
  NAND2_X1 U10237 ( .A1(n7814), .A2(n7813), .ZN(n7815) );
  NAND2_X1 U10238 ( .A1(n7816), .A2(n7815), .ZN(n15459) );
  MUX2_X1 U10239 ( .A(P3_REG2_REG_7__SCAN_IN), .B(P3_REG1_REG_7__SCAN_IN), .S(
        n12217), .Z(n7817) );
  XNOR2_X1 U10240 ( .A(n7817), .B(n15464), .ZN(n15458) );
  INV_X1 U10241 ( .A(n7817), .ZN(n7818) );
  AND2_X1 U10242 ( .A1(n7818), .A2(n15464), .ZN(n7819) );
  MUX2_X1 U10243 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12217), .Z(n7820) );
  XNOR2_X1 U10244 ( .A(n7820), .B(n15483), .ZN(n15477) );
  OAI22_X1 U10245 ( .A1(n15478), .A2(n15477), .B1(n7820), .B2(n15483), .ZN(
        n11050) );
  AND2_X1 U10246 ( .A1(n7821), .A2(n10153), .ZN(n11046) );
  AOI21_X1 U10247 ( .B1(n11048), .B2(n11050), .A(n11046), .ZN(n11159) );
  INV_X1 U10248 ( .A(n7824), .ZN(n7822) );
  OAI21_X1 U10249 ( .B1(n11164), .B2(n7823), .A(n7822), .ZN(n11160) );
  NOR2_X1 U10250 ( .A1(n7824), .A2(n11158), .ZN(n11897) );
  INV_X1 U10251 ( .A(n11906), .ZN(n10168) );
  XNOR2_X1 U10252 ( .A(n7825), .B(n10168), .ZN(n11898) );
  INV_X1 U10253 ( .A(n15500), .ZN(n8550) );
  XNOR2_X1 U10254 ( .A(n7827), .B(n8550), .ZN(n15505) );
  NAND2_X1 U10255 ( .A1(n15506), .A2(n15505), .ZN(n15503) );
  NAND2_X1 U10256 ( .A1(n7828), .A2(n15503), .ZN(n13335) );
  INV_X1 U10257 ( .A(n13334), .ZN(n7829) );
  OAI21_X1 U10258 ( .B1(n7830), .B2(n10253), .A(n7829), .ZN(n15525) );
  MUX2_X1 U10259 ( .A(n15511), .B(n15514), .S(n12217), .Z(n15526) );
  AOI21_X1 U10260 ( .B1(n15519), .B2(n7831), .A(n15524), .ZN(n7833) );
  AND2_X1 U10261 ( .A1(n7833), .A2(n13361), .ZN(n7834) );
  INV_X1 U10262 ( .A(n7834), .ZN(n7832) );
  OAI21_X1 U10263 ( .B1(n13361), .B2(n7833), .A(n7832), .ZN(n13356) );
  MUX2_X1 U10264 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12217), .Z(n13357) );
  NOR2_X1 U10265 ( .A1(n7834), .A2(n13355), .ZN(n13370) );
  AND2_X1 U10266 ( .A1(n7835), .A2(n8597), .ZN(n13369) );
  INV_X1 U10267 ( .A(n13369), .ZN(n7836) );
  OAI21_X1 U10268 ( .B1(n13368), .B2(n13370), .A(n7836), .ZN(n13393) );
  INV_X1 U10269 ( .A(n7839), .ZN(n7837) );
  OAI21_X1 U10270 ( .B1(n7838), .B2(n10531), .A(n7837), .ZN(n13394) );
  NOR2_X1 U10271 ( .A1(n13393), .A2(n13394), .ZN(n13392) );
  INV_X1 U10272 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n13540) );
  MUX2_X1 U10273 ( .A(n13540), .B(n7840), .S(n12217), .Z(n14926) );
  NAND2_X1 U10274 ( .A1(n14927), .A2(n14926), .ZN(n14925) );
  NAND2_X1 U10275 ( .A1(n14917), .A2(n7841), .ZN(n7842) );
  NAND2_X1 U10276 ( .A1(n14925), .A2(n7842), .ZN(n7848) );
  INV_X1 U10277 ( .A(n7843), .ZN(n7846) );
  MUX2_X1 U10278 ( .A(n7846), .B(n7845), .S(n7844), .Z(n7847) );
  AND2_X1 U10279 ( .A1(P3_U3897), .A2(n6812), .ZN(n15504) );
  INV_X1 U10280 ( .A(n15504), .ZN(n7858) );
  MUX2_X1 U10281 ( .A(n7850), .B(n13329), .S(n7849), .Z(n15520) );
  NAND2_X1 U10282 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(P3_U3151), .ZN(n7855) );
  INV_X1 U10283 ( .A(n7851), .ZN(n7852) );
  NAND2_X1 U10284 ( .A1(n15523), .A2(P3_ADDR_REG_19__SCAN_IN), .ZN(n7854) );
  OAI211_X1 U10285 ( .C1(n15520), .C2(n10768), .A(n7855), .B(n7854), .ZN(n7856) );
  INV_X1 U10286 ( .A(n7856), .ZN(n7857) );
  INV_X1 U10287 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n15115) );
  XOR2_X1 U10288 ( .A(P3_ADDR_REG_15__SCAN_IN), .B(n15115), .Z(n7888) );
  INV_X1 U10289 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14449) );
  XOR2_X1 U10290 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n14449), .Z(n7890) );
  INV_X1 U10291 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7891) );
  INV_X1 U10292 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n7884) );
  XOR2_X1 U10293 ( .A(P1_ADDR_REG_12__SCAN_IN), .B(n7884), .Z(n7894) );
  INV_X1 U10294 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n7882) );
  INV_X1 U10295 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n7878) );
  XOR2_X1 U10296 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n7878), .Z(n7898) );
  INV_X1 U10297 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n15493) );
  XOR2_X1 U10298 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n15493), .Z(n7900) );
  XOR2_X1 U10299 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n15453), .Z(n7917) );
  XOR2_X1 U10300 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n7862), .Z(n7904) );
  NAND2_X1 U10301 ( .A1(n7907), .A2(n7906), .ZN(n7861) );
  NAND2_X1 U10302 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n7863), .ZN(n7865) );
  NAND2_X1 U10303 ( .A1(n7903), .A2(n14393), .ZN(n7864) );
  INV_X1 U10304 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n10669) );
  NAND2_X1 U10305 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n7866), .ZN(n7867) );
  NAND2_X1 U10306 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n7869), .ZN(n7871) );
  INV_X1 U10307 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10327) );
  NAND2_X1 U10308 ( .A1(n7913), .A2(n10327), .ZN(n7870) );
  NAND2_X1 U10309 ( .A1(n7917), .A2(n7918), .ZN(n7872) );
  NAND2_X1 U10310 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n7873), .ZN(n7875) );
  INV_X1 U10311 ( .A(P3_ADDR_REG_7__SCAN_IN), .ZN(n15472) );
  XNOR2_X1 U10312 ( .A(n15472), .B(n7873), .ZN(n7924) );
  INV_X1 U10313 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n7923) );
  NAND2_X1 U10314 ( .A1(n7924), .A2(n7923), .ZN(n7874) );
  NAND2_X1 U10315 ( .A1(n7875), .A2(n7874), .ZN(n7901) );
  NAND2_X1 U10316 ( .A1(n7900), .A2(n7901), .ZN(n7876) );
  NAND2_X1 U10317 ( .A1(n7898), .A2(n7899), .ZN(n7877) );
  INV_X1 U10318 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14415) );
  INV_X1 U10319 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10431) );
  XNOR2_X1 U10320 ( .A(n10431), .B(n7882), .ZN(n7896) );
  NAND2_X1 U10321 ( .A1(n7897), .A2(n7896), .ZN(n7881) );
  NAND2_X1 U10322 ( .A1(n7894), .A2(n7895), .ZN(n7883) );
  OR2_X1 U10323 ( .A1(n7891), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n7885) );
  AOI22_X1 U10324 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n7891), .B1(n7893), .B2(
        n7885), .ZN(n7889) );
  NAND2_X1 U10325 ( .A1(n7890), .A2(n7889), .ZN(n7886) );
  OAI21_X1 U10326 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14449), .A(n7886), .ZN(
        n7887) );
  INV_X1 U10327 ( .A(n7887), .ZN(n7939) );
  XOR2_X1 U10328 ( .A(n7888), .B(n7939), .Z(n15099) );
  XNOR2_X1 U10329 ( .A(n7890), .B(n7889), .ZN(n15095) );
  XNOR2_X1 U10330 ( .A(n7891), .B(P3_ADDR_REG_13__SCAN_IN), .ZN(n7892) );
  XNOR2_X1 U10331 ( .A(n7893), .B(n7892), .ZN(n15091) );
  XNOR2_X1 U10332 ( .A(n7895), .B(n7894), .ZN(n7934) );
  XOR2_X1 U10333 ( .A(n7897), .B(n7896), .Z(n15081) );
  XOR2_X1 U10334 ( .A(n7899), .B(n7898), .Z(n7928) );
  XOR2_X1 U10335 ( .A(n7901), .B(n7900), .Z(n14897) );
  XNOR2_X1 U10336 ( .A(n10669), .B(n6694), .ZN(n7902) );
  AND2_X1 U10337 ( .A1(n7902), .A2(P2_ADDR_REG_4__SCAN_IN), .ZN(n7912) );
  XOR2_X1 U10338 ( .A(n7903), .B(n14393), .Z(n15619) );
  XOR2_X1 U10339 ( .A(n7905), .B(n7904), .Z(n14890) );
  NOR2_X1 U10340 ( .A1(n7909), .A2(n7309), .ZN(n7910) );
  AOI21_X1 U10341 ( .B1(n10957), .B2(P1_ADDR_REG_0__SCAN_IN), .A(n7907), .ZN(
        n7908) );
  INV_X1 U10342 ( .A(n7908), .ZN(n15614) );
  NAND2_X1 U10343 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(n15614), .ZN(n15624) );
  NOR2_X1 U10344 ( .A1(n15624), .A2(n15623), .ZN(n15622) );
  NAND2_X1 U10345 ( .A1(n14890), .A2(n14889), .ZN(n14888) );
  NAND2_X1 U10346 ( .A1(n15619), .A2(n15620), .ZN(n15618) );
  OAI21_X1 U10347 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(n7911), .A(n15618), .ZN(
        n15609) );
  NAND2_X1 U10348 ( .A1(n7914), .A2(n7915), .ZN(n7916) );
  INV_X1 U10349 ( .A(P2_ADDR_REG_5__SCAN_IN), .ZN(n15612) );
  NOR2_X1 U10350 ( .A1(n7919), .A2(n7005), .ZN(n7920) );
  XOR2_X1 U10351 ( .A(n7918), .B(n7917), .Z(n14894) );
  INV_X1 U10352 ( .A(P2_ADDR_REG_7__SCAN_IN), .ZN(n7921) );
  NAND2_X1 U10353 ( .A1(n7922), .A2(n7921), .ZN(n7925) );
  XNOR2_X1 U10354 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n7922), .ZN(n15617) );
  XOR2_X1 U10355 ( .A(n7924), .B(n7923), .Z(n15616) );
  NAND2_X1 U10356 ( .A1(n15617), .A2(n15616), .ZN(n15615) );
  NAND2_X1 U10357 ( .A1(n14897), .A2(n14896), .ZN(n7926) );
  NOR2_X1 U10358 ( .A1(n14897), .A2(n14896), .ZN(n14895) );
  AOI21_X2 U10359 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(n7926), .A(n14895), .ZN(
        n7927) );
  XNOR2_X1 U10360 ( .A(n7928), .B(n7927), .ZN(n14901) );
  INV_X1 U10361 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n14900) );
  NOR2_X1 U10362 ( .A1(n7930), .A2(n7929), .ZN(n7931) );
  XOR2_X1 U10363 ( .A(P3_ADDR_REG_10__SCAN_IN), .B(n7931), .Z(n14903) );
  NAND2_X1 U10364 ( .A1(n15081), .A2(n15082), .ZN(n15080) );
  OAI21_X1 U10365 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(n7932), .A(n15080), .ZN(
        n7933) );
  INV_X1 U10366 ( .A(n7933), .ZN(n7935) );
  INV_X1 U10367 ( .A(n15085), .ZN(n15086) );
  NAND2_X1 U10368 ( .A1(n7935), .A2(n7934), .ZN(n15087) );
  INV_X1 U10369 ( .A(P2_ADDR_REG_12__SCAN_IN), .ZN(n15088) );
  NAND2_X1 U10370 ( .A1(n15091), .A2(n15090), .ZN(n15089) );
  NAND2_X1 U10371 ( .A1(n15099), .A2(n15098), .ZN(n7936) );
  AOI21_X1 U10372 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(n7936), .A(n15097), .ZN(
        n7937) );
  INV_X1 U10373 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n7945) );
  XOR2_X1 U10374 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(n7945), .Z(n7943) );
  OR2_X1 U10375 ( .A1(n15115), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n7938) );
  AOI22_X1 U10376 ( .A1(P3_ADDR_REG_15__SCAN_IN), .A2(n15115), .B1(n7939), 
        .B2(n7938), .ZN(n7942) );
  XOR2_X1 U10377 ( .A(n7943), .B(n7942), .Z(n7941) );
  NAND2_X1 U10378 ( .A1(n7943), .A2(n7942), .ZN(n7944) );
  OAI21_X1 U10379 ( .B1(n7945), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n7944), .ZN(
        n7948) );
  XOR2_X1 U10380 ( .A(P1_ADDR_REG_17__SCAN_IN), .B(n7948), .Z(n7949) );
  XOR2_X1 U10381 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n7949), .Z(n7947) );
  NOR2_X1 U10382 ( .A1(P1_ADDR_REG_17__SCAN_IN), .A2(n7948), .ZN(n7951) );
  AND2_X1 U10383 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n7949), .ZN(n7950) );
  NOR2_X1 U10384 ( .A1(n7951), .A2(n7950), .ZN(n8290) );
  INV_X1 U10385 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n15129) );
  XNOR2_X1 U10386 ( .A(P3_ADDR_REG_18__SCAN_IN), .B(n15129), .ZN(n8289) );
  XOR2_X1 U10387 ( .A(n8290), .B(n8289), .Z(n7953) );
  INV_X1 U10388 ( .A(SI_13_), .ZN(n10254) );
  XNOR2_X1 U10389 ( .A(n10254), .B(keyinput_g19), .ZN(n7960) );
  AOI22_X1 U10390 ( .A1(SI_16_), .A2(keyinput_g16), .B1(
        P3_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .ZN(n7954) );
  OAI221_X1 U10391 ( .B1(SI_16_), .B2(keyinput_g16), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_g60), .A(n7954), .ZN(n7959) );
  AOI22_X1 U10392 ( .A1(P3_DATAO_REG_0__SCAN_IN), .A2(keyinput_g96), .B1(
        SI_21_), .B2(keyinput_g11), .ZN(n7955) );
  OAI221_X1 U10393 ( .B1(P3_DATAO_REG_0__SCAN_IN), .B2(keyinput_g96), .C1(
        SI_21_), .C2(keyinput_g11), .A(n7955), .ZN(n7958) );
  AOI22_X1 U10394 ( .A1(P3_DATAO_REG_4__SCAN_IN), .A2(keyinput_g92), .B1(
        P3_ADDR_REG_5__SCAN_IN), .B2(keyinput_g102), .ZN(n7956) );
  OAI221_X1 U10395 ( .B1(P3_DATAO_REG_4__SCAN_IN), .B2(keyinput_g92), .C1(
        P3_ADDR_REG_5__SCAN_IN), .C2(keyinput_g102), .A(n7956), .ZN(n7957) );
  NOR4_X1 U10396 ( .A1(n7960), .A2(n7959), .A3(n7958), .A4(n7957), .ZN(n7988)
         );
  AOI22_X1 U10397 ( .A1(P3_DATAO_REG_6__SCAN_IN), .A2(keyinput_g90), .B1(
        P3_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .ZN(n7961) );
  OAI221_X1 U10398 ( .B1(P3_DATAO_REG_6__SCAN_IN), .B2(keyinput_g90), .C1(
        P3_REG3_REG_13__SCAN_IN), .C2(keyinput_g56), .A(n7961), .ZN(n7968) );
  AOI22_X1 U10399 ( .A1(P3_DATAO_REG_21__SCAN_IN), .A2(keyinput_g75), .B1(
        SI_22_), .B2(keyinput_g10), .ZN(n7962) );
  OAI221_X1 U10400 ( .B1(P3_DATAO_REG_21__SCAN_IN), .B2(keyinput_g75), .C1(
        SI_22_), .C2(keyinput_g10), .A(n7962), .ZN(n7967) );
  AOI22_X1 U10401 ( .A1(SI_2_), .A2(keyinput_g30), .B1(P3_REG3_REG_19__SCAN_IN), .B2(keyinput_g41), .ZN(n7963) );
  OAI221_X1 U10402 ( .B1(SI_2_), .B2(keyinput_g30), .C1(
        P3_REG3_REG_19__SCAN_IN), .C2(keyinput_g41), .A(n7963), .ZN(n7966) );
  AOI22_X1 U10403 ( .A1(P3_DATAO_REG_23__SCAN_IN), .A2(keyinput_g73), .B1(
        P3_STATE_REG_SCAN_IN), .B2(keyinput_g34), .ZN(n7964) );
  OAI221_X1 U10404 ( .B1(P3_DATAO_REG_23__SCAN_IN), .B2(keyinput_g73), .C1(
        P3_STATE_REG_SCAN_IN), .C2(keyinput_g34), .A(n7964), .ZN(n7965) );
  NOR4_X1 U10405 ( .A1(n7968), .A2(n7967), .A3(n7966), .A4(n7965), .ZN(n7987)
         );
  AOI22_X1 U10406 ( .A1(P3_DATAO_REG_1__SCAN_IN), .A2(keyinput_g95), .B1(
        P3_REG3_REG_27__SCAN_IN), .B2(keyinput_g36), .ZN(n7969) );
  OAI221_X1 U10407 ( .B1(P3_DATAO_REG_1__SCAN_IN), .B2(keyinput_g95), .C1(
        P3_REG3_REG_27__SCAN_IN), .C2(keyinput_g36), .A(n7969), .ZN(n7976) );
  AOI22_X1 U10408 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(SI_3_), 
        .B2(keyinput_g29), .ZN(n7970) );
  OAI221_X1 U10409 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(SI_3_), .C2(keyinput_g29), .A(n7970), .ZN(n7975) );
  AOI22_X1 U10410 ( .A1(P3_DATAO_REG_20__SCAN_IN), .A2(keyinput_g76), .B1(
        P1_IR_REG_8__SCAN_IN), .B2(keyinput_g115), .ZN(n7971) );
  OAI221_X1 U10411 ( .B1(P3_DATAO_REG_20__SCAN_IN), .B2(keyinput_g76), .C1(
        P1_IR_REG_8__SCAN_IN), .C2(keyinput_g115), .A(n7971), .ZN(n7974) );
  AOI22_X1 U10412 ( .A1(P3_DATAO_REG_3__SCAN_IN), .A2(keyinput_g93), .B1(
        SI_24_), .B2(keyinput_g8), .ZN(n7972) );
  OAI221_X1 U10413 ( .B1(P3_DATAO_REG_3__SCAN_IN), .B2(keyinput_g93), .C1(
        SI_24_), .C2(keyinput_g8), .A(n7972), .ZN(n7973) );
  NOR4_X1 U10414 ( .A1(n7976), .A2(n7975), .A3(n7974), .A4(n7973), .ZN(n7986)
         );
  AOI22_X1 U10415 ( .A1(SI_4_), .A2(keyinput_g28), .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_g57), .ZN(n7977) );
  OAI221_X1 U10416 ( .B1(SI_4_), .B2(keyinput_g28), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_g57), .A(n7977), .ZN(n7984) );
  AOI22_X1 U10417 ( .A1(P3_DATAO_REG_19__SCAN_IN), .A2(keyinput_g77), .B1(
        P1_IR_REG_18__SCAN_IN), .B2(keyinput_g125), .ZN(n7978) );
  OAI221_X1 U10418 ( .B1(P3_DATAO_REG_19__SCAN_IN), .B2(keyinput_g77), .C1(
        P1_IR_REG_18__SCAN_IN), .C2(keyinput_g125), .A(n7978), .ZN(n7983) );
  AOI22_X1 U10419 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_g46), .B1(
        P3_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n7979) );
  OAI221_X1 U10420 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n7979), .ZN(n7982) );
  AOI22_X1 U10421 ( .A1(SI_10_), .A2(keyinput_g22), .B1(SI_17_), .B2(
        keyinput_g15), .ZN(n7980) );
  OAI221_X1 U10422 ( .B1(SI_10_), .B2(keyinput_g22), .C1(SI_17_), .C2(
        keyinput_g15), .A(n7980), .ZN(n7981) );
  NOR4_X1 U10423 ( .A1(n7984), .A2(n7983), .A3(n7982), .A4(n7981), .ZN(n7985)
         );
  NAND4_X1 U10424 ( .A1(n7988), .A2(n7987), .A3(n7986), .A4(n7985), .ZN(n8116)
         );
  AOI22_X1 U10425 ( .A1(P3_DATAO_REG_2__SCAN_IN), .A2(keyinput_g94), .B1(
        P3_REG3_REG_16__SCAN_IN), .B2(keyinput_g48), .ZN(n7989) );
  OAI221_X1 U10426 ( .B1(P3_DATAO_REG_2__SCAN_IN), .B2(keyinput_g94), .C1(
        P3_REG3_REG_16__SCAN_IN), .C2(keyinput_g48), .A(n7989), .ZN(n7996) );
  AOI22_X1 U10427 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P1_IR_REG_20__SCAN_IN), .B2(keyinput_g127), .ZN(n7990) );
  OAI221_X1 U10428 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P1_IR_REG_20__SCAN_IN), .C2(keyinput_g127), .A(n7990), .ZN(n7995) );
  AOI22_X1 U10429 ( .A1(P3_DATAO_REG_9__SCAN_IN), .A2(keyinput_g87), .B1(
        SI_23_), .B2(keyinput_g9), .ZN(n7991) );
  OAI221_X1 U10430 ( .B1(P3_DATAO_REG_9__SCAN_IN), .B2(keyinput_g87), .C1(
        SI_23_), .C2(keyinput_g9), .A(n7991), .ZN(n7994) );
  AOI22_X1 U10431 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(keyinput_g104), .B1(
        SI_18_), .B2(keyinput_g14), .ZN(n7992) );
  OAI221_X1 U10432 ( .B1(P3_ADDR_REG_7__SCAN_IN), .B2(keyinput_g104), .C1(
        SI_18_), .C2(keyinput_g14), .A(n7992), .ZN(n7993) );
  NOR4_X1 U10433 ( .A1(n7996), .A2(n7995), .A3(n7994), .A4(n7993), .ZN(n8024)
         );
  AOI22_X1 U10434 ( .A1(P3_DATAO_REG_12__SCAN_IN), .A2(keyinput_g84), .B1(
        P1_IR_REG_10__SCAN_IN), .B2(keyinput_g117), .ZN(n7997) );
  OAI221_X1 U10435 ( .B1(P3_DATAO_REG_12__SCAN_IN), .B2(keyinput_g84), .C1(
        P1_IR_REG_10__SCAN_IN), .C2(keyinput_g117), .A(n7997), .ZN(n8004) );
  AOI22_X1 U10436 ( .A1(P3_REG3_REG_9__SCAN_IN), .A2(keyinput_g53), .B1(
        P3_REG3_REG_28__SCAN_IN), .B2(keyinput_g42), .ZN(n7998) );
  OAI221_X1 U10437 ( .B1(P3_REG3_REG_9__SCAN_IN), .B2(keyinput_g53), .C1(
        P3_REG3_REG_28__SCAN_IN), .C2(keyinput_g42), .A(n7998), .ZN(n8003) );
  AOI22_X1 U10438 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(keyinput_g99), .B1(SI_31_), .B2(keyinput_g1), .ZN(n7999) );
  OAI221_X1 U10439 ( .B1(P3_ADDR_REG_2__SCAN_IN), .B2(keyinput_g99), .C1(
        SI_31_), .C2(keyinput_g1), .A(n7999), .ZN(n8002) );
  AOI22_X1 U10440 ( .A1(P3_ADDR_REG_9__SCAN_IN), .A2(keyinput_g106), .B1(
        P3_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n8000) );
  OAI221_X1 U10441 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(keyinput_g106), .C1(
        P3_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n8000), .ZN(n8001) );
  NOR4_X1 U10442 ( .A1(n8004), .A2(n8003), .A3(n8002), .A4(n8001), .ZN(n8023)
         );
  AOI22_X1 U10443 ( .A1(P3_DATAO_REG_8__SCAN_IN), .A2(keyinput_g88), .B1(
        P3_ADDR_REG_4__SCAN_IN), .B2(keyinput_g101), .ZN(n8005) );
  OAI221_X1 U10444 ( .B1(P3_DATAO_REG_8__SCAN_IN), .B2(keyinput_g88), .C1(
        P3_ADDR_REG_4__SCAN_IN), .C2(keyinput_g101), .A(n8005), .ZN(n8012) );
  AOI22_X1 U10445 ( .A1(SI_20_), .A2(keyinput_g12), .B1(SI_15_), .B2(
        keyinput_g17), .ZN(n8006) );
  OAI221_X1 U10446 ( .B1(SI_20_), .B2(keyinput_g12), .C1(SI_15_), .C2(
        keyinput_g17), .A(n8006), .ZN(n8011) );
  AOI22_X1 U10447 ( .A1(P3_DATAO_REG_29__SCAN_IN), .A2(keyinput_g67), .B1(
        P1_IR_REG_0__SCAN_IN), .B2(keyinput_g107), .ZN(n8007) );
  OAI221_X1 U10448 ( .B1(P3_DATAO_REG_29__SCAN_IN), .B2(keyinput_g67), .C1(
        P1_IR_REG_0__SCAN_IN), .C2(keyinput_g107), .A(n8007), .ZN(n8010) );
  AOI22_X1 U10449 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(keyinput_g120), .B1(SI_9_), 
        .B2(keyinput_g23), .ZN(n8008) );
  OAI221_X1 U10450 ( .B1(P1_IR_REG_13__SCAN_IN), .B2(keyinput_g120), .C1(SI_9_), .C2(keyinput_g23), .A(n8008), .ZN(n8009) );
  NOR4_X1 U10451 ( .A1(n8012), .A2(n8011), .A3(n8010), .A4(n8009), .ZN(n8022)
         );
  AOI22_X1 U10452 ( .A1(P3_DATAO_REG_14__SCAN_IN), .A2(keyinput_g82), .B1(
        P1_IR_REG_14__SCAN_IN), .B2(keyinput_g121), .ZN(n8013) );
  OAI221_X1 U10453 ( .B1(P3_DATAO_REG_14__SCAN_IN), .B2(keyinput_g82), .C1(
        P1_IR_REG_14__SCAN_IN), .C2(keyinput_g121), .A(n8013), .ZN(n8020) );
  AOI22_X1 U10454 ( .A1(P3_DATAO_REG_10__SCAN_IN), .A2(keyinput_g86), .B1(
        P3_REG3_REG_11__SCAN_IN), .B2(keyinput_g58), .ZN(n8014) );
  OAI221_X1 U10455 ( .B1(P3_DATAO_REG_10__SCAN_IN), .B2(keyinput_g86), .C1(
        P3_REG3_REG_11__SCAN_IN), .C2(keyinput_g58), .A(n8014), .ZN(n8019) );
  AOI22_X1 U10456 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_g118), .B1(
        P3_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .ZN(n8015) );
  OAI221_X1 U10457 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_g118), .C1(
        P3_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n8015), .ZN(n8018) );
  INV_X1 U10458 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n10426) );
  INV_X1 U10459 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15361) );
  AOI22_X1 U10460 ( .A1(n10426), .A2(keyinput_g78), .B1(n15361), .B2(
        keyinput_g35), .ZN(n8016) );
  OAI221_X1 U10461 ( .B1(n10426), .B2(keyinput_g78), .C1(n15361), .C2(
        keyinput_g35), .A(n8016), .ZN(n8017) );
  NOR4_X1 U10462 ( .A1(n8020), .A2(n8019), .A3(n8018), .A4(n8017), .ZN(n8021)
         );
  NAND4_X1 U10463 ( .A1(n8024), .A2(n8023), .A3(n8022), .A4(n8021), .ZN(n8115)
         );
  INV_X1 U10464 ( .A(P3_DATAO_REG_5__SCAN_IN), .ZN(n10346) );
  INV_X1 U10465 ( .A(P3_DATAO_REG_22__SCAN_IN), .ZN(n10819) );
  AOI22_X1 U10466 ( .A1(n10346), .A2(keyinput_g91), .B1(n10819), .B2(
        keyinput_g74), .ZN(n8025) );
  OAI221_X1 U10467 ( .B1(n10346), .B2(keyinput_g91), .C1(n10819), .C2(
        keyinput_g74), .A(n8025), .ZN(n8033) );
  INV_X1 U10468 ( .A(P3_DATAO_REG_27__SCAN_IN), .ZN(n11443) );
  INV_X1 U10469 ( .A(P3_REG3_REG_4__SCAN_IN), .ZN(n11099) );
  AOI22_X1 U10470 ( .A1(n11443), .A2(keyinput_g69), .B1(n11099), .B2(
        keyinput_g52), .ZN(n8026) );
  OAI221_X1 U10471 ( .B1(n11443), .B2(keyinput_g69), .C1(n11099), .C2(
        keyinput_g52), .A(n8026), .ZN(n8032) );
  XNOR2_X1 U10472 ( .A(SI_14_), .B(keyinput_g18), .ZN(n8030) );
  XNOR2_X1 U10473 ( .A(SI_5_), .B(keyinput_g27), .ZN(n8029) );
  XNOR2_X1 U10474 ( .A(P3_REG3_REG_3__SCAN_IN), .B(keyinput_g40), .ZN(n8028)
         );
  XNOR2_X1 U10475 ( .A(SI_6_), .B(keyinput_g26), .ZN(n8027) );
  NAND4_X1 U10476 ( .A1(n8030), .A2(n8029), .A3(n8028), .A4(n8027), .ZN(n8031)
         );
  NOR3_X1 U10477 ( .A1(n8033), .A2(n8032), .A3(n8031), .ZN(n8070) );
  INV_X1 U10478 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n8035) );
  AOI22_X1 U10479 ( .A1(n8035), .A2(keyinput_g124), .B1(n10167), .B2(
        keyinput_g21), .ZN(n8034) );
  OAI221_X1 U10480 ( .B1(n8035), .B2(keyinput_g124), .C1(n10167), .C2(
        keyinput_g21), .A(n8034), .ZN(n8039) );
  INV_X1 U10481 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n10121) );
  XNOR2_X1 U10482 ( .A(n10121), .B(keyinput_g111), .ZN(n8038) );
  INV_X1 U10483 ( .A(P3_B_REG_SCAN_IN), .ZN(n8036) );
  XNOR2_X1 U10484 ( .A(keyinput_g64), .B(n8036), .ZN(n8037) );
  OR3_X1 U10485 ( .A1(n8039), .A2(n8038), .A3(n8037), .ZN(n8046) );
  INV_X1 U10486 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n10370) );
  XNOR2_X1 U10487 ( .A(n10370), .B(keyinput_g79), .ZN(n8045) );
  INV_X1 U10488 ( .A(P3_DATAO_REG_30__SCAN_IN), .ZN(n8040) );
  XNOR2_X1 U10489 ( .A(keyinput_g66), .B(n8040), .ZN(n8044) );
  XNOR2_X1 U10490 ( .A(SI_1_), .B(keyinput_g31), .ZN(n8042) );
  XNOR2_X1 U10491 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_g126), .ZN(n8041)
         );
  NAND2_X1 U10492 ( .A1(n8042), .A2(n8041), .ZN(n8043) );
  NOR4_X1 U10493 ( .A1(n8046), .A2(n8045), .A3(n8044), .A4(n8043), .ZN(n8069)
         );
  INV_X1 U10494 ( .A(P3_DATAO_REG_15__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U10495 ( .A1(n8245), .A2(keyinput_g98), .B1(keyinput_g81), .B2(
        n10376), .ZN(n8047) );
  OAI221_X1 U10496 ( .B1(n8245), .B2(keyinput_g98), .C1(n10376), .C2(
        keyinput_g81), .A(n8047), .ZN(n8056) );
  INV_X1 U10497 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n8049) );
  INV_X1 U10498 ( .A(SI_25_), .ZN(n12032) );
  AOI22_X1 U10499 ( .A1(n8049), .A2(keyinput_g45), .B1(keyinput_g7), .B2(
        n12032), .ZN(n8048) );
  OAI221_X1 U10500 ( .B1(n8049), .B2(keyinput_g45), .C1(n12032), .C2(
        keyinput_g7), .A(n8048), .ZN(n8055) );
  INV_X1 U10501 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n10201) );
  AOI22_X1 U10502 ( .A1(n10201), .A2(keyinput_g116), .B1(n10180), .B2(
        keyinput_g20), .ZN(n8050) );
  OAI221_X1 U10503 ( .B1(n10201), .B2(keyinput_g116), .C1(n10180), .C2(
        keyinput_g20), .A(n8050), .ZN(n8054) );
  XNOR2_X1 U10504 ( .A(P3_REG3_REG_1__SCAN_IN), .B(keyinput_g44), .ZN(n8052)
         );
  XNOR2_X1 U10505 ( .A(SI_7_), .B(keyinput_g25), .ZN(n8051) );
  NAND2_X1 U10506 ( .A1(n8052), .A2(n8051), .ZN(n8053) );
  NOR4_X1 U10507 ( .A1(n8056), .A2(n8055), .A3(n8054), .A4(n8053), .ZN(n8068)
         );
  INV_X1 U10508 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n8058) );
  AOI22_X1 U10509 ( .A1(n8058), .A2(keyinput_g61), .B1(keyinput_g103), .B2(
        n15453), .ZN(n8057) );
  OAI221_X1 U10510 ( .B1(n8058), .B2(keyinput_g61), .C1(n15453), .C2(
        keyinput_g103), .A(n8057), .ZN(n8066) );
  INV_X1 U10511 ( .A(P3_DATAO_REG_24__SCAN_IN), .ZN(n11041) );
  INV_X1 U10512 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n11615) );
  AOI22_X1 U10513 ( .A1(n11041), .A2(keyinput_g72), .B1(keyinput_g68), .B2(
        n11615), .ZN(n8059) );
  OAI221_X1 U10514 ( .B1(n11041), .B2(keyinput_g72), .C1(n11615), .C2(
        keyinput_g68), .A(n8059), .ZN(n8065) );
  INV_X1 U10515 ( .A(P3_DATAO_REG_13__SCAN_IN), .ZN(n10374) );
  INV_X1 U10516 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n11311) );
  AOI22_X1 U10517 ( .A1(n10374), .A2(keyinput_g83), .B1(n11311), .B2(
        keyinput_g59), .ZN(n8060) );
  OAI221_X1 U10518 ( .B1(n10374), .B2(keyinput_g83), .C1(n11311), .C2(
        keyinput_g59), .A(n8060), .ZN(n8064) );
  XNOR2_X1 U10519 ( .A(SI_0_), .B(keyinput_g32), .ZN(n8062) );
  XNOR2_X1 U10520 ( .A(SI_8_), .B(keyinput_g24), .ZN(n8061) );
  NAND2_X1 U10521 ( .A1(n8062), .A2(n8061), .ZN(n8063) );
  NOR4_X1 U10522 ( .A1(n8066), .A2(n8065), .A3(n8064), .A4(n8063), .ZN(n8067)
         );
  NAND4_X1 U10523 ( .A1(n8070), .A2(n8069), .A3(n8068), .A4(n8067), .ZN(n8114)
         );
  INV_X1 U10524 ( .A(SI_27_), .ZN(n12215) );
  INV_X1 U10525 ( .A(SI_26_), .ZN(n12139) );
  AOI22_X1 U10526 ( .A1(n12215), .A2(keyinput_g5), .B1(keyinput_g6), .B2(
        n12139), .ZN(n8071) );
  OAI221_X1 U10527 ( .B1(n12215), .B2(keyinput_g5), .C1(n12139), .C2(
        keyinput_g6), .A(n8071), .ZN(n8079) );
  INV_X1 U10528 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n10368) );
  INV_X1 U10529 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15368) );
  AOI22_X1 U10530 ( .A1(n10368), .A2(keyinput_g89), .B1(n15368), .B2(
        keyinput_g39), .ZN(n8072) );
  OAI221_X1 U10531 ( .B1(n10368), .B2(keyinput_g89), .C1(n15368), .C2(
        keyinput_g39), .A(n8072), .ZN(n8078) );
  XNOR2_X1 U10532 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_g112), .ZN(n8075) );
  XNOR2_X1 U10533 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_g109), .ZN(n8074) );
  XNOR2_X1 U10534 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_g122), .ZN(n8073)
         );
  NAND3_X1 U10535 ( .A1(n8075), .A2(n8074), .A3(n8073), .ZN(n8077) );
  INV_X1 U10536 ( .A(P3_RD_REG_SCAN_IN), .ZN(n14885) );
  XNOR2_X1 U10537 ( .A(n14885), .B(keyinput_g33), .ZN(n8076) );
  NOR4_X1 U10538 ( .A1(n8079), .A2(n8078), .A3(n8077), .A4(n8076), .ZN(n8112)
         );
  INV_X1 U10539 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n10280) );
  AOI22_X1 U10540 ( .A1(n10280), .A2(keyinput_g119), .B1(n8486), .B2(
        keyinput_g43), .ZN(n8080) );
  OAI221_X1 U10541 ( .B1(n10280), .B2(keyinput_g119), .C1(n8486), .C2(
        keyinput_g43), .A(n8080), .ZN(n8083) );
  INV_X1 U10542 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n11617) );
  XNOR2_X1 U10543 ( .A(n11617), .B(keyinput_g65), .ZN(n8082) );
  INV_X1 U10544 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n10874) );
  XNOR2_X1 U10545 ( .A(n10874), .B(keyinput_g123), .ZN(n8081) );
  OR3_X1 U10546 ( .A1(n8083), .A2(n8082), .A3(n8081), .ZN(n8089) );
  INV_X1 U10547 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n10372) );
  INV_X1 U10548 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n8370) );
  AOI22_X1 U10549 ( .A1(n10372), .A2(keyinput_g80), .B1(n8370), .B2(
        keyinput_g50), .ZN(n8084) );
  OAI221_X1 U10550 ( .B1(n10372), .B2(keyinput_g80), .C1(n8370), .C2(
        keyinput_g50), .A(n8084), .ZN(n8088) );
  INV_X1 U10551 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n8086) );
  INV_X1 U10552 ( .A(SI_30_), .ZN(n13132) );
  AOI22_X1 U10553 ( .A1(n8086), .A2(keyinput_g47), .B1(keyinput_g2), .B2(
        n13132), .ZN(n8085) );
  OAI221_X1 U10554 ( .B1(n8086), .B2(keyinput_g47), .C1(n13132), .C2(
        keyinput_g2), .A(n8085), .ZN(n8087) );
  NOR3_X1 U10555 ( .A1(n8089), .A2(n8088), .A3(n8087), .ZN(n8111) );
  INV_X1 U10556 ( .A(SI_28_), .ZN(n12946) );
  INV_X1 U10557 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n8230) );
  AOI22_X1 U10558 ( .A1(n12946), .A2(keyinput_g4), .B1(n8230), .B2(
        keyinput_g51), .ZN(n8090) );
  OAI221_X1 U10559 ( .B1(n12946), .B2(keyinput_g4), .C1(n8230), .C2(
        keyinput_g51), .A(n8090), .ZN(n8099) );
  INV_X1 U10560 ( .A(SI_29_), .ZN(n13689) );
  AOI22_X1 U10561 ( .A1(n13689), .A2(keyinput_g3), .B1(keyinput_g13), .B2(
        n10767), .ZN(n8091) );
  OAI221_X1 U10562 ( .B1(n13689), .B2(keyinput_g3), .C1(n10767), .C2(
        keyinput_g13), .A(n8091), .ZN(n8098) );
  INV_X1 U10563 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n8092) );
  XOR2_X1 U10564 ( .A(n8092), .B(keyinput_g49), .Z(n8096) );
  XNOR2_X1 U10565 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_g108), .ZN(n8095) );
  XNOR2_X1 U10566 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_g113), .ZN(n8094) );
  XNOR2_X1 U10567 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_g110), .ZN(n8093) );
  NAND4_X1 U10568 ( .A1(n8096), .A2(n8095), .A3(n8094), .A4(n8093), .ZN(n8097)
         );
  NOR3_X1 U10569 ( .A1(n8099), .A2(n8098), .A3(n8097), .ZN(n8110) );
  INV_X1 U10570 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n13199) );
  INV_X1 U10571 ( .A(P3_DATAO_REG_25__SCAN_IN), .ZN(n11107) );
  AOI22_X1 U10572 ( .A1(n13199), .A2(keyinput_g38), .B1(keyinput_g71), .B2(
        n11107), .ZN(n8100) );
  OAI221_X1 U10573 ( .B1(n13199), .B2(keyinput_g38), .C1(n11107), .C2(
        keyinput_g71), .A(n8100), .ZN(n8108) );
  INV_X1 U10574 ( .A(P3_DATAO_REG_11__SCAN_IN), .ZN(n10366) );
  AOI22_X1 U10575 ( .A1(n10366), .A2(keyinput_g85), .B1(n8246), .B2(
        keyinput_g100), .ZN(n8101) );
  OAI221_X1 U10576 ( .B1(n10366), .B2(keyinput_g85), .C1(n8246), .C2(
        keyinput_g100), .A(n8101), .ZN(n8107) );
  INV_X1 U10577 ( .A(P3_DATAO_REG_26__SCAN_IN), .ZN(n11219) );
  AOI22_X1 U10578 ( .A1(n10957), .A2(keyinput_g97), .B1(keyinput_g70), .B2(
        n11219), .ZN(n8102) );
  OAI221_X1 U10579 ( .B1(n10957), .B2(keyinput_g97), .C1(n11219), .C2(
        keyinput_g70), .A(n8102), .ZN(n8106) );
  XNOR2_X1 U10580 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_g114), .ZN(n8104) );
  XNOR2_X1 U10581 ( .A(P3_REG3_REG_26__SCAN_IN), .B(keyinput_g62), .ZN(n8103)
         );
  NAND2_X1 U10582 ( .A1(n8104), .A2(n8103), .ZN(n8105) );
  NOR4_X1 U10583 ( .A1(n8108), .A2(n8107), .A3(n8106), .A4(n8105), .ZN(n8109)
         );
  NAND4_X1 U10584 ( .A1(n8112), .A2(n8111), .A3(n8110), .A4(n8109), .ZN(n8113)
         );
  NOR4_X1 U10585 ( .A1(n8116), .A2(n8115), .A3(n8114), .A4(n8113), .ZN(n8287)
         );
  AOI22_X1 U10586 ( .A1(keyinput_f75), .A2(P3_DATAO_REG_21__SCAN_IN), .B1(
        P3_ADDR_REG_5__SCAN_IN), .B2(keyinput_f102), .ZN(n8117) );
  OAI221_X1 U10587 ( .B1(keyinput_f75), .B2(P3_DATAO_REG_21__SCAN_IN), .C1(
        P3_ADDR_REG_5__SCAN_IN), .C2(keyinput_f102), .A(n8117), .ZN(n8124) );
  AOI22_X1 U10588 ( .A1(keyinput_f80), .A2(P3_DATAO_REG_16__SCAN_IN), .B1(
        SI_31_), .B2(keyinput_f1), .ZN(n8118) );
  OAI221_X1 U10589 ( .B1(keyinput_f80), .B2(P3_DATAO_REG_16__SCAN_IN), .C1(
        SI_31_), .C2(keyinput_f1), .A(n8118), .ZN(n8123) );
  AOI22_X1 U10590 ( .A1(SI_30_), .A2(keyinput_f2), .B1(P3_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n8119) );
  OAI221_X1 U10591 ( .B1(SI_30_), .B2(keyinput_f2), .C1(
        P3_REG3_REG_11__SCAN_IN), .C2(keyinput_f58), .A(n8119), .ZN(n8122) );
  AOI22_X1 U10592 ( .A1(keyinput_f81), .A2(P3_DATAO_REG_15__SCAN_IN), .B1(
        P3_REG3_REG_25__SCAN_IN), .B2(keyinput_f47), .ZN(n8120) );
  OAI221_X1 U10593 ( .B1(keyinput_f81), .B2(P3_DATAO_REG_15__SCAN_IN), .C1(
        P3_REG3_REG_25__SCAN_IN), .C2(keyinput_f47), .A(n8120), .ZN(n8121) );
  NOR4_X1 U10594 ( .A1(n8124), .A2(n8123), .A3(n8122), .A4(n8121), .ZN(n8280)
         );
  INV_X1 U10595 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n8126) );
  AOI22_X1 U10596 ( .A1(SI_0_), .A2(keyinput_f32), .B1(n8126), .B2(
        keyinput_f36), .ZN(n8125) );
  OAI221_X1 U10597 ( .B1(SI_0_), .B2(keyinput_f32), .C1(n8126), .C2(
        keyinput_f36), .A(n8125), .ZN(n8134) );
  AOI22_X1 U10598 ( .A1(SI_10_), .A2(keyinput_f22), .B1(
        P3_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .ZN(n8127) );
  OAI221_X1 U10599 ( .B1(SI_10_), .B2(keyinput_f22), .C1(
        P3_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(n8127), .ZN(n8133) );
  XNOR2_X1 U10600 ( .A(n14885), .B(keyinput_f33), .ZN(n8132) );
  XNOR2_X1 U10601 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_f123), .ZN(n8130)
         );
  XNOR2_X1 U10602 ( .A(SI_1_), .B(keyinput_f31), .ZN(n8129) );
  XNOR2_X1 U10603 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_f120), .ZN(n8128)
         );
  NAND3_X1 U10604 ( .A1(n8130), .A2(n8129), .A3(n8128), .ZN(n8131) );
  NOR4_X1 U10605 ( .A1(n8134), .A2(n8133), .A3(n8132), .A4(n8131), .ZN(n8279)
         );
  INV_X1 U10606 ( .A(SI_23_), .ZN(n11447) );
  OAI22_X1 U10607 ( .A1(n11447), .A2(keyinput_f9), .B1(n10819), .B2(
        keyinput_f74), .ZN(n8135) );
  AOI221_X1 U10608 ( .B1(n11447), .B2(keyinput_f9), .C1(keyinput_f74), .C2(
        n10819), .A(n8135), .ZN(n8144) );
  INV_X1 U10609 ( .A(P3_DATAO_REG_4__SCAN_IN), .ZN(n10344) );
  OAI22_X1 U10610 ( .A1(n8364), .A2(keyinput_f46), .B1(n10344), .B2(
        keyinput_f92), .ZN(n8136) );
  AOI221_X1 U10611 ( .B1(n8364), .B2(keyinput_f46), .C1(keyinput_f92), .C2(
        n10344), .A(n8136), .ZN(n8143) );
  INV_X1 U10612 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n8138) );
  OAI22_X1 U10613 ( .A1(n8138), .A2(keyinput_f37), .B1(n6885), .B2(
        keyinput_f10), .ZN(n8137) );
  AOI221_X1 U10614 ( .B1(n8138), .B2(keyinput_f37), .C1(keyinput_f10), .C2(
        n6885), .A(n8137), .ZN(n8142) );
  XNOR2_X1 U10615 ( .A(n10280), .B(keyinput_f119), .ZN(n8140) );
  INV_X1 U10616 ( .A(P1_IR_REG_3__SCAN_IN), .ZN(n10146) );
  XNOR2_X1 U10617 ( .A(n10146), .B(keyinput_f110), .ZN(n8139) );
  NOR2_X1 U10618 ( .A1(n8140), .A2(n8139), .ZN(n8141) );
  NAND4_X1 U10619 ( .A1(n8144), .A2(n8143), .A3(n8142), .A4(n8141), .ZN(n8156)
         );
  INV_X1 U10620 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n8146) );
  AOI22_X1 U10621 ( .A1(n8146), .A2(keyinput_f62), .B1(keyinput_f43), .B2(
        n8486), .ZN(n8145) );
  OAI221_X1 U10622 ( .B1(n8146), .B2(keyinput_f62), .C1(n8486), .C2(
        keyinput_f43), .A(n8145), .ZN(n8155) );
  INV_X1 U10623 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n13247) );
  AOI22_X1 U10624 ( .A1(n10532), .A2(keyinput_f15), .B1(n13247), .B2(
        keyinput_f48), .ZN(n8147) );
  OAI221_X1 U10625 ( .B1(n10532), .B2(keyinput_f15), .C1(n13247), .C2(
        keyinput_f48), .A(n8147), .ZN(n8154) );
  INV_X1 U10626 ( .A(SI_24_), .ZN(n12890) );
  INV_X1 U10627 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n8149) );
  OAI22_X1 U10628 ( .A1(n8149), .A2(keyinput_f122), .B1(n10374), .B2(
        keyinput_f83), .ZN(n8148) );
  AOI221_X1 U10629 ( .B1(n8149), .B2(keyinput_f122), .C1(keyinput_f83), .C2(
        n10374), .A(n8148), .ZN(n8152) );
  INV_X1 U10630 ( .A(P3_DATAO_REG_8__SCAN_IN), .ZN(n10364) );
  XNOR2_X1 U10631 ( .A(keyinput_f88), .B(n10364), .ZN(n8150) );
  AOI21_X1 U10632 ( .B1(keyinput_f8), .B2(n12890), .A(n8150), .ZN(n8151) );
  OAI211_X1 U10633 ( .C1(keyinput_f8), .C2(n12890), .A(n8152), .B(n8151), .ZN(
        n8153) );
  NOR4_X1 U10634 ( .A1(n8156), .A2(n8155), .A3(n8154), .A4(n8153), .ZN(n8278)
         );
  OAI22_X1 U10635 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(keyinput_f121), .B1(
        P3_DATAO_REG_17__SCAN_IN), .B2(keyinput_f79), .ZN(n8157) );
  AOI221_X1 U10636 ( .B1(P1_IR_REG_14__SCAN_IN), .B2(keyinput_f121), .C1(
        keyinput_f79), .C2(P3_DATAO_REG_17__SCAN_IN), .A(n8157), .ZN(n8164) );
  OAI22_X1 U10637 ( .A1(keyinput_f95), .A2(P3_DATAO_REG_1__SCAN_IN), .B1(
        keyinput_f65), .B2(P3_DATAO_REG_31__SCAN_IN), .ZN(n8158) );
  AOI221_X1 U10638 ( .B1(keyinput_f95), .B2(P3_DATAO_REG_1__SCAN_IN), .C1(
        P3_DATAO_REG_31__SCAN_IN), .C2(keyinput_f65), .A(n8158), .ZN(n8163) );
  OAI22_X1 U10639 ( .A1(P3_REG3_REG_17__SCAN_IN), .A2(keyinput_f50), .B1(
        keyinput_f86), .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n8159) );
  AOI221_X1 U10640 ( .B1(P3_REG3_REG_17__SCAN_IN), .B2(keyinput_f50), .C1(
        P3_DATAO_REG_10__SCAN_IN), .C2(keyinput_f86), .A(n8159), .ZN(n8162) );
  OAI22_X1 U10641 ( .A1(P3_ADDR_REG_0__SCAN_IN), .A2(keyinput_f97), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(keyinput_f66), .ZN(n8160) );
  AOI221_X1 U10642 ( .B1(P3_ADDR_REG_0__SCAN_IN), .B2(keyinput_f97), .C1(
        keyinput_f66), .C2(P3_DATAO_REG_30__SCAN_IN), .A(n8160), .ZN(n8161) );
  NAND4_X1 U10643 ( .A1(n8164), .A2(n8163), .A3(n8162), .A4(n8161), .ZN(n8276)
         );
  AOI22_X1 U10644 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(keyinput_f61), .B1(
        P3_REG3_REG_21__SCAN_IN), .B2(keyinput_f45), .ZN(n8165) );
  OAI221_X1 U10645 ( .B1(P3_REG3_REG_6__SCAN_IN), .B2(keyinput_f61), .C1(
        P3_REG3_REG_21__SCAN_IN), .C2(keyinput_f45), .A(n8165), .ZN(n8172) );
  AOI22_X1 U10646 ( .A1(keyinput_f89), .A2(P3_DATAO_REG_7__SCAN_IN), .B1(
        P1_IR_REG_5__SCAN_IN), .B2(keyinput_f112), .ZN(n8166) );
  OAI221_X1 U10647 ( .B1(keyinput_f89), .B2(P3_DATAO_REG_7__SCAN_IN), .C1(
        P1_IR_REG_5__SCAN_IN), .C2(keyinput_f112), .A(n8166), .ZN(n8171) );
  AOI22_X1 U10648 ( .A1(SI_14_), .A2(keyinput_f18), .B1(SI_28_), .B2(
        keyinput_f4), .ZN(n8167) );
  OAI221_X1 U10649 ( .B1(SI_14_), .B2(keyinput_f18), .C1(SI_28_), .C2(
        keyinput_f4), .A(n8167), .ZN(n8170) );
  AOI22_X1 U10650 ( .A1(SI_25_), .A2(keyinput_f7), .B1(P3_REG3_REG_9__SCAN_IN), 
        .B2(keyinput_f53), .ZN(n8168) );
  OAI221_X1 U10651 ( .B1(SI_25_), .B2(keyinput_f7), .C1(P3_REG3_REG_9__SCAN_IN), .C2(keyinput_f53), .A(n8168), .ZN(n8169) );
  NOR4_X1 U10652 ( .A1(n8172), .A2(n8171), .A3(n8170), .A4(n8169), .ZN(n8190)
         );
  AOI22_X1 U10653 ( .A1(keyinput_f87), .A2(P3_DATAO_REG_9__SCAN_IN), .B1(
        P3_ADDR_REG_4__SCAN_IN), .B2(keyinput_f101), .ZN(n8173) );
  OAI221_X1 U10654 ( .B1(keyinput_f87), .B2(P3_DATAO_REG_9__SCAN_IN), .C1(
        P3_ADDR_REG_4__SCAN_IN), .C2(keyinput_f101), .A(n8173), .ZN(n8180) );
  AOI22_X1 U10655 ( .A1(keyinput_f78), .A2(P3_DATAO_REG_18__SCAN_IN), .B1(
        P1_IR_REG_6__SCAN_IN), .B2(keyinput_f113), .ZN(n8174) );
  OAI221_X1 U10656 ( .B1(keyinput_f78), .B2(P3_DATAO_REG_18__SCAN_IN), .C1(
        P1_IR_REG_6__SCAN_IN), .C2(keyinput_f113), .A(n8174), .ZN(n8179) );
  AOI22_X1 U10657 ( .A1(SI_15_), .A2(keyinput_f17), .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_f44), .ZN(n8175) );
  OAI221_X1 U10658 ( .B1(SI_15_), .B2(keyinput_f17), .C1(
        P3_REG3_REG_1__SCAN_IN), .C2(keyinput_f44), .A(n8175), .ZN(n8178) );
  AOI22_X1 U10659 ( .A1(SI_18_), .A2(keyinput_f14), .B1(
        P3_REG3_REG_13__SCAN_IN), .B2(keyinput_f56), .ZN(n8176) );
  OAI221_X1 U10660 ( .B1(SI_18_), .B2(keyinput_f14), .C1(
        P3_REG3_REG_13__SCAN_IN), .C2(keyinput_f56), .A(n8176), .ZN(n8177) );
  NOR4_X1 U10661 ( .A1(n8180), .A2(n8179), .A3(n8178), .A4(n8177), .ZN(n8189)
         );
  OAI22_X1 U10662 ( .A1(P3_REG3_REG_23__SCAN_IN), .A2(keyinput_f38), .B1(
        keyinput_f73), .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n8181) );
  AOI221_X1 U10663 ( .B1(P3_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .C1(
        P3_DATAO_REG_23__SCAN_IN), .C2(keyinput_f73), .A(n8181), .ZN(n8187) );
  OAI22_X1 U10664 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(keyinput_f49), .B1(
        keyinput_f72), .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n8182) );
  AOI221_X1 U10665 ( .B1(P3_REG3_REG_5__SCAN_IN), .B2(keyinput_f49), .C1(
        P3_DATAO_REG_24__SCAN_IN), .C2(keyinput_f72), .A(n8182), .ZN(n8186) );
  OAI22_X1 U10666 ( .A1(P1_IR_REG_4__SCAN_IN), .A2(keyinput_f111), .B1(
        P3_DATAO_REG_2__SCAN_IN), .B2(keyinput_f94), .ZN(n8183) );
  AOI221_X1 U10667 ( .B1(P1_IR_REG_4__SCAN_IN), .B2(keyinput_f111), .C1(
        keyinput_f94), .C2(P3_DATAO_REG_2__SCAN_IN), .A(n8183), .ZN(n8185) );
  XNOR2_X1 U10668 ( .A(SI_9_), .B(keyinput_f23), .ZN(n8184) );
  AND4_X1 U10669 ( .A1(n8187), .A2(n8186), .A3(n8185), .A4(n8184), .ZN(n8188)
         );
  NAND3_X1 U10670 ( .A1(n8190), .A2(n8189), .A3(n8188), .ZN(n8275) );
  AOI22_X1 U10671 ( .A1(keyinput_f96), .A2(P3_DATAO_REG_0__SCAN_IN), .B1(SI_2_), .B2(keyinput_f30), .ZN(n8191) );
  OAI221_X1 U10672 ( .B1(keyinput_f96), .B2(P3_DATAO_REG_0__SCAN_IN), .C1(
        SI_2_), .C2(keyinput_f30), .A(n8191), .ZN(n8198) );
  AOI22_X1 U10673 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(keyinput_f99), .B1(
        P1_IR_REG_7__SCAN_IN), .B2(keyinput_f114), .ZN(n8192) );
  OAI221_X1 U10674 ( .B1(P3_ADDR_REG_2__SCAN_IN), .B2(keyinput_f99), .C1(
        P1_IR_REG_7__SCAN_IN), .C2(keyinput_f114), .A(n8192), .ZN(n8197) );
  AOI22_X1 U10675 ( .A1(P1_IR_REG_11__SCAN_IN), .A2(keyinput_f118), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(keyinput_f35), .ZN(n8193) );
  OAI221_X1 U10676 ( .B1(P1_IR_REG_11__SCAN_IN), .B2(keyinput_f118), .C1(
        P3_REG3_REG_7__SCAN_IN), .C2(keyinput_f35), .A(n8193), .ZN(n8196) );
  AOI22_X1 U10677 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(keyinput_f124), .B1(
        P1_IR_REG_19__SCAN_IN), .B2(keyinput_f126), .ZN(n8194) );
  OAI221_X1 U10678 ( .B1(P1_IR_REG_17__SCAN_IN), .B2(keyinput_f124), .C1(
        P1_IR_REG_19__SCAN_IN), .C2(keyinput_f126), .A(n8194), .ZN(n8195) );
  NOR4_X1 U10679 ( .A1(n8198), .A2(n8197), .A3(n8196), .A4(n8195), .ZN(n8226)
         );
  AOI22_X1 U10680 ( .A1(keyinput_f84), .A2(P3_DATAO_REG_12__SCAN_IN), .B1(
        P3_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .ZN(n8199) );
  OAI221_X1 U10681 ( .B1(keyinput_f84), .B2(P3_DATAO_REG_12__SCAN_IN), .C1(
        P3_REG3_REG_10__SCAN_IN), .C2(keyinput_f39), .A(n8199), .ZN(n8206) );
  AOI22_X1 U10682 ( .A1(keyinput_f90), .A2(P3_DATAO_REG_6__SCAN_IN), .B1(
        P3_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .ZN(n8200) );
  OAI221_X1 U10683 ( .B1(keyinput_f90), .B2(P3_DATAO_REG_6__SCAN_IN), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput_f55), .A(n8200), .ZN(n8205) );
  AOI22_X1 U10684 ( .A1(keyinput_f76), .A2(P3_DATAO_REG_20__SCAN_IN), .B1(
        SI_29_), .B2(keyinput_f3), .ZN(n8201) );
  OAI221_X1 U10685 ( .B1(keyinput_f76), .B2(P3_DATAO_REG_20__SCAN_IN), .C1(
        SI_29_), .C2(keyinput_f3), .A(n8201), .ZN(n8204) );
  AOI22_X1 U10686 ( .A1(keyinput_f85), .A2(P3_DATAO_REG_11__SCAN_IN), .B1(
        SI_6_), .B2(keyinput_f26), .ZN(n8202) );
  OAI221_X1 U10687 ( .B1(keyinput_f85), .B2(P3_DATAO_REG_11__SCAN_IN), .C1(
        SI_6_), .C2(keyinput_f26), .A(n8202), .ZN(n8203) );
  NOR4_X1 U10688 ( .A1(n8206), .A2(n8205), .A3(n8204), .A4(n8203), .ZN(n8225)
         );
  AOI22_X1 U10689 ( .A1(P3_ADDR_REG_9__SCAN_IN), .A2(keyinput_f106), .B1(
        SI_11_), .B2(keyinput_f21), .ZN(n8207) );
  OAI221_X1 U10690 ( .B1(P3_ADDR_REG_9__SCAN_IN), .B2(keyinput_f106), .C1(
        SI_11_), .C2(keyinput_f21), .A(n8207), .ZN(n8214) );
  AOI22_X1 U10691 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(keyinput_f104), .B1(
        P1_IR_REG_2__SCAN_IN), .B2(keyinput_f109), .ZN(n8208) );
  OAI221_X1 U10692 ( .B1(P3_ADDR_REG_7__SCAN_IN), .B2(keyinput_f104), .C1(
        P1_IR_REG_2__SCAN_IN), .C2(keyinput_f109), .A(n8208), .ZN(n8213) );
  AOI22_X1 U10693 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(keyinput_f125), .B1(
        P3_B_REG_SCAN_IN), .B2(keyinput_f64), .ZN(n8209) );
  OAI221_X1 U10694 ( .B1(P1_IR_REG_18__SCAN_IN), .B2(keyinput_f125), .C1(
        P3_B_REG_SCAN_IN), .C2(keyinput_f64), .A(n8209), .ZN(n8212) );
  AOI22_X1 U10695 ( .A1(SI_12_), .A2(keyinput_f20), .B1(SI_27_), .B2(
        keyinput_f5), .ZN(n8210) );
  OAI221_X1 U10696 ( .B1(SI_12_), .B2(keyinput_f20), .C1(SI_27_), .C2(
        keyinput_f5), .A(n8210), .ZN(n8211) );
  NOR4_X1 U10697 ( .A1(n8214), .A2(n8213), .A3(n8212), .A4(n8211), .ZN(n8224)
         );
  AOI22_X1 U10698 ( .A1(SI_7_), .A2(keyinput_f25), .B1(P3_REG3_REG_4__SCAN_IN), 
        .B2(keyinput_f52), .ZN(n8215) );
  OAI221_X1 U10699 ( .B1(SI_7_), .B2(keyinput_f25), .C1(P3_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n8215), .ZN(n8222) );
  AOI22_X1 U10700 ( .A1(keyinput_f67), .A2(P3_DATAO_REG_29__SCAN_IN), .B1(
        P3_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .ZN(n8216) );
  OAI221_X1 U10701 ( .B1(keyinput_f67), .B2(P3_DATAO_REG_29__SCAN_IN), .C1(
        P3_REG3_REG_15__SCAN_IN), .C2(keyinput_f63), .A(n8216), .ZN(n8221) );
  AOI22_X1 U10702 ( .A1(keyinput_f77), .A2(P3_DATAO_REG_19__SCAN_IN), .B1(
        SI_26_), .B2(keyinput_f6), .ZN(n8217) );
  OAI221_X1 U10703 ( .B1(keyinput_f77), .B2(P3_DATAO_REG_19__SCAN_IN), .C1(
        SI_26_), .C2(keyinput_f6), .A(n8217), .ZN(n8220) );
  AOI22_X1 U10704 ( .A1(keyinput_f70), .A2(P3_DATAO_REG_26__SCAN_IN), .B1(
        P3_STATE_REG_SCAN_IN), .B2(keyinput_f34), .ZN(n8218) );
  OAI221_X1 U10705 ( .B1(keyinput_f70), .B2(P3_DATAO_REG_26__SCAN_IN), .C1(
        P3_STATE_REG_SCAN_IN), .C2(keyinput_f34), .A(n8218), .ZN(n8219) );
  NOR4_X1 U10706 ( .A1(n8222), .A2(n8221), .A3(n8220), .A4(n8219), .ZN(n8223)
         );
  NAND4_X1 U10707 ( .A1(n8226), .A2(n8225), .A3(n8224), .A4(n8223), .ZN(n8274)
         );
  INV_X1 U10708 ( .A(keyinput_f0), .ZN(n8228) );
  AOI22_X1 U10709 ( .A1(n15453), .A2(keyinput_f103), .B1(P3_WR_REG_SCAN_IN), 
        .B2(n8228), .ZN(n8227) );
  OAI221_X1 U10710 ( .B1(n15453), .B2(keyinput_f103), .C1(n8228), .C2(
        P3_WR_REG_SCAN_IN), .A(n8227), .ZN(n8238) );
  INV_X1 U10711 ( .A(P1_IR_REG_10__SCAN_IN), .ZN(n8231) );
  AOI22_X1 U10712 ( .A1(n8231), .A2(keyinput_f117), .B1(n8230), .B2(
        keyinput_f51), .ZN(n8229) );
  OAI221_X1 U10713 ( .B1(n8231), .B2(keyinput_f117), .C1(n8230), .C2(
        keyinput_f51), .A(n8229), .ZN(n8237) );
  INV_X1 U10714 ( .A(P3_DATAO_REG_3__SCAN_IN), .ZN(n10348) );
  AOI22_X1 U10715 ( .A1(n10348), .A2(keyinput_f93), .B1(n10767), .B2(
        keyinput_f13), .ZN(n8232) );
  OAI221_X1 U10716 ( .B1(n10348), .B2(keyinput_f93), .C1(n10767), .C2(
        keyinput_f13), .A(n8232), .ZN(n8236) );
  XNOR2_X1 U10717 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_f115), .ZN(n8234) );
  XNOR2_X1 U10718 ( .A(SI_5_), .B(keyinput_f27), .ZN(n8233) );
  NAND2_X1 U10719 ( .A1(n8234), .A2(n8233), .ZN(n8235) );
  NOR4_X1 U10720 ( .A1(n8238), .A2(n8237), .A3(n8236), .A4(n8235), .ZN(n8272)
         );
  INV_X1 U10721 ( .A(SI_20_), .ZN(n11038) );
  INV_X1 U10722 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U10723 ( .A1(n11038), .A2(keyinput_f12), .B1(n10958), .B2(
        keyinput_f54), .ZN(n8239) );
  OAI221_X1 U10724 ( .B1(n11038), .B2(keyinput_f12), .C1(n10958), .C2(
        keyinput_f54), .A(n8239), .ZN(n8243) );
  XNOR2_X1 U10725 ( .A(n10346), .B(keyinput_f91), .ZN(n8242) );
  XOR2_X1 U10726 ( .A(SI_4_), .B(keyinput_f28), .Z(n8241) );
  XNOR2_X1 U10727 ( .A(n7593), .B(keyinput_f107), .ZN(n8240) );
  OR4_X1 U10728 ( .A1(n8243), .A2(n8242), .A3(n8241), .A4(n8240), .ZN(n8249)
         );
  INV_X1 U10729 ( .A(P3_DATAO_REG_14__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U10730 ( .A1(n10350), .A2(keyinput_f82), .B1(n8245), .B2(
        keyinput_f98), .ZN(n8244) );
  OAI221_X1 U10731 ( .B1(n10350), .B2(keyinput_f82), .C1(n8245), .C2(
        keyinput_f98), .A(n8244), .ZN(n8248) );
  XNOR2_X1 U10732 ( .A(n8246), .B(keyinput_f100), .ZN(n8247) );
  NOR3_X1 U10733 ( .A1(n8249), .A2(n8248), .A3(n8247), .ZN(n8271) );
  INV_X1 U10734 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n13207) );
  AOI22_X1 U10735 ( .A1(n13207), .A2(keyinput_f41), .B1(keyinput_f68), .B2(
        n11615), .ZN(n8250) );
  OAI221_X1 U10736 ( .B1(n13207), .B2(keyinput_f41), .C1(n11615), .C2(
        keyinput_f68), .A(n8250), .ZN(n8259) );
  AOI22_X1 U10737 ( .A1(n11443), .A2(keyinput_f69), .B1(n10254), .B2(
        keyinput_f19), .ZN(n8251) );
  OAI221_X1 U10738 ( .B1(n11443), .B2(keyinput_f69), .C1(n10254), .C2(
        keyinput_f19), .A(n8251), .ZN(n8258) );
  INV_X1 U10739 ( .A(P3_REG3_REG_18__SCAN_IN), .ZN(n14932) );
  AOI22_X1 U10740 ( .A1(n14932), .A2(keyinput_f60), .B1(keyinput_f59), .B2(
        n11311), .ZN(n8252) );
  OAI221_X1 U10741 ( .B1(n14932), .B2(keyinput_f60), .C1(n11311), .C2(
        keyinput_f59), .A(n8252), .ZN(n8257) );
  INV_X1 U10742 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n8253) );
  XOR2_X1 U10743 ( .A(n8253), .B(keyinput_f42), .Z(n8255) );
  XNOR2_X1 U10744 ( .A(SI_8_), .B(keyinput_f24), .ZN(n8254) );
  NAND2_X1 U10745 ( .A1(n8255), .A2(n8254), .ZN(n8256) );
  NOR4_X1 U10746 ( .A1(n8259), .A2(n8258), .A3(n8257), .A4(n8256), .ZN(n8270)
         );
  INV_X1 U10747 ( .A(SI_21_), .ZN(n11137) );
  AOI22_X1 U10748 ( .A1(n11107), .A2(keyinput_f71), .B1(n11137), .B2(
        keyinput_f11), .ZN(n8260) );
  OAI221_X1 U10749 ( .B1(n11107), .B2(keyinput_f71), .C1(n11137), .C2(
        keyinput_f11), .A(n8260), .ZN(n8268) );
  INV_X1 U10750 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n10117) );
  XNOR2_X1 U10751 ( .A(n10117), .B(keyinput_f108), .ZN(n8267) );
  INV_X1 U10752 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n11758) );
  XNOR2_X1 U10753 ( .A(n11758), .B(keyinput_f40), .ZN(n8266) );
  XNOR2_X1 U10754 ( .A(SI_3_), .B(keyinput_f29), .ZN(n8264) );
  XNOR2_X1 U10755 ( .A(SI_16_), .B(keyinput_f16), .ZN(n8263) );
  XNOR2_X1 U10756 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_f127), .ZN(n8262)
         );
  XNOR2_X1 U10757 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_f116), .ZN(n8261) );
  NAND4_X1 U10758 ( .A1(n8264), .A2(n8263), .A3(n8262), .A4(n8261), .ZN(n8265)
         );
  NOR4_X1 U10759 ( .A1(n8268), .A2(n8267), .A3(n8266), .A4(n8265), .ZN(n8269)
         );
  NAND4_X1 U10760 ( .A1(n8272), .A2(n8271), .A3(n8270), .A4(n8269), .ZN(n8273)
         );
  NOR4_X1 U10761 ( .A1(n8276), .A2(n8275), .A3(n8274), .A4(n8273), .ZN(n8277)
         );
  NAND4_X1 U10762 ( .A1(n8280), .A2(n8279), .A3(n8278), .A4(n8277), .ZN(n8282)
         );
  INV_X1 U10763 ( .A(keyinput_g105), .ZN(n8284) );
  AOI21_X1 U10764 ( .B1(keyinput_f105), .B2(n8282), .A(n8284), .ZN(n8285) );
  INV_X1 U10765 ( .A(keyinput_f105), .ZN(n8281) );
  AOI21_X1 U10766 ( .B1(n8282), .B2(n8281), .A(P3_ADDR_REG_8__SCAN_IN), .ZN(
        n8283) );
  AOI22_X1 U10767 ( .A1(P3_ADDR_REG_8__SCAN_IN), .A2(n8285), .B1(n8284), .B2(
        n8283), .ZN(n8286) );
  NOR2_X1 U10768 ( .A1(n8287), .A2(n8286), .ZN(n8288) );
  NOR2_X1 U10769 ( .A1(n8290), .A2(n8289), .ZN(n8291) );
  AOI21_X1 U10770 ( .B1(P3_ADDR_REG_18__SCAN_IN), .B2(n15129), .A(n8291), .ZN(
        n8294) );
  XNOR2_X1 U10771 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n8292) );
  XNOR2_X1 U10772 ( .A(n8292), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n8293) );
  INV_X1 U10773 ( .A(n8411), .ZN(n8296) );
  NAND2_X1 U10774 ( .A1(n8412), .A2(n8296), .ZN(n8298) );
  NAND2_X1 U10775 ( .A1(n10171), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n8297) );
  NAND2_X1 U10776 ( .A1(n8298), .A2(n8297), .ZN(n8418) );
  NAND2_X1 U10777 ( .A1(n10183), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n8300) );
  INV_X1 U10778 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n10823) );
  NAND2_X1 U10779 ( .A1(n10823), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n8299) );
  AND2_X1 U10780 ( .A1(n8300), .A2(n8299), .ZN(n8417) );
  NAND2_X1 U10781 ( .A1(n8418), .A2(n8417), .ZN(n8301) );
  NAND2_X1 U10782 ( .A1(n10979), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8302) );
  NAND2_X1 U10783 ( .A1(n8428), .A2(n8427), .ZN(n8304) );
  NAND2_X2 U10784 ( .A1(n8304), .A2(n8303), .ZN(n8440) );
  NAND2_X1 U10785 ( .A1(n11220), .A2(P1_DATAO_REG_4__SCAN_IN), .ZN(n8305) );
  NAND2_X1 U10786 ( .A1(n11326), .A2(P1_DATAO_REG_5__SCAN_IN), .ZN(n8307) );
  NAND2_X1 U10787 ( .A1(n10144), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n8309) );
  NAND2_X1 U10788 ( .A1(n10189), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n8310) );
  NAND2_X1 U10789 ( .A1(n10198), .A2(P2_DATAO_REG_7__SCAN_IN), .ZN(n8312) );
  NAND2_X1 U10790 ( .A1(n8313), .A2(n8312), .ZN(n8476) );
  NAND2_X1 U10791 ( .A1(n10175), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n8315) );
  NAND2_X1 U10792 ( .A1(n10195), .A2(P2_DATAO_REG_8__SCAN_IN), .ZN(n8314) );
  NAND2_X1 U10793 ( .A1(n10179), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n8317) );
  NAND2_X1 U10794 ( .A1(n10192), .A2(P2_DATAO_REG_9__SCAN_IN), .ZN(n8316) );
  NAND2_X1 U10795 ( .A1(n10205), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n8319) );
  NAND2_X1 U10796 ( .A1(n10200), .A2(P2_DATAO_REG_10__SCAN_IN), .ZN(n8318) );
  NAND2_X2 U10797 ( .A1(n8521), .A2(n8520), .ZN(n8523) );
  NAND2_X1 U10798 ( .A1(n10240), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n8321) );
  INV_X1 U10799 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n10233) );
  NAND2_X1 U10800 ( .A1(n10233), .A2(P2_DATAO_REG_11__SCAN_IN), .ZN(n8320) );
  NAND2_X1 U10801 ( .A1(n10259), .A2(P1_DATAO_REG_12__SCAN_IN), .ZN(n8323) );
  INV_X1 U10802 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n10261) );
  NAND2_X1 U10803 ( .A1(n10261), .A2(P2_DATAO_REG_12__SCAN_IN), .ZN(n8322) );
  INV_X1 U10804 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10536) );
  NAND2_X1 U10805 ( .A1(n10536), .A2(P1_DATAO_REG_14__SCAN_IN), .ZN(n8328) );
  INV_X1 U10806 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n10539) );
  NAND2_X1 U10807 ( .A1(n10539), .A2(P2_DATAO_REG_14__SCAN_IN), .ZN(n8327) );
  NAND2_X1 U10808 ( .A1(n10763), .A2(P1_DATAO_REG_15__SCAN_IN), .ZN(n8330) );
  NAND2_X1 U10809 ( .A1(n10766), .A2(P2_DATAO_REG_15__SCAN_IN), .ZN(n8329) );
  AND2_X1 U10810 ( .A1(n8330), .A2(n8329), .ZN(n8580) );
  NAND2_X1 U10811 ( .A1(n10879), .A2(P1_DATAO_REG_16__SCAN_IN), .ZN(n8332) );
  NAND2_X1 U10812 ( .A1(n10871), .A2(P2_DATAO_REG_16__SCAN_IN), .ZN(n8331) );
  AND2_X1 U10813 ( .A1(n8332), .A2(n8331), .ZN(n8593) );
  INV_X1 U10814 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n10974) );
  NAND2_X1 U10815 ( .A1(n10974), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n8334) );
  INV_X1 U10816 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n10971) );
  NAND2_X1 U10817 ( .A1(n10971), .A2(P2_DATAO_REG_17__SCAN_IN), .ZN(n8333) );
  AND2_X1 U10818 ( .A1(n8334), .A2(n8333), .ZN(n8607) );
  NAND2_X1 U10819 ( .A1(n11112), .A2(P1_DATAO_REG_18__SCAN_IN), .ZN(n8336) );
  NAND2_X1 U10820 ( .A1(n11113), .A2(P2_DATAO_REG_18__SCAN_IN), .ZN(n8335) );
  AND2_X1 U10821 ( .A1(n8336), .A2(n8335), .ZN(n8619) );
  INV_X1 U10822 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n11284) );
  NAND2_X1 U10823 ( .A1(n11284), .A2(P1_DATAO_REG_19__SCAN_IN), .ZN(n8338) );
  INV_X1 U10824 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n11286) );
  NAND2_X1 U10825 ( .A1(n11286), .A2(P2_DATAO_REG_19__SCAN_IN), .ZN(n8337) );
  AND2_X1 U10826 ( .A1(n8338), .A2(n8337), .ZN(n8632) );
  NAND2_X2 U10827 ( .A1(n8633), .A2(n8632), .ZN(n8635) );
  INV_X1 U10828 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n12723) );
  NAND2_X1 U10829 ( .A1(n12723), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n8341) );
  INV_X1 U10830 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n11512) );
  NAND2_X1 U10831 ( .A1(n11512), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n8340) );
  AND2_X1 U10832 ( .A1(n8341), .A2(n8340), .ZN(n8659) );
  INV_X1 U10833 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n11557) );
  XNOR2_X1 U10834 ( .A(n11557), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n8673) );
  NAND2_X1 U10835 ( .A1(n11557), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n8342) );
  XNOR2_X1 U10836 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .ZN(n8686) );
  INV_X1 U10837 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11818) );
  INV_X1 U10838 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n12142) );
  NAND2_X1 U10839 ( .A1(n8343), .A2(n12142), .ZN(n8344) );
  INV_X1 U10840 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n12327) );
  NAND2_X1 U10841 ( .A1(n12327), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n8346) );
  INV_X1 U10842 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n12772) );
  NAND2_X1 U10843 ( .A1(n12772), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n8347) );
  INV_X1 U10844 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n12383) );
  NOR2_X1 U10845 ( .A1(n12383), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8348) );
  NAND2_X1 U10846 ( .A1(n12383), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n8349) );
  INV_X1 U10847 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n12888) );
  AND2_X1 U10848 ( .A1(n12888), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n8351) );
  INV_X1 U10849 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14875) );
  NAND2_X1 U10850 ( .A1(n14875), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n8352) );
  INV_X1 U10851 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n14200) );
  NOR2_X1 U10852 ( .A1(n14200), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n8353) );
  XNOR2_X1 U10853 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n8758) );
  INV_X1 U10854 ( .A(n8758), .ZN(n8354) );
  INV_X1 U10855 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n14193) );
  INV_X1 U10856 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n13120) );
  XNOR2_X1 U10857 ( .A(n13120), .B(P2_DATAO_REG_30__SCAN_IN), .ZN(n8390) );
  XNOR2_X1 U10858 ( .A(n8391), .B(n8390), .ZN(n13130) );
  NAND3_X1 U10859 ( .A1(n14887), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n8358) );
  NAND2_X1 U10860 ( .A1(n8358), .A2(n8357), .ZN(n8359) );
  NAND2_X1 U10861 ( .A1(n13130), .A2(n8760), .ZN(n8363) );
  OR2_X1 U10862 ( .A1(n8761), .A2(n13132), .ZN(n8362) );
  INV_X1 U10863 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n8366) );
  INV_X1 U10864 ( .A(P3_REG3_REG_15__SCAN_IN), .ZN(n8368) );
  INV_X1 U10865 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n8377) );
  INV_X1 U10866 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n13676) );
  XNOR2_X2 U10867 ( .A(n8379), .B(n13676), .ZN(n13133) );
  NAND2_X1 U10868 ( .A1(n8380), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8381) );
  AND2_X2 U10869 ( .A1(n8383), .A2(n8384), .ZN(n8449) );
  NAND2_X1 U10870 ( .A1(n13123), .A2(n8757), .ZN(n8770) );
  INV_X1 U10871 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n8387) );
  NAND2_X1 U10872 ( .A1(n8736), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8386) );
  NAND2_X1 U10873 ( .A1(n8737), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8385) );
  OAI211_X1 U10874 ( .C1(n8767), .C2(n8387), .A(n8386), .B(n8385), .ZN(n8388)
         );
  INV_X1 U10875 ( .A(n8388), .ZN(n8389) );
  NOR2_X1 U10876 ( .A1(n8773), .A2(n11375), .ZN(n8930) );
  INV_X1 U10877 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n12886) );
  OAI22_X1 U10878 ( .A1(n8391), .A2(n8390), .B1(P1_DATAO_REG_30__SCAN_IN), 
        .B2(n12886), .ZN(n8393) );
  XNOR2_X1 U10879 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .ZN(n8392) );
  XNOR2_X1 U10880 ( .A(n8393), .B(n8392), .ZN(n13682) );
  NAND2_X1 U10881 ( .A1(n13682), .A2(n8760), .ZN(n8395) );
  INV_X1 U10882 ( .A(SI_31_), .ZN(n13677) );
  OR2_X1 U10883 ( .A1(n8761), .A2(n13677), .ZN(n8394) );
  NAND2_X1 U10884 ( .A1(n8600), .A2(P3_REG1_REG_31__SCAN_IN), .ZN(n8398) );
  NAND2_X1 U10885 ( .A1(n6813), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n8397) );
  NAND2_X1 U10886 ( .A1(n8752), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n8396) );
  AND3_X1 U10887 ( .A1(n8398), .A2(n8397), .A3(n8396), .ZN(n8399) );
  NAND2_X1 U10888 ( .A1(n8668), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8403) );
  NAND2_X1 U10889 ( .A1(n8764), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n8402) );
  NAND2_X1 U10890 ( .A1(n8449), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n8401) );
  NAND2_X1 U10891 ( .A1(n8600), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n8400) );
  INV_X1 U10892 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n8404) );
  NAND2_X1 U10893 ( .A1(n8404), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n8405) );
  NAND2_X1 U10894 ( .A1(n8411), .A2(n8405), .ZN(n8406) );
  MUX2_X1 U10895 ( .A(n8406), .B(SI_0_), .S(n9213), .Z(n13691) );
  MUX2_X1 U10896 ( .A(P3_IR_REG_0__SCAN_IN), .B(n13691), .S(n8361), .Z(n11011)
         );
  INV_X1 U10897 ( .A(n11011), .ZN(n10680) );
  NOR2_X2 U10898 ( .A1(n13330), .A2(n10680), .ZN(n10770) );
  NAND2_X1 U10899 ( .A1(n8764), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n8410) );
  NAND2_X1 U10900 ( .A1(n8668), .A2(P3_REG2_REG_1__SCAN_IN), .ZN(n8409) );
  NAND2_X1 U10901 ( .A1(n8449), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n8408) );
  NAND2_X1 U10902 ( .A1(n8600), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n8407) );
  AND4_X2 U10903 ( .A1(n8409), .A2(n8410), .A3(n8408), .A4(n8407), .ZN(n8955)
         );
  INV_X1 U10904 ( .A(n8955), .ZN(n13328) );
  INV_X1 U10905 ( .A(SI_1_), .ZN(n10159) );
  XNOR2_X1 U10906 ( .A(n8412), .B(n8411), .ZN(n10158) );
  INV_X1 U10907 ( .A(n10719), .ZN(n8956) );
  NAND2_X1 U10908 ( .A1(n13328), .A2(n8956), .ZN(n8804) );
  NAND2_X1 U10909 ( .A1(n8955), .A2(n10719), .ZN(n10708) );
  NAND2_X1 U10910 ( .A1(n8668), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8416) );
  NAND2_X1 U10911 ( .A1(n8764), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n8415) );
  NAND2_X1 U10912 ( .A1(n8449), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n8414) );
  NAND2_X1 U10913 ( .A1(n8600), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8413) );
  XNOR2_X1 U10914 ( .A(n8418), .B(n8417), .ZN(n10148) );
  OR2_X1 U10915 ( .A1(n8663), .A2(n10148), .ZN(n8420) );
  NAND2_X1 U10916 ( .A1(n8636), .A2(n7766), .ZN(n8419) );
  INV_X1 U10917 ( .A(n11309), .ZN(n8953) );
  NAND2_X1 U10918 ( .A1(n13327), .A2(n8953), .ZN(n8809) );
  NAND2_X1 U10919 ( .A1(n8952), .A2(n11309), .ZN(n8812) );
  NAND2_X1 U10920 ( .A1(n8668), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n8426) );
  NAND2_X1 U10921 ( .A1(n8764), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n8425) );
  NAND2_X1 U10922 ( .A1(n8449), .A2(n11758), .ZN(n8424) );
  NAND2_X1 U10923 ( .A1(n8600), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n8423) );
  OR2_X1 U10924 ( .A1(n8761), .A2(SI_3_), .ZN(n8432) );
  XNOR2_X1 U10925 ( .A(n8428), .B(n8427), .ZN(n10125) );
  OR2_X1 U10926 ( .A1(n8663), .A2(n10125), .ZN(n8431) );
  NAND2_X1 U10927 ( .A1(n8636), .A2(n8429), .ZN(n8430) );
  NAND2_X1 U10928 ( .A1(n11304), .A2(n11759), .ZN(n8813) );
  INV_X1 U10929 ( .A(n11759), .ZN(n15539) );
  NAND2_X1 U10930 ( .A1(n11750), .A2(n11753), .ZN(n8433) );
  NAND2_X1 U10931 ( .A1(n8752), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n8438) );
  NAND2_X1 U10932 ( .A1(n8668), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n8437) );
  AND2_X1 U10933 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n8434) );
  OR2_X1 U10934 ( .A1(n8434), .A2(n8447), .ZN(n11747) );
  NAND2_X1 U10935 ( .A1(n8449), .A2(n11747), .ZN(n8436) );
  NAND2_X1 U10936 ( .A1(n8600), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n8435) );
  OR2_X1 U10937 ( .A1(n8761), .A2(SI_4_), .ZN(n8443) );
  XNOR2_X1 U10938 ( .A(n8440), .B(n8439), .ZN(n10130) );
  OR2_X1 U10939 ( .A1(n8663), .A2(n10130), .ZN(n8442) );
  NAND2_X1 U10940 ( .A1(n8636), .A2(n15417), .ZN(n8441) );
  NAND2_X1 U10941 ( .A1(n11755), .A2(n15545), .ZN(n8821) );
  INV_X1 U10942 ( .A(n15545), .ZN(n8444) );
  NAND2_X1 U10943 ( .A1(n11543), .A2(n8444), .ZN(n8824) );
  INV_X1 U10944 ( .A(n11742), .ZN(n8445) );
  NAND2_X1 U10945 ( .A1(n11740), .A2(n8445), .ZN(n8446) );
  NAND2_X1 U10946 ( .A1(n8446), .A2(n8821), .ZN(n11545) );
  NAND2_X1 U10947 ( .A1(n8737), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n8453) );
  NAND2_X1 U10948 ( .A1(n8668), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n8452) );
  OR2_X1 U10949 ( .A1(n8447), .A2(n8092), .ZN(n8448) );
  NAND2_X1 U10950 ( .A1(n8459), .A2(n8448), .ZN(n11549) );
  NAND2_X1 U10951 ( .A1(n8757), .A2(n11549), .ZN(n8451) );
  NAND2_X1 U10952 ( .A1(n8600), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n8450) );
  OR2_X1 U10953 ( .A1(n8761), .A2(SI_5_), .ZN(n8458) );
  XNOR2_X1 U10954 ( .A(n8455), .B(n8454), .ZN(n10127) );
  OR2_X1 U10955 ( .A1(n6879), .A2(n15434), .ZN(n8456) );
  NAND2_X1 U10956 ( .A1(n11767), .A2(n11550), .ZN(n11763) );
  NAND2_X1 U10957 ( .A1(n11181), .A2(n15550), .ZN(n8822) );
  NAND2_X1 U10958 ( .A1(n8737), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n8464) );
  NAND2_X1 U10959 ( .A1(n8600), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8463) );
  NAND2_X1 U10960 ( .A1(n8459), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n8460) );
  AND2_X1 U10961 ( .A1(n8469), .A2(n8460), .ZN(n15402) );
  INV_X1 U10962 ( .A(n15402), .ZN(n11773) );
  NAND2_X1 U10963 ( .A1(n8757), .A2(n11773), .ZN(n8462) );
  NAND2_X1 U10964 ( .A1(n8668), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n8461) );
  INV_X1 U10965 ( .A(SI_6_), .ZN(n10161) );
  OR2_X1 U10966 ( .A1(n8761), .A2(n10161), .ZN(n8468) );
  XNOR2_X1 U10967 ( .A(n10189), .B(P2_DATAO_REG_6__SCAN_IN), .ZN(n8465) );
  XNOR2_X1 U10968 ( .A(n8466), .B(n8465), .ZN(n10162) );
  OR2_X1 U10969 ( .A1(n8663), .A2(n10162), .ZN(n8467) );
  OAI211_X1 U10970 ( .C1(n6879), .C2(n15442), .A(n8468), .B(n8467), .ZN(n15560) );
  NAND2_X1 U10971 ( .A1(n11942), .A2(n15560), .ZN(n8830) );
  AND2_X1 U10972 ( .A1(n11763), .A2(n8830), .ZN(n11935) );
  NAND2_X1 U10973 ( .A1(n8668), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n8475) );
  NAND2_X1 U10974 ( .A1(n8752), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n8474) );
  AND2_X1 U10975 ( .A1(n8469), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n8470) );
  NOR2_X1 U10976 ( .A1(n8487), .A2(n8470), .ZN(n15367) );
  INV_X1 U10977 ( .A(n15367), .ZN(n8471) );
  NAND2_X1 U10978 ( .A1(n8757), .A2(n8471), .ZN(n8473) );
  NAND2_X1 U10979 ( .A1(n8600), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n8472) );
  OR2_X1 U10980 ( .A1(n8761), .A2(SI_7_), .ZN(n8482) );
  NAND2_X1 U10981 ( .A1(n8477), .A2(n8476), .ZN(n8478) );
  AND2_X1 U10982 ( .A1(n8479), .A2(n8478), .ZN(n10123) );
  OR2_X1 U10983 ( .A1(n8663), .A2(n10123), .ZN(n8481) );
  OR2_X1 U10984 ( .A1(n6879), .A2(n15464), .ZN(n8480) );
  NAND2_X1 U10985 ( .A1(n11780), .A2(n8966), .ZN(n8834) );
  INV_X1 U10986 ( .A(n8966), .ZN(n15563) );
  NAND2_X1 U10987 ( .A1(n11714), .A2(n15563), .ZN(n8835) );
  INV_X1 U10988 ( .A(n11940), .ZN(n8781) );
  INV_X1 U10989 ( .A(n11942), .ZN(n13326) );
  INV_X1 U10990 ( .A(n15560), .ZN(n15398) );
  NAND2_X1 U10991 ( .A1(n13326), .A2(n15398), .ZN(n11937) );
  AND2_X1 U10992 ( .A1(n8781), .A2(n11937), .ZN(n8483) );
  NAND2_X1 U10993 ( .A1(n8484), .A2(n8483), .ZN(n8485) );
  NAND2_X1 U10994 ( .A1(n8764), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n8492) );
  NAND2_X1 U10995 ( .A1(n8600), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n8491) );
  NOR2_X1 U10996 ( .A1(n8487), .A2(n8486), .ZN(n8488) );
  OR2_X1 U10997 ( .A1(n8500), .A2(n8488), .ZN(n11708) );
  NAND2_X1 U10998 ( .A1(n8757), .A2(n11708), .ZN(n8490) );
  NAND2_X1 U10999 ( .A1(n6813), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n8489) );
  OR2_X1 U11000 ( .A1(n8494), .A2(n8493), .ZN(n8495) );
  NAND2_X1 U11001 ( .A1(n8496), .A2(n8495), .ZN(n10157) );
  OR2_X1 U11002 ( .A1(n8663), .A2(n10157), .ZN(n8498) );
  INV_X1 U11003 ( .A(SI_8_), .ZN(n10156) );
  OR2_X1 U11004 ( .A1(n8761), .A2(n10156), .ZN(n8497) );
  OAI211_X1 U11005 ( .C1(n6879), .C2(n15483), .A(n8498), .B(n8497), .ZN(n11721) );
  NAND2_X1 U11006 ( .A1(n12013), .A2(n11721), .ZN(n8839) );
  INV_X1 U11007 ( .A(n11721), .ZN(n15569) );
  NAND2_X1 U11008 ( .A1(n12004), .A2(n15569), .ZN(n8846) );
  NAND2_X1 U11009 ( .A1(n11776), .A2(n11778), .ZN(n8499) );
  NAND2_X1 U11010 ( .A1(n8737), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n8505) );
  NAND2_X1 U11011 ( .A1(n6813), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n8504) );
  OR2_X1 U11012 ( .A1(n8500), .A2(n12012), .ZN(n8501) );
  NAND2_X1 U11013 ( .A1(n8513), .A2(n8501), .ZN(n12016) );
  NAND2_X1 U11014 ( .A1(n8757), .A2(n12016), .ZN(n8503) );
  NAND2_X1 U11015 ( .A1(n8736), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n8502) );
  NAND4_X1 U11016 ( .A1(n8505), .A2(n8504), .A3(n8503), .A4(n8502), .ZN(n13325) );
  OR2_X1 U11017 ( .A1(n8507), .A2(n8506), .ZN(n8508) );
  AND2_X1 U11018 ( .A1(n8509), .A2(n8508), .ZN(n10152) );
  OR2_X1 U11019 ( .A1(n8663), .A2(n10152), .ZN(n8512) );
  OR2_X1 U11020 ( .A1(n8761), .A2(SI_9_), .ZN(n8511) );
  OR2_X1 U11021 ( .A1(n6879), .A2(n10153), .ZN(n8510) );
  NOR2_X1 U11022 ( .A1(n13325), .A2(n15575), .ZN(n8847) );
  NAND2_X1 U11023 ( .A1(n13325), .A2(n15575), .ZN(n8840) );
  NAND2_X1 U11024 ( .A1(n8752), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n8519) );
  NAND2_X1 U11025 ( .A1(n8736), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n8518) );
  NAND2_X1 U11026 ( .A1(n8513), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n8514) );
  AND2_X1 U11027 ( .A1(n8528), .A2(n8514), .ZN(n15380) );
  INV_X1 U11028 ( .A(n15380), .ZN(n8515) );
  NAND2_X1 U11029 ( .A1(n8757), .A2(n8515), .ZN(n8517) );
  NAND2_X1 U11030 ( .A1(n6813), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n8516) );
  OR2_X1 U11031 ( .A1(n8521), .A2(n8520), .ZN(n8522) );
  NAND2_X1 U11032 ( .A1(n8523), .A2(n8522), .ZN(n10165) );
  NAND2_X1 U11033 ( .A1(n8760), .A2(n10165), .ZN(n8526) );
  OR2_X1 U11034 ( .A1(n8761), .A2(SI_10_), .ZN(n8525) );
  NAND2_X1 U11035 ( .A1(n8636), .A2(n10163), .ZN(n8524) );
  INV_X1 U11036 ( .A(n15378), .ZN(n15581) );
  NAND2_X1 U11037 ( .A1(n13324), .A2(n15581), .ZN(n8842) );
  NAND2_X1 U11038 ( .A1(n12223), .A2(n15378), .ZN(n8850) );
  NAND2_X1 U11039 ( .A1(n8527), .A2(n8850), .ZN(n12053) );
  NAND2_X1 U11040 ( .A1(n6813), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n8533) );
  NAND2_X1 U11041 ( .A1(n8764), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n8532) );
  NAND2_X1 U11042 ( .A1(n8528), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n8529) );
  NAND2_X1 U11043 ( .A1(n8540), .A2(n8529), .ZN(n12234) );
  NAND2_X1 U11044 ( .A1(n8757), .A2(n12234), .ZN(n8531) );
  NAND2_X1 U11045 ( .A1(n8736), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n8530) );
  OR2_X1 U11046 ( .A1(n8535), .A2(n8534), .ZN(n8536) );
  NAND2_X1 U11047 ( .A1(n8537), .A2(n8536), .ZN(n10169) );
  NAND2_X1 U11048 ( .A1(n10169), .A2(n8760), .ZN(n8539) );
  AOI22_X1 U11049 ( .A1(n8637), .A2(n10167), .B1(n8636), .B2(n10168), .ZN(
        n8538) );
  NAND2_X1 U11050 ( .A1(n8539), .A2(n8538), .ZN(n14953) );
  XNOR2_X1 U11051 ( .A(n12398), .B(n12054), .ZN(n12052) );
  NAND2_X1 U11052 ( .A1(n12390), .A2(n12054), .ZN(n8843) );
  NAND2_X1 U11053 ( .A1(n8752), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U11054 ( .A1(n6813), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n8544) );
  NAND2_X1 U11055 ( .A1(n8540), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n8541) );
  NAND2_X1 U11056 ( .A1(n8559), .A2(n8541), .ZN(n12039) );
  NAND2_X1 U11057 ( .A1(n8757), .A2(n12039), .ZN(n8543) );
  NAND2_X1 U11058 ( .A1(n8736), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n8542) );
  OR2_X1 U11059 ( .A1(n8547), .A2(n8546), .ZN(n8548) );
  NAND2_X1 U11060 ( .A1(n8549), .A2(n8548), .ZN(n10181) );
  OR2_X1 U11061 ( .A1(n10181), .A2(n8663), .ZN(n8552) );
  AOI22_X1 U11062 ( .A1(n8637), .A2(SI_12_), .B1(n8636), .B2(n8550), .ZN(n8551) );
  NAND2_X1 U11063 ( .A1(n8552), .A2(n8551), .ZN(n14948) );
  OR2_X1 U11064 ( .A1(n12388), .A2(n14948), .ZN(n8856) );
  NAND2_X1 U11065 ( .A1(n14948), .A2(n12388), .ZN(n8855) );
  NAND2_X1 U11066 ( .A1(n12042), .A2(n6740), .ZN(n8553) );
  NAND2_X1 U11067 ( .A1(n8554), .A2(n10278), .ZN(n8555) );
  NAND2_X1 U11068 ( .A1(n8556), .A2(n8555), .ZN(n10255) );
  NAND2_X1 U11069 ( .A1(n10255), .A2(n8760), .ZN(n8558) );
  AOI22_X1 U11070 ( .A1(n8637), .A2(n10254), .B1(n8636), .B2(n10253), .ZN(
        n8557) );
  NAND2_X1 U11071 ( .A1(n8558), .A2(n8557), .ZN(n14943) );
  NAND2_X1 U11072 ( .A1(n6813), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n8564) );
  NAND2_X1 U11073 ( .A1(n8737), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n8563) );
  NAND2_X1 U11074 ( .A1(n8559), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n8560) );
  NAND2_X1 U11075 ( .A1(n8572), .A2(n8560), .ZN(n12438) );
  NAND2_X1 U11076 ( .A1(n8757), .A2(n12438), .ZN(n8562) );
  NAND2_X1 U11077 ( .A1(n8736), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n8561) );
  NAND4_X1 U11078 ( .A1(n8564), .A2(n8563), .A3(n8562), .A4(n8561), .ZN(n13186) );
  OR2_X1 U11079 ( .A1(n14943), .A2(n13186), .ZN(n8860) );
  INV_X1 U11080 ( .A(n8860), .ZN(n8565) );
  NAND2_X1 U11081 ( .A1(n14943), .A2(n13186), .ZN(n8861) );
  OR2_X1 U11082 ( .A1(n8567), .A2(n8566), .ZN(n8568) );
  NAND2_X1 U11083 ( .A1(n8569), .A2(n8568), .ZN(n10277) );
  NAND2_X1 U11084 ( .A1(n10277), .A2(n8760), .ZN(n8571) );
  INV_X1 U11085 ( .A(SI_14_), .ZN(n10276) );
  AOI22_X1 U11086 ( .A1(n8637), .A2(n10276), .B1(n8636), .B2(n15519), .ZN(
        n8570) );
  NAND2_X1 U11087 ( .A1(n8571), .A2(n8570), .ZN(n14938) );
  NAND2_X1 U11088 ( .A1(n6813), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8577) );
  NAND2_X1 U11089 ( .A1(n8764), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n8576) );
  NAND2_X1 U11090 ( .A1(n8572), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n8573) );
  NAND2_X1 U11091 ( .A1(n8586), .A2(n8573), .ZN(n13190) );
  NAND2_X1 U11092 ( .A1(n8757), .A2(n13190), .ZN(n8575) );
  NAND2_X1 U11093 ( .A1(n8600), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8574) );
  NAND4_X1 U11094 ( .A1(n8577), .A2(n8576), .A3(n8575), .A4(n8574), .ZN(n13312) );
  NAND2_X1 U11095 ( .A1(n14938), .A2(n13312), .ZN(n8866) );
  OR2_X1 U11096 ( .A1(n14938), .A2(n13312), .ZN(n8867) );
  OR2_X1 U11097 ( .A1(n8581), .A2(n8580), .ZN(n8582) );
  NAND2_X1 U11098 ( .A1(n8583), .A2(n8582), .ZN(n10317) );
  NAND2_X1 U11099 ( .A1(n10317), .A2(n8760), .ZN(n8585) );
  INV_X1 U11100 ( .A(n13361), .ZN(n10315) );
  AOI22_X1 U11101 ( .A1(n8637), .A2(n10316), .B1(n8636), .B2(n10315), .ZN(
        n8584) );
  NAND2_X1 U11102 ( .A1(n8737), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n8591) );
  NAND2_X1 U11103 ( .A1(n8736), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n8590) );
  NAND2_X1 U11104 ( .A1(n8586), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n8587) );
  NAND2_X1 U11105 ( .A1(n8601), .A2(n8587), .ZN(n13318) );
  NAND2_X1 U11106 ( .A1(n8757), .A2(n13318), .ZN(n8589) );
  NAND2_X1 U11107 ( .A1(n6813), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n8588) );
  NAND4_X1 U11108 ( .A1(n8591), .A2(n8590), .A3(n8589), .A4(n8588), .ZN(n13140) );
  NAND2_X1 U11109 ( .A1(n14933), .A2(n13140), .ZN(n8865) );
  NAND2_X1 U11110 ( .A1(n8873), .A2(n8865), .ZN(n12329) );
  INV_X1 U11111 ( .A(n12329), .ZN(n8863) );
  NAND2_X1 U11112 ( .A1(n12328), .A2(n8863), .ZN(n8592) );
  OR2_X1 U11113 ( .A1(n8594), .A2(n8593), .ZN(n8595) );
  NAND2_X1 U11114 ( .A1(n8596), .A2(n8595), .ZN(n10443) );
  OR2_X1 U11115 ( .A1(n10443), .A2(n8663), .ZN(n8599) );
  AOI22_X1 U11116 ( .A1(n8637), .A2(SI_16_), .B1(n8636), .B2(n8597), .ZN(n8598) );
  NAND2_X1 U11117 ( .A1(n8752), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n8606) );
  NAND2_X1 U11118 ( .A1(n8600), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n8605) );
  NAND2_X1 U11119 ( .A1(n8601), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n8602) );
  NAND2_X1 U11120 ( .A1(n8613), .A2(n8602), .ZN(n13250) );
  NAND2_X1 U11121 ( .A1(n8757), .A2(n13250), .ZN(n8604) );
  NAND2_X1 U11122 ( .A1(n6813), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n8603) );
  NAND4_X1 U11123 ( .A1(n8606), .A2(n8605), .A3(n8604), .A4(n8603), .ZN(n13256) );
  INV_X1 U11124 ( .A(n13256), .ZN(n13316) );
  OR2_X1 U11125 ( .A1(n13143), .A2(n13316), .ZN(n8875) );
  NAND2_X1 U11126 ( .A1(n13143), .A2(n13316), .ZN(n8874) );
  OR2_X1 U11127 ( .A1(n8608), .A2(n8607), .ZN(n8609) );
  NAND2_X1 U11128 ( .A1(n8610), .A2(n8609), .ZN(n10533) );
  NAND2_X1 U11129 ( .A1(n10533), .A2(n8760), .ZN(n8612) );
  AOI22_X1 U11130 ( .A1(n8637), .A2(n10532), .B1(n8636), .B2(n10531), .ZN(
        n8611) );
  NAND2_X1 U11131 ( .A1(n6813), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n8618) );
  NAND2_X1 U11132 ( .A1(n8764), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n8617) );
  NAND2_X1 U11133 ( .A1(n8613), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n8614) );
  NAND2_X1 U11134 ( .A1(n8625), .A2(n8614), .ZN(n13558) );
  NAND2_X1 U11135 ( .A1(n8757), .A2(n13558), .ZN(n8616) );
  NAND2_X1 U11136 ( .A1(n8736), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n8615) );
  NAND4_X1 U11137 ( .A1(n8618), .A2(n8617), .A3(n8616), .A4(n8615), .ZN(n13532) );
  NAND2_X1 U11138 ( .A1(n13670), .A2(n13532), .ZN(n8882) );
  INV_X1 U11139 ( .A(n13547), .ZN(n8631) );
  OR2_X1 U11140 ( .A1(n8620), .A2(n8619), .ZN(n8621) );
  NAND2_X1 U11141 ( .A1(n8622), .A2(n8621), .ZN(n10542) );
  AOI22_X1 U11142 ( .A1(n8637), .A2(SI_18_), .B1(n8636), .B2(n14917), .ZN(
        n8623) );
  NAND2_X1 U11143 ( .A1(n8737), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n8630) );
  NAND2_X1 U11144 ( .A1(n6813), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n8629) );
  NAND2_X1 U11145 ( .A1(n8625), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n8626) );
  NAND2_X1 U11146 ( .A1(n8640), .A2(n8626), .ZN(n13537) );
  NAND2_X1 U11147 ( .A1(n8757), .A2(n13537), .ZN(n8628) );
  NAND2_X1 U11148 ( .A1(n8736), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n8627) );
  NAND2_X1 U11149 ( .A1(n13544), .A2(n13517), .ZN(n8884) );
  OR2_X1 U11150 ( .A1(n8633), .A2(n8632), .ZN(n8634) );
  NAND2_X1 U11151 ( .A1(n8635), .A2(n8634), .ZN(n10769) );
  OR2_X1 U11152 ( .A1(n10769), .A2(n8663), .ZN(n8639) );
  AOI22_X1 U11153 ( .A1(n8637), .A2(SI_19_), .B1(n9014), .B2(n8636), .ZN(n8638) );
  NAND2_X1 U11154 ( .A1(n8640), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n8641) );
  NAND2_X1 U11155 ( .A1(n8654), .A2(n8641), .ZN(n13523) );
  NAND2_X1 U11156 ( .A1(n13523), .A2(n8757), .ZN(n8645) );
  NAND2_X1 U11157 ( .A1(n6813), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n8643) );
  NAND2_X1 U11158 ( .A1(n8752), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n8642) );
  AND2_X1 U11159 ( .A1(n8643), .A2(n8642), .ZN(n8644) );
  OAI211_X1 U11160 ( .C1(n8646), .C2(n13607), .A(n8645), .B(n8644), .ZN(n13534) );
  NOR2_X1 U11161 ( .A1(n13153), .A2(n13505), .ZN(n8894) );
  INV_X1 U11162 ( .A(n8894), .ZN(n8647) );
  NAND2_X1 U11163 ( .A1(n13153), .A2(n13505), .ZN(n8892) );
  NAND2_X1 U11164 ( .A1(n8648), .A2(n8892), .ZN(n13507) );
  NAND2_X1 U11165 ( .A1(n8649), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n8650) );
  NAND2_X1 U11166 ( .A1(n8651), .A2(n8650), .ZN(n11037) );
  OR2_X1 U11167 ( .A1(n8761), .A2(n11038), .ZN(n8652) );
  NAND2_X1 U11168 ( .A1(n8654), .A2(P3_REG3_REG_20__SCAN_IN), .ZN(n8655) );
  NAND2_X1 U11169 ( .A1(n8666), .A2(n8655), .ZN(n13509) );
  NAND2_X1 U11170 ( .A1(n13509), .A2(n8757), .ZN(n8658) );
  AOI22_X1 U11171 ( .A1(n6813), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n8764), .B2(
        P3_REG0_REG_20__SCAN_IN), .ZN(n8657) );
  NAND2_X1 U11172 ( .A1(n8736), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n8656) );
  NAND2_X1 U11173 ( .A1(n13274), .A2(n13519), .ZN(n8899) );
  NAND2_X1 U11174 ( .A1(n8898), .A2(n8899), .ZN(n13508) );
  OR2_X1 U11175 ( .A1(n8660), .A2(n8659), .ZN(n8661) );
  NAND2_X1 U11176 ( .A1(n8662), .A2(n8661), .ZN(n11136) );
  OR2_X1 U11177 ( .A1(n8761), .A2(n11137), .ZN(n8664) );
  NAND2_X1 U11178 ( .A1(n8666), .A2(P3_REG3_REG_21__SCAN_IN), .ZN(n8667) );
  NAND2_X1 U11179 ( .A1(n8677), .A2(n8667), .ZN(n13499) );
  NAND2_X1 U11180 ( .A1(n13499), .A2(n8757), .ZN(n8671) );
  AOI22_X1 U11181 ( .A1(n6813), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n8737), .B2(
        P3_REG0_REG_21__SCAN_IN), .ZN(n8670) );
  NAND2_X1 U11182 ( .A1(n8736), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n8669) );
  NAND2_X1 U11183 ( .A1(n13498), .A2(n13506), .ZN(n8904) );
  NAND2_X1 U11184 ( .A1(n13497), .A2(n8904), .ZN(n8672) );
  NAND2_X1 U11185 ( .A1(n8672), .A2(n8903), .ZN(n13485) );
  XNOR2_X1 U11186 ( .A(n8674), .B(n8673), .ZN(n11189) );
  NAND2_X1 U11187 ( .A1(n11189), .A2(n8760), .ZN(n8676) );
  OR2_X1 U11188 ( .A1(n8761), .A2(n6885), .ZN(n8675) );
  NAND2_X1 U11189 ( .A1(n8677), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n8678) );
  NAND2_X1 U11190 ( .A1(n8690), .A2(n8678), .ZN(n13486) );
  NAND2_X1 U11191 ( .A1(n13486), .A2(n8757), .ZN(n8684) );
  INV_X1 U11192 ( .A(P3_REG2_REG_22__SCAN_IN), .ZN(n8681) );
  NAND2_X1 U11193 ( .A1(n8736), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n8680) );
  NAND2_X1 U11194 ( .A1(n8764), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n8679) );
  OAI211_X1 U11195 ( .C1(n8767), .C2(n8681), .A(n8680), .B(n8679), .ZN(n8682)
         );
  INV_X1 U11196 ( .A(n8682), .ZN(n8683) );
  NAND2_X1 U11197 ( .A1(n13288), .A2(n13197), .ZN(n8908) );
  NAND2_X1 U11198 ( .A1(n13485), .A2(n8908), .ZN(n8685) );
  XNOR2_X1 U11199 ( .A(n8687), .B(n8686), .ZN(n11444) );
  NAND2_X1 U11200 ( .A1(n11444), .A2(n8760), .ZN(n8689) );
  OR2_X1 U11201 ( .A1(n8761), .A2(n11447), .ZN(n8688) );
  NAND2_X1 U11202 ( .A1(n8690), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n8691) );
  NAND2_X1 U11203 ( .A1(n8701), .A2(n8691), .ZN(n13475) );
  NAND2_X1 U11204 ( .A1(n13475), .A2(n8757), .ZN(n8697) );
  INV_X1 U11205 ( .A(P3_REG2_REG_23__SCAN_IN), .ZN(n8694) );
  NAND2_X1 U11206 ( .A1(n8737), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n8693) );
  NAND2_X1 U11207 ( .A1(n8736), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n8692) );
  OAI211_X1 U11208 ( .C1(n8694), .C2(n8767), .A(n8693), .B(n8692), .ZN(n8695)
         );
  INV_X1 U11209 ( .A(n8695), .ZN(n8696) );
  XNOR2_X1 U11210 ( .A(n13470), .B(n13483), .ZN(n13466) );
  INV_X1 U11211 ( .A(n13466), .ZN(n13471) );
  INV_X1 U11212 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n12747) );
  XNOR2_X1 U11213 ( .A(n8698), .B(n12747), .ZN(n12889) );
  NAND2_X1 U11214 ( .A1(n12889), .A2(n8760), .ZN(n8700) );
  OR2_X1 U11215 ( .A1(n8761), .A2(n12890), .ZN(n8699) );
  NAND2_X1 U11216 ( .A1(n8701), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n8702) );
  NAND2_X1 U11217 ( .A1(n8712), .A2(n8702), .ZN(n13461) );
  INV_X1 U11218 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n8705) );
  NAND2_X1 U11219 ( .A1(n8752), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n8704) );
  NAND2_X1 U11220 ( .A1(n8736), .A2(P3_REG1_REG_24__SCAN_IN), .ZN(n8703) );
  OAI211_X1 U11221 ( .C1(n8767), .C2(n8705), .A(n8704), .B(n8703), .ZN(n8706)
         );
  NAND2_X1 U11222 ( .A1(n13272), .A2(n13265), .ZN(n8798) );
  OR2_X1 U11223 ( .A1(n13272), .A2(n13265), .ZN(n8707) );
  NOR2_X1 U11224 ( .A1(n13470), .A2(n13483), .ZN(n13455) );
  XNOR2_X1 U11225 ( .A(n12327), .B(P2_DATAO_REG_25__SCAN_IN), .ZN(n8708) );
  XNOR2_X1 U11226 ( .A(n8709), .B(n8708), .ZN(n12031) );
  NAND2_X1 U11227 ( .A1(n12031), .A2(n8760), .ZN(n8711) );
  OR2_X1 U11228 ( .A1(n8761), .A2(n12032), .ZN(n8710) );
  NAND2_X1 U11229 ( .A1(n8712), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U11230 ( .A1(n8722), .A2(n8713), .ZN(n13449) );
  INV_X1 U11231 ( .A(P3_REG2_REG_25__SCAN_IN), .ZN(n8716) );
  NAND2_X1 U11232 ( .A1(n8752), .A2(P3_REG0_REG_25__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U11233 ( .A1(n8736), .A2(P3_REG1_REG_25__SCAN_IN), .ZN(n8714) );
  OAI211_X1 U11234 ( .C1(n8716), .C2(n8767), .A(n8715), .B(n8714), .ZN(n8717)
         );
  AOI21_X1 U11235 ( .B1(n13449), .B2(n8757), .A(n8717), .ZN(n13268) );
  OR2_X1 U11236 ( .A1(n13240), .A2(n13268), .ZN(n8796) );
  NAND2_X1 U11237 ( .A1(n13240), .A2(n13268), .ZN(n8797) );
  NAND2_X1 U11238 ( .A1(n8796), .A2(n8797), .ZN(n13447) );
  XNOR2_X1 U11239 ( .A(n12383), .B(P2_DATAO_REG_26__SCAN_IN), .ZN(n8718) );
  XNOR2_X1 U11240 ( .A(n8719), .B(n8718), .ZN(n12137) );
  NAND2_X1 U11241 ( .A1(n12137), .A2(n8760), .ZN(n8721) );
  OR2_X1 U11242 ( .A1(n8761), .A2(n12139), .ZN(n8720) );
  NAND2_X1 U11243 ( .A1(n8722), .A2(P3_REG3_REG_26__SCAN_IN), .ZN(n8723) );
  NAND2_X1 U11244 ( .A1(n8734), .A2(n8723), .ZN(n13437) );
  NAND2_X1 U11245 ( .A1(n13437), .A2(n8757), .ZN(n8729) );
  INV_X1 U11246 ( .A(P3_REG2_REG_26__SCAN_IN), .ZN(n8726) );
  NAND2_X1 U11247 ( .A1(n8736), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n8725) );
  NAND2_X1 U11248 ( .A1(n8764), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n8724) );
  OAI211_X1 U11249 ( .C1(n8767), .C2(n8726), .A(n8725), .B(n8724), .ZN(n8727)
         );
  INV_X1 U11250 ( .A(n8727), .ZN(n8728) );
  NAND2_X1 U11251 ( .A1(n13306), .A2(n13419), .ZN(n13422) );
  XNOR2_X1 U11252 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .ZN(n8730) );
  XNOR2_X1 U11253 ( .A(n8731), .B(n8730), .ZN(n12214) );
  NAND2_X1 U11254 ( .A1(n12214), .A2(n8760), .ZN(n8733) );
  OR2_X1 U11255 ( .A1(n8761), .A2(n12215), .ZN(n8732) );
  NAND2_X1 U11256 ( .A1(n8734), .A2(P3_REG3_REG_27__SCAN_IN), .ZN(n8735) );
  NAND2_X1 U11257 ( .A1(n8749), .A2(n8735), .ZN(n13426) );
  NAND2_X1 U11258 ( .A1(n13426), .A2(n8757), .ZN(n8743) );
  INV_X1 U11259 ( .A(P3_REG2_REG_27__SCAN_IN), .ZN(n8740) );
  NAND2_X1 U11260 ( .A1(n8736), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n8739) );
  NAND2_X1 U11261 ( .A1(n8737), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n8738) );
  OAI211_X1 U11262 ( .C1(n8767), .C2(n8740), .A(n8739), .B(n8738), .ZN(n8741)
         );
  INV_X1 U11263 ( .A(n8741), .ZN(n8742) );
  NAND2_X1 U11264 ( .A1(n13180), .A2(n13218), .ZN(n9040) );
  OR2_X1 U11265 ( .A1(n13180), .A2(n13218), .ZN(n8744) );
  XNOR2_X1 U11266 ( .A(n14200), .B(P2_DATAO_REG_28__SCAN_IN), .ZN(n8745) );
  XNOR2_X1 U11267 ( .A(n8746), .B(n8745), .ZN(n12945) );
  NAND2_X1 U11268 ( .A1(n12945), .A2(n8760), .ZN(n8748) );
  OR2_X1 U11269 ( .A1(n8761), .A2(n12946), .ZN(n8747) );
  NAND2_X2 U11270 ( .A1(n8748), .A2(n8747), .ZN(n13222) );
  NAND2_X1 U11271 ( .A1(n8749), .A2(P3_REG3_REG_28__SCAN_IN), .ZN(n8750) );
  NAND2_X1 U11272 ( .A1(n8751), .A2(n8750), .ZN(n13408) );
  INV_X1 U11273 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n8755) );
  NAND2_X1 U11274 ( .A1(n8736), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n8754) );
  NAND2_X1 U11275 ( .A1(n8752), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n8753) );
  OAI211_X1 U11276 ( .C1(n8767), .C2(n8755), .A(n8754), .B(n8753), .ZN(n8756)
         );
  AOI21_X1 U11277 ( .B1(n13408), .B2(n8757), .A(n8756), .ZN(n13420) );
  NAND2_X1 U11278 ( .A1(n13222), .A2(n13420), .ZN(n8777) );
  NAND2_X1 U11279 ( .A1(n8777), .A2(n9040), .ZN(n8924) );
  NAND2_X1 U11280 ( .A1(n13684), .A2(n8760), .ZN(n8763) );
  OR2_X1 U11281 ( .A1(n8761), .A2(n13689), .ZN(n8762) );
  INV_X1 U11282 ( .A(P3_REG2_REG_29__SCAN_IN), .ZN(n13124) );
  NAND2_X1 U11283 ( .A1(n8736), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8766) );
  NAND2_X1 U11284 ( .A1(n8764), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8765) );
  OAI211_X1 U11285 ( .C1(n8767), .C2(n13124), .A(n8766), .B(n8765), .ZN(n8768)
         );
  INV_X1 U11286 ( .A(n8768), .ZN(n8769) );
  NAND2_X1 U11287 ( .A1(n8773), .A2(n11375), .ZN(n8771) );
  NAND2_X1 U11288 ( .A1(n8772), .A2(n8771), .ZN(n8795) );
  NAND2_X1 U11289 ( .A1(n13128), .A2(n13219), .ZN(n8928) );
  OAI21_X1 U11290 ( .B1(n13629), .B2(n7221), .A(n8928), .ZN(n8774) );
  NAND2_X1 U11291 ( .A1(n8775), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n8776) );
  INV_X1 U11292 ( .A(n11039), .ZN(n9012) );
  NAND2_X1 U11293 ( .A1(n10704), .A2(n9012), .ZN(n8985) );
  INV_X1 U11294 ( .A(n13216), .ZN(n8926) );
  INV_X1 U11295 ( .A(n13435), .ZN(n13431) );
  XNOR2_X1 U11296 ( .A(n13153), .B(n13505), .ZN(n13521) );
  NAND2_X1 U11297 ( .A1(n8867), .A2(n8866), .ZN(n12205) );
  NOR2_X1 U11298 ( .A1(n11303), .A2(n11742), .ZN(n8779) );
  INV_X1 U11299 ( .A(n10772), .ZN(n8778) );
  NAND4_X1 U11300 ( .A1(n8779), .A2(n11753), .A3(n11765), .A4(n8778), .ZN(
        n8783) );
  NAND2_X1 U11301 ( .A1(n13330), .A2(n10680), .ZN(n8801) );
  INV_X1 U11302 ( .A(n8801), .ZN(n8780) );
  NOR2_X1 U11303 ( .A1(n10770), .A2(n8780), .ZN(n10565) );
  NAND4_X1 U11304 ( .A1(n10565), .A2(n8781), .A3(n11544), .A4(n11778), .ZN(
        n8782) );
  NOR2_X1 U11305 ( .A1(n8783), .A2(n8782), .ZN(n8784) );
  NAND2_X1 U11306 ( .A1(n8850), .A2(n8842), .ZN(n11824) );
  INV_X1 U11307 ( .A(n11824), .ZN(n11821) );
  XNOR2_X1 U11308 ( .A(n13325), .B(n11531), .ZN(n11525) );
  NAND4_X1 U11309 ( .A1(n8784), .A2(n6740), .A3(n11821), .A4(n11525), .ZN(
        n8785) );
  INV_X1 U11310 ( .A(n12052), .ZN(n12045) );
  NAND2_X1 U11311 ( .A1(n8860), .A2(n8861), .ZN(n12129) );
  OR3_X1 U11312 ( .A1(n8785), .A2(n12045), .A3(n12129), .ZN(n8786) );
  NOR2_X1 U11313 ( .A1(n12205), .A2(n8786), .ZN(n8787) );
  NAND4_X1 U11314 ( .A1(n13556), .A2(n8863), .A3(n12370), .A4(n8787), .ZN(
        n8788) );
  OR4_X1 U11315 ( .A1(n13508), .A2(n13521), .A3(n13546), .A4(n8788), .ZN(n8789) );
  NAND2_X1 U11316 ( .A1(n8903), .A2(n8904), .ZN(n13496) );
  AND2_X2 U11317 ( .A1(n8907), .A2(n8908), .ZN(n13480) );
  INV_X1 U11318 ( .A(n13480), .ZN(n13484) );
  OR4_X1 U11319 ( .A1(n13466), .A2(n8789), .A3(n13496), .A4(n13484), .ZN(n8790) );
  OR3_X1 U11320 ( .A1(n13447), .A2(n13454), .A3(n8790), .ZN(n8791) );
  NOR2_X1 U11321 ( .A1(n13431), .A2(n8791), .ZN(n8792) );
  NAND4_X1 U11322 ( .A1(n6756), .A2(n13417), .A3(n8926), .A4(n8792), .ZN(n8793) );
  INV_X1 U11323 ( .A(n10702), .ZN(n8937) );
  NAND2_X1 U11324 ( .A1(n9014), .A2(n11039), .ZN(n11314) );
  INV_X1 U11325 ( .A(n11314), .ZN(n11310) );
  INV_X1 U11326 ( .A(n10706), .ZN(n8939) );
  INV_X1 U11327 ( .A(n8795), .ZN(n8935) );
  MUX2_X1 U11328 ( .A(n8797), .B(n8796), .S(n9015), .Z(n8915) );
  XNOR2_X1 U11329 ( .A(n8798), .B(n9026), .ZN(n8799) );
  AND2_X1 U11330 ( .A1(n8800), .A2(n8799), .ZN(n8914) );
  OAI21_X1 U11331 ( .B1(n10770), .B2(n10704), .A(n8801), .ZN(n8803) );
  AND2_X1 U11332 ( .A1(n8804), .A2(n8801), .ZN(n8802) );
  MUX2_X1 U11333 ( .A(n8803), .B(n8802), .S(n9015), .Z(n8808) );
  MUX2_X1 U11334 ( .A(n8804), .B(n10708), .S(n9015), .Z(n8805) );
  NAND2_X1 U11335 ( .A1(n8806), .A2(n8805), .ZN(n8807) );
  AOI21_X1 U11336 ( .B1(n8808), .B2(n10708), .A(n8807), .ZN(n8811) );
  AOI21_X1 U11337 ( .B1(n8817), .B2(n8809), .A(n9026), .ZN(n8810) );
  OAI21_X1 U11338 ( .B1(n8811), .B2(n8810), .A(n8813), .ZN(n8816) );
  NAND2_X1 U11339 ( .A1(n8813), .A2(n8812), .ZN(n8814) );
  NAND2_X1 U11340 ( .A1(n8814), .A2(n9026), .ZN(n8815) );
  NAND2_X1 U11341 ( .A1(n8816), .A2(n8815), .ZN(n8820) );
  NOR2_X1 U11342 ( .A1(n8817), .A2(n9015), .ZN(n8818) );
  NOR2_X1 U11343 ( .A1(n11742), .A2(n8818), .ZN(n8819) );
  NAND2_X1 U11344 ( .A1(n8820), .A2(n8819), .ZN(n8825) );
  NAND3_X1 U11345 ( .A1(n8825), .A2(n11544), .A3(n8821), .ZN(n8823) );
  NAND3_X1 U11346 ( .A1(n8823), .A2(n8822), .A3(n11937), .ZN(n8829) );
  NAND3_X1 U11347 ( .A1(n8825), .A2(n11544), .A3(n8824), .ZN(n8827) );
  INV_X1 U11348 ( .A(n11937), .ZN(n8826) );
  AOI21_X1 U11349 ( .B1(n8827), .B2(n11935), .A(n8826), .ZN(n8828) );
  MUX2_X1 U11350 ( .A(n8829), .B(n8828), .S(n9015), .Z(n8833) );
  NOR2_X1 U11351 ( .A1(n8830), .A2(n9015), .ZN(n8831) );
  NOR2_X1 U11352 ( .A1(n8831), .A2(n11940), .ZN(n8832) );
  NAND2_X1 U11353 ( .A1(n8833), .A2(n8832), .ZN(n8838) );
  MUX2_X1 U11354 ( .A(n8835), .B(n8834), .S(n9015), .Z(n8836) );
  AND2_X1 U11355 ( .A1(n8836), .A2(n11778), .ZN(n8837) );
  NAND2_X1 U11356 ( .A1(n8838), .A2(n8837), .ZN(n8849) );
  NAND3_X1 U11357 ( .A1(n8849), .A2(n11525), .A3(n8839), .ZN(n8841) );
  AOI21_X1 U11358 ( .B1(n8841), .B2(n8840), .A(n11824), .ZN(n8845) );
  NAND2_X1 U11359 ( .A1(n12052), .A2(n8842), .ZN(n8844) );
  OAI211_X1 U11360 ( .C1(n8845), .C2(n8844), .A(n8855), .B(n8843), .ZN(n8854)
         );
  AND2_X1 U11361 ( .A1(n11525), .A2(n8846), .ZN(n8848) );
  AOI21_X1 U11362 ( .B1(n8849), .B2(n8848), .A(n8847), .ZN(n8851) );
  OAI211_X1 U11363 ( .C1(n8851), .C2(n11824), .A(n12052), .B(n8850), .ZN(n8852) );
  OAI211_X1 U11364 ( .C1(n12390), .C2(n12054), .A(n8852), .B(n8856), .ZN(n8853) );
  MUX2_X1 U11365 ( .A(n8854), .B(n8853), .S(n9015), .Z(n8859) );
  INV_X1 U11366 ( .A(n12129), .ZN(n8858) );
  MUX2_X1 U11367 ( .A(n8856), .B(n8855), .S(n9015), .Z(n8857) );
  NAND3_X1 U11368 ( .A1(n8859), .A2(n8858), .A3(n8857), .ZN(n8864) );
  INV_X1 U11369 ( .A(n12205), .ZN(n12203) );
  MUX2_X1 U11370 ( .A(n8861), .B(n8860), .S(n9026), .Z(n8862) );
  NAND4_X1 U11371 ( .A1(n8864), .A2(n12203), .A3(n8863), .A4(n8862), .ZN(n8872) );
  OAI211_X1 U11372 ( .C1(n8866), .C2(n12329), .A(n8875), .B(n8865), .ZN(n8869)
         );
  NOR2_X1 U11373 ( .A1(n12329), .A2(n8867), .ZN(n8868) );
  MUX2_X1 U11374 ( .A(n8869), .B(n8868), .S(n9015), .Z(n8870) );
  INV_X1 U11375 ( .A(n8870), .ZN(n8871) );
  AOI21_X1 U11376 ( .B1(n8872), .B2(n8871), .A(n7431), .ZN(n8877) );
  AOI21_X1 U11377 ( .B1(n8874), .B2(n8873), .A(n9026), .ZN(n8876) );
  OAI22_X1 U11378 ( .A1(n8877), .A2(n8876), .B1(n9026), .B2(n8875), .ZN(n8878)
         );
  NAND3_X1 U11379 ( .A1(n8878), .A2(n13528), .A3(n13556), .ZN(n8891) );
  INV_X1 U11380 ( .A(n8879), .ZN(n8880) );
  NAND2_X1 U11381 ( .A1(n13528), .A2(n8880), .ZN(n8881) );
  AND3_X1 U11382 ( .A1(n8881), .A2(n8892), .A3(n8884), .ZN(n8889) );
  INV_X1 U11383 ( .A(n8882), .ZN(n8883) );
  NAND2_X1 U11384 ( .A1(n8884), .A2(n8883), .ZN(n8886) );
  NAND2_X1 U11385 ( .A1(n8886), .A2(n8885), .ZN(n8887) );
  NOR2_X1 U11386 ( .A1(n8894), .A2(n8887), .ZN(n8888) );
  MUX2_X1 U11387 ( .A(n8889), .B(n8888), .S(n9015), .Z(n8890) );
  NAND2_X1 U11388 ( .A1(n8891), .A2(n8890), .ZN(n8897) );
  INV_X1 U11389 ( .A(n8892), .ZN(n8893) );
  MUX2_X1 U11390 ( .A(n8894), .B(n8893), .S(n9015), .Z(n8895) );
  NOR2_X1 U11391 ( .A1(n13508), .A2(n8895), .ZN(n8896) );
  NAND2_X1 U11392 ( .A1(n8897), .A2(n8896), .ZN(n8902) );
  INV_X1 U11393 ( .A(n13496), .ZN(n8901) );
  MUX2_X1 U11394 ( .A(n8899), .B(n8898), .S(n9015), .Z(n8900) );
  NAND3_X1 U11395 ( .A1(n8902), .A2(n8901), .A3(n8900), .ZN(n8906) );
  MUX2_X1 U11396 ( .A(n8904), .B(n8903), .S(n9026), .Z(n8905) );
  NAND3_X1 U11397 ( .A1(n8906), .A2(n13480), .A3(n8905), .ZN(n8910) );
  MUX2_X1 U11398 ( .A(n8908), .B(n8907), .S(n9015), .Z(n8909) );
  NAND3_X1 U11399 ( .A1(n8910), .A2(n13471), .A3(n8909), .ZN(n8912) );
  NAND3_X1 U11400 ( .A1(n13470), .A2(n13483), .A3(n9015), .ZN(n8911) );
  NAND2_X1 U11401 ( .A1(n8912), .A2(n8911), .ZN(n8913) );
  MUX2_X1 U11402 ( .A(n13422), .B(n8916), .S(n9026), .Z(n8917) );
  NAND2_X1 U11403 ( .A1(n8918), .A2(n8917), .ZN(n8919) );
  NAND2_X1 U11404 ( .A1(n13417), .A2(n8919), .ZN(n8921) );
  OR3_X1 U11405 ( .A1(n13180), .A2(n9015), .A3(n13218), .ZN(n8920) );
  OAI211_X1 U11406 ( .C1(n9026), .C2(n8924), .A(n8923), .B(n8922), .ZN(n8929)
         );
  NAND3_X1 U11407 ( .A1(n8926), .A2(n9015), .A3(n8925), .ZN(n8927) );
  NAND3_X1 U11408 ( .A1(n8929), .A2(n8928), .A3(n8927), .ZN(n8933) );
  INV_X1 U11409 ( .A(n8930), .ZN(n8932) );
  INV_X1 U11410 ( .A(n11445), .ZN(n8938) );
  NAND2_X1 U11411 ( .A1(n10562), .A2(n8939), .ZN(n10551) );
  NAND3_X1 U11412 ( .A1(n8986), .A2(n9015), .A3(n6879), .ZN(n13518) );
  NOR3_X1 U11413 ( .A1(n10551), .A2(n6812), .A3(n13518), .ZN(n8941) );
  OAI21_X1 U11414 ( .B1(n11445), .B2(n11190), .A(P3_B_REG_SCAN_IN), .ZN(n8940)
         );
  OR2_X1 U11415 ( .A1(n8941), .A2(n8940), .ZN(n8942) );
  NAND2_X1 U11416 ( .A1(n8943), .A2(n8942), .ZN(P3_U3296) );
  NAND2_X1 U11417 ( .A1(n11190), .A2(n11039), .ZN(n8944) );
  AOI21_X1 U11418 ( .B1(n9014), .B2(n8944), .A(n10704), .ZN(n8947) );
  INV_X1 U11419 ( .A(n11190), .ZN(n9013) );
  NAND2_X1 U11420 ( .A1(n11313), .A2(n11039), .ZN(n8945) );
  AND2_X1 U11421 ( .A1(n9013), .A2(n8945), .ZN(n8946) );
  OR2_X1 U11422 ( .A1(n8947), .A2(n8946), .ZN(n10555) );
  NOR2_X1 U11423 ( .A1(n10706), .A2(n15561), .ZN(n8948) );
  NAND2_X1 U11424 ( .A1(n10555), .A2(n8948), .ZN(n8950) );
  AND2_X1 U11425 ( .A1(n11190), .A2(n9012), .ZN(n8949) );
  NAND2_X1 U11426 ( .A1(n7457), .A2(n8949), .ZN(n9011) );
  AND2_X1 U11427 ( .A1(n8950), .A2(n9011), .ZN(n15557) );
  OR2_X1 U11428 ( .A1(n11314), .A2(n11190), .ZN(n15583) );
  INV_X1 U11429 ( .A(n13506), .ZN(n13284) );
  NAND2_X1 U11430 ( .A1(n8952), .A2(n8953), .ZN(n11751) );
  INV_X1 U11431 ( .A(n11751), .ZN(n8954) );
  NAND2_X1 U11432 ( .A1(n13330), .A2(n11011), .ZN(n10771) );
  NAND2_X1 U11433 ( .A1(n10772), .A2(n10771), .ZN(n8957) );
  NAND2_X1 U11434 ( .A1(n11305), .A2(n8956), .ZN(n10709) );
  NAND2_X1 U11435 ( .A1(n8957), .A2(n10709), .ZN(n11302) );
  NAND2_X1 U11436 ( .A1(n11302), .A2(n11303), .ZN(n11752) );
  NAND2_X1 U11437 ( .A1(n8958), .A2(n11752), .ZN(n11756) );
  NAND2_X1 U11438 ( .A1(n11091), .A2(n11759), .ZN(n11537) );
  NAND2_X1 U11439 ( .A1(n11543), .A2(n15545), .ZN(n11538) );
  INV_X1 U11440 ( .A(n11538), .ZN(n8959) );
  AND2_X1 U11441 ( .A1(n11537), .A2(n8961), .ZN(n8960) );
  NAND2_X1 U11442 ( .A1(n11767), .A2(n15550), .ZN(n8962) );
  AND2_X1 U11443 ( .A1(n8962), .A2(n11539), .ZN(n8963) );
  NAND2_X1 U11444 ( .A1(n13326), .A2(n15560), .ZN(n8965) );
  NAND2_X1 U11445 ( .A1(n11770), .A2(n8965), .ZN(n11941) );
  NAND2_X1 U11446 ( .A1(n11714), .A2(n8966), .ZN(n8967) );
  NAND2_X1 U11447 ( .A1(n13325), .A2(n11531), .ZN(n8968) );
  NAND2_X1 U11448 ( .A1(n11527), .A2(n8968), .ZN(n11825) );
  NAND2_X1 U11449 ( .A1(n11825), .A2(n11824), .ZN(n11823) );
  NAND2_X1 U11450 ( .A1(n13324), .A2(n15378), .ZN(n8969) );
  NAND2_X1 U11451 ( .A1(n11823), .A2(n8969), .ZN(n12046) );
  NAND2_X1 U11452 ( .A1(n12390), .A2(n14953), .ZN(n8970) );
  NAND2_X1 U11453 ( .A1(n12398), .A2(n12054), .ZN(n8971) );
  INV_X1 U11454 ( .A(n12388), .ZN(n13323) );
  NAND2_X1 U11455 ( .A1(n12130), .A2(n12129), .ZN(n8973) );
  INV_X1 U11456 ( .A(n13186), .ZN(n12433) );
  OR2_X1 U11457 ( .A1(n14943), .A2(n12433), .ZN(n8972) );
  NAND2_X1 U11458 ( .A1(n8973), .A2(n8972), .ZN(n12206) );
  NAND2_X1 U11459 ( .A1(n12206), .A2(n12205), .ZN(n8975) );
  INV_X1 U11460 ( .A(n13312), .ZN(n13137) );
  OR2_X1 U11461 ( .A1(n14938), .A2(n13137), .ZN(n8974) );
  NAND2_X1 U11462 ( .A1(n8975), .A2(n8974), .ZN(n12330) );
  NAND2_X1 U11463 ( .A1(n12330), .A2(n12329), .ZN(n8977) );
  INV_X1 U11464 ( .A(n13140), .ZN(n13188) );
  OR2_X1 U11465 ( .A1(n14933), .A2(n13188), .ZN(n8976) );
  INV_X1 U11466 ( .A(n13532), .ZN(n13294) );
  OR2_X1 U11467 ( .A1(n13670), .A2(n13294), .ZN(n8979) );
  NAND2_X1 U11468 ( .A1(n13551), .A2(n8979), .ZN(n13529) );
  INV_X1 U11469 ( .A(n13517), .ZN(n13150) );
  NOR2_X1 U11470 ( .A1(n13153), .A2(n13534), .ZN(n8980) );
  NAND2_X1 U11471 ( .A1(n13288), .A2(n13494), .ZN(n8981) );
  INV_X1 U11472 ( .A(n13288), .ZN(n13653) );
  INV_X1 U11473 ( .A(n13483), .ZN(n13322) );
  INV_X1 U11474 ( .A(n13272), .ZN(n13645) );
  NOR2_X1 U11475 ( .A1(n13645), .A2(n13265), .ZN(n13442) );
  NAND2_X1 U11476 ( .A1(n9043), .A2(n7635), .ZN(n8984) );
  XNOR2_X1 U11477 ( .A(n8984), .B(n6756), .ZN(n8990) );
  NAND2_X1 U11478 ( .A1(n9014), .A2(n11190), .ZN(n9027) );
  NAND2_X1 U11479 ( .A1(n8986), .A2(n6879), .ZN(n8987) );
  NOR2_X1 U11480 ( .A1(n6812), .A2(n8036), .ZN(n8988) );
  OR2_X1 U11481 ( .A1(n13520), .A2(n8988), .ZN(n13401) );
  OAI22_X1 U11482 ( .A1(n13420), .A2(n13518), .B1(n11375), .B2(n13401), .ZN(
        n8989) );
  NAND2_X1 U11483 ( .A1(n8991), .A2(n12033), .ZN(n8992) );
  INV_X1 U11484 ( .A(n8993), .ZN(n12138) );
  NAND2_X1 U11485 ( .A1(n12892), .A2(n12138), .ZN(n8994) );
  OR2_X1 U11486 ( .A1(n10242), .A2(P3_D_REG_1__SCAN_IN), .ZN(n8997) );
  NAND2_X1 U11487 ( .A1(n12033), .A2(n12138), .ZN(n8996) );
  XNOR2_X1 U11488 ( .A(n10703), .B(n11006), .ZN(n9010) );
  NOR2_X1 U11489 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n9001) );
  NOR4_X1 U11490 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n9000) );
  NOR4_X1 U11491 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8999) );
  NOR4_X1 U11492 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8998) );
  NAND4_X1 U11493 ( .A1(n9001), .A2(n9000), .A3(n8999), .A4(n8998), .ZN(n9007)
         );
  NOR4_X1 U11494 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n9005) );
  NOR4_X1 U11495 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n9004) );
  NOR4_X1 U11496 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n9003) );
  NOR4_X1 U11497 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n9002) );
  NAND4_X1 U11498 ( .A1(n9005), .A2(n9004), .A3(n9003), .A4(n9002), .ZN(n9006)
         );
  NOR2_X1 U11499 ( .A1(n9007), .A2(n9006), .ZN(n9008) );
  OR2_X1 U11500 ( .A1(n10242), .A2(n9008), .ZN(n9028) );
  AND2_X1 U11501 ( .A1(n10562), .A2(n9028), .ZN(n9009) );
  NAND2_X1 U11502 ( .A1(n10706), .A2(n9015), .ZN(n11002) );
  NAND2_X1 U11503 ( .A1(n9011), .A2(n9026), .ZN(n11004) );
  AND2_X1 U11504 ( .A1(n11002), .A2(n11004), .ZN(n9019) );
  OAI22_X1 U11505 ( .A1(n9014), .A2(n9013), .B1(n9012), .B2(n15582), .ZN(n9016) );
  AOI21_X1 U11506 ( .B1(n9016), .B2(n10706), .A(n9015), .ZN(n9018) );
  INV_X1 U11507 ( .A(n11006), .ZN(n9017) );
  MUX2_X1 U11508 ( .A(n9019), .B(n9018), .S(n9017), .Z(n9020) );
  INV_X1 U11509 ( .A(n13128), .ZN(n9035) );
  INV_X1 U11510 ( .A(n13623), .ZN(n9021) );
  NAND2_X1 U11511 ( .A1(n13128), .A2(n9021), .ZN(n9024) );
  INV_X1 U11512 ( .A(n10703), .ZN(n10219) );
  NAND3_X1 U11513 ( .A1(n10219), .A2(n11006), .A3(n9028), .ZN(n10556) );
  OR2_X1 U11514 ( .A1(n10706), .A2(n9026), .ZN(n10543) );
  OR2_X1 U11515 ( .A1(n9027), .A2(n10702), .ZN(n10548) );
  AND2_X1 U11516 ( .A1(n10543), .A2(n10548), .ZN(n10557) );
  NAND2_X1 U11517 ( .A1(n10703), .A2(n9028), .ZN(n9029) );
  OR2_X1 U11518 ( .A1(n11006), .A2(n9029), .ZN(n10559) );
  INV_X1 U11519 ( .A(n10555), .ZN(n9030) );
  OAI22_X1 U11520 ( .A1(n10556), .A2(n10557), .B1(n10559), .B2(n9030), .ZN(
        n9031) );
  OR2_X1 U11521 ( .A1(n15591), .A2(n9033), .ZN(n9034) );
  INV_X1 U11522 ( .A(n9036), .ZN(n9037) );
  NAND2_X1 U11523 ( .A1(n9038), .A2(n9037), .ZN(P3_U3456) );
  INV_X1 U11524 ( .A(n9040), .ZN(n9041) );
  NOR2_X1 U11525 ( .A1(n9039), .A2(n9041), .ZN(n9042) );
  XNOR2_X1 U11526 ( .A(n9042), .B(n13216), .ZN(n13412) );
  AOI21_X1 U11527 ( .B1(n13412), .B2(n14957), .A(n13407), .ZN(n9052) );
  OR2_X1 U11528 ( .A1(n9052), .A2(n15589), .ZN(n9051) );
  INV_X1 U11529 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n9048) );
  INV_X1 U11530 ( .A(n9049), .ZN(n9050) );
  NAND2_X1 U11531 ( .A1(n9051), .A2(n9050), .ZN(P3_U3455) );
  INV_X1 U11532 ( .A(P3_REG1_REG_28__SCAN_IN), .ZN(n9053) );
  MUX2_X1 U11533 ( .A(n9053), .B(n9052), .S(n15607), .Z(n9054) );
  NAND2_X1 U11534 ( .A1(n9054), .A2(n7630), .ZN(P3_U3487) );
  NOR2_X1 U11535 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), 
        .ZN(n9057) );
  NAND4_X1 U11536 ( .A1(n9057), .A2(n9056), .A3(n9055), .A4(n9313), .ZN(n9410)
         );
  NAND3_X1 U11537 ( .A1(n9059), .A2(n9254), .A3(n9058), .ZN(n9060) );
  INV_X1 U11538 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n9164) );
  NOR2_X2 U11539 ( .A1(P2_IR_REG_1__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n9087) );
  AND2_X2 U11540 ( .A1(n9087), .A2(n9063), .ZN(n9109) );
  INV_X1 U11541 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n9067) );
  NAND3_X1 U11542 ( .A1(n9078), .A2(n9067), .A3(n9080), .ZN(n9068) );
  NAND2_X1 U11543 ( .A1(n9599), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n9076) );
  INV_X1 U11544 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n11472) );
  INV_X1 U11545 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9071) );
  INV_X1 U11546 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n10075) );
  NAND2_X1 U11547 ( .A1(n9079), .A2(n9067), .ZN(n9685) );
  XNOR2_X2 U11548 ( .A(n9081), .B(n9080), .ZN(n9668) );
  MUX2_X1 U11549 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9083), .S(
        P2_IR_REG_28__SCAN_IN), .Z(n9085) );
  NAND2_X1 U11550 ( .A1(n9085), .A2(n9084), .ZN(n10070) );
  NAND2_X1 U11551 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n9086) );
  MUX2_X1 U11552 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9086), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n9089) );
  INV_X1 U11553 ( .A(n9087), .ZN(n9088) );
  NAND2_X1 U11554 ( .A1(n9089), .A2(n9088), .ZN(n15185) );
  INV_X1 U11555 ( .A(n9091), .ZN(n9090) );
  NAND2_X1 U11556 ( .A1(n9092), .A2(SI_0_), .ZN(n9103) );
  XNOR2_X1 U11557 ( .A(n9104), .B(n9103), .ZN(n10615) );
  INV_X1 U11558 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n15189) );
  NAND2_X1 U11559 ( .A1(n9213), .A2(SI_0_), .ZN(n9094) );
  XNOR2_X1 U11560 ( .A(n9094), .B(n9093), .ZN(n14202) );
  INV_X1 U11561 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n11065) );
  OR2_X1 U11562 ( .A1(n9131), .A2(n11065), .ZN(n9101) );
  INV_X1 U11563 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10047) );
  OR2_X1 U11564 ( .A1(n6666), .A2(n10047), .ZN(n9099) );
  INV_X1 U11565 ( .A(n9763), .ZN(n10698) );
  NOR2_X1 U11566 ( .A1(n11474), .A2(n9763), .ZN(n11469) );
  NAND2_X1 U11567 ( .A1(n6826), .A2(n11469), .ZN(n11467) );
  INV_X1 U11568 ( .A(n13891), .ZN(n10903) );
  NAND2_X1 U11569 ( .A1(n10903), .A2(n10725), .ZN(n9102) );
  NAND2_X1 U11570 ( .A1(n11467), .A2(n9102), .ZN(n15264) );
  OAI21_X1 U11571 ( .B1(n9147), .B2(SI_2_), .A(n9122), .ZN(n9121) );
  NOR2_X1 U11572 ( .A1(n9087), .A2(n9658), .ZN(n9107) );
  MUX2_X1 U11573 ( .A(n9658), .B(n9107), .S(P2_IR_REG_2__SCAN_IN), .Z(n9108)
         );
  INV_X1 U11574 ( .A(n9108), .ZN(n9111) );
  INV_X1 U11575 ( .A(n9109), .ZN(n9110) );
  NAND2_X1 U11576 ( .A1(n9111), .A2(n9110), .ZN(n10389) );
  OR2_X1 U11577 ( .A1(n9096), .A2(n10389), .ZN(n9113) );
  OR2_X1 U11578 ( .A1(n9948), .A2(n10183), .ZN(n9112) );
  NAND2_X1 U11579 ( .A1(n9599), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n9118) );
  INV_X1 U11580 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10377) );
  OR2_X1 U11581 ( .A1(n9131), .A2(n10377), .ZN(n9117) );
  INV_X1 U11582 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10079) );
  INV_X1 U11583 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n9114) );
  OR2_X1 U11584 ( .A1(n9420), .A2(n9114), .ZN(n9115) );
  AND4_X2 U11585 ( .A1(n9118), .A2(n9117), .A3(n9116), .A4(n9115), .ZN(n9722)
         );
  NAND2_X1 U11586 ( .A1(n15264), .A2(n15265), .ZN(n9120) );
  OR2_X1 U11587 ( .A1(n15306), .A2(n13890), .ZN(n9119) );
  NAND2_X1 U11588 ( .A1(n9120), .A2(n9119), .ZN(n11291) );
  OR2_X1 U11589 ( .A1(n9121), .A2(n9142), .ZN(n9123) );
  NAND2_X1 U11590 ( .A1(n9123), .A2(n9122), .ZN(n9125) );
  NAND2_X1 U11591 ( .A1(n9124), .A2(SI_3_), .ZN(n9148) );
  OAI21_X1 U11592 ( .B1(n9124), .B2(SI_3_), .A(n9148), .ZN(n9145) );
  INV_X2 U11593 ( .A(n9948), .ZN(n9456) );
  NOR2_X1 U11594 ( .A1(n9109), .A2(n9658), .ZN(n9126) );
  MUX2_X1 U11595 ( .A(n9658), .B(n9126), .S(P2_IR_REG_3__SCAN_IN), .Z(n9128)
         );
  AND2_X1 U11596 ( .A1(n9109), .A2(n9127), .ZN(n9139) );
  NOR2_X1 U11597 ( .A1(n9128), .A2(n9139), .ZN(n10184) );
  INV_X2 U11598 ( .A(n9131), .ZN(n9341) );
  OR2_X1 U11599 ( .A1(n9616), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9136) );
  INV_X2 U11600 ( .A(n6666), .ZN(n9923) );
  NAND2_X1 U11601 ( .A1(n9923), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9135) );
  INV_X1 U11602 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n10074) );
  OR2_X1 U11603 ( .A1(n9928), .A2(n10074), .ZN(n9134) );
  INV_X1 U11604 ( .A(n9599), .ZN(n9343) );
  INV_X1 U11605 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n9132) );
  OR2_X1 U11606 ( .A1(n9343), .A2(n9132), .ZN(n9133) );
  NAND4_X2 U11607 ( .A1(n9136), .A2(n9135), .A3(n9134), .A4(n9133), .ZN(n13889) );
  NAND2_X1 U11608 ( .A1(n11291), .A2(n11290), .ZN(n9138) );
  INV_X1 U11609 ( .A(n13889), .ZN(n10902) );
  NAND2_X1 U11610 ( .A1(n15314), .A2(n10902), .ZN(n9137) );
  INV_X1 U11611 ( .A(n9139), .ZN(n9163) );
  NAND2_X1 U11612 ( .A1(n9163), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9141) );
  INV_X1 U11613 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n9140) );
  XNOR2_X1 U11614 ( .A(n9141), .B(n9140), .ZN(n10314) );
  INV_X1 U11615 ( .A(SI_2_), .ZN(n10150) );
  NOR2_X1 U11616 ( .A1(n9143), .A2(SI_2_), .ZN(n9144) );
  MUX2_X1 U11617 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n6670), .Z(n9149) );
  NAND2_X1 U11618 ( .A1(n9149), .A2(SI_4_), .ZN(n9185) );
  OAI21_X1 U11619 ( .B1(n9149), .B2(SI_4_), .A(n9185), .ZN(n9159) );
  XNOR2_X1 U11620 ( .A(n9161), .B(n9159), .ZN(n10118) );
  OR2_X1 U11621 ( .A1(n9948), .A2(n10182), .ZN(n9151) );
  OAI211_X1 U11622 ( .C1(n9096), .C2(n10314), .A(n9152), .B(n9151), .ZN(n11116) );
  NAND2_X1 U11623 ( .A1(n9924), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9156) );
  INV_X1 U11624 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10083) );
  OR2_X1 U11625 ( .A1(n9928), .A2(n10083), .ZN(n9155) );
  INV_X1 U11626 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n11124) );
  OR2_X1 U11627 ( .A1(n6666), .A2(n11124), .ZN(n9154) );
  OAI21_X1 U11628 ( .B1(P2_REG3_REG_4__SCAN_IN), .B2(P2_REG3_REG_3__SCAN_IN), 
        .A(n9173), .ZN(n11117) );
  OR2_X1 U11629 ( .A1(n9616), .A2(n11117), .ZN(n9153) );
  NAND4_X1 U11630 ( .A1(n9156), .A2(n9155), .A3(n9154), .A4(n9153), .ZN(n13888) );
  XNOR2_X1 U11631 ( .A(n11116), .B(n9786), .ZN(n9976) );
  INV_X1 U11632 ( .A(n9976), .ZN(n11119) );
  NAND2_X1 U11633 ( .A1(n11120), .A2(n11119), .ZN(n9158) );
  NAND2_X1 U11634 ( .A1(n11116), .A2(n9786), .ZN(n9157) );
  NAND2_X1 U11635 ( .A1(n9158), .A2(n9157), .ZN(n11145) );
  INV_X1 U11636 ( .A(n9159), .ZN(n9160) );
  NAND2_X1 U11637 ( .A1(n9161), .A2(n9160), .ZN(n9187) );
  NAND2_X1 U11638 ( .A1(n9187), .A2(n9185), .ZN(n9196) );
  MUX2_X1 U11639 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n9181), .Z(n9162) );
  NAND2_X1 U11640 ( .A1(n9162), .A2(SI_5_), .ZN(n9197) );
  OAI21_X1 U11641 ( .B1(n9162), .B2(SI_5_), .A(n9197), .ZN(n9189) );
  XNOR2_X1 U11642 ( .A(n9196), .B(n9189), .ZN(n11325) );
  NAND2_X1 U11643 ( .A1(n9166), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9165) );
  MUX2_X1 U11644 ( .A(n9165), .B(P2_IR_REG_31__SCAN_IN), .S(n9164), .Z(n9168)
         );
  INV_X1 U11645 ( .A(n9166), .ZN(n9167) );
  NAND2_X1 U11646 ( .A1(n9167), .A2(n9164), .ZN(n9215) );
  NAND2_X1 U11647 ( .A1(n9168), .A2(n9215), .ZN(n10300) );
  INV_X1 U11648 ( .A(n10300), .ZN(n10087) );
  AOI22_X1 U11649 ( .A1(n9456), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n10062), 
        .B2(n10087), .ZN(n9169) );
  NAND2_X1 U11650 ( .A1(n9924), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9178) );
  INV_X1 U11651 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n11149) );
  OR2_X1 U11652 ( .A1(n6666), .A2(n11149), .ZN(n9177) );
  INV_X1 U11653 ( .A(n9173), .ZN(n9171) );
  INV_X1 U11654 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9172) );
  NAND2_X1 U11655 ( .A1(n9173), .A2(n9172), .ZN(n9174) );
  NAND2_X1 U11656 ( .A1(n9204), .A2(n9174), .ZN(n11142) );
  OR2_X1 U11657 ( .A1(n9616), .A2(n11142), .ZN(n9176) );
  INV_X1 U11658 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10084) );
  OR2_X1 U11659 ( .A1(n9928), .A2(n10084), .ZN(n9175) );
  XNOR2_X1 U11660 ( .A(n11141), .B(n13887), .ZN(n11144) );
  NAND2_X1 U11661 ( .A1(n11145), .A2(n11144), .ZN(n9180) );
  OR2_X1 U11662 ( .A1(n15332), .A2(n13887), .ZN(n9179) );
  MUX2_X1 U11663 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n6670), .Z(n9182) );
  NAND2_X1 U11664 ( .A1(n9182), .A2(SI_6_), .ZN(n9211) );
  INV_X1 U11665 ( .A(n9182), .ZN(n9183) );
  NAND2_X1 U11666 ( .A1(n9183), .A2(n10161), .ZN(n9184) );
  AND2_X1 U11667 ( .A1(n9185), .A2(n9188), .ZN(n9186) );
  NAND2_X1 U11668 ( .A1(n9187), .A2(n9186), .ZN(n9194) );
  INV_X1 U11669 ( .A(n9188), .ZN(n9192) );
  INV_X1 U11670 ( .A(n9189), .ZN(n9195) );
  AND2_X1 U11671 ( .A1(n9195), .A2(n9199), .ZN(n9191) );
  NAND2_X1 U11672 ( .A1(n9196), .A2(n9195), .ZN(n9198) );
  NAND2_X1 U11673 ( .A1(n9215), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9200) );
  XNOR2_X1 U11674 ( .A(n9200), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10090) );
  AOI22_X1 U11675 ( .A1(n9456), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n10062), 
        .B2(n10090), .ZN(n9201) );
  NAND2_X1 U11676 ( .A1(n9202), .A2(n9201), .ZN(n10945) );
  NAND2_X1 U11677 ( .A1(n9924), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9209) );
  INV_X1 U11678 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n11128) );
  OR2_X1 U11679 ( .A1(n6666), .A2(n11128), .ZN(n9208) );
  INV_X1 U11680 ( .A(n9204), .ZN(n9203) );
  INV_X1 U11681 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n10933) );
  NAND2_X1 U11682 ( .A1(n9204), .A2(n10933), .ZN(n9205) );
  NAND2_X1 U11683 ( .A1(n9221), .A2(n9205), .ZN(n11129) );
  OR2_X1 U11684 ( .A1(n9616), .A2(n11129), .ZN(n9207) );
  INV_X1 U11685 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10089) );
  OR2_X1 U11686 ( .A1(n9928), .A2(n10089), .ZN(n9206) );
  NAND4_X1 U11687 ( .A1(n9207), .A2(n9208), .A3(n9209), .A4(n9206), .ZN(n13886) );
  NAND2_X1 U11688 ( .A1(n10945), .A2(n7021), .ZN(n9210) );
  NAND2_X1 U11689 ( .A1(n9212), .A2(n9211), .ZN(n9229) );
  MUX2_X1 U11690 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n9181), .Z(n9214) );
  NAND2_X1 U11691 ( .A1(n9214), .A2(SI_7_), .ZN(n9230) );
  OAI21_X1 U11692 ( .B1(n9214), .B2(SI_7_), .A(n9230), .ZN(n9227) );
  XNOR2_X1 U11693 ( .A(n9229), .B(n9227), .ZN(n11378) );
  OAI21_X1 U11694 ( .B1(n9215), .B2(P2_IR_REG_6__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9216) );
  XNOR2_X1 U11695 ( .A(n9216), .B(P2_IR_REG_7__SCAN_IN), .ZN(n10196) );
  AOI22_X1 U11696 ( .A1(n9456), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n10062), 
        .B2(n10196), .ZN(n9217) );
  INV_X1 U11697 ( .A(n11265), .ZN(n11027) );
  NAND2_X1 U11698 ( .A1(n9923), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9226) );
  INV_X1 U11699 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9219) );
  OR2_X1 U11700 ( .A1(n9343), .A2(n9219), .ZN(n9225) );
  NAND2_X1 U11701 ( .A1(n9221), .A2(n9220), .ZN(n9222) );
  NAND2_X1 U11702 ( .A1(n9239), .A2(n9222), .ZN(n11262) );
  OR2_X1 U11703 ( .A1(n9616), .A2(n11262), .ZN(n9224) );
  INV_X1 U11704 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n10092) );
  OR2_X1 U11705 ( .A1(n9928), .A2(n10092), .ZN(n9223) );
  XNOR2_X1 U11706 ( .A(n11027), .B(n11075), .ZN(n11022) );
  INV_X1 U11707 ( .A(n11022), .ZN(n11028) );
  INV_X1 U11708 ( .A(n11075), .ZN(n13885) );
  INV_X1 U11709 ( .A(n9227), .ZN(n9228) );
  NAND2_X1 U11710 ( .A1(n9229), .A2(n9228), .ZN(n9231) );
  MUX2_X1 U11711 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n9213), .Z(n9232) );
  NAND2_X1 U11712 ( .A1(n9232), .A2(SI_8_), .ZN(n9251) );
  OAI21_X1 U11713 ( .B1(SI_8_), .B2(n9232), .A(n9251), .ZN(n9248) );
  XNOR2_X1 U11714 ( .A(n9250), .B(n9248), .ZN(n11683) );
  OR2_X1 U11715 ( .A1(n9234), .A2(n9658), .ZN(n9235) );
  XNOR2_X1 U11716 ( .A(n9235), .B(P2_IR_REG_8__SCAN_IN), .ZN(n10267) );
  AOI22_X1 U11717 ( .A1(n9456), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n10062), 
        .B2(n10267), .ZN(n9236) );
  NAND2_X1 U11718 ( .A1(n9599), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9245) );
  INV_X1 U11719 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10093) );
  OR2_X1 U11720 ( .A1(n9928), .A2(n10093), .ZN(n9244) );
  NAND2_X1 U11721 ( .A1(n9239), .A2(n9238), .ZN(n9240) );
  NAND2_X1 U11722 ( .A1(n9261), .A2(n9240), .ZN(n11210) );
  OR2_X1 U11723 ( .A1(n9616), .A2(n11210), .ZN(n9243) );
  INV_X1 U11724 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n9241) );
  OR2_X1 U11725 ( .A1(n9420), .A2(n9241), .ZN(n9242) );
  XNOR2_X1 U11726 ( .A(n11215), .B(n11198), .ZN(n11069) );
  INV_X1 U11727 ( .A(n11069), .ZN(n11073) );
  NAND2_X1 U11728 ( .A1(n11074), .A2(n11073), .ZN(n9247) );
  INV_X1 U11729 ( .A(n11198), .ZN(n13884) );
  OR2_X1 U11730 ( .A1(n11247), .A2(n13884), .ZN(n9246) );
  NAND2_X1 U11731 ( .A1(n9247), .A2(n9246), .ZN(n11172) );
  INV_X1 U11732 ( .A(n9248), .ZN(n9249) );
  NAND2_X1 U11733 ( .A1(n9250), .A2(n9249), .ZN(n9252) );
  MUX2_X1 U11734 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n9213), .Z(n9253) );
  XNOR2_X1 U11735 ( .A(n9272), .B(n9270), .ZN(n11834) );
  NAND2_X1 U11736 ( .A1(n9234), .A2(n9254), .ZN(n9256) );
  NAND2_X1 U11737 ( .A1(n9256), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9255) );
  MUX2_X1 U11738 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9255), .S(
        P2_IR_REG_9__SCAN_IN), .Z(n9257) );
  AOI22_X1 U11739 ( .A1(n9456), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n10062), 
        .B2(n10455), .ZN(n9258) );
  NAND2_X1 U11740 ( .A1(n9259), .A2(n9258), .ZN(n11272) );
  NAND2_X1 U11741 ( .A1(n9923), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9266) );
  INV_X1 U11742 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n9260) );
  OR2_X1 U11743 ( .A1(n9343), .A2(n9260), .ZN(n9265) );
  NAND2_X1 U11744 ( .A1(n9261), .A2(n11275), .ZN(n9262) );
  NAND2_X1 U11745 ( .A1(n9282), .A2(n9262), .ZN(n11254) );
  OR2_X1 U11746 ( .A1(n9616), .A2(n11254), .ZN(n9264) );
  INV_X1 U11747 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10097) );
  OR2_X1 U11748 ( .A1(n9928), .A2(n10097), .ZN(n9263) );
  NAND4_X1 U11749 ( .A1(n9266), .A2(n9265), .A3(n9264), .A4(n9263), .ZN(n13882) );
  INV_X1 U11750 ( .A(n13882), .ZN(n9812) );
  AND2_X1 U11751 ( .A1(n11272), .A2(n9812), .ZN(n9267) );
  OR2_X1 U11752 ( .A1(n11172), .A2(n9267), .ZN(n9269) );
  OR2_X1 U11753 ( .A1(n11272), .A2(n9812), .ZN(n9268) );
  NAND2_X1 U11754 ( .A1(n9269), .A2(n9268), .ZN(n11561) );
  INV_X1 U11755 ( .A(n9270), .ZN(n9271) );
  NAND2_X1 U11756 ( .A1(n9272), .A2(n9271), .ZN(n9274) );
  MUX2_X1 U11757 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n9213), .Z(n9275) );
  XNOR2_X1 U11758 ( .A(n9291), .B(n9289), .ZN(n11973) );
  NAND2_X1 U11759 ( .A1(n9411), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9276) );
  XNOR2_X1 U11760 ( .A(n9276), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10199) );
  AOI22_X1 U11761 ( .A1(n9456), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n10062), 
        .B2(n10199), .ZN(n9277) );
  NAND2_X1 U11762 ( .A1(n9278), .A2(n9277), .ZN(n11571) );
  NAND2_X1 U11763 ( .A1(n9923), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9287) );
  INV_X1 U11764 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n9279) );
  OR2_X1 U11765 ( .A1(n9343), .A2(n9279), .ZN(n9286) );
  INV_X1 U11766 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9281) );
  NAND2_X1 U11767 ( .A1(n9282), .A2(n9281), .ZN(n9283) );
  NAND2_X1 U11768 ( .A1(n9299), .A2(n9283), .ZN(n11566) );
  OR2_X1 U11769 ( .A1(n9616), .A2(n11566), .ZN(n9285) );
  INV_X1 U11770 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n10099) );
  OR2_X1 U11771 ( .A1(n9928), .A2(n10099), .ZN(n9284) );
  NAND4_X1 U11772 ( .A1(n9287), .A2(n9286), .A3(n9285), .A4(n9284), .ZN(n13881) );
  INV_X1 U11773 ( .A(n13881), .ZN(n9818) );
  NAND2_X1 U11774 ( .A1(n11571), .A2(n9818), .ZN(n11644) );
  OR2_X1 U11775 ( .A1(n11571), .A2(n9818), .ZN(n9288) );
  NAND2_X1 U11776 ( .A1(n11644), .A2(n9288), .ZN(n11562) );
  NAND2_X1 U11777 ( .A1(n11559), .A2(n11644), .ZN(n9306) );
  INV_X1 U11778 ( .A(n9289), .ZN(n9290) );
  MUX2_X1 U11779 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n9213), .Z(n9308) );
  XNOR2_X1 U11780 ( .A(n9312), .B(n9311), .ZN(n12089) );
  NOR2_X1 U11781 ( .A1(n9411), .A2(P2_IR_REG_10__SCAN_IN), .ZN(n9314) );
  OR2_X1 U11782 ( .A1(n9314), .A2(n9658), .ZN(n9294) );
  XNOR2_X1 U11783 ( .A(n9294), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10100) );
  AOI22_X1 U11784 ( .A1(n9456), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n10062), 
        .B2(n10100), .ZN(n9295) );
  NAND2_X1 U11785 ( .A1(n9923), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9305) );
  INV_X1 U11786 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n9297) );
  OR2_X1 U11787 ( .A1(n9343), .A2(n9297), .ZN(n9304) );
  INV_X1 U11788 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9298) );
  NAND2_X1 U11789 ( .A1(n9299), .A2(n9298), .ZN(n9300) );
  NAND2_X1 U11790 ( .A1(n9320), .A2(n9300), .ZN(n11674) );
  OR2_X1 U11791 ( .A1(n9616), .A2(n11674), .ZN(n9303) );
  INV_X1 U11792 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n9301) );
  OR2_X1 U11793 ( .A1(n9928), .A2(n9301), .ZN(n9302) );
  XNOR2_X1 U11794 ( .A(n11910), .B(n13880), .ZN(n11643) );
  NAND2_X1 U11795 ( .A1(n9306), .A2(n11643), .ZN(n11647) );
  OR2_X1 U11796 ( .A1(n11680), .A2(n13880), .ZN(n9307) );
  INV_X1 U11797 ( .A(n9308), .ZN(n9309) );
  NAND2_X1 U11798 ( .A1(n9309), .A2(n10167), .ZN(n9310) );
  MUX2_X1 U11799 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n9213), .Z(n9331) );
  XNOR2_X1 U11800 ( .A(n9330), .B(n9329), .ZN(n12167) );
  AND2_X1 U11801 ( .A1(n9314), .A2(n9313), .ZN(n9335) );
  OR2_X1 U11802 ( .A1(n9335), .A2(n9658), .ZN(n9315) );
  XNOR2_X1 U11803 ( .A(n9315), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10101) );
  AOI22_X1 U11804 ( .A1(n9456), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n10062), 
        .B2(n10101), .ZN(n9316) );
  NAND2_X1 U11805 ( .A1(n9924), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n9326) );
  INV_X1 U11806 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n11596) );
  OR2_X1 U11807 ( .A1(n6666), .A2(n11596), .ZN(n9325) );
  INV_X1 U11808 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9319) );
  NAND2_X1 U11809 ( .A1(n9320), .A2(n9319), .ZN(n9321) );
  NAND2_X1 U11810 ( .A1(n9339), .A2(n9321), .ZN(n11928) );
  OR2_X1 U11811 ( .A1(n9616), .A2(n11928), .ZN(n9324) );
  INV_X1 U11812 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n9322) );
  OR2_X1 U11813 ( .A1(n9928), .A2(n9322), .ZN(n9323) );
  OAI21_X1 U11814 ( .B1(n11586), .B2(n11930), .A(n11914), .ZN(n9328) );
  NAND2_X1 U11815 ( .A1(n11586), .A2(n11930), .ZN(n9327) );
  INV_X1 U11816 ( .A(n9331), .ZN(n9332) );
  MUX2_X1 U11817 ( .A(n10287), .B(n10278), .S(n9213), .Z(n9349) );
  XNOR2_X1 U11818 ( .A(n9349), .B(SI_13_), .ZN(n9333) );
  XNOR2_X1 U11819 ( .A(n9353), .B(n9333), .ZN(n12239) );
  INV_X1 U11820 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n9334) );
  AND2_X1 U11821 ( .A1(n9335), .A2(n9334), .ZN(n9357) );
  OR2_X1 U11822 ( .A1(n9357), .A2(n9658), .ZN(n9336) );
  INV_X1 U11823 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n9356) );
  XNOR2_X1 U11824 ( .A(n9336), .B(n9356), .ZN(n10279) );
  INV_X1 U11825 ( .A(n10279), .ZN(n15242) );
  AOI22_X1 U11826 ( .A1(n15242), .A2(n10062), .B1(n9456), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n9337) );
  INV_X1 U11827 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n11964) );
  NAND2_X1 U11828 ( .A1(n9339), .A2(n11964), .ZN(n9340) );
  AND2_X1 U11829 ( .A1(n9361), .A2(n9340), .ZN(n11968) );
  NAND2_X1 U11830 ( .A1(n11968), .A2(n9341), .ZN(n9347) );
  INV_X1 U11831 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10054) );
  OR2_X1 U11832 ( .A1(n9420), .A2(n10054), .ZN(n9346) );
  INV_X1 U11833 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n9342) );
  OR2_X1 U11834 ( .A1(n9343), .A2(n9342), .ZN(n9345) );
  INV_X1 U11835 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10102) );
  OR2_X1 U11836 ( .A1(n9928), .A2(n10102), .ZN(n9344) );
  NAND2_X1 U11837 ( .A1(n15021), .A2(n13878), .ZN(n9348) );
  NAND2_X1 U11838 ( .A1(n9350), .A2(SI_13_), .ZN(n9351) );
  MUX2_X1 U11839 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n9213), .Z(n9370) );
  XNOR2_X1 U11840 ( .A(n9371), .B(n9370), .ZN(n12292) );
  NAND2_X1 U11841 ( .A1(n9357), .A2(n9356), .ZN(n9375) );
  NAND2_X1 U11842 ( .A1(n9375), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9358) );
  XNOR2_X1 U11843 ( .A(n9358), .B(P2_IR_REG_14__SCAN_IN), .ZN(n15258) );
  AOI22_X1 U11844 ( .A1(n15258), .A2(n10062), .B1(n9456), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n9359) );
  INV_X1 U11845 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n12160) );
  NAND2_X1 U11846 ( .A1(n9361), .A2(n12160), .ZN(n9362) );
  AND2_X1 U11847 ( .A1(n9381), .A2(n9362), .ZN(n14990) );
  NAND2_X1 U11848 ( .A1(n14990), .A2(n9341), .ZN(n9367) );
  NAND2_X1 U11849 ( .A1(n9923), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n9364) );
  NAND2_X1 U11850 ( .A1(n9924), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n9363) );
  AND2_X1 U11851 ( .A1(n9364), .A2(n9363), .ZN(n9366) );
  NAND2_X1 U11852 ( .A1(n9097), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n9365) );
  INV_X1 U11853 ( .A(n12144), .ZN(n13877) );
  AND2_X1 U11854 ( .A1(n15014), .A2(n13877), .ZN(n9368) );
  MUX2_X1 U11855 ( .A(n10763), .B(n10766), .S(n9213), .Z(n9372) );
  INV_X1 U11856 ( .A(n9372), .ZN(n9373) );
  NAND2_X1 U11857 ( .A1(n9373), .A2(SI_15_), .ZN(n9374) );
  XNOR2_X1 U11858 ( .A(n9387), .B(n9386), .ZN(n12443) );
  OR2_X1 U11859 ( .A1(n9375), .A2(P2_IR_REG_14__SCAN_IN), .ZN(n9376) );
  NAND2_X1 U11860 ( .A1(n9376), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9393) );
  XNOR2_X1 U11861 ( .A(n9393), .B(P2_IR_REG_15__SCAN_IN), .ZN(n10764) );
  AOI22_X1 U11862 ( .A1(n10764), .A2(n10062), .B1(n9456), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n9377) );
  INV_X1 U11863 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n9380) );
  NAND2_X1 U11864 ( .A1(n9381), .A2(n9380), .ZN(n9382) );
  NAND2_X1 U11865 ( .A1(n9418), .A2(n9382), .ZN(n12064) );
  OR2_X1 U11866 ( .A1(n12064), .A2(n9616), .ZN(n9385) );
  AOI22_X1 U11867 ( .A1(n9097), .A2(P2_REG1_REG_15__SCAN_IN), .B1(n9923), .B2(
        P2_REG2_REG_15__SCAN_IN), .ZN(n9384) );
  NAND2_X1 U11868 ( .A1(n9924), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n9383) );
  MUX2_X1 U11869 ( .A(n10879), .B(n10871), .S(n9213), .Z(n9389) );
  INV_X1 U11870 ( .A(n9389), .ZN(n9390) );
  NAND2_X1 U11871 ( .A1(n9390), .A2(SI_16_), .ZN(n9391) );
  XNOR2_X1 U11872 ( .A(n9407), .B(n9406), .ZN(n12627) );
  INV_X1 U11873 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n9392) );
  NAND2_X1 U11874 ( .A1(n9393), .A2(n9392), .ZN(n9394) );
  NAND2_X1 U11875 ( .A1(n9394), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9395) );
  XNOR2_X1 U11876 ( .A(n9395), .B(P2_IR_REG_16__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U11877 ( .A1(n11958), .A2(n10062), .B1(n9456), .B2(
        P1_DATAO_REG_16__SCAN_IN), .ZN(n9396) );
  XNOR2_X1 U11878 ( .A(n9418), .B(P2_REG3_REG_16__SCAN_IN), .ZN(n14974) );
  NAND2_X1 U11879 ( .A1(n14974), .A2(n9341), .ZN(n9402) );
  INV_X1 U11880 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10073) );
  NAND2_X1 U11881 ( .A1(n9923), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n9399) );
  NAND2_X1 U11882 ( .A1(n9924), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n9398) );
  OAI211_X1 U11883 ( .C1(n10073), .C2(n9928), .A(n9399), .B(n9398), .ZN(n9400)
         );
  INV_X1 U11884 ( .A(n9400), .ZN(n9401) );
  NAND2_X1 U11885 ( .A1(n9402), .A2(n9401), .ZN(n13875) );
  INV_X1 U11886 ( .A(n13875), .ZN(n9403) );
  XNOR2_X1 U11887 ( .A(n14975), .B(n9403), .ZN(n14969) );
  NAND2_X1 U11888 ( .A1(n14970), .A2(n14979), .ZN(n9405) );
  OR2_X1 U11889 ( .A1(n14975), .A2(n9403), .ZN(n9404) );
  NAND2_X1 U11890 ( .A1(n9405), .A2(n9404), .ZN(n12282) );
  MUX2_X1 U11891 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n9213), .Z(n9430) );
  XNOR2_X1 U11892 ( .A(n9430), .B(n10532), .ZN(n9409) );
  XNOR2_X1 U11893 ( .A(n9429), .B(n9409), .ZN(n12638) );
  OAI21_X1 U11894 ( .B1(n9411), .B2(n9410), .A(P2_IR_REG_31__SCAN_IN), .ZN(
        n9412) );
  XNOR2_X1 U11895 ( .A(n9412), .B(P2_IR_REG_17__SCAN_IN), .ZN(n12337) );
  AOI22_X1 U11896 ( .A1(n9456), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n10062), 
        .B2(n12337), .ZN(n9413) );
  INV_X1 U11897 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n9416) );
  INV_X1 U11898 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9415) );
  OAI21_X1 U11899 ( .B1(n9418), .B2(n9416), .A(n9415), .ZN(n9419) );
  NAND2_X1 U11900 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_REG3_REG_16__SCAN_IN), 
        .ZN(n9417) );
  AND2_X1 U11901 ( .A1(n9419), .A2(n9443), .ZN(n13809) );
  NAND2_X1 U11902 ( .A1(n13809), .A2(n9341), .ZN(n9425) );
  INV_X1 U11903 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n12345) );
  NAND2_X1 U11904 ( .A1(n9924), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n9422) );
  INV_X1 U11905 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n12286) );
  OR2_X1 U11906 ( .A1(n6666), .A2(n12286), .ZN(n9421) );
  OAI211_X1 U11907 ( .C1(n9928), .C2(n12345), .A(n9422), .B(n9421), .ZN(n9423)
         );
  INV_X1 U11908 ( .A(n9423), .ZN(n9424) );
  NAND2_X1 U11909 ( .A1(n9425), .A2(n9424), .ZN(n13874) );
  INV_X1 U11910 ( .A(n13874), .ZN(n13840) );
  NOR2_X1 U11911 ( .A1(n13699), .A2(n13840), .ZN(n9426) );
  NAND2_X1 U11912 ( .A1(n13699), .A2(n13840), .ZN(n9427) );
  NAND2_X1 U11913 ( .A1(n9430), .A2(SI_17_), .ZN(n9428) );
  INV_X1 U11914 ( .A(n9430), .ZN(n9431) );
  NAND2_X1 U11915 ( .A1(n9431), .A2(n10532), .ZN(n9432) );
  INV_X1 U11916 ( .A(SI_18_), .ZN(n10541) );
  NAND2_X1 U11917 ( .A1(n9475), .A2(n10541), .ZN(n9434) );
  MUX2_X1 U11918 ( .A(n11112), .B(n11113), .S(n9213), .Z(n9471) );
  NAND2_X1 U11919 ( .A1(n9435), .A2(n9471), .ZN(n9436) );
  NAND2_X1 U11920 ( .A1(n9437), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9438) );
  MUX2_X1 U11921 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9438), .S(
        P2_IR_REG_18__SCAN_IN), .Z(n9439) );
  AND2_X1 U11922 ( .A1(n9655), .A2(n9439), .ZN(n13897) );
  AOI22_X1 U11923 ( .A1(n9456), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n10062), 
        .B2(n13897), .ZN(n9440) );
  INV_X1 U11924 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n12341) );
  NAND2_X1 U11925 ( .A1(n9443), .A2(n12341), .ZN(n9444) );
  NAND2_X1 U11926 ( .A1(n9460), .A2(n9444), .ZN(n14087) );
  OR2_X1 U11927 ( .A1(n14087), .A2(n9616), .ZN(n9450) );
  INV_X1 U11928 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9447) );
  NAND2_X1 U11929 ( .A1(n9923), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9446) );
  NAND2_X1 U11930 ( .A1(n9924), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n9445) );
  OAI211_X1 U11931 ( .C1(n9447), .C2(n9928), .A(n9446), .B(n9445), .ZN(n9448)
         );
  INV_X1 U11932 ( .A(n9448), .ZN(n9449) );
  NAND2_X1 U11933 ( .A1(n9450), .A2(n9449), .ZN(n13873) );
  INV_X1 U11934 ( .A(n13873), .ZN(n13758) );
  AND2_X1 U11935 ( .A1(n14161), .A2(n13758), .ZN(n9451) );
  INV_X1 U11936 ( .A(n14161), .ZN(n14095) );
  NAND2_X1 U11937 ( .A1(n14095), .A2(n13873), .ZN(n9452) );
  MUX2_X1 U11938 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n9213), .Z(n9476) );
  XNOR2_X1 U11939 ( .A(n9476), .B(SI_19_), .ZN(n9473) );
  NAND2_X1 U11940 ( .A1(n9655), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9455) );
  AOI22_X1 U11941 ( .A1(n9456), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n10062), 
        .B2(n9709), .ZN(n9457) );
  INV_X1 U11942 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9459) );
  NAND2_X1 U11943 ( .A1(n9460), .A2(n9459), .ZN(n9461) );
  NAND2_X1 U11944 ( .A1(n9485), .A2(n9461), .ZN(n14069) );
  OR2_X1 U11945 ( .A1(n14069), .A2(n9616), .ZN(n9467) );
  INV_X1 U11946 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n9464) );
  NAND2_X1 U11947 ( .A1(n9923), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n9463) );
  NAND2_X1 U11948 ( .A1(n9924), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n9462) );
  OAI211_X1 U11949 ( .C1(n9464), .C2(n9928), .A(n9463), .B(n9462), .ZN(n9465)
         );
  INV_X1 U11950 ( .A(n9465), .ZN(n9466) );
  XNOR2_X1 U11951 ( .A(n14156), .B(n13872), .ZN(n14073) );
  NAND2_X1 U11952 ( .A1(n14063), .A2(n14073), .ZN(n9469) );
  NAND2_X1 U11953 ( .A1(n14072), .A2(n13872), .ZN(n9468) );
  NAND2_X1 U11954 ( .A1(n9469), .A2(n9468), .ZN(n14053) );
  INV_X1 U11955 ( .A(n9471), .ZN(n9470) );
  NOR2_X1 U11956 ( .A1(n9471), .A2(n10541), .ZN(n9472) );
  INV_X1 U11957 ( .A(n9476), .ZN(n9477) );
  NAND2_X1 U11958 ( .A1(n9477), .A2(n10767), .ZN(n9478) );
  OR2_X1 U11959 ( .A1(n9501), .A2(n11038), .ZN(n9497) );
  NAND2_X1 U11960 ( .A1(n9501), .A2(n11038), .ZN(n9479) );
  NAND2_X1 U11961 ( .A1(n9497), .A2(n9479), .ZN(n9480) );
  MUX2_X1 U11962 ( .A(n12708), .B(n7203), .S(n9213), .Z(n9500) );
  NAND2_X1 U11963 ( .A1(n9480), .A2(n9500), .ZN(n9481) );
  OR2_X1 U11964 ( .A1(n9948), .A2(n7203), .ZN(n9482) );
  INV_X1 U11965 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9484) );
  NAND2_X1 U11966 ( .A1(n9485), .A2(n9484), .ZN(n9486) );
  NAND2_X1 U11967 ( .A1(n9529), .A2(n9486), .ZN(n14049) );
  INV_X1 U11968 ( .A(n14049), .ZN(n9487) );
  NAND2_X1 U11969 ( .A1(n9487), .A2(n9341), .ZN(n9493) );
  INV_X1 U11970 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9490) );
  NAND2_X1 U11971 ( .A1(n9924), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n9489) );
  NAND2_X1 U11972 ( .A1(n9923), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9488) );
  OAI211_X1 U11973 ( .C1(n9490), .C2(n9928), .A(n9489), .B(n9488), .ZN(n9491)
         );
  INV_X1 U11974 ( .A(n9491), .ZN(n9492) );
  NAND2_X1 U11975 ( .A1(n14151), .A2(n13759), .ZN(n9495) );
  OR2_X1 U11976 ( .A1(n14151), .A2(n13759), .ZN(n9494) );
  NAND2_X1 U11977 ( .A1(n9495), .A2(n9494), .ZN(n14054) );
  MUX2_X1 U11978 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n9213), .Z(n9496) );
  NAND2_X1 U11979 ( .A1(n9496), .A2(SI_21_), .ZN(n9517) );
  OAI21_X1 U11980 ( .B1(SI_21_), .B2(n9496), .A(n9517), .ZN(n9504) );
  AND2_X1 U11981 ( .A1(n9497), .A2(n9504), .ZN(n9498) );
  NAND2_X1 U11982 ( .A1(n9499), .A2(n9498), .ZN(n9507) );
  NOR2_X1 U11983 ( .A1(n9502), .A2(SI_20_), .ZN(n9503) );
  NOR2_X1 U11984 ( .A1(n9504), .A2(n9503), .ZN(n9505) );
  NAND2_X1 U11985 ( .A1(n9507), .A2(n9518), .ZN(n12722) );
  OR2_X1 U11986 ( .A1(n12722), .A2(n9523), .ZN(n9509) );
  OR2_X1 U11987 ( .A1(n9948), .A2(n11512), .ZN(n9508) );
  XNOR2_X1 U11988 ( .A(n9529), .B(P2_REG3_REG_21__SCAN_IN), .ZN(n14038) );
  NAND2_X1 U11989 ( .A1(n14038), .A2(n9341), .ZN(n9515) );
  INV_X1 U11990 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n9512) );
  NAND2_X1 U11991 ( .A1(n9923), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n9511) );
  NAND2_X1 U11992 ( .A1(n9924), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n9510) );
  OAI211_X1 U11993 ( .C1(n9512), .C2(n9928), .A(n9511), .B(n9510), .ZN(n9513)
         );
  INV_X1 U11994 ( .A(n9513), .ZN(n9514) );
  NAND2_X1 U11995 ( .A1(n9515), .A2(n9514), .ZN(n13870) );
  INV_X1 U11996 ( .A(n13870), .ZN(n13831) );
  AND2_X1 U11997 ( .A1(n14146), .A2(n13831), .ZN(n9516) );
  INV_X1 U11998 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9520) );
  MUX2_X1 U11999 ( .A(n9520), .B(n11557), .S(n9213), .Z(n9521) );
  NAND2_X1 U12000 ( .A1(n12736), .A2(n9521), .ZN(n9522) );
  NAND2_X1 U12001 ( .A1(n9537), .A2(n9522), .ZN(n11555) );
  OR2_X1 U12002 ( .A1(n9948), .A2(n11557), .ZN(n9524) );
  AND2_X1 U12003 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(P2_REG3_REG_21__SCAN_IN), 
        .ZN(n9526) );
  INV_X1 U12004 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n13781) );
  INV_X1 U12005 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9528) );
  OAI21_X1 U12006 ( .B1(n9529), .B2(n13781), .A(n9528), .ZN(n9530) );
  NAND2_X1 U12007 ( .A1(n9543), .A2(n9530), .ZN(n14021) );
  OR2_X1 U12008 ( .A1(n14021), .A2(n9616), .ZN(n9536) );
  INV_X1 U12009 ( .A(P2_REG1_REG_22__SCAN_IN), .ZN(n9533) );
  NAND2_X1 U12010 ( .A1(n9923), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n9532) );
  NAND2_X1 U12011 ( .A1(n9924), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n9531) );
  OAI211_X1 U12012 ( .C1(n9533), .C2(n9928), .A(n9532), .B(n9531), .ZN(n9534)
         );
  INV_X1 U12013 ( .A(n9534), .ZN(n9535) );
  NAND2_X1 U12014 ( .A1(n9536), .A2(n9535), .ZN(n13869) );
  XNOR2_X1 U12015 ( .A(n14029), .B(n13869), .ZN(n14015) );
  MUX2_X1 U12016 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n9213), .Z(n9553) );
  XNOR2_X1 U12017 ( .A(n9553), .B(SI_23_), .ZN(n9538) );
  XNOR2_X1 U12018 ( .A(n9557), .B(n9538), .ZN(n12524) );
  OR2_X1 U12019 ( .A1(n9948), .A2(n11818), .ZN(n9539) );
  INV_X1 U12020 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n9542) );
  NAND2_X1 U12021 ( .A1(n9543), .A2(n9542), .ZN(n9544) );
  NAND2_X1 U12022 ( .A1(n9565), .A2(n9544), .ZN(n14003) );
  OR2_X1 U12023 ( .A1(n14003), .A2(n9616), .ZN(n9550) );
  INV_X1 U12024 ( .A(P2_REG1_REG_23__SCAN_IN), .ZN(n9547) );
  NAND2_X1 U12025 ( .A1(n9923), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n9546) );
  NAND2_X1 U12026 ( .A1(n9924), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n9545) );
  OAI211_X1 U12027 ( .C1(n9547), .C2(n9928), .A(n9546), .B(n9545), .ZN(n9548)
         );
  INV_X1 U12028 ( .A(n9548), .ZN(n9549) );
  NAND2_X1 U12029 ( .A1(n14136), .A2(n13832), .ZN(n9552) );
  OR2_X1 U12030 ( .A1(n14136), .A2(n13832), .ZN(n9551) );
  NAND2_X1 U12031 ( .A1(n9552), .A2(n9551), .ZN(n9989) );
  NAND2_X1 U12032 ( .A1(n13999), .A2(n14000), .ZN(n13998) );
  AND2_X2 U12033 ( .A1(n13998), .A2(n9552), .ZN(n13982) );
  NOR2_X1 U12034 ( .A1(n9554), .A2(n11447), .ZN(n9556) );
  NAND2_X1 U12035 ( .A1(n9554), .A2(n11447), .ZN(n9555) );
  MUX2_X1 U12036 ( .A(n12747), .B(n12142), .S(n9213), .Z(n9560) );
  NAND2_X1 U12037 ( .A1(n9561), .A2(n9560), .ZN(n9562) );
  OR2_X1 U12038 ( .A1(n9948), .A2(n12142), .ZN(n9563) );
  INV_X1 U12039 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n13815) );
  NAND2_X1 U12040 ( .A1(n9565), .A2(n13815), .ZN(n9566) );
  AND2_X1 U12041 ( .A1(n9577), .A2(n9566), .ZN(n13988) );
  INV_X1 U12042 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9569) );
  NAND2_X1 U12043 ( .A1(n9923), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n9568) );
  NAND2_X1 U12044 ( .A1(n9599), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n9567) );
  OAI211_X1 U12045 ( .C1(n9569), .C2(n9928), .A(n9568), .B(n9567), .ZN(n9570)
         );
  AOI21_X1 U12046 ( .B1(n13988), .B2(n9341), .A(n9570), .ZN(n13788) );
  INV_X1 U12047 ( .A(n13788), .ZN(n13867) );
  MUX2_X1 U12048 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n9213), .Z(n9589) );
  XNOR2_X1 U12049 ( .A(n9589), .B(SI_25_), .ZN(n9586) );
  OR2_X1 U12050 ( .A1(n9948), .A2(n12327), .ZN(n9573) );
  INV_X1 U12051 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9576) );
  NAND2_X1 U12052 ( .A1(n9577), .A2(n9576), .ZN(n9578) );
  NAND2_X1 U12053 ( .A1(n9597), .A2(n9578), .ZN(n13973) );
  OR2_X1 U12054 ( .A1(n13973), .A2(n9616), .ZN(n9584) );
  INV_X1 U12055 ( .A(P2_REG1_REG_25__SCAN_IN), .ZN(n9581) );
  NAND2_X1 U12056 ( .A1(n9924), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n9580) );
  NAND2_X1 U12057 ( .A1(n9923), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n9579) );
  OAI211_X1 U12058 ( .C1(n9928), .C2(n9581), .A(n9580), .B(n9579), .ZN(n9582)
         );
  INV_X1 U12059 ( .A(n9582), .ZN(n9583) );
  INV_X1 U12060 ( .A(n9586), .ZN(n9587) );
  INV_X1 U12061 ( .A(n9589), .ZN(n9590) );
  NAND2_X1 U12062 ( .A1(n9590), .A2(n12032), .ZN(n9591) );
  MUX2_X1 U12063 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n9213), .Z(n9607) );
  XNOR2_X1 U12064 ( .A(n9607), .B(n12139), .ZN(n9593) );
  OR2_X1 U12065 ( .A1(n9948), .A2(n12383), .ZN(n9594) );
  INV_X1 U12066 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n9596) );
  NAND2_X1 U12067 ( .A1(n9597), .A2(n9596), .ZN(n9598) );
  NAND2_X1 U12068 ( .A1(n13955), .A2(n9341), .ZN(n9605) );
  INV_X1 U12069 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9602) );
  NAND2_X1 U12070 ( .A1(n9923), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n9601) );
  NAND2_X1 U12071 ( .A1(n9599), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n9600) );
  OAI211_X1 U12072 ( .C1(n9602), .C2(n9928), .A(n9601), .B(n9600), .ZN(n9603)
         );
  INV_X1 U12073 ( .A(n9603), .ZN(n9604) );
  NAND2_X1 U12074 ( .A1(n14122), .A2(n13789), .ZN(n9971) );
  MUX2_X1 U12075 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n9213), .Z(n9623) );
  XNOR2_X1 U12076 ( .A(n9623), .B(SI_27_), .ZN(n9609) );
  OR2_X1 U12077 ( .A1(n9948), .A2(n12888), .ZN(n9610) );
  INV_X1 U12078 ( .A(n9614), .ZN(n9612) );
  NAND2_X1 U12079 ( .A1(n9612), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n9632) );
  INV_X1 U12080 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n9613) );
  NAND2_X1 U12081 ( .A1(n9614), .A2(n9613), .ZN(n9615) );
  NAND2_X1 U12082 ( .A1(n9632), .A2(n9615), .ZN(n13737) );
  OR2_X1 U12083 ( .A1(n13737), .A2(n9616), .ZN(n9622) );
  INV_X1 U12084 ( .A(P2_REG1_REG_27__SCAN_IN), .ZN(n9619) );
  NAND2_X1 U12085 ( .A1(n9924), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n9618) );
  NAND2_X1 U12086 ( .A1(n9923), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n9617) );
  OAI211_X1 U12087 ( .C1(n9619), .C2(n9928), .A(n9618), .B(n9617), .ZN(n9620)
         );
  INV_X1 U12088 ( .A(n9620), .ZN(n9621) );
  XNOR2_X1 U12089 ( .A(n14116), .B(n9907), .ZN(n9991) );
  INV_X1 U12090 ( .A(n9623), .ZN(n9624) );
  NAND2_X1 U12091 ( .A1(n9625), .A2(n9624), .ZN(n9627) );
  MUX2_X1 U12092 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(P1_DATAO_REG_28__SCAN_IN), 
        .S(n9213), .Z(n9645) );
  XNOR2_X1 U12093 ( .A(n9645), .B(n12946), .ZN(n9643) );
  OR2_X1 U12094 ( .A1(n9948), .A2(n14200), .ZN(n9628) );
  INV_X1 U12095 ( .A(n9632), .ZN(n9630) );
  INV_X1 U12096 ( .A(n9714), .ZN(n9634) );
  INV_X1 U12097 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n9631) );
  NAND2_X1 U12098 ( .A1(n9632), .A2(n9631), .ZN(n9633) );
  NAND2_X1 U12099 ( .A1(n13934), .A2(n9341), .ZN(n9640) );
  INV_X1 U12100 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n9637) );
  NAND2_X1 U12101 ( .A1(n9923), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n9636) );
  NAND2_X1 U12102 ( .A1(n9924), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n9635) );
  OAI211_X1 U12103 ( .C1(n9637), .C2(n9928), .A(n9636), .B(n9635), .ZN(n9638)
         );
  INV_X1 U12104 ( .A(n9638), .ZN(n9639) );
  NAND2_X1 U12105 ( .A1(n14110), .A2(n13769), .ZN(n9641) );
  INV_X1 U12106 ( .A(n13923), .ZN(n13928) );
  NAND2_X1 U12107 ( .A1(n14116), .A2(n9907), .ZN(n13926) );
  NAND3_X1 U12108 ( .A1(n13925), .A2(n13928), .A3(n13926), .ZN(n13927) );
  INV_X1 U12109 ( .A(n9645), .ZN(n9646) );
  NAND2_X1 U12110 ( .A1(n9646), .A2(n12946), .ZN(n9647) );
  MUX2_X1 U12111 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n9213), .Z(n9915) );
  XNOR2_X1 U12112 ( .A(n9915), .B(n13689), .ZN(n9913) );
  OR2_X1 U12113 ( .A1(n9948), .A2(n14193), .ZN(n9649) );
  INV_X1 U12114 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n9652) );
  NAND2_X1 U12115 ( .A1(n9923), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n9651) );
  NAND2_X1 U12116 ( .A1(n9924), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n9650) );
  OAI211_X1 U12117 ( .C1(n9652), .C2(n9928), .A(n9651), .B(n9650), .ZN(n9653)
         );
  AOI21_X1 U12118 ( .B1(n9714), .B2(n9341), .A(n9653), .ZN(n13773) );
  INV_X1 U12119 ( .A(n13773), .ZN(n13862) );
  NAND2_X1 U12120 ( .A1(n9659), .A2(n9660), .ZN(n9675) );
  INV_X1 U12121 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n9656) );
  XNOR2_X2 U12122 ( .A(n9657), .B(n9656), .ZN(n11556) );
  OR2_X1 U12123 ( .A1(n11556), .A2(n9758), .ZN(n9666) );
  XNOR2_X1 U12124 ( .A(n9661), .B(n9660), .ZN(n9710) );
  INV_X1 U12125 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n9662) );
  OR2_X1 U12126 ( .A1(n11287), .A2(n9664), .ZN(n9665) );
  INV_X1 U12127 ( .A(n11556), .ZN(n10018) );
  INV_X1 U12128 ( .A(n10070), .ZN(n10066) );
  NAND2_X1 U12129 ( .A1(n10692), .A2(n10070), .ZN(n13841) );
  INV_X1 U12130 ( .A(P2_B_REG_SCAN_IN), .ZN(n9679) );
  NOR2_X1 U12131 ( .A1(n9668), .A2(n9679), .ZN(n9669) );
  NOR2_X1 U12132 ( .A1(n13841), .A2(n9669), .ZN(n13913) );
  INV_X1 U12133 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n9672) );
  NAND2_X1 U12134 ( .A1(n9923), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n9671) );
  NAND2_X1 U12135 ( .A1(n9924), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9670) );
  OAI211_X1 U12136 ( .C1(n9928), .C2(n9672), .A(n9671), .B(n9670), .ZN(n13861)
         );
  INV_X1 U12137 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n9701) );
  NAND2_X1 U12138 ( .A1(n9702), .A2(n9701), .ZN(n9677) );
  NAND2_X1 U12139 ( .A1(n9677), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9678) );
  XNOR2_X1 U12140 ( .A(n12141), .B(n9679), .ZN(n9683) );
  NAND2_X1 U12141 ( .A1(n6782), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9680) );
  MUX2_X1 U12142 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9680), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n9682) );
  NAND2_X1 U12143 ( .A1(n9682), .A2(n9681), .ZN(n12325) );
  NAND2_X1 U12144 ( .A1(n9683), .A2(n12325), .ZN(n9687) );
  NAND2_X1 U12145 ( .A1(n9681), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9684) );
  MUX2_X1 U12146 ( .A(P2_IR_REG_31__SCAN_IN), .B(n9684), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n9686) );
  NAND2_X1 U12147 ( .A1(n9686), .A2(n9685), .ZN(n12384) );
  INV_X1 U12148 ( .A(n12384), .ZN(n9704) );
  INV_X1 U12149 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n15290) );
  NAND2_X1 U12150 ( .A1(n15283), .A2(n15290), .ZN(n9689) );
  NAND2_X1 U12151 ( .A1(n12384), .A2(n12325), .ZN(n9688) );
  NAND2_X1 U12152 ( .A1(n9689), .A2(n9688), .ZN(n10939) );
  INV_X1 U12153 ( .A(n10939), .ZN(n10687) );
  NOR4_X1 U12154 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n9698) );
  OR4_X1 U12155 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n9695) );
  NOR4_X1 U12156 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n9693) );
  NOR4_X1 U12157 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n9692) );
  NOR4_X1 U12158 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n9691) );
  NOR4_X1 U12159 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n9690) );
  NAND4_X1 U12160 ( .A1(n9693), .A2(n9692), .A3(n9691), .A4(n9690), .ZN(n9694)
         );
  NOR4_X1 U12161 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        n9695), .A4(n9694), .ZN(n9697) );
  NOR4_X1 U12162 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n9696) );
  NAND3_X1 U12163 ( .A1(n9698), .A2(n9697), .A3(n9696), .ZN(n9699) );
  NOR2_X1 U12164 ( .A1(n12384), .A2(n12325), .ZN(n9700) );
  NAND2_X1 U12165 ( .A1(n12141), .A2(n9700), .ZN(n10021) );
  XNOR2_X1 U12166 ( .A(n9702), .B(n9701), .ZN(n10063) );
  NAND2_X1 U12167 ( .A1(n11287), .A2(n9758), .ZN(n10683) );
  NAND2_X1 U12168 ( .A1(n10692), .A2(n10683), .ZN(n9703) );
  AND2_X1 U12169 ( .A1(n9708), .A2(n9703), .ZN(n10750) );
  NAND2_X1 U12170 ( .A1(n10750), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10938) );
  NOR2_X1 U12171 ( .A1(n10686), .A2(n10938), .ZN(n9707) );
  INV_X1 U12172 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n15286) );
  NAND2_X1 U12173 ( .A1(n15283), .A2(n15286), .ZN(n9706) );
  OR2_X1 U12174 ( .A1(n12141), .A2(n9704), .ZN(n9705) );
  NAND3_X1 U12175 ( .A1(n10687), .A2(n9707), .A3(n15287), .ZN(n9712) );
  AND2_X2 U12176 ( .A1(n9710), .A2(n9709), .ZN(n11063) );
  INV_X1 U12177 ( .A(n11063), .ZN(n9711) );
  INV_X1 U12178 ( .A(n10688), .ZN(n10937) );
  INV_X2 U12179 ( .A(n14088), .ZN(n15269) );
  AND2_X1 U12180 ( .A1(n15275), .A2(n15306), .ZN(n15277) );
  INV_X1 U12181 ( .A(n15314), .ZN(n11297) );
  NAND2_X1 U12182 ( .A1(n15277), .A2(n11297), .ZN(n11296) );
  INV_X1 U12183 ( .A(n10945), .ZN(n11130) );
  OR2_X2 U12184 ( .A1(n11072), .A2(n11215), .ZN(n11170) );
  INV_X1 U12185 ( .A(n11571), .ZN(n15341) );
  NAND2_X1 U12186 ( .A1(n11642), .A2(n11680), .ZN(n11594) );
  OR2_X2 U12187 ( .A1(n11594), .A2(n11930), .ZN(n11885) );
  NOR2_X1 U12188 ( .A1(n14161), .A2(n14092), .ZN(n14090) );
  NAND2_X1 U12189 ( .A1(n14067), .A2(n14052), .ZN(n14048) );
  OR2_X2 U12190 ( .A1(n14048), .A2(n14146), .ZN(n14036) );
  NAND2_X1 U12191 ( .A1(n13957), .A2(n13976), .ZN(n13954) );
  AND2_X4 U12192 ( .A1(n9713), .A2(n11287), .ZN(n15274) );
  AOI211_X1 U12193 ( .C1(n14106), .C2(n13932), .A(n14091), .B(n13918), .ZN(
        n14105) );
  NOR2_X2 U12194 ( .A1(n15269), .A2(n9709), .ZN(n15279) );
  OR2_X1 U12195 ( .A1(n11062), .A2(n11287), .ZN(n10684) );
  INV_X1 U12196 ( .A(n14086), .ZN(n15268) );
  AOI22_X1 U12197 ( .A1(n9714), .A2(n15268), .B1(P2_REG2_REG_29__SCAN_IN), 
        .B2(n15269), .ZN(n9715) );
  OAI21_X1 U12198 ( .B1(n9934), .B2(n14094), .A(n9715), .ZN(n9716) );
  INV_X1 U12199 ( .A(n11290), .ZN(n11289) );
  INV_X1 U12200 ( .A(n11468), .ZN(n9719) );
  NAND2_X1 U12201 ( .A1(n9719), .A2(n11466), .ZN(n9721) );
  NAND2_X1 U12202 ( .A1(n15300), .A2(n10903), .ZN(n9720) );
  NAND2_X1 U12203 ( .A1(n9721), .A2(n9720), .ZN(n15273) );
  NAND2_X1 U12204 ( .A1(n15273), .A2(n15272), .ZN(n9724) );
  NAND2_X1 U12205 ( .A1(n15306), .A2(n9722), .ZN(n9723) );
  OR2_X1 U12206 ( .A1(n15314), .A2(n13889), .ZN(n9725) );
  NAND2_X1 U12207 ( .A1(n9726), .A2(n9725), .ZN(n11114) );
  NAND2_X1 U12208 ( .A1(n11114), .A2(n9976), .ZN(n9728) );
  OR2_X1 U12209 ( .A1(n11116), .A2(n13888), .ZN(n9727) );
  AND2_X1 U12210 ( .A1(n15332), .A2(n9794), .ZN(n9729) );
  OR2_X1 U12211 ( .A1(n11265), .A2(n11075), .ZN(n9730) );
  NAND2_X1 U12212 ( .A1(n9731), .A2(n9730), .ZN(n11070) );
  NAND2_X1 U12213 ( .A1(n11070), .A2(n11069), .ZN(n9733) );
  OR2_X1 U12214 ( .A1(n11247), .A2(n11198), .ZN(n9732) );
  XNOR2_X1 U12215 ( .A(n11272), .B(n13882), .ZN(n11171) );
  INV_X1 U12216 ( .A(n11171), .ZN(n11168) );
  NAND2_X1 U12217 ( .A1(n11272), .A2(n13882), .ZN(n9734) );
  NAND2_X1 U12218 ( .A1(n11571), .A2(n13881), .ZN(n9735) );
  NOR2_X1 U12219 ( .A1(n11680), .A2(n11587), .ZN(n9736) );
  INV_X1 U12220 ( .A(n11914), .ZN(n13879) );
  NAND2_X1 U12221 ( .A1(n11930), .A2(n13879), .ZN(n9973) );
  NAND2_X1 U12222 ( .A1(n11593), .A2(n9973), .ZN(n9737) );
  OR2_X1 U12223 ( .A1(n11930), .A2(n13879), .ZN(n9974) );
  NAND2_X1 U12224 ( .A1(n9737), .A2(n9974), .ZN(n11883) );
  OR2_X1 U12225 ( .A1(n15021), .A2(n11589), .ZN(n9738) );
  NAND2_X1 U12226 ( .A1(n11883), .A2(n9738), .ZN(n9740) );
  NAND2_X1 U12227 ( .A1(n15021), .A2(n11589), .ZN(n9739) );
  NAND2_X1 U12228 ( .A1(n9740), .A2(n9739), .ZN(n14992) );
  INV_X1 U12229 ( .A(n15014), .ZN(n14991) );
  XNOR2_X1 U12230 ( .A(n14991), .B(n12144), .ZN(n14985) );
  INV_X1 U12231 ( .A(n14985), .ZN(n14993) );
  XNOR2_X1 U12232 ( .A(n12363), .B(n12358), .ZN(n12063) );
  NAND2_X1 U12233 ( .A1(n15008), .A2(n12358), .ZN(n9742) );
  NAND2_X1 U12234 ( .A1(n14975), .A2(n13875), .ZN(n9743) );
  NAND2_X1 U12235 ( .A1(n14976), .A2(n9743), .ZN(n12278) );
  XNOR2_X1 U12236 ( .A(n13699), .B(n13874), .ZN(n9984) );
  NAND2_X1 U12237 ( .A1(n12278), .A2(n12281), .ZN(n12280) );
  NAND2_X1 U12238 ( .A1(n13699), .A2(n13874), .ZN(n9744) );
  XNOR2_X1 U12239 ( .A(n14161), .B(n13873), .ZN(n14082) );
  NAND2_X1 U12240 ( .A1(n14095), .A2(n13758), .ZN(n9745) );
  NOR2_X1 U12241 ( .A1(n14052), .A2(n13759), .ZN(n9746) );
  NAND2_X1 U12242 ( .A1(n14052), .A2(n13759), .ZN(n9747) );
  XNOR2_X1 U12243 ( .A(n14146), .B(n13870), .ZN(n14041) );
  INV_X1 U12244 ( .A(n14041), .ZN(n9748) );
  NAND2_X1 U12245 ( .A1(n14042), .A2(n9748), .ZN(n9750) );
  OR2_X1 U12246 ( .A1(n14146), .A2(n13870), .ZN(n9749) );
  NAND2_X1 U12247 ( .A1(n9750), .A2(n9749), .ZN(n14012) );
  INV_X1 U12248 ( .A(n14012), .ZN(n9752) );
  NAND2_X1 U12249 ( .A1(n14029), .A2(n13869), .ZN(n9753) );
  NAND2_X1 U12250 ( .A1(n13957), .A2(n13789), .ZN(n9754) );
  INV_X1 U12251 ( .A(n14116), .ZN(n13943) );
  AOI22_X1 U12252 ( .A1(n13924), .A2(n13923), .B1(n14110), .B2(n13863), .ZN(
        n9755) );
  INV_X1 U12253 ( .A(n9762), .ZN(n9756) );
  OR2_X1 U12254 ( .A1(n14078), .A2(n9756), .ZN(n11659) );
  OR2_X1 U12255 ( .A1(n14078), .A2(n15335), .ZN(n9760) );
  NAND2_X1 U12256 ( .A1(n11659), .A2(n9760), .ZN(n15280) );
  INV_X1 U12257 ( .A(n9764), .ZN(n9767) );
  AOI21_X1 U12258 ( .B1(n9709), .B2(n11556), .A(n10723), .ZN(n9765) );
  INV_X1 U12259 ( .A(n9768), .ZN(n9771) );
  INV_X1 U12260 ( .A(n9769), .ZN(n9770) );
  NAND2_X1 U12261 ( .A1(n9774), .A2(n9775), .ZN(n9779) );
  INV_X1 U12262 ( .A(n9774), .ZN(n9777) );
  INV_X1 U12263 ( .A(n9775), .ZN(n9776) );
  AOI22_X1 U12264 ( .A1(n9779), .A2(n9778), .B1(n9777), .B2(n9776), .ZN(n9782)
         );
  AOI22_X1 U12265 ( .A1(n15314), .A2(n9870), .B1(n9826), .B2(n13889), .ZN(
        n9781) );
  OAI22_X1 U12266 ( .A1(n11297), .A2(n9870), .B1(n10902), .B2(n10005), .ZN(
        n9780) );
  NAND2_X1 U12267 ( .A1(n9782), .A2(n9781), .ZN(n9783) );
  NAND2_X1 U12268 ( .A1(n9784), .A2(n9783), .ZN(n9789) );
  AOI22_X1 U12269 ( .A1(n11116), .A2(n9826), .B1(n13888), .B2(n9870), .ZN(
        n9790) );
  INV_X1 U12270 ( .A(n9790), .ZN(n9785) );
  NAND2_X1 U12271 ( .A1(n9789), .A2(n9785), .ZN(n9788) );
  OAI22_X1 U12272 ( .A1(n7049), .A2(n10005), .B1(n9786), .B2(n9870), .ZN(n9787) );
  NAND2_X1 U12273 ( .A1(n9788), .A2(n9787), .ZN(n9793) );
  INV_X1 U12274 ( .A(n9789), .ZN(n9791) );
  NAND2_X1 U12275 ( .A1(n9791), .A2(n9790), .ZN(n9792) );
  OAI22_X1 U12276 ( .A1(n15332), .A2(n10005), .B1(n9794), .B2(n9870), .ZN(
        n9796) );
  NAND2_X1 U12277 ( .A1(n9795), .A2(n9796), .ZN(n9800) );
  OAI22_X1 U12278 ( .A1(n15332), .A2(n9870), .B1(n9794), .B2(n9826), .ZN(n9799) );
  INV_X1 U12279 ( .A(n9795), .ZN(n9798) );
  INV_X1 U12280 ( .A(n9796), .ZN(n9797) );
  AOI22_X1 U12281 ( .A1(n10945), .A2(n9826), .B1(n13886), .B2(n9908), .ZN(
        n9802) );
  OAI22_X1 U12282 ( .A1(n11130), .A2(n9826), .B1(n7021), .B2(n9908), .ZN(n9801) );
  OAI22_X1 U12283 ( .A1(n11265), .A2(n10005), .B1(n11075), .B2(n9908), .ZN(
        n9804) );
  NAND2_X1 U12284 ( .A1(n9803), .A2(n9804), .ZN(n9808) );
  OAI22_X1 U12285 ( .A1(n11265), .A2(n9870), .B1(n11075), .B2(n10005), .ZN(
        n9807) );
  INV_X1 U12286 ( .A(n9804), .ZN(n9805) );
  OAI22_X1 U12287 ( .A1(n11247), .A2(n9826), .B1(n11198), .B2(n9870), .ZN(
        n9811) );
  AOI22_X1 U12288 ( .A1(n11272), .A2(n9870), .B1(n9826), .B2(n13882), .ZN(
        n9813) );
  INV_X1 U12289 ( .A(n11272), .ZN(n11277) );
  OAI22_X1 U12290 ( .A1(n11277), .A2(n9870), .B1(n9812), .B2(n9826), .ZN(n9816) );
  AND2_X1 U12291 ( .A1(n9814), .A2(n9813), .ZN(n9815) );
  AOI22_X1 U12292 ( .A1(n11571), .A2(n10005), .B1(n13881), .B2(n9870), .ZN(
        n9820) );
  OAI22_X1 U12293 ( .A1(n15341), .A2(n10005), .B1(n9818), .B2(n9908), .ZN(
        n9819) );
  OAI21_X1 U12294 ( .B1(n9821), .B2(n9820), .A(n9819), .ZN(n9823) );
  NAND2_X1 U12295 ( .A1(n9821), .A2(n9820), .ZN(n9822) );
  OAI22_X1 U12296 ( .A1(n11680), .A2(n10005), .B1(n11587), .B2(n9870), .ZN(
        n9825) );
  AOI22_X1 U12297 ( .A1(n11910), .A2(n9826), .B1(n13880), .B2(n9870), .ZN(
        n9824) );
  OAI22_X1 U12298 ( .A1(n15026), .A2(n9908), .B1(n11914), .B2(n9826), .ZN(
        n9829) );
  AOI22_X1 U12299 ( .A1(n11930), .A2(n9870), .B1(n9826), .B2(n13879), .ZN(
        n9827) );
  AOI21_X1 U12300 ( .B1(n9830), .B2(n9829), .A(n9827), .ZN(n9828) );
  INV_X1 U12301 ( .A(n9828), .ZN(n9831) );
  NAND2_X1 U12302 ( .A1(n9831), .A2(n7631), .ZN(n9835) );
  OAI22_X1 U12303 ( .A1(n15021), .A2(n10005), .B1(n11589), .B2(n9908), .ZN(
        n9834) );
  AOI22_X1 U12304 ( .A1(n11888), .A2(n10005), .B1(n13878), .B2(n9870), .ZN(
        n9832) );
  AOI21_X1 U12305 ( .B1(n9835), .B2(n9834), .A(n9832), .ZN(n9833) );
  INV_X1 U12306 ( .A(n9833), .ZN(n9836) );
  OAI22_X1 U12307 ( .A1(n15014), .A2(n9908), .B1(n12144), .B2(n10005), .ZN(
        n9838) );
  AOI22_X1 U12308 ( .A1(n14991), .A2(n9908), .B1(n10005), .B2(n13877), .ZN(
        n9837) );
  AND2_X1 U12309 ( .A1(n13874), .A2(n10005), .ZN(n9839) );
  AOI21_X1 U12310 ( .B1(n13699), .B2(n9908), .A(n9839), .ZN(n9857) );
  NAND2_X1 U12311 ( .A1(n13699), .A2(n10005), .ZN(n9841) );
  NAND2_X1 U12312 ( .A1(n13874), .A2(n9870), .ZN(n9840) );
  NAND2_X1 U12313 ( .A1(n9841), .A2(n9840), .ZN(n9855) );
  AND2_X1 U12314 ( .A1(n13875), .A2(n10005), .ZN(n9842) );
  AOI21_X1 U12315 ( .B1(n14975), .B2(n9908), .A(n9842), .ZN(n9852) );
  NAND2_X1 U12316 ( .A1(n14975), .A2(n10005), .ZN(n9844) );
  NAND2_X1 U12317 ( .A1(n13875), .A2(n9908), .ZN(n9843) );
  NAND2_X1 U12318 ( .A1(n9844), .A2(n9843), .ZN(n9851) );
  AOI22_X1 U12319 ( .A1(n9857), .A2(n9855), .B1(n9852), .B2(n9851), .ZN(n9850)
         );
  AOI22_X1 U12320 ( .A1(n12363), .A2(n10005), .B1(n13876), .B2(n9870), .ZN(
        n9849) );
  INV_X1 U12321 ( .A(n9849), .ZN(n9846) );
  OAI22_X1 U12322 ( .A1(n15008), .A2(n10005), .B1(n12358), .B2(n9870), .ZN(
        n9848) );
  NAND2_X1 U12323 ( .A1(n9846), .A2(n9845), .ZN(n9847) );
  NAND3_X1 U12324 ( .A1(n9850), .A2(n9849), .A3(n9848), .ZN(n9863) );
  INV_X1 U12325 ( .A(n9851), .ZN(n9854) );
  INV_X1 U12326 ( .A(n9852), .ZN(n9853) );
  NAND2_X1 U12327 ( .A1(n9854), .A2(n9853), .ZN(n9856) );
  INV_X1 U12328 ( .A(n13699), .ZN(n14167) );
  NAND3_X1 U12329 ( .A1(n9856), .A2(n13840), .A3(n14167), .ZN(n9861) );
  INV_X1 U12330 ( .A(n9855), .ZN(n9860) );
  INV_X1 U12331 ( .A(n9856), .ZN(n9859) );
  INV_X1 U12332 ( .A(n9857), .ZN(n9858) );
  AOI22_X1 U12333 ( .A1(n9861), .A2(n9860), .B1(n9859), .B2(n9858), .ZN(n9862)
         );
  AOI22_X1 U12334 ( .A1(n14161), .A2(n10005), .B1(n13873), .B2(n9870), .ZN(
        n9866) );
  OAI22_X1 U12335 ( .A1(n14095), .A2(n10005), .B1(n13758), .B2(n9908), .ZN(
        n9865) );
  OAI21_X1 U12336 ( .B1(n9867), .B2(n9866), .A(n9865), .ZN(n9869) );
  NAND2_X1 U12337 ( .A1(n9867), .A2(n9866), .ZN(n9868) );
  NAND2_X1 U12338 ( .A1(n9869), .A2(n9868), .ZN(n9871) );
  OAI22_X1 U12339 ( .A1(n14072), .A2(n10005), .B1(n13842), .B2(n9908), .ZN(
        n9872) );
  OAI22_X1 U12340 ( .A1(n14072), .A2(n9870), .B1(n13842), .B2(n10005), .ZN(
        n9874) );
  INV_X1 U12341 ( .A(n9872), .ZN(n9873) );
  OAI22_X1 U12342 ( .A1(n14052), .A2(n9908), .B1(n13759), .B2(n10005), .ZN(
        n9875) );
  OAI22_X1 U12343 ( .A1(n14052), .A2(n10005), .B1(n13759), .B2(n9908), .ZN(
        n9876) );
  AOI22_X1 U12344 ( .A1(n14146), .A2(n9870), .B1(n10005), .B2(n13870), .ZN(
        n9878) );
  INV_X1 U12345 ( .A(n14146), .ZN(n14040) );
  OAI22_X1 U12346 ( .A1(n14040), .A2(n9908), .B1(n13831), .B2(n10005), .ZN(
        n9877) );
  OAI21_X1 U12347 ( .B1(n9879), .B2(n9878), .A(n9877), .ZN(n9881) );
  NAND2_X1 U12348 ( .A1(n9879), .A2(n9878), .ZN(n9880) );
  AOI22_X1 U12349 ( .A1(n14029), .A2(n10005), .B1(n13869), .B2(n9870), .ZN(
        n9883) );
  INV_X1 U12350 ( .A(n9883), .ZN(n9882) );
  AOI22_X1 U12351 ( .A1(n14029), .A2(n9870), .B1(n10005), .B2(n13869), .ZN(
        n9884) );
  OAI22_X1 U12352 ( .A1(n14008), .A2(n9826), .B1(n13832), .B2(n9908), .ZN(
        n9885) );
  OAI22_X1 U12353 ( .A1(n14008), .A2(n9908), .B1(n13832), .B2(n10005), .ZN(
        n9886) );
  NAND2_X1 U12354 ( .A1(n9889), .A2(n9890), .ZN(n9888) );
  OAI22_X1 U12355 ( .A1(n13990), .A2(n10005), .B1(n13788), .B2(n9870), .ZN(
        n9887) );
  NAND2_X1 U12356 ( .A1(n9888), .A2(n9887), .ZN(n9894) );
  INV_X1 U12357 ( .A(n9889), .ZN(n9892) );
  INV_X1 U12358 ( .A(n9890), .ZN(n9891) );
  NAND2_X1 U12359 ( .A1(n9892), .A2(n9891), .ZN(n9893) );
  OAI22_X1 U12360 ( .A1(n13975), .A2(n10005), .B1(n9895), .B2(n9870), .ZN(
        n9899) );
  NAND2_X1 U12361 ( .A1(n9898), .A2(n9899), .ZN(n9897) );
  OAI22_X1 U12362 ( .A1(n13975), .A2(n9908), .B1(n9895), .B2(n10005), .ZN(
        n9896) );
  NAND2_X1 U12363 ( .A1(n9897), .A2(n9896), .ZN(n9903) );
  INV_X1 U12364 ( .A(n9898), .ZN(n9901) );
  INV_X1 U12365 ( .A(n9899), .ZN(n9900) );
  NAND2_X1 U12366 ( .A1(n9901), .A2(n9900), .ZN(n9902) );
  NAND2_X1 U12367 ( .A1(n9903), .A2(n9902), .ZN(n9904) );
  OAI22_X1 U12368 ( .A1(n13957), .A2(n9908), .B1(n13789), .B2(n10005), .ZN(
        n9905) );
  OAI22_X1 U12369 ( .A1(n13957), .A2(n10005), .B1(n13789), .B2(n9870), .ZN(
        n9906) );
  AOI22_X1 U12370 ( .A1(n14116), .A2(n9870), .B1(n10005), .B2(n13864), .ZN(
        n9956) );
  OAI22_X1 U12371 ( .A1(n13943), .A2(n9908), .B1(n9907), .B2(n10005), .ZN(
        n9909) );
  AND2_X1 U12372 ( .A1(n13863), .A2(n9908), .ZN(n9910) );
  AOI21_X1 U12373 ( .B1(n14110), .B2(n10005), .A(n9910), .ZN(n9961) );
  NAND2_X1 U12374 ( .A1(n14110), .A2(n9870), .ZN(n9912) );
  NAND2_X1 U12375 ( .A1(n13863), .A2(n10005), .ZN(n9911) );
  NAND2_X1 U12376 ( .A1(n9912), .A2(n9911), .ZN(n9960) );
  INV_X1 U12377 ( .A(n9915), .ZN(n9916) );
  NAND2_X1 U12378 ( .A1(n9916), .A2(n13689), .ZN(n9935) );
  MUX2_X1 U12379 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n9213), .Z(n9917) );
  NAND2_X1 U12380 ( .A1(n9917), .A2(SI_30_), .ZN(n9939) );
  INV_X1 U12381 ( .A(n9917), .ZN(n9918) );
  NAND2_X1 U12382 ( .A1(n9918), .A2(n13132), .ZN(n9936) );
  AND2_X1 U12383 ( .A1(n9939), .A2(n9936), .ZN(n9919) );
  OR2_X1 U12384 ( .A1(n9948), .A2(n13120), .ZN(n9921) );
  INV_X1 U12385 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n9927) );
  NAND2_X1 U12386 ( .A1(n9923), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n9926) );
  NAND2_X1 U12387 ( .A1(n9924), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9925) );
  OAI211_X1 U12388 ( .C1(n9928), .C2(n9927), .A(n9926), .B(n9925), .ZN(n13912)
         );
  NAND2_X1 U12389 ( .A1(n13912), .A2(n9870), .ZN(n9929) );
  NAND2_X1 U12390 ( .A1(n10018), .A2(n11063), .ZN(n10002) );
  NAND4_X1 U12391 ( .A1(n9929), .A2(n9757), .A3(n10002), .A4(n10683), .ZN(
        n9930) );
  AND2_X1 U12392 ( .A1(n9930), .A2(n13861), .ZN(n9931) );
  AOI21_X1 U12393 ( .B1(n13910), .B2(n10005), .A(n9931), .ZN(n9966) );
  NAND2_X1 U12394 ( .A1(n13910), .A2(n9870), .ZN(n9933) );
  NAND2_X1 U12395 ( .A1(n13861), .A2(n10005), .ZN(n9932) );
  NAND2_X1 U12396 ( .A1(n9933), .A2(n9932), .ZN(n9965) );
  AOI22_X1 U12397 ( .A1(n14106), .A2(n10005), .B1(n13862), .B2(n9870), .ZN(
        n9958) );
  OAI22_X1 U12398 ( .A1(n9934), .A2(n10005), .B1(n13773), .B2(n9908), .ZN(
        n9957) );
  OAI22_X1 U12399 ( .A1(n9966), .A2(n9965), .B1(n9958), .B2(n9957), .ZN(n9954)
         );
  NAND2_X1 U12400 ( .A1(n9936), .A2(n9935), .ZN(n9941) );
  MUX2_X1 U12401 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n9213), .Z(n9937) );
  XNOR2_X1 U12402 ( .A(n9937), .B(n13677), .ZN(n9940) );
  INV_X1 U12403 ( .A(n9940), .ZN(n9938) );
  NOR2_X1 U12404 ( .A1(n9941), .A2(n9938), .ZN(n9947) );
  XNOR2_X1 U12405 ( .A(n9938), .B(n9939), .ZN(n9946) );
  NOR2_X1 U12406 ( .A1(n9941), .A2(n9940), .ZN(n9942) );
  NAND2_X1 U12407 ( .A1(n9943), .A2(n9942), .ZN(n9944) );
  INV_X1 U12408 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n14188) );
  OR2_X1 U12409 ( .A1(n9948), .A2(n14188), .ZN(n9949) );
  INV_X1 U12410 ( .A(n13912), .ZN(n9951) );
  NAND2_X1 U12411 ( .A1(n9952), .A2(n9951), .ZN(n10006) );
  NAND2_X1 U12412 ( .A1(n14101), .A2(n13912), .ZN(n9953) );
  NAND2_X1 U12413 ( .A1(n9954), .A2(n9997), .ZN(n9968) );
  OAI21_X1 U12414 ( .B1(n9961), .B2(n9960), .A(n9968), .ZN(n9955) );
  INV_X1 U12415 ( .A(n9957), .ZN(n9964) );
  INV_X1 U12416 ( .A(n9958), .ZN(n9963) );
  AOI21_X1 U12417 ( .B1(n9961), .B2(n9960), .A(n9959), .ZN(n9962) );
  OAI21_X1 U12418 ( .B1(n9964), .B2(n9963), .A(n9962), .ZN(n9967) );
  AOI22_X1 U12419 ( .A1(n9968), .A2(n9967), .B1(n9966), .B2(n9965), .ZN(n9969)
         );
  NAND2_X1 U12420 ( .A1(n9970), .A2(n9969), .ZN(n10015) );
  XNOR2_X1 U12421 ( .A(n13910), .B(n13861), .ZN(n9996) );
  XNOR2_X1 U12422 ( .A(n11888), .B(n11589), .ZN(n11884) );
  NAND2_X1 U12423 ( .A1(n9974), .A2(n9973), .ZN(n11591) );
  INV_X1 U12424 ( .A(n11287), .ZN(n10000) );
  NAND2_X1 U12425 ( .A1(n10698), .A2(n11474), .ZN(n9975) );
  NAND2_X1 U12426 ( .A1(n9975), .A2(n11466), .ZN(n15291) );
  NAND4_X1 U12427 ( .A1(n6826), .A2(n10000), .A3(n15265), .A4(n15291), .ZN(
        n9977) );
  NOR2_X1 U12428 ( .A1(n9977), .A2(n9976), .ZN(n9978) );
  NAND4_X1 U12429 ( .A1(n11290), .A2(n9978), .A3(n10946), .A4(n11144), .ZN(
        n9979) );
  OR3_X1 U12430 ( .A1(n11069), .A2(n11022), .A3(n9979), .ZN(n9980) );
  NOR2_X1 U12431 ( .A1(n11562), .A2(n9980), .ZN(n9981) );
  NAND4_X1 U12432 ( .A1(n11591), .A2(n9981), .A3(n11643), .A4(n11171), .ZN(
        n9982) );
  OR4_X1 U12433 ( .A1(n12063), .A2(n14985), .A3(n11884), .A4(n9982), .ZN(n9983) );
  NOR2_X1 U12434 ( .A1(n14969), .A2(n9983), .ZN(n9985) );
  NAND3_X1 U12435 ( .A1(n14082), .A2(n9985), .A3(n9984), .ZN(n9986) );
  NOR2_X1 U12436 ( .A1(n14054), .A2(n9986), .ZN(n9987) );
  NAND4_X1 U12437 ( .A1(n14015), .A2(n9987), .A3(n14073), .A4(n14041), .ZN(
        n9988) );
  NOR2_X1 U12438 ( .A1(n9989), .A2(n9988), .ZN(n9990) );
  NAND4_X1 U12439 ( .A1(n13959), .A2(n9990), .A3(n13971), .A4(n7408), .ZN(
        n9992) );
  OR2_X1 U12440 ( .A1(n9992), .A2(n9991), .ZN(n9993) );
  NOR2_X1 U12441 ( .A1(n13923), .A2(n9993), .ZN(n9994) );
  NAND2_X1 U12442 ( .A1(n7640), .A2(n9997), .ZN(n9998) );
  XNOR2_X1 U12443 ( .A(n9998), .B(n9709), .ZN(n9999) );
  NAND2_X1 U12444 ( .A1(n9999), .A2(n9664), .ZN(n10004) );
  NAND3_X1 U12445 ( .A1(n9757), .A2(n10000), .A3(n9709), .ZN(n10001) );
  AND2_X1 U12446 ( .A1(n10002), .A2(n10001), .ZN(n10003) );
  INV_X1 U12447 ( .A(n10723), .ZN(n10008) );
  OAI21_X1 U12448 ( .B1(n9664), .B2(n9709), .A(n10683), .ZN(n10007) );
  NOR2_X1 U12449 ( .A1(n10006), .A2(n10005), .ZN(n10011) );
  AOI211_X1 U12450 ( .C1(n10008), .C2(n11556), .A(n10007), .B(n10011), .ZN(
        n10009) );
  INV_X1 U12451 ( .A(n10063), .ZN(n10020) );
  NAND2_X1 U12452 ( .A1(n10020), .A2(P2_STATE_REG_SCAN_IN), .ZN(n11816) );
  INV_X1 U12453 ( .A(n9668), .ZN(n10071) );
  INV_X1 U12454 ( .A(n10683), .ZN(n10693) );
  NAND4_X1 U12455 ( .A1(n15289), .A2(n10071), .A3(n10693), .A4(n13851), .ZN(
        n10017) );
  OAI211_X1 U12456 ( .C1(n10018), .C2(n11816), .A(n10017), .B(P2_B_REG_SCAN_IN), .ZN(n10019) );
  NOR2_X1 U12457 ( .A1(n10021), .A2(n10020), .ZN(n10065) );
  NOR2_X2 U12458 ( .A1(P1_IR_REG_7__SCAN_IN), .A2(P1_IR_REG_11__SCAN_IN), .ZN(
        n10758) );
  NOR2_X1 U12459 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_18__SCAN_IN), 
        .ZN(n10023) );
  NAND2_X1 U12460 ( .A1(n10234), .A2(n10024), .ZN(n10760) );
  NAND3_X1 U12461 ( .A1(n10137), .A2(n10027), .A3(n10140), .ZN(n10028) );
  NOR2_X2 U12462 ( .A1(n10215), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n10042) );
  NAND2_X1 U12463 ( .A1(n10042), .A2(n10044), .ZN(n10032) );
  INV_X1 U12464 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10033) );
  XNOR2_X1 U12465 ( .A(n10034), .B(n10033), .ZN(n10222) );
  NOR2_X1 U12466 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_24__SCAN_IN), 
        .ZN(n10036) );
  NAND4_X1 U12467 ( .A1(n10036), .A2(n7375), .A3(n10212), .A4(n10035), .ZN(
        n10037) );
  NAND2_X1 U12468 ( .A1(n6773), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10038) );
  MUX2_X1 U12469 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10038), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n10040) );
  NAND2_X1 U12470 ( .A1(n10040), .A2(n10209), .ZN(n12385) );
  OR2_X2 U12471 ( .A1(n10222), .A2(n12385), .ZN(n10041) );
  INV_X1 U12472 ( .A(n10042), .ZN(n10043) );
  NAND2_X1 U12473 ( .A1(n10043), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10045) );
  XNOR2_X1 U12474 ( .A(n10045), .B(n10044), .ZN(n10522) );
  INV_X1 U12475 ( .A(n10228), .ZN(n10046) );
  INV_X1 U12476 ( .A(n12337), .ZN(n12344) );
  AOI22_X1 U12477 ( .A1(n12337), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n12286), 
        .B2(n12344), .ZN(n10061) );
  INV_X1 U12478 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10059) );
  INV_X1 U12479 ( .A(n11958), .ZN(n10870) );
  AOI22_X1 U12480 ( .A1(n11958), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n10059), 
        .B2(n10870), .ZN(n11952) );
  INV_X1 U12481 ( .A(n10101), .ZN(n10864) );
  INV_X1 U12482 ( .A(n10090), .ZN(n15211) );
  INV_X1 U12483 ( .A(n10389), .ZN(n10048) );
  INV_X1 U12484 ( .A(n15185), .ZN(n10076) );
  XNOR2_X1 U12485 ( .A(n10076), .B(P2_REG2_REG_1__SCAN_IN), .ZN(n15188) );
  NOR3_X1 U12486 ( .A1(n15188), .A2(n15189), .A3(n10047), .ZN(n15187) );
  AOI21_X1 U12487 ( .B1(n10076), .B2(P2_REG2_REG_1__SCAN_IN), .A(n15187), .ZN(
        n10380) );
  MUX2_X1 U12488 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n9114), .S(n10389), .Z(
        n10379) );
  NOR2_X1 U12489 ( .A1(n10380), .A2(n10379), .ZN(n10378) );
  AOI21_X1 U12490 ( .B1(P2_REG2_REG_2__SCAN_IN), .B2(n10048), .A(n10378), .ZN(
        n15204) );
  INV_X1 U12491 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n10049) );
  MUX2_X1 U12492 ( .A(n10049), .B(P2_REG2_REG_3__SCAN_IN), .S(n10184), .Z(
        n15203) );
  OR2_X1 U12493 ( .A1(n15204), .A2(n15203), .ZN(n15206) );
  NAND2_X1 U12494 ( .A1(n10184), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n10309) );
  MUX2_X1 U12495 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n11124), .S(n10314), .Z(
        n10308) );
  AOI21_X1 U12496 ( .B1(n15206), .B2(n10309), .A(n10308), .ZN(n10307) );
  NOR2_X1 U12497 ( .A1(n10314), .A2(n11124), .ZN(n10295) );
  MUX2_X1 U12498 ( .A(n11149), .B(P2_REG2_REG_5__SCAN_IN), .S(n10300), .Z(
        n10294) );
  OAI21_X1 U12499 ( .B1(n10307), .B2(n10295), .A(n10294), .ZN(n10297) );
  OAI21_X1 U12500 ( .B1(n11149), .B2(n10300), .A(n10297), .ZN(n15216) );
  MUX2_X1 U12501 ( .A(P2_REG2_REG_6__SCAN_IN), .B(n11128), .S(n10090), .Z(
        n15215) );
  NAND2_X1 U12502 ( .A1(n15216), .A2(n15215), .ZN(n15214) );
  OAI21_X1 U12503 ( .B1(n11128), .B2(n15211), .A(n15214), .ZN(n15232) );
  INV_X1 U12504 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n10050) );
  MUX2_X1 U12505 ( .A(n10050), .B(P2_REG2_REG_7__SCAN_IN), .S(n10196), .Z(
        n10051) );
  INV_X1 U12506 ( .A(n10051), .ZN(n15231) );
  NAND2_X1 U12507 ( .A1(n15232), .A2(n15231), .ZN(n15230) );
  NAND2_X1 U12508 ( .A1(n10196), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n10263) );
  MUX2_X1 U12509 ( .A(n9241), .B(P2_REG2_REG_8__SCAN_IN), .S(n10267), .Z(
        n10262) );
  AOI21_X1 U12510 ( .B1(n15230), .B2(n10263), .A(n10262), .ZN(n10275) );
  AOI21_X1 U12511 ( .B1(P2_REG2_REG_8__SCAN_IN), .B2(n10267), .A(n10275), .ZN(
        n10453) );
  INV_X1 U12512 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n10446) );
  MUX2_X1 U12513 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n10446), .S(n10455), .Z(
        n10052) );
  NAND2_X1 U12514 ( .A1(n10453), .A2(n10052), .ZN(n10451) );
  INV_X1 U12515 ( .A(n10455), .ZN(n10190) );
  NAND2_X1 U12516 ( .A1(n10190), .A2(n10446), .ZN(n10452) );
  NAND2_X1 U12517 ( .A1(n10451), .A2(n10452), .ZN(n10843) );
  INV_X1 U12518 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10053) );
  MUX2_X1 U12519 ( .A(n10053), .B(P2_REG2_REG_10__SCAN_IN), .S(n10199), .Z(
        n10844) );
  NOR2_X1 U12520 ( .A1(n10843), .A2(n10844), .ZN(n10842) );
  AOI21_X1 U12521 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n10199), .A(n10842), 
        .ZN(n10798) );
  INV_X1 U12522 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n11655) );
  MUX2_X1 U12523 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n11655), .S(n10100), .Z(
        n10797) );
  NAND2_X1 U12524 ( .A1(n10798), .A2(n10797), .ZN(n10857) );
  INV_X1 U12525 ( .A(n10100), .ZN(n10800) );
  NAND2_X1 U12526 ( .A1(n10800), .A2(n11655), .ZN(n10855) );
  MUX2_X1 U12527 ( .A(n11596), .B(P2_REG2_REG_12__SCAN_IN), .S(n10101), .Z(
        n10856) );
  AOI21_X1 U12528 ( .B1(n10857), .B2(n10855), .A(n10856), .ZN(n10859) );
  AOI21_X1 U12529 ( .B1(n11596), .B2(n10864), .A(n10859), .ZN(n15241) );
  MUX2_X1 U12530 ( .A(n10054), .B(P2_REG2_REG_13__SCAN_IN), .S(n10279), .Z(
        n15240) );
  NAND2_X1 U12531 ( .A1(n15241), .A2(n15240), .ZN(n15239) );
  OAI21_X1 U12532 ( .B1(n10054), .B2(n10279), .A(n15239), .ZN(n10055) );
  NAND2_X1 U12533 ( .A1(n15258), .A2(n10055), .ZN(n10056) );
  INV_X1 U12534 ( .A(n15258), .ZN(n10537) );
  XNOR2_X1 U12535 ( .A(n10537), .B(n10055), .ZN(n15253) );
  NAND2_X1 U12536 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n15253), .ZN(n15251) );
  NAND2_X1 U12537 ( .A1(n10056), .A2(n15251), .ZN(n10057) );
  NAND2_X1 U12538 ( .A1(n10764), .A2(n10057), .ZN(n10058) );
  XOR2_X1 U12539 ( .A(n10764), .B(n10057), .Z(n11806) );
  NAND2_X1 U12540 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n11806), .ZN(n11805) );
  NAND2_X1 U12541 ( .A1(n10058), .A2(n11805), .ZN(n11951) );
  NAND2_X1 U12542 ( .A1(n11952), .A2(n11951), .ZN(n11950) );
  OAI21_X1 U12543 ( .B1(n10059), .B2(n10870), .A(n11950), .ZN(n10060) );
  NAND2_X1 U12544 ( .A1(n10061), .A2(n10060), .ZN(n12338) );
  OAI21_X1 U12545 ( .B1(n10061), .B2(n10060), .A(n12338), .ZN(n10069) );
  AOI21_X1 U12546 ( .B1(n10063), .B2(n10692), .A(n10062), .ZN(n10064) );
  OR2_X1 U12547 ( .A1(n10065), .A2(n10064), .ZN(n10110) );
  NAND2_X1 U12548 ( .A1(n10066), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14198) );
  INV_X1 U12549 ( .A(n14198), .ZN(n10067) );
  NAND2_X1 U12550 ( .A1(n10110), .A2(n10067), .ZN(n10072) );
  INV_X1 U12551 ( .A(n10072), .ZN(n10068) );
  NOR2_X1 U12552 ( .A1(n10069), .A2(n12354), .ZN(n10115) );
  NAND2_X1 U12553 ( .A1(n10110), .A2(n10070), .ZN(n15212) );
  OR2_X1 U12554 ( .A1(n15212), .A2(P2_U3088), .ZN(n15225) );
  NOR2_X1 U12555 ( .A1(n15225), .A2(n12344), .ZN(n10114) );
  NAND2_X1 U12556 ( .A1(n11958), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n10106) );
  MUX2_X1 U12557 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n10073), .S(n11958), .Z(
        n11954) );
  INV_X1 U12558 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n15019) );
  MUX2_X1 U12559 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n15019), .S(n15258), .Z(
        n15256) );
  MUX2_X1 U12560 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n10074), .S(n10184), .Z(
        n15201) );
  MUX2_X1 U12561 ( .A(n10079), .B(P2_REG1_REG_2__SCAN_IN), .S(n10389), .Z(
        n10078) );
  MUX2_X1 U12562 ( .A(n10075), .B(P2_REG1_REG_1__SCAN_IN), .S(n15185), .Z(
        n15193) );
  AND2_X1 U12563 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .ZN(n15194) );
  NAND2_X1 U12564 ( .A1(n15193), .A2(n15194), .ZN(n15192) );
  NAND2_X1 U12565 ( .A1(n10076), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n10384) );
  NAND2_X1 U12566 ( .A1(n15192), .A2(n10384), .ZN(n10077) );
  NAND2_X1 U12567 ( .A1(n10078), .A2(n10077), .ZN(n10386) );
  OR2_X1 U12568 ( .A1(n10389), .A2(n10079), .ZN(n10080) );
  NAND2_X1 U12569 ( .A1(n10386), .A2(n10080), .ZN(n15202) );
  NAND2_X1 U12570 ( .A1(n15201), .A2(n15202), .ZN(n15200) );
  NAND2_X1 U12571 ( .A1(n10184), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n10302) );
  NAND2_X1 U12572 ( .A1(n15200), .A2(n10302), .ZN(n10082) );
  MUX2_X1 U12573 ( .A(n10083), .B(P2_REG1_REG_4__SCAN_IN), .S(n10314), .Z(
        n10081) );
  NAND2_X1 U12574 ( .A1(n10082), .A2(n10081), .ZN(n10304) );
  OR2_X1 U12575 ( .A1(n10314), .A2(n10083), .ZN(n10288) );
  NAND2_X1 U12576 ( .A1(n10304), .A2(n10288), .ZN(n10086) );
  MUX2_X1 U12577 ( .A(n10084), .B(P2_REG1_REG_5__SCAN_IN), .S(n10300), .Z(
        n10085) );
  NAND2_X1 U12578 ( .A1(n10086), .A2(n10085), .ZN(n10291) );
  NAND2_X1 U12579 ( .A1(n10087), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n10088) );
  NAND2_X1 U12580 ( .A1(n10291), .A2(n10088), .ZN(n15219) );
  MUX2_X1 U12581 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n10089), .S(n10090), .Z(
        n15218) );
  NAND2_X1 U12582 ( .A1(n15219), .A2(n15218), .ZN(n15217) );
  NAND2_X1 U12583 ( .A1(n10090), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n10091) );
  NAND2_X1 U12584 ( .A1(n15217), .A2(n10091), .ZN(n15235) );
  MUX2_X1 U12585 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n10092), .S(n10196), .Z(
        n15234) );
  NAND2_X1 U12586 ( .A1(n15235), .A2(n15234), .ZN(n15233) );
  NAND2_X1 U12587 ( .A1(n10196), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n10269) );
  NAND2_X1 U12588 ( .A1(n15233), .A2(n10269), .ZN(n10095) );
  MUX2_X1 U12589 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n10093), .S(n10267), .Z(
        n10094) );
  NAND2_X1 U12590 ( .A1(n10095), .A2(n10094), .ZN(n10271) );
  NAND2_X1 U12591 ( .A1(n10267), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n10096) );
  NAND2_X1 U12592 ( .A1(n10271), .A2(n10096), .ZN(n10447) );
  MUX2_X1 U12593 ( .A(n10097), .B(P2_REG1_REG_9__SCAN_IN), .S(n10455), .Z(
        n10098) );
  NOR2_X1 U12594 ( .A1(n10447), .A2(n10098), .ZN(n10444) );
  AOI21_X1 U12595 ( .B1(n10097), .B2(n10190), .A(n10444), .ZN(n10848) );
  MUX2_X1 U12596 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n10099), .S(n10199), .Z(
        n10847) );
  NAND2_X1 U12597 ( .A1(n10848), .A2(n10847), .ZN(n10846) );
  NAND2_X1 U12598 ( .A1(n10199), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n10795) );
  MUX2_X1 U12599 ( .A(n9301), .B(P2_REG1_REG_11__SCAN_IN), .S(n10100), .Z(
        n10794) );
  AOI21_X1 U12600 ( .B1(n10846), .B2(n10795), .A(n10794), .ZN(n10805) );
  AOI21_X1 U12601 ( .B1(n10100), .B2(P2_REG1_REG_11__SCAN_IN), .A(n10805), 
        .ZN(n10863) );
  MUX2_X1 U12602 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n9322), .S(n10101), .Z(
        n10862) );
  AND2_X1 U12603 ( .A1(n10863), .A2(n10862), .ZN(n10860) );
  AOI21_X1 U12604 ( .B1(n9322), .B2(n10864), .A(n10860), .ZN(n15245) );
  MUX2_X1 U12605 ( .A(n10102), .B(P2_REG1_REG_13__SCAN_IN), .S(n10279), .Z(
        n15244) );
  NAND2_X1 U12606 ( .A1(n15245), .A2(n15244), .ZN(n15243) );
  OAI21_X1 U12607 ( .B1(n10102), .B2(n10279), .A(n15243), .ZN(n15257) );
  NAND2_X1 U12608 ( .A1(n15256), .A2(n15257), .ZN(n15254) );
  OAI21_X1 U12609 ( .B1(n15019), .B2(n10537), .A(n15254), .ZN(n10103) );
  NAND2_X1 U12610 ( .A1(n10764), .A2(n10103), .ZN(n10105) );
  INV_X1 U12611 ( .A(n10103), .ZN(n10104) );
  XNOR2_X1 U12612 ( .A(n10764), .B(n10104), .ZN(n11808) );
  NAND2_X1 U12613 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n11808), .ZN(n11807) );
  NAND2_X1 U12614 ( .A1(n10105), .A2(n11807), .ZN(n11955) );
  NAND2_X1 U12615 ( .A1(n11954), .A2(n11955), .ZN(n11953) );
  NAND2_X1 U12616 ( .A1(n10106), .A2(n11953), .ZN(n10108) );
  XNOR2_X1 U12617 ( .A(n12337), .B(n12345), .ZN(n10107) );
  NAND2_X1 U12618 ( .A1(n10107), .A2(n10108), .ZN(n12343) );
  OAI21_X1 U12619 ( .B1(n10108), .B2(n10107), .A(n12343), .ZN(n10109) );
  NOR2_X1 U12620 ( .A1(n13901), .A2(n10109), .ZN(n10113) );
  INV_X1 U12621 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n10111) );
  NAND2_X1 U12622 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n13806)
         );
  OAI21_X1 U12623 ( .B1(n15228), .B2(n10111), .A(n13806), .ZN(n10112) );
  OR4_X1 U12624 ( .A1(n10115), .A2(n10114), .A3(n10113), .A4(n10112), .ZN(
        P2_U3231) );
  NAND2_X1 U12625 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n10116) );
  XNOR2_X1 U12626 ( .A(n10117), .B(n10116), .ZN(n14387) );
  NAND2_X1 U12627 ( .A1(n10170), .A2(P1_U3086), .ZN(n11283) );
  AND2_X1 U12628 ( .A1(n9213), .A2(P1_U3086), .ZN(n14866) );
  INV_X2 U12629 ( .A(n14866), .ZN(n14876) );
  OAI222_X1 U12630 ( .A1(P1_U3086), .A2(n14387), .B1(n11283), .B2(n10615), 
        .C1(n6853), .C2(n14876), .ZN(P1_U3354) );
  INV_X1 U12631 ( .A(n10118), .ZN(n11221) );
  NAND2_X1 U12632 ( .A1(n10120), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10122) );
  XNOR2_X1 U12633 ( .A(n10122), .B(n10121), .ZN(n11224) );
  OAI222_X1 U12634 ( .A1(n14876), .A2(n11220), .B1(n11283), .B2(n11221), .C1(
        P1_U3086), .C2(n11224), .ZN(P1_U3351) );
  NOR2_X1 U12635 ( .A1(n9213), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13681) );
  AND2_X1 U12636 ( .A1(n9213), .A2(P3_U3151), .ZN(n10149) );
  AOI222_X1 U12637 ( .A1(n10123), .A2(n13681), .B1(SI_7_), .B2(n10149), .C1(
        n15464), .C2(P3_STATE_REG_SCAN_IN), .ZN(n10124) );
  INV_X1 U12638 ( .A(n10124), .ZN(P3_U3288) );
  AOI222_X1 U12639 ( .A1(n10125), .A2(n13681), .B1(n10594), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_3_), .C2(n10149), .ZN(n10126) );
  INV_X1 U12640 ( .A(n10126), .ZN(P3_U3292) );
  AOI222_X1 U12641 ( .A1(n10127), .A2(n13681), .B1(SI_5_), .B2(n10149), .C1(
        n15434), .C2(P3_STATE_REG_SCAN_IN), .ZN(n10128) );
  INV_X1 U12642 ( .A(n10128), .ZN(P3_U3290) );
  AOI222_X1 U12643 ( .A1(n10130), .A2(n13681), .B1(n10129), .B2(
        P3_STATE_REG_SCAN_IN), .C1(SI_4_), .C2(n10149), .ZN(n10131) );
  INV_X1 U12644 ( .A(n10131), .ZN(P3_U3291) );
  OR2_X1 U12645 ( .A1(n10132), .A2(n14864), .ZN(n10134) );
  XNOR2_X1 U12646 ( .A(n10134), .B(n10133), .ZN(n10825) );
  OAI222_X1 U12647 ( .A1(P1_U3086), .A2(n10825), .B1(n11283), .B2(n9106), .C1(
        n10823), .C2(n14876), .ZN(P1_U3353) );
  INV_X1 U12648 ( .A(n11325), .ZN(n10187) );
  INV_X1 U12649 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14864) );
  MUX2_X1 U12650 ( .A(n14864), .B(n10136), .S(P1_IR_REG_5__SCAN_IN), .Z(n10138) );
  OR2_X1 U12651 ( .A1(n10138), .A2(n10141), .ZN(n11329) );
  OAI222_X1 U12652 ( .A1(n14876), .A2(n11326), .B1(n11283), .B2(n10187), .C1(
        P1_U3086), .C2(n11329), .ZN(P1_U3350) );
  NOR2_X1 U12653 ( .A1(n10141), .A2(n14864), .ZN(n10139) );
  MUX2_X1 U12654 ( .A(n14864), .B(n10139), .S(P1_IR_REG_6__SCAN_IN), .Z(n10143) );
  INV_X1 U12655 ( .A(n10761), .ZN(n10142) );
  OAI222_X1 U12656 ( .A1(n14876), .A2(n10144), .B1(n11283), .B2(n11338), .C1(
        n10400), .C2(P1_U3086), .ZN(P1_U3349) );
  INV_X1 U12657 ( .A(n11283), .ZN(n11819) );
  INV_X1 U12658 ( .A(n11819), .ZN(n14874) );
  INV_X1 U12659 ( .A(n10977), .ZN(n10185) );
  NAND2_X1 U12660 ( .A1(n10145), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10147) );
  XNOR2_X1 U12661 ( .A(n10147), .B(n10146), .ZN(n14402) );
  OAI222_X1 U12662 ( .A1(n14876), .A2(n10979), .B1(n14874), .B2(n10185), .C1(
        P1_U3086), .C2(n14402), .ZN(P1_U3352) );
  INV_X1 U12663 ( .A(n10148), .ZN(n10151) );
  INV_X2 U12664 ( .A(n10149), .ZN(n13690) );
  OAI222_X1 U12665 ( .A1(n13688), .A2(n10151), .B1(n13690), .B2(n10150), .C1(
        n7766), .C2(P3_U3151), .ZN(P3_U3293) );
  INV_X1 U12666 ( .A(n10152), .ZN(n10155) );
  INV_X1 U12667 ( .A(SI_9_), .ZN(n10154) );
  INV_X1 U12668 ( .A(n10153), .ZN(n11054) );
  OAI222_X1 U12669 ( .A1(n13688), .A2(n10155), .B1(n13690), .B2(n10154), .C1(
        n11054), .C2(P3_U3151), .ZN(P3_U3286) );
  OAI222_X1 U12670 ( .A1(n13688), .A2(n10157), .B1(n13690), .B2(n10156), .C1(
        n15483), .C2(P3_U3151), .ZN(P3_U3287) );
  OAI222_X1 U12671 ( .A1(P3_U3151), .A2(n10160), .B1(n13690), .B2(n10159), 
        .C1(n13688), .C2(n10158), .ZN(P3_U3294) );
  OAI222_X1 U12672 ( .A1(n15442), .A2(P3_U3151), .B1(n13688), .B2(n10162), 
        .C1(n10161), .C2(n13690), .ZN(P3_U3289) );
  INV_X1 U12673 ( .A(SI_10_), .ZN(n10164) );
  OAI222_X1 U12674 ( .A1(n13688), .A2(n10165), .B1(n13690), .B2(n10164), .C1(
        n10163), .C2(P3_U3151), .ZN(P3_U3285) );
  INV_X1 U12675 ( .A(n11378), .ZN(n10197) );
  NAND2_X1 U12676 ( .A1(n10761), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10173) );
  XNOR2_X1 U12677 ( .A(n10173), .B(P1_IR_REG_7__SCAN_IN), .ZN(n11379) );
  INV_X1 U12678 ( .A(n11379), .ZN(n10475) );
  OAI222_X1 U12679 ( .A1(n14876), .A2(n10166), .B1(n11283), .B2(n10197), .C1(
        P1_U3086), .C2(n10475), .ZN(P1_U3348) );
  OAI222_X1 U12680 ( .A1(n13688), .A2(n10169), .B1(n10168), .B2(P3_U3151), 
        .C1(n13690), .C2(n10167), .ZN(P3_U3284) );
  NAND2_X2 U12681 ( .A1(n9213), .A2(P2_U3088), .ZN(n14196) );
  OAI222_X1 U12682 ( .A1(n14201), .A2(n10171), .B1(n14196), .B2(n10615), .C1(
        n15185), .C2(P2_U3088), .ZN(P2_U3326) );
  INV_X1 U12683 ( .A(n11683), .ZN(n10194) );
  INV_X1 U12684 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n10172) );
  NAND2_X1 U12685 ( .A1(n10173), .A2(n10172), .ZN(n10174) );
  NAND2_X1 U12686 ( .A1(n10174), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10177) );
  XNOR2_X1 U12687 ( .A(n10177), .B(P1_IR_REG_8__SCAN_IN), .ZN(n11684) );
  INV_X1 U12688 ( .A(n11684), .ZN(n10415) );
  OAI222_X1 U12689 ( .A1(n14876), .A2(n10175), .B1(n14874), .B2(n10194), .C1(
        P1_U3086), .C2(n10415), .ZN(P1_U3347) );
  INV_X1 U12690 ( .A(n11834), .ZN(n10191) );
  INV_X1 U12691 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n10176) );
  NAND2_X1 U12692 ( .A1(n10177), .A2(n10176), .ZN(n10178) );
  XNOR2_X1 U12693 ( .A(n10236), .B(P1_IR_REG_9__SCAN_IN), .ZN(n11835) );
  INV_X1 U12694 ( .A(n11835), .ZN(n10433) );
  OAI222_X1 U12695 ( .A1(n14876), .A2(n10179), .B1(n14874), .B2(n10191), .C1(
        P1_U3086), .C2(n10433), .ZN(P1_U3346) );
  OAI222_X1 U12696 ( .A1(n13688), .A2(n10181), .B1(n15500), .B2(P3_U3151), 
        .C1(n10180), .C2(n13690), .ZN(P3_U3283) );
  OAI222_X1 U12697 ( .A1(n14201), .A2(n10182), .B1(n14196), .B2(n11221), .C1(
        P2_U3088), .C2(n10314), .ZN(P2_U3323) );
  OAI222_X1 U12698 ( .A1(n14201), .A2(n10183), .B1(n14196), .B2(n9106), .C1(
        n10389), .C2(P2_U3088), .ZN(P2_U3325) );
  INV_X1 U12699 ( .A(n10184), .ZN(n15198) );
  OAI222_X1 U12700 ( .A1(n14201), .A2(n10186), .B1(n14196), .B2(n10185), .C1(
        P2_U3088), .C2(n15198), .ZN(P2_U3324) );
  OAI222_X1 U12701 ( .A1(n14201), .A2(n10188), .B1(n14196), .B2(n10187), .C1(
        P2_U3088), .C2(n10300), .ZN(P2_U3322) );
  OAI222_X1 U12702 ( .A1(n14201), .A2(n10189), .B1(n14196), .B2(n11338), .C1(
        n15211), .C2(P2_U3088), .ZN(P2_U3321) );
  OAI222_X1 U12703 ( .A1(n14201), .A2(n10192), .B1(n14196), .B2(n10191), .C1(
        P2_U3088), .C2(n10190), .ZN(P2_U3318) );
  INV_X1 U12704 ( .A(n10267), .ZN(n10193) );
  OAI222_X1 U12705 ( .A1(n14201), .A2(n10195), .B1(n14196), .B2(n10194), .C1(
        P2_U3088), .C2(n10193), .ZN(P2_U3319) );
  INV_X1 U12706 ( .A(n10196), .ZN(n15224) );
  OAI222_X1 U12707 ( .A1(n14201), .A2(n10198), .B1(n14196), .B2(n10197), .C1(
        P2_U3088), .C2(n15224), .ZN(P2_U3320) );
  INV_X1 U12708 ( .A(n11973), .ZN(n10204) );
  INV_X1 U12709 ( .A(n10199), .ZN(n10854) );
  OAI222_X1 U12710 ( .A1(n14201), .A2(n10200), .B1(n14196), .B2(n10204), .C1(
        P2_U3088), .C2(n10854), .ZN(P2_U3317) );
  NAND2_X1 U12711 ( .A1(n10236), .A2(n10201), .ZN(n10202) );
  NAND2_X1 U12712 ( .A1(n10202), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10203) );
  XNOR2_X1 U12713 ( .A(n10203), .B(P1_IR_REG_10__SCAN_IN), .ZN(n14418) );
  INV_X1 U12714 ( .A(n14418), .ZN(n10428) );
  OAI222_X1 U12715 ( .A1(n14876), .A2(n10205), .B1(n14874), .B2(n10204), .C1(
        P1_U3086), .C2(n10428), .ZN(P1_U3345) );
  INV_X1 U12716 ( .A(n12880), .ZN(n10206) );
  OR2_X1 U12717 ( .A1(n10522), .A2(P1_U3086), .ZN(n12883) );
  NAND2_X1 U12718 ( .A1(n10206), .A2(n12883), .ZN(n10246) );
  NAND2_X1 U12719 ( .A1(n10215), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10213) );
  NAND2_X1 U12720 ( .A1(n10489), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10214) );
  MUX2_X1 U12721 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10214), .S(
        P1_IR_REG_21__SCAN_IN), .Z(n10216) );
  NAND2_X1 U12722 ( .A1(n10216), .A2(n10215), .ZN(n12486) );
  NAND2_X1 U12723 ( .A1(n10522), .A2(n12484), .ZN(n10217) );
  NAND2_X1 U12724 ( .A1(n12738), .A2(n10217), .ZN(n10244) );
  NOR2_X1 U12725 ( .A1(n14435), .A2(n14379), .ZN(P1_U3085) );
  INV_X1 U12726 ( .A(n10218), .ZN(n10241) );
  INV_X1 U12727 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n10221) );
  NAND2_X1 U12728 ( .A1(n10219), .A2(n10241), .ZN(n10220) );
  OAI21_X1 U12729 ( .B1(n10241), .B2(n10221), .A(n10220), .ZN(P3_U3376) );
  NAND2_X1 U12730 ( .A1(n12324), .A2(P1_B_REG_SCAN_IN), .ZN(n10223) );
  MUX2_X1 U12731 ( .A(P1_B_REG_SCAN_IN), .B(n10223), .S(n10222), .Z(n10225) );
  INV_X1 U12732 ( .A(n12385), .ZN(n10224) );
  NAND2_X1 U12733 ( .A1(n10512), .A2(n12880), .ZN(n15153) );
  INV_X1 U12734 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n10227) );
  NAND2_X1 U12735 ( .A1(n12324), .A2(n12385), .ZN(n10497) );
  INV_X1 U12736 ( .A(n10497), .ZN(n10226) );
  AOI22_X1 U12737 ( .A1(n15153), .A2(n10227), .B1(n10226), .B2(n10228), .ZN(
        P1_U3446) );
  INV_X1 U12738 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10230) );
  NAND2_X1 U12739 ( .A1(n10222), .A2(n12385), .ZN(n10499) );
  INV_X1 U12740 ( .A(n10499), .ZN(n10229) );
  AOI22_X1 U12741 ( .A1(n15153), .A2(n10230), .B1(n10229), .B2(n10228), .ZN(
        P1_U3445) );
  INV_X1 U12742 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n10232) );
  NAND2_X1 U12743 ( .A1(n11006), .A2(n10241), .ZN(n10231) );
  OAI21_X1 U12744 ( .B1(n10241), .B2(n10232), .A(n10231), .ZN(P3_U3377) );
  INV_X1 U12745 ( .A(n12089), .ZN(n10238) );
  OAI222_X1 U12746 ( .A1(n14201), .A2(n10233), .B1(n14196), .B2(n10238), .C1(
        P2_U3088), .C2(n10800), .ZN(P2_U3316) );
  OR2_X1 U12747 ( .A1(n10234), .A2(n14864), .ZN(n10235) );
  NAND2_X1 U12748 ( .A1(n10236), .A2(n10235), .ZN(n10256) );
  INV_X1 U12749 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n10237) );
  XNOR2_X1 U12750 ( .A(n10256), .B(n10237), .ZN(n12090) );
  INV_X1 U12751 ( .A(n12090), .ZN(n10239) );
  OAI222_X1 U12752 ( .A1(n10240), .A2(n14876), .B1(P1_U3086), .B2(n10239), 
        .C1(n14874), .C2(n10238), .ZN(P1_U3344) );
  AND2_X1 U12753 ( .A1(n10243), .A2(P3_D_REG_10__SCAN_IN), .ZN(P3_U3255) );
  AND2_X1 U12754 ( .A1(n10243), .A2(P3_D_REG_11__SCAN_IN), .ZN(P3_U3254) );
  AND2_X1 U12755 ( .A1(n10243), .A2(P3_D_REG_13__SCAN_IN), .ZN(P3_U3252) );
  AND2_X1 U12756 ( .A1(n10243), .A2(P3_D_REG_14__SCAN_IN), .ZN(P3_U3251) );
  AND2_X1 U12757 ( .A1(n10243), .A2(P3_D_REG_12__SCAN_IN), .ZN(P3_U3253) );
  AND2_X1 U12758 ( .A1(n10243), .A2(P3_D_REG_9__SCAN_IN), .ZN(P3_U3256) );
  AND2_X1 U12759 ( .A1(n10243), .A2(P3_D_REG_17__SCAN_IN), .ZN(P3_U3248) );
  AND2_X1 U12760 ( .A1(n10243), .A2(P3_D_REG_18__SCAN_IN), .ZN(P3_U3247) );
  AND2_X1 U12761 ( .A1(n10243), .A2(P3_D_REG_26__SCAN_IN), .ZN(P3_U3239) );
  AND2_X1 U12762 ( .A1(n10243), .A2(P3_D_REG_27__SCAN_IN), .ZN(P3_U3238) );
  AND2_X1 U12763 ( .A1(n10243), .A2(P3_D_REG_28__SCAN_IN), .ZN(P3_U3237) );
  AND2_X1 U12764 ( .A1(n10243), .A2(P3_D_REG_8__SCAN_IN), .ZN(P3_U3257) );
  AND2_X1 U12765 ( .A1(n10243), .A2(P3_D_REG_30__SCAN_IN), .ZN(P3_U3235) );
  AND2_X1 U12766 ( .A1(n10243), .A2(P3_D_REG_24__SCAN_IN), .ZN(P3_U3241) );
  AND2_X1 U12767 ( .A1(n10243), .A2(P3_D_REG_25__SCAN_IN), .ZN(P3_U3240) );
  AND2_X1 U12768 ( .A1(n10243), .A2(P3_D_REG_16__SCAN_IN), .ZN(P3_U3249) );
  AND2_X1 U12769 ( .A1(n10243), .A2(P3_D_REG_20__SCAN_IN), .ZN(P3_U3245) );
  AND2_X1 U12770 ( .A1(n10243), .A2(P3_D_REG_4__SCAN_IN), .ZN(P3_U3261) );
  AND2_X1 U12771 ( .A1(n10243), .A2(P3_D_REG_29__SCAN_IN), .ZN(P3_U3236) );
  AND2_X1 U12772 ( .A1(n10243), .A2(P3_D_REG_3__SCAN_IN), .ZN(P3_U3262) );
  AND2_X1 U12773 ( .A1(n10243), .A2(P3_D_REG_31__SCAN_IN), .ZN(P3_U3234) );
  AND2_X1 U12774 ( .A1(n10243), .A2(P3_D_REG_15__SCAN_IN), .ZN(P3_U3250) );
  AND2_X1 U12775 ( .A1(n10243), .A2(P3_D_REG_2__SCAN_IN), .ZN(P3_U3263) );
  AND2_X1 U12776 ( .A1(n10243), .A2(P3_D_REG_6__SCAN_IN), .ZN(P3_U3259) );
  AND2_X1 U12777 ( .A1(n10243), .A2(P3_D_REG_7__SCAN_IN), .ZN(P3_U3258) );
  AND2_X1 U12778 ( .A1(n10243), .A2(P3_D_REG_5__SCAN_IN), .ZN(P3_U3260) );
  AND2_X1 U12779 ( .A1(n10243), .A2(P3_D_REG_23__SCAN_IN), .ZN(P3_U3242) );
  AND2_X1 U12780 ( .A1(n10243), .A2(P3_D_REG_22__SCAN_IN), .ZN(P3_U3243) );
  AND2_X1 U12781 ( .A1(n10243), .A2(P3_D_REG_19__SCAN_IN), .ZN(P3_U3246) );
  AND2_X1 U12782 ( .A1(n10243), .A2(P3_D_REG_21__SCAN_IN), .ZN(P3_U3244) );
  INV_X1 U12783 ( .A(n14435), .ZN(n15128) );
  INV_X1 U12784 ( .A(n10244), .ZN(n10245) );
  NAND2_X1 U12785 ( .A1(n10246), .A2(n10245), .ZN(n10318) );
  INV_X1 U12786 ( .A(n10318), .ZN(n10329) );
  INV_X1 U12787 ( .A(n14872), .ZN(n13102) );
  INV_X1 U12788 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10249) );
  AOI21_X1 U12789 ( .B1(n13102), .B2(n10249), .A(n10248), .ZN(n10644) );
  OAI21_X1 U12790 ( .B1(n13102), .B2(P1_REG1_REG_0__SCAN_IN), .A(n10644), .ZN(
        n10250) );
  XNOR2_X1 U12791 ( .A(n10250), .B(P1_IR_REG_0__SCAN_IN), .ZN(n10251) );
  AOI22_X1 U12792 ( .A1(n10329), .A2(n10251), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10252) );
  OAI21_X1 U12793 ( .B1(n15128), .B2(n7014), .A(n10252), .ZN(P1_U3243) );
  OAI222_X1 U12794 ( .A1(n13688), .A2(n10255), .B1(n13690), .B2(n10254), .C1(
        n10253), .C2(P3_U3151), .ZN(P3_U3282) );
  INV_X1 U12795 ( .A(n12167), .ZN(n10260) );
  NAND2_X1 U12796 ( .A1(n10257), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10281) );
  XNOR2_X1 U12797 ( .A(n10281), .B(P1_IR_REG_12__SCAN_IN), .ZN(n14440) );
  INV_X1 U12798 ( .A(n14440), .ZN(n10258) );
  OAI222_X1 U12799 ( .A1(n14876), .A2(n10259), .B1(n11283), .B2(n10260), .C1(
        n10258), .C2(P1_U3086), .ZN(P1_U3343) );
  OAI222_X1 U12800 ( .A1(n14201), .A2(n10261), .B1(n14196), .B2(n10260), .C1(
        n10864), .C2(P2_U3088), .ZN(P2_U3315) );
  NAND3_X1 U12801 ( .A1(n15230), .A2(n10263), .A3(n10262), .ZN(n10264) );
  NAND2_X1 U12802 ( .A1(n10264), .A2(n15252), .ZN(n10274) );
  INV_X1 U12803 ( .A(n15225), .ZN(n15259) );
  INV_X1 U12804 ( .A(P2_ADDR_REG_8__SCAN_IN), .ZN(n10265) );
  NAND2_X1 U12805 ( .A1(P2_U3088), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n11211) );
  OAI21_X1 U12806 ( .B1(n15228), .B2(n10265), .A(n11211), .ZN(n10266) );
  AOI21_X1 U12807 ( .B1(n10267), .B2(n15259), .A(n10266), .ZN(n10273) );
  MUX2_X1 U12808 ( .A(n10093), .B(P2_REG1_REG_8__SCAN_IN), .S(n10267), .Z(
        n10268) );
  NAND3_X1 U12809 ( .A1(n15233), .A2(n10269), .A3(n10268), .ZN(n10270) );
  NAND3_X1 U12810 ( .A1(n15255), .A2(n10271), .A3(n10270), .ZN(n10272) );
  OAI211_X1 U12811 ( .C1(n10275), .C2(n10274), .A(n10273), .B(n10272), .ZN(
        P2_U3222) );
  OAI222_X1 U12812 ( .A1(n13688), .A2(n10277), .B1(n13690), .B2(n10276), .C1(
        n15519), .C2(P3_U3151), .ZN(P3_U3281) );
  INV_X1 U12813 ( .A(n12239), .ZN(n10286) );
  OAI222_X1 U12814 ( .A1(P2_U3088), .A2(n10279), .B1(n14196), .B2(n10286), 
        .C1(n10278), .C2(n14201), .ZN(P2_U3314) );
  NAND2_X1 U12815 ( .A1(n10281), .A2(n10280), .ZN(n10282) );
  NAND2_X1 U12816 ( .A1(n10282), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10284) );
  INV_X1 U12817 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n10283) );
  NAND2_X1 U12818 ( .A1(n10284), .A2(n10283), .ZN(n10534) );
  OR2_X1 U12819 ( .A1(n10284), .A2(n10283), .ZN(n10285) );
  INV_X1 U12820 ( .A(n12240), .ZN(n11725) );
  OAI222_X1 U12821 ( .A1(n14876), .A2(n10287), .B1(n11283), .B2(n10286), .C1(
        n11725), .C2(P1_U3086), .ZN(P1_U3342) );
  INV_X1 U12822 ( .A(n15228), .ZN(n15250) );
  NAND2_X1 U12823 ( .A1(P2_U3088), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10790) );
  INV_X1 U12824 ( .A(n10790), .ZN(n10293) );
  MUX2_X1 U12825 ( .A(P2_REG1_REG_5__SCAN_IN), .B(n10084), .S(n10300), .Z(
        n10289) );
  NAND3_X1 U12826 ( .A1(n10289), .A2(n10304), .A3(n10288), .ZN(n10290) );
  AND3_X1 U12827 ( .A1(n15255), .A2(n10291), .A3(n10290), .ZN(n10292) );
  AOI211_X1 U12828 ( .C1(n15250), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n10293), .B(
        n10292), .ZN(n10299) );
  OR3_X1 U12829 ( .A1(n10307), .A2(n10295), .A3(n10294), .ZN(n10296) );
  NAND3_X1 U12830 ( .A1(n15252), .A2(n10297), .A3(n10296), .ZN(n10298) );
  OAI211_X1 U12831 ( .C1(n15225), .C2(n10300), .A(n10299), .B(n10298), .ZN(
        P2_U3219) );
  NAND2_X1 U12832 ( .A1(P2_U3088), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n10749) );
  INV_X1 U12833 ( .A(n10749), .ZN(n10306) );
  MUX2_X1 U12834 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n10083), .S(n10314), .Z(
        n10301) );
  NAND3_X1 U12835 ( .A1(n15200), .A2(n10302), .A3(n10301), .ZN(n10303) );
  AND3_X1 U12836 ( .A1(n15255), .A2(n10304), .A3(n10303), .ZN(n10305) );
  AOI211_X1 U12837 ( .C1(n15250), .C2(P2_ADDR_REG_4__SCAN_IN), .A(n10306), .B(
        n10305), .ZN(n10313) );
  INV_X1 U12838 ( .A(n10307), .ZN(n10311) );
  NAND3_X1 U12839 ( .A1(n15206), .A2(n10309), .A3(n10308), .ZN(n10310) );
  NAND3_X1 U12840 ( .A1(n15252), .A2(n10311), .A3(n10310), .ZN(n10312) );
  OAI211_X1 U12841 ( .C1(n15225), .C2(n10314), .A(n10313), .B(n10312), .ZN(
        P2_U3218) );
  OAI222_X1 U12842 ( .A1(n13688), .A2(n10317), .B1(n13690), .B2(n10316), .C1(
        n10315), .C2(P3_U3151), .ZN(P3_U3280) );
  INV_X1 U12843 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n11509) );
  MUX2_X1 U12844 ( .A(n11509), .B(P1_REG1_REG_5__SCAN_IN), .S(n11329), .Z(
        n10324) );
  INV_X1 U12845 ( .A(n11224), .ZN(n10672) );
  INV_X1 U12846 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n10632) );
  MUX2_X1 U12847 ( .A(n10632), .B(P1_REG1_REG_2__SCAN_IN), .S(n10825), .Z(
        n10320) );
  INV_X1 U12848 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10518) );
  MUX2_X1 U12849 ( .A(n10518), .B(P1_REG1_REG_1__SCAN_IN), .S(n14387), .Z(
        n14382) );
  AND2_X1 U12850 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n14383) );
  OR2_X1 U12851 ( .A1(n14387), .A2(n10518), .ZN(n10649) );
  NAND2_X1 U12852 ( .A1(n14381), .A2(n10649), .ZN(n10319) );
  NAND2_X1 U12853 ( .A1(n10320), .A2(n10319), .ZN(n14399) );
  INV_X1 U12854 ( .A(n14399), .ZN(n10322) );
  NOR2_X1 U12855 ( .A1(n10825), .A2(n10632), .ZN(n14396) );
  INV_X1 U12856 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n10833) );
  MUX2_X1 U12857 ( .A(n10833), .B(P1_REG1_REG_3__SCAN_IN), .S(n14402), .Z(
        n10321) );
  INV_X1 U12858 ( .A(n14402), .ZN(n14395) );
  NAND2_X1 U12859 ( .A1(n14395), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n10659) );
  INV_X1 U12860 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n11485) );
  MUX2_X1 U12861 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n11485), .S(n11224), .Z(
        n10658) );
  AOI21_X1 U12862 ( .B1(n14401), .B2(n10659), .A(n10658), .ZN(n10661) );
  NAND2_X1 U12863 ( .A1(n10323), .A2(n10324), .ZN(n10351) );
  OAI21_X1 U12864 ( .B1(n10324), .B2(n10323), .A(n10351), .ZN(n10341) );
  AND2_X1 U12865 ( .A1(n10329), .A2(n10248), .ZN(n14480) );
  INV_X1 U12866 ( .A(n11329), .ZN(n10354) );
  NAND2_X1 U12867 ( .A1(n14480), .A2(n10354), .ZN(n10326) );
  NAND2_X1 U12868 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n10325) );
  OAI211_X1 U12869 ( .C1(n10327), .C2(n15128), .A(n10326), .B(n10325), .ZN(
        n10340) );
  NOR2_X1 U12870 ( .A1(n10248), .A2(n14872), .ZN(n10328) );
  AND2_X1 U12871 ( .A1(n10329), .A2(n10328), .ZN(n14482) );
  INV_X1 U12872 ( .A(n14482), .ZN(n15121) );
  INV_X1 U12873 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n10645) );
  MUX2_X1 U12874 ( .A(n10645), .B(P1_REG2_REG_2__SCAN_IN), .S(n10825), .Z(
        n10331) );
  INV_X1 U12875 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n11637) );
  MUX2_X1 U12876 ( .A(n11637), .B(P1_REG2_REG_1__SCAN_IN), .S(n14387), .Z(
        n14385) );
  AND2_X1 U12877 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n14386) );
  NAND2_X1 U12878 ( .A1(n14385), .A2(n14386), .ZN(n14384) );
  OR2_X1 U12879 ( .A1(n14387), .A2(n11637), .ZN(n10646) );
  NAND2_X1 U12880 ( .A1(n14384), .A2(n10646), .ZN(n10330) );
  NAND2_X1 U12881 ( .A1(n10331), .A2(n10330), .ZN(n14405) );
  INV_X1 U12882 ( .A(n10825), .ZN(n10652) );
  NAND2_X1 U12883 ( .A1(n10652), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n14403) );
  NAND2_X1 U12884 ( .A1(n14405), .A2(n14403), .ZN(n10334) );
  INV_X1 U12885 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n10332) );
  MUX2_X1 U12886 ( .A(n10332), .B(P1_REG2_REG_3__SCAN_IN), .S(n14402), .Z(
        n10333) );
  NAND2_X1 U12887 ( .A1(n10334), .A2(n10333), .ZN(n14407) );
  OR2_X1 U12888 ( .A1(n14402), .A2(n10332), .ZN(n10664) );
  INV_X1 U12889 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n11799) );
  MUX2_X1 U12890 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n11799), .S(n11224), .Z(
        n10663) );
  AOI21_X1 U12891 ( .B1(n14407), .B2(n10664), .A(n10663), .ZN(n10662) );
  NOR2_X1 U12892 ( .A1(n11224), .A2(n11799), .ZN(n10335) );
  INV_X1 U12893 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n11232) );
  MUX2_X1 U12894 ( .A(n11232), .B(P1_REG2_REG_5__SCAN_IN), .S(n11329), .Z(
        n10336) );
  OAI21_X1 U12895 ( .B1(n10662), .B2(n10335), .A(n10336), .ZN(n10356) );
  INV_X1 U12896 ( .A(n10356), .ZN(n10338) );
  NOR3_X1 U12897 ( .A1(n10662), .A2(n10336), .A3(n10335), .ZN(n10337) );
  NOR3_X1 U12898 ( .A1(n15121), .A2(n10338), .A3(n10337), .ZN(n10339) );
  AOI211_X1 U12899 ( .C1(n14477), .C2(n10341), .A(n10340), .B(n10339), .ZN(
        n10342) );
  INV_X1 U12900 ( .A(n10342), .ZN(P1_U3248) );
  NAND2_X1 U12901 ( .A1(n11543), .A2(n6667), .ZN(n10343) );
  OAI21_X1 U12902 ( .B1(n6667), .B2(n10344), .A(n10343), .ZN(P3_U3495) );
  NAND2_X1 U12903 ( .A1(n11181), .A2(n6667), .ZN(n10345) );
  OAI21_X1 U12904 ( .B1(P3_U3897), .B2(n10346), .A(n10345), .ZN(P3_U3496) );
  NAND2_X1 U12905 ( .A1(n11091), .A2(n6667), .ZN(n10347) );
  OAI21_X1 U12906 ( .B1(P3_U3897), .B2(n10348), .A(n10347), .ZN(P3_U3494) );
  NAND2_X1 U12907 ( .A1(n13312), .A2(n6667), .ZN(n10349) );
  OAI21_X1 U12908 ( .B1(P3_U3897), .B2(n10350), .A(n10349), .ZN(P3_U3505) );
  OAI21_X1 U12909 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n10354), .A(n10351), .ZN(
        n10353) );
  INV_X1 U12910 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n15178) );
  MUX2_X1 U12911 ( .A(P1_REG1_REG_6__SCAN_IN), .B(n15178), .S(n10400), .Z(
        n10352) );
  NOR2_X1 U12912 ( .A1(n10353), .A2(n10352), .ZN(n10472) );
  AOI211_X1 U12913 ( .C1(n10353), .C2(n10352), .A(n10472), .B(n15124), .ZN(
        n10360) );
  NAND2_X1 U12914 ( .A1(n10354), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n10355) );
  MUX2_X1 U12915 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n11367), .S(n10400), .Z(
        n10357) );
  AOI21_X1 U12916 ( .B1(n10356), .B2(n10355), .A(n10357), .ZN(n10395) );
  AND3_X1 U12917 ( .A1(n10357), .A2(n10356), .A3(n10355), .ZN(n10358) );
  NOR3_X1 U12918 ( .A1(n15121), .A2(n10395), .A3(n10358), .ZN(n10359) );
  NOR2_X1 U12919 ( .A1(n10360), .A2(n10359), .ZN(n10362) );
  AND2_X1 U12920 ( .A1(P1_U3086), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n14325) );
  AOI21_X1 U12921 ( .B1(n14435), .B2(P1_ADDR_REG_6__SCAN_IN), .A(n14325), .ZN(
        n10361) );
  OAI211_X1 U12922 ( .C1(n10400), .C2(n15122), .A(n10362), .B(n10361), .ZN(
        P1_U3249) );
  NAND2_X1 U12923 ( .A1(n12004), .A2(n6667), .ZN(n10363) );
  OAI21_X1 U12924 ( .B1(P3_U3897), .B2(n10364), .A(n10363), .ZN(P3_U3499) );
  NAND2_X1 U12925 ( .A1(n12398), .A2(n6667), .ZN(n10365) );
  OAI21_X1 U12926 ( .B1(P3_U3897), .B2(n10366), .A(n10365), .ZN(P3_U3502) );
  NAND2_X1 U12927 ( .A1(n11714), .A2(n6667), .ZN(n10367) );
  OAI21_X1 U12928 ( .B1(P3_U3897), .B2(n10368), .A(n10367), .ZN(P3_U3498) );
  NAND2_X1 U12929 ( .A1(n13532), .A2(n6667), .ZN(n10369) );
  OAI21_X1 U12930 ( .B1(n6667), .B2(n10370), .A(n10369), .ZN(P3_U3508) );
  NAND2_X1 U12931 ( .A1(n13256), .A2(n6667), .ZN(n10371) );
  OAI21_X1 U12932 ( .B1(n6667), .B2(n10372), .A(n10371), .ZN(P3_U3507) );
  NAND2_X1 U12933 ( .A1(n13186), .A2(n6667), .ZN(n10373) );
  OAI21_X1 U12934 ( .B1(P3_U3897), .B2(n10374), .A(n10373), .ZN(P3_U3504) );
  NAND2_X1 U12935 ( .A1(n13140), .A2(n6667), .ZN(n10375) );
  OAI21_X1 U12936 ( .B1(P3_U3897), .B2(n10376), .A(n10375), .ZN(P3_U3506) );
  NOR2_X1 U12937 ( .A1(n10377), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10382) );
  AOI211_X1 U12938 ( .C1(n10380), .C2(n10379), .A(n10378), .B(n12354), .ZN(
        n10381) );
  AOI211_X1 U12939 ( .C1(n15250), .C2(P2_ADDR_REG_2__SCAN_IN), .A(n10382), .B(
        n10381), .ZN(n10388) );
  MUX2_X1 U12940 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n10079), .S(n10389), .Z(
        n10383) );
  NAND3_X1 U12941 ( .A1(n15192), .A2(n10384), .A3(n10383), .ZN(n10385) );
  NAND3_X1 U12942 ( .A1(n15255), .A2(n10386), .A3(n10385), .ZN(n10387) );
  OAI211_X1 U12943 ( .C1(n15225), .C2(n10389), .A(n10388), .B(n10387), .ZN(
        P2_U3216) );
  INV_X1 U12944 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n15348) );
  AOI22_X1 U12945 ( .A1(n15255), .A2(P2_REG1_REG_0__SCAN_IN), .B1(n15252), 
        .B2(P2_REG2_REG_0__SCAN_IN), .ZN(n10392) );
  OAI21_X1 U12946 ( .B1(n12354), .B2(P2_REG2_REG_0__SCAN_IN), .A(n15225), .ZN(
        n10390) );
  AOI21_X1 U12947 ( .B1(n15255), .B2(n15348), .A(n10390), .ZN(n10391) );
  MUX2_X1 U12948 ( .A(n10392), .B(n10391), .S(P2_IR_REG_0__SCAN_IN), .Z(n10394) );
  AOI22_X1 U12949 ( .A1(n15250), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(P2_U3088), 
        .B2(P2_REG3_REG_0__SCAN_IN), .ZN(n10393) );
  NAND2_X1 U12950 ( .A1(n10394), .A2(n10393), .ZN(P2_U3214) );
  INV_X1 U12951 ( .A(n10400), .ZN(n11337) );
  AOI21_X1 U12952 ( .B1(n11337), .B2(P1_REG2_REG_6__SCAN_IN), .A(n10395), .ZN(
        n10463) );
  INV_X1 U12953 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10396) );
  MUX2_X1 U12954 ( .A(n10396), .B(P1_REG2_REG_7__SCAN_IN), .S(n11379), .Z(
        n10462) );
  NOR2_X1 U12955 ( .A1(n10463), .A2(n10462), .ZN(n10461) );
  NOR2_X1 U12956 ( .A1(n10475), .A2(n10396), .ZN(n10419) );
  INV_X1 U12957 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n11703) );
  MUX2_X1 U12958 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n11703), .S(n11684), .Z(
        n10418) );
  OAI21_X1 U12959 ( .B1(n10461), .B2(n10419), .A(n10418), .ZN(n10421) );
  NAND2_X1 U12960 ( .A1(n11684), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n10398) );
  INV_X1 U12961 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10432) );
  MUX2_X1 U12962 ( .A(n10432), .B(P1_REG2_REG_9__SCAN_IN), .S(n11835), .Z(
        n10397) );
  AOI21_X1 U12963 ( .B1(n10421), .B2(n10398), .A(n10397), .ZN(n14421) );
  NAND3_X1 U12964 ( .A1(n10421), .A2(n10398), .A3(n10397), .ZN(n10399) );
  NAND2_X1 U12965 ( .A1(n10399), .A2(n14482), .ZN(n10411) );
  INV_X1 U12966 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n11622) );
  NOR2_X1 U12967 ( .A1(n10400), .A2(n15178), .ZN(n10467) );
  MUX2_X1 U12968 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n11622), .S(n11379), .Z(
        n10401) );
  OAI21_X1 U12969 ( .B1(n11622), .B2(n10475), .A(n10470), .ZN(n10413) );
  INV_X1 U12970 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n11383) );
  MUX2_X1 U12971 ( .A(n11383), .B(P1_REG1_REG_8__SCAN_IN), .S(n11684), .Z(
        n10414) );
  NOR2_X1 U12972 ( .A1(n11684), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n10403) );
  INV_X1 U12973 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10402) );
  MUX2_X1 U12974 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n10402), .S(n11835), .Z(
        n10404) );
  OAI21_X1 U12975 ( .B1(n10412), .B2(n10403), .A(n10404), .ZN(n10427) );
  INV_X1 U12976 ( .A(n10427), .ZN(n10406) );
  NOR3_X1 U12977 ( .A1(n10412), .A2(n10404), .A3(n10403), .ZN(n10405) );
  OAI21_X1 U12978 ( .B1(n10406), .B2(n10405), .A(n14477), .ZN(n10410) );
  INV_X1 U12979 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n12121) );
  NOR2_X1 U12980 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n12121), .ZN(n10408) );
  NOR2_X1 U12981 ( .A1(n15122), .A2(n10433), .ZN(n10407) );
  AOI211_X1 U12982 ( .C1(n14435), .C2(P1_ADDR_REG_9__SCAN_IN), .A(n10408), .B(
        n10407), .ZN(n10409) );
  OAI211_X1 U12983 ( .C1(n14421), .C2(n10411), .A(n10410), .B(n10409), .ZN(
        P1_U3252) );
  AOI21_X1 U12984 ( .B1(n10414), .B2(n10413), .A(n10412), .ZN(n10424) );
  AND2_X1 U12985 ( .A1(P1_U3086), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n10417) );
  NOR2_X1 U12986 ( .A1(n15122), .A2(n10415), .ZN(n10416) );
  AOI211_X1 U12987 ( .C1(n14435), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10417), .B(
        n10416), .ZN(n10423) );
  OR3_X1 U12988 ( .A1(n10461), .A2(n10419), .A3(n10418), .ZN(n10420) );
  NAND3_X1 U12989 ( .A1(n14482), .A2(n10421), .A3(n10420), .ZN(n10422) );
  OAI211_X1 U12990 ( .C1(n10424), .C2(n15124), .A(n10423), .B(n10422), .ZN(
        P1_U3251) );
  NAND2_X1 U12991 ( .A1(n13150), .A2(n6667), .ZN(n10425) );
  OAI21_X1 U12992 ( .B1(P3_U3897), .B2(n10426), .A(n10425), .ZN(P3_U3509) );
  INV_X1 U12993 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n11985) );
  MUX2_X1 U12994 ( .A(n11985), .B(P1_REG1_REG_11__SCAN_IN), .S(n12090), .Z(
        n10430) );
  INV_X1 U12995 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n15182) );
  OAI21_X1 U12996 ( .B1(n11835), .B2(P1_REG1_REG_9__SCAN_IN), .A(n10427), .ZN(
        n14412) );
  MUX2_X1 U12997 ( .A(n15182), .B(P1_REG1_REG_10__SCAN_IN), .S(n14418), .Z(
        n14411) );
  OR2_X1 U12998 ( .A1(n14412), .A2(n14411), .ZN(n14413) );
  OAI21_X1 U12999 ( .B1(n15182), .B2(n10428), .A(n14413), .ZN(n10429) );
  AOI21_X1 U13000 ( .B1(n10430), .B2(n10429), .A(n14430), .ZN(n10441) );
  NAND2_X1 U13001 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n15069)
         );
  OAI21_X1 U13002 ( .B1(n15128), .B2(n10431), .A(n15069), .ZN(n10439) );
  NOR2_X1 U13003 ( .A1(n10433), .A2(n10432), .ZN(n14420) );
  INV_X1 U13004 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n11991) );
  MUX2_X1 U13005 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n11991), .S(n14418), .Z(
        n14419) );
  OAI21_X1 U13006 ( .B1(n14421), .B2(n14420), .A(n14419), .ZN(n14423) );
  NAND2_X1 U13007 ( .A1(n14418), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n10436) );
  INV_X1 U13008 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10434) );
  MUX2_X1 U13009 ( .A(n10434), .B(P1_REG2_REG_11__SCAN_IN), .S(n12090), .Z(
        n10435) );
  AOI21_X1 U13010 ( .B1(n14423), .B2(n10436), .A(n10435), .ZN(n10809) );
  AND3_X1 U13011 ( .A1(n14423), .A2(n10436), .A3(n10435), .ZN(n10437) );
  NOR3_X1 U13012 ( .A1(n10809), .A2(n10437), .A3(n15121), .ZN(n10438) );
  AOI211_X1 U13013 ( .C1(n14480), .C2(n12090), .A(n10439), .B(n10438), .ZN(
        n10440) );
  OAI21_X1 U13014 ( .B1(n10441), .B2(n15124), .A(n10440), .ZN(P1_U3254) );
  OAI222_X1 U13015 ( .A1(n13688), .A2(n10443), .B1(n13690), .B2(n10442), .C1(
        n13374), .C2(P3_U3151), .ZN(P3_U3279) );
  NOR2_X1 U13016 ( .A1(n10455), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n10445) );
  AOI21_X1 U13017 ( .B1(n10445), .B2(n10447), .A(n10444), .ZN(n10460) );
  NOR3_X1 U13018 ( .A1(n10453), .A2(n10446), .A3(n12354), .ZN(n10450) );
  INV_X1 U13019 ( .A(n10447), .ZN(n10448) );
  NOR3_X1 U13020 ( .A1(n13901), .A2(n10448), .A3(n10097), .ZN(n10449) );
  OR3_X1 U13021 ( .A1(n10450), .A2(n15259), .A3(n10449), .ZN(n10456) );
  OAI21_X1 U13022 ( .B1(n10453), .B2(n10452), .A(n10451), .ZN(n10454) );
  AOI22_X1 U13023 ( .A1(n10456), .A2(n10455), .B1(n15252), .B2(n10454), .ZN(
        n10459) );
  AND2_X1 U13024 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n10457) );
  AOI21_X1 U13025 ( .B1(n15250), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n10457), .ZN(
        n10458) );
  OAI211_X1 U13026 ( .C1(n10460), .C2(n13901), .A(n10459), .B(n10458), .ZN(
        P2_U3223) );
  NAND2_X1 U13027 ( .A1(P1_REG3_REG_7__SCAN_IN), .A2(P1_U3086), .ZN(n11872) );
  AOI211_X1 U13028 ( .C1(n10463), .C2(n10462), .A(n10461), .B(n15121), .ZN(
        n10464) );
  INV_X1 U13029 ( .A(n10464), .ZN(n10465) );
  NAND2_X1 U13030 ( .A1(n11872), .A2(n10465), .ZN(n10466) );
  AOI21_X1 U13031 ( .B1(n14435), .B2(P1_ADDR_REG_7__SCAN_IN), .A(n10466), .ZN(
        n10474) );
  MUX2_X1 U13032 ( .A(n11622), .B(P1_REG1_REG_7__SCAN_IN), .S(n11379), .Z(
        n10469) );
  INV_X1 U13033 ( .A(n10467), .ZN(n10468) );
  NAND2_X1 U13034 ( .A1(n10469), .A2(n10468), .ZN(n10471) );
  OAI211_X1 U13035 ( .C1(n10472), .C2(n10471), .A(n14477), .B(n10470), .ZN(
        n10473) );
  OAI211_X1 U13036 ( .C1(n15122), .C2(n10475), .A(n10474), .B(n10473), .ZN(
        P1_U3250) );
  NAND2_X1 U13037 ( .A1(n10478), .A2(n10479), .ZN(n14862) );
  XNOR2_X2 U13038 ( .A(n10477), .B(n10476), .ZN(n10481) );
  XNOR2_X2 U13039 ( .A(n10480), .B(n10479), .ZN(n12951) );
  NAND2_X1 U13040 ( .A1(n12702), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n10486) );
  INV_X1 U13041 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n11785) );
  OR2_X1 U13042 ( .A1(n12753), .A2(n11785), .ZN(n10485) );
  OR2_X1 U13043 ( .A1(n10989), .A2(n10249), .ZN(n10484) );
  INV_X1 U13044 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10493) );
  OR2_X1 U13045 ( .A1(n10832), .A2(n10493), .ZN(n10483) );
  AND4_X2 U13046 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n11320) );
  INV_X1 U13047 ( .A(n11320), .ZN(n14380) );
  INV_X1 U13048 ( .A(n10487), .ZN(n10496) );
  NAND2_X1 U13049 ( .A1(n10496), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10488) );
  MUX2_X1 U13050 ( .A(P1_IR_REG_31__SCAN_IN), .B(n10488), .S(
        P1_IR_REG_20__SCAN_IN), .Z(n10490) );
  NAND2_X1 U13051 ( .A1(n10490), .A2(n10489), .ZN(n12478) );
  AND2_X2 U13052 ( .A1(n10523), .A2(n12540), .ZN(n10616) );
  INV_X1 U13053 ( .A(n10616), .ZN(n12975) );
  INV_X2 U13054 ( .A(n12975), .ZN(n13038) );
  INV_X1 U13055 ( .A(SI_0_), .ZN(n10491) );
  NOR2_X1 U13056 ( .A1(n9213), .A2(n10491), .ZN(n10492) );
  XNOR2_X1 U13057 ( .A(n10492), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14879) );
  AND2_X2 U13058 ( .A1(n10523), .A2(n10620), .ZN(n10617) );
  OAI22_X1 U13059 ( .A1(n11786), .A2(n11858), .B1(n10523), .B2(n10493), .ZN(
        n10494) );
  NAND2_X1 U13060 ( .A1(n14811), .A2(n12475), .ZN(n12465) );
  OAI222_X1 U13061 ( .A1(n11786), .A2(n12975), .B1(n12974), .B2(n11320), .C1(
        n10523), .C2(n7593), .ZN(n10628) );
  XOR2_X1 U13062 ( .A(n10627), .B(n10628), .Z(n10640) );
  OR2_X1 U13063 ( .A1(n10512), .A2(P1_D_REG_1__SCAN_IN), .ZN(n10498) );
  OR2_X1 U13064 ( .A1(n10512), .A2(P1_D_REG_0__SCAN_IN), .ZN(n10500) );
  NOR2_X1 U13065 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n10504) );
  NOR4_X1 U13066 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n10503) );
  NOR4_X1 U13067 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n10502) );
  NOR4_X1 U13068 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n10501) );
  NAND4_X1 U13069 ( .A1(n10504), .A2(n10503), .A3(n10502), .A4(n10501), .ZN(
        n10510) );
  NOR4_X1 U13070 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n10508) );
  NOR4_X1 U13071 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n10507) );
  NOR4_X1 U13072 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n10506) );
  NOR4_X1 U13073 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n10505) );
  NAND4_X1 U13074 ( .A1(n10508), .A2(n10507), .A3(n10506), .A4(n10505), .ZN(
        n10509) );
  NOR2_X1 U13075 ( .A1(n10510), .A2(n10509), .ZN(n10511) );
  OR2_X1 U13076 ( .A1(n10512), .A2(n10511), .ZN(n10891) );
  AND2_X1 U13077 ( .A1(n10891), .A2(n12880), .ZN(n10513) );
  INV_X1 U13078 ( .A(n10888), .ZN(n10514) );
  OR2_X1 U13079 ( .A1(n10514), .A2(n12478), .ZN(n11369) );
  OR2_X1 U13080 ( .A1(n10514), .A2(n12475), .ZN(n10515) );
  NAND2_X1 U13081 ( .A1(n11369), .A2(n10515), .ZN(n15157) );
  NOR2_X1 U13082 ( .A1(n15157), .A2(n12484), .ZN(n10516) );
  NAND2_X1 U13083 ( .A1(n12475), .A2(n12478), .ZN(n10517) );
  NAND2_X1 U13084 ( .A1(n12484), .A2(n10517), .ZN(n12879) );
  NAND2_X1 U13085 ( .A1(n14349), .A2(n14771), .ZN(n15055) );
  INV_X1 U13086 ( .A(n15055), .ZN(n14321) );
  OR2_X1 U13087 ( .A1(n10832), .A2(n10518), .ZN(n10520) );
  INV_X1 U13088 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n11629) );
  NAND2_X1 U13089 ( .A1(n12702), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n10519) );
  NAND3_X1 U13090 ( .A1(n11514), .A2(n11345), .A3(n10891), .ZN(n10521) );
  NAND2_X1 U13091 ( .A1(n14811), .A2(n14483), .ZN(n10892) );
  NAND2_X1 U13092 ( .A1(n10521), .A2(n10892), .ZN(n10525) );
  AND3_X1 U13093 ( .A1(n10523), .A2(n10522), .A3(n12879), .ZN(n10524) );
  NAND2_X1 U13094 ( .A1(n10525), .A2(n10524), .ZN(n10987) );
  OR2_X1 U13095 ( .A1(n10987), .A2(P1_U3086), .ZN(n10839) );
  AOI22_X1 U13096 ( .A1(n14321), .A2(n14378), .B1(P1_REG3_REG_0__SCAN_IN), 
        .B2(n10839), .ZN(n10530) );
  INV_X1 U13097 ( .A(n11369), .ZN(n10526) );
  NAND2_X1 U13098 ( .A1(n10527), .A2(n10526), .ZN(n10528) );
  INV_X1 U13099 ( .A(n10892), .ZN(n11513) );
  INV_X1 U13100 ( .A(n11786), .ZN(n11422) );
  NAND2_X1 U13101 ( .A1(n15067), .A2(n11422), .ZN(n10529) );
  OAI211_X1 U13102 ( .C1(n10640), .C2(n15062), .A(n10530), .B(n10529), .ZN(
        P1_U3232) );
  OAI222_X1 U13103 ( .A1(n13688), .A2(n10533), .B1(n13690), .B2(n10532), .C1(
        n10531), .C2(P3_U3151), .ZN(P3_U3278) );
  INV_X1 U13104 ( .A(n12292), .ZN(n10538) );
  NAND2_X1 U13105 ( .A1(n10534), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10535) );
  INV_X1 U13106 ( .A(n14451), .ZN(n11727) );
  OAI222_X1 U13107 ( .A1(n14876), .A2(n10536), .B1(n11283), .B2(n10538), .C1(
        n11727), .C2(P1_U3086), .ZN(P1_U3341) );
  OAI222_X1 U13108 ( .A1(n14201), .A2(n10539), .B1(n14196), .B2(n10538), .C1(
        n10537), .C2(P2_U3088), .ZN(P2_U3313) );
  OAI222_X1 U13109 ( .A1(n13688), .A2(n10542), .B1(n13690), .B2(n10541), .C1(
        n10540), .C2(P3_U3151), .ZN(P3_U3277) );
  NAND2_X1 U13110 ( .A1(n10543), .A2(n15582), .ZN(n10544) );
  OAI22_X1 U13111 ( .A1(n10565), .A2(n10544), .B1(n11305), .B2(n13520), .ZN(
        n11009) );
  NOR2_X1 U13112 ( .A1(n15607), .A2(n10545), .ZN(n10546) );
  AOI21_X1 U13113 ( .B1(n11009), .B2(n15607), .A(n10546), .ZN(n10547) );
  OAI21_X1 U13114 ( .B1(n10680), .B2(n13623), .A(n10547), .ZN(P3_U3459) );
  NAND2_X1 U13115 ( .A1(n10555), .A2(n15582), .ZN(n10549) );
  OAI22_X1 U13116 ( .A1(n10556), .A2(n10549), .B1(n10559), .B2(n10548), .ZN(
        n10550) );
  NAND2_X1 U13117 ( .A1(n15393), .A2(n13533), .ZN(n13315) );
  INV_X1 U13118 ( .A(n13315), .ZN(n13278) );
  INV_X1 U13119 ( .A(n10553), .ZN(n10552) );
  OR2_X1 U13120 ( .A1(n10552), .A2(n10556), .ZN(n10554) );
  AOI22_X1 U13121 ( .A1(n13278), .A2(n13328), .B1(n11011), .B2(n15377), .ZN(
        n10564) );
  NAND2_X1 U13122 ( .A1(n10556), .A2(n10555), .ZN(n10561) );
  INV_X1 U13123 ( .A(n10557), .ZN(n10558) );
  NAND2_X1 U13124 ( .A1(n10559), .A2(n10558), .ZN(n10560) );
  AND3_X1 U13125 ( .A1(n10561), .A2(n10560), .A3(n11002), .ZN(n11084) );
  NAND2_X1 U13126 ( .A1(n11084), .A2(n10562), .ZN(n10899) );
  NAND2_X1 U13127 ( .A1(n10899), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n10563) );
  OAI211_X1 U13128 ( .C1(n10565), .C2(n15381), .A(n10564), .B(n10563), .ZN(
        P3_U3172) );
  XOR2_X1 U13129 ( .A(n10567), .B(n10566), .Z(n10580) );
  INV_X1 U13130 ( .A(n15520), .ZN(n15485) );
  AOI21_X1 U13131 ( .B1(n10570), .B2(n10569), .A(n10568), .ZN(n10571) );
  NOR2_X1 U13132 ( .A1(n15530), .A2(n10571), .ZN(n10578) );
  AOI21_X1 U13133 ( .B1(n10574), .B2(n10573), .A(n10572), .ZN(n10576) );
  AOI22_X1 U13134 ( .A1(n15523), .A2(P3_ADDR_REG_2__SCAN_IN), .B1(
        P3_REG3_REG_2__SCAN_IN), .B2(P3_U3151), .ZN(n10575) );
  OAI21_X1 U13135 ( .B1(n10576), .B2(n15516), .A(n10575), .ZN(n10577) );
  AOI211_X1 U13136 ( .C1(n15485), .C2(n7768), .A(n10578), .B(n10577), .ZN(
        n10579) );
  OAI21_X1 U13137 ( .B1(n10580), .B2(n7858), .A(n10579), .ZN(P3_U3184) );
  XOR2_X1 U13138 ( .A(n10581), .B(n10582), .Z(n10596) );
  INV_X1 U13139 ( .A(n15530), .ZN(n13387) );
  OAI21_X1 U13140 ( .B1(n10584), .B2(P3_REG2_REG_3__SCAN_IN), .A(n10583), .ZN(
        n10585) );
  NAND2_X1 U13141 ( .A1(n13387), .A2(n10585), .ZN(n10592) );
  INV_X1 U13142 ( .A(n15516), .ZN(n10603) );
  OAI21_X1 U13143 ( .B1(n10587), .B2(P3_REG1_REG_3__SCAN_IN), .A(n10586), .ZN(
        n10588) );
  NAND2_X1 U13144 ( .A1(n10603), .A2(n10588), .ZN(n10591) );
  NAND2_X1 U13145 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_U3151), .ZN(n10590) );
  NAND2_X1 U13146 ( .A1(n15523), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n10589) );
  NAND4_X1 U13147 ( .A1(n10592), .A2(n10591), .A3(n10590), .A4(n10589), .ZN(
        n10593) );
  AOI21_X1 U13148 ( .B1(n10594), .B2(n15485), .A(n10593), .ZN(n10595) );
  OAI21_X1 U13149 ( .B1(n10596), .B2(n7858), .A(n10595), .ZN(P3_U3185) );
  INV_X1 U13150 ( .A(n10597), .ZN(n10600) );
  NAND2_X1 U13151 ( .A1(n10598), .A2(n11665), .ZN(n10599) );
  NAND2_X1 U13152 ( .A1(n10600), .A2(n10599), .ZN(n10601) );
  NAND2_X1 U13153 ( .A1(n13387), .A2(n10601), .ZN(n10611) );
  NOR2_X1 U13154 ( .A1(n10602), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n10604) );
  OAI21_X1 U13155 ( .B1(n10605), .B2(n10604), .A(n10603), .ZN(n10610) );
  AOI22_X1 U13156 ( .A1(n15523), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n10609) );
  XNOR2_X1 U13157 ( .A(n10606), .B(n10962), .ZN(n10607) );
  NAND2_X1 U13158 ( .A1(n10607), .A2(n15504), .ZN(n10608) );
  NAND4_X1 U13159 ( .A1(n10611), .A2(n10610), .A3(n10609), .A4(n10608), .ZN(
        n10612) );
  AOI21_X1 U13160 ( .B1(n10613), .B2(n15485), .A(n10612), .ZN(n10614) );
  INV_X1 U13161 ( .A(n10614), .ZN(P3_U3183) );
  NAND2_X1 U13162 ( .A1(n11355), .A2(n10616), .ZN(n10619) );
  NAND2_X1 U13163 ( .A1(n12530), .A2(n10617), .ZN(n10618) );
  NAND2_X1 U13164 ( .A1(n10619), .A2(n10618), .ZN(n10621) );
  NAND2_X1 U13165 ( .A1(n14878), .A2(n12475), .ZN(n10884) );
  XNOR2_X1 U13166 ( .A(n10621), .B(n10886), .ZN(n10623) );
  NAND2_X1 U13167 ( .A1(n10622), .A2(n10623), .ZN(n10626) );
  INV_X1 U13168 ( .A(n10623), .ZN(n10624) );
  NAND2_X1 U13169 ( .A1(n10625), .A2(n10624), .ZN(n10820) );
  NAND2_X1 U13170 ( .A1(n10626), .A2(n10820), .ZN(n10630) );
  MUX2_X1 U13171 ( .A(n10628), .B(n13057), .S(n10627), .Z(n10629) );
  NOR2_X2 U13172 ( .A1(n10630), .A2(n10629), .ZN(n10822) );
  AOI21_X1 U13173 ( .B1(n10630), .B2(n10629), .A(n10822), .ZN(n10639) );
  INV_X1 U13174 ( .A(n10248), .ZN(n10641) );
  NAND2_X1 U13175 ( .A1(n14349), .A2(n14620), .ZN(n15056) );
  INV_X1 U13176 ( .A(n15056), .ZN(n14322) );
  AOI22_X1 U13177 ( .A1(n14322), .A2(n14380), .B1(n12530), .B2(n15067), .ZN(
        n10638) );
  INV_X1 U13178 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10631) );
  OR2_X1 U13179 ( .A1(n12753), .A2(n10631), .ZN(n10636) );
  OR2_X1 U13180 ( .A1(n10832), .A2(n10632), .ZN(n10633) );
  AOI22_X1 U13181 ( .A1(n14321), .A2(n14377), .B1(P1_REG3_REG_1__SCAN_IN), 
        .B2(n10839), .ZN(n10637) );
  OAI211_X1 U13182 ( .C1(n10639), .C2(n15062), .A(n10638), .B(n10637), .ZN(
        P1_U3222) );
  MUX2_X1 U13183 ( .A(n14386), .B(n10640), .S(n14872), .Z(n10642) );
  NAND2_X1 U13184 ( .A1(n10642), .A2(n10641), .ZN(n10643) );
  OAI211_X1 U13185 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n10644), .A(n10643), .B(
        n14379), .ZN(n10674) );
  MUX2_X1 U13186 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n10645), .S(n10825), .Z(
        n10647) );
  NAND3_X1 U13187 ( .A1(n10647), .A2(n14384), .A3(n10646), .ZN(n10648) );
  NAND3_X1 U13188 ( .A1(n14482), .A2(n14405), .A3(n10648), .ZN(n10656) );
  MUX2_X1 U13189 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n10632), .S(n10825), .Z(
        n10650) );
  NAND3_X1 U13190 ( .A1(n10650), .A2(n14381), .A3(n10649), .ZN(n10651) );
  NAND3_X1 U13191 ( .A1(n14477), .A2(n14399), .A3(n10651), .ZN(n10655) );
  NAND2_X1 U13192 ( .A1(n14480), .A2(n10652), .ZN(n10654) );
  AOI22_X1 U13193 ( .A1(n14435), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10653) );
  AND4_X1 U13194 ( .A1(n10656), .A2(n10655), .A3(n10654), .A4(n10653), .ZN(
        n10657) );
  NAND2_X1 U13195 ( .A1(n10674), .A2(n10657), .ZN(P1_U3245) );
  AND3_X1 U13196 ( .A1(n14401), .A2(n10659), .A3(n10658), .ZN(n10660) );
  NOR3_X1 U13197 ( .A1(n15124), .A2(n10661), .A3(n10660), .ZN(n10671) );
  INV_X1 U13198 ( .A(n10662), .ZN(n10666) );
  NAND3_X1 U13199 ( .A1(n14407), .A2(n10664), .A3(n10663), .ZN(n10665) );
  NAND3_X1 U13200 ( .A1(n14482), .A2(n10666), .A3(n10665), .ZN(n10668) );
  NAND2_X1 U13201 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n10667) );
  OAI211_X1 U13202 ( .C1(n10669), .C2(n15128), .A(n10668), .B(n10667), .ZN(
        n10670) );
  AOI211_X1 U13203 ( .C1(n14480), .C2(n10672), .A(n10671), .B(n10670), .ZN(
        n10673) );
  NAND2_X1 U13204 ( .A1(n10674), .A2(n10673), .ZN(P1_U3247) );
  INV_X1 U13205 ( .A(P3_DATAO_REG_21__SCAN_IN), .ZN(n10676) );
  NAND2_X1 U13206 ( .A1(n13284), .A2(n6667), .ZN(n10675) );
  OAI21_X1 U13207 ( .B1(n6667), .B2(n10676), .A(n10675), .ZN(P3_U3512) );
  INV_X1 U13208 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10677) );
  NOR2_X1 U13209 ( .A1(n15591), .A2(n10677), .ZN(n10678) );
  AOI21_X1 U13210 ( .B1(n11009), .B2(n15591), .A(n10678), .ZN(n10679) );
  OAI21_X1 U13211 ( .B1(n10680), .B2(n13674), .A(n10679), .ZN(P3_U3390) );
  OR2_X1 U13212 ( .A1(n10939), .A2(n15285), .ZN(n15288) );
  INV_X1 U13213 ( .A(n15288), .ZN(n10682) );
  NOR2_X1 U13214 ( .A1(n15287), .A2(n10686), .ZN(n10681) );
  NAND2_X1 U13215 ( .A1(n10682), .A2(n10681), .ZN(n10696) );
  NAND2_X1 U13216 ( .A1(n13852), .A2(n13891), .ZN(n11060) );
  OR2_X1 U13217 ( .A1(n10696), .A2(n10684), .ZN(n10685) );
  INV_X1 U13218 ( .A(n15287), .ZN(n10967) );
  NAND3_X1 U13219 ( .A1(n10967), .A2(n10687), .A3(n10941), .ZN(n10689) );
  NAND2_X1 U13220 ( .A1(n10689), .A2(n10688), .ZN(n10751) );
  INV_X1 U13221 ( .A(n10938), .ZN(n10690) );
  NAND2_X1 U13222 ( .A1(n10751), .A2(n10690), .ZN(n10912) );
  AOI22_X1 U13223 ( .A1(n13857), .A2(n10691), .B1(n10912), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n10701) );
  INV_X1 U13224 ( .A(n10692), .ZN(n10694) );
  NAND2_X1 U13225 ( .A1(n10694), .A2(n15340), .ZN(n10695) );
  OR2_X1 U13226 ( .A1(n11466), .A2(n10697), .ZN(n10729) );
  OAI21_X1 U13227 ( .B1(n10697), .B2(n10698), .A(n11474), .ZN(n10699) );
  NAND3_X1 U13228 ( .A1(n6908), .A2(n10729), .A3(n10699), .ZN(n10700) );
  OAI211_X1 U13229 ( .C1(n13855), .C2(n11060), .A(n10701), .B(n10700), .ZN(
        P2_U3204) );
  INV_X1 U13230 ( .A(n10899), .ZN(n10722) );
  INV_X1 U13231 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n11664) );
  NAND2_X1 U13232 ( .A1(n10704), .A2(n11039), .ZN(n10705) );
  AND2_X1 U13233 ( .A1(n10706), .A2(n10705), .ZN(n10707) );
  NAND3_X1 U13234 ( .A1(n13328), .A2(n13174), .A3(n10719), .ZN(n10710) );
  NAND2_X1 U13235 ( .A1(n10771), .A2(n13174), .ZN(n10711) );
  NAND2_X1 U13236 ( .A1(n10712), .A2(n10711), .ZN(n10713) );
  INV_X1 U13237 ( .A(n10770), .ZN(n10714) );
  NAND3_X1 U13238 ( .A1(n10714), .A2(n10772), .A3(n12432), .ZN(n10715) );
  OAI211_X1 U13239 ( .C1(n10716), .C2(n10771), .A(n10896), .B(n10715), .ZN(
        n10717) );
  NAND2_X1 U13240 ( .A1(n10717), .A2(n15390), .ZN(n10721) );
  INV_X1 U13241 ( .A(n13330), .ZN(n10718) );
  OAI22_X1 U13242 ( .A1(n10718), .A2(n13518), .B1(n8952), .B2(n13520), .ZN(
        n10773) );
  AOI22_X1 U13243 ( .A1(n10773), .A2(n15393), .B1(n10719), .B2(n15377), .ZN(
        n10720) );
  OAI211_X1 U13244 ( .C1(n10722), .C2(n11664), .A(n10721), .B(n10720), .ZN(
        P3_U3162) );
  INV_X1 U13245 ( .A(n10726), .ZN(n10727) );
  XNOR2_X1 U13246 ( .A(n13729), .B(n11116), .ZN(n10778) );
  AND2_X1 U13247 ( .A1(n10734), .A2(n13888), .ZN(n10779) );
  XNOR2_X1 U13248 ( .A(n10778), .B(n10779), .ZN(n10748) );
  NAND2_X1 U13249 ( .A1(n10734), .A2(n13891), .ZN(n10731) );
  XNOR2_X1 U13250 ( .A(n10731), .B(n10730), .ZN(n10914) );
  NAND2_X1 U13251 ( .A1(n10727), .A2(n11474), .ZN(n10728) );
  NAND2_X1 U13252 ( .A1(n10914), .A2(n10915), .ZN(n10913) );
  INV_X1 U13253 ( .A(n10730), .ZN(n10732) );
  NAND2_X1 U13254 ( .A1(n10732), .A2(n10731), .ZN(n10733) );
  INV_X1 U13255 ( .A(n10735), .ZN(n10736) );
  NAND2_X1 U13256 ( .A1(n10737), .A2(n10736), .ZN(n10738) );
  XNOR2_X1 U13257 ( .A(n10726), .B(n15314), .ZN(n10742) );
  INV_X1 U13258 ( .A(n10742), .ZN(n10740) );
  AND2_X1 U13259 ( .A1(n10734), .A2(n13889), .ZN(n10741) );
  INV_X1 U13260 ( .A(n10741), .ZN(n10739) );
  NAND2_X1 U13261 ( .A1(n10740), .A2(n10739), .ZN(n10743) );
  NAND2_X1 U13262 ( .A1(n10742), .A2(n10741), .ZN(n10744) );
  INV_X1 U13263 ( .A(n10747), .ZN(n10746) );
  INV_X1 U13264 ( .A(n10748), .ZN(n10745) );
  NAND2_X1 U13265 ( .A1(n10746), .A2(n10745), .ZN(n10785) );
  INV_X1 U13266 ( .A(n10785), .ZN(n10783) );
  AOI21_X1 U13267 ( .B1(n10748), .B2(n10747), .A(n10783), .ZN(n10756) );
  AOI22_X1 U13268 ( .A1(n13887), .A2(n13852), .B1(n13851), .B2(n13889), .ZN(
        n11121) );
  OAI21_X1 U13269 ( .B1(n13855), .B2(n11121), .A(n10749), .ZN(n10754) );
  NAND2_X1 U13270 ( .A1(n10751), .A2(n10750), .ZN(n10752) );
  NOR2_X1 U13271 ( .A1(n13845), .A2(n11117), .ZN(n10753) );
  AOI211_X1 U13272 ( .C1(n11116), .C2(n13857), .A(n10754), .B(n10753), .ZN(
        n10755) );
  OAI21_X1 U13273 ( .B1(n10756), .B2(n13859), .A(n10755), .ZN(P2_U3202) );
  INV_X1 U13274 ( .A(n12443), .ZN(n10765) );
  NAND2_X1 U13275 ( .A1(n10758), .A2(n10757), .ZN(n10759) );
  OR3_X1 U13276 ( .A1(n10761), .A2(n10760), .A3(n10759), .ZN(n10872) );
  NAND2_X1 U13277 ( .A1(n10872), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n10762) );
  XNOR2_X1 U13278 ( .A(n10762), .B(P1_IR_REG_15__SCAN_IN), .ZN(n12444) );
  INV_X1 U13279 ( .A(n12444), .ZN(n15111) );
  OAI222_X1 U13280 ( .A1(n14876), .A2(n10763), .B1(n11283), .B2(n10765), .C1(
        n15111), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U13281 ( .A(n10764), .ZN(n11812) );
  OAI222_X1 U13282 ( .A1(n14201), .A2(n10766), .B1(n14196), .B2(n10765), .C1(
        n11812), .C2(P2_U3088), .ZN(P2_U3312) );
  OAI222_X1 U13283 ( .A1(n13688), .A2(n10769), .B1(n10768), .B2(P3_U3151), 
        .C1(n10767), .C2(n13690), .ZN(P3_U3276) );
  XNOR2_X1 U13284 ( .A(n10772), .B(n10770), .ZN(n11669) );
  XNOR2_X1 U13285 ( .A(n10772), .B(n10771), .ZN(n10774) );
  AOI21_X1 U13286 ( .B1(n10774), .B2(n13552), .A(n10773), .ZN(n11662) );
  OAI21_X1 U13287 ( .B1(n15570), .B2(n11669), .A(n11662), .ZN(n10882) );
  INV_X1 U13288 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n10775) );
  OAI22_X1 U13289 ( .A1(n13623), .A2(n8956), .B1(n15607), .B2(n10775), .ZN(
        n10776) );
  AOI21_X1 U13290 ( .B1(n10882), .B2(n15607), .A(n10776), .ZN(n10777) );
  INV_X1 U13291 ( .A(n10777), .ZN(P3_U3460) );
  INV_X1 U13292 ( .A(n10778), .ZN(n10781) );
  INV_X1 U13293 ( .A(n10779), .ZN(n10780) );
  NAND2_X1 U13294 ( .A1(n10781), .A2(n10780), .ZN(n10784) );
  INV_X1 U13295 ( .A(n10784), .ZN(n10782) );
  XNOR2_X1 U13296 ( .A(n15332), .B(n13729), .ZN(n10921) );
  AND2_X1 U13297 ( .A1(n13887), .A2(n10734), .ZN(n10919) );
  XNOR2_X1 U13298 ( .A(n10921), .B(n10919), .ZN(n10786) );
  NOR3_X1 U13299 ( .A1(n10783), .A2(n10782), .A3(n10786), .ZN(n10789) );
  NAND2_X1 U13300 ( .A1(n10785), .A2(n10784), .ZN(n10787) );
  NAND2_X1 U13301 ( .A1(n10787), .A2(n10786), .ZN(n10923) );
  INV_X1 U13302 ( .A(n10923), .ZN(n10788) );
  OAI21_X1 U13303 ( .B1(n10789), .B2(n10788), .A(n6908), .ZN(n10793) );
  AOI22_X1 U13304 ( .A1(n13852), .A2(n13886), .B1(n13851), .B2(n13888), .ZN(
        n11146) );
  OAI21_X1 U13305 ( .B1(n13855), .B2(n11146), .A(n10790), .ZN(n10791) );
  AOI21_X1 U13306 ( .B1(n11141), .B2(n13857), .A(n10791), .ZN(n10792) );
  OAI211_X1 U13307 ( .C1(n13845), .C2(n11142), .A(n10793), .B(n10792), .ZN(
        P2_U3199) );
  NAND3_X1 U13308 ( .A1(n10846), .A2(n10795), .A3(n10794), .ZN(n10796) );
  NAND2_X1 U13309 ( .A1(n10796), .A2(n15255), .ZN(n10804) );
  OAI21_X1 U13310 ( .B1(n10798), .B2(n10797), .A(n10857), .ZN(n10799) );
  NAND2_X1 U13311 ( .A1(n10799), .A2(n15252), .ZN(n10803) );
  AND2_X1 U13312 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3088), .ZN(n11676) );
  NOR2_X1 U13313 ( .A1(n15225), .A2(n10800), .ZN(n10801) );
  AOI211_X1 U13314 ( .C1(n15250), .C2(P2_ADDR_REG_11__SCAN_IN), .A(n11676), 
        .B(n10801), .ZN(n10802) );
  OAI211_X1 U13315 ( .C1(n10805), .C2(n10804), .A(n10803), .B(n10802), .ZN(
        P2_U3225) );
  NOR2_X1 U13316 ( .A1(n12090), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n14428) );
  INV_X1 U13317 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n14912) );
  MUX2_X1 U13318 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n14912), .S(n14440), .Z(
        n14429) );
  OAI21_X1 U13319 ( .B1(n14430), .B2(n14428), .A(n14429), .ZN(n14427) );
  OAI21_X1 U13320 ( .B1(n14440), .B2(P1_REG1_REG_12__SCAN_IN), .A(n14427), 
        .ZN(n10807) );
  INV_X1 U13321 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n12379) );
  MUX2_X1 U13322 ( .A(n12379), .B(P1_REG1_REG_13__SCAN_IN), .S(n12240), .Z(
        n10806) );
  NOR2_X1 U13323 ( .A1(n10807), .A2(n10806), .ZN(n11732) );
  AOI211_X1 U13324 ( .C1(n10807), .C2(n10806), .A(n15124), .B(n11732), .ZN(
        n10808) );
  INV_X1 U13325 ( .A(n10808), .ZN(n10817) );
  NAND2_X1 U13326 ( .A1(P1_REG3_REG_13__SCAN_IN), .A2(P1_U3086), .ZN(n14293)
         );
  INV_X1 U13327 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n11724) );
  MUX2_X1 U13328 ( .A(n11724), .B(P1_REG2_REG_13__SCAN_IN), .S(n12240), .Z(
        n10812) );
  AOI21_X1 U13329 ( .B1(n12090), .B2(P1_REG2_REG_11__SCAN_IN), .A(n10809), 
        .ZN(n14437) );
  INV_X1 U13330 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n10810) );
  MUX2_X1 U13331 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n10810), .S(n14440), .Z(
        n14438) );
  NAND2_X1 U13332 ( .A1(n14437), .A2(n14438), .ZN(n14436) );
  OAI21_X1 U13333 ( .B1(n14440), .B2(P1_REG2_REG_12__SCAN_IN), .A(n14436), 
        .ZN(n10811) );
  NOR2_X1 U13334 ( .A1(n10811), .A2(n10812), .ZN(n14458) );
  AOI211_X1 U13335 ( .C1(n10812), .C2(n10811), .A(n14458), .B(n15121), .ZN(
        n10813) );
  INV_X1 U13336 ( .A(n10813), .ZN(n10814) );
  NAND2_X1 U13337 ( .A1(n14293), .A2(n10814), .ZN(n10815) );
  AOI21_X1 U13338 ( .B1(n14435), .B2(P1_ADDR_REG_13__SCAN_IN), .A(n10815), 
        .ZN(n10816) );
  OAI211_X1 U13339 ( .C1(n15122), .C2(n11725), .A(n10817), .B(n10816), .ZN(
        P1_U3256) );
  NAND2_X1 U13340 ( .A1(n13494), .A2(n6667), .ZN(n10818) );
  OAI21_X1 U13341 ( .B1(P3_U3897), .B2(n10819), .A(n10818), .ZN(P3_U3513) );
  OR2_X1 U13342 ( .A1(n12820), .A2(n10823), .ZN(n10824) );
  AOI22_X1 U13343 ( .A1(n14377), .A2(n13059), .B1(n13070), .B2(n11434), .ZN(
        n10976) );
  NAND2_X1 U13344 ( .A1(n14377), .A2(n13038), .ZN(n10827) );
  NAND2_X1 U13345 ( .A1(n11434), .A2(n10617), .ZN(n10826) );
  NAND2_X1 U13346 ( .A1(n10827), .A2(n10826), .ZN(n10828) );
  XNOR2_X1 U13347 ( .A(n10828), .B(n10886), .ZN(n10975) );
  AOI21_X1 U13348 ( .B1(n10830), .B2(n10829), .A(n6801), .ZN(n10841) );
  INV_X1 U13349 ( .A(n11434), .ZN(n12533) );
  INV_X1 U13350 ( .A(n15067), .ZN(n14352) );
  INV_X1 U13351 ( .A(n14349), .ZN(n14306) );
  NAND2_X1 U13352 ( .A1(n12812), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n10837) );
  OR2_X1 U13353 ( .A1(n12786), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n10836) );
  INV_X2 U13354 ( .A(n12702), .ZN(n10990) );
  INV_X1 U13355 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n10831) );
  OR2_X1 U13356 ( .A1(n10990), .A2(n10831), .ZN(n10835) );
  OR2_X1 U13357 ( .A1(n12670), .A2(n10833), .ZN(n10834) );
  AOI22_X1 U13358 ( .A1(n14620), .A2(n14378), .B1(n14376), .B2(n14771), .ZN(
        n11438) );
  OAI22_X1 U13359 ( .A1(n12533), .A2(n14352), .B1(n14306), .B2(n11438), .ZN(
        n10838) );
  AOI21_X1 U13360 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n10839), .A(n10838), .ZN(
        n10840) );
  OAI21_X1 U13361 ( .B1(n10841), .B2(n15062), .A(n10840), .ZN(P1_U3237) );
  AOI211_X1 U13362 ( .C1(n10844), .C2(n10843), .A(n10842), .B(n12354), .ZN(
        n10845) );
  INV_X1 U13363 ( .A(n10845), .ZN(n10850) );
  OAI211_X1 U13364 ( .C1(n10848), .C2(n10847), .A(n15255), .B(n10846), .ZN(
        n10849) );
  NAND2_X1 U13365 ( .A1(n10850), .A2(n10849), .ZN(n10852) );
  NAND2_X1 U13366 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3088), .ZN(n11461)
         );
  INV_X1 U13367 ( .A(n11461), .ZN(n10851) );
  AOI211_X1 U13368 ( .C1(n15250), .C2(P2_ADDR_REG_10__SCAN_IN), .A(n10852), 
        .B(n10851), .ZN(n10853) );
  OAI21_X1 U13369 ( .B1(n10854), .B2(n15225), .A(n10853), .ZN(P2_U3224) );
  AND3_X1 U13370 ( .A1(n10857), .A2(n10856), .A3(n10855), .ZN(n10858) );
  OAI21_X1 U13371 ( .B1(n10859), .B2(n10858), .A(n15252), .ZN(n10869) );
  INV_X1 U13372 ( .A(n10860), .ZN(n10861) );
  OAI21_X1 U13373 ( .B1(n10863), .B2(n10862), .A(n10861), .ZN(n10867) );
  NOR2_X1 U13374 ( .A1(n15225), .A2(n10864), .ZN(n10866) );
  NAND2_X1 U13375 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3088), .ZN(n11927)
         );
  OAI21_X1 U13376 ( .B1(n15228), .B2(n15088), .A(n11927), .ZN(n10865) );
  AOI211_X1 U13377 ( .C1(n10867), .C2(n15255), .A(n10866), .B(n10865), .ZN(
        n10868) );
  NAND2_X1 U13378 ( .A1(n10869), .A2(n10868), .ZN(P2_U3226) );
  INV_X1 U13379 ( .A(n12627), .ZN(n10878) );
  OAI222_X1 U13380 ( .A1(n14201), .A2(n10871), .B1(n14196), .B2(n10878), .C1(
        n10870), .C2(P2_U3088), .ZN(P2_U3311) );
  NOR2_X1 U13381 ( .A1(n10872), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n10875) );
  NOR2_X1 U13382 ( .A1(n10875), .A2(n14864), .ZN(n10873) );
  MUX2_X1 U13383 ( .A(n14864), .B(n10873), .S(P1_IR_REG_16__SCAN_IN), .Z(
        n10877) );
  NAND2_X1 U13384 ( .A1(n10875), .A2(n10874), .ZN(n10972) );
  INV_X1 U13385 ( .A(n10972), .ZN(n10876) );
  NOR2_X1 U13386 ( .A1(n10877), .A2(n10876), .ZN(n12628) );
  INV_X1 U13387 ( .A(n12628), .ZN(n12022) );
  OAI222_X1 U13388 ( .A1(n14876), .A2(n10879), .B1(n11283), .B2(n10878), .C1(
        n12022), .C2(P1_U3086), .ZN(P1_U3339) );
  INV_X1 U13389 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n10880) );
  OAI22_X1 U13390 ( .A1(n13674), .A2(n8956), .B1(n15591), .B2(n10880), .ZN(
        n10881) );
  AOI21_X1 U13391 ( .B1(n10882), .B2(n15591), .A(n10881), .ZN(n10883) );
  INV_X1 U13392 ( .A(n10883), .ZN(P3_U3393) );
  OR2_X1 U13393 ( .A1(n11320), .A2(n11422), .ZN(n12541) );
  NAND2_X1 U13394 ( .A1(n11320), .A2(n11422), .ZN(n12539) );
  NAND2_X1 U13395 ( .A1(n12541), .A2(n12539), .ZN(n12840) );
  INV_X1 U13396 ( .A(n10884), .ZN(n10885) );
  NAND2_X1 U13397 ( .A1(n10885), .A2(n12540), .ZN(n10887) );
  NAND2_X1 U13398 ( .A1(n10887), .A2(n10886), .ZN(n11605) );
  OR2_X1 U13399 ( .A1(n11605), .A2(n14483), .ZN(n11347) );
  AND2_X1 U13400 ( .A1(n12474), .A2(n12478), .ZN(n12483) );
  NAND2_X1 U13401 ( .A1(n12483), .A2(n14483), .ZN(n15161) );
  NAND2_X1 U13402 ( .A1(n14878), .A2(n14483), .ZN(n12477) );
  INV_X1 U13403 ( .A(n12478), .ZN(n12485) );
  NAND2_X1 U13404 ( .A1(n12500), .A2(n12485), .ZN(n12492) );
  NAND2_X1 U13405 ( .A1(n12477), .A2(n12492), .ZN(n14618) );
  NAND2_X1 U13406 ( .A1(n14815), .A2(n14699), .ZN(n10889) );
  AOI222_X1 U13407 ( .A1(n12840), .A2(n10889), .B1(n10888), .B2(n11422), .C1(
        n14378), .C2(n14771), .ZN(n15155) );
  AND2_X1 U13408 ( .A1(n12880), .A2(n12879), .ZN(n10890) );
  NAND2_X1 U13409 ( .A1(n10891), .A2(n10890), .ZN(n11343) );
  OR2_X1 U13410 ( .A1(n11345), .A2(n11343), .ZN(n11516) );
  NAND2_X1 U13411 ( .A1(n11514), .A2(n10892), .ZN(n10893) );
  NAND2_X1 U13412 ( .A1(n15181), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n10894) );
  OAI21_X1 U13413 ( .B1(n15155), .B2(n15181), .A(n10894), .ZN(P1_U3528) );
  XNOR2_X1 U13414 ( .A(n11713), .B(n11309), .ZN(n11088) );
  XNOR2_X1 U13415 ( .A(n11088), .B(n13327), .ZN(n11087) );
  NAND2_X1 U13416 ( .A1(n10896), .A2(n10895), .ZN(n11086) );
  XOR2_X1 U13417 ( .A(n11086), .B(n11087), .Z(n10901) );
  NAND2_X1 U13418 ( .A1(n15393), .A2(n13531), .ZN(n13295) );
  AOI22_X1 U13419 ( .A1(n13278), .A2(n11091), .B1(n11309), .B2(n15377), .ZN(
        n10897) );
  OAI21_X1 U13420 ( .B1(n11305), .B2(n13295), .A(n10897), .ZN(n10898) );
  AOI21_X1 U13421 ( .B1(P3_REG3_REG_2__SCAN_IN), .B2(n10899), .A(n10898), .ZN(
        n10900) );
  OAI21_X1 U13422 ( .B1(n10901), .B2(n15381), .A(n10900), .ZN(P3_U3177) );
  INV_X1 U13423 ( .A(n13857), .ZN(n13812) );
  OAI22_X1 U13424 ( .A1(n10903), .A2(n13839), .B1(n10902), .B2(n13841), .ZN(
        n15266) );
  AOI22_X1 U13425 ( .A1(n13843), .A2(n15266), .B1(P2_REG3_REG_2__SCAN_IN), 
        .B2(n10912), .ZN(n10909) );
  OAI21_X1 U13426 ( .B1(n10906), .B2(n10905), .A(n10904), .ZN(n10907) );
  NAND2_X1 U13427 ( .A1(n6908), .A2(n10907), .ZN(n10908) );
  OAI211_X1 U13428 ( .C1(n15306), .C2(n13812), .A(n10909), .B(n10908), .ZN(
        P2_U3209) );
  OR2_X1 U13429 ( .A1(n9722), .A2(n13841), .ZN(n10911) );
  NAND2_X1 U13430 ( .A1(n13851), .A2(n9763), .ZN(n10910) );
  NAND2_X1 U13431 ( .A1(n10911), .A2(n10910), .ZN(n11470) );
  AOI22_X1 U13432 ( .A1(n13843), .A2(n11470), .B1(n10912), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n10918) );
  OAI21_X1 U13433 ( .B1(n10915), .B2(n10914), .A(n10913), .ZN(n10916) );
  NAND2_X1 U13434 ( .A1(n6908), .A2(n10916), .ZN(n10917) );
  OAI211_X1 U13435 ( .C1(n15300), .C2(n13812), .A(n10918), .B(n10917), .ZN(
        P2_U3194) );
  INV_X1 U13436 ( .A(n10919), .ZN(n10920) );
  NAND2_X1 U13437 ( .A1(n10921), .A2(n10920), .ZN(n10922) );
  XNOR2_X1 U13438 ( .A(n10945), .B(n13734), .ZN(n10924) );
  AND2_X1 U13439 ( .A1(n10734), .A2(n13886), .ZN(n10925) );
  NAND2_X1 U13440 ( .A1(n10924), .A2(n10925), .ZN(n11015) );
  INV_X1 U13441 ( .A(n10924), .ZN(n10927) );
  INV_X1 U13442 ( .A(n10925), .ZN(n10926) );
  NAND2_X1 U13443 ( .A1(n10927), .A2(n10926), .ZN(n10928) );
  NAND2_X1 U13444 ( .A1(n11015), .A2(n10928), .ZN(n10930) );
  AOI21_X1 U13445 ( .B1(n10929), .B2(n10930), .A(n13859), .ZN(n10932) );
  NAND2_X1 U13446 ( .A1(n10932), .A2(n11016), .ZN(n10936) );
  AOI22_X1 U13447 ( .A1(n13852), .A2(n13885), .B1(n13887), .B2(n13851), .ZN(
        n10948) );
  OAI22_X1 U13448 ( .A1(n13855), .A2(n10948), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10933), .ZN(n10934) );
  AOI21_X1 U13449 ( .B1(n10945), .B2(n13857), .A(n10934), .ZN(n10935) );
  OAI211_X1 U13450 ( .C1(n13845), .C2(n11129), .A(n10936), .B(n10935), .ZN(
        P2_U3211) );
  NOR2_X1 U13451 ( .A1(n10938), .A2(n10937), .ZN(n10940) );
  INV_X1 U13452 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10953) );
  NAND2_X1 U13453 ( .A1(n11556), .A2(n11063), .ZN(n15334) );
  XNOR2_X1 U13454 ( .A(n10943), .B(n10942), .ZN(n11135) );
  INV_X1 U13455 ( .A(n11139), .ZN(n10944) );
  AOI211_X1 U13456 ( .C1(n10945), .C2(n10944), .A(n14091), .B(n11024), .ZN(
        n11132) );
  AOI21_X1 U13457 ( .B1(n15313), .B2(n10945), .A(n11132), .ZN(n10951) );
  XNOR2_X1 U13458 ( .A(n10947), .B(n10946), .ZN(n10950) );
  INV_X1 U13459 ( .A(n10948), .ZN(n10949) );
  AOI21_X1 U13460 ( .B1(n10950), .B2(n14065), .A(n10949), .ZN(n11127) );
  OAI211_X1 U13461 ( .C1(n15000), .C2(n11135), .A(n10951), .B(n11127), .ZN(
        n10969) );
  NAND2_X1 U13462 ( .A1(n10969), .A2(n15347), .ZN(n10952) );
  OAI21_X1 U13463 ( .B1(n15347), .B2(n10953), .A(n10952), .ZN(P2_U3448) );
  NAND3_X1 U13464 ( .A1(n15530), .A2(n15516), .A3(n7858), .ZN(n10961) );
  INV_X1 U13465 ( .A(n10954), .ZN(n10956) );
  OAI22_X1 U13466 ( .A1(n15530), .A2(n10956), .B1(n15516), .B2(n10955), .ZN(
        n10960) );
  INV_X1 U13467 ( .A(n15523), .ZN(n15492) );
  OAI22_X1 U13468 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n10958), .B1(n10957), .B2(
        n15492), .ZN(n10959) );
  AOI211_X1 U13469 ( .C1(n10962), .C2(n10961), .A(n10960), .B(n10959), .ZN(
        n10966) );
  OR2_X1 U13470 ( .A1(n7858), .A2(n10963), .ZN(n10964) );
  MUX2_X1 U13471 ( .A(n10964), .B(n15520), .S(P3_IR_REG_0__SCAN_IN), .Z(n10965) );
  NAND2_X1 U13472 ( .A1(n10966), .A2(n10965), .ZN(P3_U3182) );
  NAND2_X1 U13473 ( .A1(n10969), .A2(n15357), .ZN(n10970) );
  OAI21_X1 U13474 ( .B1(n15357), .B2(n10089), .A(n10970), .ZN(P2_U3505) );
  INV_X1 U13475 ( .A(n12638), .ZN(n10973) );
  OAI222_X1 U13476 ( .A1(n14201), .A2(n10971), .B1(n14196), .B2(n10973), .C1(
        n12344), .C2(P2_U3088), .ZN(P2_U3310) );
  NAND2_X1 U13477 ( .A1(n10972), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11109) );
  XNOR2_X1 U13478 ( .A(n11109), .B(P1_IR_REG_17__SCAN_IN), .ZN(n14467) );
  INV_X1 U13479 ( .A(n14467), .ZN(n14463) );
  OAI222_X1 U13480 ( .A1(n14876), .A2(n10974), .B1(n11283), .B2(n10973), .C1(
        n14463), .C2(P1_U3086), .ZN(P1_U3338) );
  NAND2_X1 U13481 ( .A1(n14376), .A2(n13070), .ZN(n10982) );
  OR2_X1 U13482 ( .A1(n12820), .A2(n10979), .ZN(n10980) );
  NAND2_X1 U13483 ( .A1(n15139), .A2(n13086), .ZN(n10981) );
  NAND2_X1 U13484 ( .A1(n10982), .A2(n10981), .ZN(n10983) );
  XNOR2_X1 U13485 ( .A(n10983), .B(n10886), .ZN(n11227) );
  AND2_X1 U13486 ( .A1(n15139), .A2(n13085), .ZN(n10984) );
  AOI21_X1 U13487 ( .B1(n14376), .B2(n13087), .A(n10984), .ZN(n11230) );
  XNOR2_X1 U13488 ( .A(n11227), .B(n11230), .ZN(n10985) );
  OAI211_X1 U13489 ( .C1(n10986), .C2(n10985), .A(n11228), .B(n14341), .ZN(
        n11001) );
  INV_X1 U13490 ( .A(n15072), .ZN(n14338) );
  INV_X1 U13491 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n15141) );
  INV_X1 U13492 ( .A(n10988), .ZN(n11578) );
  NAND2_X1 U13493 ( .A1(n14377), .A2(n14620), .ZN(n10997) );
  INV_X4 U13494 ( .A(n12670), .ZN(n12811) );
  NAND2_X1 U13495 ( .A1(n12811), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n10995) );
  OR2_X1 U13496 ( .A1(n12664), .A2(n11799), .ZN(n10994) );
  XNOR2_X1 U13497 ( .A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n11798) );
  OR2_X1 U13498 ( .A1(n12753), .A2(n11798), .ZN(n10993) );
  INV_X1 U13499 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10991) );
  NAND2_X1 U13500 ( .A1(n14375), .A2(n14771), .ZN(n10996) );
  NAND2_X1 U13501 ( .A1(n10997), .A2(n10996), .ZN(n11494) );
  AOI22_X1 U13502 ( .A1(n14349), .A2(n11494), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(P1_U3086), .ZN(n10998) );
  OAI21_X1 U13503 ( .B1(n14352), .B2(n11578), .A(n10998), .ZN(n10999) );
  AOI21_X1 U13504 ( .B1(n14338), .B2(n15141), .A(n10999), .ZN(n11000) );
  NAND2_X1 U13505 ( .A1(n11001), .A2(n11000), .ZN(P1_U3218) );
  INV_X1 U13506 ( .A(n11002), .ZN(n11003) );
  NOR2_X1 U13507 ( .A1(n11006), .A2(n11003), .ZN(n11005) );
  MUX2_X1 U13508 ( .A(n11006), .B(n11005), .S(n11004), .Z(n11007) );
  NAND2_X1 U13509 ( .A1(n11008), .A2(n11007), .ZN(n11010) );
  NAND2_X1 U13510 ( .A1(n11009), .A2(n13541), .ZN(n11013) );
  NAND2_X1 U13511 ( .A1(n11314), .A2(n15561), .ZN(n11663) );
  AOI22_X1 U13512 ( .A1(n13543), .A2(n11011), .B1(n13559), .B2(
        P3_REG3_REG_0__SCAN_IN), .ZN(n11012) );
  OAI211_X1 U13513 ( .C1(n11014), .C2(n13541), .A(n11013), .B(n11012), .ZN(
        P3_U3233) );
  XNOR2_X1 U13514 ( .A(n11265), .B(n10727), .ZN(n11195) );
  OR2_X1 U13515 ( .A1(n10697), .A2(n11075), .ZN(n11193) );
  XNOR2_X1 U13516 ( .A(n11195), .B(n11193), .ZN(n11017) );
  OAI211_X1 U13517 ( .C1(n11018), .C2(n11017), .A(n11197), .B(n6908), .ZN(
        n11021) );
  AOI22_X1 U13518 ( .A1(n13884), .A2(n13852), .B1(n13851), .B2(n13886), .ZN(
        n11030) );
  NAND2_X1 U13519 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n15226) );
  OAI21_X1 U13520 ( .B1(n13855), .B2(n11030), .A(n15226), .ZN(n11019) );
  AOI21_X1 U13521 ( .B1(n11027), .B2(n13857), .A(n11019), .ZN(n11020) );
  OAI211_X1 U13522 ( .C1(n13845), .C2(n11262), .A(n11021), .B(n11020), .ZN(
        P2_U3185) );
  XNOR2_X1 U13523 ( .A(n11023), .B(n11022), .ZN(n11266) );
  INV_X1 U13524 ( .A(n11024), .ZN(n11026) );
  INV_X1 U13525 ( .A(n11072), .ZN(n11025) );
  AOI211_X1 U13526 ( .C1(n11027), .C2(n11026), .A(n14091), .B(n11025), .ZN(
        n11269) );
  AOI21_X1 U13527 ( .B1(n15313), .B2(n11027), .A(n11269), .ZN(n11033) );
  XNOR2_X1 U13528 ( .A(n11029), .B(n11028), .ZN(n11032) );
  INV_X1 U13529 ( .A(n11030), .ZN(n11031) );
  AOI21_X1 U13530 ( .B1(n11032), .B2(n14065), .A(n11031), .ZN(n11271) );
  OAI211_X1 U13531 ( .C1(n15000), .C2(n11266), .A(n11033), .B(n11271), .ZN(
        n11035) );
  NAND2_X1 U13532 ( .A1(n11035), .A2(n15347), .ZN(n11034) );
  OAI21_X1 U13533 ( .B1(n15347), .B2(n9219), .A(n11034), .ZN(P2_U3451) );
  NAND2_X1 U13534 ( .A1(n11035), .A2(n15357), .ZN(n11036) );
  OAI21_X1 U13535 ( .B1(n15357), .B2(n10092), .A(n11036), .ZN(P2_U3506) );
  OAI222_X1 U13536 ( .A1(P3_U3151), .A2(n11039), .B1(n13690), .B2(n11038), 
        .C1(n13688), .C2(n11037), .ZN(P3_U3275) );
  INV_X1 U13537 ( .A(n13265), .ZN(n13237) );
  NAND2_X1 U13538 ( .A1(n13237), .A2(n6667), .ZN(n11040) );
  OAI21_X1 U13539 ( .B1(n6667), .B2(n11041), .A(n11040), .ZN(P3_U3515) );
  AOI21_X1 U13540 ( .B1(n15604), .B2(n11043), .A(n11042), .ZN(n11059) );
  AOI21_X1 U13541 ( .B1(n11533), .B2(n11045), .A(n11044), .ZN(n11052) );
  INV_X1 U13542 ( .A(n11046), .ZN(n11047) );
  NAND2_X1 U13543 ( .A1(n11048), .A2(n11047), .ZN(n11049) );
  XNOR2_X1 U13544 ( .A(n11050), .B(n11049), .ZN(n11051) );
  OAI22_X1 U13545 ( .A1(n11052), .A2(n15530), .B1(n7858), .B2(n11051), .ZN(
        n11053) );
  INV_X1 U13546 ( .A(n11053), .ZN(n11058) );
  AND2_X1 U13547 ( .A1(P3_U3151), .A2(P3_REG3_REG_9__SCAN_IN), .ZN(n11056) );
  NOR2_X1 U13548 ( .A1(n15520), .A2(n11054), .ZN(n11055) );
  AOI211_X1 U13549 ( .C1(n15523), .C2(P3_ADDR_REG_9__SCAN_IN), .A(n11056), .B(
        n11055), .ZN(n11057) );
  OAI211_X1 U13550 ( .C1(n11059), .C2(n15516), .A(n11058), .B(n11057), .ZN(
        P3_U3191) );
  AND2_X1 U13551 ( .A1(n15335), .A2(n13962), .ZN(n11061) );
  OAI21_X1 U13552 ( .B1(n15291), .B2(n11061), .A(n11060), .ZN(n15293) );
  OR2_X1 U13553 ( .A1(n11474), .A2(n11062), .ZN(n15292) );
  NOR2_X1 U13554 ( .A1(n15292), .A2(n11063), .ZN(n11064) );
  NOR2_X1 U13555 ( .A1(n15293), .A2(n11064), .ZN(n11066) );
  OAI22_X1 U13556 ( .A1(n15269), .A2(n11066), .B1(n11065), .B2(n14086), .ZN(
        n11067) );
  AOI21_X1 U13557 ( .B1(n15269), .B2(P2_REG2_REG_0__SCAN_IN), .A(n11067), .ZN(
        n11068) );
  OAI21_X1 U13558 ( .B1(n15291), .B2(n11659), .A(n11068), .ZN(P2_U3265) );
  INV_X1 U13559 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n11082) );
  XNOR2_X1 U13560 ( .A(n11070), .B(n11069), .ZN(n11248) );
  INV_X1 U13561 ( .A(n11170), .ZN(n11071) );
  AOI211_X1 U13562 ( .C1(n11215), .C2(n11072), .A(n14091), .B(n11071), .ZN(
        n11251) );
  AOI21_X1 U13563 ( .B1(n15313), .B2(n11215), .A(n11251), .ZN(n11080) );
  XNOR2_X1 U13564 ( .A(n11074), .B(n11073), .ZN(n11079) );
  OR2_X1 U13565 ( .A1(n13839), .A2(n11075), .ZN(n11077) );
  NAND2_X1 U13566 ( .A1(n13852), .A2(n13882), .ZN(n11076) );
  AND2_X1 U13567 ( .A1(n11077), .A2(n11076), .ZN(n11213) );
  INV_X1 U13568 ( .A(n11213), .ZN(n11078) );
  AOI21_X1 U13569 ( .B1(n11079), .B2(n14065), .A(n11078), .ZN(n11253) );
  OAI211_X1 U13570 ( .C1(n15000), .C2(n11248), .A(n11080), .B(n11253), .ZN(
        n11104) );
  NAND2_X1 U13571 ( .A1(n11104), .A2(n15347), .ZN(n11081) );
  OAI21_X1 U13572 ( .B1(n15347), .B2(n11082), .A(n11081), .ZN(P2_U3454) );
  INV_X1 U13573 ( .A(n11747), .ZN(n11103) );
  NAND2_X1 U13574 ( .A1(n11084), .A2(n11083), .ZN(n11085) );
  XNOR2_X1 U13575 ( .A(n12432), .B(n15545), .ZN(n11182) );
  XNOR2_X1 U13576 ( .A(n11182), .B(n11543), .ZN(n11095) );
  NAND2_X1 U13577 ( .A1(n11088), .A2(n8952), .ZN(n11089) );
  XNOR2_X1 U13578 ( .A(n11090), .B(n11304), .ZN(n15382) );
  INV_X1 U13579 ( .A(n11090), .ZN(n11092) );
  NAND2_X1 U13580 ( .A1(n11092), .A2(n11091), .ZN(n11093) );
  OAI21_X1 U13581 ( .B1(n11095), .B2(n11094), .A(n11184), .ZN(n11096) );
  NAND2_X1 U13582 ( .A1(n11096), .A2(n15390), .ZN(n11102) );
  INV_X1 U13583 ( .A(n15393), .ZN(n15370) );
  OR2_X1 U13584 ( .A1(n11304), .A2(n13518), .ZN(n11098) );
  OR2_X1 U13585 ( .A1(n11767), .A2(n13520), .ZN(n11097) );
  AND2_X1 U13586 ( .A1(n11098), .A2(n11097), .ZN(n11744) );
  OAI22_X1 U13587 ( .A1(n15370), .A2(n11744), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n11099), .ZN(n11100) );
  AOI21_X1 U13588 ( .B1(n15545), .B2(n15377), .A(n11100), .ZN(n11101) );
  OAI211_X1 U13589 ( .C1(n11103), .C2(n15401), .A(n11102), .B(n11101), .ZN(
        P3_U3170) );
  NAND2_X1 U13590 ( .A1(n11104), .A2(n15357), .ZN(n11105) );
  OAI21_X1 U13591 ( .B1(n15357), .B2(n10093), .A(n11105), .ZN(P2_U3507) );
  INV_X1 U13592 ( .A(n13268), .ZN(n13302) );
  NAND2_X1 U13593 ( .A1(n13302), .A2(n6667), .ZN(n11106) );
  OAI21_X1 U13594 ( .B1(n6667), .B2(n11107), .A(n11106), .ZN(P3_U3516) );
  NAND2_X1 U13595 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), 
        .ZN(n11108) );
  NAND2_X1 U13596 ( .A1(n11109), .A2(n11108), .ZN(n11111) );
  INV_X1 U13597 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n11110) );
  XNOR2_X1 U13598 ( .A(n11111), .B(n11110), .ZN(n14474) );
  OAI222_X1 U13599 ( .A1(n14876), .A2(n11112), .B1(P1_U3086), .B2(n6818), .C1(
        n12659), .C2(n14874), .ZN(P1_U3337) );
  INV_X1 U13600 ( .A(n13897), .ZN(n12351) );
  OAI222_X1 U13601 ( .A1(P2_U3088), .A2(n12351), .B1(n14196), .B2(n12659), 
        .C1(n11113), .C2(n14201), .ZN(P2_U3309) );
  XNOR2_X1 U13602 ( .A(n11114), .B(n11119), .ZN(n15325) );
  INV_X1 U13603 ( .A(n11140), .ZN(n11115) );
  AOI211_X1 U13604 ( .C1(n11116), .C2(n11296), .A(n14091), .B(n11115), .ZN(
        n15322) );
  OAI22_X1 U13605 ( .A1(n14094), .A2(n7049), .B1(n11117), .B2(n14086), .ZN(
        n11118) );
  AOI21_X1 U13606 ( .B1(n15279), .B2(n15322), .A(n11118), .ZN(n11126) );
  XNOR2_X1 U13607 ( .A(n11120), .B(n11119), .ZN(n11123) );
  INV_X1 U13608 ( .A(n11121), .ZN(n11122) );
  AOI21_X1 U13609 ( .B1(n11123), .B2(n14065), .A(n11122), .ZN(n15323) );
  MUX2_X1 U13610 ( .A(n11124), .B(n15323), .S(n14088), .Z(n11125) );
  OAI211_X1 U13611 ( .C1(n14099), .C2(n15325), .A(n11126), .B(n11125), .ZN(
        P2_U3261) );
  MUX2_X1 U13612 ( .A(n11128), .B(n11127), .S(n14088), .Z(n11134) );
  OAI22_X1 U13613 ( .A1(n14094), .A2(n11130), .B1(n14086), .B2(n11129), .ZN(
        n11131) );
  AOI21_X1 U13614 ( .B1(n11132), .B2(n15279), .A(n11131), .ZN(n11133) );
  OAI211_X1 U13615 ( .C1(n14099), .C2(n11135), .A(n11134), .B(n11133), .ZN(
        P2_U3259) );
  OAI222_X1 U13616 ( .A1(P3_U3151), .A2(n11313), .B1(n13690), .B2(n11137), 
        .C1(n13688), .C2(n11136), .ZN(P3_U3274) );
  XNOR2_X1 U13617 ( .A(n11138), .B(n11144), .ZN(n15333) );
  AOI211_X1 U13618 ( .C1(n11141), .C2(n11140), .A(n14091), .B(n11139), .ZN(
        n15329) );
  OAI22_X1 U13619 ( .A1(n14094), .A2(n15332), .B1(n14086), .B2(n11142), .ZN(
        n11143) );
  AOI21_X1 U13620 ( .B1(n15329), .B2(n15279), .A(n11143), .ZN(n11151) );
  XNOR2_X1 U13621 ( .A(n11145), .B(n11144), .ZN(n11148) );
  INV_X1 U13622 ( .A(n11146), .ZN(n11147) );
  AOI21_X1 U13623 ( .B1(n11148), .B2(n14065), .A(n11147), .ZN(n15330) );
  MUX2_X1 U13624 ( .A(n11149), .B(n15330), .S(n14088), .Z(n11150) );
  OAI211_X1 U13625 ( .C1(n14099), .C2(n15333), .A(n11151), .B(n11150), .ZN(
        P2_U3260) );
  AOI21_X1 U13626 ( .B1(n6791), .B2(n11153), .A(n11152), .ZN(n11167) );
  AOI21_X1 U13627 ( .B1(n6792), .B2(n11155), .A(n11154), .ZN(n11156) );
  OAI22_X1 U13628 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15368), .B1(n11156), .B2(
        n15530), .ZN(n11157) );
  INV_X1 U13629 ( .A(n11157), .ZN(n11166) );
  INV_X1 U13630 ( .A(P3_ADDR_REG_10__SCAN_IN), .ZN(n11162) );
  AOI21_X1 U13631 ( .B1(n11160), .B2(n11159), .A(n11158), .ZN(n11161) );
  OAI22_X1 U13632 ( .A1(n15492), .A2(n11162), .B1(n11161), .B2(n7858), .ZN(
        n11163) );
  AOI21_X1 U13633 ( .B1(n11164), .B2(n15485), .A(n11163), .ZN(n11165) );
  OAI211_X1 U13634 ( .C1(n11167), .C2(n15516), .A(n11166), .B(n11165), .ZN(
        P3_U3192) );
  XNOR2_X1 U13635 ( .A(n11169), .B(n11168), .ZN(n11256) );
  AOI211_X1 U13636 ( .C1(n11272), .C2(n11170), .A(n14091), .B(n11568), .ZN(
        n11259) );
  AOI21_X1 U13637 ( .B1(n15313), .B2(n11272), .A(n11259), .ZN(n11177) );
  XNOR2_X1 U13638 ( .A(n11172), .B(n11171), .ZN(n11176) );
  OR2_X1 U13639 ( .A1(n13839), .A2(n11198), .ZN(n11174) );
  NAND2_X1 U13640 ( .A1(n13852), .A2(n13881), .ZN(n11173) );
  AND2_X1 U13641 ( .A1(n11174), .A2(n11173), .ZN(n11276) );
  INV_X1 U13642 ( .A(n11276), .ZN(n11175) );
  AOI21_X1 U13643 ( .B1(n11176), .B2(n14065), .A(n11175), .ZN(n11261) );
  OAI211_X1 U13644 ( .C1(n15000), .C2(n11256), .A(n11177), .B(n11261), .ZN(
        n11179) );
  NAND2_X1 U13645 ( .A1(n11179), .A2(n15347), .ZN(n11178) );
  OAI21_X1 U13646 ( .B1(n15347), .B2(n9260), .A(n11178), .ZN(P2_U3457) );
  NAND2_X1 U13647 ( .A1(n11179), .A2(n15357), .ZN(n11180) );
  OAI21_X1 U13648 ( .B1(n15357), .B2(n10097), .A(n11180), .ZN(P2_U3508) );
  XNOR2_X1 U13649 ( .A(n12432), .B(n11550), .ZN(n11709) );
  XNOR2_X1 U13650 ( .A(n11181), .B(n11709), .ZN(n11710) );
  NAND2_X1 U13651 ( .A1(n11182), .A2(n11755), .ZN(n11183) );
  XOR2_X1 U13652 ( .A(n11711), .B(n11710), .Z(n11188) );
  INV_X1 U13653 ( .A(n15377), .ZN(n15397) );
  OAI22_X1 U13654 ( .A1(n15397), .A2(n15550), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n8092), .ZN(n11186) );
  OAI22_X1 U13655 ( .A1(n11755), .A2(n13295), .B1(n13315), .B2(n11942), .ZN(
        n11185) );
  AOI211_X1 U13656 ( .C1(n13319), .C2(n11549), .A(n11186), .B(n11185), .ZN(
        n11187) );
  OAI21_X1 U13657 ( .B1(n11188), .B2(n15381), .A(n11187), .ZN(P3_U3167) );
  INV_X1 U13658 ( .A(n11189), .ZN(n11192) );
  OAI22_X1 U13659 ( .A1(n11190), .A2(P3_U3151), .B1(SI_22_), .B2(n13690), .ZN(
        n11191) );
  AOI21_X1 U13660 ( .B1(n11192), .B2(n13681), .A(n11191), .ZN(P3_U3273) );
  OAI222_X1 U13661 ( .A1(n14876), .A2(n12708), .B1(n11283), .B2(n12707), .C1(
        n12478), .C2(P1_U3086), .ZN(P1_U3335) );
  INV_X1 U13662 ( .A(n11193), .ZN(n11194) );
  NAND2_X1 U13663 ( .A1(n11195), .A2(n11194), .ZN(n11196) );
  XNOR2_X1 U13664 ( .A(n11247), .B(n13734), .ZN(n11199) );
  OR2_X1 U13665 ( .A1(n10697), .A2(n11198), .ZN(n11200) );
  NAND2_X1 U13666 ( .A1(n11199), .A2(n11200), .ZN(n11208) );
  INV_X1 U13667 ( .A(n11199), .ZN(n11202) );
  INV_X1 U13668 ( .A(n11200), .ZN(n11201) );
  NAND2_X1 U13669 ( .A1(n11202), .A2(n11201), .ZN(n11204) );
  INV_X1 U13670 ( .A(n11273), .ZN(n11209) );
  INV_X1 U13671 ( .A(n11203), .ZN(n11205) );
  NAND2_X1 U13672 ( .A1(n11205), .A2(n11204), .ZN(n11207) );
  AOI22_X1 U13673 ( .A1(n11209), .A2(n11208), .B1(n11207), .B2(n11206), .ZN(
        n11217) );
  INV_X1 U13674 ( .A(n11210), .ZN(n11245) );
  NAND2_X1 U13675 ( .A1(n13853), .A2(n11245), .ZN(n11212) );
  OAI211_X1 U13676 ( .C1(n11213), .C2(n13855), .A(n11212), .B(n11211), .ZN(
        n11214) );
  AOI21_X1 U13677 ( .B1(n11215), .B2(n13857), .A(n11214), .ZN(n11216) );
  OAI21_X1 U13678 ( .B1(n11217), .B2(n13859), .A(n11216), .ZN(P2_U3193) );
  NAND2_X1 U13679 ( .A1(n13238), .A2(n6667), .ZN(n11218) );
  OAI21_X1 U13680 ( .B1(P3_U3897), .B2(n11219), .A(n11218), .ZN(P3_U3517) );
  OAI222_X1 U13681 ( .A1(n14876), .A2(n12723), .B1(n14874), .B2(n12722), .C1(
        n12486), .C2(P1_U3086), .ZN(P1_U3334) );
  INV_X2 U13682 ( .A(n11858), .ZN(n13086) );
  OR2_X1 U13683 ( .A1(n12820), .A2(n11220), .ZN(n11223) );
  OR2_X1 U13684 ( .A1(n12721), .A2(n11221), .ZN(n11222) );
  AOI22_X1 U13685 ( .A1(n14375), .A2(n13038), .B1(n13086), .B2(n12555), .ZN(
        n11225) );
  XOR2_X1 U13686 ( .A(n10886), .B(n11225), .Z(n11411) );
  AND2_X1 U13687 ( .A1(n12555), .A2(n13085), .ZN(n11226) );
  AOI21_X1 U13688 ( .B1(n14375), .B2(n13087), .A(n11226), .ZN(n11408) );
  INV_X1 U13689 ( .A(n11227), .ZN(n11229) );
  OAI21_X1 U13690 ( .B1(n11230), .B2(n11229), .A(n11228), .ZN(n11409) );
  XOR2_X1 U13691 ( .A(n11408), .B(n11409), .Z(n11412) );
  XOR2_X1 U13692 ( .A(n11411), .B(n11412), .Z(n11244) );
  INV_X1 U13693 ( .A(n11798), .ZN(n11242) );
  NAND2_X1 U13694 ( .A1(n14376), .A2(n14620), .ZN(n11239) );
  AOI21_X1 U13695 ( .B1(P1_REG3_REG_4__SCAN_IN), .B2(P1_REG3_REG_3__SCAN_IN), 
        .A(P1_REG3_REG_5__SCAN_IN), .ZN(n11231) );
  NOR2_X1 U13696 ( .A1(n11231), .A2(n11331), .ZN(n15130) );
  NAND2_X1 U13697 ( .A1(n12810), .A2(n15130), .ZN(n11237) );
  OR2_X1 U13698 ( .A1(n12664), .A2(n11232), .ZN(n11236) );
  OR2_X1 U13699 ( .A1(n12670), .A2(n11509), .ZN(n11235) );
  INV_X1 U13700 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n11233) );
  OR2_X1 U13701 ( .A1(n10990), .A2(n11233), .ZN(n11234) );
  NAND4_X1 U13702 ( .A1(n11237), .A2(n11236), .A3(n11235), .A4(n11234), .ZN(
        n14374) );
  NAND2_X1 U13703 ( .A1(n14374), .A2(n14771), .ZN(n11238) );
  NAND2_X1 U13704 ( .A1(n11239), .A2(n11238), .ZN(n11795) );
  AOI22_X1 U13705 ( .A1(n14349), .A2(n11795), .B1(P1_REG3_REG_4__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11240) );
  OAI21_X1 U13706 ( .B1(n14352), .B2(n11797), .A(n11240), .ZN(n11241) );
  AOI21_X1 U13707 ( .B1(n11242), .B2(n14338), .A(n11241), .ZN(n11243) );
  OAI21_X1 U13708 ( .B1(n11244), .B2(n15062), .A(n11243), .ZN(P1_U3230) );
  AOI22_X1 U13709 ( .A1(n15269), .A2(P2_REG2_REG_8__SCAN_IN), .B1(n11245), 
        .B2(n15268), .ZN(n11246) );
  OAI21_X1 U13710 ( .B1(n14094), .B2(n11247), .A(n11246), .ZN(n11250) );
  NOR2_X1 U13711 ( .A1(n11248), .A2(n14099), .ZN(n11249) );
  AOI211_X1 U13712 ( .C1(n11251), .C2(n15279), .A(n11250), .B(n11249), .ZN(
        n11252) );
  OAI21_X1 U13713 ( .B1(n14078), .B2(n11253), .A(n11252), .ZN(P2_U3257) );
  INV_X1 U13714 ( .A(n11254), .ZN(n11280) );
  AOI22_X1 U13715 ( .A1(n15269), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n11280), 
        .B2(n15268), .ZN(n11255) );
  OAI21_X1 U13716 ( .B1(n14094), .B2(n11277), .A(n11255), .ZN(n11258) );
  NOR2_X1 U13717 ( .A1(n11256), .A2(n14099), .ZN(n11257) );
  AOI211_X1 U13718 ( .C1(n11259), .C2(n15279), .A(n11258), .B(n11257), .ZN(
        n11260) );
  OAI21_X1 U13719 ( .B1(n14078), .B2(n11261), .A(n11260), .ZN(P2_U3256) );
  INV_X1 U13720 ( .A(n11262), .ZN(n11263) );
  AOI22_X1 U13721 ( .A1(n15269), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n11263), 
        .B2(n15268), .ZN(n11264) );
  OAI21_X1 U13722 ( .B1(n14094), .B2(n11265), .A(n11264), .ZN(n11268) );
  NOR2_X1 U13723 ( .A1(n11266), .A2(n14099), .ZN(n11267) );
  AOI211_X1 U13724 ( .C1(n11269), .C2(n15279), .A(n11268), .B(n11267), .ZN(
        n11270) );
  OAI21_X1 U13725 ( .B1(n14078), .B2(n11271), .A(n11270), .ZN(P2_U3258) );
  XNOR2_X1 U13726 ( .A(n11272), .B(n10727), .ZN(n11449) );
  NAND2_X1 U13727 ( .A1(n10734), .A2(n13882), .ZN(n11448) );
  XNOR2_X1 U13728 ( .A(n11449), .B(n11448), .ZN(n11274) );
  AOI21_X1 U13729 ( .B1(n11274), .B2(n11273), .A(n11450), .ZN(n11282) );
  OAI22_X1 U13730 ( .A1(n13855), .A2(n11276), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11275), .ZN(n11279) );
  NOR2_X1 U13731 ( .A1(n13812), .A2(n11277), .ZN(n11278) );
  AOI211_X1 U13732 ( .C1(n13853), .C2(n11280), .A(n11279), .B(n11278), .ZN(
        n11281) );
  OAI21_X1 U13733 ( .B1(n11282), .B2(n13859), .A(n11281), .ZN(P2_U3203) );
  INV_X1 U13734 ( .A(n12649), .ZN(n11285) );
  OAI222_X1 U13735 ( .A1(n14876), .A2(n11284), .B1(n11283), .B2(n11285), .C1(
        P1_U3086), .C2(n12475), .ZN(P1_U3336) );
  OAI222_X1 U13736 ( .A1(n14201), .A2(n11286), .B1(n14196), .B2(n11285), .C1(
        n9758), .C2(P2_U3088), .ZN(P2_U3308) );
  OAI222_X1 U13737 ( .A1(n14201), .A2(n7203), .B1(P2_U3088), .B2(n11287), .C1(
        n14196), .C2(n12707), .ZN(P2_U3307) );
  XNOR2_X1 U13738 ( .A(n11289), .B(n11288), .ZN(n15317) );
  XNOR2_X1 U13739 ( .A(n11290), .B(n11291), .ZN(n11294) );
  OR2_X1 U13740 ( .A1(n13839), .A2(n9722), .ZN(n11293) );
  NAND2_X1 U13741 ( .A1(n13852), .A2(n13888), .ZN(n11292) );
  NAND2_X1 U13742 ( .A1(n11293), .A2(n11292), .ZN(n13748) );
  AOI21_X1 U13743 ( .B1(n11294), .B2(n14065), .A(n13748), .ZN(n15321) );
  OAI21_X1 U13744 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(n14086), .A(n15321), .ZN(
        n11295) );
  MUX2_X1 U13745 ( .A(n11295), .B(P2_REG2_REG_3__SCAN_IN), .S(n14078), .Z(
        n11299) );
  OAI211_X1 U13746 ( .C1(n15277), .C2(n11297), .A(n15274), .B(n11296), .ZN(
        n15316) );
  OAI22_X1 U13747 ( .A1(n14026), .A2(n15316), .B1(n11297), .B2(n14094), .ZN(
        n11298) );
  AOI211_X1 U13748 ( .C1(n15317), .C2(n15280), .A(n11299), .B(n11298), .ZN(
        n11300) );
  INV_X1 U13749 ( .A(n11300), .ZN(P2_U3262) );
  INV_X1 U13750 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n11318) );
  XNOR2_X1 U13751 ( .A(n11301), .B(n11303), .ZN(n11315) );
  XNOR2_X1 U13752 ( .A(n11303), .B(n11302), .ZN(n11307) );
  OAI22_X1 U13753 ( .A1(n11305), .A2(n13518), .B1(n11304), .B2(n13520), .ZN(
        n11306) );
  AOI21_X1 U13754 ( .B1(n11307), .B2(n13552), .A(n11306), .ZN(n11308) );
  OAI21_X1 U13755 ( .B1(n15557), .B2(n11315), .A(n11308), .ZN(n15533) );
  NAND2_X1 U13756 ( .A1(n11309), .A2(n15561), .ZN(n15532) );
  OAI22_X1 U13757 ( .A1(n13538), .A2(n11311), .B1(n11310), .B2(n15532), .ZN(
        n11312) );
  OAI21_X1 U13758 ( .B1(n15533), .B2(n11312), .A(n13541), .ZN(n11317) );
  OR2_X1 U13759 ( .A1(n11314), .A2(n11313), .ZN(n11660) );
  NOR2_X1 U13760 ( .A1(n13560), .A2(n11660), .ZN(n13464) );
  INV_X1 U13761 ( .A(n11315), .ZN(n15535) );
  NAND2_X1 U13762 ( .A1(n13464), .A2(n15535), .ZN(n11316) );
  OAI211_X1 U13763 ( .C1(n11318), .C2(n13541), .A(n11317), .B(n11316), .ZN(
        P3_U3231) );
  NAND2_X1 U13764 ( .A1(n11355), .A2(n12530), .ZN(n11319) );
  OR2_X1 U13765 ( .A1(n11320), .A2(n11786), .ZN(n11421) );
  NAND2_X1 U13766 ( .A1(n14377), .A2(n11434), .ZN(n11321) );
  NAND2_X1 U13767 ( .A1(n11432), .A2(n11322), .ZN(n11489) );
  NAND2_X1 U13768 ( .A1(n11489), .A2(n11490), .ZN(n11488) );
  OR2_X1 U13769 ( .A1(n14376), .A2(n15139), .ZN(n11323) );
  NAND2_X1 U13770 ( .A1(n11488), .A2(n11323), .ZN(n11480) );
  NAND2_X1 U13771 ( .A1(n11480), .A2(n11479), .ZN(n11478) );
  OR2_X1 U13772 ( .A1(n14375), .A2(n12555), .ZN(n11324) );
  NAND2_X1 U13773 ( .A1(n11478), .A2(n11324), .ZN(n11501) );
  NAND2_X1 U13774 ( .A1(n12819), .A2(n11325), .ZN(n11328) );
  OR2_X1 U13775 ( .A1(n12820), .A2(n11326), .ZN(n11327) );
  OAI211_X1 U13776 ( .C1(n12738), .C2(n11329), .A(n11328), .B(n11327), .ZN(
        n15131) );
  XNOR2_X1 U13777 ( .A(n14374), .B(n11582), .ZN(n12843) );
  NAND2_X1 U13778 ( .A1(n11501), .A2(n12843), .ZN(n11500) );
  OR2_X1 U13779 ( .A1(n14374), .A2(n15131), .ZN(n11330) );
  NAND2_X1 U13780 ( .A1(n11500), .A2(n11330), .ZN(n11342) );
  NAND2_X1 U13781 ( .A1(n12811), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n11336) );
  INV_X1 U13782 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n11367) );
  OR2_X1 U13783 ( .A1(n12664), .A2(n11367), .ZN(n11335) );
  OAI21_X1 U13784 ( .B1(n11331), .B2(P1_REG3_REG_6__SCAN_IN), .A(n11386), .ZN(
        n14323) );
  OR2_X1 U13785 ( .A1(n12786), .A2(n14323), .ZN(n11334) );
  INV_X1 U13786 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n11332) );
  OR2_X1 U13787 ( .A1(n10990), .A2(n11332), .ZN(n11333) );
  NAND4_X1 U13788 ( .A1(n11336), .A2(n11335), .A3(n11334), .A4(n11333), .ZN(
        n14373) );
  INV_X2 U13789 ( .A(n12820), .ZN(n12661) );
  AOI22_X1 U13790 ( .A1(n12661), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n12660), 
        .B2(n11337), .ZN(n11340) );
  OR2_X1 U13791 ( .A1(n11338), .A2(n12721), .ZN(n11339) );
  INV_X1 U13792 ( .A(n15158), .ZN(n11370) );
  OR2_X1 U13793 ( .A1(n14373), .A2(n11370), .ZN(n11394) );
  NAND2_X1 U13794 ( .A1(n14373), .A2(n11370), .ZN(n11341) );
  NAND2_X1 U13795 ( .A1(n11394), .A2(n11341), .ZN(n12838) );
  NAND2_X1 U13796 ( .A1(n11342), .A2(n12838), .ZN(n11377) );
  OAI21_X1 U13797 ( .B1(n11342), .B2(n12838), .A(n11377), .ZN(n11366) );
  INV_X1 U13798 ( .A(n11366), .ZN(n15162) );
  INV_X1 U13799 ( .A(n11514), .ZN(n11346) );
  INV_X1 U13800 ( .A(n11343), .ZN(n11344) );
  NAND3_X1 U13801 ( .A1(n11346), .A2(n11345), .A3(n11344), .ZN(n13103) );
  NAND2_X1 U13802 ( .A1(n12540), .A2(n14483), .ZN(n12482) );
  OR2_X1 U13803 ( .A1(n15143), .A2(n12482), .ZN(n14673) );
  INV_X1 U13804 ( .A(n11347), .ZN(n14665) );
  INV_X1 U13805 ( .A(n14374), .ZN(n11354) );
  INV_X1 U13806 ( .A(n14620), .ZN(n14700) );
  NAND2_X1 U13807 ( .A1(n12811), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n11353) );
  OR2_X1 U13808 ( .A1(n12664), .A2(n10396), .ZN(n11352) );
  INV_X1 U13809 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n11348) );
  XNOR2_X1 U13810 ( .A(n11386), .B(n11348), .ZN(n11874) );
  OR2_X1 U13811 ( .A1(n12753), .A2(n11874), .ZN(n11351) );
  INV_X1 U13812 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n11349) );
  OR2_X1 U13813 ( .A1(n10990), .A2(n11349), .ZN(n11350) );
  NAND4_X1 U13814 ( .A1(n11353), .A2(n11352), .A3(n11351), .A4(n11350), .ZN(
        n14372) );
  OAI22_X1 U13815 ( .A1(n11354), .A2(n14700), .B1(n12080), .B2(n14702), .ZN(
        n11365) );
  NAND2_X1 U13816 ( .A1(n11355), .A2(n11632), .ZN(n12546) );
  NAND2_X1 U13817 ( .A1(n12542), .A2(n12546), .ZN(n11437) );
  OR2_X1 U13818 ( .A1(n14376), .A2(n11578), .ZN(n11357) );
  INV_X1 U13819 ( .A(n11479), .ZN(n12841) );
  NAND2_X1 U13820 ( .A1(n11481), .A2(n12841), .ZN(n11359) );
  OR2_X1 U13821 ( .A1(n14375), .A2(n11797), .ZN(n11358) );
  NAND2_X1 U13822 ( .A1(n11359), .A2(n11358), .ZN(n11502) );
  NOR2_X1 U13823 ( .A1(n14374), .A2(n11582), .ZN(n11361) );
  NAND2_X1 U13824 ( .A1(n14374), .A2(n11582), .ZN(n11360) );
  OR2_X2 U13825 ( .A1(n11362), .A2(n12838), .ZN(n11395) );
  NAND2_X1 U13826 ( .A1(n11362), .A2(n12838), .ZN(n11363) );
  AOI21_X1 U13827 ( .B1(n11395), .B2(n11363), .A(n14699), .ZN(n11364) );
  AOI211_X1 U13828 ( .C1(n14665), .C2(n11366), .A(n11365), .B(n11364), .ZN(
        n15160) );
  INV_X2 U13829 ( .A(n15143), .ZN(n14708) );
  MUX2_X1 U13830 ( .A(n11367), .B(n15160), .S(n14708), .Z(n11373) );
  NAND2_X1 U13831 ( .A1(n11507), .A2(n11582), .ZN(n11506) );
  AOI21_X1 U13832 ( .B1(n11506), .B2(n15158), .A(n14781), .ZN(n11368) );
  AND2_X1 U13833 ( .A1(n11368), .A2(n11400), .ZN(n15156) );
  OR2_X1 U13834 ( .A1(n13103), .A2(n14483), .ZN(n15146) );
  OAI22_X1 U13835 ( .A1(n14709), .A2(n11370), .B1(n14323), .B2(n14706), .ZN(
        n11371) );
  AOI21_X1 U13836 ( .B1(n15156), .B2(n14713), .A(n11371), .ZN(n11372) );
  OAI211_X1 U13837 ( .C1(n15162), .C2(n14673), .A(n11373), .B(n11372), .ZN(
        P1_U3287) );
  NAND2_X1 U13838 ( .A1(n13329), .A2(P3_DATAO_REG_30__SCAN_IN), .ZN(n11374) );
  OAI21_X1 U13839 ( .B1(n11375), .B2(n13329), .A(n11374), .ZN(P3_U3521) );
  OR2_X1 U13840 ( .A1(n14373), .A2(n15158), .ZN(n11376) );
  NAND2_X1 U13841 ( .A1(n11377), .A2(n11376), .ZN(n11382) );
  NAND2_X1 U13842 ( .A1(n11378), .A2(n12819), .ZN(n11381) );
  AOI22_X1 U13843 ( .A1(n12661), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n12660), 
        .B2(n11379), .ZN(n11380) );
  XNOR2_X1 U13844 ( .A(n12080), .B(n12577), .ZN(n12844) );
  NAND2_X1 U13845 ( .A1(n11382), .A2(n12844), .ZN(n11700) );
  OAI21_X1 U13846 ( .B1(n11382), .B2(n12844), .A(n11700), .ZN(n11621) );
  INV_X1 U13847 ( .A(n11621), .ZN(n11404) );
  INV_X1 U13848 ( .A(n14373), .ZN(n11873) );
  NAND2_X1 U13849 ( .A1(n12702), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n11391) );
  OR2_X1 U13850 ( .A1(n12670), .A2(n11383), .ZN(n11390) );
  OR2_X1 U13851 ( .A1(n12664), .A2(n11703), .ZN(n11389) );
  INV_X1 U13852 ( .A(n11386), .ZN(n11384) );
  AOI21_X1 U13853 ( .B1(n11384), .B2(P1_REG3_REG_7__SCAN_IN), .A(
        P1_REG3_REG_8__SCAN_IN), .ZN(n11387) );
  NAND2_X1 U13854 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_REG3_REG_7__SCAN_IN), 
        .ZN(n11385) );
  OR2_X1 U13855 ( .A1(n11387), .A2(n11690), .ZN(n12081) );
  OR2_X1 U13856 ( .A1(n12786), .A2(n12081), .ZN(n11388) );
  NAND4_X1 U13857 ( .A1(n11391), .A2(n11390), .A3(n11389), .A4(n11388), .ZN(
        n14371) );
  OAI22_X1 U13858 ( .A1(n11873), .A2(n14700), .B1(n12123), .B2(n14702), .ZN(
        n11399) );
  NAND2_X1 U13859 ( .A1(n11395), .A2(n11394), .ZN(n11393) );
  INV_X1 U13860 ( .A(n12844), .ZN(n11392) );
  CLKBUF_X1 U13861 ( .A(n11682), .Z(n11397) );
  NAND3_X1 U13862 ( .A1(n11395), .A2(n12844), .A3(n11394), .ZN(n11396) );
  AOI21_X1 U13863 ( .B1(n11397), .B2(n11396), .A(n14699), .ZN(n11398) );
  AOI211_X1 U13864 ( .C1(n14665), .C2(n11621), .A(n11399), .B(n11398), .ZN(
        n11618) );
  MUX2_X1 U13865 ( .A(n10396), .B(n11618), .S(n14708), .Z(n11403) );
  AOI211_X1 U13866 ( .C1(n12577), .C2(n11400), .A(n14781), .B(n11702), .ZN(
        n11620) );
  INV_X1 U13867 ( .A(n12577), .ZN(n11625) );
  OAI22_X1 U13868 ( .A1(n14709), .A2(n11625), .B1(n11874), .B2(n14706), .ZN(
        n11401) );
  AOI21_X1 U13869 ( .B1(n11620), .B2(n14713), .A(n11401), .ZN(n11402) );
  OAI211_X1 U13870 ( .C1(n11404), .C2(n14673), .A(n11403), .B(n11402), .ZN(
        P1_U3286) );
  NAND2_X1 U13871 ( .A1(n14374), .A2(n13085), .ZN(n11406) );
  NAND2_X1 U13872 ( .A1(n15131), .A2(n13086), .ZN(n11405) );
  NAND2_X1 U13873 ( .A1(n11406), .A2(n11405), .ZN(n11407) );
  XNOR2_X1 U13874 ( .A(n11407), .B(n10886), .ZN(n11860) );
  AOI22_X1 U13875 ( .A1(n14374), .A2(n13087), .B1(n13085), .B2(n15131), .ZN(
        n11861) );
  XNOR2_X1 U13876 ( .A(n11860), .B(n11861), .ZN(n11863) );
  INV_X1 U13877 ( .A(n11408), .ZN(n11410) );
  OAI22_X1 U13878 ( .A1(n11412), .A2(n11411), .B1(n11410), .B2(n11409), .ZN(
        n11864) );
  XOR2_X1 U13879 ( .A(n11863), .B(n11864), .Z(n11418) );
  NAND2_X1 U13880 ( .A1(n14375), .A2(n14620), .ZN(n11414) );
  NAND2_X1 U13881 ( .A1(n14373), .A2(n14771), .ZN(n11413) );
  NAND2_X1 U13882 ( .A1(n11414), .A2(n11413), .ZN(n11505) );
  AOI22_X1 U13883 ( .A1(n14349), .A2(n11505), .B1(P1_REG3_REG_5__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11415) );
  OAI21_X1 U13884 ( .B1(n14352), .B2(n11582), .A(n11415), .ZN(n11416) );
  AOI21_X1 U13885 ( .B1(n15130), .B2(n14338), .A(n11416), .ZN(n11417) );
  OAI21_X1 U13886 ( .B1(n11418), .B2(n15062), .A(n11417), .ZN(P1_U3227) );
  OAI21_X1 U13887 ( .B1(n11419), .B2(n11421), .A(n11420), .ZN(n11635) );
  INV_X1 U13888 ( .A(n14377), .ZN(n11631) );
  NAND2_X1 U13889 ( .A1(n11422), .A2(n12530), .ZN(n11423) );
  NAND2_X1 U13890 ( .A1(n11435), .A2(n11423), .ZN(n11630) );
  OAI22_X1 U13891 ( .A1(n11631), .A2(n14702), .B1(n11630), .B2(n14781), .ZN(
        n11429) );
  INV_X1 U13892 ( .A(n11419), .ZN(n11424) );
  AOI21_X1 U13893 ( .B1(n11424), .B2(n14380), .A(n14699), .ZN(n11427) );
  XOR2_X1 U13894 ( .A(n14378), .B(n11630), .Z(n11425) );
  OAI21_X1 U13895 ( .B1(n11425), .B2(n14699), .A(n11320), .ZN(n11426) );
  OAI21_X1 U13896 ( .B1(n11427), .B2(n14620), .A(n11426), .ZN(n11636) );
  INV_X1 U13897 ( .A(n11636), .ZN(n11428) );
  AOI211_X1 U13898 ( .C1(n15175), .C2(n11635), .A(n11429), .B(n11428), .ZN(
        n11520) );
  OAI22_X1 U13899 ( .A1(n14804), .A2(n11632), .B1(n15184), .B2(n10518), .ZN(
        n11430) );
  INV_X1 U13900 ( .A(n11430), .ZN(n11431) );
  OAI21_X1 U13901 ( .B1(n11520), .B2(n15181), .A(n11431), .ZN(P1_U3529) );
  OAI21_X1 U13902 ( .B1(n11433), .B2(n6859), .A(n11432), .ZN(n11610) );
  AOI21_X1 U13903 ( .B1(n11435), .B2(n11434), .A(n14781), .ZN(n11436) );
  AND2_X1 U13904 ( .A1(n11436), .A2(n11495), .ZN(n11606) );
  INV_X1 U13905 ( .A(n6859), .ZN(n12547) );
  XNOR2_X1 U13906 ( .A(n11437), .B(n12547), .ZN(n11439) );
  OAI21_X1 U13907 ( .B1(n11439), .B2(n14699), .A(n11438), .ZN(n11604) );
  AOI211_X1 U13908 ( .C1(n15175), .C2(n11610), .A(n11606), .B(n11604), .ZN(
        n11524) );
  OAI22_X1 U13909 ( .A1(n14804), .A2(n12533), .B1(n15184), .B2(n10632), .ZN(
        n11440) );
  INV_X1 U13910 ( .A(n11440), .ZN(n11441) );
  OAI21_X1 U13911 ( .B1(n11524), .B2(n15181), .A(n11441), .ZN(P1_U3530) );
  NAND2_X1 U13912 ( .A1(n13303), .A2(n6667), .ZN(n11442) );
  OAI21_X1 U13913 ( .B1(n6667), .B2(n11443), .A(n11442), .ZN(P3_U3518) );
  NAND2_X1 U13914 ( .A1(n11444), .A2(n13681), .ZN(n11446) );
  OAI211_X1 U13915 ( .C1(n11447), .C2(n13690), .A(n11446), .B(n11445), .ZN(
        P3_U3272) );
  XNOR2_X1 U13916 ( .A(n11571), .B(n13734), .ZN(n11451) );
  AND2_X1 U13917 ( .A1(n13735), .A2(n13881), .ZN(n11452) );
  NAND2_X1 U13918 ( .A1(n11451), .A2(n11452), .ZN(n11670) );
  INV_X1 U13919 ( .A(n11451), .ZN(n11454) );
  INV_X1 U13920 ( .A(n11452), .ZN(n11453) );
  NAND2_X1 U13921 ( .A1(n11454), .A2(n11453), .ZN(n11455) );
  AND2_X1 U13922 ( .A1(n11670), .A2(n11455), .ZN(n11456) );
  OAI211_X1 U13923 ( .C1(n11457), .C2(n11456), .A(n11671), .B(n6908), .ZN(
        n11465) );
  OR2_X1 U13924 ( .A1(n11587), .A2(n13841), .ZN(n11459) );
  NAND2_X1 U13925 ( .A1(n13851), .A2(n13882), .ZN(n11458) );
  AND2_X1 U13926 ( .A1(n11459), .A2(n11458), .ZN(n11564) );
  INV_X1 U13927 ( .A(n11566), .ZN(n11460) );
  NAND2_X1 U13928 ( .A1(n13853), .A2(n11460), .ZN(n11462) );
  OAI211_X1 U13929 ( .C1(n11564), .C2(n13855), .A(n11462), .B(n11461), .ZN(
        n11463) );
  AOI21_X1 U13930 ( .B1(n11571), .B2(n13857), .A(n11463), .ZN(n11464) );
  NAND2_X1 U13931 ( .A1(n11465), .A2(n11464), .ZN(P2_U3189) );
  XNOR2_X1 U13932 ( .A(n6826), .B(n11466), .ZN(n15297) );
  OAI21_X1 U13933 ( .B1(n11469), .B2(n6826), .A(n11467), .ZN(n11471) );
  AOI21_X1 U13934 ( .B1(n11471), .B2(n14065), .A(n11470), .ZN(n15299) );
  OAI22_X1 U13935 ( .A1(n15269), .A2(n15299), .B1(n11472), .B2(n14086), .ZN(
        n11476) );
  INV_X1 U13936 ( .A(n15275), .ZN(n11473) );
  OAI211_X1 U13937 ( .C1(n15300), .C2(n11474), .A(n11473), .B(n15274), .ZN(
        n15298) );
  OAI22_X1 U13938 ( .A1(n14026), .A2(n15298), .B1(n15300), .B2(n14094), .ZN(
        n11475) );
  AOI211_X1 U13939 ( .C1(P2_REG2_REG_1__SCAN_IN), .C2(n15269), .A(n11476), .B(
        n11475), .ZN(n11477) );
  OAI21_X1 U13940 ( .B1(n14099), .B2(n15297), .A(n11477), .ZN(P2_U3264) );
  OAI21_X1 U13941 ( .B1(n11480), .B2(n11479), .A(n11478), .ZN(n11802) );
  AOI211_X1 U13942 ( .C1(n12555), .C2(n11496), .A(n14781), .B(n11507), .ZN(
        n11796) );
  AOI211_X1 U13943 ( .C1(n11802), .C2(n15175), .A(n11795), .B(n11796), .ZN(
        n11484) );
  XNOR2_X1 U13944 ( .A(n12841), .B(n11482), .ZN(n11483) );
  NAND2_X1 U13945 ( .A1(n11483), .A2(n14618), .ZN(n11793) );
  NAND2_X1 U13946 ( .A1(n11484), .A2(n11793), .ZN(n11576) );
  OAI22_X1 U13947 ( .A1(n14804), .A2(n11797), .B1(n15184), .B2(n11485), .ZN(
        n11486) );
  AOI21_X1 U13948 ( .B1(n11576), .B2(n15184), .A(n11486), .ZN(n11487) );
  INV_X1 U13949 ( .A(n11487), .ZN(P1_U3532) );
  OAI21_X1 U13950 ( .B1(n11489), .B2(n11490), .A(n11488), .ZN(n15150) );
  INV_X1 U13951 ( .A(n15150), .ZN(n11497) );
  XNOR2_X1 U13952 ( .A(n11491), .B(n11490), .ZN(n11492) );
  NOR2_X1 U13953 ( .A1(n11492), .A2(n14699), .ZN(n11493) );
  AOI211_X1 U13954 ( .C1(n14665), .C2(n15150), .A(n11494), .B(n11493), .ZN(
        n15152) );
  OAI211_X1 U13955 ( .C1(n7032), .C2(n11578), .A(n14811), .B(n11496), .ZN(
        n15147) );
  OAI211_X1 U13956 ( .C1(n11497), .C2(n15161), .A(n15152), .B(n15147), .ZN(
        n11580) );
  OAI22_X1 U13957 ( .A1(n14804), .A2(n11578), .B1(n15184), .B2(n10833), .ZN(
        n11498) );
  AOI21_X1 U13958 ( .B1(n11580), .B2(n15184), .A(n11498), .ZN(n11499) );
  INV_X1 U13959 ( .A(n11499), .ZN(P1_U3531) );
  OAI21_X1 U13960 ( .B1(n11501), .B2(n12843), .A(n11500), .ZN(n15136) );
  INV_X1 U13961 ( .A(n15136), .ZN(n11508) );
  XNOR2_X1 U13962 ( .A(n11502), .B(n12843), .ZN(n11503) );
  NOR2_X1 U13963 ( .A1(n11503), .A2(n14699), .ZN(n11504) );
  AOI211_X1 U13964 ( .C1(n14665), .C2(n15136), .A(n11505), .B(n11504), .ZN(
        n15138) );
  OAI211_X1 U13965 ( .C1(n11507), .C2(n11582), .A(n11506), .B(n14811), .ZN(
        n15134) );
  OAI211_X1 U13966 ( .C1(n11508), .C2(n15161), .A(n15138), .B(n15134), .ZN(
        n11584) );
  OAI22_X1 U13967 ( .A1(n14804), .A2(n11582), .B1(n15184), .B2(n11509), .ZN(
        n11510) );
  AOI21_X1 U13968 ( .B1(n11584), .B2(n15184), .A(n11510), .ZN(n11511) );
  INV_X1 U13969 ( .A(n11511), .ZN(P1_U3533) );
  OAI222_X1 U13970 ( .A1(n14201), .A2(n11512), .B1(P2_U3088), .B2(n9664), .C1(
        n14196), .C2(n12722), .ZN(P2_U3306) );
  OR2_X1 U13971 ( .A1(n11514), .A2(n11513), .ZN(n11515) );
  NOR2_X4 U13972 ( .A1(n11516), .A2(n11515), .ZN(n14854) );
  INV_X1 U13973 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n11517) );
  OAI22_X1 U13974 ( .A1(n14858), .A2(n11632), .B1(n14854), .B2(n11517), .ZN(
        n11518) );
  INV_X1 U13975 ( .A(n11518), .ZN(n11519) );
  OAI21_X1 U13976 ( .B1(n11520), .B2(n15177), .A(n11519), .ZN(P1_U3462) );
  INV_X1 U13977 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n11521) );
  OAI22_X1 U13978 ( .A1(n14858), .A2(n12533), .B1(n14854), .B2(n11521), .ZN(
        n11522) );
  INV_X1 U13979 ( .A(n11522), .ZN(n11523) );
  OAI21_X1 U13980 ( .B1(n11524), .B2(n15177), .A(n11523), .ZN(P1_U3465) );
  XNOR2_X1 U13981 ( .A(n11526), .B(n7108), .ZN(n11530) );
  OAI211_X1 U13982 ( .C1(n6794), .C2(n7108), .A(n13552), .B(n11527), .ZN(
        n11529) );
  AOI22_X1 U13983 ( .A1(n13531), .A2(n12004), .B1(n13324), .B2(n13533), .ZN(
        n11528) );
  OAI211_X1 U13984 ( .C1(n15557), .C2(n11530), .A(n11529), .B(n11528), .ZN(
        n15576) );
  INV_X1 U13985 ( .A(n15576), .ZN(n11536) );
  INV_X1 U13986 ( .A(n11530), .ZN(n15579) );
  AOI22_X1 U13987 ( .A1(n13543), .A2(n11531), .B1(n13559), .B2(n12016), .ZN(
        n11532) );
  OAI21_X1 U13988 ( .B1(n11533), .B2(n13541), .A(n11532), .ZN(n11534) );
  AOI21_X1 U13989 ( .B1(n15579), .B2(n13464), .A(n11534), .ZN(n11535) );
  OAI21_X1 U13990 ( .B1(n11536), .B2(n13566), .A(n11535), .ZN(P3_U3224) );
  NAND2_X1 U13991 ( .A1(n11756), .A2(n11537), .ZN(n11743) );
  NAND2_X1 U13992 ( .A1(n11743), .A2(n11742), .ZN(n11741) );
  NAND2_X1 U13993 ( .A1(n11741), .A2(n11538), .ZN(n11542) );
  NAND2_X1 U13994 ( .A1(n11540), .A2(n11539), .ZN(n11541) );
  AOI21_X1 U13995 ( .B1(n11544), .B2(n11542), .A(n11541), .ZN(n11548) );
  AOI22_X1 U13996 ( .A1(n13531), .A2(n11543), .B1(n13326), .B2(n13533), .ZN(
        n11547) );
  XNOR2_X1 U13997 ( .A(n11545), .B(n11544), .ZN(n15553) );
  INV_X1 U13998 ( .A(n15557), .ZN(n15588) );
  NAND2_X1 U13999 ( .A1(n15553), .A2(n15588), .ZN(n11546) );
  OAI211_X1 U14000 ( .C1(n11548), .C2(n13515), .A(n11547), .B(n11546), .ZN(
        n15551) );
  INV_X1 U14001 ( .A(n15551), .ZN(n11554) );
  AOI22_X1 U14002 ( .A1(n13543), .A2(n11550), .B1(n13559), .B2(n11549), .ZN(
        n11551) );
  OAI21_X1 U14003 ( .B1(n15424), .B2(n13541), .A(n11551), .ZN(n11552) );
  AOI21_X1 U14004 ( .B1(n15553), .B2(n13464), .A(n11552), .ZN(n11553) );
  OAI21_X1 U14005 ( .B1(n11554), .B2(n13566), .A(n11553), .ZN(P3_U3228) );
  OAI222_X1 U14006 ( .A1(n14201), .A2(n11557), .B1(P2_U3088), .B2(n11556), 
        .C1(n14196), .C2(n11555), .ZN(P2_U3305) );
  XOR2_X1 U14007 ( .A(n11558), .B(n11562), .Z(n15344) );
  INV_X1 U14008 ( .A(n15344), .ZN(n11574) );
  INV_X1 U14009 ( .A(n11559), .ZN(n11560) );
  AOI21_X1 U14010 ( .B1(n11562), .B2(n11561), .A(n11560), .ZN(n11565) );
  INV_X1 U14011 ( .A(n15335), .ZN(n15318) );
  NAND2_X1 U14012 ( .A1(n15344), .A2(n15318), .ZN(n11563) );
  OAI211_X1 U14013 ( .C1(n11565), .C2(n13962), .A(n11564), .B(n11563), .ZN(
        n15342) );
  NAND2_X1 U14014 ( .A1(n15342), .A2(n14088), .ZN(n11573) );
  OAI22_X1 U14015 ( .A1(n14088), .A2(n10053), .B1(n11566), .B2(n14086), .ZN(
        n11570) );
  INV_X1 U14016 ( .A(n11642), .ZN(n11567) );
  OAI211_X1 U14017 ( .C1(n15341), .C2(n11568), .A(n11567), .B(n15274), .ZN(
        n15339) );
  NOR2_X1 U14018 ( .A1(n15339), .A2(n14026), .ZN(n11569) );
  AOI211_X1 U14019 ( .C1(n15270), .C2(n11571), .A(n11570), .B(n11569), .ZN(
        n11572) );
  OAI211_X1 U14020 ( .C1(n11574), .C2(n11659), .A(n11573), .B(n11572), .ZN(
        P2_U3255) );
  OAI22_X1 U14021 ( .A1(n14858), .A2(n11797), .B1(n14854), .B2(n10991), .ZN(
        n11575) );
  AOI21_X1 U14022 ( .B1(n11576), .B2(n14854), .A(n11575), .ZN(n11577) );
  INV_X1 U14023 ( .A(n11577), .ZN(P1_U3471) );
  OAI22_X1 U14024 ( .A1(n14858), .A2(n11578), .B1(n14854), .B2(n10831), .ZN(
        n11579) );
  AOI21_X1 U14025 ( .B1(n11580), .B2(n14854), .A(n11579), .ZN(n11581) );
  INV_X1 U14026 ( .A(n11581), .ZN(P1_U3468) );
  OAI22_X1 U14027 ( .A1(n14858), .A2(n11582), .B1(n14854), .B2(n11233), .ZN(
        n11583) );
  AOI21_X1 U14028 ( .B1(n11584), .B2(n14854), .A(n11583), .ZN(n11585) );
  INV_X1 U14029 ( .A(n11585), .ZN(P1_U3474) );
  XNOR2_X1 U14030 ( .A(n11586), .B(n11591), .ZN(n11590) );
  OR2_X1 U14031 ( .A1(n13839), .A2(n11587), .ZN(n11588) );
  OAI21_X1 U14032 ( .B1(n11589), .B2(n13841), .A(n11588), .ZN(n11925) );
  AOI21_X1 U14033 ( .B1(n11590), .B2(n14065), .A(n11925), .ZN(n15030) );
  INV_X1 U14034 ( .A(n11591), .ZN(n11592) );
  XNOR2_X1 U14035 ( .A(n11593), .B(n11592), .ZN(n15028) );
  AOI21_X1 U14036 ( .B1(n11594), .B2(n11930), .A(n14091), .ZN(n11595) );
  NAND2_X1 U14037 ( .A1(n11595), .A2(n11885), .ZN(n15025) );
  OAI22_X1 U14038 ( .A1(n14088), .A2(n11596), .B1(n11928), .B2(n14086), .ZN(
        n11597) );
  AOI21_X1 U14039 ( .B1(n11930), .B2(n15270), .A(n11597), .ZN(n11598) );
  OAI21_X1 U14040 ( .B1(n15025), .B2(n14026), .A(n11598), .ZN(n11599) );
  AOI21_X1 U14041 ( .B1(n15028), .B2(n15280), .A(n11599), .ZN(n11600) );
  OAI21_X1 U14042 ( .B1(n15030), .B2(n14078), .A(n11600), .ZN(P2_U3253) );
  INV_X1 U14043 ( .A(P3_DATAO_REG_29__SCAN_IN), .ZN(n11603) );
  INV_X1 U14044 ( .A(n13219), .ZN(n11601) );
  NAND2_X1 U14045 ( .A1(n11601), .A2(n6667), .ZN(n11602) );
  OAI21_X1 U14046 ( .B1(P3_U3897), .B2(n11603), .A(n11602), .ZN(P3_U3520) );
  INV_X1 U14047 ( .A(n11604), .ZN(n11612) );
  INV_X1 U14048 ( .A(n14706), .ZN(n15142) );
  AOI22_X1 U14049 ( .A1(n14713), .A2(n11606), .B1(P1_REG3_REG_2__SCAN_IN), 
        .B2(n15142), .ZN(n11608) );
  NAND2_X1 U14050 ( .A1(n15143), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n11607) );
  OAI211_X1 U14051 ( .C1(n12533), .C2(n14709), .A(n11608), .B(n11607), .ZN(
        n11609) );
  AOI21_X1 U14052 ( .B1(n14649), .B2(n11610), .A(n11609), .ZN(n11611) );
  OAI21_X1 U14053 ( .B1(n15143), .B2(n11612), .A(n11611), .ZN(P1_U3291) );
  INV_X1 U14054 ( .A(n13420), .ZN(n11613) );
  NAND2_X1 U14055 ( .A1(n11613), .A2(n6667), .ZN(n11614) );
  OAI21_X1 U14056 ( .B1(P3_U3897), .B2(n11615), .A(n11614), .ZN(P3_U3519) );
  NAND2_X1 U14057 ( .A1(n7221), .A2(n6667), .ZN(n11616) );
  OAI21_X1 U14058 ( .B1(P3_U3897), .B2(n11617), .A(n11616), .ZN(P3_U3522) );
  INV_X1 U14059 ( .A(n15161), .ZN(n14910) );
  INV_X1 U14060 ( .A(n11618), .ZN(n11619) );
  AOI211_X1 U14061 ( .C1(n14910), .C2(n11621), .A(n11620), .B(n11619), .ZN(
        n11628) );
  OAI22_X1 U14062 ( .A1(n14804), .A2(n11625), .B1(n15184), .B2(n11622), .ZN(
        n11623) );
  INV_X1 U14063 ( .A(n11623), .ZN(n11624) );
  OAI21_X1 U14064 ( .B1(n11628), .B2(n15181), .A(n11624), .ZN(P1_U3535) );
  OAI22_X1 U14065 ( .A1(n14858), .A2(n11625), .B1(n14854), .B2(n11349), .ZN(
        n11626) );
  INV_X1 U14066 ( .A(n11626), .ZN(n11627) );
  OAI21_X1 U14067 ( .B1(n11628), .B2(n15177), .A(n11627), .ZN(P1_U3480) );
  NAND2_X1 U14068 ( .A1(n14713), .A2(n14811), .ZN(n14635) );
  OAI22_X1 U14069 ( .A1(n14635), .A2(n11630), .B1(n11629), .B2(n14706), .ZN(
        n11634) );
  OR2_X1 U14070 ( .A1(n15143), .A2(n14702), .ZN(n14606) );
  OAI22_X1 U14071 ( .A1(n11632), .A2(n14709), .B1(n14606), .B2(n11631), .ZN(
        n11633) );
  AOI211_X1 U14072 ( .C1(n14649), .C2(n11635), .A(n11634), .B(n11633), .ZN(
        n11639) );
  MUX2_X1 U14073 ( .A(n11637), .B(n11636), .S(n14708), .Z(n11638) );
  NAND2_X1 U14074 ( .A1(n11639), .A2(n11638), .ZN(P1_U3292) );
  XOR2_X1 U14075 ( .A(n11643), .B(n11640), .Z(n11912) );
  NOR2_X1 U14076 ( .A1(n11912), .A2(n11641), .ZN(n11654) );
  XNOR2_X1 U14077 ( .A(n11642), .B(n11680), .ZN(n11651) );
  INV_X1 U14078 ( .A(n11643), .ZN(n11645) );
  NAND3_X1 U14079 ( .A1(n11559), .A2(n11645), .A3(n11644), .ZN(n11646) );
  AOI21_X1 U14080 ( .B1(n11647), .B2(n11646), .A(n13962), .ZN(n11650) );
  OR2_X1 U14081 ( .A1(n11914), .A2(n13841), .ZN(n11649) );
  NAND2_X1 U14082 ( .A1(n13851), .A2(n13881), .ZN(n11648) );
  NAND2_X1 U14083 ( .A1(n11649), .A2(n11648), .ZN(n11677) );
  NOR2_X1 U14084 ( .A1(n11650), .A2(n11677), .ZN(n11652) );
  OAI21_X1 U14085 ( .B1(n14091), .B2(n11651), .A(n11652), .ZN(n11909) );
  OAI21_X1 U14086 ( .B1(n11652), .B2(n15269), .A(n14026), .ZN(n11653) );
  OAI21_X1 U14087 ( .B1(n11654), .B2(n11909), .A(n11653), .ZN(n11658) );
  OAI22_X1 U14088 ( .A1(n14088), .A2(n11655), .B1(n11674), .B2(n14086), .ZN(
        n11656) );
  AOI21_X1 U14089 ( .B1(n11910), .B2(n15270), .A(n11656), .ZN(n11657) );
  OAI211_X1 U14090 ( .C1(n11912), .C2(n11659), .A(n11658), .B(n11657), .ZN(
        P2_U3254) );
  AND2_X1 U14091 ( .A1(n15557), .A2(n11660), .ZN(n11661) );
  OAI21_X1 U14092 ( .B1(n8956), .B2(n11663), .A(n11662), .ZN(n11667) );
  OAI22_X1 U14093 ( .A1(n13541), .A2(n11665), .B1(n11664), .B2(n13538), .ZN(
        n11666) );
  AOI21_X1 U14094 ( .B1(n11667), .B2(n13541), .A(n11666), .ZN(n11668) );
  OAI21_X1 U14095 ( .B1(n13125), .B2(n11669), .A(n11668), .ZN(P3_U3232) );
  NAND2_X1 U14096 ( .A1(n11671), .A2(n11670), .ZN(n11673) );
  XNOR2_X1 U14097 ( .A(n11680), .B(n13734), .ZN(n11919) );
  AND2_X1 U14098 ( .A1(n13880), .A2(n13735), .ZN(n11920) );
  XNOR2_X1 U14099 ( .A(n11919), .B(n11920), .ZN(n11672) );
  OAI211_X1 U14100 ( .C1(n11673), .C2(n11672), .A(n11923), .B(n6908), .ZN(
        n11679) );
  NOR2_X1 U14101 ( .A1(n13845), .A2(n11674), .ZN(n11675) );
  AOI211_X1 U14102 ( .C1(n13843), .C2(n11677), .A(n11676), .B(n11675), .ZN(
        n11678) );
  OAI211_X1 U14103 ( .C1(n11680), .C2(n13812), .A(n11679), .B(n11678), .ZN(
        P2_U3208) );
  NAND2_X1 U14104 ( .A1(n12080), .A2(n12577), .ZN(n11681) );
  NAND2_X1 U14105 ( .A1(n11683), .A2(n12819), .ZN(n11686) );
  AOI22_X1 U14106 ( .A1(n12661), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n12660), 
        .B2(n11684), .ZN(n11685) );
  XNOR2_X1 U14107 ( .A(n12580), .B(n12123), .ZN(n12845) );
  AOI21_X1 U14108 ( .B1(n11687), .B2(n12845), .A(n14699), .ZN(n11698) );
  INV_X1 U14109 ( .A(n12845), .ZN(n11688) );
  NAND2_X1 U14110 ( .A1(n12812), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n11696) );
  OR2_X1 U14111 ( .A1(n12670), .A2(n10402), .ZN(n11695) );
  OR2_X1 U14112 ( .A1(n11690), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n11691) );
  NAND2_X1 U14113 ( .A1(n11982), .A2(n11691), .ZN(n12122) );
  OR2_X1 U14114 ( .A1(n12786), .A2(n12122), .ZN(n11694) );
  INV_X1 U14115 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11692) );
  OR2_X1 U14116 ( .A1(n10990), .A2(n11692), .ZN(n11693) );
  NAND4_X1 U14117 ( .A1(n11696), .A2(n11695), .A3(n11694), .A4(n11693), .ZN(
        n14370) );
  OAI22_X1 U14118 ( .A1(n12080), .A2(n14700), .B1(n12082), .B2(n14702), .ZN(
        n11697) );
  AOI21_X1 U14119 ( .B1(n11698), .B2(n11840), .A(n11697), .ZN(n15165) );
  OR2_X1 U14120 ( .A1(n12577), .A2(n14372), .ZN(n11699) );
  NAND2_X1 U14121 ( .A1(n11700), .A2(n11699), .ZN(n11701) );
  NAND2_X1 U14122 ( .A1(n11701), .A2(n12845), .ZN(n11833) );
  OAI21_X1 U14123 ( .B1(n11701), .B2(n12845), .A(n11833), .ZN(n15168) );
  INV_X1 U14124 ( .A(n12580), .ZN(n15166) );
  OAI211_X1 U14125 ( .C1(n15166), .C2(n11702), .A(n6692), .B(n14811), .ZN(
        n15164) );
  OAI22_X1 U14126 ( .A1(n14708), .A2(n11703), .B1(n12081), .B2(n14706), .ZN(
        n11704) );
  AOI21_X1 U14127 ( .B1(n15140), .B2(n12580), .A(n11704), .ZN(n11705) );
  OAI21_X1 U14128 ( .B1(n15164), .B2(n15146), .A(n11705), .ZN(n11706) );
  AOI21_X1 U14129 ( .B1(n15168), .B2(n14649), .A(n11706), .ZN(n11707) );
  OAI21_X1 U14130 ( .B1(n15143), .B2(n15165), .A(n11707), .ZN(P1_U3285) );
  INV_X1 U14131 ( .A(n11708), .ZN(n11781) );
  XNOR2_X1 U14132 ( .A(n12432), .B(n15398), .ZN(n11712) );
  XNOR2_X1 U14133 ( .A(n11712), .B(n11942), .ZN(n15392) );
  XNOR2_X1 U14134 ( .A(n11940), .B(n13174), .ZN(n15359) );
  INV_X1 U14135 ( .A(n15359), .ZN(n11715) );
  NAND2_X1 U14136 ( .A1(n11715), .A2(n11714), .ZN(n11716) );
  XNOR2_X1 U14137 ( .A(n12432), .B(n15569), .ZN(n12005) );
  XNOR2_X1 U14138 ( .A(n12005), .B(n12013), .ZN(n11717) );
  OAI211_X1 U14139 ( .C1(n11718), .C2(n11717), .A(n12007), .B(n15390), .ZN(
        n11723) );
  NAND2_X1 U14140 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n15490) );
  INV_X1 U14141 ( .A(n15490), .ZN(n11720) );
  INV_X1 U14142 ( .A(n13325), .ZN(n12219) );
  OAI22_X1 U14143 ( .A1(n11780), .A2(n13295), .B1(n13315), .B2(n12219), .ZN(
        n11719) );
  AOI211_X1 U14144 ( .C1(n11721), .C2(n15377), .A(n11720), .B(n11719), .ZN(
        n11722) );
  OAI211_X1 U14145 ( .C1(n11781), .C2(n15401), .A(n11723), .B(n11722), .ZN(
        P3_U3161) );
  INV_X1 U14146 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n14452) );
  NOR2_X1 U14147 ( .A1(n11725), .A2(n11724), .ZN(n14453) );
  MUX2_X1 U14148 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n14452), .S(n14451), .Z(
        n11726) );
  OAI21_X1 U14149 ( .B1(n14458), .B2(n14453), .A(n11726), .ZN(n14456) );
  OAI21_X1 U14150 ( .B1(n14452), .B2(n11727), .A(n14456), .ZN(n11728) );
  NOR2_X1 U14151 ( .A1(n11728), .A2(n12444), .ZN(n11730) );
  XNOR2_X1 U14152 ( .A(n11728), .B(n12444), .ZN(n15106) );
  NOR2_X1 U14153 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n15106), .ZN(n15105) );
  INV_X1 U14154 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n12020) );
  MUX2_X1 U14155 ( .A(n12020), .B(P1_REG2_REG_16__SCAN_IN), .S(n12628), .Z(
        n11729) );
  OAI21_X1 U14156 ( .B1(n11730), .B2(n15105), .A(n11729), .ZN(n11731) );
  NAND3_X1 U14157 ( .A1(n11731), .A2(n14482), .A3(n12019), .ZN(n11739) );
  NAND2_X1 U14158 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n14259)
         );
  XOR2_X1 U14159 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n12628), .Z(n11735) );
  INV_X1 U14160 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n15078) );
  MUX2_X1 U14161 ( .A(P1_REG1_REG_14__SCAN_IN), .B(n15078), .S(n14451), .Z(
        n14447) );
  NAND2_X1 U14162 ( .A1(n14446), .A2(n14447), .ZN(n14445) );
  OAI21_X1 U14163 ( .B1(n14451), .B2(P1_REG1_REG_14__SCAN_IN), .A(n14445), 
        .ZN(n11733) );
  XNOR2_X1 U14164 ( .A(n11733), .B(n15111), .ZN(n15108) );
  NOR2_X1 U14165 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n15108), .ZN(n15107) );
  OAI211_X1 U14166 ( .C1(n11735), .C2(n11734), .A(n14477), .B(n12021), .ZN(
        n11736) );
  NAND2_X1 U14167 ( .A1(n14259), .A2(n11736), .ZN(n11737) );
  AOI21_X1 U14168 ( .B1(n14435), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n11737), 
        .ZN(n11738) );
  OAI211_X1 U14169 ( .C1(n15122), .C2(n12022), .A(n11739), .B(n11738), .ZN(
        P1_U3259) );
  XNOR2_X1 U14170 ( .A(n11740), .B(n11742), .ZN(n15543) );
  INV_X1 U14171 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n11746) );
  OAI211_X1 U14172 ( .C1(n11743), .C2(n11742), .A(n11741), .B(n13552), .ZN(
        n11745) );
  AND2_X1 U14173 ( .A1(n11745), .A2(n11744), .ZN(n15548) );
  MUX2_X1 U14174 ( .A(n11746), .B(n15548), .S(n13541), .Z(n11749) );
  AOI22_X1 U14175 ( .A1(n13543), .A2(n15545), .B1(n13559), .B2(n11747), .ZN(
        n11748) );
  OAI211_X1 U14176 ( .C1(n13125), .C2(n15543), .A(n11749), .B(n11748), .ZN(
        P3_U3229) );
  XNOR2_X1 U14177 ( .A(n11750), .B(n11753), .ZN(n15541) );
  INV_X1 U14178 ( .A(n15541), .ZN(n11762) );
  NAND2_X1 U14179 ( .A1(n11752), .A2(n11751), .ZN(n11754) );
  AOI21_X1 U14180 ( .B1(n11754), .B2(n11753), .A(n13515), .ZN(n11757) );
  OAI22_X1 U14181 ( .A1(n8952), .A2(n13518), .B1(n11755), .B2(n13520), .ZN(
        n15384) );
  AOI21_X1 U14182 ( .B1(n11757), .B2(n11756), .A(n15384), .ZN(n15538) );
  MUX2_X1 U14183 ( .A(n7158), .B(n15538), .S(n13541), .Z(n11761) );
  AOI22_X1 U14184 ( .A1(n13543), .A2(n11759), .B1(n13559), .B2(n11758), .ZN(
        n11760) );
  OAI211_X1 U14185 ( .C1(n13125), .C2(n11762), .A(n11761), .B(n11760), .ZN(
        P3_U3230) );
  NAND2_X1 U14186 ( .A1(n11936), .A2(n11763), .ZN(n11764) );
  XOR2_X1 U14187 ( .A(n11765), .B(n11764), .Z(n15556) );
  AOI21_X1 U14188 ( .B1(n11766), .B2(n11765), .A(n13515), .ZN(n11771) );
  OR2_X1 U14189 ( .A1(n11767), .A2(n13518), .ZN(n11769) );
  OR2_X1 U14190 ( .A1(n11780), .A2(n13520), .ZN(n11768) );
  NAND2_X1 U14191 ( .A1(n11769), .A2(n11768), .ZN(n15394) );
  AOI21_X1 U14192 ( .B1(n11771), .B2(n11770), .A(n15394), .ZN(n15555) );
  INV_X1 U14193 ( .A(P3_REG2_REG_6__SCAN_IN), .ZN(n11772) );
  MUX2_X1 U14194 ( .A(n15555), .B(n11772), .S(n13560), .Z(n11775) );
  AOI22_X1 U14195 ( .A1(n13543), .A2(n15560), .B1(n13559), .B2(n11773), .ZN(
        n11774) );
  OAI211_X1 U14196 ( .C1(n13125), .C2(n15556), .A(n11775), .B(n11774), .ZN(
        P3_U3227) );
  XOR2_X1 U14197 ( .A(n11776), .B(n11778), .Z(n15571) );
  XOR2_X1 U14198 ( .A(n11778), .B(n11777), .Z(n11779) );
  OAI222_X1 U14199 ( .A1(n13520), .A2(n12219), .B1(n13518), .B2(n11780), .C1(
        n11779), .C2(n13515), .ZN(n15573) );
  NAND2_X1 U14200 ( .A1(n15573), .A2(n13541), .ZN(n11784) );
  OAI22_X1 U14201 ( .A1(n13562), .A2(n15569), .B1(n11781), .B2(n13538), .ZN(
        n11782) );
  AOI21_X1 U14202 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n13560), .A(n11782), .ZN(
        n11783) );
  OAI211_X1 U14203 ( .C1(n13125), .C2(n15571), .A(n11784), .B(n11783), .ZN(
        P3_U3225) );
  INV_X1 U14204 ( .A(n12840), .ZN(n11792) );
  AOI21_X1 U14205 ( .B1(n14618), .B2(n14708), .A(n14649), .ZN(n11791) );
  INV_X1 U14206 ( .A(n14606), .ZN(n11789) );
  OAI22_X1 U14207 ( .A1(n14708), .A2(n10249), .B1(n11785), .B2(n14706), .ZN(
        n11788) );
  AOI21_X1 U14208 ( .B1(n14635), .B2(n14709), .A(n11786), .ZN(n11787) );
  AOI211_X1 U14209 ( .C1(n11789), .C2(n14378), .A(n11788), .B(n11787), .ZN(
        n11790) );
  OAI21_X1 U14210 ( .B1(n11792), .B2(n11791), .A(n11790), .ZN(P1_U3293) );
  INV_X1 U14211 ( .A(n11793), .ZN(n11794) );
  AOI211_X1 U14212 ( .C1(n11796), .C2(n12475), .A(n11795), .B(n11794), .ZN(
        n11804) );
  NOR2_X1 U14213 ( .A1(n14709), .A2(n11797), .ZN(n11801) );
  OAI22_X1 U14214 ( .A1(n14708), .A2(n11799), .B1(n11798), .B2(n14706), .ZN(
        n11800) );
  AOI211_X1 U14215 ( .C1(n11802), .C2(n14649), .A(n11801), .B(n11800), .ZN(
        n11803) );
  OAI21_X1 U14216 ( .B1(n11804), .B2(n15143), .A(n11803), .ZN(P1_U3289) );
  OAI21_X1 U14217 ( .B1(P2_REG2_REG_15__SCAN_IN), .B2(n11806), .A(n11805), 
        .ZN(n11815) );
  AND2_X1 U14218 ( .A1(P2_U3088), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n12361) );
  AOI21_X1 U14219 ( .B1(n15250), .B2(P2_ADDR_REG_15__SCAN_IN), .A(n12361), 
        .ZN(n11811) );
  OAI21_X1 U14220 ( .B1(n11808), .B2(P2_REG1_REG_15__SCAN_IN), .A(n11807), 
        .ZN(n11809) );
  OR2_X1 U14221 ( .A1(n13901), .A2(n11809), .ZN(n11810) );
  OAI211_X1 U14222 ( .C1(n15225), .C2(n11812), .A(n11811), .B(n11810), .ZN(
        n11813) );
  INV_X1 U14223 ( .A(n11813), .ZN(n11814) );
  OAI21_X1 U14224 ( .B1(n11815), .B2(n12354), .A(n11814), .ZN(P2_U3229) );
  INV_X1 U14225 ( .A(n14196), .ZN(n14197) );
  NAND2_X1 U14226 ( .A1(n12524), .A2(n14197), .ZN(n11817) );
  OAI211_X1 U14227 ( .C1(n11818), .C2(n14201), .A(n11817), .B(n11816), .ZN(
        P2_U3304) );
  INV_X1 U14228 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n12525) );
  NAND2_X1 U14229 ( .A1(n12524), .A2(n11819), .ZN(n11820) );
  OAI211_X1 U14230 ( .C1(n12525), .C2(n14876), .A(n11820), .B(n12883), .ZN(
        P1_U3332) );
  XNOR2_X1 U14231 ( .A(n11822), .B(n11821), .ZN(n15584) );
  OAI211_X1 U14232 ( .C1(n11825), .C2(n11824), .A(n11823), .B(n13552), .ZN(
        n11828) );
  OR2_X1 U14233 ( .A1(n12390), .A2(n13520), .ZN(n11827) );
  NAND2_X1 U14234 ( .A1(n13325), .A2(n13531), .ZN(n11826) );
  AND2_X1 U14235 ( .A1(n11827), .A2(n11826), .ZN(n15369) );
  NAND2_X1 U14236 ( .A1(n11828), .A2(n15369), .ZN(n15585) );
  NAND2_X1 U14237 ( .A1(n15585), .A2(n13541), .ZN(n11831) );
  OAI22_X1 U14238 ( .A1(n13562), .A2(n15581), .B1(n15380), .B2(n13538), .ZN(
        n11829) );
  AOI21_X1 U14239 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n13560), .A(n11829), 
        .ZN(n11830) );
  OAI211_X1 U14240 ( .C1(n15584), .C2(n13125), .A(n11831), .B(n11830), .ZN(
        P3_U3223) );
  OR2_X1 U14241 ( .A1(n12580), .A2(n14371), .ZN(n11832) );
  NAND2_X1 U14242 ( .A1(n11834), .A2(n12819), .ZN(n11837) );
  AOI22_X1 U14243 ( .A1(n12661), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n12660), 
        .B2(n11835), .ZN(n11836) );
  XNOR2_X1 U14244 ( .A(n12589), .B(n12082), .ZN(n12847) );
  OAI21_X1 U14245 ( .B1(n11838), .B2(n12847), .A(n11972), .ZN(n11998) );
  INV_X1 U14246 ( .A(n11998), .ZN(n11857) );
  OR2_X1 U14247 ( .A1(n12580), .A2(n12123), .ZN(n11839) );
  CLKBUF_X1 U14248 ( .A(n11841), .Z(n11844) );
  CLKBUF_X1 U14249 ( .A(n11977), .Z(n11842) );
  INV_X1 U14250 ( .A(n11842), .ZN(n11843) );
  AOI21_X1 U14251 ( .B1(n12847), .B2(n11844), .A(n11843), .ZN(n11852) );
  NAND2_X1 U14252 ( .A1(n12811), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n11849) );
  OR2_X1 U14253 ( .A1(n12664), .A2(n11991), .ZN(n11848) );
  XNOR2_X1 U14254 ( .A(n11982), .B(n11981), .ZN(n12274) );
  OR2_X1 U14255 ( .A1(n12786), .A2(n12274), .ZN(n11847) );
  INV_X1 U14256 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n11845) );
  OR2_X1 U14257 ( .A1(n10990), .A2(n11845), .ZN(n11846) );
  NAND4_X1 U14258 ( .A1(n11849), .A2(n11848), .A3(n11847), .A4(n11846), .ZN(
        n14369) );
  AOI22_X1 U14259 ( .A1(n14771), .A2(n14369), .B1(n14371), .B2(n14620), .ZN(
        n11851) );
  NAND2_X1 U14260 ( .A1(n11998), .A2(n14665), .ZN(n11850) );
  OAI211_X1 U14261 ( .C1(n11852), .C2(n14699), .A(n11851), .B(n11850), .ZN(
        n11996) );
  NAND2_X1 U14262 ( .A1(n11996), .A2(n14708), .ZN(n11856) );
  INV_X1 U14263 ( .A(n12589), .ZN(n11999) );
  AOI211_X1 U14264 ( .C1(n12589), .C2(n6692), .A(n14781), .B(n6788), .ZN(
        n11997) );
  NOR2_X1 U14265 ( .A1(n14709), .A2(n11999), .ZN(n11854) );
  OAI22_X1 U14266 ( .A1(n14708), .A2(n10432), .B1(n12122), .B2(n14706), .ZN(
        n11853) );
  AOI211_X1 U14267 ( .C1(n11997), .C2(n14713), .A(n11854), .B(n11853), .ZN(
        n11855) );
  OAI211_X1 U14268 ( .C1(n11857), .C2(n14673), .A(n11856), .B(n11855), .ZN(
        P1_U3284) );
  AOI22_X1 U14269 ( .A1(n14373), .A2(n13087), .B1(n13085), .B2(n15158), .ZN(
        n11866) );
  AOI22_X1 U14270 ( .A1(n14373), .A2(n13085), .B1(n13086), .B2(n15158), .ZN(
        n11859) );
  XNOR2_X1 U14271 ( .A(n11859), .B(n10886), .ZN(n11865) );
  INV_X1 U14272 ( .A(n11860), .ZN(n11862) );
  XOR2_X1 U14273 ( .A(n11866), .B(n11865), .Z(n14319) );
  NAND2_X1 U14274 ( .A1(n14320), .A2(n14319), .ZN(n14318) );
  NAND2_X1 U14275 ( .A1(n12577), .A2(n13086), .ZN(n11868) );
  NAND2_X1 U14276 ( .A1(n14372), .A2(n13070), .ZN(n11867) );
  NAND2_X1 U14277 ( .A1(n11868), .A2(n11867), .ZN(n11869) );
  XNOR2_X1 U14278 ( .A(n11869), .B(n10886), .ZN(n12071) );
  AOI22_X1 U14279 ( .A1(n12577), .A2(n13038), .B1(n14372), .B2(n13087), .ZN(
        n12072) );
  XNOR2_X1 U14280 ( .A(n12071), .B(n12072), .ZN(n11870) );
  OAI211_X1 U14281 ( .C1(n11871), .C2(n11870), .A(n12075), .B(n14341), .ZN(
        n11878) );
  OAI21_X1 U14282 ( .B1(n15056), .B2(n11873), .A(n11872), .ZN(n11876) );
  OAI22_X1 U14283 ( .A1(n15055), .A2(n12123), .B1(n15072), .B2(n11874), .ZN(
        n11875) );
  AOI211_X1 U14284 ( .C1(n12577), .C2(n15067), .A(n11876), .B(n11875), .ZN(
        n11877) );
  NAND2_X1 U14285 ( .A1(n11878), .A2(n11877), .ZN(P1_U3213) );
  XNOR2_X1 U14286 ( .A(n11879), .B(n11884), .ZN(n11882) );
  OR2_X1 U14287 ( .A1(n12144), .A2(n13841), .ZN(n11881) );
  OR2_X1 U14288 ( .A1(n13839), .A2(n11914), .ZN(n11880) );
  AND2_X1 U14289 ( .A1(n11881), .A2(n11880), .ZN(n11965) );
  OAI21_X1 U14290 ( .B1(n11882), .B2(n13962), .A(n11965), .ZN(n15022) );
  INV_X1 U14291 ( .A(n15022), .ZN(n11893) );
  XNOR2_X1 U14292 ( .A(n11883), .B(n11884), .ZN(n15024) );
  INV_X1 U14293 ( .A(n11885), .ZN(n11887) );
  INV_X1 U14294 ( .A(n14996), .ZN(n11886) );
  OAI211_X1 U14295 ( .C1(n15021), .C2(n11887), .A(n11886), .B(n15274), .ZN(
        n15020) );
  AOI22_X1 U14296 ( .A1(n15269), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n11968), 
        .B2(n15268), .ZN(n11890) );
  NAND2_X1 U14297 ( .A1(n11888), .A2(n15270), .ZN(n11889) );
  OAI211_X1 U14298 ( .C1(n15020), .C2(n14026), .A(n11890), .B(n11889), .ZN(
        n11891) );
  AOI21_X1 U14299 ( .B1(n15024), .B2(n15280), .A(n11891), .ZN(n11892) );
  OAI21_X1 U14300 ( .B1(n11893), .B2(n14078), .A(n11892), .ZN(P2_U3252) );
  AOI21_X1 U14301 ( .B1(n12056), .B2(n11895), .A(n11894), .ZN(n11908) );
  AOI21_X1 U14302 ( .B1(n11898), .B2(n11897), .A(n11896), .ZN(n11900) );
  NAND2_X1 U14303 ( .A1(n15523), .A2(P3_ADDR_REG_11__SCAN_IN), .ZN(n11899) );
  NAND2_X1 U14304 ( .A1(P3_U3151), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n12232)
         );
  OAI211_X1 U14305 ( .C1(n11900), .C2(n7858), .A(n11899), .B(n12232), .ZN(
        n11905) );
  AOI21_X1 U14306 ( .B1(n14958), .B2(n11902), .A(n11901), .ZN(n11903) );
  NOR2_X1 U14307 ( .A1(n11903), .A2(n15516), .ZN(n11904) );
  AOI211_X1 U14308 ( .C1(n15485), .C2(n11906), .A(n11905), .B(n11904), .ZN(
        n11907) );
  OAI21_X1 U14309 ( .B1(n11908), .B2(n15530), .A(n11907), .ZN(P3_U3193) );
  AOI21_X1 U14310 ( .B1(n15313), .B2(n11910), .A(n11909), .ZN(n11911) );
  OAI21_X1 U14311 ( .B1(n15000), .B2(n11912), .A(n11911), .ZN(n11933) );
  NAND2_X1 U14312 ( .A1(n11933), .A2(n15347), .ZN(n11913) );
  OAI21_X1 U14313 ( .B1(n15347), .B2(n9297), .A(n11913), .ZN(P2_U3463) );
  XNOR2_X1 U14314 ( .A(n15026), .B(n13734), .ZN(n11915) );
  OR2_X1 U14315 ( .A1(n10697), .A2(n11914), .ZN(n11916) );
  NAND2_X1 U14316 ( .A1(n11915), .A2(n11916), .ZN(n11961) );
  INV_X1 U14317 ( .A(n11915), .ZN(n11918) );
  INV_X1 U14318 ( .A(n11916), .ZN(n11917) );
  NAND2_X1 U14319 ( .A1(n11918), .A2(n11917), .ZN(n11963) );
  NAND2_X1 U14320 ( .A1(n11961), .A2(n11963), .ZN(n11924) );
  INV_X1 U14321 ( .A(n11919), .ZN(n11921) );
  NAND2_X1 U14322 ( .A1(n11921), .A2(n11920), .ZN(n11922) );
  XOR2_X1 U14323 ( .A(n11924), .B(n11962), .Z(n11932) );
  NAND2_X1 U14324 ( .A1(n13843), .A2(n11925), .ZN(n11926) );
  OAI211_X1 U14325 ( .C1(n13845), .C2(n11928), .A(n11927), .B(n11926), .ZN(
        n11929) );
  AOI21_X1 U14326 ( .B1(n11930), .B2(n13857), .A(n11929), .ZN(n11931) );
  OAI21_X1 U14327 ( .B1(n11932), .B2(n13859), .A(n11931), .ZN(P2_U3196) );
  NAND2_X1 U14328 ( .A1(n11933), .A2(n15357), .ZN(n11934) );
  OAI21_X1 U14329 ( .B1(n15357), .B2(n9301), .A(n11934), .ZN(P2_U3510) );
  AND2_X1 U14330 ( .A1(n8484), .A2(n11937), .ZN(n11938) );
  XNOR2_X1 U14331 ( .A(n11938), .B(n11940), .ZN(n15564) );
  OAI211_X1 U14332 ( .C1(n11941), .C2(n11940), .A(n11939), .B(n13552), .ZN(
        n11946) );
  OR2_X1 U14333 ( .A1(n11942), .A2(n13518), .ZN(n11944) );
  OR2_X1 U14334 ( .A1(n12013), .A2(n13520), .ZN(n11943) );
  NAND2_X1 U14335 ( .A1(n11944), .A2(n11943), .ZN(n15362) );
  INV_X1 U14336 ( .A(n15362), .ZN(n11945) );
  NAND2_X1 U14337 ( .A1(n11946), .A2(n11945), .ZN(n15565) );
  NAND2_X1 U14338 ( .A1(n15565), .A2(n13541), .ZN(n11949) );
  OAI22_X1 U14339 ( .A1(n13562), .A2(n15563), .B1(n15367), .B2(n13538), .ZN(
        n11947) );
  AOI21_X1 U14340 ( .B1(n13560), .B2(P3_REG2_REG_7__SCAN_IN), .A(n11947), .ZN(
        n11948) );
  OAI211_X1 U14341 ( .C1(n13125), .C2(n15564), .A(n11949), .B(n11948), .ZN(
        P3_U3226) );
  OAI21_X1 U14342 ( .B1(n11952), .B2(n11951), .A(n11950), .ZN(n11960) );
  INV_X1 U14343 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n15104) );
  NAND2_X1 U14344 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n13798)
         );
  OAI211_X1 U14345 ( .C1(n11955), .C2(n11954), .A(n11953), .B(n15255), .ZN(
        n11956) );
  OAI211_X1 U14346 ( .C1(n15104), .C2(n15228), .A(n13798), .B(n11956), .ZN(
        n11957) );
  AOI21_X1 U14347 ( .B1(n15259), .B2(n11958), .A(n11957), .ZN(n11959) );
  OAI21_X1 U14348 ( .B1(n11960), .B2(n12354), .A(n11959), .ZN(P2_U3230) );
  XNOR2_X1 U14349 ( .A(n15021), .B(n13734), .ZN(n12152) );
  AND2_X1 U14350 ( .A1(n13878), .A2(n13735), .ZN(n12153) );
  XNOR2_X1 U14351 ( .A(n12152), .B(n12153), .ZN(n12150) );
  XNOR2_X1 U14352 ( .A(n12151), .B(n12150), .ZN(n11970) );
  OAI22_X1 U14353 ( .A1(n13855), .A2(n11965), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11964), .ZN(n11967) );
  NOR2_X1 U14354 ( .A1(n15021), .A2(n13812), .ZN(n11966) );
  AOI211_X1 U14355 ( .C1(n13853), .C2(n11968), .A(n11967), .B(n11966), .ZN(
        n11969) );
  OAI21_X1 U14356 ( .B1(n11970), .B2(n13859), .A(n11969), .ZN(P2_U3206) );
  OR2_X1 U14357 ( .A1(n12589), .A2(n14370), .ZN(n11971) );
  NAND2_X1 U14358 ( .A1(n11973), .A2(n12819), .ZN(n11975) );
  AOI22_X1 U14359 ( .A1(n12661), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n12660), 
        .B2(n14418), .ZN(n11974) );
  XNOR2_X1 U14360 ( .A(n12592), .B(n15057), .ZN(n12087) );
  XNOR2_X1 U14361 ( .A(n12088), .B(n12087), .ZN(n15176) );
  INV_X1 U14362 ( .A(n15176), .ZN(n11995) );
  NAND2_X1 U14363 ( .A1(n12589), .A2(n12082), .ZN(n11976) );
  AND2_X2 U14364 ( .A1(n11977), .A2(n11976), .ZN(n11978) );
  OAI211_X1 U14365 ( .C1(n11978), .C2(n7610), .A(n12101), .B(n14618), .ZN(
        n11979) );
  OAI21_X1 U14366 ( .B1(n12082), .B2(n14700), .A(n11979), .ZN(n15173) );
  OAI211_X1 U14367 ( .C1(n6788), .C2(n7042), .A(n14811), .B(n12105), .ZN(
        n15171) );
  NAND2_X1 U14368 ( .A1(n12812), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n11989) );
  INV_X1 U14369 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n11980) );
  OAI21_X1 U14370 ( .B1(n11982), .B2(n11981), .A(n11980), .ZN(n11983) );
  NAND2_X1 U14371 ( .A1(n11983), .A2(n12094), .ZN(n15071) );
  OR2_X1 U14372 ( .A1(n12786), .A2(n15071), .ZN(n11988) );
  INV_X1 U14373 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n11984) );
  OR2_X1 U14374 ( .A1(n10990), .A2(n11984), .ZN(n11987) );
  OR2_X1 U14375 ( .A1(n12670), .A2(n11985), .ZN(n11986) );
  NAND4_X1 U14376 ( .A1(n11989), .A2(n11988), .A3(n11987), .A4(n11986), .ZN(
        n14368) );
  NAND2_X1 U14377 ( .A1(n14368), .A2(n14771), .ZN(n15170) );
  AOI21_X1 U14378 ( .B1(n15171), .B2(n15170), .A(n14483), .ZN(n11990) );
  OAI21_X1 U14379 ( .B1(n15173), .B2(n11990), .A(n14708), .ZN(n11994) );
  OAI22_X1 U14380 ( .A1(n14708), .A2(n11991), .B1(n12274), .B2(n14706), .ZN(
        n11992) );
  AOI21_X1 U14381 ( .B1(n15140), .B2(n12592), .A(n11992), .ZN(n11993) );
  OAI211_X1 U14382 ( .C1(n11995), .C2(n14716), .A(n11994), .B(n11993), .ZN(
        P1_U3283) );
  AOI211_X1 U14383 ( .C1(n14910), .C2(n11998), .A(n11997), .B(n11996), .ZN(
        n12003) );
  OAI22_X1 U14384 ( .A1(n11999), .A2(n14858), .B1(n14854), .B2(n11692), .ZN(
        n12000) );
  INV_X1 U14385 ( .A(n12000), .ZN(n12001) );
  OAI21_X1 U14386 ( .B1(n12003), .B2(n15177), .A(n12001), .ZN(P1_U3486) );
  INV_X1 U14387 ( .A(n14804), .ZN(n12200) );
  AOI22_X1 U14388 ( .A1(n12200), .A2(n12589), .B1(n15181), .B2(
        P1_REG1_REG_9__SCAN_IN), .ZN(n12002) );
  OAI21_X1 U14389 ( .B1(n12003), .B2(n15181), .A(n12002), .ZN(P1_U3537) );
  XNOR2_X1 U14390 ( .A(n12432), .B(n15575), .ZN(n12218) );
  XNOR2_X1 U14391 ( .A(n12218), .B(n13325), .ZN(n12011) );
  NAND2_X1 U14392 ( .A1(n12005), .A2(n12004), .ZN(n12006) );
  INV_X1 U14393 ( .A(n12222), .ZN(n12009) );
  AOI21_X1 U14394 ( .B1(n12011), .B2(n12010), .A(n12009), .ZN(n12018) );
  OAI22_X1 U14395 ( .A1(n15397), .A2(n15575), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12012), .ZN(n12015) );
  OAI22_X1 U14396 ( .A1(n12013), .A2(n13295), .B1(n13315), .B2(n12223), .ZN(
        n12014) );
  AOI211_X1 U14397 ( .C1(n13319), .C2(n12016), .A(n12015), .B(n12014), .ZN(
        n12017) );
  OAI21_X1 U14398 ( .B1(n12018), .B2(n15381), .A(n12017), .ZN(P3_U3171) );
  MUX2_X1 U14399 ( .A(n14685), .B(P1_REG2_REG_17__SCAN_IN), .S(n14467), .Z(
        n14468) );
  OAI21_X1 U14400 ( .B1(n12020), .B2(n12022), .A(n12019), .ZN(n14470) );
  XOR2_X1 U14401 ( .A(n14468), .B(n14470), .Z(n12030) );
  NAND2_X1 U14402 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n14268)
         );
  INV_X1 U14403 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n14802) );
  XNOR2_X1 U14404 ( .A(n14467), .B(n14802), .ZN(n12025) );
  INV_X1 U14405 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n12023) );
  OAI21_X1 U14406 ( .B1(n12023), .B2(n12022), .A(n12021), .ZN(n12024) );
  NAND2_X1 U14407 ( .A1(n12024), .A2(n12025), .ZN(n14462) );
  OAI211_X1 U14408 ( .C1(n12025), .C2(n12024), .A(n14477), .B(n14462), .ZN(
        n12026) );
  NAND2_X1 U14409 ( .A1(n14268), .A2(n12026), .ZN(n12028) );
  NOR2_X1 U14410 ( .A1(n15122), .A2(n14463), .ZN(n12027) );
  AOI211_X1 U14411 ( .C1(n14435), .C2(P1_ADDR_REG_17__SCAN_IN), .A(n12028), 
        .B(n12027), .ZN(n12029) );
  OAI21_X1 U14412 ( .B1(n12030), .B2(n15121), .A(n12029), .ZN(P1_U3260) );
  INV_X1 U14413 ( .A(n12031), .ZN(n12034) );
  OAI222_X1 U14414 ( .A1(n13688), .A2(n12034), .B1(n12033), .B2(P3_U3151), 
        .C1(n12032), .C2(n13690), .ZN(P3_U3270) );
  XNOR2_X1 U14415 ( .A(n12035), .B(n6740), .ZN(n12038) );
  NAND2_X1 U14416 ( .A1(n13186), .A2(n13533), .ZN(n12036) );
  OAI21_X1 U14417 ( .B1(n12390), .B2(n13518), .A(n12036), .ZN(n12037) );
  AOI21_X1 U14418 ( .B1(n12038), .B2(n13552), .A(n12037), .ZN(n14951) );
  INV_X1 U14419 ( .A(n14948), .ZN(n12040) );
  INV_X1 U14420 ( .A(n12039), .ZN(n12403) );
  OAI22_X1 U14421 ( .A1(n13562), .A2(n12040), .B1(n12403), .B2(n13538), .ZN(
        n12041) );
  AOI21_X1 U14422 ( .B1(P3_REG2_REG_12__SCAN_IN), .B2(n13560), .A(n12041), 
        .ZN(n12044) );
  XNOR2_X1 U14423 ( .A(n12042), .B(n6740), .ZN(n14949) );
  NAND2_X1 U14424 ( .A1(n14949), .A2(n13564), .ZN(n12043) );
  OAI211_X1 U14425 ( .C1(n14951), .C2(n13560), .A(n12044), .B(n12043), .ZN(
        P3_U3221) );
  XNOR2_X1 U14426 ( .A(n12046), .B(n12045), .ZN(n12050) );
  OR2_X1 U14427 ( .A1(n12223), .A2(n13518), .ZN(n12048) );
  OR2_X1 U14428 ( .A1(n12388), .A2(n13520), .ZN(n12047) );
  NAND2_X1 U14429 ( .A1(n12048), .A2(n12047), .ZN(n12230) );
  INV_X1 U14430 ( .A(n12230), .ZN(n12049) );
  OAI21_X1 U14431 ( .B1(n12050), .B2(n13515), .A(n12049), .ZN(n14954) );
  INV_X1 U14432 ( .A(n14954), .ZN(n12059) );
  OAI21_X1 U14433 ( .B1(n12053), .B2(n12052), .A(n12051), .ZN(n14956) );
  AOI22_X1 U14434 ( .A1(n13543), .A2(n12054), .B1(n13559), .B2(n12234), .ZN(
        n12055) );
  OAI21_X1 U14435 ( .B1(n12056), .B2(n13541), .A(n12055), .ZN(n12057) );
  AOI21_X1 U14436 ( .B1(n14956), .B2(n13564), .A(n12057), .ZN(n12058) );
  OAI21_X1 U14437 ( .B1(n12059), .B2(n13566), .A(n12058), .ZN(P3_U3222) );
  XNOR2_X1 U14438 ( .A(n12060), .B(n12063), .ZN(n12061) );
  AOI22_X1 U14439 ( .A1(n13875), .A2(n13852), .B1(n13877), .B2(n13851), .ZN(
        n12359) );
  OAI21_X1 U14440 ( .B1(n12061), .B2(n13962), .A(n12359), .ZN(n15009) );
  INV_X1 U14441 ( .A(n15009), .ZN(n12069) );
  OAI21_X1 U14442 ( .B1(n7641), .B2(n12063), .A(n12062), .ZN(n15011) );
  OAI211_X1 U14443 ( .C1(n15008), .C2(n14994), .A(n15274), .B(n14980), .ZN(
        n15007) );
  INV_X1 U14444 ( .A(n12064), .ZN(n12362) );
  AOI22_X1 U14445 ( .A1(n15269), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n12362), 
        .B2(n15268), .ZN(n12066) );
  NAND2_X1 U14446 ( .A1(n12363), .A2(n15270), .ZN(n12065) );
  OAI211_X1 U14447 ( .C1(n15007), .C2(n14026), .A(n12066), .B(n12065), .ZN(
        n12067) );
  AOI21_X1 U14448 ( .B1(n15011), .B2(n15280), .A(n12067), .ZN(n12068) );
  OAI21_X1 U14449 ( .B1(n12069), .B2(n14078), .A(n12068), .ZN(P2_U3250) );
  AOI22_X1 U14450 ( .A1(n12580), .A2(n13086), .B1(n13085), .B2(n14371), .ZN(
        n12070) );
  XNOR2_X1 U14451 ( .A(n12070), .B(n10886), .ZN(n12111) );
  AOI22_X1 U14452 ( .A1(n12580), .A2(n13038), .B1(n13087), .B2(n14371), .ZN(
        n12112) );
  XNOR2_X1 U14453 ( .A(n12111), .B(n12112), .ZN(n12078) );
  INV_X1 U14454 ( .A(n12072), .ZN(n12073) );
  INV_X1 U14455 ( .A(n12114), .ZN(n12076) );
  AOI21_X1 U14456 ( .B1(n12078), .B2(n12077), .A(n12076), .ZN(n12086) );
  INV_X1 U14457 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n12079) );
  OAI22_X1 U14458 ( .A1(n15056), .A2(n12080), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12079), .ZN(n12084) );
  OAI22_X1 U14459 ( .A1(n15055), .A2(n12082), .B1(n15072), .B2(n12081), .ZN(
        n12083) );
  AOI211_X1 U14460 ( .C1(n12580), .C2(n15067), .A(n12084), .B(n12083), .ZN(
        n12085) );
  OAI21_X1 U14461 ( .B1(n12086), .B2(n15062), .A(n12085), .ZN(P1_U3221) );
  NAND2_X1 U14462 ( .A1(n12089), .A2(n12819), .ZN(n12092) );
  AOI22_X1 U14463 ( .A1(n12661), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n12660), 
        .B2(n12090), .ZN(n12091) );
  XNOR2_X1 U14464 ( .A(n15068), .B(n12424), .ZN(n12102) );
  OAI21_X1 U14465 ( .B1(n12093), .B2(n12102), .A(n12166), .ZN(n12196) );
  INV_X1 U14466 ( .A(n12196), .ZN(n12110) );
  NAND2_X1 U14467 ( .A1(n12702), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n12099) );
  OR2_X1 U14468 ( .A1(n12670), .A2(n14912), .ZN(n12098) );
  OR2_X1 U14469 ( .A1(n12664), .A2(n10810), .ZN(n12097) );
  INV_X1 U14470 ( .A(n12175), .ZN(n12177) );
  NAND2_X1 U14471 ( .A1(n12094), .A2(n14433), .ZN(n12095) );
  NAND2_X1 U14472 ( .A1(n12177), .A2(n12095), .ZN(n12425) );
  OR2_X1 U14473 ( .A1(n12786), .A2(n12425), .ZN(n12096) );
  NAND4_X1 U14474 ( .A1(n12099), .A2(n12098), .A3(n12097), .A4(n12096), .ZN(
        n14367) );
  OR2_X1 U14475 ( .A1(n12592), .A2(n15057), .ZN(n12100) );
  CLKBUF_X1 U14476 ( .A(n12171), .Z(n12103) );
  INV_X1 U14477 ( .A(n12102), .ZN(n12849) );
  XNOR2_X1 U14478 ( .A(n12103), .B(n12849), .ZN(n12104) );
  OAI222_X1 U14479 ( .A1(n14702), .A2(n15054), .B1(n14700), .B2(n15057), .C1(
        n12104), .C2(n14699), .ZN(n12194) );
  NAND2_X1 U14480 ( .A1(n12194), .A2(n14708), .ZN(n12109) );
  INV_X1 U14481 ( .A(n12187), .ZN(n12188) );
  AOI211_X1 U14482 ( .C1(n15068), .C2(n12105), .A(n14781), .B(n12188), .ZN(
        n12195) );
  NOR2_X1 U14483 ( .A1(n7041), .A2(n14709), .ZN(n12107) );
  OAI22_X1 U14484 ( .A1(n14708), .A2(n10434), .B1(n15071), .B2(n14706), .ZN(
        n12106) );
  AOI211_X1 U14485 ( .C1(n12195), .C2(n14713), .A(n12107), .B(n12106), .ZN(
        n12108) );
  OAI211_X1 U14486 ( .C1(n12110), .C2(n14716), .A(n12109), .B(n12108), .ZN(
        P1_U3282) );
  NAND2_X1 U14487 ( .A1(n12111), .A2(n12112), .ZN(n12113) );
  NAND2_X1 U14488 ( .A1(n12589), .A2(n13086), .ZN(n12116) );
  NAND2_X1 U14489 ( .A1(n14370), .A2(n13085), .ZN(n12115) );
  NAND2_X1 U14490 ( .A1(n12116), .A2(n12115), .ZN(n12117) );
  XNOR2_X1 U14491 ( .A(n12117), .B(n10886), .ZN(n12265) );
  NAND2_X1 U14492 ( .A1(n12589), .A2(n13085), .ZN(n12119) );
  NAND2_X1 U14493 ( .A1(n14370), .A2(n13087), .ZN(n12118) );
  NAND2_X1 U14494 ( .A1(n12119), .A2(n12118), .ZN(n12264) );
  XNOR2_X1 U14495 ( .A(n12265), .B(n12264), .ZN(n12120) );
  XNOR2_X1 U14496 ( .A(n12269), .B(n12120), .ZN(n12127) );
  OAI22_X1 U14497 ( .A1(n15055), .A2(n15057), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n12121), .ZN(n12125) );
  OAI22_X1 U14498 ( .A1(n15056), .A2(n12123), .B1(n12122), .B2(n15072), .ZN(
        n12124) );
  AOI211_X1 U14499 ( .C1(n12589), .C2(n15067), .A(n12125), .B(n12124), .ZN(
        n12126) );
  OAI21_X1 U14500 ( .B1(n12127), .B2(n15062), .A(n12126), .ZN(P1_U3231) );
  XNOR2_X1 U14501 ( .A(n12128), .B(n12129), .ZN(n14944) );
  XNOR2_X1 U14502 ( .A(n12130), .B(n12129), .ZN(n12131) );
  OAI222_X1 U14503 ( .A1(n13520), .A2(n13137), .B1(n13518), .B2(n12388), .C1(
        n12131), .C2(n13515), .ZN(n14946) );
  NAND2_X1 U14504 ( .A1(n14946), .A2(n13541), .ZN(n12136) );
  INV_X1 U14505 ( .A(n14943), .ZN(n12134) );
  INV_X1 U14506 ( .A(n12438), .ZN(n12132) );
  OAI22_X1 U14507 ( .A1(n13541), .A2(n13333), .B1(n12132), .B2(n13538), .ZN(
        n12133) );
  AOI21_X1 U14508 ( .B1(n12134), .B2(n13543), .A(n12133), .ZN(n12135) );
  OAI211_X1 U14509 ( .C1(n13125), .C2(n14944), .A(n12136), .B(n12135), .ZN(
        P3_U3220) );
  INV_X1 U14510 ( .A(n12137), .ZN(n12140) );
  OAI222_X1 U14511 ( .A1(n13688), .A2(n12140), .B1(n13690), .B2(n12139), .C1(
        P3_U3151), .C2(n12138), .ZN(P3_U3269) );
  INV_X1 U14512 ( .A(n12141), .ZN(n12143) );
  INV_X1 U14513 ( .A(n12746), .ZN(n12470) );
  OAI222_X1 U14514 ( .A1(n12143), .A2(P2_U3088), .B1(n14196), .B2(n12470), 
        .C1(n12142), .C2(n14201), .ZN(P2_U3303) );
  XNOR2_X1 U14515 ( .A(n15014), .B(n13734), .ZN(n12145) );
  OR2_X1 U14516 ( .A1(n12144), .A2(n10697), .ZN(n12146) );
  NAND2_X1 U14517 ( .A1(n12145), .A2(n12146), .ZN(n12356) );
  INV_X1 U14518 ( .A(n12145), .ZN(n12148) );
  INV_X1 U14519 ( .A(n12146), .ZN(n12147) );
  NAND2_X1 U14520 ( .A1(n12148), .A2(n12147), .ZN(n12149) );
  NAND2_X1 U14521 ( .A1(n12356), .A2(n12149), .ZN(n12159) );
  INV_X1 U14522 ( .A(n12152), .ZN(n12154) );
  NAND2_X1 U14523 ( .A1(n12154), .A2(n12153), .ZN(n12155) );
  INV_X1 U14524 ( .A(n12357), .ZN(n12157) );
  AOI21_X1 U14525 ( .B1(n12159), .B2(n12158), .A(n12157), .ZN(n12164) );
  AOI22_X1 U14526 ( .A1(n13876), .A2(n13852), .B1(n13851), .B2(n13878), .ZN(
        n14987) );
  OAI22_X1 U14527 ( .A1(n13855), .A2(n14987), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12160), .ZN(n12162) );
  NOR2_X1 U14528 ( .A1(n15014), .A2(n13812), .ZN(n12161) );
  AOI211_X1 U14529 ( .C1(n13853), .C2(n14990), .A(n12162), .B(n12161), .ZN(
        n12163) );
  OAI21_X1 U14530 ( .B1(n12164), .B2(n13859), .A(n12163), .ZN(P2_U3187) );
  OR2_X1 U14531 ( .A1(n15068), .A2(n14368), .ZN(n12165) );
  NAND2_X1 U14532 ( .A1(n12166), .A2(n12165), .ZN(n12170) );
  NAND2_X1 U14533 ( .A1(n12167), .A2(n12819), .ZN(n12169) );
  AOI22_X1 U14534 ( .A1(n12661), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n14440), 
        .B2(n12660), .ZN(n12168) );
  XNOR2_X1 U14535 ( .A(n12608), .B(n15054), .ZN(n12851) );
  NAND2_X1 U14536 ( .A1(n12170), .A2(n12851), .ZN(n12238) );
  OAI21_X1 U14537 ( .B1(n12170), .B2(n12851), .A(n12238), .ZN(n14909) );
  INV_X1 U14538 ( .A(n14909), .ZN(n12193) );
  NAND2_X1 U14539 ( .A1(n12171), .A2(n12849), .ZN(n12173) );
  OR2_X1 U14540 ( .A1(n15068), .A2(n12424), .ZN(n12172) );
  NAND2_X1 U14541 ( .A1(n12173), .A2(n12172), .ZN(n12253) );
  INV_X1 U14542 ( .A(n12851), .ZN(n12252) );
  XNOR2_X1 U14543 ( .A(n12174), .B(n12252), .ZN(n12186) );
  NAND2_X1 U14544 ( .A1(n12811), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n12183) );
  OR2_X1 U14545 ( .A1(n12664), .A2(n11724), .ZN(n12182) );
  NAND2_X1 U14546 ( .A1(n12175), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n12245) );
  INV_X1 U14547 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n12176) );
  NAND2_X1 U14548 ( .A1(n12177), .A2(n12176), .ZN(n12178) );
  NAND2_X1 U14549 ( .A1(n12245), .A2(n12178), .ZN(n14294) );
  OR2_X1 U14550 ( .A1(n12753), .A2(n14294), .ZN(n12181) );
  INV_X1 U14551 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n12179) );
  OR2_X1 U14552 ( .A1(n10990), .A2(n12179), .ZN(n12180) );
  NAND4_X1 U14553 ( .A1(n12183), .A2(n12182), .A3(n12181), .A4(n12180), .ZN(
        n14366) );
  OAI22_X1 U14554 ( .A1(n15041), .A2(n14702), .B1(n12424), .B2(n14700), .ZN(
        n12184) );
  AOI21_X1 U14555 ( .B1(n14909), .B2(n14665), .A(n12184), .ZN(n12185) );
  OAI21_X1 U14556 ( .B1(n14699), .B2(n12186), .A(n12185), .ZN(n14907) );
  NAND2_X1 U14557 ( .A1(n14907), .A2(n14708), .ZN(n12192) );
  OAI22_X1 U14558 ( .A1(n14708), .A2(n10810), .B1(n12425), .B2(n14706), .ZN(
        n12190) );
  INV_X1 U14559 ( .A(n12608), .ZN(n14906) );
  NOR2_X1 U14560 ( .A1(n12187), .A2(n12608), .ZN(n12257) );
  INV_X1 U14561 ( .A(n12257), .ZN(n12258) );
  OAI211_X1 U14562 ( .C1(n14906), .C2(n12188), .A(n12258), .B(n14811), .ZN(
        n14905) );
  NOR2_X1 U14563 ( .A1(n14905), .A2(n15146), .ZN(n12189) );
  AOI211_X1 U14564 ( .C1(n15140), .C2(n12608), .A(n12190), .B(n12189), .ZN(
        n12191) );
  OAI211_X1 U14565 ( .C1(n12193), .C2(n14673), .A(n12192), .B(n12191), .ZN(
        P1_U3281) );
  AOI211_X1 U14566 ( .C1(n15175), .C2(n12196), .A(n12195), .B(n12194), .ZN(
        n12202) );
  INV_X1 U14567 ( .A(n14858), .ZN(n12198) );
  NOR2_X1 U14568 ( .A1(n14854), .A2(n11984), .ZN(n12197) );
  AOI21_X1 U14569 ( .B1(n15068), .B2(n12198), .A(n12197), .ZN(n12199) );
  OAI21_X1 U14570 ( .B1(n12202), .B2(n15177), .A(n12199), .ZN(P1_U3492) );
  AOI22_X1 U14571 ( .A1(n15068), .A2(n12200), .B1(n15181), .B2(
        P1_REG1_REG_11__SCAN_IN), .ZN(n12201) );
  OAI21_X1 U14572 ( .B1(n12202), .B2(n15181), .A(n12201), .ZN(P1_U3539) );
  XNOR2_X1 U14573 ( .A(n12204), .B(n12203), .ZN(n14939) );
  XNOR2_X1 U14574 ( .A(n12206), .B(n12205), .ZN(n12207) );
  OAI222_X1 U14575 ( .A1(n13518), .A2(n12433), .B1(n13520), .B2(n13188), .C1(
        n12207), .C2(n13515), .ZN(n14941) );
  NAND2_X1 U14576 ( .A1(n14941), .A2(n13541), .ZN(n12213) );
  INV_X1 U14577 ( .A(n14938), .ZN(n12211) );
  INV_X1 U14578 ( .A(P3_REG2_REG_14__SCAN_IN), .ZN(n12209) );
  INV_X1 U14579 ( .A(n13190), .ZN(n12208) );
  OAI22_X1 U14580 ( .A1(n13541), .A2(n12209), .B1(n12208), .B2(n13538), .ZN(
        n12210) );
  AOI21_X1 U14581 ( .B1(n12211), .B2(n13543), .A(n12210), .ZN(n12212) );
  OAI211_X1 U14582 ( .C1(n14939), .C2(n13125), .A(n12213), .B(n12212), .ZN(
        P3_U3219) );
  INV_X1 U14583 ( .A(n12214), .ZN(n12216) );
  OAI222_X1 U14584 ( .A1(n12217), .A2(P3_U3151), .B1(n13688), .B2(n12216), 
        .C1(n12215), .C2(n13690), .ZN(P3_U3268) );
  INV_X1 U14585 ( .A(n12218), .ZN(n12220) );
  NAND2_X1 U14586 ( .A1(n12220), .A2(n12219), .ZN(n12221) );
  XNOR2_X1 U14587 ( .A(n12432), .B(n15378), .ZN(n12224) );
  XNOR2_X1 U14588 ( .A(n12224), .B(n12223), .ZN(n15374) );
  INV_X1 U14589 ( .A(n12224), .ZN(n12225) );
  NAND2_X1 U14590 ( .A1(n12225), .A2(n13324), .ZN(n12226) );
  XNOR2_X1 U14591 ( .A(n12432), .B(n14953), .ZN(n12227) );
  NAND2_X1 U14592 ( .A1(n12392), .A2(n12391), .ZN(n12229) );
  XNOR2_X1 U14593 ( .A(n12229), .B(n12390), .ZN(n12236) );
  NAND2_X1 U14594 ( .A1(n12230), .A2(n15393), .ZN(n12231) );
  OAI211_X1 U14595 ( .C1(n15397), .C2(n14953), .A(n12232), .B(n12231), .ZN(
        n12233) );
  AOI21_X1 U14596 ( .B1(n13319), .B2(n12234), .A(n12233), .ZN(n12235) );
  OAI21_X1 U14597 ( .B1(n12236), .B2(n15381), .A(n12235), .ZN(P3_U3176) );
  OR2_X1 U14598 ( .A1(n12608), .A2(n14367), .ZN(n12237) );
  NAND2_X1 U14599 ( .A1(n12238), .A2(n12237), .ZN(n12243) );
  NAND2_X1 U14600 ( .A1(n12239), .A2(n12819), .ZN(n12242) );
  AOI22_X1 U14601 ( .A1(n12240), .A2(n12660), .B1(n12661), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n12241) );
  XNOR2_X1 U14602 ( .A(n12957), .B(n15041), .ZN(n12852) );
  OAI21_X1 U14603 ( .B1(n12243), .B2(n12852), .A(n12296), .ZN(n12378) );
  INV_X1 U14604 ( .A(n12378), .ZN(n12263) );
  NAND2_X1 U14605 ( .A1(n12812), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n12251) );
  INV_X1 U14606 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n12244) );
  NAND2_X1 U14607 ( .A1(n12245), .A2(n12244), .ZN(n12246) );
  NAND2_X1 U14608 ( .A1(n12309), .A2(n12246), .ZN(n15053) );
  OR2_X1 U14609 ( .A1(n12753), .A2(n15053), .ZN(n12250) );
  INV_X1 U14610 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n12247) );
  OR2_X1 U14611 ( .A1(n10990), .A2(n12247), .ZN(n12249) );
  OR2_X1 U14612 ( .A1(n12670), .A2(n15078), .ZN(n12248) );
  NAND4_X1 U14613 ( .A1(n12251), .A2(n12250), .A3(n12249), .A4(n12248), .ZN(
        n14365) );
  INV_X1 U14614 ( .A(n14365), .ZN(n14295) );
  NAND2_X1 U14615 ( .A1(n12253), .A2(n12252), .ZN(n12255) );
  OR2_X1 U14616 ( .A1(n12608), .A2(n15054), .ZN(n12254) );
  INV_X1 U14617 ( .A(n12852), .ZN(n12299) );
  XNOR2_X1 U14618 ( .A(n12300), .B(n12299), .ZN(n12256) );
  OAI222_X1 U14619 ( .A1(n14700), .A2(n15054), .B1(n14702), .B2(n14295), .C1(
        n12256), .C2(n14699), .ZN(n12376) );
  NAND2_X1 U14620 ( .A1(n12376), .A2(n14708), .ZN(n12262) );
  AOI211_X1 U14621 ( .C1(n12957), .C2(n12258), .A(n14781), .B(n12318), .ZN(
        n12377) );
  NOR2_X1 U14622 ( .A1(n14300), .A2(n14709), .ZN(n12260) );
  OAI22_X1 U14623 ( .A1(n14708), .A2(n11724), .B1(n14294), .B2(n14706), .ZN(
        n12259) );
  AOI211_X1 U14624 ( .C1(n12377), .C2(n14713), .A(n12260), .B(n12259), .ZN(
        n12261) );
  OAI211_X1 U14625 ( .C1(n12263), .C2(n14716), .A(n12262), .B(n12261), .ZN(
        P1_U3280) );
  NOR2_X1 U14626 ( .A1(n12265), .A2(n12264), .ZN(n12268) );
  INV_X1 U14627 ( .A(n12264), .ZN(n12267) );
  INV_X1 U14628 ( .A(n12265), .ZN(n12266) );
  AND2_X1 U14629 ( .A1(n14369), .A2(n13059), .ZN(n12270) );
  AOI21_X1 U14630 ( .B1(n12592), .B2(n13038), .A(n12270), .ZN(n12409) );
  AOI22_X1 U14631 ( .A1(n12592), .A2(n13086), .B1(n13085), .B2(n14369), .ZN(
        n12271) );
  XNOR2_X1 U14632 ( .A(n12271), .B(n10886), .ZN(n12408) );
  XOR2_X1 U14633 ( .A(n12409), .B(n12408), .Z(n12272) );
  OAI211_X1 U14634 ( .C1(n12273), .C2(n12272), .A(n15060), .B(n14341), .ZN(
        n12277) );
  NOR2_X1 U14635 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n11981), .ZN(n14417) );
  OAI22_X1 U14636 ( .A1(n15055), .A2(n12424), .B1(n15072), .B2(n12274), .ZN(
        n12275) );
  AOI211_X1 U14637 ( .C1(n14322), .C2(n14370), .A(n14417), .B(n12275), .ZN(
        n12276) );
  OAI211_X1 U14638 ( .C1(n7042), .C2(n14352), .A(n12277), .B(n12276), .ZN(
        P1_U3217) );
  OR2_X1 U14639 ( .A1(n12278), .A2(n12281), .ZN(n12279) );
  NAND2_X1 U14640 ( .A1(n12280), .A2(n12279), .ZN(n14165) );
  XNOR2_X1 U14641 ( .A(n12282), .B(n12281), .ZN(n12283) );
  NAND2_X1 U14642 ( .A1(n12283), .A2(n14065), .ZN(n12284) );
  AOI22_X1 U14643 ( .A1(n13873), .A2(n13852), .B1(n13851), .B2(n13875), .ZN(
        n13807) );
  NAND2_X1 U14644 ( .A1(n12284), .A2(n13807), .ZN(n14169) );
  NAND2_X1 U14645 ( .A1(n14169), .A2(n14088), .ZN(n12291) );
  INV_X1 U14646 ( .A(n13809), .ZN(n12285) );
  OAI22_X1 U14647 ( .A1(n14088), .A2(n12286), .B1(n12285), .B2(n14086), .ZN(
        n12289) );
  AOI21_X1 U14648 ( .B1(n13699), .B2(n14981), .A(n14091), .ZN(n12287) );
  NAND2_X1 U14649 ( .A1(n12287), .A2(n14092), .ZN(n14166) );
  NOR2_X1 U14650 ( .A1(n14166), .A2(n14026), .ZN(n12288) );
  AOI211_X1 U14651 ( .C1(n15270), .C2(n13699), .A(n12289), .B(n12288), .ZN(
        n12290) );
  OAI211_X1 U14652 ( .C1(n14099), .C2(n14165), .A(n12291), .B(n12290), .ZN(
        P2_U3248) );
  NAND2_X1 U14653 ( .A1(n12292), .A2(n12819), .ZN(n12294) );
  AOI22_X1 U14654 ( .A1(n14451), .A2(n12660), .B1(n12661), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n12293) );
  NAND2_X1 U14655 ( .A1(n15050), .A2(n14295), .ZN(n12615) );
  OR2_X1 U14656 ( .A1(n12957), .A2(n14366), .ZN(n12295) );
  INV_X1 U14657 ( .A(n12442), .ZN(n12297) );
  AOI21_X1 U14658 ( .B1(n12854), .B2(n12298), .A(n12297), .ZN(n15077) );
  INV_X1 U14659 ( .A(n15077), .ZN(n12323) );
  AOI22_X1 U14660 ( .A1(n15050), .A2(n15140), .B1(P1_REG2_REG_14__SCAN_IN), 
        .B2(n15143), .ZN(n12322) );
  NAND2_X1 U14661 ( .A1(n12300), .A2(n12299), .ZN(n12302) );
  OR2_X1 U14662 ( .A1(n12957), .A2(n15041), .ZN(n12301) );
  NAND2_X1 U14663 ( .A1(n12302), .A2(n12301), .ZN(n12447) );
  INV_X1 U14664 ( .A(n12854), .ZN(n12303) );
  XNOR2_X1 U14665 ( .A(n12304), .B(n12303), .ZN(n12305) );
  NAND2_X1 U14666 ( .A1(n12305), .A2(n14618), .ZN(n12317) );
  NAND2_X1 U14667 ( .A1(n12811), .A2(P1_REG1_REG_15__SCAN_IN), .ZN(n12315) );
  INV_X1 U14668 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n12306) );
  OR2_X1 U14669 ( .A1(n12664), .A2(n12306), .ZN(n12314) );
  INV_X1 U14670 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n12308) );
  NAND2_X1 U14671 ( .A1(n12309), .A2(n12308), .ZN(n12310) );
  NAND2_X1 U14672 ( .A1(n12452), .A2(n12310), .ZN(n14345) );
  OR2_X1 U14673 ( .A1(n12786), .A2(n14345), .ZN(n12313) );
  INV_X1 U14674 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n12311) );
  OR2_X1 U14675 ( .A1(n10990), .A2(n12311), .ZN(n12312) );
  NAND4_X1 U14676 ( .A1(n12315), .A2(n12314), .A3(n12313), .A4(n12312), .ZN(
        n14364) );
  AOI22_X1 U14677 ( .A1(n14620), .A2(n14366), .B1(n14364), .B2(n14771), .ZN(
        n12316) );
  NAND2_X1 U14678 ( .A1(n12317), .A2(n12316), .ZN(n15076) );
  INV_X1 U14679 ( .A(n15050), .ZN(n15074) );
  OAI21_X1 U14680 ( .B1(n12318), .B2(n15074), .A(n14811), .ZN(n12319) );
  OR2_X1 U14681 ( .A1(n12462), .A2(n12319), .ZN(n15073) );
  OAI22_X1 U14682 ( .A1(n15073), .A2(n14483), .B1(n14706), .B2(n15053), .ZN(
        n12320) );
  OAI21_X1 U14683 ( .B1(n15076), .B2(n12320), .A(n14708), .ZN(n12321) );
  OAI211_X1 U14684 ( .C1(n12323), .C2(n14716), .A(n12322), .B(n12321), .ZN(
        P1_U3279) );
  INV_X1 U14685 ( .A(n12771), .ZN(n12326) );
  OAI222_X1 U14686 ( .A1(n14876), .A2(n12772), .B1(n14874), .B2(n12326), .C1(
        P1_U3086), .C2(n12324), .ZN(P1_U3330) );
  OAI222_X1 U14687 ( .A1(n14201), .A2(n12327), .B1(n14196), .B2(n12326), .C1(
        n12325), .C2(P2_U3088), .ZN(P2_U3302) );
  XNOR2_X1 U14688 ( .A(n12328), .B(n12329), .ZN(n14934) );
  XNOR2_X1 U14689 ( .A(n12330), .B(n12329), .ZN(n12331) );
  OAI222_X1 U14690 ( .A1(n13520), .A2(n13316), .B1(n13518), .B2(n13137), .C1(
        n12331), .C2(n13515), .ZN(n14936) );
  NAND2_X1 U14691 ( .A1(n14936), .A2(n13541), .ZN(n12336) );
  INV_X1 U14692 ( .A(n14933), .ZN(n12334) );
  INV_X1 U14693 ( .A(n13318), .ZN(n12332) );
  OAI22_X1 U14694 ( .A1(n13541), .A2(n13351), .B1(n12332), .B2(n13538), .ZN(
        n12333) );
  AOI21_X1 U14695 ( .B1(n12334), .B2(n13543), .A(n12333), .ZN(n12335) );
  OAI211_X1 U14696 ( .C1(n13125), .C2(n14934), .A(n12336), .B(n12335), .ZN(
        P3_U3218) );
  NAND2_X1 U14697 ( .A1(n12337), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n12339) );
  NAND2_X1 U14698 ( .A1(n12339), .A2(n12338), .ZN(n13892) );
  XNOR2_X1 U14699 ( .A(n13897), .B(n13892), .ZN(n12340) );
  NOR2_X1 U14700 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n12340), .ZN(n13894) );
  AOI21_X1 U14701 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n12340), .A(n13894), 
        .ZN(n12355) );
  NOR2_X1 U14702 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n12341), .ZN(n12342) );
  AOI21_X1 U14703 ( .B1(n15250), .B2(P2_ADDR_REG_18__SCAN_IN), .A(n12342), 
        .ZN(n12350) );
  OAI21_X1 U14704 ( .B1(n12345), .B2(n12344), .A(n12343), .ZN(n13896) );
  INV_X1 U14705 ( .A(n13896), .ZN(n12346) );
  XNOR2_X1 U14706 ( .A(n13897), .B(n12346), .ZN(n12347) );
  NAND2_X1 U14707 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n12347), .ZN(n13899) );
  OAI21_X1 U14708 ( .B1(n12347), .B2(P2_REG1_REG_18__SCAN_IN), .A(n13899), 
        .ZN(n12348) );
  OR2_X1 U14709 ( .A1(n13901), .A2(n12348), .ZN(n12349) );
  OAI211_X1 U14710 ( .C1(n15225), .C2(n12351), .A(n12350), .B(n12349), .ZN(
        n12352) );
  INV_X1 U14711 ( .A(n12352), .ZN(n12353) );
  OAI21_X1 U14712 ( .B1(n12355), .B2(n12354), .A(n12353), .ZN(P2_U3232) );
  XNOR2_X1 U14713 ( .A(n12363), .B(n13729), .ZN(n13692) );
  NOR2_X1 U14714 ( .A1(n12358), .A2(n10697), .ZN(n13693) );
  XNOR2_X1 U14715 ( .A(n13694), .B(n13693), .ZN(n12366) );
  NOR2_X1 U14716 ( .A1(n13855), .A2(n12359), .ZN(n12360) );
  AOI211_X1 U14717 ( .C1(n13853), .C2(n12362), .A(n12361), .B(n12360), .ZN(
        n12365) );
  NAND2_X1 U14718 ( .A1(n12363), .A2(n13857), .ZN(n12364) );
  OAI211_X1 U14719 ( .C1(n12366), .C2(n13859), .A(n12365), .B(n12364), .ZN(
        P2_U3213) );
  XOR2_X1 U14720 ( .A(n12367), .B(n12370), .Z(n12368) );
  AOI22_X1 U14721 ( .A1(n13531), .A2(n13140), .B1(n13532), .B2(n13533), .ZN(
        n13248) );
  OAI21_X1 U14722 ( .B1(n12368), .B2(n13515), .A(n13248), .ZN(n13619) );
  INV_X1 U14723 ( .A(n13619), .ZN(n12375) );
  OAI21_X1 U14724 ( .B1(n12371), .B2(n12370), .A(n12369), .ZN(n13620) );
  INV_X1 U14725 ( .A(n13143), .ZN(n13675) );
  AOI22_X1 U14726 ( .A1(n13566), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n13559), 
        .B2(n13250), .ZN(n12372) );
  OAI21_X1 U14727 ( .B1(n13675), .B2(n13562), .A(n12372), .ZN(n12373) );
  AOI21_X1 U14728 ( .B1(n13620), .B2(n13564), .A(n12373), .ZN(n12374) );
  OAI21_X1 U14729 ( .B1(n12375), .B2(n13566), .A(n12374), .ZN(P3_U3217) );
  AOI211_X1 U14730 ( .C1(n15175), .C2(n12378), .A(n12377), .B(n12376), .ZN(
        n12381) );
  MUX2_X1 U14731 ( .A(n12379), .B(n12381), .S(n14801), .Z(n12380) );
  OAI21_X1 U14732 ( .B1(n14300), .B2(n14804), .A(n12380), .ZN(P1_U3541) );
  MUX2_X1 U14733 ( .A(n12179), .B(n12381), .S(n14854), .Z(n12382) );
  OAI21_X1 U14734 ( .B1(n14300), .B2(n14858), .A(n12382), .ZN(P1_U3498) );
  INV_X1 U14735 ( .A(n12792), .ZN(n12386) );
  OAI222_X1 U14736 ( .A1(n12384), .A2(P2_U3088), .B1(n14196), .B2(n12386), 
        .C1(n12383), .C2(n14201), .ZN(P2_U3301) );
  INV_X1 U14737 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n12793) );
  OAI222_X1 U14738 ( .A1(n14876), .A2(n12793), .B1(n14874), .B2(n12386), .C1(
        n12385), .C2(P1_U3086), .ZN(P1_U3329) );
  XNOR2_X1 U14739 ( .A(n14948), .B(n12432), .ZN(n12389) );
  INV_X1 U14740 ( .A(n12389), .ZN(n12387) );
  NAND2_X1 U14741 ( .A1(n12387), .A2(n13323), .ZN(n12430) );
  NAND2_X1 U14742 ( .A1(n12389), .A2(n12388), .ZN(n12393) );
  AOI21_X1 U14743 ( .B1(n12430), .B2(n12393), .A(n12394), .ZN(n12396) );
  INV_X1 U14744 ( .A(n12431), .ZN(n12395) );
  OAI22_X1 U14745 ( .A1(n12396), .A2(n12395), .B1(n12430), .B2(n7145), .ZN(
        n12397) );
  NAND2_X1 U14746 ( .A1(n12397), .A2(n15390), .ZN(n12402) );
  INV_X1 U14747 ( .A(n13295), .ZN(n13313) );
  NAND2_X1 U14748 ( .A1(n13313), .A2(n12398), .ZN(n12399) );
  NAND2_X1 U14749 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(P3_U3151), .ZN(n15499)
         );
  OAI211_X1 U14750 ( .C1(n12433), .C2(n13315), .A(n12399), .B(n15499), .ZN(
        n12400) );
  AOI21_X1 U14751 ( .B1(n14948), .B2(n15377), .A(n12400), .ZN(n12401) );
  OAI211_X1 U14752 ( .C1(n12403), .C2(n15401), .A(n12402), .B(n12401), .ZN(
        P3_U3164) );
  NAND2_X1 U14753 ( .A1(n15068), .A2(n13086), .ZN(n12405) );
  NAND2_X1 U14754 ( .A1(n14368), .A2(n13070), .ZN(n12404) );
  NAND2_X1 U14755 ( .A1(n12405), .A2(n12404), .ZN(n12406) );
  XNOR2_X1 U14756 ( .A(n12406), .B(n10886), .ZN(n12415) );
  AND2_X1 U14757 ( .A1(n14368), .A2(n13059), .ZN(n12407) );
  AOI21_X1 U14758 ( .B1(n15068), .B2(n13085), .A(n12407), .ZN(n12413) );
  XNOR2_X1 U14759 ( .A(n12415), .B(n12413), .ZN(n15058) );
  INV_X1 U14760 ( .A(n12408), .ZN(n12411) );
  INV_X1 U14761 ( .A(n12409), .ZN(n12410) );
  NAND2_X1 U14762 ( .A1(n12411), .A2(n12410), .ZN(n15059) );
  INV_X1 U14763 ( .A(n12413), .ZN(n12414) );
  AND2_X1 U14764 ( .A1(n14367), .A2(n13059), .ZN(n12417) );
  AOI21_X1 U14765 ( .B1(n12608), .B2(n13085), .A(n12417), .ZN(n12953) );
  NAND2_X1 U14766 ( .A1(n12608), .A2(n13086), .ZN(n12419) );
  NAND2_X1 U14767 ( .A1(n14367), .A2(n13070), .ZN(n12418) );
  NAND2_X1 U14768 ( .A1(n12419), .A2(n12418), .ZN(n12420) );
  XNOR2_X1 U14769 ( .A(n12420), .B(n10886), .ZN(n12952) );
  XOR2_X1 U14770 ( .A(n12953), .B(n12952), .Z(n12422) );
  AOI21_X1 U14771 ( .B1(n12421), .B2(n12422), .A(n15062), .ZN(n12423) );
  NAND2_X1 U14772 ( .A1(n12423), .A2(n12955), .ZN(n12429) );
  OAI22_X1 U14773 ( .A1(n15056), .A2(n12424), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14433), .ZN(n12427) );
  OAI22_X1 U14774 ( .A1(n15055), .A2(n15041), .B1(n12425), .B2(n15072), .ZN(
        n12426) );
  AOI211_X1 U14775 ( .C1(n12608), .C2(n15067), .A(n12427), .B(n12426), .ZN(
        n12428) );
  NAND2_X1 U14776 ( .A1(n12429), .A2(n12428), .ZN(P1_U3224) );
  XNOR2_X1 U14777 ( .A(n14943), .B(n12432), .ZN(n13134) );
  XNOR2_X1 U14778 ( .A(n13134), .B(n12433), .ZN(n12434) );
  NAND2_X1 U14779 ( .A1(n12435), .A2(n12434), .ZN(n13136) );
  OAI211_X1 U14780 ( .C1(n12435), .C2(n12434), .A(n13136), .B(n15390), .ZN(
        n12440) );
  NAND2_X1 U14781 ( .A1(n13313), .A2(n13323), .ZN(n12436) );
  NAND2_X1 U14782 ( .A1(P3_REG3_REG_13__SCAN_IN), .A2(P3_U3151), .ZN(n13337)
         );
  OAI211_X1 U14783 ( .C1(n13137), .C2(n13315), .A(n12436), .B(n13337), .ZN(
        n12437) );
  AOI21_X1 U14784 ( .B1(n13319), .B2(n12438), .A(n12437), .ZN(n12439) );
  OAI211_X1 U14785 ( .C1(n15397), .C2(n14943), .A(n12440), .B(n12439), .ZN(
        P3_U3174) );
  NAND2_X1 U14786 ( .A1(n15050), .A2(n14365), .ZN(n12441) );
  NAND2_X1 U14787 ( .A1(n12442), .A2(n12441), .ZN(n12914) );
  NAND2_X1 U14788 ( .A1(n12443), .A2(n12819), .ZN(n12446) );
  AOI22_X1 U14789 ( .A1(n12661), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n12660), 
        .B2(n12444), .ZN(n12445) );
  NAND2_X1 U14790 ( .A1(n14810), .A2(n15040), .ZN(n12624) );
  XOR2_X1 U14791 ( .A(n12914), .B(n12915), .Z(n14816) );
  NAND2_X1 U14792 ( .A1(n12447), .A2(n12854), .ZN(n12448) );
  INV_X1 U14793 ( .A(n12450), .ZN(n12449) );
  AOI21_X1 U14794 ( .B1(n12449), .B2(n12916), .A(n14699), .ZN(n12461) );
  NAND2_X1 U14795 ( .A1(n12811), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n12458) );
  OR2_X1 U14796 ( .A1(n12664), .A2(n12020), .ZN(n12457) );
  INV_X1 U14797 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n12451) );
  NAND2_X1 U14798 ( .A1(n12452), .A2(n12451), .ZN(n12453) );
  NAND2_X1 U14799 ( .A1(n12632), .A2(n12453), .ZN(n14707) );
  OR2_X1 U14800 ( .A1(n12786), .A2(n14707), .ZN(n12456) );
  INV_X1 U14801 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n12454) );
  OR2_X1 U14802 ( .A1(n10990), .A2(n12454), .ZN(n12455) );
  NAND4_X1 U14803 ( .A1(n12458), .A2(n12457), .A3(n12456), .A4(n12455), .ZN(
        n14363) );
  NAND2_X1 U14804 ( .A1(n14363), .A2(n14771), .ZN(n12460) );
  NAND2_X1 U14805 ( .A1(n14365), .A2(n14620), .ZN(n12459) );
  NAND2_X1 U14806 ( .A1(n12460), .A2(n12459), .ZN(n14348) );
  AOI21_X1 U14807 ( .B1(n12461), .B2(n12894), .A(n14348), .ZN(n14814) );
  INV_X1 U14808 ( .A(n12462), .ZN(n12464) );
  INV_X1 U14809 ( .A(n14810), .ZN(n14353) );
  INV_X1 U14810 ( .A(n14703), .ZN(n12463) );
  AOI21_X1 U14811 ( .B1(n14810), .B2(n12464), .A(n12463), .ZN(n14812) );
  INV_X1 U14812 ( .A(n12465), .ZN(n14538) );
  NAND2_X1 U14813 ( .A1(n14812), .A2(n14538), .ZN(n12466) );
  OAI211_X1 U14814 ( .C1(n14706), .C2(n14345), .A(n14814), .B(n12466), .ZN(
        n12467) );
  NAND2_X1 U14815 ( .A1(n12467), .A2(n14708), .ZN(n12469) );
  AOI22_X1 U14816 ( .A1(n14810), .A2(n15140), .B1(n15143), .B2(
        P1_REG2_REG_15__SCAN_IN), .ZN(n12468) );
  OAI211_X1 U14817 ( .C1(n14816), .C2(n14716), .A(n12469), .B(n12468), .ZN(
        P1_U3278) );
  OAI222_X1 U14818 ( .A1(n14876), .A2(n12747), .B1(n14874), .B2(n12470), .C1(
        n10222), .C2(P1_U3086), .ZN(P1_U3331) );
  NAND2_X1 U14819 ( .A1(n14186), .A2(n12819), .ZN(n12473) );
  INV_X1 U14820 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n12471) );
  OR2_X1 U14821 ( .A1(n12820), .A2(n12471), .ZN(n12472) );
  NAND2_X1 U14822 ( .A1(n12475), .A2(n12474), .ZN(n12476) );
  NAND2_X1 U14823 ( .A1(n12477), .A2(n12476), .ZN(n12499) );
  CLKBUF_X3 U14824 ( .A(n12496), .Z(n12827) );
  NOR2_X1 U14825 ( .A1(n14488), .A2(n12823), .ZN(n12867) );
  INV_X1 U14826 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n14718) );
  INV_X1 U14827 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n12479) );
  OR2_X1 U14828 ( .A1(n12664), .A2(n12479), .ZN(n12481) );
  NAND2_X1 U14829 ( .A1(n12702), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n12480) );
  OAI211_X1 U14830 ( .C1(n12670), .C2(n14718), .A(n12481), .B(n12480), .ZN(
        n14491) );
  OAI21_X1 U14831 ( .B1(n12484), .B2(n12483), .A(n12482), .ZN(n12874) );
  NAND2_X1 U14832 ( .A1(n12486), .A2(n12485), .ZN(n12871) );
  NAND2_X1 U14833 ( .A1(n12874), .A2(n12871), .ZN(n12863) );
  NAND2_X1 U14834 ( .A1(n14488), .A2(n12823), .ZN(n12865) );
  NOR2_X1 U14835 ( .A1(n12865), .A2(n14491), .ZN(n12487) );
  AOI211_X1 U14836 ( .C1(n12867), .C2(n14491), .A(n12863), .B(n12487), .ZN(
        n12488) );
  INV_X1 U14837 ( .A(n12488), .ZN(n12877) );
  INV_X1 U14838 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n14722) );
  NAND2_X1 U14839 ( .A1(n12702), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n12491) );
  INV_X1 U14840 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n12489) );
  OR2_X1 U14841 ( .A1(n12664), .A2(n12489), .ZN(n12490) );
  OAI211_X1 U14842 ( .C1(n12670), .C2(n14722), .A(n12491), .B(n12490), .ZN(
        n14354) );
  OAI21_X1 U14843 ( .B1(n14491), .B2(n12492), .A(n14354), .ZN(n12493) );
  INV_X1 U14844 ( .A(n12493), .ZN(n12497) );
  NAND2_X1 U14845 ( .A1(n12885), .A2(n12819), .ZN(n12495) );
  OR2_X1 U14846 ( .A1(n12820), .A2(n12886), .ZN(n12494) );
  INV_X1 U14847 ( .A(n12496), .ZN(n12823) );
  MUX2_X1 U14848 ( .A(n12497), .B(n14497), .S(n12823), .Z(n12835) );
  INV_X1 U14849 ( .A(n12835), .ZN(n12504) );
  NAND2_X1 U14850 ( .A1(n14491), .A2(n12823), .ZN(n12498) );
  OAI21_X1 U14851 ( .B1(n12500), .B2(n12499), .A(n12498), .ZN(n12501) );
  AND2_X1 U14852 ( .A1(n12501), .A2(n14354), .ZN(n12502) );
  AOI21_X1 U14853 ( .B1(n14497), .B2(n12827), .A(n12502), .ZN(n12834) );
  INV_X1 U14854 ( .A(n12834), .ZN(n12503) );
  INV_X1 U14855 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n12665) );
  INV_X1 U14856 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n12652) );
  INV_X1 U14857 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n14305) );
  INV_X1 U14858 ( .A(n12751), .ZN(n12509) );
  AND2_X1 U14859 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(P1_REG3_REG_23__SCAN_IN), 
        .ZN(n12508) );
  NAND2_X1 U14860 ( .A1(n12509), .A2(n12508), .ZN(n12763) );
  INV_X1 U14861 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n14250) );
  INV_X1 U14862 ( .A(n12784), .ZN(n12510) );
  NAND2_X1 U14863 ( .A1(n12510), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n12798) );
  INV_X1 U14864 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n14210) );
  INV_X1 U14865 ( .A(n13105), .ZN(n12516) );
  INV_X1 U14866 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n13104) );
  NOR2_X1 U14867 ( .A1(n12786), .A2(n13104), .ZN(n12515) );
  INV_X1 U14868 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n12513) );
  NAND2_X1 U14869 ( .A1(n12811), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n12512) );
  NAND2_X1 U14870 ( .A1(n12812), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n12511) );
  OAI211_X1 U14871 ( .C1(n12513), .C2(n6668), .A(n12512), .B(n12511), .ZN(
        n12514) );
  AOI21_X1 U14872 ( .B1(n12516), .B2(n12515), .A(n12514), .ZN(n13092) );
  INV_X1 U14873 ( .A(n13092), .ZN(n14355) );
  NAND2_X1 U14874 ( .A1(n12949), .A2(n12819), .ZN(n12518) );
  INV_X1 U14875 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n12950) );
  OR2_X1 U14876 ( .A1(n12820), .A2(n12950), .ZN(n12517) );
  INV_X1 U14877 ( .A(n12496), .ZN(n12691) );
  MUX2_X1 U14878 ( .A(n14355), .B(n13101), .S(n12691), .Z(n12829) );
  INV_X1 U14879 ( .A(n12829), .ZN(n12833) );
  XNOR2_X1 U14880 ( .A(n12751), .B(P1_REG3_REG_23__SCAN_IN), .ZN(n14572) );
  NAND2_X1 U14881 ( .A1(n14572), .A2(n12810), .ZN(n12523) );
  INV_X1 U14882 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n14837) );
  NAND2_X1 U14883 ( .A1(n12811), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n12520) );
  NAND2_X1 U14884 ( .A1(n12812), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n12519) );
  OAI211_X1 U14885 ( .C1(n14837), .C2(n10990), .A(n12520), .B(n12519), .ZN(
        n12521) );
  INV_X1 U14886 ( .A(n12521), .ZN(n12522) );
  NAND2_X1 U14887 ( .A1(n12523), .A2(n12522), .ZN(n14360) );
  NAND2_X1 U14888 ( .A1(n12524), .A2(n12819), .ZN(n12527) );
  OR2_X1 U14889 ( .A1(n12820), .A2(n12525), .ZN(n12526) );
  MUX2_X1 U14890 ( .A(n14360), .B(n13039), .S(n12691), .Z(n12745) );
  INV_X1 U14891 ( .A(n12528), .ZN(n12529) );
  NOR2_X1 U14892 ( .A1(n6859), .A2(n12529), .ZN(n12538) );
  MUX2_X1 U14893 ( .A(n14378), .B(n12530), .S(n12827), .Z(n12531) );
  INV_X1 U14894 ( .A(n12531), .ZN(n12537) );
  OR3_X1 U14895 ( .A1(n14377), .A2(n12532), .A3(n12827), .ZN(n12535) );
  NAND3_X1 U14896 ( .A1(n14377), .A2(n12533), .A3(n12496), .ZN(n12534) );
  NAND2_X1 U14897 ( .A1(n12535), .A2(n12534), .ZN(n12536) );
  AOI21_X1 U14898 ( .B1(n12538), .B2(n12537), .A(n12536), .ZN(n12550) );
  INV_X1 U14899 ( .A(n12539), .ZN(n12545) );
  AND2_X1 U14900 ( .A1(n12541), .A2(n12540), .ZN(n12543) );
  NOR2_X1 U14901 ( .A1(n12543), .A2(n12542), .ZN(n12544) );
  MUX2_X1 U14902 ( .A(n12545), .B(n12544), .S(n12827), .Z(n12548) );
  NAND3_X1 U14903 ( .A1(n12548), .A2(n12547), .A3(n12546), .ZN(n12549) );
  AND2_X1 U14904 ( .A1(n14376), .A2(n12691), .ZN(n12552) );
  NOR2_X1 U14905 ( .A1(n14376), .A2(n12691), .ZN(n12551) );
  MUX2_X1 U14906 ( .A(n12555), .B(n14375), .S(n12827), .Z(n12554) );
  INV_X1 U14907 ( .A(n12554), .ZN(n12557) );
  MUX2_X1 U14908 ( .A(n14375), .B(n12555), .S(n12827), .Z(n12556) );
  NAND2_X1 U14909 ( .A1(n12558), .A2(n12557), .ZN(n12559) );
  NAND2_X1 U14910 ( .A1(n12560), .A2(n12559), .ZN(n12563) );
  MUX2_X1 U14911 ( .A(n15131), .B(n14374), .S(n12691), .Z(n12564) );
  NAND2_X1 U14912 ( .A1(n12563), .A2(n12564), .ZN(n12562) );
  MUX2_X1 U14913 ( .A(n14374), .B(n15131), .S(n12691), .Z(n12561) );
  NAND2_X1 U14914 ( .A1(n12562), .A2(n12561), .ZN(n12568) );
  INV_X1 U14915 ( .A(n12563), .ZN(n12566) );
  INV_X1 U14916 ( .A(n12564), .ZN(n12565) );
  NAND2_X1 U14917 ( .A1(n12566), .A2(n12565), .ZN(n12567) );
  NAND2_X1 U14918 ( .A1(n12568), .A2(n12567), .ZN(n12571) );
  MUX2_X1 U14919 ( .A(n15158), .B(n14373), .S(n12827), .Z(n12572) );
  NAND2_X1 U14920 ( .A1(n12571), .A2(n12572), .ZN(n12570) );
  MUX2_X1 U14921 ( .A(n14373), .B(n15158), .S(n12827), .Z(n12569) );
  NAND2_X1 U14922 ( .A1(n12570), .A2(n12569), .ZN(n12576) );
  INV_X1 U14923 ( .A(n12571), .ZN(n12574) );
  INV_X1 U14924 ( .A(n12572), .ZN(n12573) );
  NAND2_X1 U14925 ( .A1(n12574), .A2(n12573), .ZN(n12575) );
  MUX2_X1 U14926 ( .A(n14372), .B(n12577), .S(n12827), .Z(n12579) );
  MUX2_X1 U14927 ( .A(n14372), .B(n12577), .S(n12691), .Z(n12578) );
  MUX2_X1 U14928 ( .A(n14371), .B(n12580), .S(n12691), .Z(n12584) );
  NAND2_X1 U14929 ( .A1(n12583), .A2(n12584), .ZN(n12582) );
  MUX2_X1 U14930 ( .A(n14371), .B(n12580), .S(n12496), .Z(n12581) );
  NAND2_X1 U14931 ( .A1(n12582), .A2(n12581), .ZN(n12588) );
  INV_X1 U14932 ( .A(n12583), .ZN(n12586) );
  INV_X1 U14933 ( .A(n12584), .ZN(n12585) );
  NAND2_X1 U14934 ( .A1(n12586), .A2(n12585), .ZN(n12587) );
  MUX2_X1 U14935 ( .A(n14370), .B(n12589), .S(n12496), .Z(n12591) );
  MUX2_X1 U14936 ( .A(n14370), .B(n12589), .S(n12691), .Z(n12590) );
  MUX2_X1 U14937 ( .A(n14369), .B(n12592), .S(n12691), .Z(n12596) );
  NAND2_X1 U14938 ( .A1(n12595), .A2(n12596), .ZN(n12594) );
  MUX2_X1 U14939 ( .A(n14369), .B(n12592), .S(n12496), .Z(n12593) );
  NAND2_X1 U14940 ( .A1(n12594), .A2(n12593), .ZN(n12600) );
  INV_X1 U14941 ( .A(n12595), .ZN(n12598) );
  INV_X1 U14942 ( .A(n12596), .ZN(n12597) );
  NAND2_X1 U14943 ( .A1(n12598), .A2(n12597), .ZN(n12599) );
  NAND2_X1 U14944 ( .A1(n12600), .A2(n12599), .ZN(n12603) );
  MUX2_X1 U14945 ( .A(n14368), .B(n15068), .S(n12496), .Z(n12604) );
  NAND2_X1 U14946 ( .A1(n12603), .A2(n12604), .ZN(n12602) );
  MUX2_X1 U14947 ( .A(n14368), .B(n15068), .S(n12823), .Z(n12601) );
  INV_X1 U14948 ( .A(n12603), .ZN(n12606) );
  INV_X1 U14949 ( .A(n12604), .ZN(n12605) );
  NAND2_X1 U14950 ( .A1(n12606), .A2(n12605), .ZN(n12607) );
  MUX2_X1 U14951 ( .A(n14367), .B(n12608), .S(n12823), .Z(n12612) );
  MUX2_X1 U14952 ( .A(n14367), .B(n12608), .S(n12827), .Z(n12609) );
  MUX2_X1 U14953 ( .A(n14366), .B(n12957), .S(n12827), .Z(n12617) );
  NAND2_X1 U14954 ( .A1(n14366), .A2(n12496), .ZN(n12610) );
  OAI211_X1 U14955 ( .C1(n14300), .C2(n12827), .A(n12617), .B(n12610), .ZN(
        n12611) );
  NAND2_X1 U14956 ( .A1(n12893), .A2(n12613), .ZN(n12614) );
  NAND2_X1 U14957 ( .A1(n12614), .A2(n12496), .ZN(n12622) );
  NAND2_X1 U14958 ( .A1(n12624), .A2(n12615), .ZN(n12616) );
  NAND2_X1 U14959 ( .A1(n12616), .A2(n12823), .ZN(n12621) );
  INV_X1 U14960 ( .A(n12617), .ZN(n12619) );
  MUX2_X1 U14961 ( .A(n14366), .B(n12957), .S(n12823), .Z(n12618) );
  NAND3_X1 U14962 ( .A1(n12854), .A2(n12619), .A3(n12618), .ZN(n12620) );
  NAND2_X1 U14963 ( .A1(n12623), .A2(n7638), .ZN(n12626) );
  MUX2_X1 U14964 ( .A(n12893), .B(n12624), .S(n12827), .Z(n12625) );
  NAND2_X1 U14965 ( .A1(n12626), .A2(n12625), .ZN(n12648) );
  NAND2_X1 U14966 ( .A1(n12627), .A2(n12819), .ZN(n12630) );
  AOI22_X1 U14967 ( .A1(n12661), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n12660), 
        .B2(n12628), .ZN(n12629) );
  MUX2_X1 U14968 ( .A(n14363), .B(n14807), .S(n12827), .Z(n12684) );
  NAND2_X1 U14969 ( .A1(n12702), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n12637) );
  INV_X1 U14970 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n14685) );
  OR2_X1 U14971 ( .A1(n12664), .A2(n14685), .ZN(n12636) );
  INV_X1 U14972 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n12631) );
  NAND2_X1 U14973 ( .A1(n12632), .A2(n12631), .ZN(n12633) );
  NAND2_X1 U14974 ( .A1(n12666), .A2(n12633), .ZN(n14684) );
  OR2_X1 U14975 ( .A1(n12786), .A2(n14684), .ZN(n12635) );
  OR2_X1 U14976 ( .A1(n12670), .A2(n14802), .ZN(n12634) );
  NAND4_X1 U14977 ( .A1(n12637), .A2(n12636), .A3(n12635), .A4(n12634), .ZN(
        n14362) );
  NOR2_X1 U14978 ( .A1(n14363), .A2(n12823), .ZN(n12679) );
  AOI21_X1 U14979 ( .B1(n12684), .B2(n14362), .A(n12679), .ZN(n12646) );
  NAND2_X1 U14980 ( .A1(n12638), .A2(n12819), .ZN(n12640) );
  AOI22_X1 U14981 ( .A1(n12661), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n12660), 
        .B2(n14467), .ZN(n12639) );
  INV_X1 U14982 ( .A(n14683), .ZN(n14859) );
  NAND2_X1 U14983 ( .A1(n14362), .A2(n12823), .ZN(n12676) );
  OR2_X1 U14984 ( .A1(n14807), .A2(n12676), .ZN(n12642) );
  INV_X1 U14985 ( .A(n14362), .ZN(n14701) );
  NAND2_X1 U14986 ( .A1(n12679), .A2(n14701), .ZN(n12641) );
  AND2_X1 U14987 ( .A1(n12642), .A2(n12641), .ZN(n12682) );
  NAND2_X1 U14988 ( .A1(n12684), .A2(n14701), .ZN(n12643) );
  OR2_X1 U14989 ( .A1(n14807), .A2(n12827), .ZN(n12675) );
  NAND2_X1 U14990 ( .A1(n12643), .A2(n12675), .ZN(n12644) );
  NAND2_X1 U14991 ( .A1(n12644), .A2(n14859), .ZN(n12645) );
  OAI211_X1 U14992 ( .C1(n12646), .C2(n14859), .A(n12682), .B(n12645), .ZN(
        n12647) );
  NAND2_X1 U14993 ( .A1(n12648), .A2(n12647), .ZN(n12690) );
  NAND2_X1 U14994 ( .A1(n12649), .A2(n12819), .ZN(n12651) );
  AOI22_X1 U14995 ( .A1(n12661), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n14483), 
        .B2(n12660), .ZN(n12650) );
  NAND2_X1 U14996 ( .A1(n12668), .A2(n12652), .ZN(n12653) );
  NAND2_X1 U14997 ( .A1(n12700), .A2(n12653), .ZN(n14646) );
  INV_X1 U14998 ( .A(n14646), .ZN(n14231) );
  NAND2_X1 U14999 ( .A1(n12810), .A2(n14231), .ZN(n12658) );
  INV_X1 U15000 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n12654) );
  OR2_X1 U15001 ( .A1(n12664), .A2(n12654), .ZN(n12657) );
  INV_X1 U15002 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14790) );
  OR2_X1 U15003 ( .A1(n12670), .A2(n14790), .ZN(n12656) );
  INV_X1 U15004 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n14850) );
  OR2_X1 U15005 ( .A1(n10990), .A2(n14850), .ZN(n12655) );
  NAND4_X1 U15006 ( .A1(n12658), .A2(n12657), .A3(n12656), .A4(n12655), .ZN(
        n14619) );
  AOI22_X1 U15007 ( .A1(n12661), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n12660), 
        .B2(n14474), .ZN(n12662) );
  NAND2_X1 U15008 ( .A1(n12702), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n12674) );
  INV_X1 U15009 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n14670) );
  OR2_X1 U15010 ( .A1(n12664), .A2(n14670), .ZN(n12673) );
  NAND2_X1 U15011 ( .A1(n12666), .A2(n12665), .ZN(n12667) );
  NAND2_X1 U15012 ( .A1(n12668), .A2(n12667), .ZN(n14669) );
  OR2_X1 U15013 ( .A1(n12753), .A2(n14669), .ZN(n12672) );
  INV_X1 U15014 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n12669) );
  OR2_X1 U15015 ( .A1(n12670), .A2(n12669), .ZN(n12671) );
  NAND4_X1 U15016 ( .A1(n12674), .A2(n12673), .A3(n12672), .A4(n12671), .ZN(
        n14361) );
  INV_X1 U15017 ( .A(n14361), .ZN(n14680) );
  XNOR2_X1 U15018 ( .A(n14794), .B(n14680), .ZN(n14662) );
  INV_X1 U15019 ( .A(n12675), .ZN(n12678) );
  INV_X1 U15020 ( .A(n12676), .ZN(n12677) );
  AOI21_X1 U15021 ( .B1(n12684), .B2(n12678), .A(n12677), .ZN(n12687) );
  NAND2_X1 U15022 ( .A1(n12684), .A2(n12679), .ZN(n12680) );
  OAI21_X1 U15023 ( .B1(n12823), .B2(n14362), .A(n12680), .ZN(n12681) );
  NAND2_X1 U15024 ( .A1(n12681), .A2(n14683), .ZN(n12686) );
  INV_X1 U15025 ( .A(n12682), .ZN(n12683) );
  NAND2_X1 U15026 ( .A1(n12684), .A2(n12683), .ZN(n12685) );
  OAI211_X1 U15027 ( .C1(n12687), .C2(n14683), .A(n12686), .B(n12685), .ZN(
        n12688) );
  NAND2_X1 U15028 ( .A1(n12690), .A2(n12689), .ZN(n12699) );
  NAND2_X1 U15029 ( .A1(n14668), .A2(n14361), .ZN(n12899) );
  NAND3_X1 U15030 ( .A1(n14794), .A2(n14680), .A3(n12691), .ZN(n12692) );
  OAI21_X1 U15031 ( .B1(n12899), .B2(n12823), .A(n12692), .ZN(n12696) );
  AND2_X1 U15032 ( .A1(n14619), .A2(n12827), .ZN(n12694) );
  NOR2_X1 U15033 ( .A1(n14619), .A2(n12827), .ZN(n12693) );
  MUX2_X1 U15034 ( .A(n12694), .B(n12693), .S(n14650), .Z(n12695) );
  NAND2_X1 U15035 ( .A1(n12699), .A2(n12698), .ZN(n12713) );
  INV_X1 U15036 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n14285) );
  NAND2_X1 U15037 ( .A1(n12700), .A2(n14285), .ZN(n12701) );
  NAND2_X1 U15038 ( .A1(n12716), .A2(n12701), .ZN(n14631) );
  NAND2_X1 U15039 ( .A1(n12812), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n12704) );
  NAND2_X1 U15040 ( .A1(n12702), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n12703) );
  AND2_X1 U15041 ( .A1(n12704), .A2(n12703), .ZN(n12706) );
  NAND2_X1 U15042 ( .A1(n12811), .A2(P1_REG1_REG_20__SCAN_IN), .ZN(n12705) );
  OAI211_X1 U15043 ( .C1(n14631), .C2(n12786), .A(n12706), .B(n12705), .ZN(
        n14610) );
  INV_X1 U15044 ( .A(n14610), .ZN(n14239) );
  OR2_X1 U15045 ( .A1(n12820), .A2(n12708), .ZN(n12709) );
  INV_X1 U15046 ( .A(n14633), .ZN(n14780) );
  MUX2_X1 U15047 ( .A(n14239), .B(n14780), .S(n12827), .Z(n12712) );
  MUX2_X1 U15048 ( .A(n14610), .B(n14633), .S(n12823), .Z(n12711) );
  NAND2_X1 U15049 ( .A1(n12713), .A2(n12712), .ZN(n12714) );
  NAND2_X1 U15050 ( .A1(n12715), .A2(n12714), .ZN(n12727) );
  INV_X1 U15051 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n12720) );
  INV_X1 U15052 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n14238) );
  NAND2_X1 U15053 ( .A1(n12716), .A2(n14238), .ZN(n12717) );
  NAND2_X1 U15054 ( .A1(n12729), .A2(n12717), .ZN(n14602) );
  OR2_X1 U15055 ( .A1(n14602), .A2(n12786), .ZN(n12719) );
  AOI22_X1 U15056 ( .A1(n12811), .A2(P1_REG1_REG_21__SCAN_IN), .B1(n12812), 
        .B2(P1_REG2_REG_21__SCAN_IN), .ZN(n12718) );
  OAI211_X1 U15057 ( .C1(n10990), .C2(n12720), .A(n12719), .B(n12718), .ZN(
        n14621) );
  OR2_X1 U15058 ( .A1(n12722), .A2(n12721), .ZN(n12725) );
  OR2_X1 U15059 ( .A1(n12820), .A2(n12723), .ZN(n12724) );
  MUX2_X1 U15060 ( .A(n14621), .B(n14601), .S(n12823), .Z(n12728) );
  MUX2_X1 U15061 ( .A(n14621), .B(n14601), .S(n12827), .Z(n12726) );
  NAND2_X1 U15062 ( .A1(n12729), .A2(n14305), .ZN(n12730) );
  AND2_X1 U15063 ( .A1(n12751), .A2(n12730), .ZN(n14592) );
  NAND2_X1 U15064 ( .A1(n14592), .A2(n12810), .ZN(n12735) );
  INV_X1 U15065 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n14841) );
  NAND2_X1 U15066 ( .A1(n12811), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n12732) );
  NAND2_X1 U15067 ( .A1(n12812), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n12731) );
  OAI211_X1 U15068 ( .C1(n14841), .C2(n10990), .A(n12732), .B(n12731), .ZN(
        n12733) );
  INV_X1 U15069 ( .A(n12733), .ZN(n12734) );
  OR2_X1 U15070 ( .A1(n12736), .A2(n9213), .ZN(n12737) );
  XNOR2_X1 U15071 ( .A(n12737), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14877) );
  INV_X1 U15072 ( .A(n14843), .ZN(n14591) );
  MUX2_X1 U15073 ( .A(n14772), .B(n14591), .S(n12827), .Z(n12740) );
  MUX2_X1 U15074 ( .A(n14607), .B(n14843), .S(n12823), .Z(n12739) );
  MUX2_X1 U15075 ( .A(n14360), .B(n13039), .S(n12827), .Z(n12742) );
  OAI21_X1 U15076 ( .B1(n12745), .B2(n12744), .A(n12743), .ZN(n12761) );
  NAND2_X1 U15077 ( .A1(n12746), .A2(n12819), .ZN(n12749) );
  OR2_X1 U15078 ( .A1(n12820), .A2(n12747), .ZN(n12748) );
  INV_X1 U15079 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n14220) );
  INV_X1 U15080 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n12750) );
  OAI21_X1 U15081 ( .B1(n12751), .B2(n14220), .A(n12750), .ZN(n12752) );
  NAND2_X1 U15082 ( .A1(n12763), .A2(n12752), .ZN(n14554) );
  OR2_X1 U15083 ( .A1(n14554), .A2(n12753), .ZN(n12759) );
  INV_X1 U15084 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n12756) );
  NAND2_X1 U15085 ( .A1(n12812), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n12755) );
  NAND2_X1 U15086 ( .A1(n12811), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n12754) );
  OAI211_X1 U15087 ( .C1(n6668), .C2(n12756), .A(n12755), .B(n12754), .ZN(
        n12757) );
  INV_X1 U15088 ( .A(n12757), .ZN(n12758) );
  NAND2_X1 U15089 ( .A1(n12759), .A2(n12758), .ZN(n14359) );
  MUX2_X1 U15090 ( .A(n14757), .B(n14359), .S(n12823), .Z(n12762) );
  MUX2_X1 U15091 ( .A(n14359), .B(n14757), .S(n12823), .Z(n12760) );
  NAND2_X1 U15092 ( .A1(n12763), .A2(n14250), .ZN(n12764) );
  AND2_X1 U15093 ( .A1(n12784), .A2(n12764), .ZN(n14537) );
  NAND2_X1 U15094 ( .A1(n14537), .A2(n12810), .ZN(n12770) );
  INV_X1 U15095 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n12767) );
  NAND2_X1 U15096 ( .A1(n12812), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n12766) );
  NAND2_X1 U15097 ( .A1(n12811), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n12765) );
  OAI211_X1 U15098 ( .C1(n10990), .C2(n12767), .A(n12766), .B(n12765), .ZN(
        n12768) );
  INV_X1 U15099 ( .A(n12768), .ZN(n12769) );
  NAND2_X1 U15100 ( .A1(n12770), .A2(n12769), .ZN(n14524) );
  NAND2_X1 U15101 ( .A1(n12771), .A2(n12819), .ZN(n12774) );
  OR2_X1 U15102 ( .A1(n12820), .A2(n12772), .ZN(n12773) );
  MUX2_X1 U15103 ( .A(n14524), .B(n14751), .S(n12823), .Z(n12778) );
  MUX2_X1 U15104 ( .A(n14751), .B(n14524), .S(n12823), .Z(n12775) );
  NAND2_X1 U15105 ( .A1(n12776), .A2(n12775), .ZN(n12782) );
  INV_X1 U15106 ( .A(n12777), .ZN(n12780) );
  INV_X1 U15107 ( .A(n12778), .ZN(n12779) );
  NAND2_X1 U15108 ( .A1(n12780), .A2(n12779), .ZN(n12781) );
  INV_X1 U15109 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n12783) );
  NAND2_X1 U15110 ( .A1(n12784), .A2(n12783), .ZN(n12785) );
  NAND2_X1 U15111 ( .A1(n12798), .A2(n12785), .ZN(n14334) );
  OR2_X1 U15112 ( .A1(n14334), .A2(n12786), .ZN(n12791) );
  INV_X1 U15113 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n14832) );
  NAND2_X1 U15114 ( .A1(n12811), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n12788) );
  NAND2_X1 U15115 ( .A1(n12812), .A2(P1_REG2_REG_26__SCAN_IN), .ZN(n12787) );
  OAI211_X1 U15116 ( .C1(n14832), .C2(n6668), .A(n12788), .B(n12787), .ZN(
        n12789) );
  INV_X1 U15117 ( .A(n12789), .ZN(n12790) );
  NAND2_X1 U15118 ( .A1(n12792), .A2(n12819), .ZN(n12795) );
  OR2_X1 U15119 ( .A1(n12820), .A2(n12793), .ZN(n12794) );
  MUX2_X1 U15120 ( .A(n14358), .B(n14329), .S(n12827), .Z(n12797) );
  MUX2_X1 U15121 ( .A(n14358), .B(n14329), .S(n12823), .Z(n12796) );
  NAND2_X1 U15122 ( .A1(n12798), .A2(n14210), .ZN(n12799) );
  NAND2_X1 U15123 ( .A1(n14511), .A2(n12810), .ZN(n12804) );
  INV_X1 U15124 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n14828) );
  NAND2_X1 U15125 ( .A1(n12811), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n12801) );
  NAND2_X1 U15126 ( .A1(n12812), .A2(P1_REG2_REG_27__SCAN_IN), .ZN(n12800) );
  OAI211_X1 U15127 ( .C1(n14828), .C2(n10990), .A(n12801), .B(n12800), .ZN(
        n12802) );
  INV_X1 U15128 ( .A(n12802), .ZN(n12803) );
  NAND2_X1 U15129 ( .A1(n12887), .A2(n12819), .ZN(n12806) );
  OR2_X1 U15130 ( .A1(n12820), .A2(n14875), .ZN(n12805) );
  MUX2_X1 U15131 ( .A(n14357), .B(n14508), .S(n12823), .Z(n12808) );
  MUX2_X1 U15132 ( .A(n14357), .B(n14508), .S(n12827), .Z(n12807) );
  INV_X1 U15133 ( .A(n12808), .ZN(n12809) );
  XNOR2_X1 U15134 ( .A(n13105), .B(P1_REG3_REG_28__SCAN_IN), .ZN(n13093) );
  NAND2_X1 U15135 ( .A1(n13093), .A2(n12810), .ZN(n12818) );
  INV_X1 U15136 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n12815) );
  NAND2_X1 U15137 ( .A1(n12811), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n12814) );
  NAND2_X1 U15138 ( .A1(n12812), .A2(P1_REG2_REG_28__SCAN_IN), .ZN(n12813) );
  OAI211_X1 U15139 ( .C1(n12815), .C2(n10990), .A(n12814), .B(n12813), .ZN(
        n12816) );
  INV_X1 U15140 ( .A(n12816), .ZN(n12817) );
  NAND2_X1 U15141 ( .A1(n14869), .A2(n12819), .ZN(n12822) );
  INV_X1 U15142 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n14871) );
  OR2_X1 U15143 ( .A1(n12820), .A2(n14871), .ZN(n12821) );
  MUX2_X1 U15144 ( .A(n14356), .B(n14734), .S(n12827), .Z(n12825) );
  MUX2_X1 U15145 ( .A(n14356), .B(n14734), .S(n12823), .Z(n12824) );
  INV_X1 U15146 ( .A(n12825), .ZN(n12826) );
  INV_X1 U15147 ( .A(n12830), .ZN(n12832) );
  INV_X1 U15148 ( .A(n13101), .ZN(n14726) );
  MUX2_X1 U15149 ( .A(n13092), .B(n14726), .S(n12827), .Z(n12828) );
  AOI21_X1 U15150 ( .B1(n12830), .B2(n12829), .A(n12828), .ZN(n12831) );
  AOI21_X1 U15151 ( .B1(n12833), .B2(n12832), .A(n12831), .ZN(n12836) );
  XOR2_X1 U15152 ( .A(n14491), .B(n14488), .Z(n12875) );
  XOR2_X1 U15153 ( .A(n14354), .B(n14497), .Z(n12861) );
  XNOR2_X1 U15154 ( .A(n13101), .B(n13092), .ZN(n13114) );
  XNOR2_X2 U15155 ( .A(n14734), .B(n14356), .ZN(n12939) );
  NAND2_X1 U15156 ( .A1(n14751), .A2(n14546), .ZN(n12907) );
  OR2_X1 U15157 ( .A1(n14751), .A2(n14546), .ZN(n12837) );
  XNOR2_X1 U15158 ( .A(n13039), .B(n14360), .ZN(n14569) );
  INV_X1 U15159 ( .A(n14569), .ZN(n14562) );
  XNOR2_X1 U15160 ( .A(n14843), .B(n14772), .ZN(n14587) );
  INV_X1 U15161 ( .A(n14587), .ZN(n14580) );
  XNOR2_X1 U15162 ( .A(n14633), .B(n14610), .ZN(n14627) );
  INV_X1 U15163 ( .A(n14627), .ZN(n12856) );
  XNOR2_X1 U15164 ( .A(n14807), .B(n14681), .ZN(n14697) );
  OR2_X1 U15165 ( .A1(n14683), .A2(n14362), .ZN(n12920) );
  NAND2_X1 U15166 ( .A1(n14683), .A2(n14362), .ZN(n12919) );
  NAND2_X1 U15167 ( .A1(n12920), .A2(n12919), .ZN(n14677) );
  NOR4_X1 U15168 ( .A1(n11419), .A2(n12840), .A3(n6859), .A4(n12838), .ZN(
        n12842) );
  NOR4_X1 U15169 ( .A1(n12846), .A2(n12845), .A3(n12844), .A4(n12843), .ZN(
        n12848) );
  NAND4_X1 U15170 ( .A1(n12849), .A2(n12848), .A3(n7610), .A4(n7607), .ZN(
        n12850) );
  NOR3_X1 U15171 ( .A1(n12852), .A2(n12851), .A3(n12850), .ZN(n12853) );
  NAND4_X1 U15172 ( .A1(n14677), .A2(n12854), .A3(n12915), .A4(n12853), .ZN(
        n12855) );
  NOR4_X1 U15173 ( .A1(n12856), .A2(n14662), .A3(n14697), .A4(n12855), .ZN(
        n12857) );
  XNOR2_X1 U15174 ( .A(n14601), .B(n14621), .ZN(n14609) );
  NAND4_X1 U15175 ( .A1(n14580), .A2(n12857), .A3(n12697), .A4(n14609), .ZN(
        n12858) );
  NOR4_X1 U15176 ( .A1(n14531), .A2(n14550), .A3(n14562), .A4(n12858), .ZN(
        n12859) );
  INV_X1 U15177 ( .A(n14358), .ZN(n12908) );
  XNOR2_X1 U15178 ( .A(n14329), .B(n12908), .ZN(n12932) );
  NAND4_X1 U15179 ( .A1(n12939), .A2(n12859), .A3(n14504), .A4(n14520), .ZN(
        n12860) );
  XNOR2_X1 U15180 ( .A(n12862), .B(n14483), .ZN(n12872) );
  NOR3_X1 U15181 ( .A1(n14820), .A2(n14491), .A3(n12863), .ZN(n12866) );
  NOR3_X1 U15182 ( .A1(n12865), .A2(n14491), .A3(n12874), .ZN(n12864) );
  AOI21_X1 U15183 ( .B1(n12866), .B2(n12865), .A(n12864), .ZN(n12870) );
  XOR2_X1 U15184 ( .A(n12874), .B(n12867), .Z(n12868) );
  NAND4_X1 U15185 ( .A1(n12868), .A2(n14820), .A3(n14491), .A4(n12871), .ZN(
        n12869) );
  OAI211_X1 U15186 ( .C1(n12872), .C2(n12871), .A(n12870), .B(n12869), .ZN(
        n12873) );
  INV_X1 U15187 ( .A(n12873), .ZN(n12876) );
  INV_X1 U15188 ( .A(n12878), .ZN(n12884) );
  NAND4_X1 U15189 ( .A1(n12880), .A2(n13102), .A3(n14620), .A4(n12879), .ZN(
        n12881) );
  OAI211_X1 U15190 ( .C1(n14878), .C2(n12883), .A(n12881), .B(P1_B_REG_SCAN_IN), .ZN(n12882) );
  OAI21_X1 U15191 ( .B1(n12884), .B2(n12883), .A(n12882), .ZN(P1_U3242) );
  INV_X1 U15192 ( .A(n12885), .ZN(n13122) );
  OAI222_X1 U15193 ( .A1(n14874), .A2(n13122), .B1(P1_U3086), .B2(n10481), 
        .C1(n12886), .C2(n14876), .ZN(P1_U3325) );
  INV_X1 U15194 ( .A(n12887), .ZN(n14873) );
  OAI222_X1 U15195 ( .A1(n14201), .A2(n12888), .B1(n14196), .B2(n14873), .C1(
        P2_U3088), .C2(n9668), .ZN(P2_U3300) );
  INV_X1 U15196 ( .A(n12889), .ZN(n12891) );
  OAI222_X1 U15197 ( .A1(n12892), .A2(P3_U3151), .B1(n13688), .B2(n12891), 
        .C1(n12890), .C2(n13690), .ZN(P3_U3271) );
  NAND2_X1 U15198 ( .A1(n14807), .A2(n14681), .ZN(n12895) );
  OR2_X1 U15199 ( .A1(n14683), .A2(n14701), .ZN(n12896) );
  NAND2_X1 U15200 ( .A1(n14683), .A2(n14701), .ZN(n12897) );
  INV_X1 U15201 ( .A(n14662), .ZN(n12898) );
  NAND2_X1 U15202 ( .A1(n14650), .A2(n14658), .ZN(n12901) );
  INV_X1 U15203 ( .A(n14621), .ZN(n14286) );
  OR2_X1 U15204 ( .A1(n14601), .A2(n14286), .ZN(n14581) );
  AND2_X1 U15205 ( .A1(n14580), .A2(n14581), .ZN(n12902) );
  OR2_X1 U15206 ( .A1(n14843), .A2(n14772), .ZN(n12903) );
  INV_X1 U15207 ( .A(n14360), .ZN(n14545) );
  NAND2_X1 U15208 ( .A1(n13039), .A2(n14545), .ZN(n12904) );
  OR2_X1 U15209 ( .A1(n14757), .A2(n6822), .ZN(n12906) );
  AND2_X1 U15210 ( .A1(n14329), .A2(n12908), .ZN(n12909) );
  AOI21_X2 U15211 ( .B1(n14521), .B2(n14520), .A(n12909), .ZN(n14501) );
  NAND2_X1 U15212 ( .A1(n14355), .A2(n14771), .ZN(n12911) );
  NAND2_X1 U15213 ( .A1(n14357), .A2(n14620), .ZN(n12910) );
  INV_X1 U15214 ( .A(n12915), .ZN(n12916) );
  OR2_X1 U15215 ( .A1(n14810), .A2(n14364), .ZN(n12917) );
  OR2_X1 U15216 ( .A1(n14807), .A2(n14363), .ZN(n12918) );
  NAND2_X1 U15217 ( .A1(n14794), .A2(n14361), .ZN(n12921) );
  NAND2_X1 U15218 ( .A1(n14668), .A2(n14680), .ZN(n12922) );
  NAND2_X1 U15219 ( .A1(n14648), .A2(n14642), .ZN(n12924) );
  OR2_X1 U15220 ( .A1(n14650), .A2(n14619), .ZN(n12923) );
  NAND2_X1 U15221 ( .A1(n12924), .A2(n12923), .ZN(n14626) );
  INV_X1 U15222 ( .A(n14626), .ZN(n12925) );
  NAND2_X1 U15223 ( .A1(n14633), .A2(n14610), .ZN(n12926) );
  INV_X1 U15224 ( .A(n14609), .ZN(n12927) );
  OR2_X1 U15225 ( .A1(n14601), .A2(n14621), .ZN(n12928) );
  NAND2_X1 U15226 ( .A1(n14843), .A2(n14607), .ZN(n12929) );
  NAND2_X1 U15227 ( .A1(n14586), .A2(n12929), .ZN(n14566) );
  NAND2_X1 U15228 ( .A1(n13039), .A2(n14360), .ZN(n12930) );
  OR2_X1 U15229 ( .A1(n14757), .A2(n14359), .ZN(n12931) );
  NAND2_X1 U15230 ( .A1(n14516), .A2(n12932), .ZN(n12934) );
  NAND2_X1 U15231 ( .A1(n14329), .A2(n14358), .ZN(n12933) );
  NAND2_X1 U15232 ( .A1(n12934), .A2(n12933), .ZN(n14505) );
  INV_X1 U15233 ( .A(n14505), .ZN(n12936) );
  INV_X1 U15234 ( .A(n14734), .ZN(n13110) );
  INV_X1 U15235 ( .A(n14751), .ZN(n14254) );
  NOR2_X1 U15236 ( .A1(n14651), .A2(n14633), .ZN(n14628) );
  INV_X1 U15237 ( .A(n14601), .ZN(n14847) );
  AOI21_X1 U15238 ( .B1(n14734), .B2(n14509), .A(n14781), .ZN(n12940) );
  AND2_X1 U15239 ( .A1(n13100), .A2(n12940), .ZN(n14733) );
  NAND2_X1 U15240 ( .A1(n14733), .A2(n14713), .ZN(n12942) );
  AOI22_X1 U15241 ( .A1(n13093), .A2(n15142), .B1(P1_REG2_REG_28__SCAN_IN), 
        .B2(n15143), .ZN(n12941) );
  OAI211_X1 U15242 ( .C1(n13110), .C2(n14709), .A(n12942), .B(n12941), .ZN(
        n12943) );
  AOI21_X1 U15243 ( .B1(n14732), .B2(n14649), .A(n12943), .ZN(n12944) );
  OAI21_X1 U15244 ( .B1(n14736), .B2(n15143), .A(n12944), .ZN(P1_U3265) );
  INV_X1 U15245 ( .A(n12945), .ZN(n12948) );
  OAI222_X1 U15246 ( .A1(n13688), .A2(n12948), .B1(n6812), .B2(P3_U3151), .C1(
        n12946), .C2(n13690), .ZN(P3_U3267) );
  INV_X1 U15247 ( .A(n12949), .ZN(n14195) );
  INV_X1 U15248 ( .A(n12952), .ZN(n12954) );
  NAND2_X1 U15249 ( .A1(n12955), .A2(n6778), .ZN(n14292) );
  AND2_X1 U15250 ( .A1(n14366), .A2(n13059), .ZN(n12956) );
  AOI21_X1 U15251 ( .B1(n12957), .B2(n13038), .A(n12956), .ZN(n12964) );
  AOI22_X1 U15252 ( .A1(n12957), .A2(n13086), .B1(n13085), .B2(n14366), .ZN(
        n12958) );
  XNOR2_X1 U15253 ( .A(n12958), .B(n10886), .ZN(n12963) );
  XOR2_X1 U15254 ( .A(n12964), .B(n12963), .Z(n14291) );
  NAND2_X1 U15255 ( .A1(n15050), .A2(n13086), .ZN(n12960) );
  NAND2_X1 U15256 ( .A1(n14365), .A2(n13085), .ZN(n12959) );
  NAND2_X1 U15257 ( .A1(n12960), .A2(n12959), .ZN(n12961) );
  XNOR2_X1 U15258 ( .A(n12961), .B(n10886), .ZN(n12970) );
  AND2_X1 U15259 ( .A1(n14365), .A2(n13059), .ZN(n12962) );
  AOI21_X1 U15260 ( .B1(n15050), .B2(n13038), .A(n12962), .ZN(n12968) );
  XNOR2_X1 U15261 ( .A(n12970), .B(n12968), .ZN(n15042) );
  INV_X1 U15262 ( .A(n12963), .ZN(n12966) );
  INV_X1 U15263 ( .A(n12964), .ZN(n12965) );
  NAND2_X1 U15264 ( .A1(n12966), .A2(n12965), .ZN(n15043) );
  INV_X1 U15265 ( .A(n12968), .ZN(n12969) );
  NAND2_X1 U15266 ( .A1(n14810), .A2(n13086), .ZN(n12972) );
  NAND2_X1 U15267 ( .A1(n14364), .A2(n13085), .ZN(n12971) );
  NAND2_X1 U15268 ( .A1(n12972), .A2(n12971), .ZN(n12973) );
  XNOR2_X1 U15269 ( .A(n12973), .B(n10886), .ZN(n12976) );
  OAI22_X1 U15270 ( .A1(n14353), .A2(n12975), .B1(n15040), .B2(n12974), .ZN(
        n14343) );
  INV_X1 U15271 ( .A(n12976), .ZN(n12977) );
  OR2_X1 U15272 ( .A1(n12978), .A2(n12977), .ZN(n12979) );
  NAND2_X1 U15273 ( .A1(n14342), .A2(n12979), .ZN(n14257) );
  AOI22_X1 U15274 ( .A1(n14807), .A2(n13086), .B1(n13085), .B2(n14363), .ZN(
        n12980) );
  XNOR2_X1 U15275 ( .A(n12980), .B(n10886), .ZN(n12982) );
  AOI22_X1 U15276 ( .A1(n14807), .A2(n13070), .B1(n13087), .B2(n14363), .ZN(
        n12981) );
  XNOR2_X1 U15277 ( .A(n12982), .B(n12981), .ZN(n14258) );
  NAND2_X1 U15278 ( .A1(n12982), .A2(n12981), .ZN(n12983) );
  NAND2_X1 U15279 ( .A1(n14683), .A2(n13086), .ZN(n12985) );
  NAND2_X1 U15280 ( .A1(n14362), .A2(n13085), .ZN(n12984) );
  NAND2_X1 U15281 ( .A1(n12985), .A2(n12984), .ZN(n12986) );
  XNOR2_X1 U15282 ( .A(n12986), .B(n10886), .ZN(n12989) );
  NAND2_X1 U15283 ( .A1(n14683), .A2(n13085), .ZN(n12988) );
  NAND2_X1 U15284 ( .A1(n14362), .A2(n13087), .ZN(n12987) );
  NAND2_X1 U15285 ( .A1(n12988), .A2(n12987), .ZN(n12990) );
  NAND2_X1 U15286 ( .A1(n12989), .A2(n12990), .ZN(n14264) );
  INV_X1 U15287 ( .A(n12989), .ZN(n12992) );
  INV_X1 U15288 ( .A(n12990), .ZN(n12991) );
  NAND2_X1 U15289 ( .A1(n12992), .A2(n12991), .ZN(n14265) );
  NAND2_X1 U15290 ( .A1(n14794), .A2(n13086), .ZN(n12994) );
  NAND2_X1 U15291 ( .A1(n14361), .A2(n13070), .ZN(n12993) );
  NAND2_X1 U15292 ( .A1(n12994), .A2(n12993), .ZN(n12995) );
  XNOR2_X1 U15293 ( .A(n12995), .B(n10886), .ZN(n13000) );
  AOI22_X1 U15294 ( .A1(n14794), .A2(n13070), .B1(n13059), .B2(n14361), .ZN(
        n12998) );
  XNOR2_X1 U15295 ( .A(n13000), .B(n12998), .ZN(n14312) );
  NAND2_X1 U15296 ( .A1(n14310), .A2(n14312), .ZN(n14224) );
  AOI22_X1 U15297 ( .A1(n14650), .A2(n13086), .B1(n13085), .B2(n14619), .ZN(
        n12996) );
  XNOR2_X1 U15298 ( .A(n12996), .B(n10886), .ZN(n13017) );
  AND2_X1 U15299 ( .A1(n14619), .A2(n13059), .ZN(n12997) );
  AOI21_X1 U15300 ( .B1(n14650), .B2(n13085), .A(n12997), .ZN(n13018) );
  XNOR2_X1 U15301 ( .A(n13017), .B(n13018), .ZN(n14225) );
  INV_X1 U15302 ( .A(n12998), .ZN(n12999) );
  NOR2_X1 U15303 ( .A1(n13000), .A2(n12999), .ZN(n14226) );
  NOR2_X1 U15304 ( .A1(n14225), .A2(n14226), .ZN(n14228) );
  NAND2_X1 U15305 ( .A1(n14633), .A2(n13086), .ZN(n13002) );
  NAND2_X1 U15306 ( .A1(n14610), .A2(n13085), .ZN(n13001) );
  NAND2_X1 U15307 ( .A1(n13002), .A2(n13001), .ZN(n13003) );
  XNOR2_X1 U15308 ( .A(n13003), .B(n10886), .ZN(n13007) );
  AND2_X1 U15309 ( .A1(n14610), .A2(n13059), .ZN(n13004) );
  AOI21_X1 U15310 ( .B1(n14633), .B2(n13085), .A(n13004), .ZN(n13006) );
  INV_X1 U15311 ( .A(n13006), .ZN(n13005) );
  NAND2_X1 U15312 ( .A1(n13007), .A2(n13005), .ZN(n13021) );
  INV_X1 U15313 ( .A(n13021), .ZN(n13008) );
  XNOR2_X1 U15314 ( .A(n13007), .B(n13006), .ZN(n14283) );
  AND2_X1 U15315 ( .A1(n14228), .A2(n13016), .ZN(n13009) );
  NAND2_X1 U15316 ( .A1(n14601), .A2(n13086), .ZN(n13011) );
  NAND2_X1 U15317 ( .A1(n14621), .A2(n13070), .ZN(n13010) );
  NAND2_X1 U15318 ( .A1(n13011), .A2(n13010), .ZN(n13012) );
  XNOR2_X1 U15319 ( .A(n13012), .B(n13057), .ZN(n13015) );
  AND2_X1 U15320 ( .A1(n14621), .A2(n13059), .ZN(n13013) );
  AOI21_X1 U15321 ( .B1(n14601), .B2(n13085), .A(n13013), .ZN(n13014) );
  NAND2_X1 U15322 ( .A1(n13015), .A2(n13014), .ZN(n14301) );
  OAI21_X1 U15323 ( .B1(n13015), .B2(n13014), .A(n14301), .ZN(n14236) );
  INV_X1 U15324 ( .A(n14236), .ZN(n13024) );
  INV_X1 U15325 ( .A(n13016), .ZN(n13023) );
  INV_X1 U15326 ( .A(n13017), .ZN(n13020) );
  INV_X1 U15327 ( .A(n13018), .ZN(n13019) );
  NAND2_X1 U15328 ( .A1(n13020), .A2(n13019), .ZN(n14281) );
  AND2_X1 U15329 ( .A1(n14281), .A2(n13021), .ZN(n13022) );
  AND2_X1 U15330 ( .A1(n13024), .A2(n14234), .ZN(n13025) );
  OAI22_X1 U15331 ( .A1(n14843), .A2(n11858), .B1(n14607), .B2(n13026), .ZN(
        n13027) );
  XNOR2_X1 U15332 ( .A(n13027), .B(n13057), .ZN(n13029) );
  AND2_X1 U15333 ( .A1(n14772), .A2(n13059), .ZN(n13028) );
  AOI21_X1 U15334 ( .B1(n14591), .B2(n13038), .A(n13028), .ZN(n13030) );
  NAND2_X1 U15335 ( .A1(n13029), .A2(n13030), .ZN(n14215) );
  INV_X1 U15336 ( .A(n13029), .ZN(n13032) );
  INV_X1 U15337 ( .A(n13030), .ZN(n13031) );
  NAND2_X1 U15338 ( .A1(n13032), .A2(n13031), .ZN(n13033) );
  NAND2_X1 U15339 ( .A1(n14214), .A2(n14215), .ZN(n13045) );
  NAND2_X1 U15340 ( .A1(n13039), .A2(n13086), .ZN(n13035) );
  NAND2_X1 U15341 ( .A1(n14360), .A2(n13070), .ZN(n13034) );
  NAND2_X1 U15342 ( .A1(n13035), .A2(n13034), .ZN(n13036) );
  XNOR2_X1 U15343 ( .A(n13036), .B(n13057), .ZN(n13040) );
  AND2_X1 U15344 ( .A1(n14360), .A2(n13059), .ZN(n13037) );
  AOI21_X1 U15345 ( .B1(n13039), .B2(n13038), .A(n13037), .ZN(n13041) );
  NAND2_X1 U15346 ( .A1(n13040), .A2(n13041), .ZN(n14273) );
  INV_X1 U15347 ( .A(n13040), .ZN(n13043) );
  INV_X1 U15348 ( .A(n13041), .ZN(n13042) );
  NAND2_X1 U15349 ( .A1(n13043), .A2(n13042), .ZN(n13044) );
  NAND2_X1 U15350 ( .A1(n13045), .A2(n14216), .ZN(n14218) );
  NAND2_X1 U15351 ( .A1(n14757), .A2(n13086), .ZN(n13047) );
  NAND2_X1 U15352 ( .A1(n14359), .A2(n13070), .ZN(n13046) );
  NAND2_X1 U15353 ( .A1(n13047), .A2(n13046), .ZN(n13048) );
  XNOR2_X1 U15354 ( .A(n13048), .B(n13057), .ZN(n13050) );
  AND2_X1 U15355 ( .A1(n14359), .A2(n13059), .ZN(n13049) );
  AOI21_X1 U15356 ( .B1(n14757), .B2(n13085), .A(n13049), .ZN(n13051) );
  NAND2_X1 U15357 ( .A1(n13050), .A2(n13051), .ZN(n14244) );
  INV_X1 U15358 ( .A(n13050), .ZN(n13053) );
  INV_X1 U15359 ( .A(n13051), .ZN(n13052) );
  NAND2_X1 U15360 ( .A1(n13053), .A2(n13052), .ZN(n13054) );
  NAND2_X1 U15361 ( .A1(n14751), .A2(n13086), .ZN(n13056) );
  NAND2_X1 U15362 ( .A1(n14524), .A2(n13070), .ZN(n13055) );
  NAND2_X1 U15363 ( .A1(n13056), .A2(n13055), .ZN(n13058) );
  XNOR2_X1 U15364 ( .A(n13058), .B(n13057), .ZN(n13061) );
  AND2_X1 U15365 ( .A1(n14524), .A2(n13059), .ZN(n13060) );
  AOI21_X1 U15366 ( .B1(n14751), .B2(n13085), .A(n13060), .ZN(n13062) );
  NAND2_X1 U15367 ( .A1(n13061), .A2(n13062), .ZN(n13066) );
  INV_X1 U15368 ( .A(n13061), .ZN(n13064) );
  INV_X1 U15369 ( .A(n13062), .ZN(n13063) );
  NAND2_X1 U15370 ( .A1(n13064), .A2(n13063), .ZN(n13065) );
  NAND2_X1 U15371 ( .A1(n14246), .A2(n13066), .ZN(n14331) );
  NAND2_X1 U15372 ( .A1(n14329), .A2(n13086), .ZN(n13068) );
  NAND2_X1 U15373 ( .A1(n14358), .A2(n13070), .ZN(n13067) );
  NAND2_X1 U15374 ( .A1(n13068), .A2(n13067), .ZN(n13069) );
  XNOR2_X1 U15375 ( .A(n13069), .B(n10886), .ZN(n13074) );
  NAND2_X1 U15376 ( .A1(n14329), .A2(n13070), .ZN(n13072) );
  NAND2_X1 U15377 ( .A1(n14358), .A2(n13087), .ZN(n13071) );
  NAND2_X1 U15378 ( .A1(n13072), .A2(n13071), .ZN(n13073) );
  NOR2_X1 U15379 ( .A1(n13074), .A2(n13073), .ZN(n13075) );
  AOI21_X1 U15380 ( .B1(n13074), .B2(n13073), .A(n13075), .ZN(n14332) );
  NAND2_X1 U15381 ( .A1(n14331), .A2(n14332), .ZN(n14330) );
  INV_X1 U15382 ( .A(n13075), .ZN(n13076) );
  NAND2_X1 U15383 ( .A1(n14330), .A2(n13076), .ZN(n14205) );
  NAND2_X1 U15384 ( .A1(n14508), .A2(n13086), .ZN(n13078) );
  NAND2_X1 U15385 ( .A1(n14357), .A2(n13085), .ZN(n13077) );
  NAND2_X1 U15386 ( .A1(n13078), .A2(n13077), .ZN(n13079) );
  XNOR2_X1 U15387 ( .A(n13079), .B(n10886), .ZN(n13083) );
  NAND2_X1 U15388 ( .A1(n14508), .A2(n13085), .ZN(n13081) );
  NAND2_X1 U15389 ( .A1(n14357), .A2(n13087), .ZN(n13080) );
  NAND2_X1 U15390 ( .A1(n13081), .A2(n13080), .ZN(n13082) );
  NOR2_X1 U15391 ( .A1(n13083), .A2(n13082), .ZN(n13084) );
  AOI21_X1 U15392 ( .B1(n13083), .B2(n13082), .A(n13084), .ZN(n14206) );
  NAND2_X1 U15393 ( .A1(n14205), .A2(n14206), .ZN(n14204) );
  AOI22_X1 U15394 ( .A1(n14734), .A2(n13086), .B1(n13085), .B2(n14356), .ZN(
        n13090) );
  AOI22_X1 U15395 ( .A1(n14734), .A2(n13070), .B1(n13087), .B2(n14356), .ZN(
        n13088) );
  XNOR2_X1 U15396 ( .A(n13088), .B(n10886), .ZN(n13089) );
  XOR2_X1 U15397 ( .A(n13090), .B(n13089), .Z(n13091) );
  OAI22_X1 U15398 ( .A1(n13092), .A2(n15055), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13104), .ZN(n13096) );
  INV_X1 U15399 ( .A(n14357), .ZN(n14335) );
  INV_X1 U15400 ( .A(n13093), .ZN(n13094) );
  OAI22_X1 U15401 ( .A1(n14335), .A2(n15056), .B1(n15072), .B2(n13094), .ZN(
        n13095) );
  AOI211_X1 U15402 ( .C1(n14734), .C2(n15067), .A(n13096), .B(n13095), .ZN(
        n13097) );
  AOI211_X1 U15403 ( .C1(n13101), .C2(n13100), .A(n14781), .B(n14495), .ZN(
        n14728) );
  AOI21_X1 U15404 ( .B1(n13102), .B2(P1_B_REG_SCAN_IN), .A(n14702), .ZN(n14490) );
  NAND2_X1 U15405 ( .A1(n14354), .A2(n14490), .ZN(n14724) );
  NOR2_X1 U15406 ( .A1(n13103), .A2(n14724), .ZN(n13107) );
  NOR3_X1 U15407 ( .A1(n13105), .A2(n14706), .A3(n13104), .ZN(n13106) );
  AOI211_X1 U15408 ( .C1(n15143), .C2(P1_REG2_REG_29__SCAN_IN), .A(n13107), 
        .B(n13106), .ZN(n13108) );
  OAI21_X1 U15409 ( .B1(n14726), .B2(n14709), .A(n13108), .ZN(n13109) );
  AOI21_X1 U15410 ( .B1(n14728), .B2(n14713), .A(n13109), .ZN(n13119) );
  NOR2_X1 U15411 ( .A1(n13110), .A2(n14356), .ZN(n13112) );
  INV_X1 U15412 ( .A(n14356), .ZN(n13111) );
  XNOR2_X1 U15413 ( .A(n13115), .B(n13114), .ZN(n13116) );
  NAND2_X1 U15414 ( .A1(n14356), .A2(n14620), .ZN(n14725) );
  AOI21_X1 U15415 ( .B1(n14730), .B2(n14725), .A(n15143), .ZN(n13117) );
  INV_X1 U15416 ( .A(n13117), .ZN(n13118) );
  OAI211_X1 U15417 ( .C1(n14731), .C2(n14716), .A(n13119), .B(n13118), .ZN(
        P1_U3356) );
  OAI222_X1 U15418 ( .A1(n14196), .A2(n13122), .B1(P2_U3088), .B2(n13121), 
        .C1(n13120), .C2(n14201), .ZN(P2_U3297) );
  NAND2_X1 U15419 ( .A1(n13123), .A2(n13559), .ZN(n13403) );
  OAI21_X1 U15420 ( .B1(n13541), .B2(n13124), .A(n13403), .ZN(n13127) );
  OAI21_X1 U15421 ( .B1(n13129), .B2(n13566), .A(n6765), .ZN(P3_U3204) );
  INV_X1 U15422 ( .A(n13130), .ZN(n13131) );
  OAI222_X1 U15423 ( .A1(P3_U3151), .A2(n13133), .B1(n13690), .B2(n13132), 
        .C1(n13688), .C2(n13131), .ZN(P3_U3265) );
  XNOR2_X1 U15424 ( .A(n13180), .B(n13174), .ZN(n13212) );
  XNOR2_X1 U15425 ( .A(n13212), .B(n13303), .ZN(n13213) );
  NAND2_X1 U15426 ( .A1(n13134), .A2(n13186), .ZN(n13135) );
  NAND2_X1 U15427 ( .A1(n13136), .A2(n13135), .ZN(n13185) );
  XNOR2_X1 U15428 ( .A(n14938), .B(n13215), .ZN(n13138) );
  XNOR2_X1 U15429 ( .A(n13138), .B(n13137), .ZN(n13184) );
  NAND2_X1 U15430 ( .A1(n13138), .A2(n13312), .ZN(n13139) );
  XNOR2_X1 U15431 ( .A(n14933), .B(n13215), .ZN(n13141) );
  XNOR2_X1 U15432 ( .A(n13141), .B(n13188), .ZN(n13310) );
  NAND2_X1 U15433 ( .A1(n13311), .A2(n13310), .ZN(n13309) );
  NAND2_X1 U15434 ( .A1(n13141), .A2(n13140), .ZN(n13142) );
  NAND2_X1 U15435 ( .A1(n13309), .A2(n13142), .ZN(n13246) );
  XNOR2_X1 U15436 ( .A(n13143), .B(n13215), .ZN(n13144) );
  XNOR2_X1 U15437 ( .A(n13144), .B(n13256), .ZN(n13245) );
  INV_X1 U15438 ( .A(n13144), .ZN(n13145) );
  NAND2_X1 U15439 ( .A1(n13145), .A2(n13256), .ZN(n13146) );
  XNOR2_X1 U15440 ( .A(n13670), .B(n13215), .ZN(n13147) );
  XNOR2_X1 U15441 ( .A(n13147), .B(n13294), .ZN(n13254) );
  NAND2_X1 U15442 ( .A1(n13255), .A2(n13254), .ZN(n13253) );
  NAND2_X1 U15443 ( .A1(n13147), .A2(n13532), .ZN(n13148) );
  XNOR2_X1 U15444 ( .A(n13544), .B(n13215), .ZN(n13149) );
  XNOR2_X1 U15445 ( .A(n13149), .B(n13150), .ZN(n13292) );
  INV_X1 U15446 ( .A(n13149), .ZN(n13151) );
  NAND2_X1 U15447 ( .A1(n13151), .A2(n13150), .ZN(n13152) );
  NAND2_X1 U15448 ( .A1(n13291), .A2(n13152), .ZN(n13206) );
  XNOR2_X1 U15449 ( .A(n13153), .B(n13215), .ZN(n13154) );
  XNOR2_X1 U15450 ( .A(n13154), .B(n13534), .ZN(n13205) );
  NAND2_X1 U15451 ( .A1(n13206), .A2(n13205), .ZN(n13204) );
  INV_X1 U15452 ( .A(n13154), .ZN(n13155) );
  NAND2_X1 U15453 ( .A1(n13155), .A2(n13534), .ZN(n13156) );
  XNOR2_X1 U15454 ( .A(n13274), .B(n13215), .ZN(n13157) );
  XNOR2_X1 U15455 ( .A(n13157), .B(n13493), .ZN(n13276) );
  INV_X1 U15456 ( .A(n13157), .ZN(n13158) );
  NAND2_X1 U15457 ( .A1(n13158), .A2(n13493), .ZN(n13159) );
  XNOR2_X1 U15458 ( .A(n13498), .B(n13215), .ZN(n13161) );
  XNOR2_X1 U15459 ( .A(n13161), .B(n13506), .ZN(n13229) );
  NAND2_X1 U15460 ( .A1(n13161), .A2(n13506), .ZN(n13162) );
  XNOR2_X1 U15461 ( .A(n13288), .B(n6816), .ZN(n13193) );
  XNOR2_X1 U15462 ( .A(n13272), .B(n13215), .ZN(n13266) );
  OR2_X1 U15463 ( .A1(n13266), .A2(n13265), .ZN(n13164) );
  XNOR2_X1 U15464 ( .A(n13470), .B(n13215), .ZN(n13262) );
  OR2_X1 U15465 ( .A1(n13262), .A2(n13483), .ZN(n13163) );
  NAND2_X1 U15466 ( .A1(n13164), .A2(n13163), .ZN(n13165) );
  AOI21_X1 U15467 ( .B1(n13193), .B2(n13494), .A(n13165), .ZN(n13171) );
  INV_X1 U15468 ( .A(n13266), .ZN(n13169) );
  AOI21_X1 U15469 ( .B1(n13262), .B2(n13483), .A(n13265), .ZN(n13168) );
  OR3_X1 U15470 ( .A1(n13165), .A2(n13193), .A3(n13494), .ZN(n13167) );
  NAND3_X1 U15471 ( .A1(n13262), .A2(n13483), .A3(n13265), .ZN(n13166) );
  OAI211_X1 U15472 ( .C1(n13169), .C2(n13168), .A(n13167), .B(n13166), .ZN(
        n13170) );
  XNOR2_X1 U15473 ( .A(n13240), .B(n13215), .ZN(n13172) );
  XNOR2_X1 U15474 ( .A(n13172), .B(n13268), .ZN(n13236) );
  INV_X1 U15475 ( .A(n13172), .ZN(n13173) );
  XNOR2_X1 U15476 ( .A(n13306), .B(n13174), .ZN(n13175) );
  XNOR2_X1 U15477 ( .A(n13175), .B(n13419), .ZN(n13301) );
  INV_X1 U15478 ( .A(n13175), .ZN(n13176) );
  XOR2_X1 U15479 ( .A(n13213), .B(n13214), .Z(n13182) );
  AOI22_X1 U15480 ( .A1(n13238), .A2(n13313), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13178) );
  NAND2_X1 U15481 ( .A1(n13426), .A2(n13319), .ZN(n13177) );
  OAI211_X1 U15482 ( .C1(n13420), .C2(n13315), .A(n13178), .B(n13177), .ZN(
        n13179) );
  AOI21_X1 U15483 ( .B1(n13180), .B2(n15377), .A(n13179), .ZN(n13181) );
  OAI21_X1 U15484 ( .B1(n13182), .B2(n15381), .A(n13181), .ZN(P3_U3154) );
  OAI211_X1 U15485 ( .C1(n13185), .C2(n13184), .A(n13183), .B(n15390), .ZN(
        n13192) );
  NAND2_X1 U15486 ( .A1(n13313), .A2(n13186), .ZN(n13187) );
  NAND2_X1 U15487 ( .A1(P3_REG3_REG_14__SCAN_IN), .A2(P3_U3151), .ZN(n15518)
         );
  OAI211_X1 U15488 ( .C1(n13188), .C2(n13315), .A(n13187), .B(n15518), .ZN(
        n13189) );
  AOI21_X1 U15489 ( .B1(n13319), .B2(n13190), .A(n13189), .ZN(n13191) );
  OAI211_X1 U15490 ( .C1(n15397), .C2(n14938), .A(n13192), .B(n13191), .ZN(
        P3_U3155) );
  INV_X1 U15491 ( .A(n13193), .ZN(n13194) );
  XNOR2_X1 U15492 ( .A(n13264), .B(n13483), .ZN(n13203) );
  AOI22_X1 U15493 ( .A1(n13237), .A2(n13533), .B1(n13531), .B2(n13494), .ZN(
        n13468) );
  OAI22_X1 U15494 ( .A1(n13468), .A2(n15370), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13199), .ZN(n13200) );
  AOI21_X1 U15495 ( .B1(n13319), .B2(n13475), .A(n13200), .ZN(n13202) );
  NAND2_X1 U15496 ( .A1(n13470), .A2(n15377), .ZN(n13201) );
  OAI211_X1 U15497 ( .C1(n13203), .C2(n15381), .A(n13202), .B(n13201), .ZN(
        P3_U3156) );
  OAI211_X1 U15498 ( .C1(n13206), .C2(n13205), .A(n13204), .B(n15390), .ZN(
        n13211) );
  NOR2_X1 U15499 ( .A1(n13295), .A2(n13517), .ZN(n13209) );
  OAI22_X1 U15500 ( .A1(n13315), .A2(n13519), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n13207), .ZN(n13208) );
  AOI211_X1 U15501 ( .C1(n13319), .C2(n13523), .A(n13209), .B(n13208), .ZN(
        n13210) );
  OAI211_X1 U15502 ( .C1(n13665), .C2(n15397), .A(n13211), .B(n13210), .ZN(
        P3_U3159) );
  XNOR2_X1 U15503 ( .A(n13216), .B(n13215), .ZN(n13217) );
  OAI22_X1 U15504 ( .A1(n13218), .A2(n13295), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n8253), .ZN(n13221) );
  NOR2_X1 U15505 ( .A1(n13219), .A2(n13315), .ZN(n13220) );
  AOI211_X1 U15506 ( .C1(n13319), .C2(n13408), .A(n13221), .B(n13220), .ZN(
        n13224) );
  NAND2_X1 U15507 ( .A1(n13222), .A2(n15377), .ZN(n13223) );
  OAI211_X1 U15508 ( .C1(n13225), .C2(n15381), .A(n13224), .B(n13223), .ZN(
        P3_U3160) );
  INV_X1 U15509 ( .A(n13226), .ZN(n13227) );
  AOI21_X1 U15510 ( .B1(n13229), .B2(n13228), .A(n13227), .ZN(n13234) );
  NAND2_X1 U15511 ( .A1(n13319), .A2(n13499), .ZN(n13231) );
  AOI22_X1 U15512 ( .A1(n13494), .A2(n13278), .B1(P3_REG3_REG_21__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13230) );
  OAI211_X1 U15513 ( .C1(n13519), .C2(n13295), .A(n13231), .B(n13230), .ZN(
        n13232) );
  AOI21_X1 U15514 ( .B1(n13498), .B2(n15377), .A(n13232), .ZN(n13233) );
  OAI21_X1 U15515 ( .B1(n13234), .B2(n15381), .A(n13233), .ZN(P3_U3163) );
  XOR2_X1 U15516 ( .A(n13236), .B(n13235), .Z(n13243) );
  AOI22_X1 U15517 ( .A1(n13238), .A2(n13533), .B1(n13237), .B2(n13531), .ZN(
        n13445) );
  OAI22_X1 U15518 ( .A1(n13445), .A2(n15370), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n8086), .ZN(n13239) );
  AOI21_X1 U15519 ( .B1(n13319), .B2(n13449), .A(n13239), .ZN(n13242) );
  NAND2_X1 U15520 ( .A1(n13240), .A2(n15377), .ZN(n13241) );
  OAI211_X1 U15521 ( .C1(n13243), .C2(n15381), .A(n13242), .B(n13241), .ZN(
        P3_U3165) );
  OAI211_X1 U15522 ( .C1(n13246), .C2(n13245), .A(n13244), .B(n15390), .ZN(
        n13252) );
  NOR2_X1 U15523 ( .A1(n13247), .A2(P3_STATE_REG_SCAN_IN), .ZN(n13372) );
  NOR2_X1 U15524 ( .A1(n15370), .A2(n13248), .ZN(n13249) );
  AOI211_X1 U15525 ( .C1(n13319), .C2(n13250), .A(n13372), .B(n13249), .ZN(
        n13251) );
  OAI211_X1 U15526 ( .C1(n13675), .C2(n15397), .A(n13252), .B(n13251), .ZN(
        P3_U3166) );
  OAI211_X1 U15527 ( .C1(n13255), .C2(n13254), .A(n13253), .B(n15390), .ZN(
        n13261) );
  OR2_X1 U15528 ( .A1(n13517), .A2(n13520), .ZN(n13258) );
  NAND2_X1 U15529 ( .A1(n13256), .A2(n13531), .ZN(n13257) );
  AND2_X1 U15530 ( .A1(n13258), .A2(n13257), .ZN(n13554) );
  NAND2_X1 U15531 ( .A1(P3_U3151), .A2(P3_REG3_REG_17__SCAN_IN), .ZN(n13390)
         );
  OAI21_X1 U15532 ( .B1(n15370), .B2(n13554), .A(n13390), .ZN(n13259) );
  AOI21_X1 U15533 ( .B1(n13319), .B2(n13558), .A(n13259), .ZN(n13260) );
  OAI211_X1 U15534 ( .C1(n15397), .C2(n13670), .A(n13261), .B(n13260), .ZN(
        P3_U3168) );
  XNOR2_X1 U15535 ( .A(n13266), .B(n13265), .ZN(n13267) );
  INV_X1 U15536 ( .A(n13461), .ZN(n13270) );
  OAI22_X1 U15537 ( .A1(n13268), .A2(n13520), .B1(n13483), .B2(n13518), .ZN(
        n13460) );
  AOI22_X1 U15538 ( .A1(n13460), .A2(n15393), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13269) );
  OAI21_X1 U15539 ( .B1(n13270), .B2(n15401), .A(n13269), .ZN(n13271) );
  AOI21_X1 U15540 ( .B1(n13272), .B2(n15377), .A(n13271), .ZN(n13273) );
  INV_X1 U15541 ( .A(n13274), .ZN(n13661) );
  OAI211_X1 U15542 ( .C1(n13277), .C2(n13276), .A(n13275), .B(n15390), .ZN(
        n13282) );
  AOI22_X1 U15543 ( .A1(n13284), .A2(n13278), .B1(P3_REG3_REG_20__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13279) );
  OAI21_X1 U15544 ( .B1(n13505), .B2(n13295), .A(n13279), .ZN(n13280) );
  AOI21_X1 U15545 ( .B1(n13319), .B2(n13509), .A(n13280), .ZN(n13281) );
  OAI211_X1 U15546 ( .C1(n13661), .C2(n15397), .A(n13282), .B(n13281), .ZN(
        P3_U3173) );
  XNOR2_X1 U15547 ( .A(n13283), .B(n13494), .ZN(n13290) );
  NAND2_X1 U15548 ( .A1(n13319), .A2(n13486), .ZN(n13286) );
  AOI22_X1 U15549 ( .A1(n13284), .A2(n13313), .B1(P3_REG3_REG_22__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13285) );
  OAI211_X1 U15550 ( .C1(n13483), .C2(n13315), .A(n13286), .B(n13285), .ZN(
        n13287) );
  AOI21_X1 U15551 ( .B1(n13288), .B2(n15377), .A(n13287), .ZN(n13289) );
  OAI21_X1 U15552 ( .B1(n13290), .B2(n15381), .A(n13289), .ZN(P3_U3175) );
  INV_X1 U15553 ( .A(n13544), .ZN(n13612) );
  OAI211_X1 U15554 ( .C1(n13293), .C2(n13292), .A(n13291), .B(n15390), .ZN(
        n13299) );
  NOR2_X1 U15555 ( .A1(n13295), .A2(n13294), .ZN(n13297) );
  OAI22_X1 U15556 ( .A1(n13315), .A2(n13505), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n14932), .ZN(n13296) );
  AOI211_X1 U15557 ( .C1(n13319), .C2(n13537), .A(n13297), .B(n13296), .ZN(
        n13298) );
  OAI211_X1 U15558 ( .C1(n13612), .C2(n15397), .A(n13299), .B(n13298), .ZN(
        P3_U3178) );
  XOR2_X1 U15559 ( .A(n13301), .B(n13300), .Z(n13308) );
  AOI22_X1 U15560 ( .A1(n13303), .A2(n13533), .B1(n13531), .B2(n13302), .ZN(
        n13433) );
  AOI22_X1 U15561 ( .A1(n13437), .A2(n13319), .B1(P3_REG3_REG_26__SCAN_IN), 
        .B2(P3_U3151), .ZN(n13304) );
  OAI21_X1 U15562 ( .B1(n13433), .B2(n15370), .A(n13304), .ZN(n13305) );
  AOI21_X1 U15563 ( .B1(n13306), .B2(n15377), .A(n13305), .ZN(n13307) );
  OAI21_X1 U15564 ( .B1(n13308), .B2(n15381), .A(n13307), .ZN(P3_U3180) );
  OAI211_X1 U15565 ( .C1(n13311), .C2(n13310), .A(n13309), .B(n15390), .ZN(
        n13321) );
  NAND2_X1 U15566 ( .A1(n13313), .A2(n13312), .ZN(n13314) );
  NAND2_X1 U15567 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(P3_U3151), .ZN(n13353)
         );
  OAI211_X1 U15568 ( .C1(n13316), .C2(n13315), .A(n13314), .B(n13353), .ZN(
        n13317) );
  AOI21_X1 U15569 ( .B1(n13319), .B2(n13318), .A(n13317), .ZN(n13320) );
  OAI211_X1 U15570 ( .C1(n15397), .C2(n14933), .A(n13321), .B(n13320), .ZN(
        P3_U3181) );
  MUX2_X1 U15571 ( .A(n13322), .B(P3_DATAO_REG_23__SCAN_IN), .S(n13329), .Z(
        P3_U3514) );
  MUX2_X1 U15572 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n13493), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U15573 ( .A(n13534), .B(P3_DATAO_REG_19__SCAN_IN), .S(n13329), .Z(
        P3_U3510) );
  MUX2_X1 U15574 ( .A(P3_DATAO_REG_12__SCAN_IN), .B(n13323), .S(P3_U3897), .Z(
        P3_U3503) );
  MUX2_X1 U15575 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n13324), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U15576 ( .A(n13325), .B(P3_DATAO_REG_9__SCAN_IN), .S(n13329), .Z(
        P3_U3500) );
  MUX2_X1 U15577 ( .A(P3_DATAO_REG_6__SCAN_IN), .B(n13326), .S(P3_U3897), .Z(
        P3_U3497) );
  MUX2_X1 U15578 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n13327), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U15579 ( .A(P3_DATAO_REG_1__SCAN_IN), .B(n13328), .S(P3_U3897), .Z(
        P3_U3492) );
  MUX2_X1 U15580 ( .A(n13330), .B(P3_DATAO_REG_0__SCAN_IN), .S(n13329), .Z(
        P3_U3491) );
  AOI21_X1 U15581 ( .B1(n13333), .B2(n13332), .A(n13331), .ZN(n13346) );
  AOI21_X1 U15582 ( .B1(n13336), .B2(n13335), .A(n13334), .ZN(n13339) );
  NAND2_X1 U15583 ( .A1(n15523), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n13338) );
  OAI211_X1 U15584 ( .C1(n13339), .C2(n7858), .A(n13338), .B(n13337), .ZN(
        n13344) );
  AOI21_X1 U15585 ( .B1(n14947), .B2(n13341), .A(n13340), .ZN(n13342) );
  NOR2_X1 U15586 ( .A1(n13342), .A2(n15516), .ZN(n13343) );
  AOI211_X1 U15587 ( .C1(n15485), .C2(n6870), .A(n13344), .B(n13343), .ZN(
        n13345) );
  OAI21_X1 U15588 ( .B1(n13346), .B2(n15530), .A(n13345), .ZN(P3_U3195) );
  AOI21_X1 U15589 ( .B1(n14937), .B2(n13348), .A(n13347), .ZN(n13364) );
  AOI21_X1 U15590 ( .B1(n13351), .B2(n13350), .A(n13349), .ZN(n13352) );
  OR2_X1 U15591 ( .A1(n13352), .A2(n15530), .ZN(n13363) );
  NAND2_X1 U15592 ( .A1(n15523), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n13354) );
  NAND2_X1 U15593 ( .A1(n13354), .A2(n13353), .ZN(n13360) );
  AOI21_X1 U15594 ( .B1(n13357), .B2(n13356), .A(n13355), .ZN(n13358) );
  NOR2_X1 U15595 ( .A1(n13358), .A2(n7858), .ZN(n13359) );
  AOI211_X1 U15596 ( .C1(n15485), .C2(n13361), .A(n13360), .B(n13359), .ZN(
        n13362) );
  OAI211_X1 U15597 ( .C1(n13364), .C2(n15516), .A(n13363), .B(n13362), .ZN(
        P3_U3197) );
  AOI21_X1 U15598 ( .B1(n13367), .B2(n13366), .A(n13365), .ZN(n13382) );
  NOR2_X1 U15599 ( .A1(n13369), .A2(n13368), .ZN(n13371) );
  XOR2_X1 U15600 ( .A(n13371), .B(n13370), .Z(n13380) );
  AOI21_X1 U15601 ( .B1(n15523), .B2(P3_ADDR_REG_16__SCAN_IN), .A(n13372), 
        .ZN(n13373) );
  OAI21_X1 U15602 ( .B1(n15520), .B2(n13374), .A(n13373), .ZN(n13379) );
  AOI21_X1 U15603 ( .B1(n6719), .B2(n13376), .A(n13375), .ZN(n13377) );
  NOR2_X1 U15604 ( .A1(n13377), .A2(n15516), .ZN(n13378) );
  AOI211_X1 U15605 ( .C1(n15504), .C2(n13380), .A(n13379), .B(n13378), .ZN(
        n13381) );
  OAI21_X1 U15606 ( .B1(n13382), .B2(n15530), .A(n13381), .ZN(P3_U3198) );
  AOI21_X1 U15607 ( .B1(n13617), .B2(n13384), .A(n13383), .ZN(n13400) );
  INV_X1 U15608 ( .A(n13385), .ZN(n13386) );
  NOR2_X1 U15609 ( .A1(n13386), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n13389) );
  OAI21_X1 U15610 ( .B1(n13389), .B2(n13388), .A(n13387), .ZN(n13399) );
  INV_X1 U15611 ( .A(P3_ADDR_REG_17__SCAN_IN), .ZN(n13391) );
  OAI21_X1 U15612 ( .B1(n15492), .B2(n13391), .A(n13390), .ZN(n13396) );
  AOI211_X1 U15613 ( .C1(n13394), .C2(n13393), .A(n7858), .B(n13392), .ZN(
        n13395) );
  AOI211_X1 U15614 ( .C1(n15485), .C2(n13397), .A(n13396), .B(n13395), .ZN(
        n13398) );
  OAI211_X1 U15615 ( .C1(n13400), .C2(n15516), .A(n13399), .B(n13398), .ZN(
        P3_U3199) );
  AOI21_X1 U15616 ( .B1(n13403), .B2(n13624), .A(n13560), .ZN(n13405) );
  AOI21_X1 U15617 ( .B1(n13560), .B2(P3_REG2_REG_31__SCAN_IN), .A(n13405), 
        .ZN(n13404) );
  OAI21_X1 U15618 ( .B1(n13626), .B2(n13562), .A(n13404), .ZN(P3_U3202) );
  AOI21_X1 U15619 ( .B1(n13560), .B2(P3_REG2_REG_30__SCAN_IN), .A(n13405), 
        .ZN(n13406) );
  OAI21_X1 U15620 ( .B1(n13629), .B2(n13562), .A(n13406), .ZN(P3_U3203) );
  INV_X1 U15621 ( .A(n13407), .ZN(n13414) );
  AOI22_X1 U15622 ( .A1(n13408), .A2(n13559), .B1(P3_REG2_REG_28__SCAN_IN), 
        .B2(n13566), .ZN(n13409) );
  OAI21_X1 U15623 ( .B1(n13410), .B2(n13562), .A(n13409), .ZN(n13411) );
  AOI21_X1 U15624 ( .B1(n13412), .B2(n13564), .A(n13411), .ZN(n13413) );
  OAI21_X1 U15625 ( .B1(n13414), .B2(n13566), .A(n13413), .ZN(P3_U3205) );
  AOI21_X1 U15626 ( .B1(n13417), .B2(n13416), .A(n13415), .ZN(n13418) );
  OAI222_X1 U15627 ( .A1(n13520), .A2(n13420), .B1(n13518), .B2(n13419), .C1(
        n13418), .C2(n13515), .ZN(n13571) );
  INV_X1 U15628 ( .A(n13571), .ZN(n13430) );
  INV_X1 U15629 ( .A(n9039), .ZN(n13425) );
  NAND3_X1 U15630 ( .A1(n13423), .A2(n13422), .A3(n13421), .ZN(n13424) );
  NAND2_X1 U15631 ( .A1(n13425), .A2(n13424), .ZN(n13572) );
  AOI22_X1 U15632 ( .A1(n13426), .A2(n13559), .B1(P3_REG2_REG_27__SCAN_IN), 
        .B2(n13566), .ZN(n13427) );
  OAI21_X1 U15633 ( .B1(n13633), .B2(n13562), .A(n13427), .ZN(n13428) );
  AOI21_X1 U15634 ( .B1(n13572), .B2(n13564), .A(n13428), .ZN(n13429) );
  OAI21_X1 U15635 ( .B1(n13430), .B2(n13560), .A(n13429), .ZN(P3_U3206) );
  XNOR2_X1 U15636 ( .A(n13432), .B(n13431), .ZN(n13434) );
  OAI21_X1 U15637 ( .B1(n13434), .B2(n13515), .A(n13433), .ZN(n13575) );
  INV_X1 U15638 ( .A(n13575), .ZN(n13441) );
  XNOR2_X1 U15639 ( .A(n13436), .B(n13435), .ZN(n13576) );
  AOI22_X1 U15640 ( .A1(n13437), .A2(n13559), .B1(P3_REG2_REG_26__SCAN_IN), 
        .B2(n13566), .ZN(n13438) );
  OAI21_X1 U15641 ( .B1(n13637), .B2(n13562), .A(n13438), .ZN(n13439) );
  AOI21_X1 U15642 ( .B1(n13576), .B2(n13564), .A(n13439), .ZN(n13440) );
  OAI21_X1 U15643 ( .B1(n13441), .B2(n13566), .A(n13440), .ZN(P3_U3207) );
  OR3_X1 U15644 ( .A1(n6705), .A2(n13442), .A3(n13447), .ZN(n13443) );
  NAND3_X1 U15645 ( .A1(n13444), .A2(n13552), .A3(n13443), .ZN(n13446) );
  NAND2_X1 U15646 ( .A1(n13446), .A2(n13445), .ZN(n13579) );
  INV_X1 U15647 ( .A(n13579), .ZN(n13453) );
  XNOR2_X1 U15648 ( .A(n13448), .B(n13447), .ZN(n13580) );
  AOI22_X1 U15649 ( .A1(n13449), .A2(n13559), .B1(P3_REG2_REG_25__SCAN_IN), 
        .B2(n13566), .ZN(n13450) );
  OAI21_X1 U15650 ( .B1(n13641), .B2(n13562), .A(n13450), .ZN(n13451) );
  AOI21_X1 U15651 ( .B1(n13580), .B2(n13564), .A(n13451), .ZN(n13452) );
  OAI21_X1 U15652 ( .B1(n13453), .B2(n13566), .A(n13452), .ZN(P3_U3208) );
  OAI21_X1 U15653 ( .B1(n13474), .B2(n13455), .A(n13454), .ZN(n13456) );
  NAND2_X1 U15654 ( .A1(n7471), .A2(n13456), .ZN(n13585) );
  AOI211_X1 U15655 ( .C1(n13458), .C2(n13457), .A(n13515), .B(n6705), .ZN(
        n13459) );
  AOI211_X1 U15656 ( .C1(n15588), .C2(n13585), .A(n13460), .B(n13459), .ZN(
        n13583) );
  AOI22_X1 U15657 ( .A1(n13461), .A2(n13559), .B1(n13560), .B2(
        P3_REG2_REG_24__SCAN_IN), .ZN(n13462) );
  OAI21_X1 U15658 ( .B1(n13645), .B2(n13562), .A(n13462), .ZN(n13463) );
  AOI21_X1 U15659 ( .B1(n13585), .B2(n13464), .A(n13463), .ZN(n13465) );
  OAI21_X1 U15660 ( .B1(n13583), .B2(n13566), .A(n13465), .ZN(P3_U3209) );
  XNOR2_X1 U15661 ( .A(n13467), .B(n13466), .ZN(n13469) );
  OAI21_X1 U15662 ( .B1(n13469), .B2(n13515), .A(n13468), .ZN(n13588) );
  INV_X1 U15663 ( .A(n13470), .ZN(n13649) );
  NOR2_X1 U15664 ( .A1(n13472), .A2(n13471), .ZN(n13473) );
  NOR2_X1 U15665 ( .A1(n13474), .A2(n13473), .ZN(n13589) );
  NAND2_X1 U15666 ( .A1(n13589), .A2(n13564), .ZN(n13477) );
  AOI22_X1 U15667 ( .A1(n13560), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n13559), 
        .B2(n13475), .ZN(n13476) );
  OAI211_X1 U15668 ( .C1(n13649), .C2(n13562), .A(n13477), .B(n13476), .ZN(
        n13478) );
  AOI21_X1 U15669 ( .B1(n13588), .B2(n13541), .A(n13478), .ZN(n13479) );
  INV_X1 U15670 ( .A(n13479), .ZN(P3_U3210) );
  XNOR2_X1 U15671 ( .A(n13481), .B(n13480), .ZN(n13482) );
  OAI222_X1 U15672 ( .A1(n13520), .A2(n13483), .B1(n13518), .B2(n13506), .C1(
        n13515), .C2(n13482), .ZN(n13592) );
  INV_X1 U15673 ( .A(n13592), .ZN(n13490) );
  XNOR2_X1 U15674 ( .A(n13485), .B(n13484), .ZN(n13593) );
  AOI22_X1 U15675 ( .A1(n13560), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n13559), 
        .B2(n13486), .ZN(n13487) );
  OAI21_X1 U15676 ( .B1(n13653), .B2(n13562), .A(n13487), .ZN(n13488) );
  AOI21_X1 U15677 ( .B1(n13593), .B2(n13564), .A(n13488), .ZN(n13489) );
  OAI21_X1 U15678 ( .B1(n13490), .B2(n13566), .A(n13489), .ZN(P3_U3211) );
  OAI21_X1 U15679 ( .B1(n13492), .B2(n13496), .A(n13491), .ZN(n13495) );
  AOI222_X1 U15680 ( .A1(n13552), .A2(n13495), .B1(n13494), .B2(n13533), .C1(
        n13493), .C2(n13531), .ZN(n13596) );
  XNOR2_X1 U15681 ( .A(n13497), .B(n13496), .ZN(n13598) );
  INV_X1 U15682 ( .A(n13498), .ZN(n13657) );
  AOI22_X1 U15683 ( .A1(n13560), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n13559), 
        .B2(n13499), .ZN(n13500) );
  OAI21_X1 U15684 ( .B1(n13657), .B2(n13562), .A(n13500), .ZN(n13501) );
  AOI21_X1 U15685 ( .B1(n13598), .B2(n13564), .A(n13501), .ZN(n13502) );
  OAI21_X1 U15686 ( .B1(n13596), .B2(n13566), .A(n13502), .ZN(P3_U3212) );
  XNOR2_X1 U15687 ( .A(n13503), .B(n13508), .ZN(n13504) );
  OAI222_X1 U15688 ( .A1(n13520), .A2(n13506), .B1(n13518), .B2(n13505), .C1(
        n13504), .C2(n13515), .ZN(n13601) );
  INV_X1 U15689 ( .A(n13601), .ZN(n13513) );
  XOR2_X1 U15690 ( .A(n13508), .B(n13507), .Z(n13602) );
  AOI22_X1 U15691 ( .A1(n13560), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n13559), 
        .B2(n13509), .ZN(n13510) );
  OAI21_X1 U15692 ( .B1(n13661), .B2(n13562), .A(n13510), .ZN(n13511) );
  AOI21_X1 U15693 ( .B1(n13602), .B2(n13564), .A(n13511), .ZN(n13512) );
  OAI21_X1 U15694 ( .B1(n13513), .B2(n13566), .A(n13512), .ZN(P3_U3213) );
  XOR2_X1 U15695 ( .A(n13521), .B(n13514), .Z(n13516) );
  OAI222_X1 U15696 ( .A1(n13520), .A2(n13519), .B1(n13518), .B2(n13517), .C1(
        n13516), .C2(n13515), .ZN(n13605) );
  INV_X1 U15697 ( .A(n13605), .ZN(n13527) );
  XNOR2_X1 U15698 ( .A(n13522), .B(n13521), .ZN(n13606) );
  AOI22_X1 U15699 ( .A1(n13560), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n13559), 
        .B2(n13523), .ZN(n13524) );
  OAI21_X1 U15700 ( .B1(n13665), .B2(n13562), .A(n13524), .ZN(n13525) );
  AOI21_X1 U15701 ( .B1(n13606), .B2(n13564), .A(n13525), .ZN(n13526) );
  OAI21_X1 U15702 ( .B1(n13527), .B2(n13566), .A(n13526), .ZN(P3_U3214) );
  XNOR2_X1 U15703 ( .A(n13529), .B(n13528), .ZN(n13530) );
  NAND2_X1 U15704 ( .A1(n13530), .A2(n13552), .ZN(n13536) );
  AOI22_X1 U15705 ( .A1(n13534), .A2(n13533), .B1(n13532), .B2(n13531), .ZN(
        n13535) );
  NAND2_X1 U15706 ( .A1(n13536), .A2(n13535), .ZN(n13614) );
  INV_X1 U15707 ( .A(n13614), .ZN(n13550) );
  INV_X1 U15708 ( .A(n13537), .ZN(n13539) );
  OAI22_X1 U15709 ( .A1(n13541), .A2(n13540), .B1(n13539), .B2(n13538), .ZN(
        n13542) );
  AOI21_X1 U15710 ( .B1(n13544), .B2(n13543), .A(n13542), .ZN(n13549) );
  NAND2_X1 U15711 ( .A1(n13547), .A2(n13546), .ZN(n13609) );
  NAND3_X1 U15712 ( .A1(n13610), .A2(n13609), .A3(n13564), .ZN(n13548) );
  OAI211_X1 U15713 ( .C1(n13550), .C2(n13560), .A(n13549), .B(n13548), .ZN(
        P3_U3215) );
  OAI211_X1 U15714 ( .C1(n13553), .C2(n8978), .A(n13552), .B(n13551), .ZN(
        n13555) );
  NAND2_X1 U15715 ( .A1(n13555), .A2(n13554), .ZN(n13615) );
  INV_X1 U15716 ( .A(n13615), .ZN(n13567) );
  XNOR2_X1 U15717 ( .A(n13557), .B(n13556), .ZN(n13616) );
  AOI22_X1 U15718 ( .A1(n13560), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n13559), 
        .B2(n13558), .ZN(n13561) );
  OAI21_X1 U15719 ( .B1(n13670), .B2(n13562), .A(n13561), .ZN(n13563) );
  AOI21_X1 U15720 ( .B1(n13616), .B2(n13564), .A(n13563), .ZN(n13565) );
  OAI21_X1 U15721 ( .B1(n13567), .B2(n13566), .A(n13565), .ZN(P3_U3216) );
  NOR2_X1 U15722 ( .A1(n13624), .A2(n9022), .ZN(n13569) );
  AOI21_X1 U15723 ( .B1(P3_REG1_REG_31__SCAN_IN), .B2(n9022), .A(n13569), .ZN(
        n13568) );
  OAI21_X1 U15724 ( .B1(n13626), .B2(n13623), .A(n13568), .ZN(P3_U3490) );
  AOI21_X1 U15725 ( .B1(P3_REG1_REG_30__SCAN_IN), .B2(n9022), .A(n13569), .ZN(
        n13570) );
  OAI21_X1 U15726 ( .B1(n13629), .B2(n13623), .A(n13570), .ZN(P3_U3489) );
  INV_X1 U15727 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n13573) );
  AOI21_X1 U15728 ( .B1(n14957), .B2(n13572), .A(n13571), .ZN(n13630) );
  OAI21_X1 U15729 ( .B1(n13633), .B2(n13623), .A(n13574), .ZN(P3_U3486) );
  INV_X1 U15730 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n13577) );
  AOI21_X1 U15731 ( .B1(n13576), .B2(n14957), .A(n13575), .ZN(n13634) );
  MUX2_X1 U15732 ( .A(n13577), .B(n13634), .S(n15607), .Z(n13578) );
  OAI21_X1 U15733 ( .B1(n13637), .B2(n13623), .A(n13578), .ZN(P3_U3485) );
  INV_X1 U15734 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n13581) );
  AOI21_X1 U15735 ( .B1(n13580), .B2(n14957), .A(n13579), .ZN(n13638) );
  MUX2_X1 U15736 ( .A(n13581), .B(n13638), .S(n15607), .Z(n13582) );
  OAI21_X1 U15737 ( .B1(n13641), .B2(n13623), .A(n13582), .ZN(P3_U3484) );
  INV_X1 U15738 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n13586) );
  INV_X1 U15739 ( .A(n15583), .ZN(n15578) );
  INV_X1 U15740 ( .A(n13583), .ZN(n13584) );
  AOI21_X1 U15741 ( .B1(n15578), .B2(n13585), .A(n13584), .ZN(n13642) );
  MUX2_X1 U15742 ( .A(n13586), .B(n13642), .S(n15607), .Z(n13587) );
  OAI21_X1 U15743 ( .B1(n13645), .B2(n13623), .A(n13587), .ZN(P3_U3483) );
  INV_X1 U15744 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n13590) );
  AOI21_X1 U15745 ( .B1(n13589), .B2(n14957), .A(n13588), .ZN(n13646) );
  MUX2_X1 U15746 ( .A(n13590), .B(n13646), .S(n15607), .Z(n13591) );
  OAI21_X1 U15747 ( .B1(n13649), .B2(n13623), .A(n13591), .ZN(P3_U3482) );
  INV_X1 U15748 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n13594) );
  AOI21_X1 U15749 ( .B1(n14957), .B2(n13593), .A(n13592), .ZN(n13650) );
  MUX2_X1 U15750 ( .A(n13594), .B(n13650), .S(n15607), .Z(n13595) );
  OAI21_X1 U15751 ( .B1(n13653), .B2(n13623), .A(n13595), .ZN(P3_U3481) );
  INV_X1 U15752 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n13599) );
  INV_X1 U15753 ( .A(n13596), .ZN(n13597) );
  AOI21_X1 U15754 ( .B1(n14957), .B2(n13598), .A(n13597), .ZN(n13654) );
  MUX2_X1 U15755 ( .A(n13599), .B(n13654), .S(n15607), .Z(n13600) );
  OAI21_X1 U15756 ( .B1(n13657), .B2(n13623), .A(n13600), .ZN(P3_U3480) );
  INV_X1 U15757 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n13603) );
  AOI21_X1 U15758 ( .B1(n13602), .B2(n14957), .A(n13601), .ZN(n13658) );
  MUX2_X1 U15759 ( .A(n13603), .B(n13658), .S(n15607), .Z(n13604) );
  OAI21_X1 U15760 ( .B1(n13661), .B2(n13623), .A(n13604), .ZN(P3_U3479) );
  AOI21_X1 U15761 ( .B1(n13606), .B2(n14957), .A(n13605), .ZN(n13662) );
  MUX2_X1 U15762 ( .A(n13607), .B(n13662), .S(n15607), .Z(n13608) );
  OAI21_X1 U15763 ( .B1(n13665), .B2(n13623), .A(n13608), .ZN(P3_U3478) );
  NAND3_X1 U15764 ( .A1(n13610), .A2(n13609), .A3(n14957), .ZN(n13611) );
  OAI21_X1 U15765 ( .B1(n13612), .B2(n15582), .A(n13611), .ZN(n13613) );
  MUX2_X1 U15766 ( .A(P3_REG1_REG_18__SCAN_IN), .B(n13666), .S(n15607), .Z(
        P3_U3477) );
  AOI21_X1 U15767 ( .B1(n13616), .B2(n14957), .A(n13615), .ZN(n13667) );
  MUX2_X1 U15768 ( .A(n13617), .B(n13667), .S(n15607), .Z(n13618) );
  OAI21_X1 U15769 ( .B1(n13623), .B2(n13670), .A(n13618), .ZN(P3_U3476) );
  AOI21_X1 U15770 ( .B1(n14957), .B2(n13620), .A(n13619), .ZN(n13671) );
  MUX2_X1 U15771 ( .A(n13621), .B(n13671), .S(n15607), .Z(n13622) );
  OAI21_X1 U15772 ( .B1(n13675), .B2(n13623), .A(n13622), .ZN(P3_U3475) );
  NOR2_X1 U15773 ( .A1(n13624), .A2(n15589), .ZN(n13627) );
  AOI21_X1 U15774 ( .B1(P3_REG0_REG_31__SCAN_IN), .B2(n15589), .A(n13627), 
        .ZN(n13625) );
  OAI21_X1 U15775 ( .B1(n13626), .B2(n13674), .A(n13625), .ZN(P3_U3458) );
  AOI21_X1 U15776 ( .B1(P3_REG0_REG_30__SCAN_IN), .B2(n15589), .A(n13627), 
        .ZN(n13628) );
  OAI21_X1 U15777 ( .B1(n13629), .B2(n13674), .A(n13628), .ZN(P3_U3457) );
  INV_X1 U15778 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n13631) );
  OAI21_X1 U15779 ( .B1(n13633), .B2(n13674), .A(n13632), .ZN(P3_U3454) );
  INV_X1 U15780 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n13635) );
  MUX2_X1 U15781 ( .A(n13635), .B(n13634), .S(n15591), .Z(n13636) );
  OAI21_X1 U15782 ( .B1(n13637), .B2(n13674), .A(n13636), .ZN(P3_U3453) );
  INV_X1 U15783 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n13639) );
  MUX2_X1 U15784 ( .A(n13639), .B(n13638), .S(n15591), .Z(n13640) );
  OAI21_X1 U15785 ( .B1(n13641), .B2(n13674), .A(n13640), .ZN(P3_U3452) );
  INV_X1 U15786 ( .A(P3_REG0_REG_24__SCAN_IN), .ZN(n13643) );
  MUX2_X1 U15787 ( .A(n13643), .B(n13642), .S(n15591), .Z(n13644) );
  OAI21_X1 U15788 ( .B1(n13645), .B2(n13674), .A(n13644), .ZN(P3_U3451) );
  INV_X1 U15789 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n13647) );
  MUX2_X1 U15790 ( .A(n13647), .B(n13646), .S(n15591), .Z(n13648) );
  OAI21_X1 U15791 ( .B1(n13649), .B2(n13674), .A(n13648), .ZN(P3_U3450) );
  INV_X1 U15792 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n13651) );
  MUX2_X1 U15793 ( .A(n13651), .B(n13650), .S(n15591), .Z(n13652) );
  OAI21_X1 U15794 ( .B1(n13653), .B2(n13674), .A(n13652), .ZN(P3_U3449) );
  INV_X1 U15795 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n13655) );
  MUX2_X1 U15796 ( .A(n13655), .B(n13654), .S(n15591), .Z(n13656) );
  OAI21_X1 U15797 ( .B1(n13657), .B2(n13674), .A(n13656), .ZN(P3_U3448) );
  INV_X1 U15798 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n13659) );
  MUX2_X1 U15799 ( .A(n13659), .B(n13658), .S(n15591), .Z(n13660) );
  OAI21_X1 U15800 ( .B1(n13661), .B2(n13674), .A(n13660), .ZN(P3_U3447) );
  INV_X1 U15801 ( .A(P3_REG0_REG_19__SCAN_IN), .ZN(n13663) );
  MUX2_X1 U15802 ( .A(n13663), .B(n13662), .S(n15591), .Z(n13664) );
  OAI21_X1 U15803 ( .B1(n13665), .B2(n13674), .A(n13664), .ZN(P3_U3446) );
  MUX2_X1 U15804 ( .A(P3_REG0_REG_18__SCAN_IN), .B(n13666), .S(n15591), .Z(
        P3_U3444) );
  INV_X1 U15805 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n13668) );
  MUX2_X1 U15806 ( .A(n13668), .B(n13667), .S(n15591), .Z(n13669) );
  OAI21_X1 U15807 ( .B1(n13674), .B2(n13670), .A(n13669), .ZN(P3_U3441) );
  INV_X1 U15808 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n13672) );
  MUX2_X1 U15809 ( .A(n13672), .B(n13671), .S(n15591), .Z(n13673) );
  OAI21_X1 U15810 ( .B1(n13675), .B2(n13674), .A(n13673), .ZN(P3_U3438) );
  NAND3_X1 U15811 ( .A1(n13676), .A2(P3_IR_REG_31__SCAN_IN), .A3(
        P3_STATE_REG_SCAN_IN), .ZN(n13678) );
  OAI22_X1 U15812 ( .A1(n13679), .A2(n13678), .B1(n13677), .B2(n13690), .ZN(
        n13680) );
  AOI21_X1 U15813 ( .B1(n13682), .B2(n13681), .A(n13680), .ZN(n13683) );
  INV_X1 U15814 ( .A(n13683), .ZN(P3_U3264) );
  INV_X1 U15815 ( .A(n13684), .ZN(n13687) );
  OAI222_X1 U15816 ( .A1(n13690), .A2(n13689), .B1(n13688), .B2(n13687), .C1(
        P3_U3151), .C2(n13685), .ZN(P3_U3266) );
  MUX2_X1 U15817 ( .A(n13691), .B(P3_IR_REG_0__SCAN_IN), .S(
        P3_STATE_REG_SCAN_IN), .Z(P3_U3295) );
  AND2_X1 U15818 ( .A1(n13875), .A2(n13735), .ZN(n13696) );
  XNOR2_X1 U15819 ( .A(n14975), .B(n13734), .ZN(n13695) );
  NOR2_X1 U15820 ( .A1(n13695), .A2(n13696), .ZN(n13697) );
  AOI21_X1 U15821 ( .B1(n13696), .B2(n13695), .A(n13697), .ZN(n13796) );
  NAND2_X1 U15822 ( .A1(n13795), .A2(n13796), .ZN(n13794) );
  INV_X1 U15823 ( .A(n13697), .ZN(n13698) );
  NAND2_X1 U15824 ( .A1(n13794), .A2(n13698), .ZN(n13803) );
  AND2_X1 U15825 ( .A1(n13874), .A2(n13735), .ZN(n13701) );
  XNOR2_X1 U15826 ( .A(n13699), .B(n13729), .ZN(n13700) );
  NOR2_X1 U15827 ( .A1(n13700), .A2(n13701), .ZN(n13702) );
  AOI21_X1 U15828 ( .B1(n13701), .B2(n13700), .A(n13702), .ZN(n13804) );
  INV_X1 U15829 ( .A(n13702), .ZN(n13703) );
  NAND2_X1 U15830 ( .A1(n13873), .A2(n13735), .ZN(n13705) );
  XNOR2_X1 U15831 ( .A(n14161), .B(n13729), .ZN(n13704) );
  XOR2_X1 U15832 ( .A(n13705), .B(n13704), .Z(n13837) );
  XNOR2_X1 U15833 ( .A(n14072), .B(n13734), .ZN(n13707) );
  NAND2_X1 U15834 ( .A1(n13872), .A2(n13735), .ZN(n13706) );
  NAND2_X1 U15835 ( .A1(n13707), .A2(n13706), .ZN(n13708) );
  OAI21_X1 U15836 ( .B1(n13707), .B2(n13706), .A(n13708), .ZN(n13756) );
  INV_X1 U15837 ( .A(n13708), .ZN(n13709) );
  XNOR2_X1 U15838 ( .A(n14052), .B(n13729), .ZN(n13711) );
  INV_X1 U15839 ( .A(n13759), .ZN(n13871) );
  NAND2_X1 U15840 ( .A1(n13871), .A2(n13735), .ZN(n13710) );
  NAND2_X1 U15841 ( .A1(n13711), .A2(n13710), .ZN(n13712) );
  OAI21_X1 U15842 ( .B1(n13711), .B2(n13710), .A(n13712), .ZN(n13821) );
  INV_X1 U15843 ( .A(n13712), .ZN(n13713) );
  XNOR2_X1 U15844 ( .A(n14146), .B(n13734), .ZN(n13716) );
  NAND2_X1 U15845 ( .A1(n13870), .A2(n13735), .ZN(n13714) );
  XNOR2_X1 U15846 ( .A(n13716), .B(n13714), .ZN(n13779) );
  INV_X1 U15847 ( .A(n13714), .ZN(n13715) );
  AND2_X1 U15848 ( .A1(n13716), .A2(n13715), .ZN(n13717) );
  AOI21_X1 U15849 ( .B1(n13780), .B2(n13779), .A(n13717), .ZN(n13718) );
  XNOR2_X1 U15850 ( .A(n14029), .B(n13729), .ZN(n13719) );
  XNOR2_X1 U15851 ( .A(n13718), .B(n13719), .ZN(n13829) );
  NAND2_X1 U15852 ( .A1(n13869), .A2(n13735), .ZN(n13828) );
  INV_X1 U15853 ( .A(n13718), .ZN(n13720) );
  XNOR2_X1 U15854 ( .A(n14008), .B(n13729), .ZN(n13721) );
  INV_X1 U15855 ( .A(n13832), .ZN(n13868) );
  NAND2_X1 U15856 ( .A1(n13868), .A2(n13735), .ZN(n13743) );
  OAI21_X2 U15857 ( .B1(n13742), .B2(n13743), .A(n13723), .ZN(n13814) );
  XNOR2_X1 U15858 ( .A(n13990), .B(n13734), .ZN(n13724) );
  NOR2_X1 U15859 ( .A1(n13788), .A2(n10697), .ZN(n13726) );
  XNOR2_X1 U15860 ( .A(n13724), .B(n13726), .ZN(n13813) );
  INV_X1 U15861 ( .A(n13724), .ZN(n13725) );
  XNOR2_X1 U15862 ( .A(n13975), .B(n13734), .ZN(n13728) );
  NAND2_X1 U15863 ( .A1(n13866), .A2(n13735), .ZN(n13727) );
  XNOR2_X1 U15864 ( .A(n13728), .B(n13727), .ZN(n13786) );
  XNOR2_X1 U15865 ( .A(n13957), .B(n13729), .ZN(n13731) );
  NAND2_X1 U15866 ( .A1(n13865), .A2(n13735), .ZN(n13730) );
  NAND2_X1 U15867 ( .A1(n13731), .A2(n13730), .ZN(n13732) );
  OAI21_X1 U15868 ( .B1(n13731), .B2(n13730), .A(n13732), .ZN(n13849) );
  INV_X1 U15869 ( .A(n13732), .ZN(n13733) );
  XNOR2_X1 U15870 ( .A(n14116), .B(n13734), .ZN(n13766) );
  NAND2_X1 U15871 ( .A1(n13864), .A2(n13735), .ZN(n13764) );
  XNOR2_X1 U15872 ( .A(n13766), .B(n13764), .ZN(n13767) );
  XNOR2_X1 U15873 ( .A(n13768), .B(n13767), .ZN(n13741) );
  NOR2_X1 U15874 ( .A1(n13789), .A2(n13839), .ZN(n13736) );
  AOI21_X1 U15875 ( .B1(n13863), .B2(n13852), .A(n13736), .ZN(n13946) );
  INV_X1 U15876 ( .A(n13737), .ZN(n13941) );
  AOI22_X1 U15877 ( .A1(n13941), .A2(n13853), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13738) );
  OAI21_X1 U15878 ( .B1(n13946), .B2(n13855), .A(n13738), .ZN(n13739) );
  AOI21_X1 U15879 ( .B1(n14116), .B2(n13857), .A(n13739), .ZN(n13740) );
  OAI21_X1 U15880 ( .B1(n13741), .B2(n13859), .A(n13740), .ZN(P2_U3186) );
  XNOR2_X1 U15881 ( .A(n13742), .B(n13743), .ZN(n13747) );
  OAI22_X1 U15882 ( .A1(n13788), .A2(n13841), .B1(n7273), .B2(n13839), .ZN(
        n14001) );
  AOI22_X1 U15883 ( .A1(n14001), .A2(n13843), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13744) );
  OAI21_X1 U15884 ( .B1(n14003), .B2(n13845), .A(n13744), .ZN(n13745) );
  AOI21_X1 U15885 ( .B1(n14136), .B2(n13857), .A(n13745), .ZN(n13746) );
  OAI21_X1 U15886 ( .B1(n13747), .B2(n13859), .A(n13746), .ZN(P2_U3188) );
  MUX2_X1 U15887 ( .A(n13845), .B(P2_STATE_REG_SCAN_IN), .S(
        P2_REG3_REG_3__SCAN_IN), .Z(n13755) );
  AOI22_X1 U15888 ( .A1(n13843), .A2(n13748), .B1(n13857), .B2(n15314), .ZN(
        n13754) );
  AOI21_X1 U15889 ( .B1(n13750), .B2(n13749), .A(n13859), .ZN(n13752) );
  NAND2_X1 U15890 ( .A1(n13752), .A2(n13751), .ZN(n13753) );
  NAND3_X1 U15891 ( .A1(n13755), .A2(n13754), .A3(n13753), .ZN(P2_U3190) );
  AOI21_X1 U15892 ( .B1(n13757), .B2(n13756), .A(n6781), .ZN(n13763) );
  NAND2_X1 U15893 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13908)
         );
  OAI22_X1 U15894 ( .A1(n13759), .A2(n13841), .B1(n13758), .B2(n13839), .ZN(
        n14064) );
  NAND2_X1 U15895 ( .A1(n13843), .A2(n14064), .ZN(n13760) );
  OAI211_X1 U15896 ( .C1(n13845), .C2(n14069), .A(n13908), .B(n13760), .ZN(
        n13761) );
  AOI21_X1 U15897 ( .B1(n14156), .B2(n13857), .A(n13761), .ZN(n13762) );
  OAI21_X1 U15898 ( .B1(n13763), .B2(n13859), .A(n13762), .ZN(P2_U3191) );
  INV_X1 U15899 ( .A(n13764), .ZN(n13765) );
  NOR2_X1 U15900 ( .A1(n13769), .A2(n10697), .ZN(n13770) );
  XNOR2_X1 U15901 ( .A(n13770), .B(n13734), .ZN(n13771) );
  XNOR2_X1 U15902 ( .A(n14110), .B(n13771), .ZN(n13772) );
  OR2_X1 U15903 ( .A1(n13773), .A2(n13841), .ZN(n13775) );
  NAND2_X1 U15904 ( .A1(n13864), .A2(n13851), .ZN(n13774) );
  AND2_X1 U15905 ( .A1(n13775), .A2(n13774), .ZN(n13930) );
  AOI22_X1 U15906 ( .A1(n13934), .A2(n13853), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13776) );
  OAI21_X1 U15907 ( .B1(n13930), .B2(n13855), .A(n13776), .ZN(n13777) );
  AOI21_X1 U15908 ( .B1(n14110), .B2(n13857), .A(n13777), .ZN(n13778) );
  XNOR2_X1 U15909 ( .A(n13780), .B(n13779), .ZN(n13785) );
  AOI22_X1 U15910 ( .A1(n13851), .A2(n13871), .B1(n13869), .B2(n13852), .ZN(
        n14033) );
  OAI22_X1 U15911 ( .A1(n14033), .A2(n13855), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13781), .ZN(n13782) );
  AOI21_X1 U15912 ( .B1(n14038), .B2(n13853), .A(n13782), .ZN(n13784) );
  NAND2_X1 U15913 ( .A1(n14146), .A2(n13857), .ZN(n13783) );
  OAI211_X1 U15914 ( .C1(n13785), .C2(n13859), .A(n13784), .B(n13783), .ZN(
        P2_U3195) );
  XNOR2_X1 U15915 ( .A(n13787), .B(n13786), .ZN(n13793) );
  OAI22_X1 U15916 ( .A1(n13789), .A2(n13841), .B1(n13788), .B2(n13839), .ZN(
        n13967) );
  AOI22_X1 U15917 ( .A1(n13967), .A2(n13843), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13790) );
  OAI21_X1 U15918 ( .B1(n13973), .B2(n13845), .A(n13790), .ZN(n13791) );
  AOI21_X1 U15919 ( .B1(n14126), .B2(n13857), .A(n13791), .ZN(n13792) );
  OAI21_X1 U15920 ( .B1(n13793), .B2(n13859), .A(n13792), .ZN(P2_U3197) );
  INV_X1 U15921 ( .A(n14975), .ZN(n15002) );
  OAI21_X1 U15922 ( .B1(n13796), .B2(n13795), .A(n13794), .ZN(n13797) );
  NAND2_X1 U15923 ( .A1(n13797), .A2(n6908), .ZN(n13801) );
  AOI22_X1 U15924 ( .A1(n13851), .A2(n13876), .B1(n13874), .B2(n13852), .ZN(
        n14971) );
  OAI21_X1 U15925 ( .B1(n13855), .B2(n14971), .A(n13798), .ZN(n13799) );
  AOI21_X1 U15926 ( .B1(n14974), .B2(n13853), .A(n13799), .ZN(n13800) );
  OAI211_X1 U15927 ( .C1(n15002), .C2(n13812), .A(n13801), .B(n13800), .ZN(
        P2_U3198) );
  OAI21_X1 U15928 ( .B1(n13804), .B2(n13803), .A(n13802), .ZN(n13805) );
  NAND2_X1 U15929 ( .A1(n13805), .A2(n6908), .ZN(n13811) );
  OAI21_X1 U15930 ( .B1(n13855), .B2(n13807), .A(n13806), .ZN(n13808) );
  AOI21_X1 U15931 ( .B1(n13809), .B2(n13853), .A(n13808), .ZN(n13810) );
  OAI211_X1 U15932 ( .C1(n14167), .C2(n13812), .A(n13811), .B(n13810), .ZN(
        P2_U3200) );
  XNOR2_X1 U15933 ( .A(n13814), .B(n13813), .ZN(n13819) );
  AOI22_X1 U15934 ( .A1(n13866), .A2(n13852), .B1(n13851), .B2(n13868), .ZN(
        n13983) );
  OAI22_X1 U15935 ( .A1(n13983), .A2(n13855), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13815), .ZN(n13816) );
  AOI21_X1 U15936 ( .B1(n13988), .B2(n13853), .A(n13816), .ZN(n13818) );
  NAND2_X1 U15937 ( .A1(n14131), .A2(n13857), .ZN(n13817) );
  OAI211_X1 U15938 ( .C1(n13819), .C2(n13859), .A(n13818), .B(n13817), .ZN(
        P2_U3201) );
  AOI21_X1 U15939 ( .B1(n13822), .B2(n13821), .A(n13820), .ZN(n13826) );
  OAI22_X1 U15940 ( .A1(n13831), .A2(n13841), .B1(n13842), .B2(n13839), .ZN(
        n14058) );
  AOI22_X1 U15941 ( .A1(n14058), .A2(n13843), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13823) );
  OAI21_X1 U15942 ( .B1(n14049), .B2(n13845), .A(n13823), .ZN(n13824) );
  AOI21_X1 U15943 ( .B1(n14151), .B2(n13857), .A(n13824), .ZN(n13825) );
  OAI21_X1 U15944 ( .B1(n13826), .B2(n13859), .A(n13825), .ZN(P2_U3205) );
  OAI21_X1 U15945 ( .B1(n13829), .B2(n13828), .A(n13827), .ZN(n13830) );
  INV_X1 U15946 ( .A(n13830), .ZN(n13836) );
  OAI22_X1 U15947 ( .A1(n13832), .A2(n13841), .B1(n13831), .B2(n13839), .ZN(
        n14018) );
  AOI22_X1 U15948 ( .A1(n14018), .A2(n13843), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13833) );
  OAI21_X1 U15949 ( .B1(n14021), .B2(n13845), .A(n13833), .ZN(n13834) );
  AOI21_X1 U15950 ( .B1(n14029), .B2(n13857), .A(n13834), .ZN(n13835) );
  OAI21_X1 U15951 ( .B1(n13836), .B2(n13859), .A(n13835), .ZN(P2_U3207) );
  XNOR2_X1 U15952 ( .A(n13838), .B(n13837), .ZN(n13848) );
  OAI22_X1 U15953 ( .A1(n13842), .A2(n13841), .B1(n13840), .B2(n13839), .ZN(
        n14084) );
  AOI22_X1 U15954 ( .A1(n13843), .A2(n14084), .B1(P2_REG3_REG_18__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13844) );
  OAI21_X1 U15955 ( .B1(n14087), .B2(n13845), .A(n13844), .ZN(n13846) );
  AOI21_X1 U15956 ( .B1(n14161), .B2(n13857), .A(n13846), .ZN(n13847) );
  OAI21_X1 U15957 ( .B1(n13848), .B2(n13859), .A(n13847), .ZN(P2_U3210) );
  AOI21_X1 U15958 ( .B1(n13850), .B2(n13849), .A(n6728), .ZN(n13860) );
  AOI22_X1 U15959 ( .A1(n13864), .A2(n13852), .B1(n13851), .B2(n13866), .ZN(
        n13961) );
  AOI22_X1 U15960 ( .A1(n13955), .A2(n13853), .B1(P2_REG3_REG_26__SCAN_IN), 
        .B2(P2_U3088), .ZN(n13854) );
  OAI21_X1 U15961 ( .B1(n13961), .B2(n13855), .A(n13854), .ZN(n13856) );
  AOI21_X1 U15962 ( .B1(n14122), .B2(n13857), .A(n13856), .ZN(n13858) );
  OAI21_X1 U15963 ( .B1(n13860), .B2(n13859), .A(n13858), .ZN(P2_U3212) );
  INV_X2 U15964 ( .A(P2_U3947), .ZN(n13883) );
  MUX2_X1 U15965 ( .A(n13912), .B(P2_DATAO_REG_31__SCAN_IN), .S(n13883), .Z(
        P2_U3562) );
  MUX2_X1 U15966 ( .A(n13861), .B(P2_DATAO_REG_30__SCAN_IN), .S(n13883), .Z(
        P2_U3561) );
  MUX2_X1 U15967 ( .A(n13862), .B(P2_DATAO_REG_29__SCAN_IN), .S(n13883), .Z(
        P2_U3560) );
  MUX2_X1 U15968 ( .A(n13863), .B(P2_DATAO_REG_28__SCAN_IN), .S(n13883), .Z(
        P2_U3559) );
  MUX2_X1 U15969 ( .A(n13864), .B(P2_DATAO_REG_27__SCAN_IN), .S(n13883), .Z(
        P2_U3558) );
  MUX2_X1 U15970 ( .A(n13865), .B(P2_DATAO_REG_26__SCAN_IN), .S(n13883), .Z(
        P2_U3557) );
  MUX2_X1 U15971 ( .A(n13866), .B(P2_DATAO_REG_25__SCAN_IN), .S(n13883), .Z(
        P2_U3556) );
  MUX2_X1 U15972 ( .A(n13867), .B(P2_DATAO_REG_24__SCAN_IN), .S(n13883), .Z(
        P2_U3555) );
  MUX2_X1 U15973 ( .A(n13868), .B(P2_DATAO_REG_23__SCAN_IN), .S(n13883), .Z(
        P2_U3554) );
  MUX2_X1 U15974 ( .A(n13869), .B(P2_DATAO_REG_22__SCAN_IN), .S(n13883), .Z(
        P2_U3553) );
  MUX2_X1 U15975 ( .A(n13870), .B(P2_DATAO_REG_21__SCAN_IN), .S(n13883), .Z(
        P2_U3552) );
  MUX2_X1 U15976 ( .A(n13871), .B(P2_DATAO_REG_20__SCAN_IN), .S(n13883), .Z(
        P2_U3551) );
  MUX2_X1 U15977 ( .A(n13872), .B(P2_DATAO_REG_19__SCAN_IN), .S(n13883), .Z(
        P2_U3550) );
  MUX2_X1 U15978 ( .A(n13873), .B(P2_DATAO_REG_18__SCAN_IN), .S(n13883), .Z(
        P2_U3549) );
  MUX2_X1 U15979 ( .A(n13874), .B(P2_DATAO_REG_17__SCAN_IN), .S(n13883), .Z(
        P2_U3548) );
  MUX2_X1 U15980 ( .A(n13875), .B(P2_DATAO_REG_16__SCAN_IN), .S(n13883), .Z(
        P2_U3547) );
  MUX2_X1 U15981 ( .A(n13876), .B(P2_DATAO_REG_15__SCAN_IN), .S(n13883), .Z(
        P2_U3546) );
  MUX2_X1 U15982 ( .A(n13877), .B(P2_DATAO_REG_14__SCAN_IN), .S(n13883), .Z(
        P2_U3545) );
  MUX2_X1 U15983 ( .A(n13878), .B(P2_DATAO_REG_13__SCAN_IN), .S(n13883), .Z(
        P2_U3544) );
  MUX2_X1 U15984 ( .A(n13879), .B(P2_DATAO_REG_12__SCAN_IN), .S(n13883), .Z(
        P2_U3543) );
  MUX2_X1 U15985 ( .A(n13880), .B(P2_DATAO_REG_11__SCAN_IN), .S(n13883), .Z(
        P2_U3542) );
  MUX2_X1 U15986 ( .A(n13881), .B(P2_DATAO_REG_10__SCAN_IN), .S(n13883), .Z(
        P2_U3541) );
  MUX2_X1 U15987 ( .A(n13882), .B(P2_DATAO_REG_9__SCAN_IN), .S(n13883), .Z(
        P2_U3540) );
  MUX2_X1 U15988 ( .A(n13884), .B(P2_DATAO_REG_8__SCAN_IN), .S(n13883), .Z(
        P2_U3539) );
  MUX2_X1 U15989 ( .A(n13885), .B(P2_DATAO_REG_7__SCAN_IN), .S(n13883), .Z(
        P2_U3538) );
  MUX2_X1 U15990 ( .A(n13886), .B(P2_DATAO_REG_6__SCAN_IN), .S(n13883), .Z(
        P2_U3537) );
  MUX2_X1 U15991 ( .A(n13887), .B(P2_DATAO_REG_5__SCAN_IN), .S(n13883), .Z(
        P2_U3536) );
  MUX2_X1 U15992 ( .A(n13888), .B(P2_DATAO_REG_4__SCAN_IN), .S(n13883), .Z(
        P2_U3535) );
  MUX2_X1 U15993 ( .A(n13889), .B(P2_DATAO_REG_3__SCAN_IN), .S(n13883), .Z(
        P2_U3534) );
  MUX2_X1 U15994 ( .A(n13890), .B(P2_DATAO_REG_2__SCAN_IN), .S(n13883), .Z(
        P2_U3533) );
  MUX2_X1 U15995 ( .A(n13891), .B(P2_DATAO_REG_1__SCAN_IN), .S(n13883), .Z(
        P2_U3532) );
  MUX2_X1 U15996 ( .A(n9763), .B(P2_DATAO_REG_0__SCAN_IN), .S(n13883), .Z(
        P2_U3531) );
  NOR2_X1 U15997 ( .A1(n13897), .A2(n13892), .ZN(n13893) );
  NOR2_X1 U15998 ( .A1(n13894), .A2(n13893), .ZN(n13895) );
  XOR2_X1 U15999 ( .A(n13895), .B(P2_REG2_REG_19__SCAN_IN), .Z(n13905) );
  INV_X1 U16000 ( .A(n13905), .ZN(n13903) );
  NAND2_X1 U16001 ( .A1(n13897), .A2(n13896), .ZN(n13898) );
  NAND2_X1 U16002 ( .A1(n13899), .A2(n13898), .ZN(n13900) );
  XOR2_X1 U16003 ( .A(n13900), .B(P2_REG1_REG_19__SCAN_IN), .Z(n13904) );
  OAI21_X1 U16004 ( .B1(n13904), .B2(n13901), .A(n15225), .ZN(n13902) );
  AOI21_X1 U16005 ( .B1(n13903), .B2(n15252), .A(n13902), .ZN(n13907) );
  AOI22_X1 U16006 ( .A1(n13905), .A2(n15252), .B1(n15255), .B2(n13904), .ZN(
        n13906) );
  MUX2_X1 U16007 ( .A(n13907), .B(n13906), .S(n9758), .Z(n13909) );
  OAI211_X1 U16008 ( .C1(n8356), .C2(n15228), .A(n13909), .B(n13908), .ZN(
        P2_U3233) );
  XNOR2_X1 U16009 ( .A(n13917), .B(n14101), .ZN(n13911) );
  NAND2_X1 U16010 ( .A1(n13911), .A2(n15274), .ZN(n14100) );
  NAND2_X1 U16011 ( .A1(n15269), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n13914) );
  NAND2_X1 U16012 ( .A1(n13913), .A2(n13912), .ZN(n14102) );
  OR2_X1 U16013 ( .A1(n14078), .A2(n14102), .ZN(n13919) );
  OAI211_X1 U16014 ( .C1(n14101), .C2(n14094), .A(n13914), .B(n13919), .ZN(
        n13915) );
  INV_X1 U16015 ( .A(n13915), .ZN(n13916) );
  OAI21_X1 U16016 ( .B1(n14100), .B2(n14026), .A(n13916), .ZN(P2_U3234) );
  OAI211_X1 U16017 ( .C1(n13918), .C2(n14104), .A(n15274), .B(n13917), .ZN(
        n14103) );
  INV_X1 U16018 ( .A(n13919), .ZN(n13921) );
  NOR2_X1 U16019 ( .A1(n14104), .A2(n14094), .ZN(n13920) );
  AOI211_X1 U16020 ( .C1(n14078), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13921), 
        .B(n13920), .ZN(n13922) );
  OAI21_X1 U16021 ( .B1(n14026), .B2(n14103), .A(n13922), .ZN(P2_U3235) );
  XNOR2_X1 U16022 ( .A(n13924), .B(n13923), .ZN(n14114) );
  AOI22_X1 U16023 ( .A1(n14110), .A2(n15270), .B1(n15269), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n13938) );
  AND2_X1 U16024 ( .A1(n13925), .A2(n13926), .ZN(n13929) );
  OAI211_X1 U16025 ( .C1(n13929), .C2(n13928), .A(n13927), .B(n14065), .ZN(
        n13931) );
  INV_X1 U16026 ( .A(n13932), .ZN(n13933) );
  AOI21_X1 U16027 ( .B1(n14110), .B2(n13940), .A(n13933), .ZN(n14111) );
  AOI22_X1 U16028 ( .A1(n14111), .A2(n10697), .B1(n13934), .B2(n15268), .ZN(
        n13935) );
  AOI21_X1 U16029 ( .B1(n14113), .B2(n13935), .A(n15269), .ZN(n13936) );
  INV_X1 U16030 ( .A(n13936), .ZN(n13937) );
  OAI211_X1 U16031 ( .C1(n14114), .C2(n14099), .A(n13938), .B(n13937), .ZN(
        P2_U3237) );
  XNOR2_X1 U16032 ( .A(n13939), .B(n13944), .ZN(n14119) );
  AOI211_X1 U16033 ( .C1(n14116), .C2(n13954), .A(n14091), .B(n7058), .ZN(
        n14115) );
  AOI22_X1 U16034 ( .A1(n13941), .A2(n15268), .B1(P2_REG2_REG_27__SCAN_IN), 
        .B2(n15269), .ZN(n13942) );
  OAI21_X1 U16035 ( .B1(n13943), .B2(n14094), .A(n13942), .ZN(n13950) );
  OAI21_X1 U16036 ( .B1(n13945), .B2(n13944), .A(n13925), .ZN(n13948) );
  INV_X1 U16037 ( .A(n13946), .ZN(n13947) );
  AOI21_X1 U16038 ( .B1(n13948), .B2(n14065), .A(n13947), .ZN(n14118) );
  NOR2_X1 U16039 ( .A1(n14118), .A2(n15269), .ZN(n13949) );
  AOI211_X1 U16040 ( .C1(n14115), .C2(n15279), .A(n13950), .B(n13949), .ZN(
        n13951) );
  OAI21_X1 U16041 ( .B1(n14099), .B2(n14119), .A(n13951), .ZN(P2_U3238) );
  XOR2_X1 U16042 ( .A(n13959), .B(n13952), .Z(n14124) );
  OR2_X1 U16043 ( .A1(n13976), .A2(n13957), .ZN(n13953) );
  AND3_X1 U16044 ( .A1(n13954), .A2(n13953), .A3(n15274), .ZN(n14121) );
  AOI22_X1 U16045 ( .A1(n13955), .A2(n15268), .B1(P2_REG2_REG_26__SCAN_IN), 
        .B2(n15269), .ZN(n13956) );
  OAI21_X1 U16046 ( .B1(n13957), .B2(n14094), .A(n13956), .ZN(n13958) );
  AOI21_X1 U16047 ( .B1(n14121), .B2(n15279), .A(n13958), .ZN(n13965) );
  XNOR2_X1 U16048 ( .A(n13960), .B(n13959), .ZN(n13963) );
  OAI21_X1 U16049 ( .B1(n13963), .B2(n13962), .A(n13961), .ZN(n14120) );
  NAND2_X1 U16050 ( .A1(n14120), .A2(n14088), .ZN(n13964) );
  OAI211_X1 U16051 ( .C1(n14124), .C2(n14099), .A(n13965), .B(n13964), .ZN(
        P2_U3239) );
  XNOR2_X1 U16052 ( .A(n13966), .B(n13971), .ZN(n13968) );
  AOI21_X1 U16053 ( .B1(n13968), .B2(n14065), .A(n13967), .ZN(n14128) );
  AOI21_X1 U16054 ( .B1(n13971), .B2(n13970), .A(n13969), .ZN(n14129) );
  INV_X1 U16055 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n13972) );
  OAI22_X1 U16056 ( .A1(n13973), .A2(n14086), .B1(n14088), .B2(n13972), .ZN(
        n13974) );
  AOI21_X1 U16057 ( .B1(n14126), .B2(n15270), .A(n13974), .ZN(n13979) );
  OAI21_X1 U16058 ( .B1(n13975), .B2(n13986), .A(n15274), .ZN(n13977) );
  NOR2_X1 U16059 ( .A1(n13977), .A2(n13976), .ZN(n14125) );
  NAND2_X1 U16060 ( .A1(n14125), .A2(n15279), .ZN(n13978) );
  OAI211_X1 U16061 ( .C1(n14129), .C2(n14099), .A(n13979), .B(n13978), .ZN(
        n13980) );
  INV_X1 U16062 ( .A(n13980), .ZN(n13981) );
  OAI21_X1 U16063 ( .B1(n14078), .B2(n14128), .A(n13981), .ZN(P2_U3240) );
  XNOR2_X1 U16064 ( .A(n13982), .B(n13992), .ZN(n13985) );
  INV_X1 U16065 ( .A(n13983), .ZN(n13984) );
  AOI21_X1 U16066 ( .B1(n13985), .B2(n14065), .A(n13984), .ZN(n14133) );
  OAI21_X1 U16067 ( .B1(n13990), .B2(n14005), .A(n15274), .ZN(n13987) );
  NOR2_X1 U16068 ( .A1(n13987), .A2(n13986), .ZN(n14130) );
  AOI22_X1 U16069 ( .A1(n13988), .A2(n15268), .B1(n15269), .B2(
        P2_REG2_REG_24__SCAN_IN), .ZN(n13989) );
  OAI21_X1 U16070 ( .B1(n13990), .B2(n14094), .A(n13989), .ZN(n13994) );
  OAI21_X1 U16071 ( .B1(n6764), .B2(n13992), .A(n13991), .ZN(n14134) );
  NOR2_X1 U16072 ( .A1(n14134), .A2(n14099), .ZN(n13993) );
  AOI211_X1 U16073 ( .C1(n14130), .C2(n15279), .A(n13994), .B(n13993), .ZN(
        n13995) );
  OAI21_X1 U16074 ( .B1(n14078), .B2(n14133), .A(n13995), .ZN(P2_U3241) );
  AOI21_X1 U16075 ( .B1(n14000), .B2(n13997), .A(n13996), .ZN(n14139) );
  OAI21_X1 U16076 ( .B1(n14000), .B2(n13999), .A(n13998), .ZN(n14002) );
  AOI21_X1 U16077 ( .B1(n14002), .B2(n14065), .A(n14001), .ZN(n14138) );
  OAI21_X1 U16078 ( .B1(n14003), .B2(n14086), .A(n14138), .ZN(n14004) );
  NAND2_X1 U16079 ( .A1(n14004), .A2(n14088), .ZN(n14011) );
  INV_X1 U16080 ( .A(n14025), .ZN(n14006) );
  AOI211_X1 U16081 ( .C1(n14136), .C2(n14006), .A(n14091), .B(n14005), .ZN(
        n14135) );
  INV_X1 U16082 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n14007) );
  OAI22_X1 U16083 ( .A1(n14008), .A2(n14094), .B1(n14088), .B2(n14007), .ZN(
        n14009) );
  AOI21_X1 U16084 ( .B1(n14135), .B2(n15279), .A(n14009), .ZN(n14010) );
  OAI211_X1 U16085 ( .C1(n14099), .C2(n14139), .A(n14011), .B(n14010), .ZN(
        P2_U3242) );
  NAND2_X1 U16086 ( .A1(n14012), .A2(n14015), .ZN(n14013) );
  NAND2_X1 U16087 ( .A1(n14014), .A2(n14013), .ZN(n14140) );
  XNOR2_X1 U16088 ( .A(n14016), .B(n9751), .ZN(n14017) );
  NAND2_X1 U16089 ( .A1(n14017), .A2(n14065), .ZN(n14020) );
  INV_X1 U16090 ( .A(n14018), .ZN(n14019) );
  NAND2_X1 U16091 ( .A1(n14020), .A2(n14019), .ZN(n14143) );
  NAND2_X1 U16092 ( .A1(n14143), .A2(n14088), .ZN(n14031) );
  INV_X1 U16093 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n14022) );
  OAI22_X1 U16094 ( .A1(n14088), .A2(n14022), .B1(n14021), .B2(n14086), .ZN(
        n14028) );
  NAND2_X1 U16095 ( .A1(n14036), .A2(n14029), .ZN(n14023) );
  NAND2_X1 U16096 ( .A1(n14023), .A2(n15274), .ZN(n14024) );
  OR2_X1 U16097 ( .A1(n14025), .A2(n14024), .ZN(n14141) );
  NOR2_X1 U16098 ( .A1(n14141), .A2(n14026), .ZN(n14027) );
  AOI211_X1 U16099 ( .C1(n15270), .C2(n14029), .A(n14028), .B(n14027), .ZN(
        n14030) );
  OAI211_X1 U16100 ( .C1(n14099), .C2(n14140), .A(n14031), .B(n14030), .ZN(
        P2_U3243) );
  XNOR2_X1 U16101 ( .A(n14032), .B(n14041), .ZN(n14035) );
  INV_X1 U16102 ( .A(n14033), .ZN(n14034) );
  AOI21_X1 U16103 ( .B1(n14035), .B2(n14065), .A(n14034), .ZN(n14147) );
  INV_X1 U16104 ( .A(n14036), .ZN(n14037) );
  AOI211_X1 U16105 ( .C1(n14146), .C2(n14048), .A(n14091), .B(n14037), .ZN(
        n14145) );
  AOI22_X1 U16106 ( .A1(n15269), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n14038), 
        .B2(n15268), .ZN(n14039) );
  OAI21_X1 U16107 ( .B1(n14040), .B2(n14094), .A(n14039), .ZN(n14044) );
  XNOR2_X1 U16108 ( .A(n14042), .B(n14041), .ZN(n14149) );
  NOR2_X1 U16109 ( .A1(n14149), .A2(n14099), .ZN(n14043) );
  AOI211_X1 U16110 ( .C1(n14145), .C2(n15279), .A(n14044), .B(n14043), .ZN(
        n14045) );
  OAI21_X1 U16111 ( .B1(n14078), .B2(n14147), .A(n14045), .ZN(P2_U3244) );
  XNOR2_X1 U16112 ( .A(n14046), .B(n14054), .ZN(n14154) );
  OR2_X1 U16113 ( .A1(n14067), .A2(n14052), .ZN(n14047) );
  AND3_X1 U16114 ( .A1(n14048), .A2(n14047), .A3(n15274), .ZN(n14150) );
  NOR2_X1 U16115 ( .A1(n14049), .A2(n14086), .ZN(n14050) );
  AOI21_X1 U16116 ( .B1(n14078), .B2(P2_REG2_REG_20__SCAN_IN), .A(n14050), 
        .ZN(n14051) );
  OAI21_X1 U16117 ( .B1(n14052), .B2(n14094), .A(n14051), .ZN(n14061) );
  INV_X1 U16118 ( .A(n14053), .ZN(n14057) );
  INV_X1 U16119 ( .A(n14054), .ZN(n14056) );
  OAI21_X1 U16120 ( .B1(n14057), .B2(n14056), .A(n14055), .ZN(n14059) );
  AOI21_X1 U16121 ( .B1(n14059), .B2(n14065), .A(n14058), .ZN(n14153) );
  NOR2_X1 U16122 ( .A1(n14153), .A2(n15269), .ZN(n14060) );
  AOI211_X1 U16123 ( .C1(n14150), .C2(n15279), .A(n14061), .B(n14060), .ZN(
        n14062) );
  OAI21_X1 U16124 ( .B1(n14099), .B2(n14154), .A(n14062), .ZN(P2_U3245) );
  XOR2_X1 U16125 ( .A(n14063), .B(n14073), .Z(n14066) );
  AOI21_X1 U16126 ( .B1(n14066), .B2(n14065), .A(n14064), .ZN(n14158) );
  INV_X1 U16127 ( .A(n14090), .ZN(n14068) );
  AOI211_X1 U16128 ( .C1(n14156), .C2(n14068), .A(n14091), .B(n14067), .ZN(
        n14155) );
  INV_X1 U16129 ( .A(n14069), .ZN(n14070) );
  AOI22_X1 U16130 ( .A1(n15269), .A2(P2_REG2_REG_19__SCAN_IN), .B1(n14070), 
        .B2(n15268), .ZN(n14071) );
  OAI21_X1 U16131 ( .B1(n14072), .B2(n14094), .A(n14071), .ZN(n14076) );
  XNOR2_X1 U16132 ( .A(n14074), .B(n14073), .ZN(n14159) );
  NOR2_X1 U16133 ( .A1(n14159), .A2(n14099), .ZN(n14075) );
  AOI211_X1 U16134 ( .C1(n14155), .C2(n15279), .A(n14076), .B(n14075), .ZN(
        n14077) );
  OAI21_X1 U16135 ( .B1(n14078), .B2(n14158), .A(n14077), .ZN(P2_U3246) );
  INV_X1 U16136 ( .A(n14079), .ZN(n14080) );
  AOI21_X1 U16137 ( .B1(n14082), .B2(n14081), .A(n14080), .ZN(n14164) );
  XNOR2_X1 U16138 ( .A(n14083), .B(n14082), .ZN(n14085) );
  AOI21_X1 U16139 ( .B1(n14085), .B2(n14065), .A(n14084), .ZN(n14163) );
  OAI21_X1 U16140 ( .B1(n14087), .B2(n14086), .A(n14163), .ZN(n14089) );
  NAND2_X1 U16141 ( .A1(n14089), .A2(n14088), .ZN(n14098) );
  AOI211_X1 U16142 ( .C1(n14161), .C2(n14092), .A(n14091), .B(n14090), .ZN(
        n14160) );
  INV_X1 U16143 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n14093) );
  OAI22_X1 U16144 ( .A1(n14095), .A2(n14094), .B1(n14088), .B2(n14093), .ZN(
        n14096) );
  AOI21_X1 U16145 ( .B1(n14160), .B2(n15279), .A(n14096), .ZN(n14097) );
  OAI211_X1 U16146 ( .C1(n14099), .C2(n14164), .A(n14098), .B(n14097), .ZN(
        P2_U3247) );
  OAI211_X1 U16147 ( .C1(n14101), .C2(n15340), .A(n14100), .B(n14102), .ZN(
        n14171) );
  MUX2_X1 U16148 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n14171), .S(n15357), .Z(
        P2_U3530) );
  OAI211_X1 U16149 ( .C1(n14104), .C2(n15340), .A(n14103), .B(n14102), .ZN(
        n14172) );
  MUX2_X1 U16150 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n14172), .S(n15357), .Z(
        P2_U3529) );
  AOI21_X1 U16151 ( .B1(n15313), .B2(n14106), .A(n14105), .ZN(n14107) );
  AOI22_X1 U16152 ( .A1(n14111), .A2(n15274), .B1(n15313), .B2(n14110), .ZN(
        n14112) );
  OAI211_X1 U16153 ( .C1(n14114), .C2(n15000), .A(n14113), .B(n14112), .ZN(
        n14174) );
  MUX2_X1 U16154 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n14174), .S(n15357), .Z(
        P2_U3527) );
  AOI21_X1 U16155 ( .B1(n15313), .B2(n14116), .A(n14115), .ZN(n14117) );
  OAI211_X1 U16156 ( .C1(n14119), .C2(n15000), .A(n14118), .B(n14117), .ZN(
        n14175) );
  MUX2_X1 U16157 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n14175), .S(n15357), .Z(
        P2_U3526) );
  AOI211_X1 U16158 ( .C1(n15313), .C2(n14122), .A(n14121), .B(n14120), .ZN(
        n14123) );
  OAI21_X1 U16159 ( .B1(n14124), .B2(n15000), .A(n14123), .ZN(n14176) );
  MUX2_X1 U16160 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n14176), .S(n15357), .Z(
        P2_U3525) );
  AOI21_X1 U16161 ( .B1(n15313), .B2(n14126), .A(n14125), .ZN(n14127) );
  OAI211_X1 U16162 ( .C1(n14129), .C2(n15000), .A(n14128), .B(n14127), .ZN(
        n14177) );
  MUX2_X1 U16163 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n14177), .S(n15357), .Z(
        P2_U3524) );
  AOI21_X1 U16164 ( .B1(n15313), .B2(n14131), .A(n14130), .ZN(n14132) );
  OAI211_X1 U16165 ( .C1(n14134), .C2(n15000), .A(n14133), .B(n14132), .ZN(
        n14178) );
  MUX2_X1 U16166 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n14178), .S(n15357), .Z(
        P2_U3523) );
  AOI21_X1 U16167 ( .B1(n15313), .B2(n14136), .A(n14135), .ZN(n14137) );
  OAI211_X1 U16168 ( .C1(n14139), .C2(n15000), .A(n14138), .B(n14137), .ZN(
        n14179) );
  MUX2_X1 U16169 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n14179), .S(n15357), .Z(
        P2_U3522) );
  NOR2_X1 U16170 ( .A1(n14140), .A2(n15000), .ZN(n14144) );
  OAI21_X1 U16171 ( .B1(n7056), .B2(n15340), .A(n14141), .ZN(n14142) );
  MUX2_X1 U16172 ( .A(n14180), .B(P2_REG1_REG_22__SCAN_IN), .S(n15355), .Z(
        P2_U3521) );
  AOI21_X1 U16173 ( .B1(n15313), .B2(n14146), .A(n14145), .ZN(n14148) );
  OAI211_X1 U16174 ( .C1(n15000), .C2(n14149), .A(n14148), .B(n14147), .ZN(
        n14181) );
  MUX2_X1 U16175 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n14181), .S(n15357), .Z(
        P2_U3520) );
  AOI21_X1 U16176 ( .B1(n15313), .B2(n14151), .A(n14150), .ZN(n14152) );
  OAI211_X1 U16177 ( .C1(n15000), .C2(n14154), .A(n14153), .B(n14152), .ZN(
        n14182) );
  MUX2_X1 U16178 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n14182), .S(n15357), .Z(
        P2_U3519) );
  AOI21_X1 U16179 ( .B1(n15313), .B2(n14156), .A(n14155), .ZN(n14157) );
  OAI211_X1 U16180 ( .C1(n15000), .C2(n14159), .A(n14158), .B(n14157), .ZN(
        n14183) );
  MUX2_X1 U16181 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n14183), .S(n15357), .Z(
        P2_U3518) );
  AOI21_X1 U16182 ( .B1(n15313), .B2(n14161), .A(n14160), .ZN(n14162) );
  OAI211_X1 U16183 ( .C1(n14164), .C2(n15000), .A(n14163), .B(n14162), .ZN(
        n14184) );
  MUX2_X1 U16184 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n14184), .S(n15357), .Z(
        P2_U3517) );
  NOR2_X1 U16185 ( .A1(n14165), .A2(n15000), .ZN(n14170) );
  OAI21_X1 U16186 ( .B1(n14167), .B2(n15340), .A(n14166), .ZN(n14168) );
  MUX2_X1 U16187 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n14185), .S(n15357), .Z(
        P2_U3516) );
  MUX2_X1 U16188 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n14171), .S(n15347), .Z(
        P2_U3498) );
  MUX2_X1 U16189 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n14172), .S(n15347), .Z(
        P2_U3497) );
  MUX2_X1 U16190 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n14174), .S(n15347), .Z(
        P2_U3495) );
  MUX2_X1 U16191 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n14175), .S(n15347), .Z(
        P2_U3494) );
  MUX2_X1 U16192 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n14176), .S(n15347), .Z(
        P2_U3493) );
  MUX2_X1 U16193 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n14177), .S(n15347), .Z(
        P2_U3492) );
  MUX2_X1 U16194 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n14178), .S(n15347), .Z(
        P2_U3491) );
  MUX2_X1 U16195 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n14179), .S(n15347), .Z(
        P2_U3490) );
  MUX2_X1 U16196 ( .A(n14180), .B(P2_REG0_REG_22__SCAN_IN), .S(n15346), .Z(
        P2_U3489) );
  MUX2_X1 U16197 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n14181), .S(n15347), .Z(
        P2_U3488) );
  MUX2_X1 U16198 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n14182), .S(n15347), .Z(
        P2_U3487) );
  MUX2_X1 U16199 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n14183), .S(n15347), .Z(
        P2_U3486) );
  MUX2_X1 U16200 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n14184), .S(n15347), .Z(
        P2_U3484) );
  MUX2_X1 U16201 ( .A(n14185), .B(P2_REG0_REG_17__SCAN_IN), .S(n15346), .Z(
        P2_U3481) );
  INV_X1 U16202 ( .A(n14186), .ZN(n14868) );
  NAND3_X1 U16203 ( .A1(n14187), .A2(P2_IR_REG_31__SCAN_IN), .A3(
        P2_STATE_REG_SCAN_IN), .ZN(n14189) );
  OAI22_X1 U16204 ( .A1(n14190), .A2(n14189), .B1(n14188), .B2(n14201), .ZN(
        n14191) );
  INV_X1 U16205 ( .A(n14191), .ZN(n14192) );
  OAI21_X1 U16206 ( .B1(n14868), .B2(n14196), .A(n14192), .ZN(P2_U3296) );
  OAI222_X1 U16207 ( .A1(n14196), .A2(n14195), .B1(P2_U3088), .B2(n14194), 
        .C1(n14193), .C2(n14201), .ZN(P2_U3298) );
  NAND2_X1 U16208 ( .A1(n14869), .A2(n14197), .ZN(n14199) );
  OAI211_X1 U16209 ( .C1(n14201), .C2(n14200), .A(n14199), .B(n14198), .ZN(
        P2_U3299) );
  INV_X1 U16210 ( .A(n14202), .ZN(n14203) );
  MUX2_X1 U16211 ( .A(n14203), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  OAI21_X1 U16212 ( .B1(n14206), .B2(n14205), .A(n14204), .ZN(n14207) );
  NAND2_X1 U16213 ( .A1(n14356), .A2(n14771), .ZN(n14209) );
  NAND2_X1 U16214 ( .A1(n14358), .A2(n14620), .ZN(n14208) );
  NAND2_X1 U16215 ( .A1(n14209), .A2(n14208), .ZN(n14502) );
  INV_X1 U16216 ( .A(n14511), .ZN(n14211) );
  OAI22_X1 U16217 ( .A1(n14211), .A2(n15072), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14210), .ZN(n14212) );
  AOI21_X1 U16218 ( .B1(n14502), .B2(n14349), .A(n14212), .ZN(n14213) );
  INV_X1 U16219 ( .A(n14214), .ZN(n14303) );
  INV_X1 U16220 ( .A(n14215), .ZN(n14217) );
  NOR3_X1 U16221 ( .A1(n14303), .A2(n14217), .A3(n14216), .ZN(n14219) );
  INV_X1 U16222 ( .A(n14218), .ZN(n14275) );
  OAI21_X1 U16223 ( .B1(n14219), .B2(n14275), .A(n14341), .ZN(n14223) );
  AOI22_X1 U16224 ( .A1(n14620), .A2(n14772), .B1(n14359), .B2(n14771), .ZN(
        n14564) );
  OAI22_X1 U16225 ( .A1(n14564), .A2(n14306), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14220), .ZN(n14221) );
  AOI21_X1 U16226 ( .B1(n14572), .B2(n14338), .A(n14221), .ZN(n14222) );
  OAI211_X1 U16227 ( .C1(n14839), .C2(n14352), .A(n14223), .B(n14222), .ZN(
        P1_U3216) );
  INV_X1 U16228 ( .A(n14650), .ZN(n14852) );
  INV_X1 U16229 ( .A(n14311), .ZN(n14227) );
  OAI21_X1 U16230 ( .B1(n14227), .B2(n14226), .A(n14225), .ZN(n14229) );
  NAND2_X1 U16231 ( .A1(n14311), .A2(n14228), .ZN(n14282) );
  NAND3_X1 U16232 ( .A1(n14229), .A2(n14341), .A3(n14282), .ZN(n14233) );
  AOI22_X1 U16233 ( .A1(n14610), .A2(n14771), .B1(n14620), .B2(n14361), .ZN(
        n14643) );
  NAND2_X1 U16234 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n14486)
         );
  OAI21_X1 U16235 ( .B1(n14306), .B2(n14643), .A(n14486), .ZN(n14230) );
  AOI21_X1 U16236 ( .B1(n14231), .B2(n14338), .A(n14230), .ZN(n14232) );
  OAI211_X1 U16237 ( .C1(n14852), .C2(n14352), .A(n14233), .B(n14232), .ZN(
        P1_U3219) );
  NAND2_X1 U16238 ( .A1(n14235), .A2(n14234), .ZN(n14237) );
  AOI21_X1 U16239 ( .B1(n14237), .B2(n14236), .A(n6697), .ZN(n14243) );
  OAI22_X1 U16240 ( .A1(n15056), .A2(n14239), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14238), .ZN(n14241) );
  OAI22_X1 U16241 ( .A1(n15055), .A2(n14607), .B1(n15072), .B2(n14602), .ZN(
        n14240) );
  AOI211_X1 U16242 ( .C1(n14601), .C2(n15067), .A(n14241), .B(n14240), .ZN(
        n14242) );
  OAI21_X1 U16243 ( .B1(n14243), .B2(n15062), .A(n14242), .ZN(P1_U3223) );
  NOR3_X1 U16244 ( .A1(n6698), .A2(n7346), .A3(n14245), .ZN(n14248) );
  INV_X1 U16245 ( .A(n14246), .ZN(n14247) );
  OAI21_X1 U16246 ( .B1(n14248), .B2(n14247), .A(n14341), .ZN(n14253) );
  AND2_X1 U16247 ( .A1(n14359), .A2(n14620), .ZN(n14249) );
  AOI21_X1 U16248 ( .B1(n14358), .B2(n14771), .A(n14249), .ZN(n14534) );
  OAI22_X1 U16249 ( .A1(n14534), .A2(n14306), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14250), .ZN(n14251) );
  AOI21_X1 U16250 ( .B1(n14537), .B2(n14338), .A(n14251), .ZN(n14252) );
  OAI211_X1 U16251 ( .C1(n14254), .C2(n14352), .A(n14253), .B(n14252), .ZN(
        P1_U3225) );
  INV_X1 U16252 ( .A(n14255), .ZN(n14256) );
  AOI21_X1 U16253 ( .B1(n14258), .B2(n14257), .A(n14256), .ZN(n14263) );
  OAI21_X1 U16254 ( .B1(n15056), .B2(n15040), .A(n14259), .ZN(n14261) );
  OAI22_X1 U16255 ( .A1(n15055), .A2(n14701), .B1(n15072), .B2(n14707), .ZN(
        n14260) );
  AOI211_X1 U16256 ( .C1(n14807), .C2(n15067), .A(n14261), .B(n14260), .ZN(
        n14262) );
  OAI21_X1 U16257 ( .B1(n14263), .B2(n15062), .A(n14262), .ZN(P1_U3226) );
  NAND2_X1 U16258 ( .A1(n14265), .A2(n14264), .ZN(n14266) );
  XNOR2_X1 U16259 ( .A(n14267), .B(n14266), .ZN(n14272) );
  OAI21_X1 U16260 ( .B1(n15056), .B2(n14681), .A(n14268), .ZN(n14270) );
  OAI22_X1 U16261 ( .A1(n15055), .A2(n14680), .B1(n14684), .B2(n15072), .ZN(
        n14269) );
  AOI211_X1 U16262 ( .C1(n14683), .C2(n15067), .A(n14270), .B(n14269), .ZN(
        n14271) );
  OAI21_X1 U16263 ( .B1(n14272), .B2(n15062), .A(n14271), .ZN(P1_U3228) );
  INV_X1 U16264 ( .A(n14757), .ZN(n14557) );
  NOR3_X1 U16265 ( .A1(n14275), .A2(n7347), .A3(n14274), .ZN(n14276) );
  OAI21_X1 U16266 ( .B1(n14276), .B2(n6698), .A(n14341), .ZN(n14280) );
  NOR2_X1 U16267 ( .A1(n14545), .A2(n15056), .ZN(n14278) );
  OAI22_X1 U16268 ( .A1(n14546), .A2(n15055), .B1(n15072), .B2(n14554), .ZN(
        n14277) );
  AOI211_X1 U16269 ( .C1(P1_REG3_REG_24__SCAN_IN), .C2(P1_U3086), .A(n14278), 
        .B(n14277), .ZN(n14279) );
  OAI211_X1 U16270 ( .C1(n14557), .C2(n14352), .A(n14280), .B(n14279), .ZN(
        P1_U3229) );
  NAND2_X1 U16271 ( .A1(n14282), .A2(n14281), .ZN(n14284) );
  XNOR2_X1 U16272 ( .A(n14284), .B(n14283), .ZN(n14290) );
  OAI22_X1 U16273 ( .A1(n15056), .A2(n14658), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14285), .ZN(n14288) );
  OAI22_X1 U16274 ( .A1(n15055), .A2(n14286), .B1(n15072), .B2(n14631), .ZN(
        n14287) );
  AOI211_X1 U16275 ( .C1(n14633), .C2(n15067), .A(n14288), .B(n14287), .ZN(
        n14289) );
  OAI21_X1 U16276 ( .B1(n14290), .B2(n15062), .A(n14289), .ZN(P1_U3233) );
  OAI211_X1 U16277 ( .C1(n14292), .C2(n14291), .A(n15044), .B(n14341), .ZN(
        n14299) );
  INV_X1 U16278 ( .A(n14293), .ZN(n14297) );
  OAI22_X1 U16279 ( .A1(n15055), .A2(n14295), .B1(n14294), .B2(n15072), .ZN(
        n14296) );
  AOI211_X1 U16280 ( .C1(n14322), .C2(n14367), .A(n14297), .B(n14296), .ZN(
        n14298) );
  OAI211_X1 U16281 ( .C1(n14300), .C2(n14352), .A(n14299), .B(n14298), .ZN(
        P1_U3234) );
  NOR3_X1 U16282 ( .A1(n6697), .A2(n7353), .A3(n14302), .ZN(n14304) );
  OAI21_X1 U16283 ( .B1(n14304), .B2(n14303), .A(n14341), .ZN(n14309) );
  AOI22_X1 U16284 ( .A1(n14360), .A2(n14771), .B1(n14620), .B2(n14621), .ZN(
        n14584) );
  OAI22_X1 U16285 ( .A1(n14584), .A2(n14306), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n14305), .ZN(n14307) );
  AOI21_X1 U16286 ( .B1(n14592), .B2(n14338), .A(n14307), .ZN(n14308) );
  OAI211_X1 U16287 ( .C1(n14352), .C2(n14843), .A(n14309), .B(n14308), .ZN(
        P1_U3235) );
  OAI21_X1 U16288 ( .B1(n14312), .B2(n14310), .A(n14311), .ZN(n14313) );
  NAND2_X1 U16289 ( .A1(n14313), .A2(n14341), .ZN(n14317) );
  NAND2_X1 U16290 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n15126)
         );
  INV_X1 U16291 ( .A(n15126), .ZN(n14315) );
  OAI22_X1 U16292 ( .A1(n15055), .A2(n14658), .B1(n15072), .B2(n14669), .ZN(
        n14314) );
  AOI211_X1 U16293 ( .C1(n14322), .C2(n14362), .A(n14315), .B(n14314), .ZN(
        n14316) );
  OAI211_X1 U16294 ( .C1(n14668), .C2(n14352), .A(n14317), .B(n14316), .ZN(
        P1_U3238) );
  OAI211_X1 U16295 ( .C1(n14320), .C2(n14319), .A(n14318), .B(n14341), .ZN(
        n14328) );
  AOI22_X1 U16296 ( .A1(n14322), .A2(n14374), .B1(n14321), .B2(n14372), .ZN(
        n14327) );
  NOR2_X1 U16297 ( .A1(n15072), .A2(n14323), .ZN(n14324) );
  AOI211_X1 U16298 ( .C1(n15158), .C2(n15067), .A(n14325), .B(n14324), .ZN(
        n14326) );
  NAND3_X1 U16299 ( .A1(n14328), .A2(n14327), .A3(n14326), .ZN(P1_U3239) );
  OAI21_X1 U16300 ( .B1(n14332), .B2(n14331), .A(n14330), .ZN(n14333) );
  NAND2_X1 U16301 ( .A1(n14333), .A2(n14341), .ZN(n14340) );
  INV_X1 U16302 ( .A(n14334), .ZN(n14518) );
  NOR2_X1 U16303 ( .A1(n14335), .A2(n14702), .ZN(n14522) );
  AOI22_X1 U16304 ( .A1(n14522), .A2(n14349), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n14336) );
  OAI21_X1 U16305 ( .B1(n14546), .B2(n15056), .A(n14336), .ZN(n14337) );
  AOI21_X1 U16306 ( .B1(n14518), .B2(n14338), .A(n14337), .ZN(n14339) );
  OAI211_X1 U16307 ( .C1(n7044), .C2(n14352), .A(n14340), .B(n14339), .ZN(
        P1_U3240) );
  OAI211_X1 U16308 ( .C1(n14344), .C2(n14343), .A(n14342), .B(n14341), .ZN(
        n14351) );
  NAND2_X1 U16309 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n15113)
         );
  INV_X1 U16310 ( .A(n15113), .ZN(n14347) );
  NOR2_X1 U16311 ( .A1(n15072), .A2(n14345), .ZN(n14346) );
  AOI211_X1 U16312 ( .C1(n14349), .C2(n14348), .A(n14347), .B(n14346), .ZN(
        n14350) );
  OAI211_X1 U16313 ( .C1(n14353), .C2(n14352), .A(n14351), .B(n14350), .ZN(
        P1_U3241) );
  MUX2_X1 U16314 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(n14491), .S(n14379), .Z(
        P1_U3591) );
  MUX2_X1 U16315 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n14354), .S(P1_U4016), .Z(
        P1_U3590) );
  MUX2_X1 U16316 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n14355), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U16317 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n14356), .S(P1_U4016), .Z(
        P1_U3588) );
  MUX2_X1 U16318 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n14357), .S(P1_U4016), .Z(
        P1_U3587) );
  MUX2_X1 U16319 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n14358), .S(P1_U4016), .Z(
        P1_U3586) );
  MUX2_X1 U16320 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n14524), .S(P1_U4016), .Z(
        P1_U3585) );
  MUX2_X1 U16321 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n14359), .S(P1_U4016), .Z(
        P1_U3584) );
  MUX2_X1 U16322 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(n14360), .S(P1_U4016), .Z(
        P1_U3583) );
  MUX2_X1 U16323 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n14772), .S(n14379), .Z(
        P1_U3582) );
  MUX2_X1 U16324 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n14621), .S(n14379), .Z(
        P1_U3581) );
  MUX2_X1 U16325 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n14610), .S(n14379), .Z(
        P1_U3580) );
  MUX2_X1 U16326 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n14619), .S(n14379), .Z(
        P1_U3579) );
  MUX2_X1 U16327 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n14361), .S(n14379), .Z(
        P1_U3578) );
  MUX2_X1 U16328 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n14362), .S(P1_U4016), .Z(
        P1_U3577) );
  MUX2_X1 U16329 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n14363), .S(P1_U4016), .Z(
        P1_U3576) );
  MUX2_X1 U16330 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14364), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U16331 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n14365), .S(P1_U4016), .Z(
        P1_U3574) );
  MUX2_X1 U16332 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n14366), .S(P1_U4016), .Z(
        P1_U3573) );
  MUX2_X1 U16333 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n14367), .S(P1_U4016), .Z(
        P1_U3572) );
  MUX2_X1 U16334 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n14368), .S(P1_U4016), .Z(
        P1_U3571) );
  MUX2_X1 U16335 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n14369), .S(P1_U4016), .Z(
        P1_U3570) );
  MUX2_X1 U16336 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n14370), .S(n14379), .Z(
        P1_U3569) );
  MUX2_X1 U16337 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n14371), .S(n14379), .Z(
        P1_U3568) );
  MUX2_X1 U16338 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n14372), .S(n14379), .Z(
        P1_U3567) );
  MUX2_X1 U16339 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n14373), .S(P1_U4016), .Z(
        P1_U3566) );
  MUX2_X1 U16340 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n14374), .S(n14379), .Z(
        P1_U3565) );
  MUX2_X1 U16341 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n14375), .S(n14379), .Z(
        P1_U3564) );
  MUX2_X1 U16342 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n14376), .S(n14379), .Z(
        P1_U3563) );
  MUX2_X1 U16343 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n14377), .S(n14379), .Z(
        P1_U3562) );
  MUX2_X1 U16344 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n14378), .S(n14379), .Z(
        P1_U3561) );
  MUX2_X1 U16345 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n14380), .S(n14379), .Z(
        P1_U3560) );
  OAI211_X1 U16346 ( .C1(n14383), .C2(n14382), .A(n14477), .B(n14381), .ZN(
        n14392) );
  OAI211_X1 U16347 ( .C1(n14386), .C2(n14385), .A(n14482), .B(n14384), .ZN(
        n14391) );
  AOI22_X1 U16348 ( .A1(n14435), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n14390) );
  INV_X1 U16349 ( .A(n14387), .ZN(n14388) );
  NAND2_X1 U16350 ( .A1(n14480), .A2(n14388), .ZN(n14389) );
  NAND4_X1 U16351 ( .A1(n14392), .A2(n14391), .A3(n14390), .A4(n14389), .ZN(
        P1_U3244) );
  OAI22_X1 U16352 ( .A1(n15128), .A2(n14393), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n15141), .ZN(n14394) );
  AOI21_X1 U16353 ( .B1(n14395), .B2(n14480), .A(n14394), .ZN(n14410) );
  MUX2_X1 U16354 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n10833), .S(n14402), .Z(
        n14398) );
  INV_X1 U16355 ( .A(n14396), .ZN(n14397) );
  NAND3_X1 U16356 ( .A1(n14399), .A2(n14398), .A3(n14397), .ZN(n14400) );
  NAND3_X1 U16357 ( .A1(n14477), .A2(n14401), .A3(n14400), .ZN(n14409) );
  MUX2_X1 U16358 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n10332), .S(n14402), .Z(
        n14404) );
  NAND3_X1 U16359 ( .A1(n14405), .A2(n14404), .A3(n14403), .ZN(n14406) );
  NAND3_X1 U16360 ( .A1(n14482), .A2(n14407), .A3(n14406), .ZN(n14408) );
  NAND3_X1 U16361 ( .A1(n14410), .A2(n14409), .A3(n14408), .ZN(P1_U3246) );
  AOI21_X1 U16362 ( .B1(n14412), .B2(n14411), .A(n15124), .ZN(n14414) );
  NAND2_X1 U16363 ( .A1(n14414), .A2(n14413), .ZN(n14426) );
  NOR2_X1 U16364 ( .A1(n15128), .A2(n14415), .ZN(n14416) );
  AOI211_X1 U16365 ( .C1(n14480), .C2(n14418), .A(n14417), .B(n14416), .ZN(
        n14425) );
  OR3_X1 U16366 ( .A1(n14421), .A2(n14420), .A3(n14419), .ZN(n14422) );
  NAND3_X1 U16367 ( .A1(n14423), .A2(n14482), .A3(n14422), .ZN(n14424) );
  NAND3_X1 U16368 ( .A1(n14426), .A2(n14425), .A3(n14424), .ZN(P1_U3253) );
  INV_X1 U16369 ( .A(n14427), .ZN(n14432) );
  NOR3_X1 U16370 ( .A1(n14430), .A2(n14429), .A3(n14428), .ZN(n14431) );
  OAI21_X1 U16371 ( .B1(n14432), .B2(n14431), .A(n14477), .ZN(n14444) );
  NOR2_X1 U16372 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n14433), .ZN(n14434) );
  AOI21_X1 U16373 ( .B1(n14435), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n14434), 
        .ZN(n14443) );
  OAI21_X1 U16374 ( .B1(n14438), .B2(n14437), .A(n14436), .ZN(n14439) );
  NAND2_X1 U16375 ( .A1(n14439), .A2(n14482), .ZN(n14442) );
  NAND2_X1 U16376 ( .A1(n14480), .A2(n14440), .ZN(n14441) );
  NAND4_X1 U16377 ( .A1(n14444), .A2(n14443), .A3(n14442), .A4(n14441), .ZN(
        P1_U3255) );
  OAI21_X1 U16378 ( .B1(n14447), .B2(n14446), .A(n14445), .ZN(n14448) );
  NAND2_X1 U16379 ( .A1(n14448), .A2(n14477), .ZN(n14461) );
  NAND2_X1 U16380 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n15051)
         );
  OAI21_X1 U16381 ( .B1(n15128), .B2(n14449), .A(n15051), .ZN(n14450) );
  AOI21_X1 U16382 ( .B1(n14451), .B2(n14480), .A(n14450), .ZN(n14460) );
  MUX2_X1 U16383 ( .A(n14452), .B(P1_REG2_REG_14__SCAN_IN), .S(n14451), .Z(
        n14455) );
  INV_X1 U16384 ( .A(n14453), .ZN(n14454) );
  NAND2_X1 U16385 ( .A1(n14455), .A2(n14454), .ZN(n14457) );
  OAI211_X1 U16386 ( .C1(n14458), .C2(n14457), .A(n14456), .B(n14482), .ZN(
        n14459) );
  NAND3_X1 U16387 ( .A1(n14461), .A2(n14460), .A3(n14459), .ZN(P1_U3257) );
  OAI21_X1 U16388 ( .B1(n14802), .B2(n14463), .A(n14462), .ZN(n14464) );
  NAND2_X1 U16389 ( .A1(n14474), .A2(n14464), .ZN(n14465) );
  NAND2_X1 U16390 ( .A1(n15116), .A2(n14465), .ZN(n14466) );
  XOR2_X1 U16391 ( .A(n14466), .B(P1_REG1_REG_19__SCAN_IN), .Z(n14479) );
  NAND2_X1 U16392 ( .A1(n14467), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n14472) );
  INV_X1 U16393 ( .A(n14468), .ZN(n14469) );
  NAND2_X1 U16394 ( .A1(n14470), .A2(n14469), .ZN(n14471) );
  NAND2_X1 U16395 ( .A1(n14472), .A2(n14471), .ZN(n14473) );
  XOR2_X1 U16396 ( .A(n14474), .B(n14473), .Z(n15119) );
  NAND2_X1 U16397 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n15119), .ZN(n15118) );
  NAND2_X1 U16398 ( .A1(n14474), .A2(n14473), .ZN(n14475) );
  NAND2_X1 U16399 ( .A1(n15118), .A2(n14475), .ZN(n14476) );
  XOR2_X1 U16400 ( .A(n14476), .B(P1_REG2_REG_19__SCAN_IN), .Z(n14478) );
  AOI22_X1 U16401 ( .A1(n14479), .A2(n14477), .B1(n14482), .B2(n14478), .ZN(
        n14485) );
  INV_X1 U16402 ( .A(n14478), .ZN(n14481) );
  MUX2_X1 U16403 ( .A(n14485), .B(n14484), .S(n14483), .Z(n14487) );
  OAI211_X1 U16404 ( .C1(n8355), .C2(n15128), .A(n14487), .B(n14486), .ZN(
        P1_U3262) );
  NAND2_X1 U16405 ( .A1(n14717), .A2(n14713), .ZN(n14494) );
  AND2_X1 U16406 ( .A1(n14491), .A2(n14490), .ZN(n14720) );
  INV_X1 U16407 ( .A(n14720), .ZN(n14492) );
  NOR2_X1 U16408 ( .A1(n15143), .A2(n14492), .ZN(n14498) );
  AOI21_X1 U16409 ( .B1(n15143), .B2(P1_REG2_REG_31__SCAN_IN), .A(n14498), 
        .ZN(n14493) );
  OAI211_X1 U16410 ( .C1(n14820), .C2(n14709), .A(n14494), .B(n14493), .ZN(
        P1_U3263) );
  INV_X1 U16411 ( .A(n14495), .ZN(n14496) );
  NAND2_X1 U16412 ( .A1(n14721), .A2(n14713), .ZN(n14500) );
  AOI21_X1 U16413 ( .B1(n15143), .B2(P1_REG2_REG_30__SCAN_IN), .A(n14498), 
        .ZN(n14499) );
  OAI211_X1 U16414 ( .C1(n14824), .C2(n14709), .A(n14500), .B(n14499), .ZN(
        P1_U3264) );
  XNOR2_X1 U16415 ( .A(n14501), .B(n12935), .ZN(n14503) );
  AOI21_X1 U16416 ( .B1(n14503), .B2(n14618), .A(n14502), .ZN(n14741) );
  NAND2_X1 U16417 ( .A1(n14505), .A2(n14504), .ZN(n14506) );
  NAND2_X1 U16418 ( .A1(n14507), .A2(n14506), .ZN(n14739) );
  AOI21_X1 U16419 ( .B1(n14508), .B2(n14517), .A(n14781), .ZN(n14510) );
  NAND2_X1 U16420 ( .A1(n14738), .A2(n14713), .ZN(n14513) );
  AOI22_X1 U16421 ( .A1(n14511), .A2(n15142), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n15143), .ZN(n14512) );
  OAI211_X1 U16422 ( .C1(n14830), .C2(n14709), .A(n14513), .B(n14512), .ZN(
        n14514) );
  AOI21_X1 U16423 ( .B1(n14739), .B2(n14649), .A(n14514), .ZN(n14515) );
  OAI21_X1 U16424 ( .B1(n14741), .B2(n15143), .A(n14515), .ZN(P1_U3266) );
  XNOR2_X1 U16425 ( .A(n14516), .B(n14520), .ZN(n14748) );
  INV_X1 U16426 ( .A(n14748), .ZN(n14529) );
  OAI211_X1 U16427 ( .C1(n7044), .C2(n6679), .A(n14811), .B(n14517), .ZN(
        n14744) );
  INV_X1 U16428 ( .A(n14744), .ZN(n14527) );
  AOI22_X1 U16429 ( .A1(n14518), .A2(n15142), .B1(P1_REG2_REG_26__SCAN_IN), 
        .B2(n15143), .ZN(n14519) );
  OAI21_X1 U16430 ( .B1(n7044), .B2(n14709), .A(n14519), .ZN(n14526) );
  XNOR2_X1 U16431 ( .A(n14521), .B(n14520), .ZN(n14523) );
  AOI21_X1 U16432 ( .B1(n14523), .B2(n14618), .A(n14522), .ZN(n14746) );
  NAND2_X1 U16433 ( .A1(n14524), .A2(n14620), .ZN(n14745) );
  AOI21_X1 U16434 ( .B1(n14746), .B2(n14745), .A(n15143), .ZN(n14525) );
  AOI211_X1 U16435 ( .C1(n14527), .C2(n14713), .A(n14526), .B(n14525), .ZN(
        n14528) );
  OAI21_X1 U16436 ( .B1(n14529), .B2(n14716), .A(n14528), .ZN(P1_U3267) );
  OAI21_X1 U16437 ( .B1(n6724), .B2(n14531), .A(n14530), .ZN(n14755) );
  OAI21_X1 U16438 ( .B1(n6722), .B2(n14533), .A(n14532), .ZN(n14536) );
  INV_X1 U16439 ( .A(n14534), .ZN(n14535) );
  AOI21_X1 U16440 ( .B1(n14536), .B2(n14618), .A(n14535), .ZN(n14754) );
  AOI21_X1 U16441 ( .B1(n14751), .B2(n7048), .A(n6679), .ZN(n14752) );
  AOI22_X1 U16442 ( .A1(n14752), .A2(n14538), .B1(n14537), .B2(n15142), .ZN(
        n14539) );
  AOI21_X1 U16443 ( .B1(n14754), .B2(n14539), .A(n15143), .ZN(n14540) );
  INV_X1 U16444 ( .A(n14540), .ZN(n14542) );
  AOI22_X1 U16445 ( .A1(n14751), .A2(n15140), .B1(P1_REG2_REG_25__SCAN_IN), 
        .B2(n15143), .ZN(n14541) );
  OAI211_X1 U16446 ( .C1(n14755), .C2(n14716), .A(n14542), .B(n14541), .ZN(
        P1_U3268) );
  OAI21_X1 U16447 ( .B1(n14544), .B2(n14550), .A(n14543), .ZN(n14558) );
  OAI22_X1 U16448 ( .A1(n14546), .A2(n14702), .B1(n14545), .B2(n14700), .ZN(
        n14552) );
  INV_X1 U16449 ( .A(n14547), .ZN(n14548) );
  AOI211_X1 U16450 ( .C1(n14550), .C2(n14549), .A(n14699), .B(n14548), .ZN(
        n14551) );
  AOI211_X1 U16451 ( .C1(n14665), .C2(n14558), .A(n14552), .B(n14551), .ZN(
        n14759) );
  AOI211_X1 U16452 ( .C1(n14757), .C2(n14571), .A(n14781), .B(n14553), .ZN(
        n14756) );
  INV_X1 U16453 ( .A(n14554), .ZN(n14555) );
  AOI22_X1 U16454 ( .A1(n15143), .A2(P1_REG2_REG_24__SCAN_IN), .B1(n14555), 
        .B2(n15142), .ZN(n14556) );
  OAI21_X1 U16455 ( .B1(n14557), .B2(n14709), .A(n14556), .ZN(n14560) );
  INV_X1 U16456 ( .A(n14558), .ZN(n14760) );
  NOR2_X1 U16457 ( .A1(n14760), .A2(n14673), .ZN(n14559) );
  AOI211_X1 U16458 ( .C1(n14756), .C2(n14713), .A(n14560), .B(n14559), .ZN(
        n14561) );
  OAI21_X1 U16459 ( .B1(n14759), .B2(n15143), .A(n14561), .ZN(P1_U3269) );
  XNOR2_X1 U16460 ( .A(n14563), .B(n14562), .ZN(n14565) );
  OAI21_X1 U16461 ( .B1(n14565), .B2(n14699), .A(n14564), .ZN(n14761) );
  INV_X1 U16462 ( .A(n14761), .ZN(n14577) );
  INV_X1 U16463 ( .A(n14567), .ZN(n14568) );
  AOI21_X1 U16464 ( .B1(n14569), .B2(n14566), .A(n14568), .ZN(n14763) );
  OR2_X1 U16465 ( .A1(n14839), .A2(n14589), .ZN(n14570) );
  AND3_X1 U16466 ( .A1(n14571), .A2(n14811), .A3(n14570), .ZN(n14762) );
  NAND2_X1 U16467 ( .A1(n14762), .A2(n14713), .ZN(n14574) );
  AOI22_X1 U16468 ( .A1(n15143), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n14572), 
        .B2(n15142), .ZN(n14573) );
  OAI211_X1 U16469 ( .C1(n14839), .C2(n14709), .A(n14574), .B(n14573), .ZN(
        n14575) );
  AOI21_X1 U16470 ( .B1(n14763), .B2(n14649), .A(n14575), .ZN(n14576) );
  OAI21_X1 U16471 ( .B1(n15143), .B2(n14577), .A(n14576), .ZN(P1_U3270) );
  INV_X1 U16472 ( .A(n14578), .ZN(n14583) );
  AOI21_X1 U16473 ( .B1(n14579), .B2(n14581), .A(n14580), .ZN(n14582) );
  OAI21_X1 U16474 ( .B1(n14583), .B2(n14582), .A(n14618), .ZN(n14585) );
  NAND2_X1 U16475 ( .A1(n14585), .A2(n14584), .ZN(n14766) );
  INV_X1 U16476 ( .A(n14766), .ZN(n14597) );
  OAI21_X1 U16477 ( .B1(n14588), .B2(n14587), .A(n14586), .ZN(n14768) );
  INV_X1 U16478 ( .A(n14599), .ZN(n14590) );
  AOI211_X1 U16479 ( .C1(n14591), .C2(n14590), .A(n14781), .B(n14589), .ZN(
        n14767) );
  NAND2_X1 U16480 ( .A1(n14767), .A2(n14713), .ZN(n14594) );
  AOI22_X1 U16481 ( .A1(n15143), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n14592), 
        .B2(n15142), .ZN(n14593) );
  OAI211_X1 U16482 ( .C1(n14709), .C2(n14843), .A(n14594), .B(n14593), .ZN(
        n14595) );
  AOI21_X1 U16483 ( .B1(n14768), .B2(n14649), .A(n14595), .ZN(n14596) );
  OAI21_X1 U16484 ( .B1(n14597), .B2(n15143), .A(n14596), .ZN(P1_U3271) );
  XNOR2_X1 U16485 ( .A(n14598), .B(n12927), .ZN(n14777) );
  OAI21_X1 U16486 ( .B1(n14628), .B2(n14847), .A(n14811), .ZN(n14600) );
  OR2_X1 U16487 ( .A1(n14600), .A2(n14599), .ZN(n14774) );
  INV_X1 U16488 ( .A(n14774), .ZN(n14615) );
  NAND2_X1 U16489 ( .A1(n14601), .A2(n15140), .ZN(n14605) );
  NOR2_X1 U16490 ( .A1(n14602), .A2(n14706), .ZN(n14603) );
  AOI21_X1 U16491 ( .B1(n15143), .B2(P1_REG2_REG_21__SCAN_IN), .A(n14603), 
        .ZN(n14604) );
  OAI211_X1 U16492 ( .C1(n14607), .C2(n14606), .A(n14605), .B(n14604), .ZN(
        n14614) );
  OAI211_X1 U16493 ( .C1(n14609), .C2(n14608), .A(n14579), .B(n14618), .ZN(
        n14612) );
  NAND2_X1 U16494 ( .A1(n14610), .A2(n14620), .ZN(n14611) );
  AND2_X1 U16495 ( .A1(n14612), .A2(n14611), .ZN(n14776) );
  NOR2_X1 U16496 ( .A1(n14776), .A2(n15143), .ZN(n14613) );
  AOI211_X1 U16497 ( .C1(n14615), .C2(n14713), .A(n14614), .B(n14613), .ZN(
        n14616) );
  OAI21_X1 U16498 ( .B1(n14777), .B2(n14716), .A(n14616), .ZN(P1_U3272) );
  OAI211_X1 U16499 ( .C1(n6769), .C2(n14627), .A(n14617), .B(n14618), .ZN(
        n14623) );
  AOI22_X1 U16500 ( .A1(n14621), .A2(n14771), .B1(n14620), .B2(n14619), .ZN(
        n14622) );
  NAND2_X1 U16501 ( .A1(n14623), .A2(n14622), .ZN(n14783) );
  INV_X1 U16502 ( .A(n14783), .ZN(n14638) );
  INV_X1 U16503 ( .A(n14624), .ZN(n14625) );
  AOI21_X1 U16504 ( .B1(n14627), .B2(n14626), .A(n14625), .ZN(n14785) );
  AND2_X1 U16505 ( .A1(n14651), .A2(n14633), .ZN(n14629) );
  OR2_X1 U16506 ( .A1(n14629), .A2(n14628), .ZN(n14782) );
  NAND2_X1 U16507 ( .A1(n15143), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n14630) );
  OAI21_X1 U16508 ( .B1(n14706), .B2(n14631), .A(n14630), .ZN(n14632) );
  AOI21_X1 U16509 ( .B1(n14633), .B2(n15140), .A(n14632), .ZN(n14634) );
  OAI21_X1 U16510 ( .B1(n14782), .B2(n14635), .A(n14634), .ZN(n14636) );
  AOI21_X1 U16511 ( .B1(n14785), .B2(n14649), .A(n14636), .ZN(n14637) );
  OAI21_X1 U16512 ( .B1(n15143), .B2(n14638), .A(n14637), .ZN(P1_U3273) );
  INV_X1 U16513 ( .A(n14639), .ZN(n14640) );
  AOI21_X1 U16514 ( .B1(n14642), .B2(n6860), .A(n14640), .ZN(n14644) );
  OAI21_X1 U16515 ( .B1(n14644), .B2(n14699), .A(n14643), .ZN(n14787) );
  NAND2_X1 U16516 ( .A1(n14787), .A2(n14708), .ZN(n14656) );
  NAND2_X1 U16517 ( .A1(n15143), .A2(P1_REG2_REG_19__SCAN_IN), .ZN(n14645) );
  OAI21_X1 U16518 ( .B1(n14706), .B2(n14646), .A(n14645), .ZN(n14647) );
  AOI21_X1 U16519 ( .B1(n14650), .B2(n15140), .A(n14647), .ZN(n14655) );
  XNOR2_X1 U16520 ( .A(n14648), .B(n14642), .ZN(n14789) );
  NAND2_X1 U16521 ( .A1(n14789), .A2(n14649), .ZN(n14654) );
  AOI21_X1 U16522 ( .B1(n14650), .B2(n14666), .A(n14781), .ZN(n14652) );
  AND2_X1 U16523 ( .A1(n14652), .A2(n14651), .ZN(n14788) );
  NAND2_X1 U16524 ( .A1(n14788), .A2(n14713), .ZN(n14653) );
  NAND4_X1 U16525 ( .A1(n14656), .A2(n14655), .A3(n14654), .A4(n14653), .ZN(
        P1_U3274) );
  XNOR2_X1 U16526 ( .A(n14657), .B(n14662), .ZN(n14792) );
  OAI22_X1 U16527 ( .A1(n14658), .A2(n14702), .B1(n14701), .B2(n14700), .ZN(
        n14664) );
  INV_X1 U16528 ( .A(n14659), .ZN(n14660) );
  AOI211_X1 U16529 ( .C1(n14662), .C2(n14661), .A(n14699), .B(n14660), .ZN(
        n14663) );
  AOI211_X1 U16530 ( .C1(n14792), .C2(n14665), .A(n14664), .B(n14663), .ZN(
        n14796) );
  INV_X1 U16531 ( .A(n14666), .ZN(n14667) );
  AOI211_X1 U16532 ( .C1(n14794), .C2(n7035), .A(n14781), .B(n14667), .ZN(
        n14793) );
  NOR2_X1 U16533 ( .A1(n14668), .A2(n14709), .ZN(n14672) );
  OAI22_X1 U16534 ( .A1(n14708), .A2(n14670), .B1(n14669), .B2(n14706), .ZN(
        n14671) );
  AOI211_X1 U16535 ( .C1(n14793), .C2(n14713), .A(n14672), .B(n14671), .ZN(
        n14675) );
  INV_X1 U16536 ( .A(n14673), .ZN(n15149) );
  NAND2_X1 U16537 ( .A1(n14792), .A2(n15149), .ZN(n14674) );
  OAI211_X1 U16538 ( .C1(n14796), .C2(n15143), .A(n14675), .B(n14674), .ZN(
        P1_U3275) );
  XOR2_X1 U16539 ( .A(n14677), .B(n14676), .Z(n14800) );
  INV_X1 U16540 ( .A(n14800), .ZN(n14690) );
  XOR2_X1 U16541 ( .A(n14678), .B(n14677), .Z(n14679) );
  OAI222_X1 U16542 ( .A1(n14700), .A2(n14681), .B1(n14702), .B2(n14680), .C1(
        n14699), .C2(n14679), .ZN(n14798) );
  NAND2_X1 U16543 ( .A1(n14798), .A2(n14708), .ZN(n14689) );
  AOI211_X1 U16544 ( .C1(n14683), .C2(n14704), .A(n14781), .B(n14682), .ZN(
        n14799) );
  NOR2_X1 U16545 ( .A1(n14859), .A2(n14709), .ZN(n14687) );
  OAI22_X1 U16546 ( .A1(n14708), .A2(n14685), .B1(n14684), .B2(n14706), .ZN(
        n14686) );
  AOI211_X1 U16547 ( .C1(n14799), .C2(n14713), .A(n14687), .B(n14686), .ZN(
        n14688) );
  OAI211_X1 U16548 ( .C1(n14690), .C2(n14716), .A(n14689), .B(n14688), .ZN(
        P1_U3276) );
  OAI21_X1 U16549 ( .B1(n14692), .B2(n14697), .A(n14691), .ZN(n14693) );
  INV_X1 U16550 ( .A(n14693), .ZN(n14809) );
  INV_X1 U16551 ( .A(n14694), .ZN(n14695) );
  AOI21_X1 U16552 ( .B1(n14697), .B2(n14696), .A(n14695), .ZN(n14698) );
  OAI222_X1 U16553 ( .A1(n14702), .A2(n14701), .B1(n14700), .B2(n15040), .C1(
        n14699), .C2(n14698), .ZN(n14805) );
  NAND2_X1 U16554 ( .A1(n14805), .A2(n14708), .ZN(n14715) );
  AOI21_X1 U16555 ( .B1(n14703), .B2(n14807), .A(n14781), .ZN(n14705) );
  AND2_X1 U16556 ( .A1(n14705), .A2(n14704), .ZN(n14806) );
  OAI22_X1 U16557 ( .A1(n14708), .A2(n12020), .B1(n14707), .B2(n14706), .ZN(
        n14712) );
  INV_X1 U16558 ( .A(n14807), .ZN(n14710) );
  NOR2_X1 U16559 ( .A1(n14710), .A2(n14709), .ZN(n14711) );
  AOI211_X1 U16560 ( .C1(n14806), .C2(n14713), .A(n14712), .B(n14711), .ZN(
        n14714) );
  OAI211_X1 U16561 ( .C1(n14809), .C2(n14716), .A(n14715), .B(n14714), .ZN(
        P1_U3277) );
  NOR2_X1 U16562 ( .A1(n14717), .A2(n14720), .ZN(n14817) );
  MUX2_X1 U16563 ( .A(n14718), .B(n14817), .S(n14801), .Z(n14719) );
  OAI21_X1 U16564 ( .B1(n14820), .B2(n14804), .A(n14719), .ZN(P1_U3559) );
  NOR2_X1 U16565 ( .A1(n14721), .A2(n14720), .ZN(n14821) );
  MUX2_X1 U16566 ( .A(n14722), .B(n14821), .S(n14801), .Z(n14723) );
  OAI21_X1 U16567 ( .B1(n14824), .B2(n14804), .A(n14723), .ZN(P1_U3558) );
  INV_X1 U16568 ( .A(n15157), .ZN(n15172) );
  OAI211_X1 U16569 ( .C1(n14726), .C2(n15172), .A(n14725), .B(n14724), .ZN(
        n14727) );
  NOR2_X1 U16570 ( .A1(n14728), .A2(n14727), .ZN(n14729) );
  OAI211_X1 U16571 ( .C1(n14731), .C2(n14815), .A(n14730), .B(n14729), .ZN(
        n14825) );
  MUX2_X1 U16572 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n14825), .S(n15184), .Z(
        P1_U3557) );
  AOI21_X1 U16573 ( .B1(n14734), .B2(n15157), .A(n14733), .ZN(n14735) );
  OAI211_X1 U16574 ( .C1(n14737), .C2(n14815), .A(n14736), .B(n14735), .ZN(
        n14826) );
  MUX2_X1 U16575 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14826), .S(n15184), .Z(
        P1_U3556) );
  INV_X1 U16576 ( .A(P1_REG1_REG_27__SCAN_IN), .ZN(n14742) );
  AOI21_X1 U16577 ( .B1(n14739), .B2(n15175), .A(n14738), .ZN(n14740) );
  AND2_X1 U16578 ( .A1(n14741), .A2(n14740), .ZN(n14827) );
  MUX2_X1 U16579 ( .A(n14742), .B(n14827), .S(n14801), .Z(n14743) );
  OAI21_X1 U16580 ( .B1(n14830), .B2(n14804), .A(n14743), .ZN(P1_U3555) );
  INV_X1 U16581 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n14749) );
  NAND3_X1 U16582 ( .A1(n14746), .A2(n14745), .A3(n14744), .ZN(n14747) );
  AOI21_X1 U16583 ( .B1(n15175), .B2(n14748), .A(n14747), .ZN(n14831) );
  MUX2_X1 U16584 ( .A(n14749), .B(n14831), .S(n14801), .Z(n14750) );
  OAI21_X1 U16585 ( .B1(n7044), .B2(n14804), .A(n14750), .ZN(P1_U3554) );
  AOI22_X1 U16586 ( .A1(n14752), .A2(n14811), .B1(n14751), .B2(n15157), .ZN(
        n14753) );
  OAI211_X1 U16587 ( .C1(n14755), .C2(n14815), .A(n14754), .B(n14753), .ZN(
        n14834) );
  MUX2_X1 U16588 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14834), .S(n15184), .Z(
        P1_U3553) );
  AOI21_X1 U16589 ( .B1(n14757), .B2(n15157), .A(n14756), .ZN(n14758) );
  OAI211_X1 U16590 ( .C1(n14760), .C2(n15161), .A(n14759), .B(n14758), .ZN(
        n14835) );
  MUX2_X1 U16591 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14835), .S(n15184), .Z(
        P1_U3552) );
  INV_X1 U16592 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n14764) );
  AOI211_X1 U16593 ( .C1(n14763), .C2(n15175), .A(n14762), .B(n14761), .ZN(
        n14836) );
  MUX2_X1 U16594 ( .A(n14764), .B(n14836), .S(n14801), .Z(n14765) );
  OAI21_X1 U16595 ( .B1(n14839), .B2(n14804), .A(n14765), .ZN(P1_U3551) );
  INV_X1 U16596 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n14769) );
  AOI211_X1 U16597 ( .C1(n15175), .C2(n14768), .A(n14767), .B(n14766), .ZN(
        n14840) );
  MUX2_X1 U16598 ( .A(n14769), .B(n14840), .S(n14801), .Z(n14770) );
  OAI21_X1 U16599 ( .B1(n14804), .B2(n14843), .A(n14770), .ZN(P1_U3550) );
  NAND2_X1 U16600 ( .A1(n14772), .A2(n14771), .ZN(n14773) );
  AND2_X1 U16601 ( .A1(n14774), .A2(n14773), .ZN(n14775) );
  OAI211_X1 U16602 ( .C1(n14815), .C2(n14777), .A(n14776), .B(n14775), .ZN(
        n14844) );
  MUX2_X1 U16603 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14844), .S(n15184), .Z(
        n14778) );
  INV_X1 U16604 ( .A(n14778), .ZN(n14779) );
  OAI21_X1 U16605 ( .B1(n14847), .B2(n14804), .A(n14779), .ZN(P1_U3549) );
  OAI22_X1 U16606 ( .A1(n14782), .A2(n14781), .B1(n14780), .B2(n15172), .ZN(
        n14784) );
  AOI211_X1 U16607 ( .C1(n14785), .C2(n15175), .A(n14784), .B(n14783), .ZN(
        n14786) );
  INV_X1 U16608 ( .A(n14786), .ZN(n14848) );
  MUX2_X1 U16609 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14848), .S(n15184), .Z(
        P1_U3548) );
  AOI211_X1 U16610 ( .C1(n14789), .C2(n15175), .A(n14788), .B(n14787), .ZN(
        n14849) );
  MUX2_X1 U16611 ( .A(n14790), .B(n14849), .S(n14801), .Z(n14791) );
  OAI21_X1 U16612 ( .B1(n14852), .B2(n14804), .A(n14791), .ZN(P1_U3547) );
  INV_X1 U16613 ( .A(n14792), .ZN(n14797) );
  AOI21_X1 U16614 ( .B1(n14794), .B2(n15157), .A(n14793), .ZN(n14795) );
  OAI211_X1 U16615 ( .C1(n15161), .C2(n14797), .A(n14796), .B(n14795), .ZN(
        n14853) );
  MUX2_X1 U16616 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n14853), .S(n15184), .Z(
        P1_U3546) );
  AOI211_X1 U16617 ( .C1(n14800), .C2(n15175), .A(n14799), .B(n14798), .ZN(
        n14855) );
  MUX2_X1 U16618 ( .A(n14802), .B(n14855), .S(n14801), .Z(n14803) );
  OAI21_X1 U16619 ( .B1(n14859), .B2(n14804), .A(n14803), .ZN(P1_U3545) );
  AOI211_X1 U16620 ( .C1(n14807), .C2(n15157), .A(n14806), .B(n14805), .ZN(
        n14808) );
  OAI21_X1 U16621 ( .B1(n14815), .B2(n14809), .A(n14808), .ZN(n14860) );
  MUX2_X1 U16622 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n14860), .S(n15184), .Z(
        P1_U3544) );
  AOI22_X1 U16623 ( .A1(n14812), .A2(n14811), .B1(n14810), .B2(n15157), .ZN(
        n14813) );
  OAI211_X1 U16624 ( .C1(n14816), .C2(n14815), .A(n14814), .B(n14813), .ZN(
        n14861) );
  MUX2_X1 U16625 ( .A(P1_REG1_REG_15__SCAN_IN), .B(n14861), .S(n15184), .Z(
        P1_U3543) );
  INV_X1 U16626 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n14818) );
  MUX2_X1 U16627 ( .A(n14818), .B(n14817), .S(n14854), .Z(n14819) );
  OAI21_X1 U16628 ( .B1(n14820), .B2(n14858), .A(n14819), .ZN(P1_U3527) );
  INV_X1 U16629 ( .A(P1_REG0_REG_30__SCAN_IN), .ZN(n14822) );
  MUX2_X1 U16630 ( .A(n14822), .B(n14821), .S(n14854), .Z(n14823) );
  OAI21_X1 U16631 ( .B1(n14824), .B2(n14858), .A(n14823), .ZN(P1_U3526) );
  MUX2_X1 U16632 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14825), .S(n14854), .Z(
        P1_U3525) );
  MUX2_X1 U16633 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14826), .S(n14854), .Z(
        P1_U3524) );
  MUX2_X1 U16634 ( .A(n14828), .B(n14827), .S(n14854), .Z(n14829) );
  OAI21_X1 U16635 ( .B1(n14830), .B2(n14858), .A(n14829), .ZN(P1_U3523) );
  MUX2_X1 U16636 ( .A(n14832), .B(n14831), .S(n14854), .Z(n14833) );
  OAI21_X1 U16637 ( .B1(n7044), .B2(n14858), .A(n14833), .ZN(P1_U3522) );
  MUX2_X1 U16638 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14834), .S(n14854), .Z(
        P1_U3521) );
  MUX2_X1 U16639 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14835), .S(n14854), .Z(
        P1_U3520) );
  MUX2_X1 U16640 ( .A(n14837), .B(n14836), .S(n14854), .Z(n14838) );
  OAI21_X1 U16641 ( .B1(n14839), .B2(n14858), .A(n14838), .ZN(P1_U3519) );
  MUX2_X1 U16642 ( .A(n14841), .B(n14840), .S(n14854), .Z(n14842) );
  OAI21_X1 U16643 ( .B1(n14858), .B2(n14843), .A(n14842), .ZN(P1_U3518) );
  MUX2_X1 U16644 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14844), .S(n14854), .Z(
        n14845) );
  INV_X1 U16645 ( .A(n14845), .ZN(n14846) );
  OAI21_X1 U16646 ( .B1(n14847), .B2(n14858), .A(n14846), .ZN(P1_U3517) );
  MUX2_X1 U16647 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14848), .S(n14854), .Z(
        P1_U3516) );
  MUX2_X1 U16648 ( .A(n14850), .B(n14849), .S(n14854), .Z(n14851) );
  OAI21_X1 U16649 ( .B1(n14852), .B2(n14858), .A(n14851), .ZN(P1_U3515) );
  MUX2_X1 U16650 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n14853), .S(n14854), .Z(
        P1_U3513) );
  INV_X1 U16651 ( .A(P1_REG0_REG_17__SCAN_IN), .ZN(n14856) );
  MUX2_X1 U16652 ( .A(n14856), .B(n14855), .S(n14854), .Z(n14857) );
  OAI21_X1 U16653 ( .B1(n14859), .B2(n14858), .A(n14857), .ZN(P1_U3510) );
  MUX2_X1 U16654 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n14860), .S(n14854), .Z(
        P1_U3507) );
  MUX2_X1 U16655 ( .A(P1_REG0_REG_15__SCAN_IN), .B(n14861), .S(n14854), .Z(
        P1_U3504) );
  NOR4_X1 U16656 ( .A1(n14862), .A2(P1_IR_REG_30__SCAN_IN), .A3(n14864), .A4(
        P1_U3086), .ZN(n14865) );
  AOI21_X1 U16657 ( .B1(n14866), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14865), 
        .ZN(n14867) );
  OAI21_X1 U16658 ( .B1(n14868), .B2(n14874), .A(n14867), .ZN(P1_U3324) );
  INV_X1 U16659 ( .A(n14869), .ZN(n14870) );
  OAI222_X1 U16660 ( .A1(n14876), .A2(n14871), .B1(n14874), .B2(n14870), .C1(
        n10248), .C2(P1_U3086), .ZN(P1_U3327) );
  OAI222_X1 U16661 ( .A1(n14876), .A2(n14875), .B1(n14874), .B2(n14873), .C1(
        P1_U3086), .C2(n14872), .ZN(P1_U3328) );
  MUX2_X1 U16662 ( .A(n14878), .B(n14877), .S(P1_U3086), .Z(P1_U3333) );
  INV_X1 U16663 ( .A(n14879), .ZN(n14880) );
  MUX2_X1 U16664 ( .A(n14880), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U16665 ( .A1(n14882), .A2(n14881), .ZN(n14883) );
  XOR2_X1 U16666 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14883), .Z(SUB_1596_U62)
         );
  AOI21_X1 U16667 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14884) );
  OAI21_X1 U16668 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14884), 
        .ZN(U28) );
  INV_X1 U16669 ( .A(P1_RD_REG_SCAN_IN), .ZN(n14886) );
  INV_X1 U16670 ( .A(P2_RD_REG_SCAN_IN), .ZN(n14887) );
  OAI221_X1 U16671 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(
        n14887), .C2(n14886), .A(n14885), .ZN(U29) );
  OAI21_X1 U16672 ( .B1(n14890), .B2(n14889), .A(n14888), .ZN(n14891) );
  XNOR2_X1 U16673 ( .A(n14891), .B(P2_ADDR_REG_2__SCAN_IN), .ZN(SUB_1596_U61)
         );
  AOI21_X1 U16674 ( .B1(n14894), .B2(n14893), .A(n14892), .ZN(SUB_1596_U57) );
  AOI21_X1 U16675 ( .B1(n14897), .B2(n14896), .A(n14895), .ZN(n14898) );
  XOR2_X1 U16676 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n14898), .Z(SUB_1596_U55) );
  AOI21_X1 U16677 ( .B1(n14901), .B2(n14900), .A(n14899), .ZN(SUB_1596_U54) );
  OAI21_X1 U16678 ( .B1(n14903), .B2(n6796), .A(n14902), .ZN(n14904) );
  XNOR2_X1 U16679 ( .A(n14904), .B(P2_ADDR_REG_10__SCAN_IN), .ZN(SUB_1596_U70)
         );
  OAI21_X1 U16680 ( .B1(n14906), .B2(n15172), .A(n14905), .ZN(n14908) );
  AOI211_X1 U16681 ( .C1(n14910), .C2(n14909), .A(n14908), .B(n14907), .ZN(
        n14913) );
  INV_X1 U16682 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14911) );
  AOI22_X1 U16683 ( .A1(n14854), .A2(n14913), .B1(n14911), .B2(n15177), .ZN(
        P1_U3495) );
  AOI22_X1 U16684 ( .A1(n15184), .A2(n14913), .B1(n14912), .B2(n15181), .ZN(
        P1_U3540) );
  NOR2_X1 U16685 ( .A1(n14915), .A2(n14914), .ZN(n14916) );
  XOR2_X1 U16686 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(n14916), .Z(SUB_1596_U63)
         );
  AOI22_X1 U16687 ( .A1(n15485), .A2(n14917), .B1(n15523), .B2(
        P3_ADDR_REG_18__SCAN_IN), .ZN(n14931) );
  AOI21_X1 U16688 ( .B1(n14920), .B2(n14919), .A(n14918), .ZN(n14930) );
  AOI21_X1 U16689 ( .B1(n14923), .B2(n14922), .A(n14921), .ZN(n14924) );
  OAI21_X1 U16690 ( .B1(n14927), .B2(n14926), .A(n14925), .ZN(n14928) );
  NAND2_X1 U16691 ( .A1(n15504), .A2(n14928), .ZN(n14929) );
  OAI22_X1 U16692 ( .A1(n14934), .A2(n15570), .B1(n15582), .B2(n14933), .ZN(
        n14935) );
  NOR2_X1 U16693 ( .A1(n14936), .A2(n14935), .ZN(n14960) );
  AOI22_X1 U16694 ( .A1(n15607), .A2(n14960), .B1(n14937), .B2(n9022), .ZN(
        P3_U3474) );
  OAI22_X1 U16695 ( .A1(n14939), .A2(n15570), .B1(n15582), .B2(n14938), .ZN(
        n14940) );
  NOR2_X1 U16696 ( .A1(n14941), .A2(n14940), .ZN(n14962) );
  INV_X1 U16697 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n14942) );
  AOI22_X1 U16698 ( .A1(n15607), .A2(n14962), .B1(n14942), .B2(n9022), .ZN(
        P3_U3473) );
  OAI22_X1 U16699 ( .A1(n14944), .A2(n15570), .B1(n15582), .B2(n14943), .ZN(
        n14945) );
  NOR2_X1 U16700 ( .A1(n14946), .A2(n14945), .ZN(n14964) );
  AOI22_X1 U16701 ( .A1(n15607), .A2(n14964), .B1(n14947), .B2(n9022), .ZN(
        P3_U3472) );
  AOI22_X1 U16702 ( .A1(n14949), .A2(n14957), .B1(n15561), .B2(n14948), .ZN(
        n14950) );
  AND2_X1 U16703 ( .A1(n14951), .A2(n14950), .ZN(n14966) );
  INV_X1 U16704 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14952) );
  AOI22_X1 U16705 ( .A1(n15607), .A2(n14966), .B1(n14952), .B2(n9022), .ZN(
        P3_U3471) );
  NOR2_X1 U16706 ( .A1(n14953), .A2(n15582), .ZN(n14955) );
  AOI211_X1 U16707 ( .C1(n14957), .C2(n14956), .A(n14955), .B(n14954), .ZN(
        n14968) );
  AOI22_X1 U16708 ( .A1(n15607), .A2(n14968), .B1(n14958), .B2(n9022), .ZN(
        P3_U3470) );
  INV_X1 U16709 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n14959) );
  AOI22_X1 U16710 ( .A1(n15591), .A2(n14960), .B1(n14959), .B2(n15589), .ZN(
        P3_U3435) );
  INV_X1 U16711 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14961) );
  AOI22_X1 U16712 ( .A1(n15591), .A2(n14962), .B1(n14961), .B2(n15589), .ZN(
        P3_U3432) );
  INV_X1 U16713 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14963) );
  AOI22_X1 U16714 ( .A1(n15591), .A2(n14964), .B1(n14963), .B2(n15589), .ZN(
        P3_U3429) );
  INV_X1 U16715 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14965) );
  AOI22_X1 U16716 ( .A1(n15591), .A2(n14966), .B1(n14965), .B2(n15589), .ZN(
        P3_U3426) );
  INV_X1 U16717 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14967) );
  AOI22_X1 U16718 ( .A1(n15591), .A2(n14968), .B1(n14967), .B2(n15589), .ZN(
        P3_U3423) );
  XNOR2_X1 U16719 ( .A(n14970), .B(n14969), .ZN(n14973) );
  INV_X1 U16720 ( .A(n14971), .ZN(n14972) );
  AOI21_X1 U16721 ( .B1(n14973), .B2(n14065), .A(n14972), .ZN(n15003) );
  AOI222_X1 U16722 ( .A1(n14975), .A2(n15270), .B1(P2_REG2_REG_16__SCAN_IN), 
        .B2(n15269), .C1(n15268), .C2(n14974), .ZN(n14984) );
  INV_X1 U16723 ( .A(n14976), .ZN(n14977) );
  AOI21_X1 U16724 ( .B1(n14979), .B2(n14978), .A(n14977), .ZN(n15006) );
  OAI211_X1 U16725 ( .C1(n15002), .C2(n7059), .A(n15274), .B(n14981), .ZN(
        n15001) );
  INV_X1 U16726 ( .A(n15001), .ZN(n14982) );
  AOI22_X1 U16727 ( .A1(n15006), .A2(n15280), .B1(n14982), .B2(n15279), .ZN(
        n14983) );
  OAI211_X1 U16728 ( .C1(n14078), .C2(n15003), .A(n14984), .B(n14983), .ZN(
        P2_U3249) );
  XNOR2_X1 U16729 ( .A(n14986), .B(n14985), .ZN(n14989) );
  INV_X1 U16730 ( .A(n14987), .ZN(n14988) );
  AOI21_X1 U16731 ( .B1(n14989), .B2(n14065), .A(n14988), .ZN(n15015) );
  AOI222_X1 U16732 ( .A1(n14991), .A2(n15270), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n15269), .C1(n15268), .C2(n14990), .ZN(n14999) );
  AOI21_X1 U16733 ( .B1(n14993), .B2(n14992), .A(n9741), .ZN(n15018) );
  INV_X1 U16734 ( .A(n14994), .ZN(n14995) );
  OAI211_X1 U16735 ( .C1(n15014), .C2(n14996), .A(n14995), .B(n15274), .ZN(
        n15013) );
  INV_X1 U16736 ( .A(n15013), .ZN(n14997) );
  AOI22_X1 U16737 ( .A1(n15018), .A2(n15280), .B1(n14997), .B2(n15279), .ZN(
        n14998) );
  OAI211_X1 U16738 ( .C1(n14078), .C2(n15015), .A(n14999), .B(n14998), .ZN(
        P2_U3251) );
  INV_X1 U16739 ( .A(n15000), .ZN(n15310) );
  OAI21_X1 U16740 ( .B1(n15002), .B2(n15340), .A(n15001), .ZN(n15005) );
  INV_X1 U16741 ( .A(n15003), .ZN(n15004) );
  AOI211_X1 U16742 ( .C1(n15006), .C2(n15310), .A(n15005), .B(n15004), .ZN(
        n15032) );
  AOI22_X1 U16743 ( .A1(n15357), .A2(n15032), .B1(n10073), .B2(n15355), .ZN(
        P2_U3515) );
  OAI21_X1 U16744 ( .B1(n15008), .B2(n15340), .A(n15007), .ZN(n15010) );
  AOI211_X1 U16745 ( .C1(n15310), .C2(n15011), .A(n15010), .B(n15009), .ZN(
        n15034) );
  INV_X1 U16746 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n15012) );
  AOI22_X1 U16747 ( .A1(n15357), .A2(n15034), .B1(n15012), .B2(n15355), .ZN(
        P2_U3514) );
  OAI21_X1 U16748 ( .B1(n15014), .B2(n15340), .A(n15013), .ZN(n15017) );
  INV_X1 U16749 ( .A(n15015), .ZN(n15016) );
  AOI211_X1 U16750 ( .C1(n15018), .C2(n15310), .A(n15017), .B(n15016), .ZN(
        n15036) );
  AOI22_X1 U16751 ( .A1(n15357), .A2(n15036), .B1(n15019), .B2(n15355), .ZN(
        P2_U3513) );
  OAI21_X1 U16752 ( .B1(n15021), .B2(n15340), .A(n15020), .ZN(n15023) );
  AOI211_X1 U16753 ( .C1(n15024), .C2(n15310), .A(n15023), .B(n15022), .ZN(
        n15037) );
  AOI22_X1 U16754 ( .A1(n15357), .A2(n15037), .B1(n10102), .B2(n15355), .ZN(
        P2_U3512) );
  OAI21_X1 U16755 ( .B1(n15026), .B2(n15340), .A(n15025), .ZN(n15027) );
  AOI21_X1 U16756 ( .B1(n15028), .B2(n15310), .A(n15027), .ZN(n15029) );
  AND2_X1 U16757 ( .A1(n15030), .A2(n15029), .ZN(n15039) );
  AOI22_X1 U16758 ( .A1(n15357), .A2(n15039), .B1(n9322), .B2(n15355), .ZN(
        P2_U3511) );
  INV_X1 U16759 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n15031) );
  AOI22_X1 U16760 ( .A1(n15347), .A2(n15032), .B1(n15031), .B2(n15346), .ZN(
        P2_U3478) );
  INV_X1 U16761 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n15033) );
  AOI22_X1 U16762 ( .A1(n15347), .A2(n15034), .B1(n15033), .B2(n15346), .ZN(
        P2_U3475) );
  INV_X1 U16763 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n15035) );
  AOI22_X1 U16764 ( .A1(n15347), .A2(n15036), .B1(n15035), .B2(n15346), .ZN(
        P2_U3472) );
  AOI22_X1 U16765 ( .A1(n15347), .A2(n15037), .B1(n9342), .B2(n15346), .ZN(
        P2_U3469) );
  INV_X1 U16766 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n15038) );
  AOI22_X1 U16767 ( .A1(n15347), .A2(n15039), .B1(n15038), .B2(n15346), .ZN(
        P2_U3466) );
  OAI22_X1 U16768 ( .A1(n15041), .A2(n15056), .B1(n15055), .B2(n15040), .ZN(
        n15049) );
  AOI21_X1 U16769 ( .B1(n15044), .B2(n15043), .A(n15042), .ZN(n15045) );
  INV_X1 U16770 ( .A(n15045), .ZN(n15047) );
  AOI21_X1 U16771 ( .B1(n15047), .B2(n15046), .A(n15062), .ZN(n15048) );
  AOI211_X1 U16772 ( .C1(n15050), .C2(n15067), .A(n15049), .B(n15048), .ZN(
        n15052) );
  OAI211_X1 U16773 ( .C1(n15072), .C2(n15053), .A(n15052), .B(n15051), .ZN(
        P1_U3215) );
  OAI22_X1 U16774 ( .A1(n15057), .A2(n15056), .B1(n15055), .B2(n15054), .ZN(
        n15066) );
  AOI21_X1 U16775 ( .B1(n15060), .B2(n15059), .A(n15058), .ZN(n15061) );
  INV_X1 U16776 ( .A(n15061), .ZN(n15064) );
  AOI21_X1 U16777 ( .B1(n15064), .B2(n15063), .A(n15062), .ZN(n15065) );
  AOI211_X1 U16778 ( .C1(n15068), .C2(n15067), .A(n15066), .B(n15065), .ZN(
        n15070) );
  OAI211_X1 U16779 ( .C1(n15072), .C2(n15071), .A(n15070), .B(n15069), .ZN(
        P1_U3236) );
  OAI21_X1 U16780 ( .B1(n15074), .B2(n15172), .A(n15073), .ZN(n15075) );
  AOI211_X1 U16781 ( .C1(n15077), .C2(n15175), .A(n15076), .B(n15075), .ZN(
        n15079) );
  AOI22_X1 U16782 ( .A1(n15184), .A2(n15079), .B1(n15078), .B2(n15181), .ZN(
        P1_U3542) );
  AOI22_X1 U16783 ( .A1(n14854), .A2(n15079), .B1(n12247), .B2(n15177), .ZN(
        P1_U3501) );
  OAI21_X1 U16784 ( .B1(n15082), .B2(n15081), .A(n15080), .ZN(n15083) );
  XNOR2_X1 U16785 ( .A(n15083), .B(P2_ADDR_REG_11__SCAN_IN), .ZN(SUB_1596_U69)
         );
  OAI222_X1 U16786 ( .A1(n15088), .A2(n15087), .B1(n15088), .B2(n15086), .C1(
        n15085), .C2(n15084), .ZN(SUB_1596_U68) );
  OAI21_X1 U16787 ( .B1(n15091), .B2(n15090), .A(n15089), .ZN(n15092) );
  XNOR2_X1 U16788 ( .A(n15092), .B(P2_ADDR_REG_13__SCAN_IN), .ZN(SUB_1596_U67)
         );
  OAI21_X1 U16789 ( .B1(n15095), .B2(n15094), .A(n15093), .ZN(n15096) );
  XNOR2_X1 U16790 ( .A(n15096), .B(P2_ADDR_REG_14__SCAN_IN), .ZN(SUB_1596_U66)
         );
  AOI21_X1 U16791 ( .B1(n15099), .B2(n15098), .A(n15097), .ZN(n15100) );
  XOR2_X1 U16792 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(n15100), .Z(SUB_1596_U65)
         );
  NOR2_X1 U16793 ( .A1(n15102), .A2(n15101), .ZN(n15103) );
  XNOR2_X1 U16794 ( .A(n15104), .B(n15103), .ZN(SUB_1596_U64) );
  AOI21_X1 U16795 ( .B1(n15106), .B2(P1_REG2_REG_15__SCAN_IN), .A(n15105), 
        .ZN(n15110) );
  AOI21_X1 U16796 ( .B1(n15108), .B2(P1_REG1_REG_15__SCAN_IN), .A(n15107), 
        .ZN(n15109) );
  OAI222_X1 U16797 ( .A1(n15122), .A2(n15111), .B1(n15121), .B2(n15110), .C1(
        n15124), .C2(n15109), .ZN(n15112) );
  INV_X1 U16798 ( .A(n15112), .ZN(n15114) );
  OAI211_X1 U16799 ( .C1(n15115), .C2(n15128), .A(n15114), .B(n15113), .ZN(
        P1_U3258) );
  OAI21_X1 U16800 ( .B1(P1_REG1_REG_18__SCAN_IN), .B2(n15117), .A(n15116), 
        .ZN(n15123) );
  OAI21_X1 U16801 ( .B1(P1_REG2_REG_18__SCAN_IN), .B2(n15119), .A(n15118), 
        .ZN(n15120) );
  OAI222_X1 U16802 ( .A1(n15124), .A2(n15123), .B1(n15122), .B2(n6818), .C1(
        n15121), .C2(n15120), .ZN(n15125) );
  INV_X1 U16803 ( .A(n15125), .ZN(n15127) );
  OAI211_X1 U16804 ( .C1(n15129), .C2(n15128), .A(n15127), .B(n15126), .ZN(
        P1_U3261) );
  AOI22_X1 U16805 ( .A1(n15143), .A2(P1_REG2_REG_5__SCAN_IN), .B1(n15130), 
        .B2(n15142), .ZN(n15133) );
  NAND2_X1 U16806 ( .A1(n15140), .A2(n15131), .ZN(n15132) );
  OAI211_X1 U16807 ( .C1(n15134), .C2(n15146), .A(n15133), .B(n15132), .ZN(
        n15135) );
  AOI21_X1 U16808 ( .B1(n15136), .B2(n15149), .A(n15135), .ZN(n15137) );
  OAI21_X1 U16809 ( .B1(n15143), .B2(n15138), .A(n15137), .ZN(P1_U3288) );
  NAND2_X1 U16810 ( .A1(n15140), .A2(n15139), .ZN(n15145) );
  AOI22_X1 U16811 ( .A1(n15143), .A2(P1_REG2_REG_3__SCAN_IN), .B1(n15142), 
        .B2(n15141), .ZN(n15144) );
  OAI211_X1 U16812 ( .C1(n15147), .C2(n15146), .A(n15145), .B(n15144), .ZN(
        n15148) );
  AOI21_X1 U16813 ( .B1(n15150), .B2(n15149), .A(n15148), .ZN(n15151) );
  OAI21_X1 U16814 ( .B1(n15143), .B2(n15152), .A(n15151), .ZN(P1_U3290) );
  AND2_X1 U16815 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n15153), .ZN(P1_U3294) );
  AND2_X1 U16816 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n15153), .ZN(P1_U3295) );
  AND2_X1 U16817 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n15153), .ZN(P1_U3296) );
  AND2_X1 U16818 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n15153), .ZN(P1_U3297) );
  AND2_X1 U16819 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n15153), .ZN(P1_U3298) );
  AND2_X1 U16820 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n15153), .ZN(P1_U3299) );
  AND2_X1 U16821 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n15153), .ZN(P1_U3300) );
  AND2_X1 U16822 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n15153), .ZN(P1_U3301) );
  AND2_X1 U16823 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n15153), .ZN(P1_U3302) );
  AND2_X1 U16824 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n15153), .ZN(P1_U3303) );
  AND2_X1 U16825 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n15153), .ZN(P1_U3304) );
  AND2_X1 U16826 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n15153), .ZN(P1_U3305) );
  AND2_X1 U16827 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n15153), .ZN(P1_U3306) );
  AND2_X1 U16828 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n15153), .ZN(P1_U3307) );
  AND2_X1 U16829 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n15153), .ZN(P1_U3308) );
  AND2_X1 U16830 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n15153), .ZN(P1_U3309) );
  AND2_X1 U16831 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n15153), .ZN(P1_U3310) );
  AND2_X1 U16832 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n15153), .ZN(P1_U3311) );
  AND2_X1 U16833 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n15153), .ZN(P1_U3312) );
  AND2_X1 U16834 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n15153), .ZN(P1_U3313) );
  AND2_X1 U16835 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n15153), .ZN(P1_U3314) );
  AND2_X1 U16836 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n15153), .ZN(P1_U3315) );
  AND2_X1 U16837 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n15153), .ZN(P1_U3316) );
  AND2_X1 U16838 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n15153), .ZN(P1_U3317) );
  AND2_X1 U16839 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n15153), .ZN(P1_U3318) );
  AND2_X1 U16840 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n15153), .ZN(P1_U3319) );
  AND2_X1 U16841 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n15153), .ZN(P1_U3320) );
  AND2_X1 U16842 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n15153), .ZN(P1_U3321) );
  AND2_X1 U16843 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n15153), .ZN(P1_U3322) );
  AND2_X1 U16844 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n15153), .ZN(P1_U3323) );
  INV_X1 U16845 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n15154) );
  AOI22_X1 U16846 ( .A1(n14854), .A2(n15155), .B1(n15154), .B2(n15177), .ZN(
        P1_U3459) );
  AOI21_X1 U16847 ( .B1(n15158), .B2(n15157), .A(n15156), .ZN(n15159) );
  OAI211_X1 U16848 ( .C1(n15162), .C2(n15161), .A(n15160), .B(n15159), .ZN(
        n15163) );
  INV_X1 U16849 ( .A(n15163), .ZN(n15179) );
  AOI22_X1 U16850 ( .A1(n14854), .A2(n15179), .B1(n11332), .B2(n15177), .ZN(
        P1_U3477) );
  OAI211_X1 U16851 ( .C1(n15166), .C2(n15172), .A(n15165), .B(n15164), .ZN(
        n15167) );
  AOI21_X1 U16852 ( .B1(n15175), .B2(n15168), .A(n15167), .ZN(n15180) );
  INV_X1 U16853 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n15169) );
  AOI22_X1 U16854 ( .A1(n14854), .A2(n15180), .B1(n15169), .B2(n15177), .ZN(
        P1_U3483) );
  OAI211_X1 U16855 ( .C1(n7042), .C2(n15172), .A(n15171), .B(n15170), .ZN(
        n15174) );
  AOI211_X1 U16856 ( .C1(n15176), .C2(n15175), .A(n15174), .B(n15173), .ZN(
        n15183) );
  AOI22_X1 U16857 ( .A1(n14854), .A2(n15183), .B1(n11845), .B2(n15177), .ZN(
        P1_U3489) );
  AOI22_X1 U16858 ( .A1(n15184), .A2(n15179), .B1(n15178), .B2(n15181), .ZN(
        P1_U3534) );
  AOI22_X1 U16859 ( .A1(n15184), .A2(n15180), .B1(n11383), .B2(n15181), .ZN(
        P1_U3536) );
  AOI22_X1 U16860 ( .A1(n15184), .A2(n15183), .B1(n15182), .B2(n15181), .ZN(
        P1_U3538) );
  NOR2_X1 U16861 ( .A1(n15250), .A2(P2_U3947), .ZN(P2_U3087) );
  OAI22_X1 U16862 ( .A1(n15225), .A2(n15185), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n11472), .ZN(n15186) );
  AOI21_X1 U16863 ( .B1(P2_ADDR_REG_1__SCAN_IN), .B2(n15250), .A(n15186), .ZN(
        n15197) );
  INV_X1 U16864 ( .A(n15187), .ZN(n15191) );
  OAI21_X1 U16865 ( .B1(n10047), .B2(n15189), .A(n15188), .ZN(n15190) );
  NAND3_X1 U16866 ( .A1(n15252), .A2(n15191), .A3(n15190), .ZN(n15196) );
  OAI211_X1 U16867 ( .C1(n15194), .C2(n15193), .A(n15255), .B(n15192), .ZN(
        n15195) );
  NAND3_X1 U16868 ( .A1(n15197), .A2(n15196), .A3(n15195), .ZN(P2_U3215) );
  OAI21_X1 U16869 ( .B1(n15212), .B2(n15198), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15199) );
  OAI21_X1 U16870 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15199), .ZN(n15210) );
  OAI211_X1 U16871 ( .C1(n15202), .C2(n15201), .A(n15255), .B(n15200), .ZN(
        n15209) );
  NAND2_X1 U16872 ( .A1(n15204), .A2(n15203), .ZN(n15205) );
  NAND3_X1 U16873 ( .A1(n15252), .A2(n15206), .A3(n15205), .ZN(n15208) );
  NAND2_X1 U16874 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(n15250), .ZN(n15207) );
  NAND4_X1 U16875 ( .A1(n15210), .A2(n15209), .A3(n15208), .A4(n15207), .ZN(
        P2_U3217) );
  OAI21_X1 U16876 ( .B1(n15212), .B2(n15211), .A(P2_STATE_REG_SCAN_IN), .ZN(
        n15213) );
  OAI21_X1 U16877 ( .B1(P2_REG3_REG_6__SCAN_IN), .B2(P2_STATE_REG_SCAN_IN), 
        .A(n15213), .ZN(n15223) );
  OAI211_X1 U16878 ( .C1(n15216), .C2(n15215), .A(n15214), .B(n15252), .ZN(
        n15222) );
  OAI211_X1 U16879 ( .C1(n15219), .C2(n15218), .A(n15255), .B(n15217), .ZN(
        n15221) );
  NAND2_X1 U16880 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n15250), .ZN(n15220) );
  NAND4_X1 U16881 ( .A1(n15223), .A2(n15222), .A3(n15221), .A4(n15220), .ZN(
        P2_U3220) );
  OR2_X1 U16882 ( .A1(n15225), .A2(n15224), .ZN(n15227) );
  OAI211_X1 U16883 ( .C1(n15228), .C2(n7921), .A(n15227), .B(n15226), .ZN(
        n15229) );
  INV_X1 U16884 ( .A(n15229), .ZN(n15238) );
  OAI211_X1 U16885 ( .C1(n15232), .C2(n15231), .A(n15230), .B(n15252), .ZN(
        n15237) );
  OAI211_X1 U16886 ( .C1(n15235), .C2(n15234), .A(n15255), .B(n15233), .ZN(
        n15236) );
  NAND3_X1 U16887 ( .A1(n15238), .A2(n15237), .A3(n15236), .ZN(P2_U3221) );
  AOI22_X1 U16888 ( .A1(n15250), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n15249) );
  OAI211_X1 U16889 ( .C1(n15241), .C2(n15240), .A(n15239), .B(n15252), .ZN(
        n15248) );
  NAND2_X1 U16890 ( .A1(n15259), .A2(n15242), .ZN(n15247) );
  OAI211_X1 U16891 ( .C1(n15245), .C2(n15244), .A(n15243), .B(n15255), .ZN(
        n15246) );
  NAND4_X1 U16892 ( .A1(n15249), .A2(n15248), .A3(n15247), .A4(n15246), .ZN(
        P2_U3227) );
  AOI22_X1 U16893 ( .A1(n15250), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(
        P2_REG3_REG_14__SCAN_IN), .B2(P2_U3088), .ZN(n15263) );
  OAI211_X1 U16894 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n15253), .A(n15252), 
        .B(n15251), .ZN(n15262) );
  OAI211_X1 U16895 ( .C1(n15257), .C2(n15256), .A(n15255), .B(n15254), .ZN(
        n15261) );
  NAND2_X1 U16896 ( .A1(n15259), .A2(n15258), .ZN(n15260) );
  NAND4_X1 U16897 ( .A1(n15263), .A2(n15262), .A3(n15261), .A4(n15260), .ZN(
        P2_U3228) );
  XNOR2_X1 U16898 ( .A(n15265), .B(n15264), .ZN(n15267) );
  AOI21_X1 U16899 ( .B1(n15267), .B2(n14065), .A(n15266), .ZN(n15307) );
  AOI222_X1 U16900 ( .A1(n15271), .A2(n15270), .B1(P2_REG2_REG_2__SCAN_IN), 
        .B2(n15269), .C1(n15268), .C2(P2_REG3_REG_2__SCAN_IN), .ZN(n15282) );
  XNOR2_X1 U16901 ( .A(n15273), .B(n15272), .ZN(n15311) );
  OAI21_X1 U16902 ( .B1(n15275), .B2(n15306), .A(n15274), .ZN(n15276) );
  OR2_X1 U16903 ( .A1(n15277), .A2(n15276), .ZN(n15305) );
  INV_X1 U16904 ( .A(n15305), .ZN(n15278) );
  AOI22_X1 U16905 ( .A1(n15311), .A2(n15280), .B1(n15279), .B2(n15278), .ZN(
        n15281) );
  OAI211_X1 U16906 ( .C1(n14078), .C2(n15307), .A(n15282), .B(n15281), .ZN(
        P2_U3263) );
  AND2_X1 U16907 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n15284), .ZN(P2_U3266) );
  AND2_X1 U16908 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n15284), .ZN(P2_U3267) );
  AND2_X1 U16909 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n15284), .ZN(P2_U3268) );
  AND2_X1 U16910 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n15284), .ZN(P2_U3269) );
  AND2_X1 U16911 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n15284), .ZN(P2_U3270) );
  AND2_X1 U16912 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n15284), .ZN(P2_U3271) );
  AND2_X1 U16913 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n15284), .ZN(P2_U3272) );
  AND2_X1 U16914 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n15284), .ZN(P2_U3273) );
  AND2_X1 U16915 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n15284), .ZN(P2_U3274) );
  AND2_X1 U16916 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n15284), .ZN(P2_U3275) );
  AND2_X1 U16917 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n15284), .ZN(P2_U3276) );
  AND2_X1 U16918 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n15284), .ZN(P2_U3277) );
  AND2_X1 U16919 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n15284), .ZN(P2_U3278) );
  AND2_X1 U16920 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n15284), .ZN(P2_U3279) );
  AND2_X1 U16921 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n15284), .ZN(P2_U3280) );
  AND2_X1 U16922 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n15284), .ZN(P2_U3281) );
  AND2_X1 U16923 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n15284), .ZN(P2_U3282) );
  AND2_X1 U16924 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n15284), .ZN(P2_U3283) );
  AND2_X1 U16925 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n15284), .ZN(P2_U3284) );
  AND2_X1 U16926 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n15284), .ZN(P2_U3285) );
  AND2_X1 U16927 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n15284), .ZN(P2_U3286) );
  AND2_X1 U16928 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n15284), .ZN(P2_U3287) );
  AND2_X1 U16929 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n15284), .ZN(P2_U3288) );
  AND2_X1 U16930 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n15284), .ZN(P2_U3289) );
  AND2_X1 U16931 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n15284), .ZN(P2_U3290) );
  AND2_X1 U16932 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n15284), .ZN(P2_U3291) );
  AND2_X1 U16933 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n15284), .ZN(P2_U3292) );
  AND2_X1 U16934 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n15284), .ZN(P2_U3293) );
  AND2_X1 U16935 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n15284), .ZN(P2_U3294) );
  AND2_X1 U16936 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n15284), .ZN(P2_U3295) );
  AOI22_X1 U16937 ( .A1(n15289), .A2(n15287), .B1(n15286), .B2(n15285), .ZN(
        P2_U3416) );
  OAI21_X1 U16938 ( .B1(n15290), .B2(n15289), .A(n15288), .ZN(P2_U3417) );
  INV_X1 U16939 ( .A(n15334), .ZN(n15345) );
  INV_X1 U16940 ( .A(n15291), .ZN(n15295) );
  INV_X1 U16941 ( .A(n15292), .ZN(n15294) );
  AOI211_X1 U16942 ( .C1(n15345), .C2(n15295), .A(n15294), .B(n15293), .ZN(
        n15349) );
  INV_X1 U16943 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n15296) );
  AOI22_X1 U16944 ( .A1(n15347), .A2(n15349), .B1(n15296), .B2(n15346), .ZN(
        P2_U3430) );
  INV_X1 U16945 ( .A(n15297), .ZN(n15303) );
  NOR2_X1 U16946 ( .A1(n15297), .A2(n15334), .ZN(n15302) );
  OAI211_X1 U16947 ( .C1(n15300), .C2(n15340), .A(n15299), .B(n15298), .ZN(
        n15301) );
  AOI211_X1 U16948 ( .C1(n15303), .C2(n15318), .A(n15302), .B(n15301), .ZN(
        n15350) );
  INV_X1 U16949 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n15304) );
  AOI22_X1 U16950 ( .A1(n15347), .A2(n15350), .B1(n15304), .B2(n15346), .ZN(
        P2_U3433) );
  OAI21_X1 U16951 ( .B1(n15306), .B2(n15340), .A(n15305), .ZN(n15309) );
  INV_X1 U16952 ( .A(n15307), .ZN(n15308) );
  AOI211_X1 U16953 ( .C1(n15311), .C2(n15310), .A(n15309), .B(n15308), .ZN(
        n15351) );
  INV_X1 U16954 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n15312) );
  AOI22_X1 U16955 ( .A1(n15347), .A2(n15351), .B1(n15312), .B2(n15346), .ZN(
        P2_U3436) );
  NAND2_X1 U16956 ( .A1(n15314), .A2(n15313), .ZN(n15315) );
  AND2_X1 U16957 ( .A1(n15316), .A2(n15315), .ZN(n15320) );
  OAI21_X1 U16958 ( .B1(n15318), .B2(n15345), .A(n15317), .ZN(n15319) );
  AND3_X1 U16959 ( .A1(n15321), .A2(n15320), .A3(n15319), .ZN(n15352) );
  AOI22_X1 U16960 ( .A1(n15347), .A2(n15352), .B1(n9132), .B2(n15346), .ZN(
        P2_U3439) );
  INV_X1 U16961 ( .A(n15322), .ZN(n15324) );
  OAI211_X1 U16962 ( .C1(n7049), .C2(n15340), .A(n15324), .B(n15323), .ZN(
        n15327) );
  AOI21_X1 U16963 ( .B1(n15335), .B2(n15334), .A(n15325), .ZN(n15326) );
  NOR2_X1 U16964 ( .A1(n15327), .A2(n15326), .ZN(n15353) );
  INV_X1 U16965 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n15328) );
  AOI22_X1 U16966 ( .A1(n15347), .A2(n15353), .B1(n15328), .B2(n15346), .ZN(
        P2_U3442) );
  INV_X1 U16967 ( .A(n15329), .ZN(n15331) );
  OAI211_X1 U16968 ( .C1(n15332), .C2(n15340), .A(n15331), .B(n15330), .ZN(
        n15337) );
  AOI21_X1 U16969 ( .B1(n15335), .B2(n15334), .A(n15333), .ZN(n15336) );
  NOR2_X1 U16970 ( .A1(n15337), .A2(n15336), .ZN(n15354) );
  INV_X1 U16971 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n15338) );
  AOI22_X1 U16972 ( .A1(n15347), .A2(n15354), .B1(n15338), .B2(n15346), .ZN(
        P2_U3445) );
  OAI21_X1 U16973 ( .B1(n15341), .B2(n15340), .A(n15339), .ZN(n15343) );
  AOI211_X1 U16974 ( .C1(n15345), .C2(n15344), .A(n15343), .B(n15342), .ZN(
        n15356) );
  AOI22_X1 U16975 ( .A1(n15347), .A2(n15356), .B1(n9279), .B2(n15346), .ZN(
        P2_U3460) );
  AOI22_X1 U16976 ( .A1(n15357), .A2(n15349), .B1(n15348), .B2(n15355), .ZN(
        P2_U3499) );
  AOI22_X1 U16977 ( .A1(n15357), .A2(n15350), .B1(n10075), .B2(n15355), .ZN(
        P2_U3500) );
  AOI22_X1 U16978 ( .A1(n15357), .A2(n15351), .B1(n10079), .B2(n15355), .ZN(
        P2_U3501) );
  AOI22_X1 U16979 ( .A1(n15357), .A2(n15352), .B1(n10074), .B2(n15355), .ZN(
        P2_U3502) );
  AOI22_X1 U16980 ( .A1(n15357), .A2(n15353), .B1(n10083), .B2(n15355), .ZN(
        P2_U3503) );
  AOI22_X1 U16981 ( .A1(n15357), .A2(n15354), .B1(n10084), .B2(n15355), .ZN(
        P2_U3504) );
  AOI22_X1 U16982 ( .A1(n15357), .A2(n15356), .B1(n10099), .B2(n15355), .ZN(
        P2_U3509) );
  NOR2_X1 U16983 ( .A1(P3_U3897), .A2(n15523), .ZN(P3_U3150) );
  OAI211_X1 U16984 ( .C1(n15360), .C2(n15359), .A(n15358), .B(n15390), .ZN(
        n15364) );
  NOR2_X1 U16985 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15361), .ZN(n15469) );
  AOI21_X1 U16986 ( .B1(n15362), .B2(n15393), .A(n15469), .ZN(n15363) );
  OAI211_X1 U16987 ( .C1(n15397), .C2(n15563), .A(n15364), .B(n15363), .ZN(
        n15365) );
  INV_X1 U16988 ( .A(n15365), .ZN(n15366) );
  OAI21_X1 U16989 ( .B1(n15367), .B2(n15401), .A(n15366), .ZN(P3_U3153) );
  OAI22_X1 U16990 ( .A1(n15370), .A2(n15369), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15368), .ZN(n15376) );
  INV_X1 U16991 ( .A(n15371), .ZN(n15372) );
  AOI211_X1 U16992 ( .C1(n15374), .C2(n15373), .A(n15381), .B(n15372), .ZN(
        n15375) );
  AOI211_X1 U16993 ( .C1(n15378), .C2(n15377), .A(n15376), .B(n15375), .ZN(
        n15379) );
  OAI21_X1 U16994 ( .B1(n15380), .B2(n15401), .A(n15379), .ZN(P3_U3157) );
  AOI21_X1 U16995 ( .B1(n15383), .B2(n15382), .A(n15381), .ZN(n15388) );
  AOI22_X1 U16996 ( .A1(n15384), .A2(n15393), .B1(P3_REG3_REG_3__SCAN_IN), 
        .B2(P3_U3151), .ZN(n15385) );
  OAI21_X1 U16997 ( .B1(n15397), .B2(n15539), .A(n15385), .ZN(n15386) );
  AOI21_X1 U16998 ( .B1(n15388), .B2(n15387), .A(n15386), .ZN(n15389) );
  OAI21_X1 U16999 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(n15401), .A(n15389), .ZN(
        P3_U3158) );
  OAI211_X1 U17000 ( .C1(n6797), .C2(n15392), .A(n15391), .B(n15390), .ZN(
        n15396) );
  AOI22_X1 U17001 ( .A1(n15394), .A2(n15393), .B1(P3_REG3_REG_6__SCAN_IN), 
        .B2(P3_U3151), .ZN(n15395) );
  OAI211_X1 U17002 ( .C1(n15398), .C2(n15397), .A(n15396), .B(n15395), .ZN(
        n15399) );
  INV_X1 U17003 ( .A(n15399), .ZN(n15400) );
  OAI21_X1 U17004 ( .B1(n15402), .B2(n15401), .A(n15400), .ZN(P3_U3179) );
  INV_X1 U17005 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n15421) );
  AOI21_X1 U17006 ( .B1(n15405), .B2(n15404), .A(n15403), .ZN(n15410) );
  AOI21_X1 U17007 ( .B1(n15406), .B2(n15408), .A(n15407), .ZN(n15409) );
  OAI22_X1 U17008 ( .A1(n15410), .A2(n15530), .B1(n15516), .B2(n15409), .ZN(
        n15411) );
  INV_X1 U17009 ( .A(n15411), .ZN(n15416) );
  XNOR2_X1 U17010 ( .A(n15413), .B(n15412), .ZN(n15414) );
  NAND2_X1 U17011 ( .A1(n15414), .A2(n15504), .ZN(n15415) );
  OAI211_X1 U17012 ( .C1(n15520), .C2(n15417), .A(n15416), .B(n15415), .ZN(
        n15418) );
  INV_X1 U17013 ( .A(n15418), .ZN(n15420) );
  NAND2_X1 U17014 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_U3151), .ZN(n15419) );
  OAI211_X1 U17015 ( .C1(n15421), .C2(n15492), .A(n15420), .B(n15419), .ZN(
        P3_U3186) );
  AOI21_X1 U17016 ( .B1(n15424), .B2(n15423), .A(n15422), .ZN(n15428) );
  AOI21_X1 U17017 ( .B1(n15596), .B2(n15426), .A(n15425), .ZN(n15427) );
  OAI22_X1 U17018 ( .A1(n15428), .A2(n15530), .B1(n15516), .B2(n15427), .ZN(
        n15433) );
  XOR2_X1 U17019 ( .A(n15429), .B(n15430), .Z(n15431) );
  NOR2_X1 U17020 ( .A1(n15431), .A2(n7858), .ZN(n15432) );
  AOI211_X1 U17021 ( .C1(n15485), .C2(n15434), .A(n15433), .B(n15432), .ZN(
        n15436) );
  NAND2_X1 U17022 ( .A1(P3_REG3_REG_5__SCAN_IN), .A2(P3_U3151), .ZN(n15435) );
  OAI211_X1 U17023 ( .C1(n7868), .C2(n15492), .A(n15436), .B(n15435), .ZN(
        P3_U3187) );
  XNOR2_X1 U17024 ( .A(n15438), .B(n15437), .ZN(n15450) );
  AOI21_X1 U17025 ( .B1(n15441), .B2(n15440), .A(n15439), .ZN(n15443) );
  OAI22_X1 U17026 ( .A1(n15443), .A2(n15516), .B1(n15442), .B2(n15520), .ZN(
        n15449) );
  AOI21_X1 U17027 ( .B1(n15446), .B2(n15445), .A(n15444), .ZN(n15447) );
  NOR2_X1 U17028 ( .A1(n15447), .A2(n15530), .ZN(n15448) );
  AOI211_X1 U17029 ( .C1(n15504), .C2(n15450), .A(n15449), .B(n15448), .ZN(
        n15452) );
  NAND2_X1 U17030 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n15451) );
  OAI211_X1 U17031 ( .C1(n15453), .C2(n15492), .A(n15452), .B(n15451), .ZN(
        P3_U3188) );
  AOI21_X1 U17032 ( .B1(n15456), .B2(n15455), .A(n15454), .ZN(n15457) );
  OR2_X1 U17033 ( .A1(n15457), .A2(n15530), .ZN(n15468) );
  XNOR2_X1 U17034 ( .A(n15459), .B(n15458), .ZN(n15460) );
  NAND2_X1 U17035 ( .A1(n15460), .A2(n15504), .ZN(n15467) );
  AOI21_X1 U17036 ( .B1(n15600), .B2(n15462), .A(n15461), .ZN(n15463) );
  OR2_X1 U17037 ( .A1(n15463), .A2(n15516), .ZN(n15466) );
  NAND2_X1 U17038 ( .A1(n15485), .A2(n15464), .ZN(n15465) );
  AND4_X1 U17039 ( .A1(n15468), .A2(n15467), .A3(n15466), .A4(n15465), .ZN(
        n15471) );
  INV_X1 U17040 ( .A(n15469), .ZN(n15470) );
  OAI211_X1 U17041 ( .C1(n15472), .C2(n15492), .A(n15471), .B(n15470), .ZN(
        P3_U3189) );
  AOI21_X1 U17042 ( .B1(n15475), .B2(n15474), .A(n15473), .ZN(n15476) );
  OR2_X1 U17043 ( .A1(n15476), .A2(n15530), .ZN(n15489) );
  XNOR2_X1 U17044 ( .A(n15478), .B(n15477), .ZN(n15479) );
  NAND2_X1 U17045 ( .A1(n15479), .A2(n15504), .ZN(n15488) );
  AOI21_X1 U17046 ( .B1(n6793), .B2(n15481), .A(n15480), .ZN(n15482) );
  OR2_X1 U17047 ( .A1(n15482), .A2(n15516), .ZN(n15487) );
  INV_X1 U17048 ( .A(n15483), .ZN(n15484) );
  NAND2_X1 U17049 ( .A1(n15485), .A2(n15484), .ZN(n15486) );
  AND4_X1 U17050 ( .A1(n15489), .A2(n15488), .A3(n15487), .A4(n15486), .ZN(
        n15491) );
  OAI211_X1 U17051 ( .C1(n15493), .C2(n15492), .A(n15491), .B(n15490), .ZN(
        P3_U3190) );
  AOI21_X1 U17052 ( .B1(n6780), .B2(n15495), .A(n15494), .ZN(n15509) );
  AOI21_X1 U17053 ( .B1(n6779), .B2(n15497), .A(n15496), .ZN(n15498) );
  NOR2_X1 U17054 ( .A1(n15498), .A2(n15516), .ZN(n15502) );
  OAI21_X1 U17055 ( .B1(n15520), .B2(n15500), .A(n15499), .ZN(n15501) );
  AOI211_X1 U17056 ( .C1(P3_ADDR_REG_12__SCAN_IN), .C2(n15523), .A(n15502), 
        .B(n15501), .ZN(n15508) );
  OAI211_X1 U17057 ( .C1(n15506), .C2(n15505), .A(n15504), .B(n15503), .ZN(
        n15507) );
  OAI211_X1 U17058 ( .C1(n15509), .C2(n15530), .A(n15508), .B(n15507), .ZN(
        P3_U3194) );
  AOI21_X1 U17059 ( .B1(n15512), .B2(n15511), .A(n15510), .ZN(n15531) );
  AOI21_X1 U17060 ( .B1(n15515), .B2(n15514), .A(n15513), .ZN(n15517) );
  NOR2_X1 U17061 ( .A1(n15517), .A2(n15516), .ZN(n15522) );
  OAI21_X1 U17062 ( .B1(n15520), .B2(n15519), .A(n15518), .ZN(n15521) );
  AOI211_X1 U17063 ( .C1(P3_ADDR_REG_14__SCAN_IN), .C2(n15523), .A(n15522), 
        .B(n15521), .ZN(n15529) );
  AOI211_X1 U17064 ( .C1(n15526), .C2(n15525), .A(n15524), .B(n7858), .ZN(
        n15527) );
  INV_X1 U17065 ( .A(n15527), .ZN(n15528) );
  OAI211_X1 U17066 ( .C1(n15531), .C2(n15530), .A(n15529), .B(n15528), .ZN(
        P3_U3196) );
  INV_X1 U17067 ( .A(n15532), .ZN(n15534) );
  AOI211_X1 U17068 ( .C1(n15535), .C2(n15578), .A(n15534), .B(n15533), .ZN(
        n15592) );
  INV_X1 U17069 ( .A(P3_REG0_REG_2__SCAN_IN), .ZN(n15536) );
  AOI22_X1 U17070 ( .A1(n15591), .A2(n15592), .B1(n15536), .B2(n15589), .ZN(
        P3_U3396) );
  NAND2_X1 U17071 ( .A1(n15541), .A2(n15578), .ZN(n15537) );
  OAI211_X1 U17072 ( .C1(n15539), .C2(n15582), .A(n15538), .B(n15537), .ZN(
        n15540) );
  AOI21_X1 U17073 ( .B1(n15541), .B2(n15588), .A(n15540), .ZN(n15593) );
  INV_X1 U17074 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n15542) );
  AOI22_X1 U17075 ( .A1(n15591), .A2(n15593), .B1(n15542), .B2(n15589), .ZN(
        P3_U3399) );
  INV_X1 U17076 ( .A(n15543), .ZN(n15544) );
  OAI21_X1 U17077 ( .B1(n15578), .B2(n15588), .A(n15544), .ZN(n15547) );
  NAND2_X1 U17078 ( .A1(n15545), .A2(n15561), .ZN(n15546) );
  AND3_X1 U17079 ( .A1(n15548), .A2(n15547), .A3(n15546), .ZN(n15595) );
  INV_X1 U17080 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n15549) );
  AOI22_X1 U17081 ( .A1(n15591), .A2(n15595), .B1(n15549), .B2(n15589), .ZN(
        P3_U3402) );
  NOR2_X1 U17082 ( .A1(n15550), .A2(n15582), .ZN(n15552) );
  AOI211_X1 U17083 ( .C1(n15553), .C2(n15578), .A(n15552), .B(n15551), .ZN(
        n15597) );
  INV_X1 U17084 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n15554) );
  AOI22_X1 U17085 ( .A1(n15591), .A2(n15597), .B1(n15554), .B2(n15589), .ZN(
        P3_U3405) );
  INV_X1 U17086 ( .A(n15555), .ZN(n15559) );
  AOI21_X1 U17087 ( .B1(n15557), .B2(n15583), .A(n15556), .ZN(n15558) );
  AOI211_X1 U17088 ( .C1(n15561), .C2(n15560), .A(n15559), .B(n15558), .ZN(
        n15599) );
  INV_X1 U17089 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15562) );
  AOI22_X1 U17090 ( .A1(n15591), .A2(n15599), .B1(n15562), .B2(n15589), .ZN(
        P3_U3408) );
  INV_X1 U17091 ( .A(n15564), .ZN(n15567) );
  OAI22_X1 U17092 ( .A1(n15564), .A2(n15583), .B1(n15582), .B2(n15563), .ZN(
        n15566) );
  AOI211_X1 U17093 ( .C1(n15567), .C2(n15588), .A(n15566), .B(n15565), .ZN(
        n15601) );
  INV_X1 U17094 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15568) );
  AOI22_X1 U17095 ( .A1(n15591), .A2(n15601), .B1(n15568), .B2(n15589), .ZN(
        P3_U3411) );
  OAI22_X1 U17096 ( .A1(n15571), .A2(n15570), .B1(n15569), .B2(n15582), .ZN(
        n15572) );
  NOR2_X1 U17097 ( .A1(n15573), .A2(n15572), .ZN(n15603) );
  INV_X1 U17098 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15574) );
  AOI22_X1 U17099 ( .A1(n15591), .A2(n15603), .B1(n15574), .B2(n15589), .ZN(
        P3_U3414) );
  NOR2_X1 U17100 ( .A1(n15575), .A2(n15582), .ZN(n15577) );
  AOI211_X1 U17101 ( .C1(n15579), .C2(n15578), .A(n15577), .B(n15576), .ZN(
        n15605) );
  INV_X1 U17102 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15580) );
  AOI22_X1 U17103 ( .A1(n15591), .A2(n15605), .B1(n15580), .B2(n15589), .ZN(
        P3_U3417) );
  INV_X1 U17104 ( .A(n15584), .ZN(n15587) );
  OAI22_X1 U17105 ( .A1(n15584), .A2(n15583), .B1(n15582), .B2(n15581), .ZN(
        n15586) );
  AOI211_X1 U17106 ( .C1(n15588), .C2(n15587), .A(n15586), .B(n15585), .ZN(
        n15606) );
  INV_X1 U17107 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15590) );
  AOI22_X1 U17108 ( .A1(n15591), .A2(n15606), .B1(n15590), .B2(n15589), .ZN(
        P3_U3420) );
  AOI22_X1 U17109 ( .A1(n15607), .A2(n15592), .B1(n7767), .B2(n9022), .ZN(
        P3_U3461) );
  AOI22_X1 U17110 ( .A1(n15607), .A2(n15593), .B1(n7519), .B2(n9022), .ZN(
        P3_U3462) );
  INV_X1 U17111 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n15594) );
  AOI22_X1 U17112 ( .A1(n15607), .A2(n15595), .B1(n15594), .B2(n9022), .ZN(
        P3_U3463) );
  AOI22_X1 U17113 ( .A1(n15607), .A2(n15597), .B1(n15596), .B2(n9022), .ZN(
        P3_U3464) );
  INV_X1 U17114 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15598) );
  AOI22_X1 U17115 ( .A1(n15607), .A2(n15599), .B1(n15598), .B2(n9022), .ZN(
        P3_U3465) );
  AOI22_X1 U17116 ( .A1(n15607), .A2(n15601), .B1(n15600), .B2(n9022), .ZN(
        P3_U3466) );
  INV_X1 U17117 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15602) );
  AOI22_X1 U17118 ( .A1(n15607), .A2(n15603), .B1(n15602), .B2(n9022), .ZN(
        P3_U3467) );
  AOI22_X1 U17119 ( .A1(n15607), .A2(n15605), .B1(n15604), .B2(n9022), .ZN(
        P3_U3468) );
  AOI22_X1 U17120 ( .A1(n15607), .A2(n15606), .B1(n7790), .B2(n9022), .ZN(
        P3_U3469) );
  AOI21_X1 U17121 ( .B1(n15610), .B2(n15609), .A(n15608), .ZN(SUB_1596_U59) );
  OAI21_X1 U17122 ( .B1(n15613), .B2(n15612), .A(n15611), .ZN(SUB_1596_U58) );
  XOR2_X1 U17123 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(n15614), .Z(SUB_1596_U53) );
  OAI21_X1 U17124 ( .B1(n15617), .B2(n15616), .A(n15615), .ZN(SUB_1596_U56) );
  OAI21_X1 U17125 ( .B1(n15620), .B2(n15619), .A(n15618), .ZN(n15621) );
  XNOR2_X1 U17126 ( .A(n15621), .B(P2_ADDR_REG_3__SCAN_IN), .ZN(SUB_1596_U60)
         );
  AOI21_X1 U17127 ( .B1(n15624), .B2(n15623), .A(n15622), .ZN(SUB_1596_U5) );
  BUF_X2 U7418 ( .A(n10832), .Z(n12670) );
  CLKBUF_X2 U7419 ( .A(n10989), .Z(n12664) );
  OAI21_X1 U7521 ( .B1(n8775), .B2(n7102), .A(P3_IR_REG_31__SCAN_IN), .ZN(
        n7753) );
  NAND2_X2 U7525 ( .A1(n15274), .A2(n9758), .ZN(n10734) );
  CLKBUF_X2 U7630 ( .A(n8361), .Z(n6879) );
  CLKBUF_X1 U9461 ( .A(n9105), .Z(n9523) );
  NOR2_X2 U9499 ( .A1(n10495), .A2(n10028), .ZN(n10029) );
endmodule

