

module b20_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, 
        SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, 
        SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, 
        SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_, 
        P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN, 
        P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN, 
        P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN, 
        P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN, 
        P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN, 
        P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN, 
        P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN, 
        P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN, 
        P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN, 
        P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, 
        P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, 
        P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, 
        P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, 
        P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, 
        P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, 
        P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, 
        P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, 
        P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, 
        P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, 
        P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, 
        P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, 
        P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, 
        P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, 
        P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, 
        P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, 
        P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, 
        P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, 
        P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, 
        P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, 
        P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, 
        P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, 
        P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, 
        P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, 
        P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, 
        P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN, 
        P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN, 
        P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN, 
        P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN, 
        P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN, 
        P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN, 
        P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN, 
        P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN, 
        P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN, 
        P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN, 
        P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN, 
        P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN, 
        P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN, 
        P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN, 
        P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN, 
        P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN, 
        P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN, 
        P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN, 
        P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN, 
        P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN, 
        P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN, 
        P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN, 
        P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN, 
        P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN, 
        P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN, 
        P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN, 
        P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, 
        P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, 
        P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, 
        P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN, 
        P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN, 
        P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN, 
        P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN, 
        P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN, 
        P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN, 
        P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN, 
        P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN, 
        P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN, 
        P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN, 
        P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN, 
        P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN, 
        P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN, 
        P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN, 
        P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN, 
        P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN, 
        P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN, 
        P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN, 
        P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN, 
        P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, 
        P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN, 
        P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN, 
        P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN, 
        P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN, 
        P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN, 
        P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, ADD_1068_U4, 
        ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58, ADD_1068_U59, 
        ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63, ADD_1068_U47, 
        ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51, ADD_1068_U52, 
        ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46, U126, U123, 
        P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, 
        P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, 
        P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, 
        P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, 
        P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440, P1_U3323, 
        P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, 
        P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, 
        P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, 
        P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, 
        P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465, P1_U3468, 
        P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, 
        P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3509, 
        P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516, 
        P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, 
        P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, 
        P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, 
        P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, 
        P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, 
        P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290, P1_U3289, 
        P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, 
        P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, 
        P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, 
        P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263, P1_U3262, 
        P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, 
        P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, 
        P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554, P1_U3555, 
        P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562, 
        P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, 
        P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, 
        P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, 
        P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239, P1_U3238, 
        P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, 
        P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, 
        P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, 
        P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085, P1_U3973, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377, P2_U3263, 
        P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, 
        P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, 
        P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, 
        P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, 
        P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402, P2_U3405, 
        P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423, P2_U3426, 
        P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444, P2_U3446, 
        P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452, P2_U3453, 
        P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459, P2_U3460, 
        P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466, P2_U3467, 
        P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473, P2_U3474, 
        P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480, P2_U3481, 
        P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487, P2_U3488, 
        P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, 
        P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, 
        P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, 
        P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491, P2_U3492, 
        P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499, 
        P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506, 
        P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513, 
        P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520, 
        P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179, P2_U3178, 
        P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, 
        P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, 
        P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, 
        P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150, P2_U3893
 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
         ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
         ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
         ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
         U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351,
         P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344,
         P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337,
         P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330,
         P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439,
         P1_U3440, P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318,
         P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311,
         P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304,
         P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297,
         P1_U3296, P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462,
         P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483,
         P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504,
         P1_U3507, P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291,
         P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284,
         P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277,
         P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270,
         P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264,
         P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257,
         P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250,
         P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243,
         P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240,
         P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233,
         P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226,
         P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219,
         P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086,
         P1_U3085, P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291,
         P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284,
         P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277,
         P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270,
         P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376,
         P2_U3377, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
         P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
         P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244,
         P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237,
         P2_U3236, P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399,
         P2_U3402, P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420,
         P2_U3423, P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441,
         P2_U3444, P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451,
         P2_U3452, P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458,
         P2_U3459, P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465,
         P2_U3466, P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472,
         P2_U3473, P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479,
         P2_U3480, P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486,
         P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231,
         P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224,
         P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217,
         P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210,
         P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203,
         P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196,
         P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189,
         P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182,
         P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497,
         P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504,
         P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511,
         P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518,
         P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180,
         P2_U3179, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173,
         P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166,
         P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159,
         P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151,
         P2_U3150, P2_U3893;
  wire   n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211,
         n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221,
         n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231,
         n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241,
         n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251,
         n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261,
         n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271,
         n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281,
         n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291,
         n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301,
         n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311,
         n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321,
         n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331,
         n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341,
         n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351,
         n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
         n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
         n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381,
         n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391,
         n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401,
         n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411,
         n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421,
         n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431,
         n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441,
         n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451,
         n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461,
         n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
         n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
         n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
         n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
         n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
         n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
         n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531,
         n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541,
         n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551,
         n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
         n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571,
         n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581,
         n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
         n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
         n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
         n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
         n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
         n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
         n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
         n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
         n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
         n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
         n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
         n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701,
         n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711,
         n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721,
         n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731,
         n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741,
         n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781,
         n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791,
         n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801,
         n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811,
         n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821,
         n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831,
         n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841,
         n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851,
         n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861,
         n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871,
         n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881,
         n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891,
         n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
         n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
         n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
         n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
         n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941,
         n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951,
         n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961,
         n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971,
         n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981,
         n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991,
         n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
         n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011,
         n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
         n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031,
         n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041,
         n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051,
         n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061,
         n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071,
         n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081,
         n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091,
         n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101,
         n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111,
         n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121,
         n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141,
         n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151,
         n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161,
         n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
         n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191,
         n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201,
         n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211,
         n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221,
         n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231,
         n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241,
         n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251,
         n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261,
         n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271,
         n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281,
         n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291,
         n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301,
         n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311,
         n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321,
         n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331,
         n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341,
         n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351,
         n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361,
         n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371,
         n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381,
         n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391,
         n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401,
         n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411,
         n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421,
         n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431,
         n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441,
         n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
         n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471,
         n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481,
         n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491,
         n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501,
         n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
         n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521,
         n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531,
         n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541,
         n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551,
         n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561,
         n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571,
         n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581,
         n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591,
         n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601,
         n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611,
         n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621,
         n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631,
         n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641,
         n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651,
         n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661,
         n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671,
         n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681,
         n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701,
         n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711,
         n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721,
         n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731,
         n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751,
         n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761,
         n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
         n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781,
         n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791,
         n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801,
         n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811,
         n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821,
         n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831,
         n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841,
         n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851,
         n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861,
         n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871,
         n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881,
         n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891,
         n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901,
         n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
         n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921,
         n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931,
         n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941,
         n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951,
         n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961,
         n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971,
         n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981,
         n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991,
         n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001,
         n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011,
         n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021,
         n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031,
         n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041,
         n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051,
         n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061,
         n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071,
         n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081,
         n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091,
         n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101,
         n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111,
         n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121,
         n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131,
         n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141,
         n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151,
         n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161,
         n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171,
         n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181,
         n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191,
         n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201,
         n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211,
         n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221,
         n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231,
         n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241,
         n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251,
         n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261,
         n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271,
         n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281,
         n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291,
         n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301,
         n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311,
         n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321,
         n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331,
         n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341,
         n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351,
         n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361,
         n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371,
         n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381,
         n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391,
         n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401,
         n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411,
         n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421,
         n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431,
         n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441,
         n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
         n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461,
         n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471,
         n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
         n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
         n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
         n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
         n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
         n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
         n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
         n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
         n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
         n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
         n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
         n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
         n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
         n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
         n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
         n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
         n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
         n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
         n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
         n9672, n9673, n9674, n9675, n9676, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11212;

  INV_X4 U5194 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  AOI21_X1 U5195 ( .B1(n6090), .B2(n5814), .A(n5728), .ZN(n6100) );
  BUF_X1 U5196 ( .A(n8389), .Z(n5144) );
  INV_X1 U5197 ( .A(n5891), .ZN(n5914) );
  BUF_X2 U5198 ( .A(n5915), .Z(n7377) );
  AND3_X1 U5199 ( .A1(n6964), .A2(n6963), .A3(n6962), .ZN(n11023) );
  OR2_X4 U5200 ( .A1(n6522), .A2(n6520), .ZN(n6968) );
  XNOR2_X1 U5201 ( .A(n6784), .B(P1_IR_REG_19__SCAN_IN), .ZN(n10158) );
  INV_X1 U5203 ( .A(n11212), .ZN(n5131) );
  INV_X1 U5204 ( .A(n8676), .ZN(n8663) );
  INV_X1 U5205 ( .A(n8330), .ZN(n8388) );
  NOR2_X1 U5206 ( .A1(n5622), .A2(n6889), .ZN(n6892) );
  INV_X1 U5207 ( .A(n8389), .ZN(n8264) );
  OR2_X1 U5208 ( .A1(n6996), .A2(n6997), .ZN(n7014) );
  INV_X2 U5209 ( .A(n7325), .ZN(n8387) );
  CLKBUF_X3 U5210 ( .A(n6949), .Z(n8346) );
  NAND2_X2 U5213 ( .A1(n5912), .A2(n6884), .ZN(n5926) );
  NAND2_X1 U5214 ( .A1(n8673), .A2(n8962), .ZN(n7119) );
  OR2_X1 U5215 ( .A1(n9252), .A2(n9253), .ZN(n5757) );
  NAND2_X1 U5216 ( .A1(n7460), .A2(n7459), .ZN(n7681) );
  NAND2_X1 U5217 ( .A1(n5633), .A2(n5631), .ZN(n7866) );
  INV_X1 U5218 ( .A(n8390), .ZN(n8349) );
  AND2_X1 U5219 ( .A1(n7675), .A2(n10158), .ZN(n9663) );
  AND3_X1 U5220 ( .A1(n7003), .A2(n7002), .A3(n7001), .ZN(n7394) );
  INV_X1 U5221 ( .A(n9409), .ZN(n10983) );
  OAI21_X2 U5222 ( .B1(n6461), .B2(P1_IR_REG_21__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6537) );
  AND2_X1 U5223 ( .A1(n6279), .A2(n6278), .ZN(n9015) );
  AOI21_X1 U5224 ( .B1(n8292), .B2(n8468), .A(n6223), .ZN(n9174) );
  NAND2_X1 U5225 ( .A1(n6003), .A2(n6002), .ZN(n7628) );
  OAI21_X1 U5226 ( .B1(n9301), .B2(n5628), .A(n5626), .ZN(n5629) );
  INV_X1 U5227 ( .A(n6959), .ZN(n8029) );
  NAND2_X1 U5228 ( .A1(n9623), .A2(n10185), .ZN(n10262) );
  NAND4_X1 U5229 ( .A1(n5920), .A2(n5919), .A3(n5918), .A4(n5917), .ZN(n8843)
         );
  BUF_X1 U5230 ( .A(n8525), .Z(n5140) );
  INV_X2 U5232 ( .A(n8387), .ZN(n8390) );
  NAND2_X1 U5233 ( .A1(n6787), .A2(n10522), .ZN(n5132) );
  NAND2_X1 U5234 ( .A1(n6787), .A2(n10522), .ZN(n5133) );
  NAND2_X1 U5235 ( .A1(n6787), .A2(n10522), .ZN(n7322) );
  NAND2_X2 U5236 ( .A1(n6329), .A2(n8585), .ZN(n7817) );
  OAI21_X2 U5237 ( .B1(n7590), .B2(n7585), .A(n6033), .ZN(n7730) );
  NAND2_X1 U5238 ( .A1(n6783), .A2(n6460), .ZN(n6461) );
  OAI21_X2 U5239 ( .B1(n6174), .B2(P2_IR_REG_18__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6293) );
  XNOR2_X2 U5240 ( .A(n6347), .B(n6346), .ZN(n6354) );
  AOI21_X2 U5241 ( .B1(P1_REG1_REG_14__SCAN_IN), .B2(n10699), .A(n10701), .ZN(
        n10114) );
  OAI21_X2 U5242 ( .B1(n7960), .B2(n5471), .A(n5469), .ZN(n9139) );
  BUF_X4 U5243 ( .A(n5872), .Z(n5134) );
  NAND2_X1 U5244 ( .A1(n5323), .A2(n5324), .ZN(n5872) );
  XNOR2_X2 U5245 ( .A(n8844), .B(n8539), .ZN(n8541) );
  BUF_X1 U5246 ( .A(n5889), .Z(n5135) );
  BUF_X2 U5247 ( .A(n5889), .Z(n5137) );
  INV_X1 U5248 ( .A(n5916), .ZN(n5889) );
  NAND2_X1 U5250 ( .A1(n6808), .A2(n6807), .ZN(n5622) );
  NAND2_X1 U5251 ( .A1(n5132), .A2(n5134), .ZN(n5138) );
  NAND2_X1 U5252 ( .A1(n5132), .A2(n5134), .ZN(n5139) );
  OAI21_X4 U5253 ( .B1(n9068), .B2(n8472), .A(n8642), .ZN(n9056) );
  OAI21_X2 U5254 ( .B1(n9094), .B2(n5465), .A(n5462), .ZN(n9068) );
  AOI22_X2 U5255 ( .A1(n9678), .A2(n9679), .B1(n7525), .B2(
        P1_REG1_REG_10__SCAN_IN), .ZN(n10684) );
  NAND4_X2 U5256 ( .A1(n5174), .A2(n6900), .A3(n6899), .A4(n6898), .ZN(n11020)
         );
  XNOR2_X1 U5257 ( .A(n6296), .B(n6295), .ZN(n8525) );
  OR2_X4 U5258 ( .A1(n6800), .A2(n6799), .ZN(n7325) );
  AOI22_X2 U5259 ( .A1(n10371), .A2(n10370), .B1(n10364), .B2(n10483), .ZN(
        n10353) );
  OAI22_X2 U5260 ( .A1(n10192), .A2(n10191), .B1(n10190), .B2(n10378), .ZN(
        n10371) );
  NAND2_X1 U5261 ( .A1(n7975), .A2(n7974), .ZN(n8058) );
  AOI21_X1 U5262 ( .B1(n7197), .B2(n7179), .A(n5731), .ZN(n7270) );
  NAND2_X1 U5263 ( .A1(n6933), .A2(n5898), .ZN(n6923) );
  INV_X1 U5264 ( .A(n8843), .ZN(n7137) );
  INV_X1 U5265 ( .A(n8842), .ZN(n7047) );
  INV_X1 U5266 ( .A(n8838), .ZN(n7570) );
  INV_X1 U5267 ( .A(n8837), .ZN(n7510) );
  INV_X1 U5268 ( .A(n6730), .ZN(n8539) );
  INV_X2 U5270 ( .A(n6949), .ZN(n8314) );
  INV_X4 U5271 ( .A(n5134), .ZN(n6884) );
  OAI21_X1 U5272 ( .B1(n9271), .B2(n5171), .A(n9376), .ZN(n9276) );
  AND2_X1 U5273 ( .A1(n6438), .A2(n7448), .ZN(n6439) );
  AOI21_X1 U5274 ( .B1(n10404), .B2(n11181), .A(n5333), .ZN(n10405) );
  OR2_X1 U5275 ( .A1(n10414), .A2(n11104), .ZN(n5288) );
  OAI21_X1 U5276 ( .B1(n8510), .B2(n8509), .A(n5732), .ZN(n8511) );
  NAND2_X1 U5277 ( .A1(n10235), .A2(n10187), .ZN(n10218) );
  AND2_X1 U5278 ( .A1(n5508), .A2(n5181), .ZN(n6404) );
  NAND2_X1 U5279 ( .A1(n10284), .A2(n10283), .ZN(n10282) );
  AND2_X1 U5280 ( .A1(n10222), .A2(n10221), .ZN(n10407) );
  NOR2_X1 U5281 ( .A1(n10305), .A2(n5343), .ZN(n5338) );
  NAND2_X1 U5282 ( .A1(n10234), .A2(n10199), .ZN(n5722) );
  OR2_X1 U5283 ( .A1(n10403), .A2(n10402), .ZN(n5333) );
  AOI21_X1 U5284 ( .B1(n5723), .B2(n5627), .A(n8374), .ZN(n5626) );
  INV_X1 U5285 ( .A(n5723), .ZN(n5628) );
  NOR2_X1 U5286 ( .A1(n9089), .A2(n9093), .ZN(n5402) );
  NAND2_X1 U5287 ( .A1(n5290), .A2(n10184), .ZN(n5537) );
  NAND2_X1 U5288 ( .A1(n8058), .A2(n5725), .ZN(n8171) );
  OAI22_X1 U5289 ( .A1(n10194), .A2(n5707), .B1(n10306), .B2(n10463), .ZN(
        n5706) );
  AOI21_X2 U5290 ( .B1(n8319), .B2(n8029), .A(n5239), .ZN(n10435) );
  NAND2_X1 U5291 ( .A1(n7799), .A2(n7798), .ZN(n7986) );
  NAND2_X1 U5292 ( .A1(n7758), .A2(n7757), .ZN(n7799) );
  OR2_X1 U5293 ( .A1(n10382), .A2(n10483), .ZN(n10379) );
  NAND2_X1 U5294 ( .A1(n6202), .A2(n6201), .ZN(n9179) );
  NAND2_X1 U5295 ( .A1(n6220), .A2(n6219), .ZN(n6222) );
  NOR2_X1 U5296 ( .A1(n7791), .A2(n5325), .ZN(n7792) );
  NAND2_X1 U5297 ( .A1(n8032), .A2(n8031), .ZN(n9400) );
  NAND2_X1 U5298 ( .A1(n7989), .A2(n7988), .ZN(n8121) );
  NAND2_X1 U5299 ( .A1(n6103), .A2(n6102), .ZN(n8115) );
  NAND2_X1 U5300 ( .A1(n5284), .A2(n5283), .ZN(n6126) );
  NAND2_X1 U5301 ( .A1(n6074), .A2(n6073), .ZN(n7908) );
  NAND2_X1 U5302 ( .A1(n7527), .A2(n7526), .ZN(n11148) );
  NAND2_X2 U5303 ( .A1(n7134), .A2(n8545), .ZN(n7133) );
  INV_X1 U5304 ( .A(n9554), .ZN(n11062) );
  INV_X2 U5305 ( .A(n9145), .ZN(n9150) );
  NAND2_X1 U5306 ( .A1(n6021), .A2(n6020), .ZN(n7664) );
  XNOR2_X1 U5307 ( .A(n5396), .B(n5997), .ZN(n7539) );
  NAND2_X1 U5308 ( .A1(n5990), .A2(n5257), .ZN(n7400) );
  AND2_X1 U5309 ( .A1(n9543), .A2(n9541), .ZN(n7269) );
  NAND2_X1 U5310 ( .A1(n5897), .A2(n6682), .ZN(n8537) );
  AND3_X1 U5311 ( .A1(n6947), .A2(n6946), .A3(n6945), .ZN(n11010) );
  NAND4_X2 U5312 ( .A1(n6767), .A2(n6766), .A3(n6765), .A4(n6764), .ZN(n11007)
         );
  NAND4_X1 U5313 ( .A1(n5941), .A2(n5940), .A3(n5939), .A4(n5938), .ZN(n8842)
         );
  CLKBUF_X3 U5314 ( .A(n6752), .Z(n8440) );
  NAND4_X1 U5315 ( .A1(n6987), .A2(n6986), .A3(n6985), .A4(n6984), .ZN(n11019)
         );
  NAND2_X1 U5316 ( .A1(n5914), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5902) );
  CLKBUF_X1 U5317 ( .A(n6426), .Z(n7372) );
  AND4_X1 U5318 ( .A1(n5895), .A2(n5894), .A3(n5893), .A4(n5892), .ZN(n8168)
         );
  NAND2_X1 U5319 ( .A1(n6426), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5901) );
  OAI211_X1 U5320 ( .C1(n5912), .C2(n6613), .A(n5911), .B(n5910), .ZN(n6730)
         );
  NAND2_X1 U5321 ( .A1(n8699), .A2(n5762), .ZN(n5891) );
  CLKBUF_X1 U5322 ( .A(n6800), .Z(n6806) );
  OR2_X2 U5323 ( .A1(n6800), .A2(n6791), .ZN(n6949) );
  OAI211_X1 U5325 ( .C1(n5926), .C2(n5769), .A(n5881), .B(n5724), .ZN(n6682)
         );
  NAND2_X1 U5326 ( .A1(n5761), .A2(n5762), .ZN(n5916) );
  CLKBUF_X1 U5327 ( .A(n5909), .Z(n6070) );
  NAND2_X1 U5328 ( .A1(n10508), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5550) );
  NAND2_X1 U5329 ( .A1(n9655), .A2(n9663), .ZN(n10995) );
  INV_X1 U5331 ( .A(n9260), .ZN(n5762) );
  XNOR2_X1 U5332 ( .A(n5760), .B(n5759), .ZN(n9260) );
  XNOR2_X1 U5333 ( .A(n6518), .B(n10093), .ZN(n6520) );
  XNOR2_X1 U5334 ( .A(n6472), .B(n10084), .ZN(n8155) );
  INV_X1 U5335 ( .A(n10158), .ZN(n10163) );
  INV_X1 U5336 ( .A(n9652), .ZN(n7675) );
  NAND2_X1 U5337 ( .A1(n6461), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6538) );
  OR2_X1 U5338 ( .A1(n6345), .A2(n9253), .ZN(n6347) );
  NAND2_X1 U5339 ( .A1(n6471), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6784) );
  NAND2_X1 U5341 ( .A1(n5778), .A2(n5777), .ZN(n5780) );
  OR2_X1 U5342 ( .A1(n6884), .A2(n5776), .ZN(n5778) );
  AND2_X1 U5343 ( .A1(n6482), .A2(n6485), .ZN(n6863) );
  INV_X1 U5344 ( .A(n6094), .ZN(n5666) );
  INV_X1 U5345 ( .A(n7489), .ZN(n5141) );
  NAND2_X1 U5346 ( .A1(n5382), .A2(n5379), .ZN(n10600) );
  AND2_X1 U5347 ( .A1(n5879), .A2(n5748), .ZN(n5924) );
  NAND2_X1 U5348 ( .A1(n5254), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n5324) );
  NAND4_X1 U5349 ( .A1(n6157), .A2(n5752), .A3(n6292), .A4(n6161), .ZN(n5753)
         );
  NAND2_X1 U5350 ( .A1(n5255), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5254) );
  OAI21_X1 U5351 ( .B1(P1_RD_REG_SCAN_IN), .B2(P2_ADDR_REG_19__SCAN_IN), .A(
        n5444), .ZN(n5323) );
  AND2_X1 U5352 ( .A1(n5247), .A2(n5246), .ZN(n6481) );
  AND2_X1 U5353 ( .A1(n5751), .A2(n5750), .ZN(n6157) );
  NOR2_X1 U5354 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_16__SCAN_IN), .ZN(
        n5751) );
  NOR2_X1 U5355 ( .A1(P2_IR_REG_15__SCAN_IN), .A2(P2_IR_REG_14__SCAN_IN), .ZN(
        n5750) );
  INV_X1 U5356 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n10062) );
  NOR2_X1 U5357 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6453) );
  NOR2_X1 U5358 ( .A1(P1_IR_REG_17__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n6452) );
  NOR2_X1 U5359 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_5__SCAN_IN), .ZN(
        n6451) );
  INV_X1 U5360 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n9846) );
  INV_X4 U5361 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3151) );
  NOR2_X1 U5362 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6544) );
  NOR2_X1 U5363 ( .A1(P1_IR_REG_2__SCAN_IN), .A2(P1_IR_REG_3__SCAN_IN), .ZN(
        n5533) );
  INV_X1 U5364 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n6013) );
  INV_X1 U5365 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6015) );
  INV_X1 U5366 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n5352) );
  INV_X1 U5367 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n5353) );
  INV_X1 U5368 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n6056) );
  INV_X1 U5369 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5444) );
  NOR2_X1 U5370 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_6__SCAN_IN), .ZN(
        n6016) );
  INV_X1 U5371 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n6053) );
  NAND4_X2 U5372 ( .A1(n5885), .A2(n5886), .A3(n5884), .A4(n5887), .ZN(n6695)
         );
  NAND2_X1 U5373 ( .A1(n5135), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5887) );
  OR2_X2 U5374 ( .A1(n7879), .A2(n7880), .ZN(n7931) );
  NAND2_X1 U5375 ( .A1(n6533), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n5695) );
  NAND2_X2 U5376 ( .A1(n9099), .A2(n8631), .ZN(n9094) );
  NAND4_X2 U5377 ( .A1(n6798), .A2(n6797), .A3(n6796), .A4(n6795), .ZN(n7175)
         );
  CLKBUF_X2 U5378 ( .A(n11006), .Z(n5142) );
  NAND4_X1 U5379 ( .A1(n6972), .A2(n6971), .A3(n6970), .A4(n6969), .ZN(n11006)
         );
  BUF_X4 U5380 ( .A(n7558), .Z(n5143) );
  NAND2_X1 U5381 ( .A1(n6522), .A2(n6520), .ZN(n7558) );
  OR2_X1 U5382 ( .A1(n5142), .A2(n11023), .ZN(n9543) );
  OAI22_X1 U5383 ( .A1(n7270), .A2(n7269), .B1(n7268), .B2(n5142), .ZN(n7395)
         );
  OR2_X1 U5384 ( .A1(n6800), .A2(n6793), .ZN(n8389) );
  AOI21_X2 U5385 ( .B1(n7922), .B2(n8594), .A(n5186), .ZN(n7960) );
  OAI21_X2 U5386 ( .B1(n7817), .B2(n8591), .A(n7816), .ZN(n7922) );
  NOR2_X2 U5387 ( .A1(n6489), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6492) );
  XNOR2_X1 U5388 ( .A(n5695), .B(n10089), .ZN(n6787) );
  OR2_X1 U5389 ( .A1(n6800), .A2(n6793), .ZN(n5146) );
  OAI21_X2 U5390 ( .B1(n9389), .B2(n8193), .A(n8192), .ZN(n9325) );
  NAND2_X2 U5391 ( .A1(n8176), .A2(n8175), .ZN(n9389) );
  AND2_X1 U5392 ( .A1(n5588), .A2(n6139), .ZN(n5587) );
  NAND2_X1 U5393 ( .A1(n6125), .A2(n5826), .ZN(n5588) );
  OAI21_X1 U5394 ( .B1(n7347), .B2(n5980), .A(n5979), .ZN(n7590) );
  OAI21_X1 U5395 ( .B1(n10806), .B2(n5610), .A(n5609), .ZN(n10822) );
  NAND2_X1 U5396 ( .A1(n5613), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5610) );
  NAND2_X1 U5397 ( .A1(n8925), .A2(n5613), .ZN(n5609) );
  INV_X1 U5398 ( .A(n10823), .ZN(n5613) );
  NAND2_X1 U5399 ( .A1(n5722), .A2(n5193), .ZN(n10222) );
  OR2_X1 U5400 ( .A1(n8121), .A2(n8062), .ZN(n9587) );
  INV_X1 U5401 ( .A(n8641), .ZN(n5434) );
  NAND2_X1 U5402 ( .A1(n5435), .A2(n5432), .ZN(n5431) );
  NAND2_X1 U5403 ( .A1(n9034), .A2(n8649), .ZN(n5433) );
  NAND2_X1 U5404 ( .A1(n5601), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5600) );
  INV_X1 U5405 ( .A(n10888), .ZN(n5371) );
  AND2_X1 U5406 ( .A1(n6403), .A2(n5181), .ZN(n5507) );
  NOR2_X1 U5407 ( .A1(n9058), .A2(n5525), .ZN(n5524) );
  INV_X1 U5408 ( .A(n5527), .ZN(n5525) );
  OR2_X1 U5409 ( .A1(n9175), .A2(n8727), .ZN(n8642) );
  NAND2_X1 U5410 ( .A1(n9175), .A2(n9075), .ZN(n5531) );
  OR2_X1 U5411 ( .A1(n9237), .A2(n9120), .ZN(n8631) );
  NOR2_X1 U5412 ( .A1(n6032), .A2(n6031), .ZN(n7586) );
  AND2_X1 U5413 ( .A1(n7593), .A2(n7591), .ZN(n6032) );
  OR2_X1 U5414 ( .A1(n8806), .A2(n9025), .ZN(n6260) );
  AND2_X1 U5415 ( .A1(n5755), .A2(n6346), .ZN(n5481) );
  NOR2_X1 U5416 ( .A1(n5753), .A2(n5665), .ZN(n5664) );
  NAND2_X1 U5417 ( .A1(n5754), .A2(n5749), .ZN(n5665) );
  INV_X1 U5418 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n5754) );
  INV_X1 U5419 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n6292) );
  INV_X1 U5420 ( .A(P2_IR_REG_8__SCAN_IN), .ZN(n6014) );
  OR2_X1 U5421 ( .A1(n9467), .A2(n9466), .ZN(n9642) );
  OR2_X1 U5422 ( .A1(n10257), .A2(n10269), .ZN(n9628) );
  INV_X1 U5423 ( .A(n10262), .ZN(n5290) );
  INV_X1 U5424 ( .A(n5309), .ZN(n5307) );
  NAND2_X1 U5425 ( .A1(n5309), .A2(n5305), .ZN(n5304) );
  INV_X1 U5426 ( .A(n5310), .ZN(n5305) );
  INV_X1 U5427 ( .A(n5341), .ZN(n5340) );
  NOR2_X1 U5428 ( .A1(n5706), .A2(n10195), .ZN(n5703) );
  OAI21_X1 U5429 ( .B1(n9456), .B2(n5543), .A(n5542), .ZN(n5541) );
  NAND2_X1 U5430 ( .A1(n10361), .A2(n5544), .ZN(n5540) );
  INV_X1 U5431 ( .A(n9516), .ZN(n5543) );
  OR2_X1 U5432 ( .A1(n9322), .A2(n9390), .ZN(n9595) );
  OR2_X1 U5433 ( .A1(n11175), .A2(n8119), .ZN(n5729) );
  OR2_X1 U5434 ( .A1(n11137), .A2(n11108), .ZN(n9523) );
  OR2_X1 U5435 ( .A1(n11088), .A2(n11110), .ZN(n9560) );
  NAND2_X1 U5436 ( .A1(n11088), .A2(n11110), .ZN(n11102) );
  INV_X1 U5437 ( .A(n10964), .ZN(n6814) );
  OAI21_X1 U5438 ( .B1(n8453), .B2(n9687), .A(n8452), .ZN(n8465) );
  OR2_X1 U5439 ( .A1(n8451), .A2(n8450), .ZN(n8452) );
  XNOR2_X1 U5440 ( .A(n8451), .B(n8450), .ZN(n8453) );
  AND2_X1 U5441 ( .A1(n5157), .A2(n10084), .ZN(n5160) );
  NAND2_X1 U5442 ( .A1(n5564), .A2(n5562), .ZN(n6263) );
  AOI21_X1 U5443 ( .B1(n5565), .B2(n5568), .A(n5563), .ZN(n5562) );
  INV_X1 U5444 ( .A(n5864), .ZN(n5563) );
  INV_X1 U5445 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U5446 ( .A1(n5592), .A2(n5232), .ZN(n6210) );
  INV_X1 U5447 ( .A(SI_21_), .ZN(n5841) );
  OAI21_X2 U5448 ( .B1(n6471), .B2(P1_IR_REG_19__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6783) );
  AND2_X1 U5449 ( .A1(n5839), .A2(n5838), .ZN(n6187) );
  AOI21_X1 U5450 ( .B1(n5587), .B2(n5584), .A(n5583), .ZN(n5582) );
  INV_X1 U5451 ( .A(n5830), .ZN(n5583) );
  INV_X1 U5452 ( .A(n5826), .ZN(n5584) );
  AND2_X1 U5453 ( .A1(n5830), .A2(n5829), .ZN(n6139) );
  AOI21_X1 U5454 ( .B1(n6099), .B2(n5285), .A(n5233), .ZN(n5283) );
  NAND2_X1 U5455 ( .A1(n6100), .A2(n5285), .ZN(n5284) );
  INV_X1 U5456 ( .A(n6051), .ZN(n5291) );
  OAI21_X1 U5457 ( .B1(n5134), .B2(n5597), .A(n5596), .ZN(n5770) );
  NAND2_X1 U5458 ( .A1(n5134), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n5596) );
  NAND2_X1 U5459 ( .A1(n8779), .A2(n8428), .ZN(n8430) );
  OR2_X1 U5460 ( .A1(n10822), .A2(n5241), .ZN(n5364) );
  NAND2_X1 U5461 ( .A1(n10899), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n10898) );
  NOR2_X1 U5462 ( .A1(n9123), .A2(n5461), .ZN(n5460) );
  INV_X1 U5463 ( .A(n6332), .ZN(n5461) );
  AOI21_X1 U5464 ( .B1(n5514), .B2(n5517), .A(n5511), .ZN(n5510) );
  INV_X1 U5465 ( .A(n9119), .ZN(n9136) );
  NAND2_X1 U5466 ( .A1(n6163), .A2(n6162), .ZN(n8786) );
  INV_X1 U5467 ( .A(n5926), .ZN(n6176) );
  INV_X1 U5468 ( .A(n6479), .ZN(n6175) );
  NAND2_X1 U5469 ( .A1(n6353), .A2(n6379), .ZN(n6494) );
  OAI21_X1 U5470 ( .B1(n10983), .B2(n8330), .A(n6890), .ZN(n6891) );
  INV_X1 U5471 ( .A(n6966), .ZN(n8377) );
  NOR2_X1 U5472 ( .A1(n10917), .A2(n5385), .ZN(n10614) );
  AND2_X1 U5473 ( .A1(n6863), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n5385) );
  AND2_X1 U5474 ( .A1(n5378), .A2(n5377), .ZN(n10642) );
  NAND2_X1 U5475 ( .A1(n6869), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n5377) );
  OR2_X1 U5476 ( .A1(n10642), .A2(n10641), .ZN(n5376) );
  OR2_X1 U5477 ( .A1(n10265), .A2(n5488), .ZN(n10224) );
  AND4_X1 U5478 ( .A1(n8367), .A2(n8366), .A3(n8365), .A4(n8364), .ZN(n10409)
         );
  INV_X1 U5479 ( .A(n6968), .ZN(n8357) );
  NAND2_X1 U5480 ( .A1(n10466), .A2(n10350), .ZN(n5707) );
  NAND2_X1 U5481 ( .A1(n8149), .A2(n9595), .ZN(n8150) );
  INV_X1 U5482 ( .A(n5345), .ZN(n5344) );
  INV_X1 U5483 ( .A(n9587), .ZN(n5346) );
  OR2_X1 U5484 ( .A1(n11137), .A2(n9673), .ZN(n5719) );
  INV_X1 U5485 ( .A(n5138), .ZN(n8215) );
  OR2_X1 U5486 ( .A1(n8465), .A2(n8464), .ZN(n8467) );
  NAND2_X1 U5487 ( .A1(n6319), .A2(n6318), .ZN(n8990) );
  NOR2_X1 U5488 ( .A1(n6317), .A2(n6316), .ZN(n6318) );
  NAND2_X1 U5489 ( .A1(n6304), .A2(n9130), .ZN(n6319) );
  INV_X1 U5490 ( .A(n10244), .ZN(n10419) );
  NAND2_X1 U5491 ( .A1(n5443), .A2(n5442), .ZN(n8572) );
  NAND2_X1 U5492 ( .A1(n8517), .A2(n8663), .ZN(n5443) );
  OAI21_X1 U5493 ( .B1(n8514), .B2(n8513), .A(n8676), .ZN(n5442) );
  AOI21_X1 U5494 ( .B1(n5408), .B2(n8593), .A(n8592), .ZN(n8605) );
  NAND2_X1 U5495 ( .A1(n5411), .A2(n5409), .ZN(n5408) );
  NAND2_X1 U5496 ( .A1(n9589), .A2(n9590), .ZN(n5276) );
  INV_X1 U5497 ( .A(n9619), .ZN(n5271) );
  NAND2_X1 U5498 ( .A1(n5269), .A2(n9640), .ZN(n5268) );
  INV_X1 U5499 ( .A(n10181), .ZN(n5269) );
  MUX2_X1 U5500 ( .A(n8623), .B(n8622), .S(n8663), .Z(n8634) );
  NAND2_X1 U5501 ( .A1(n9058), .A2(n5428), .ZN(n5425) );
  AOI21_X1 U5502 ( .B1(n5424), .B2(n9058), .A(n8650), .ZN(n5423) );
  INV_X1 U5503 ( .A(n5426), .ZN(n5424) );
  OR2_X1 U5504 ( .A1(n7628), .A2(n7570), .ZN(n8515) );
  OR2_X1 U5505 ( .A1(n9162), .A2(n9044), .ZN(n8651) );
  INV_X1 U5506 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5756) );
  AND2_X1 U5507 ( .A1(n10398), .A2(n10408), .ZN(n9473) );
  INV_X1 U5508 ( .A(SI_14_), .ZN(n9714) );
  INV_X1 U5509 ( .A(n5802), .ZN(n5418) );
  INV_X1 U5510 ( .A(n5997), .ZN(n5420) );
  AND2_X1 U5511 ( .A1(n8407), .A2(n8105), .ZN(n5689) );
  NAND2_X2 U5512 ( .A1(n6678), .A2(n6677), .ZN(n6752) );
  AND2_X1 U5513 ( .A1(n8525), .A2(n7119), .ZN(n6674) );
  AOI21_X1 U5514 ( .B1(n5211), .B2(n8666), .A(n5439), .ZN(n5438) );
  NOR2_X1 U5515 ( .A1(n8662), .A2(n8668), .ZN(n5439) );
  NAND2_X1 U5516 ( .A1(n8507), .A2(n8506), .ZN(n8509) );
  NAND2_X1 U5517 ( .A1(n9214), .A2(n8675), .ZN(n8506) );
  NAND2_X1 U5518 ( .A1(n5614), .A2(n8941), .ZN(n8953) );
  NAND2_X1 U5519 ( .A1(n5370), .A2(n5369), .ZN(n5614) );
  AOI21_X1 U5520 ( .B1(n5507), .B2(n5150), .A(n5209), .ZN(n5506) );
  NOR2_X1 U5521 ( .A1(n5402), .A2(n5401), .ZN(n5518) );
  INV_X1 U5522 ( .A(n6198), .ZN(n5401) );
  INV_X1 U5523 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n9752) );
  INV_X1 U5524 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n9767) );
  NAND2_X1 U5525 ( .A1(n8448), .A2(n8468), .ZN(n5591) );
  INV_X1 U5526 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5868) );
  INV_X1 U5527 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n5755) );
  INV_X1 U5528 ( .A(n5637), .ZN(n5636) );
  OAI21_X1 U5529 ( .B1(n7826), .B2(n5638), .A(n7825), .ZN(n5637) );
  NAND2_X1 U5530 ( .A1(n5641), .A2(n5640), .ZN(n5638) );
  NAND2_X1 U5531 ( .A1(n5630), .A2(n5185), .ZN(n5633) );
  INV_X1 U5532 ( .A(n7782), .ZN(n5630) );
  NAND2_X1 U5533 ( .A1(n7781), .A2(n7780), .ZN(n5640) );
  NAND2_X1 U5534 ( .A1(n5266), .A2(n5264), .ZN(n5263) );
  NOR2_X1 U5535 ( .A1(n10203), .A2(n5265), .ZN(n5264) );
  NAND2_X1 U5536 ( .A1(n9635), .A2(n5184), .ZN(n5266) );
  INV_X1 U5537 ( .A(n9637), .ZN(n5265) );
  NOR2_X1 U5538 ( .A1(n5201), .A2(n5262), .ZN(n5261) );
  NAND2_X1 U5539 ( .A1(n9643), .A2(n9642), .ZN(n5262) );
  NAND2_X1 U5540 ( .A1(n10171), .A2(n9466), .ZN(n9643) );
  NAND2_X1 U5541 ( .A1(n9649), .A2(n9641), .ZN(n5558) );
  INV_X1 U5542 ( .A(n10600), .ZN(n6846) );
  OR2_X1 U5543 ( .A1(n10244), .A2(n10409), .ZN(n9633) );
  INV_X1 U5544 ( .A(n9476), .ZN(n9623) );
  AOI21_X1 U5545 ( .B1(n5310), .B2(n5149), .A(n5207), .ZN(n5309) );
  NAND2_X1 U5546 ( .A1(n10341), .A2(n10355), .ZN(n5485) );
  OR2_X1 U5547 ( .A1(n10483), .A2(n9432), .ZN(n9602) );
  OR2_X1 U5548 ( .A1(n10488), .A2(n10378), .ZN(n9601) );
  OR2_X1 U5549 ( .A1(n9400), .A2(n8178), .ZN(n9591) );
  NOR2_X1 U5550 ( .A1(n7874), .A2(n7929), .ZN(n5487) );
  OR2_X1 U5551 ( .A1(n7929), .A2(n7981), .ZN(n9577) );
  NAND2_X1 U5552 ( .A1(n7632), .A2(n7884), .ZN(n5718) );
  INV_X1 U5553 ( .A(n9560), .ZN(n7543) );
  NAND2_X1 U5554 ( .A1(n5202), .A2(n5348), .ZN(n7547) );
  NOR2_X2 U5555 ( .A1(n7555), .A2(n11148), .ZN(n7637) );
  OR2_X1 U5556 ( .A1(n11148), .A2(n7884), .ZN(n9568) );
  NAND2_X1 U5557 ( .A1(n5549), .A2(n5547), .ZN(n7546) );
  NOR2_X1 U5558 ( .A1(n9483), .A2(n5548), .ZN(n5547) );
  INV_X1 U5559 ( .A(n9415), .ZN(n5548) );
  NAND2_X1 U5560 ( .A1(n7404), .A2(n9552), .ZN(n5549) );
  NAND2_X1 U5561 ( .A1(n5287), .A2(n5580), .ZN(n6173) );
  AOI21_X1 U5562 ( .B1(n5152), .B2(n5585), .A(n5234), .ZN(n5580) );
  NAND2_X1 U5563 ( .A1(n6126), .A2(n5152), .ZN(n5287) );
  AND2_X1 U5564 ( .A1(n6089), .A2(n5811), .ZN(n5814) );
  AOI21_X1 U5565 ( .B1(n5575), .B2(n5577), .A(n5574), .ZN(n5573) );
  INV_X1 U5566 ( .A(n5808), .ZN(n5574) );
  NAND2_X1 U5567 ( .A1(n5419), .A2(n5802), .ZN(n6012) );
  NAND2_X1 U5568 ( .A1(n5495), .A2(n5153), .ZN(n5419) );
  NAND2_X1 U5569 ( .A1(n6011), .A2(n5418), .ZN(n5417) );
  NAND2_X1 U5570 ( .A1(n5315), .A2(n5316), .ZN(n5496) );
  NAND2_X1 U5571 ( .A1(n5318), .A2(n5313), .ZN(n5315) );
  NAND2_X1 U5572 ( .A1(n5317), .A2(n5799), .ZN(n5316) );
  NOR2_X1 U5573 ( .A1(n5499), .A2(n5497), .ZN(n5313) );
  INV_X1 U5574 ( .A(n5973), .ZN(n5318) );
  OAI211_X1 U5575 ( .C1(n5324), .C2(n5322), .A(n5320), .B(n5319), .ZN(n5792)
         );
  NAND2_X1 U5576 ( .A1(n5321), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n5320) );
  OAI21_X1 U5577 ( .B1(n5134), .B2(n5399), .A(n5398), .ZN(n5400) );
  NAND2_X1 U5578 ( .A1(n5134), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n5398) );
  INV_X1 U5579 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6722) );
  NAND2_X1 U5580 ( .A1(n7891), .A2(n7890), .ZN(n5662) );
  NAND2_X1 U5581 ( .A1(n5681), .A2(n9045), .ZN(n5680) );
  INV_X1 U5582 ( .A(n8429), .ZN(n5681) );
  AOI21_X1 U5583 ( .B1(n5684), .B2(n7238), .A(n5243), .ZN(n5683) );
  INV_X1 U5584 ( .A(n8732), .ZN(n5673) );
  OR2_X1 U5585 ( .A1(n5678), .A2(n8432), .ZN(n5675) );
  NOR2_X1 U5586 ( .A1(n5679), .A2(n5148), .ZN(n5678) );
  INV_X1 U5587 ( .A(n8762), .ZN(n5679) );
  BUF_X1 U5588 ( .A(n5891), .Z(n7374) );
  NAND2_X1 U5589 ( .A1(n5137), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5894) );
  OAI21_X1 U5590 ( .B1(n6661), .B2(n6611), .A(n6612), .ZN(n6663) );
  XNOR2_X1 U5591 ( .A(n6613), .B(n7122), .ZN(n8854) );
  NAND2_X1 U5592 ( .A1(n5603), .A2(n5602), .ZN(n5601) );
  NAND2_X1 U5593 ( .A1(n6615), .A2(n6651), .ZN(n5604) );
  NAND2_X1 U5594 ( .A1(n5360), .A2(n5359), .ZN(n5354) );
  NAND2_X1 U5595 ( .A1(n6712), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n10758) );
  NAND2_X1 U5596 ( .A1(n10762), .A2(n10763), .ZN(n10761) );
  AND2_X1 U5597 ( .A1(n5331), .A2(n5330), .ZN(n8861) );
  NAND2_X1 U5598 ( .A1(n7257), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5330) );
  INV_X1 U5599 ( .A(n7255), .ZN(n5331) );
  OR2_X1 U5600 ( .A1(n10806), .A2(n8890), .ZN(n5612) );
  INV_X1 U5601 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n9967) );
  NAND2_X1 U5602 ( .A1(n5237), .A2(n5366), .ZN(n5365) );
  NAND2_X1 U5603 ( .A1(n10822), .A2(n5366), .ZN(n5363) );
  NAND3_X1 U5604 ( .A1(n5173), .A2(n5155), .A3(n5924), .ZN(n6094) );
  NOR2_X1 U5605 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_12__SCAN_IN), .ZN(
        n5747) );
  XNOR2_X1 U5606 ( .A(n8868), .B(n10829), .ZN(n10831) );
  AND2_X1 U5607 ( .A1(n5178), .A2(n5367), .ZN(n10856) );
  XNOR2_X1 U5608 ( .A(n8870), .B(n8933), .ZN(n10865) );
  NAND2_X1 U5609 ( .A1(n10865), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n10864) );
  NOR2_X1 U5610 ( .A1(n5473), .A2(n5478), .ZN(n9017) );
  INV_X1 U5611 ( .A(n5479), .ZN(n5474) );
  AOI21_X1 U5612 ( .B1(n5524), .B2(n5522), .A(n5212), .ZN(n5521) );
  INV_X1 U5613 ( .A(n5528), .ZN(n5522) );
  INV_X1 U5614 ( .A(n9174), .ZN(n5530) );
  INV_X1 U5615 ( .A(n5524), .ZN(n5523) );
  NAND2_X1 U5616 ( .A1(n5215), .A2(n5531), .ZN(n5527) );
  AND2_X1 U5617 ( .A1(n5531), .A2(n6336), .ZN(n5528) );
  NAND2_X1 U5618 ( .A1(n9094), .A2(n9093), .ZN(n5466) );
  INV_X1 U5619 ( .A(n5518), .ZN(n9074) );
  NOR2_X1 U5620 ( .A1(n6334), .A2(n8417), .ZN(n5458) );
  NAND2_X1 U5621 ( .A1(n9131), .A2(n6154), .ZN(n9115) );
  AOI21_X1 U5622 ( .B1(n5472), .B2(n8607), .A(n5470), .ZN(n5469) );
  INV_X1 U5623 ( .A(n5472), .ZN(n5471) );
  INV_X1 U5624 ( .A(n8611), .ZN(n5470) );
  AND2_X1 U5625 ( .A1(n8489), .A2(n8599), .ZN(n5472) );
  NAND2_X1 U5626 ( .A1(n7960), .A2(n6330), .ZN(n7959) );
  INV_X1 U5627 ( .A(n8834), .ZN(n7947) );
  NOR2_X1 U5628 ( .A1(n7586), .A2(n5169), .ZN(n6033) );
  AND4_X1 U5629 ( .A1(n6048), .A2(n6047), .A3(n6046), .A4(n6045), .ZN(n7849)
         );
  AND2_X1 U5630 ( .A1(n8579), .A2(n8580), .ZN(n8486) );
  OR2_X1 U5631 ( .A1(n7664), .A2(n7510), .ZN(n8516) );
  NAND2_X1 U5632 ( .A1(n7477), .A2(n8573), .ZN(n5452) );
  NAND2_X1 U5633 ( .A1(n6629), .A2(n6500), .ZN(n7099) );
  NAND2_X1 U5634 ( .A1(n6686), .A2(n8663), .ZN(n9121) );
  OR2_X1 U5635 ( .A1(n6686), .A2(n8676), .ZN(n9119) );
  INV_X1 U5636 ( .A(n9121), .ZN(n9133) );
  OR2_X1 U5637 ( .A1(n8168), .A2(n6679), .ZN(n8534) );
  NAND2_X1 U5638 ( .A1(n8168), .A2(n6679), .ZN(n8526) );
  NAND2_X1 U5639 ( .A1(n8463), .A2(n8462), .ZN(n8689) );
  NAND2_X1 U5640 ( .A1(n5591), .A2(n6270), .ZN(n9155) );
  AOI21_X1 U5641 ( .B1(n9001), .B2(n9130), .A(n5405), .ZN(n9157) );
  NAND2_X1 U5642 ( .A1(n5407), .A2(n5406), .ZN(n5405) );
  NAND2_X1 U5643 ( .A1(n9025), .A2(n9136), .ZN(n5406) );
  NAND2_X1 U5644 ( .A1(n6190), .A2(n6189), .ZN(n8768) );
  NAND2_X1 U5645 ( .A1(n6116), .A2(n6115), .ZN(n8404) );
  INV_X1 U5646 ( .A(n9173), .ZN(n9180) );
  XNOR2_X1 U5647 ( .A(n6352), .B(P2_IR_REG_26__SCAN_IN), .ZN(n6379) );
  OR2_X1 U5648 ( .A1(n6351), .A2(n9253), .ZN(n6352) );
  NAND2_X1 U5649 ( .A1(n6294), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6298) );
  INV_X1 U5650 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n6297) );
  NAND2_X1 U5651 ( .A1(n6298), .A2(n6297), .ZN(n6300) );
  AND2_X1 U5652 ( .A1(n9253), .A2(n5748), .ZN(n5350) );
  AND2_X2 U5653 ( .A1(n6571), .A2(n6475), .ZN(n6800) );
  NAND2_X1 U5654 ( .A1(n5645), .A2(n5646), .ZN(n9302) );
  AND2_X1 U5655 ( .A1(n5647), .A2(n9335), .ZN(n5646) );
  NAND2_X1 U5656 ( .A1(n5726), .A2(n5651), .ZN(n5647) );
  NOR2_X1 U5657 ( .A1(n7781), .A2(n7780), .ZN(n5641) );
  INV_X1 U5658 ( .A(n5640), .ZN(n5639) );
  NOR2_X1 U5659 ( .A1(n9296), .A2(n5657), .ZN(n5656) );
  INV_X1 U5660 ( .A(n8249), .ZN(n5657) );
  NAND2_X1 U5661 ( .A1(n5656), .A2(n5654), .ZN(n5653) );
  INV_X1 U5662 ( .A(n9344), .ZN(n5654) );
  INV_X1 U5663 ( .A(n7055), .ZN(n6953) );
  OR2_X1 U5664 ( .A1(n6968), .A2(n10992), .ZN(n6765) );
  INV_X1 U5665 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6450) );
  NOR2_X1 U5666 ( .A1(n10654), .A2(n5227), .ZN(n10671) );
  NOR2_X1 U5667 ( .A1(n10670), .A2(n10671), .ZN(n10669) );
  NOR3_X1 U5668 ( .A1(n10265), .A2(n10398), .A3(n5488), .ZN(n10206) );
  AOI21_X1 U5669 ( .B1(n5200), .B2(n5339), .A(n5279), .ZN(n5278) );
  INV_X1 U5670 ( .A(n10186), .ZN(n5279) );
  AOI21_X1 U5671 ( .B1(n5339), .B2(n5340), .A(n5336), .ZN(n5335) );
  INV_X1 U5672 ( .A(n5534), .ZN(n5336) );
  AOI21_X1 U5673 ( .B1(n5538), .B2(n5536), .A(n5535), .ZN(n5534) );
  INV_X1 U5674 ( .A(n10185), .ZN(n5535) );
  NAND2_X1 U5675 ( .A1(n9628), .A2(n10186), .ZN(n10249) );
  INV_X1 U5676 ( .A(n5537), .ZN(n5538) );
  NOR2_X1 U5677 ( .A1(n5338), .A2(n5340), .ZN(n10284) );
  AOI21_X1 U5678 ( .B1(n5703), .B2(n5700), .A(n5213), .ZN(n5699) );
  INV_X1 U5679 ( .A(n5708), .ZN(n5700) );
  INV_X1 U5680 ( .A(n5703), .ZN(n5701) );
  AND2_X1 U5681 ( .A1(n10182), .A2(n10181), .ZN(n10290) );
  NOR2_X1 U5682 ( .A1(n10194), .A2(n10319), .ZN(n5708) );
  AND4_X1 U5683 ( .A1(n8283), .A2(n8282), .A3(n8281), .A4(n8280), .ZN(n10329)
         );
  AND2_X1 U5684 ( .A1(n5159), .A2(n9455), .ZN(n5546) );
  NAND2_X1 U5685 ( .A1(n5308), .A2(n5309), .ZN(n10320) );
  NAND2_X1 U5686 ( .A1(n10353), .A2(n5310), .ZN(n5308) );
  INV_X1 U5687 ( .A(n10454), .ZN(n10350) );
  NAND2_X1 U5688 ( .A1(n10372), .A2(n9602), .ZN(n10363) );
  AND2_X1 U5689 ( .A1(n9455), .A2(n9608), .ZN(n10362) );
  NOR2_X1 U5690 ( .A1(n8039), .A2(n9400), .ZN(n8091) );
  AND4_X1 U5691 ( .A1(n8027), .A2(n8026), .A3(n8025), .A4(n8024), .ZN(n9390)
         );
  OR2_X1 U5692 ( .A1(n8036), .A2(n5301), .ZN(n5298) );
  NAND2_X1 U5693 ( .A1(n5216), .A2(n5302), .ZN(n5297) );
  NAND2_X1 U5694 ( .A1(n5303), .A2(n5729), .ZN(n5300) );
  AND2_X1 U5695 ( .A1(n9591), .A2(n9593), .ZN(n9496) );
  INV_X1 U5696 ( .A(n5729), .ZN(n5301) );
  NAND2_X1 U5697 ( .A1(n7986), .A2(n5176), .ZN(n8028) );
  AND4_X1 U5698 ( .A1(n7808), .A2(n7807), .A3(n7806), .A4(n7805), .ZN(n8062)
         );
  AND2_X1 U5699 ( .A1(n7929), .A2(n11171), .ZN(n5325) );
  AND4_X1 U5700 ( .A1(n7562), .A2(n7561), .A3(n7560), .A4(n7559), .ZN(n7872)
         );
  NAND2_X1 U5701 ( .A1(n5716), .A2(n5718), .ZN(n5715) );
  NAND2_X1 U5702 ( .A1(n9489), .A2(n5717), .ZN(n5716) );
  NAND2_X1 U5703 ( .A1(n9569), .A2(n5719), .ZN(n5717) );
  NAND2_X1 U5704 ( .A1(n5718), .A2(n5719), .ZN(n5714) );
  NAND2_X1 U5705 ( .A1(n9533), .A2(n9568), .ZN(n9489) );
  AND4_X1 U5706 ( .A1(n7418), .A2(n7417), .A3(n7416), .A4(n7415), .ZN(n11084)
         );
  NAND2_X1 U5707 ( .A1(n7385), .A2(n11035), .ZN(n5697) );
  OR2_X1 U5708 ( .A1(n5133), .A2(n10600), .ZN(n5467) );
  AND2_X1 U5709 ( .A1(n7168), .A2(n7167), .ZN(n7714) );
  AOI21_X1 U5710 ( .B1(n9452), .B2(n8029), .A(n9451), .ZN(n10393) );
  INV_X1 U5711 ( .A(n10176), .ZN(n10396) );
  AND2_X1 U5712 ( .A1(n8253), .A2(n8252), .ZN(n10466) );
  OR2_X1 U5713 ( .A1(n5145), .A2(n9469), .ZN(n11109) );
  NAND2_X1 U5714 ( .A1(n7187), .A2(n5145), .ZN(n11107) );
  NAND2_X1 U5715 ( .A1(n7183), .A2(n7182), .ZN(n11181) );
  INV_X1 U5716 ( .A(n11181), .ZN(n11104) );
  AND2_X1 U5717 ( .A1(n6573), .A2(n6576), .ZN(n6780) );
  NAND2_X1 U5718 ( .A1(n8467), .A2(n8466), .ZN(n9446) );
  NAND2_X1 U5719 ( .A1(n6532), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6535) );
  INV_X1 U5720 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n10084) );
  NAND2_X1 U5721 ( .A1(n5561), .A2(n5565), .ZN(n5865) );
  XNOR2_X1 U5722 ( .A(n5277), .B(n6248), .ZN(n8319) );
  NAND2_X1 U5723 ( .A1(n6245), .A2(n6244), .ZN(n5277) );
  NAND2_X1 U5724 ( .A1(n6233), .A2(n6232), .ZN(n6245) );
  INV_X1 U5725 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n10082) );
  XNOR2_X1 U5726 ( .A(n6464), .B(P1_IR_REG_23__SCAN_IN), .ZN(n7913) );
  INV_X1 U5727 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6460) );
  NAND2_X1 U5728 ( .A1(n5581), .A2(n5582), .ZN(n6156) );
  OR2_X1 U5729 ( .A1(n6126), .A2(n5585), .ZN(n5581) );
  NAND2_X1 U5730 ( .A1(n5586), .A2(n5826), .ZN(n6140) );
  OR2_X1 U5731 ( .A1(n6068), .A2(n6067), .ZN(n6090) );
  NAND2_X1 U5732 ( .A1(n6012), .A2(n6011), .ZN(n5578) );
  NAND2_X1 U5733 ( .A1(n5961), .A2(n5791), .ZN(n5974) );
  NAND2_X1 U5734 ( .A1(n5974), .A2(n5973), .ZN(n5976) );
  NAND2_X1 U5735 ( .A1(n5959), .A2(n5958), .ZN(n5961) );
  INV_X1 U5736 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n5246) );
  NAND2_X1 U5737 ( .A1(n5134), .A2(n5772), .ZN(n5259) );
  NAND2_X1 U5738 ( .A1(n5770), .A2(SI_1_), .ZN(n5773) );
  INV_X1 U5739 ( .A(n5770), .ZN(n5260) );
  AND2_X1 U5740 ( .A1(n8434), .A2(n8735), .ZN(n8435) );
  INV_X1 U5741 ( .A(n9025), .ZN(n8735) );
  XOR2_X1 U5742 ( .A(n8828), .B(n8433), .Z(n8732) );
  NAND2_X1 U5743 ( .A1(n6235), .A2(n6234), .ZN(n9039) );
  NAND2_X1 U5744 ( .A1(n8426), .A2(n8425), .ZN(n8779) );
  NAND2_X1 U5745 ( .A1(n6243), .A2(n6242), .ZN(n9054) );
  INV_X1 U5746 ( .A(n7849), .ZN(n8836) );
  NAND2_X1 U5747 ( .A1(n8874), .A2(n10898), .ZN(n8951) );
  NOR2_X1 U5748 ( .A1(n8973), .A2(n5618), .ZN(n5617) );
  NAND2_X1 U5749 ( .A1(n8963), .A2(n5619), .ZN(n5618) );
  NAND2_X1 U5750 ( .A1(n5621), .A2(n10790), .ZN(n5620) );
  XNOR2_X1 U5751 ( .A(n8960), .B(n8969), .ZN(n5621) );
  AOI21_X1 U5752 ( .B1(n10907), .B2(n8959), .A(n8958), .ZN(n8960) );
  XNOR2_X1 U5753 ( .A(n9007), .B(n9006), .ZN(n9156) );
  NAND2_X1 U5754 ( .A1(n6041), .A2(n6040), .ZN(n7741) );
  NAND2_X1 U5755 ( .A1(n5140), .A2(n7857), .ZN(n9173) );
  AND2_X1 U5756 ( .A1(n8995), .A2(n9204), .ZN(n6344) );
  NAND2_X1 U5757 ( .A1(n7403), .A2(n7402), .ZN(n11088) );
  NAND2_X1 U5758 ( .A1(n5256), .A2(n8029), .ZN(n7403) );
  INV_X1 U5759 ( .A(n7400), .ZN(n5256) );
  OR2_X1 U5760 ( .A1(n8057), .A2(n8056), .ZN(n5725) );
  AND4_X1 U5761 ( .A1(n8311), .A2(n8310), .A3(n8309), .A4(n8308), .ZN(n10297)
         );
  NAND2_X1 U5762 ( .A1(n8302), .A2(n8301), .ZN(n10442) );
  INV_X1 U5763 ( .A(n7394), .ZN(n7004) );
  NAND2_X1 U5764 ( .A1(n7530), .A2(n7529), .ZN(n11137) );
  INV_X1 U5765 ( .A(n10341), .ZN(n10473) );
  INV_X1 U5766 ( .A(n7992), .ZN(n11175) );
  NAND2_X1 U5767 ( .A1(n8274), .A2(n8273), .ZN(n10306) );
  NAND2_X1 U5768 ( .A1(n6942), .A2(n6941), .ZN(n5625) );
  INV_X1 U5769 ( .A(n11064), .ZN(n11035) );
  NAND2_X1 U5770 ( .A1(n6813), .A2(n6811), .ZN(n9402) );
  NAND2_X1 U5771 ( .A1(n6815), .A2(n10968), .ZN(n9399) );
  NAND2_X1 U5772 ( .A1(n9656), .A2(n9651), .ZN(n9653) );
  NAND2_X1 U5773 ( .A1(n5554), .A2(n6816), .ZN(n5553) );
  INV_X1 U5774 ( .A(n9665), .ZN(n5554) );
  INV_X1 U5775 ( .A(n10329), .ZN(n10463) );
  INV_X1 U5776 ( .A(n5384), .ZN(n10612) );
  INV_X1 U5777 ( .A(n5376), .ZN(n10640) );
  NAND2_X1 U5778 ( .A1(n6855), .A2(n6856), .ZN(n7355) );
  AOI21_X1 U5779 ( .B1(n10744), .B2(n10730), .A(n5251), .ZN(n5250) );
  OAI21_X1 U5780 ( .B1(n10733), .B2(n10732), .A(n10731), .ZN(n5251) );
  NOR2_X1 U5781 ( .A1(n10723), .A2(n10724), .ZN(n10722) );
  XNOR2_X1 U5782 ( .A(n10218), .B(n5289), .ZN(n10414) );
  NAND2_X1 U5783 ( .A1(n5722), .A2(n10200), .ZN(n10219) );
  AND2_X1 U5784 ( .A1(n10224), .A2(n10223), .ZN(n10410) );
  INV_X2 U5785 ( .A(n11123), .ZN(n10968) );
  OR2_X1 U5786 ( .A1(n6574), .A2(n6806), .ZN(n10506) );
  INV_X1 U5787 ( .A(n8572), .ZN(n8521) );
  INV_X1 U5788 ( .A(n5410), .ZN(n5409) );
  OAI21_X1 U5789 ( .B1(n8584), .B2(n8676), .A(n5511), .ZN(n5410) );
  NAND2_X1 U5790 ( .A1(n5412), .A2(n8676), .ZN(n5411) );
  NAND2_X1 U5791 ( .A1(n5413), .A2(n8579), .ZN(n5412) );
  NAND2_X1 U5792 ( .A1(n8576), .A2(n8575), .ZN(n5413) );
  OAI21_X1 U5793 ( .B1(n5276), .B2(n9592), .A(n9594), .ZN(n5273) );
  INV_X1 U5794 ( .A(n8637), .ZN(n5432) );
  AND3_X1 U5795 ( .A1(n5274), .A2(n5272), .A3(n10191), .ZN(n9600) );
  NAND2_X1 U5796 ( .A1(n5275), .A2(n9640), .ZN(n5274) );
  NAND2_X1 U5797 ( .A1(n5273), .A2(n9644), .ZN(n5272) );
  OAI21_X1 U5798 ( .B1(n5276), .B2(n9596), .A(n9595), .ZN(n5275) );
  AOI21_X1 U5799 ( .B1(n8616), .B2(n8615), .A(n8614), .ZN(n8624) );
  MUX2_X1 U5800 ( .A(n8604), .B(n8603), .S(n8663), .Z(n8616) );
  AOI21_X1 U5801 ( .B1(n5428), .B2(n5430), .A(n5427), .ZN(n5426) );
  INV_X1 U5802 ( .A(n8644), .ZN(n5427) );
  OAI21_X1 U5803 ( .B1(n5270), .B2(n5180), .A(n5267), .ZN(n9625) );
  AND2_X1 U5804 ( .A1(n10283), .A2(n5268), .ZN(n5267) );
  AOI21_X1 U5805 ( .B1(n9614), .B2(n9615), .A(n5271), .ZN(n5270) );
  INV_X1 U5806 ( .A(SI_17_), .ZN(n9913) );
  INV_X1 U5807 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n10032) );
  AOI21_X1 U5808 ( .B1(n5423), .B2(n5425), .A(n5433), .ZN(n5422) );
  OAI211_X1 U5809 ( .C1(n8634), .C2(n8633), .A(n9093), .B(n8632), .ZN(n8638)
         );
  INV_X1 U5810 ( .A(n8662), .ZN(n5441) );
  INV_X1 U5811 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n9951) );
  NAND2_X1 U5812 ( .A1(n6932), .A2(n6695), .ZN(n8535) );
  NAND2_X1 U5813 ( .A1(n7860), .A2(n8110), .ZN(n5395) );
  NOR2_X1 U5814 ( .A1(n5532), .A2(n5394), .ZN(n5393) );
  INV_X1 U5815 ( .A(n6081), .ZN(n5394) );
  NOR2_X1 U5816 ( .A1(n7860), .A2(n8110), .ZN(n5532) );
  INV_X1 U5817 ( .A(n5348), .ZN(n9486) );
  INV_X1 U5818 ( .A(n9638), .ZN(n5560) );
  AOI21_X1 U5819 ( .B1(n10290), .B2(n5342), .A(n10183), .ZN(n5341) );
  INV_X1 U5820 ( .A(n10180), .ZN(n5342) );
  AND2_X1 U5821 ( .A1(n10299), .A2(n10312), .ZN(n10183) );
  NOR2_X1 U5822 ( .A1(n5545), .A2(n9514), .ZN(n5544) );
  NAND2_X1 U5823 ( .A1(n9532), .A2(n11102), .ZN(n5348) );
  NAND2_X1 U5824 ( .A1(n6411), .A2(n6410), .ZN(n8451) );
  INV_X1 U5825 ( .A(SI_18_), .ZN(n9912) );
  NOR2_X1 U5826 ( .A1(n5821), .A2(n5286), .ZN(n5285) );
  INV_X1 U5827 ( .A(n5818), .ZN(n5286) );
  NAND2_X1 U5828 ( .A1(n5989), .A2(n5499), .ZN(n5317) );
  INV_X1 U5829 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n9966) );
  NAND2_X1 U5830 ( .A1(n8677), .A2(n8689), .ZN(n8508) );
  AND3_X1 U5831 ( .A1(n5605), .A2(n5606), .A3(n5236), .ZN(n8919) );
  NAND2_X1 U5832 ( .A1(n10813), .A2(n8867), .ZN(n8868) );
  OR2_X1 U5833 ( .A1(n8665), .A2(n8664), .ZN(n6417) );
  OAI21_X1 U5834 ( .B1(n5154), .B2(n8646), .A(n5210), .ZN(n5478) );
  NOR2_X1 U5835 ( .A1(n5154), .A2(n9052), .ZN(n5479) );
  INV_X1 U5836 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n7258) );
  NAND2_X1 U5837 ( .A1(n5397), .A2(n6029), .ZN(n7589) );
  NAND2_X1 U5838 ( .A1(n8519), .A2(n7500), .ZN(n7616) );
  OR2_X1 U5839 ( .A1(n5965), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5982) );
  INV_X1 U5840 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n9975) );
  AND2_X1 U5841 ( .A1(n8660), .A2(n8661), .ZN(n8998) );
  NAND2_X1 U5842 ( .A1(n9000), .A2(n9133), .ZN(n5407) );
  NOR2_X1 U5843 ( .A1(n5523), .A2(n9048), .ZN(n5520) );
  OAI21_X1 U5844 ( .B1(n5521), .B2(n9048), .A(n5203), .ZN(n5519) );
  NAND2_X1 U5845 ( .A1(n5392), .A2(n5390), .ZN(n7917) );
  NOR2_X1 U5846 ( .A1(n8594), .A2(n5391), .ZN(n5390) );
  INV_X1 U5847 ( .A(n5395), .ZN(n5391) );
  OR2_X1 U5848 ( .A1(n6494), .A2(n6369), .ZN(n6388) );
  XNOR2_X1 U5849 ( .A(n5869), .B(n5868), .ZN(n6305) );
  INV_X1 U5850 ( .A(n9337), .ZN(n5651) );
  AND2_X1 U5851 ( .A1(P1_REG3_REG_20__SCAN_IN), .A2(n8238), .ZN(n8237) );
  AND2_X1 U5852 ( .A1(n8255), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n6735) );
  AND2_X1 U5853 ( .A1(n8237), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8255) );
  NAND2_X1 U5854 ( .A1(n9325), .A2(n9327), .ZN(n5644) );
  AND2_X1 U5855 ( .A1(n8304), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8321) );
  AND2_X1 U5856 ( .A1(n8336), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n8359) );
  OR2_X1 U5857 ( .A1(n5489), .A2(n10412), .ZN(n5488) );
  NAND2_X1 U5858 ( .A1(n10419), .A2(n5490), .ZN(n5489) );
  INV_X1 U5859 ( .A(n10249), .ZN(n5281) );
  INV_X1 U5860 ( .A(n10283), .ZN(n5536) );
  INV_X1 U5861 ( .A(n10424), .ZN(n10196) );
  AND2_X1 U5862 ( .A1(n6837), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8304) );
  AND2_X1 U5863 ( .A1(n6735), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n6837) );
  NAND2_X1 U5864 ( .A1(n10290), .A2(n10194), .ZN(n5343) );
  NAND2_X1 U5865 ( .A1(n5484), .A2(n10466), .ZN(n5483) );
  INV_X1 U5866 ( .A(n5485), .ZN(n5484) );
  NOR2_X1 U5867 ( .A1(n10346), .A2(n5311), .ZN(n5310) );
  NOR2_X1 U5868 ( .A1(n5149), .A2(n10193), .ZN(n5311) );
  AND2_X1 U5869 ( .A1(n8091), .A2(n11196), .ZN(n8135) );
  AND2_X1 U5870 ( .A1(n5298), .A2(n5175), .ZN(n5294) );
  NOR2_X1 U5871 ( .A1(n11188), .A2(n8178), .ZN(n5293) );
  AND2_X1 U5872 ( .A1(n9535), .A2(n9532), .ZN(n11101) );
  NAND2_X1 U5873 ( .A1(n11061), .A2(n9674), .ZN(n9561) );
  AND2_X1 U5874 ( .A1(n9559), .A2(n9561), .ZN(n9554) );
  NOR2_X1 U5875 ( .A1(n7268), .A2(n7004), .ZN(n5493) );
  OR2_X1 U5876 ( .A1(n11019), .A2(n7394), .ZN(n9544) );
  INV_X1 U5877 ( .A(n7179), .ZN(n7180) );
  AND2_X1 U5878 ( .A1(n6262), .A2(n5863), .ZN(n5864) );
  INV_X1 U5879 ( .A(n5566), .ZN(n5565) );
  OAI21_X1 U5880 ( .B1(n5568), .B2(n5852), .A(n5567), .ZN(n5566) );
  OR2_X1 U5881 ( .A1(n5859), .A2(n5860), .ZN(n5567) );
  NAND2_X1 U5882 ( .A1(n6246), .A2(n6232), .ZN(n5568) );
  NAND2_X1 U5883 ( .A1(n6222), .A2(n5852), .ZN(n6233) );
  NOR2_X1 U5884 ( .A1(n5842), .A2(n5594), .ZN(n5593) );
  INV_X1 U5885 ( .A(n5839), .ZN(n5594) );
  INV_X1 U5886 ( .A(n5587), .ZN(n5585) );
  INV_X1 U5887 ( .A(SI_16_), .ZN(n5822) );
  INV_X1 U5888 ( .A(SI_10_), .ZN(n9923) );
  NAND2_X1 U5889 ( .A1(n5400), .A2(SI_2_), .ZN(n5775) );
  INV_X1 U5890 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5255) );
  NAND2_X1 U5891 ( .A1(n8424), .A2(n6680), .ZN(n6681) );
  AOI21_X1 U5892 ( .B1(n5668), .B2(n8418), .A(n5230), .ZN(n5667) );
  OR2_X1 U5893 ( .A1(n5690), .A2(n5687), .ZN(n5686) );
  INV_X1 U5894 ( .A(n8407), .ZN(n5687) );
  NAND2_X1 U5895 ( .A1(n5743), .A2(n9966), .ZN(n6213) );
  INV_X1 U5896 ( .A(n6203), .ZN(n5743) );
  NAND2_X1 U5897 ( .A1(n7705), .A2(n7704), .ZN(n7844) );
  XNOR2_X1 U5898 ( .A(n6682), .B(n6752), .ZN(n6724) );
  AND2_X1 U5899 ( .A1(n8812), .A2(n8402), .ZN(n5690) );
  INV_X1 U5900 ( .A(n8672), .ZN(n8507) );
  NAND2_X1 U5901 ( .A1(n5437), .A2(n5436), .ZN(n8681) );
  AOI21_X1 U5902 ( .B1(n5438), .B2(n5440), .A(n8669), .ZN(n5436) );
  NOR2_X1 U5903 ( .A1(n8667), .A2(n8666), .ZN(n5440) );
  AND2_X1 U5904 ( .A1(n9217), .A2(n8825), .ZN(n8677) );
  NAND2_X1 U5905 ( .A1(n5914), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5919) );
  XNOR2_X1 U5906 ( .A(n5871), .B(n5870), .ZN(n6580) );
  NAND2_X1 U5907 ( .A1(n5482), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5871) );
  AND2_X1 U5908 ( .A1(n5481), .A2(n5691), .ZN(n5480) );
  OR2_X1 U5909 ( .A1(n6663), .A2(n6662), .ZN(n6665) );
  INV_X1 U5910 ( .A(n5600), .ZN(n5599) );
  NAND2_X1 U5911 ( .A1(n5600), .A2(n5604), .ZN(n6616) );
  NAND2_X1 U5912 ( .A1(n6616), .A2(n6617), .ZN(n6709) );
  NAND2_X1 U5913 ( .A1(n5354), .A2(n5199), .ZN(n5356) );
  OR2_X1 U5914 ( .A1(n7220), .A2(n7221), .ZN(n5606) );
  NAND2_X1 U5915 ( .A1(n5356), .A2(n5355), .ZN(n7220) );
  NAND2_X1 U5916 ( .A1(n10761), .A2(n5195), .ZN(n5328) );
  XNOR2_X1 U5917 ( .A(n5328), .B(n7215), .ZN(n7209) );
  XNOR2_X1 U5918 ( .A(n8919), .B(n8920), .ZN(n8922) );
  NAND2_X1 U5919 ( .A1(n8862), .A2(n8863), .ZN(n10785) );
  NAND2_X1 U5920 ( .A1(n10801), .A2(n8866), .ZN(n10814) );
  NAND2_X1 U5921 ( .A1(n10814), .A2(n10815), .ZN(n10813) );
  AND2_X1 U5922 ( .A1(n5363), .A2(n5362), .ZN(n5361) );
  AND2_X1 U5923 ( .A1(n5365), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5362) );
  OR2_X1 U5924 ( .A1(n10856), .A2(n10857), .ZN(n10854) );
  NAND2_X1 U5925 ( .A1(n10864), .A2(n8872), .ZN(n10881) );
  INV_X1 U5926 ( .A(n8870), .ZN(n8871) );
  OAI22_X1 U5927 ( .A1(n10872), .A2(n5368), .B1(n5242), .B2(n5371), .ZN(n8939)
         );
  OR2_X1 U5928 ( .A1(n8935), .A2(n5242), .ZN(n5368) );
  XNOR2_X1 U5929 ( .A(n8873), .B(n10897), .ZN(n10899) );
  NAND2_X1 U5930 ( .A1(n10880), .A2(n5326), .ZN(n8873) );
  OR2_X1 U5931 ( .A1(n10879), .A2(n9207), .ZN(n5326) );
  NAND2_X1 U5932 ( .A1(n10895), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n5619) );
  NAND2_X1 U5933 ( .A1(n8955), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n8956) );
  NAND2_X1 U5934 ( .A1(n8954), .A2(n8965), .ZN(n8957) );
  NOR2_X1 U5935 ( .A1(n10908), .A2(n9144), .ZN(n10907) );
  NAND2_X1 U5936 ( .A1(n8669), .A2(n5506), .ZN(n5505) );
  OAI21_X1 U5937 ( .B1(n5509), .B2(n5158), .A(n5501), .ZN(n5500) );
  NAND2_X1 U5938 ( .A1(n5509), .A2(n5506), .ZN(n5501) );
  INV_X1 U5939 ( .A(n5507), .ZN(n5502) );
  NAND2_X1 U5940 ( .A1(n5591), .A2(n5589), .ZN(n8660) );
  NOR2_X1 U5941 ( .A1(n9015), .A2(n5590), .ZN(n5589) );
  INV_X1 U5942 ( .A(n6270), .ZN(n5590) );
  OAI21_X1 U5943 ( .B1(n9056), .B2(n5476), .A(n5475), .ZN(n9005) );
  NAND2_X1 U5944 ( .A1(n5479), .A2(n5477), .ZN(n5476) );
  NAND2_X1 U5945 ( .A1(n5478), .A2(n5477), .ZN(n5475) );
  INV_X1 U5946 ( .A(n8656), .ZN(n5477) );
  OR2_X1 U5947 ( .A1(n8656), .A2(n9004), .ZN(n9016) );
  NAND2_X1 U5948 ( .A1(n9057), .A2(n8646), .ZN(n9049) );
  NAND2_X1 U5949 ( .A1(n5744), .A2(n9979), .ZN(n6251) );
  INV_X1 U5950 ( .A(n6236), .ZN(n5744) );
  OR2_X1 U5951 ( .A1(n6224), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6236) );
  OR2_X1 U5952 ( .A1(n9056), .A2(n9052), .ZN(n9057) );
  AOI21_X1 U5953 ( .B1(n5464), .B2(n5463), .A(n5217), .ZN(n5462) );
  INV_X1 U5954 ( .A(n6179), .ZN(n5742) );
  NAND2_X1 U5955 ( .A1(n5494), .A2(n6171), .ZN(n9101) );
  INV_X1 U5956 ( .A(n6147), .ZN(n5741) );
  NAND2_X1 U5957 ( .A1(n5740), .A2(n10000), .ZN(n6132) );
  INV_X1 U5958 ( .A(n6117), .ZN(n5740) );
  OR2_X1 U5959 ( .A1(n6132), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6147) );
  NAND2_X1 U5960 ( .A1(n5739), .A2(n5738), .ZN(n6104) );
  OR2_X1 U5961 ( .A1(n8590), .A2(n8591), .ZN(n8589) );
  NAND2_X1 U5962 ( .A1(n5737), .A2(n9967), .ZN(n6083) );
  INV_X1 U5963 ( .A(n6075), .ZN(n5737) );
  AOI21_X1 U5964 ( .B1(n5515), .B2(n5151), .A(n5182), .ZN(n5514) );
  NOR2_X1 U5965 ( .A1(n5516), .A2(n6049), .ZN(n5515) );
  INV_X1 U5966 ( .A(n6050), .ZN(n5516) );
  NAND2_X1 U5967 ( .A1(n5151), .A2(n6050), .ZN(n5517) );
  OR2_X1 U5968 ( .A1(n6043), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U5969 ( .A1(n5736), .A2(n7258), .ZN(n6043) );
  INV_X1 U5970 ( .A(n6023), .ZN(n5736) );
  AOI21_X1 U5971 ( .B1(n7133), .B2(n6324), .A(n6323), .ZN(n7350) );
  INV_X1 U5972 ( .A(n8841), .ZN(n7349) );
  INV_X1 U5973 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n5733) );
  AND2_X1 U5974 ( .A1(n8552), .A2(n8548), .ZN(n8545) );
  OR2_X1 U5975 ( .A1(n6494), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6357) );
  NAND2_X1 U5976 ( .A1(n8470), .A2(n8469), .ZN(n8675) );
  AND3_X1 U5977 ( .A1(n6355), .A2(n7095), .A3(n6388), .ZN(n6687) );
  INV_X1 U5978 ( .A(n7099), .ZN(n6495) );
  CLKBUF_X1 U5979 ( .A(n6305), .Z(n6306) );
  INV_X1 U5980 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n6346) );
  OR2_X1 U5981 ( .A1(n6018), .A2(n6017), .ZN(n6038) );
  INV_X1 U5982 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5991) );
  AND2_X1 U5983 ( .A1(n5636), .A2(n5632), .ZN(n5631) );
  INV_X1 U5984 ( .A(n7831), .ZN(n5632) );
  OAI21_X1 U5985 ( .B1(n11023), .B2(n8330), .A(n6973), .ZN(n6974) );
  INV_X1 U5986 ( .A(n8142), .ZN(n8219) );
  NAND2_X1 U5987 ( .A1(n5658), .A2(n5656), .ZN(n9294) );
  NAND2_X1 U5988 ( .A1(n9345), .A2(n9344), .ZN(n5658) );
  INV_X1 U5989 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9317) );
  NOR2_X1 U5990 ( .A1(n8020), .A2(n9317), .ZN(n8021) );
  NOR2_X1 U5991 ( .A1(n7532), .A2(n7531), .ZN(n7533) );
  OAI21_X1 U5992 ( .B1(n10982), .B2(n8330), .A(n6801), .ZN(n6888) );
  OR2_X1 U5993 ( .A1(n7760), .A2(n7979), .ZN(n7803) );
  NAND2_X1 U5994 ( .A1(n5644), .A2(n5642), .ZN(n9364) );
  NOR2_X1 U5995 ( .A1(n5643), .A2(n8210), .ZN(n5642) );
  INV_X1 U5996 ( .A(n9326), .ZN(n5643) );
  AND2_X1 U5997 ( .A1(n6902), .A2(n6901), .ZN(n9394) );
  NOR4_X1 U5998 ( .A1(n9507), .A2(n9506), .A3(n10203), .A4(n9505), .ZN(n9654)
         );
  NAND3_X1 U5999 ( .A1(n9646), .A2(n5559), .A3(n5557), .ZN(n9656) );
  NAND2_X1 U6000 ( .A1(n5558), .A2(n9643), .ZN(n5557) );
  NAND2_X1 U6001 ( .A1(n5263), .A2(n5261), .ZN(n5559) );
  INV_X1 U6002 ( .A(n9650), .ZN(n9651) );
  OR2_X1 U6003 ( .A1(n10614), .A2(n10613), .ZN(n5384) );
  AOI21_X1 U6004 ( .B1(n10620), .B2(P1_REG1_REG_3__SCAN_IN), .A(n10615), .ZN(
        n10951) );
  AND2_X1 U6005 ( .A1(n5384), .A2(n5383), .ZN(n10943) );
  NAND2_X1 U6006 ( .A1(n10620), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n5383) );
  NOR2_X1 U6007 ( .A1(n10943), .A2(n10944), .ZN(n10945) );
  AOI21_X1 U6008 ( .B1(n6869), .B2(P1_REG1_REG_5__SCAN_IN), .A(n10629), .ZN(
        n10645) );
  AOI21_X1 U6009 ( .B1(n10648), .B2(P1_REG1_REG_6__SCAN_IN), .A(n10643), .ZN(
        n10659) );
  NAND2_X1 U6010 ( .A1(n10648), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n5375) );
  INV_X1 U6011 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n7676) );
  AOI21_X1 U6012 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n10677), .A(n10672), .ZN(
        n6874) );
  AOI21_X1 U6013 ( .B1(n10690), .B2(P1_REG1_REG_11__SCAN_IN), .A(n10682), .ZN(
        n7363) );
  AOI21_X1 U6014 ( .B1(n10743), .B2(P1_REG1_REG_13__SCAN_IN), .A(n10735), .ZN(
        n10702) );
  NOR2_X1 U6015 ( .A1(n10738), .A2(n5389), .ZN(n10694) );
  AND2_X1 U6016 ( .A1(n10743), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n5389) );
  NOR2_X1 U6017 ( .A1(n10694), .A2(n10695), .ZN(n10696) );
  NOR2_X1 U6018 ( .A1(n10696), .A2(n5388), .ZN(n10125) );
  AND2_X1 U6019 ( .A1(n10699), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n5388) );
  NAND2_X1 U6020 ( .A1(n10117), .A2(n10116), .ZN(n10139) );
  NAND2_X1 U6021 ( .A1(n10139), .A2(n5252), .ZN(n10141) );
  OR2_X1 U6022 ( .A1(n10140), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n5252) );
  NAND2_X1 U6023 ( .A1(n9408), .A2(n9407), .ZN(n10398) );
  OR2_X1 U6024 ( .A1(n10265), .A2(n5489), .ZN(n10238) );
  AND2_X1 U6025 ( .A1(n9633), .A2(n10187), .ZN(n10236) );
  AND4_X1 U6026 ( .A1(n8343), .A2(n8342), .A3(n8341), .A4(n8340), .ZN(n10269)
         );
  NAND2_X1 U6027 ( .A1(n5312), .A2(n5190), .ZN(n10261) );
  NOR2_X1 U6028 ( .A1(n10442), .A2(n10292), .ZN(n10276) );
  NOR3_X1 U6029 ( .A1(n10379), .A2(n5483), .A3(n10306), .ZN(n10309) );
  INV_X1 U6030 ( .A(n10453), .ZN(n10312) );
  NOR2_X1 U6031 ( .A1(n10379), .A2(n5485), .ZN(n10339) );
  NOR2_X1 U6032 ( .A1(n10379), .A2(n10478), .ZN(n10354) );
  AND2_X1 U6033 ( .A1(n9602), .A2(n9604), .ZN(n10373) );
  AND4_X1 U6034 ( .A1(n8148), .A2(n8147), .A3(n8146), .A4(n8145), .ZN(n9432)
         );
  OAI21_X1 U6035 ( .B1(n5296), .B2(n5295), .A(n5292), .ZN(n8131) );
  NAND2_X1 U6036 ( .A1(n5297), .A2(n5175), .ZN(n5295) );
  AOI21_X1 U6037 ( .B1(n5297), .B2(n5294), .A(n5293), .ZN(n5292) );
  INV_X1 U6038 ( .A(n7991), .ZN(n5296) );
  AND2_X1 U6039 ( .A1(n9595), .A2(n9594), .ZN(n9497) );
  NAND2_X1 U6040 ( .A1(n7637), .A2(n5196), .ZN(n8039) );
  INV_X1 U6041 ( .A(n8121), .ZN(n5486) );
  NAND2_X1 U6042 ( .A1(n7637), .A2(n5170), .ZN(n8003) );
  AND2_X1 U6043 ( .A1(n7637), .A2(n5487), .ZN(n7801) );
  NAND2_X1 U6044 ( .A1(n7753), .A2(n9517), .ZN(n7759) );
  OAI211_X1 U6045 ( .C1(n5715), .C2(n5156), .A(n5189), .B(n5712), .ZN(n7791)
         );
  AND2_X1 U6046 ( .A1(n7533), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n7642) );
  AND4_X1 U6047 ( .A1(n7649), .A2(n7648), .A3(n7647), .A4(n7646), .ZN(n7981)
         );
  NAND2_X1 U6048 ( .A1(n7546), .A2(n7545), .ZN(n7548) );
  INV_X1 U6049 ( .A(n9489), .ZN(n7553) );
  NAND2_X1 U6050 ( .A1(n11113), .A2(n7554), .ZN(n7555) );
  INV_X1 U6051 ( .A(n7637), .ZN(n7638) );
  AND4_X1 U6052 ( .A1(n7538), .A2(n7537), .A3(n7536), .A4(n7535), .ZN(n11108)
         );
  NOR2_X1 U6053 ( .A1(n11059), .A2(n11088), .ZN(n11116) );
  AND2_X1 U6054 ( .A1(n11116), .A2(n11117), .ZN(n11113) );
  INV_X1 U6055 ( .A(n9562), .ZN(n9553) );
  NAND2_X1 U6056 ( .A1(n9560), .A2(n11102), .ZN(n9562) );
  NAND2_X1 U6057 ( .A1(n5549), .A2(n9415), .ZN(n11063) );
  NAND3_X1 U6058 ( .A1(n5492), .A2(n5161), .A3(n11061), .ZN(n11059) );
  AOI21_X1 U6059 ( .B1(n7395), .B2(n9481), .A(n5214), .ZN(n7399) );
  NAND2_X1 U6060 ( .A1(n5161), .A2(n5492), .ZN(n11058) );
  NOR2_X1 U6061 ( .A1(n7199), .A2(n5491), .ZN(n7386) );
  INV_X1 U6062 ( .A(n5493), .ZN(n5491) );
  AND2_X1 U6063 ( .A1(n9544), .A2(n9546), .ZN(n7393) );
  NAND2_X1 U6064 ( .A1(n5492), .A2(n11023), .ZN(n7271) );
  NAND2_X1 U6066 ( .A1(n9663), .A2(n6814), .ZN(n7711) );
  OR2_X1 U6067 ( .A1(n6792), .A2(n9655), .ZN(n10964) );
  AND2_X1 U6068 ( .A1(n8294), .A2(n8293), .ZN(n10448) );
  AND4_X1 U6069 ( .A1(n7765), .A2(n7764), .A3(n7763), .A4(n7762), .ZN(n8119)
         );
  AND4_X1 U6070 ( .A1(n7305), .A2(n7304), .A3(n7303), .A4(n7302), .ZN(n11085)
         );
  INV_X1 U6071 ( .A(n11109), .ZN(n11172) );
  INV_X1 U6072 ( .A(n11107), .ZN(n11169) );
  AND2_X1 U6073 ( .A1(n7169), .A2(n7714), .ZN(n7722) );
  INV_X1 U6074 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n10093) );
  XNOR2_X1 U6075 ( .A(n8453), .B(SI_29_), .ZN(n9405) );
  NAND2_X1 U6076 ( .A1(n6281), .A2(n6280), .ZN(n6406) );
  INV_X1 U6077 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n10089) );
  INV_X1 U6078 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6534) );
  INV_X1 U6079 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6458) );
  INV_X1 U6080 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6467) );
  NAND2_X1 U6081 ( .A1(n6210), .A2(n5848), .ZN(n6220) );
  NAND2_X1 U6082 ( .A1(n5840), .A2(n5839), .ZN(n6200) );
  OAI21_X1 U6083 ( .B1(n6100), .B2(n6099), .A(n5818), .ZN(n6112) );
  AOI21_X1 U6084 ( .B1(n5218), .B2(n5576), .A(n5164), .ZN(n5570) );
  OR2_X1 U6085 ( .A1(n6645), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6721) );
  NAND2_X1 U6086 ( .A1(n5571), .A2(n5573), .ZN(n6052) );
  NAND2_X1 U6087 ( .A1(n5572), .A2(n5577), .ZN(n5571) );
  INV_X1 U6088 ( .A(n6012), .ZN(n5572) );
  OAI211_X1 U6089 ( .C1(n5495), .C2(n5168), .A(n5415), .B(n5414), .ZN(n6541)
         );
  INV_X1 U6090 ( .A(n5416), .ZN(n5415) );
  OAI21_X1 U6091 ( .B1(n5153), .B2(n5168), .A(n5417), .ZN(n5416) );
  NAND2_X1 U6092 ( .A1(n5495), .A2(n5496), .ZN(n5396) );
  NAND2_X1 U6093 ( .A1(n5253), .A2(n5786), .ZN(n5959) );
  OAI21_X1 U6094 ( .B1(n5400), .B2(SI_2_), .A(n5775), .ZN(n5905) );
  NAND2_X1 U6095 ( .A1(n5878), .A2(n5773), .ZN(n5904) );
  MUX2_X1 U6096 ( .A(n6722), .B(n6483), .S(P1_IR_REG_2__SCAN_IN), .Z(n6484) );
  AND2_X1 U6097 ( .A1(n6593), .A2(n6478), .ZN(n6594) );
  AND2_X1 U6098 ( .A1(n7428), .A2(n7427), .ZN(n7430) );
  NAND2_X1 U6099 ( .A1(n8700), .A2(n8702), .ZN(n8701) );
  CLKBUF_X1 U6100 ( .A(n6910), .Z(n6754) );
  CLKBUF_X1 U6101 ( .A(n8722), .Z(n8723) );
  NOR2_X1 U6102 ( .A1(n7896), .A2(n5661), .ZN(n5660) );
  INV_X1 U6103 ( .A(n7894), .ZN(n5661) );
  NAND2_X1 U6104 ( .A1(n8430), .A2(n5676), .ZN(n5674) );
  NAND2_X1 U6105 ( .A1(n6250), .A2(n6249), .ZN(n9162) );
  INV_X1 U6106 ( .A(n8816), .ZN(n8800) );
  NAND2_X1 U6107 ( .A1(n6146), .A2(n6145), .ZN(n8758) );
  NAND2_X1 U6108 ( .A1(n6753), .A2(n6755), .ZN(n6910) );
  NAND2_X1 U6109 ( .A1(n7573), .A2(n7572), .ZN(n7574) );
  AND4_X1 U6110 ( .A1(n6184), .A2(n6183), .A3(n6182), .A4(n6181), .ZN(n9120)
         );
  NAND2_X1 U6111 ( .A1(n8714), .A2(n5668), .ZN(n8769) );
  AND2_X1 U6112 ( .A1(n8714), .A2(n8419), .ZN(n8771) );
  INV_X1 U6113 ( .A(n8830), .ZN(n9118) );
  AND2_X1 U6114 ( .A1(n6642), .A2(n6641), .ZN(n8805) );
  INV_X1 U6115 ( .A(n5672), .ZN(n5671) );
  AOI21_X1 U6116 ( .B1(n5672), .B2(n5677), .A(n5162), .ZN(n5670) );
  AND2_X1 U6117 ( .A1(n5675), .A2(n5673), .ZN(n5672) );
  NAND2_X1 U6118 ( .A1(n5874), .A2(n5873), .ZN(n8806) );
  AND2_X1 U6119 ( .A1(n8403), .A2(n8402), .ZN(n8813) );
  NAND2_X1 U6120 ( .A1(n8403), .A2(n5690), .ZN(n8811) );
  INV_X1 U6121 ( .A(n8808), .ZN(n8810) );
  NAND2_X1 U6122 ( .A1(n6635), .A2(n6634), .ZN(n8819) );
  XNOR2_X1 U6123 ( .A(n6301), .B(P2_IR_REG_22__SCAN_IN), .ZN(n8694) );
  NOR2_X1 U6124 ( .A1(n5753), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n5663) );
  INV_X1 U6125 ( .A(n8664), .ZN(n9000) );
  NAND2_X1 U6126 ( .A1(n5768), .A2(n5767), .ZN(n9025) );
  NAND4_X1 U6127 ( .A1(n6010), .A2(n6009), .A3(n6008), .A4(n6007), .ZN(n8838)
         );
  INV_X2 U6128 ( .A(P2_U3893), .ZN(n8913) );
  NAND2_X1 U6129 ( .A1(n5601), .A2(n5604), .ZN(n6653) );
  INV_X1 U6130 ( .A(n5354), .ZN(n10760) );
  NOR2_X1 U6131 ( .A1(n7218), .A2(n7070), .ZN(n7071) );
  AND2_X1 U6132 ( .A1(n7069), .A2(n7215), .ZN(n7070) );
  INV_X1 U6133 ( .A(n7220), .ZN(n7218) );
  INV_X1 U6134 ( .A(n5356), .ZN(n7069) );
  NAND2_X1 U6135 ( .A1(n7071), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n7222) );
  AOI21_X1 U6136 ( .B1(n7209), .B2(P2_REG1_REG_7__SCAN_IN), .A(n5327), .ZN(
        n7210) );
  AND2_X1 U6137 ( .A1(n5328), .A2(n5355), .ZN(n5327) );
  XNOR2_X1 U6138 ( .A(n8861), .B(n5329), .ZN(n7256) );
  INV_X1 U6139 ( .A(n8920), .ZN(n5329) );
  NAND2_X1 U6140 ( .A1(n7256), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n8862) );
  AND2_X1 U6141 ( .A1(n10789), .A2(n10788), .ZN(n10791) );
  INV_X1 U6142 ( .A(n5612), .ZN(n10805) );
  INV_X1 U6143 ( .A(n8925), .ZN(n5611) );
  CLKBUF_X1 U6144 ( .A(n6094), .Z(n6095) );
  NOR2_X1 U6145 ( .A1(n10872), .A2(n8935), .ZN(n10889) );
  INV_X1 U6146 ( .A(n8974), .ZN(n10905) );
  INV_X1 U6147 ( .A(n10772), .ZN(n10904) );
  MUX2_X1 U6148 ( .A(n6424), .B(n6423), .S(n8669), .Z(n8989) );
  OAI21_X1 U6149 ( .B1(n9074), .B2(n5523), .A(n5521), .ZN(n9042) );
  NAND2_X1 U6150 ( .A1(n5526), .A2(n5527), .ZN(n9053) );
  NAND2_X1 U6151 ( .A1(n9074), .A2(n5528), .ZN(n5526) );
  NAND2_X1 U6152 ( .A1(n6212), .A2(n6211), .ZN(n9175) );
  NAND2_X1 U6153 ( .A1(n9074), .A2(n6336), .ZN(n5529) );
  NAND2_X1 U6154 ( .A1(n5466), .A2(n5464), .ZN(n9083) );
  NAND2_X1 U6155 ( .A1(n5466), .A2(n6335), .ZN(n9081) );
  AND2_X1 U6156 ( .A1(n5459), .A2(n8618), .ZN(n9100) );
  NAND2_X1 U6157 ( .A1(n7959), .A2(n5472), .ZN(n8010) );
  AND2_X1 U6158 ( .A1(n7959), .A2(n8599), .ZN(n8011) );
  NAND2_X1 U6159 ( .A1(n6131), .A2(n6130), .ZN(n8739) );
  OR2_X1 U6160 ( .A1(n9173), .A2(n6372), .ZN(n9040) );
  NAND2_X1 U6161 ( .A1(n5513), .A2(n6050), .ZN(n7667) );
  NAND2_X1 U6162 ( .A1(n7730), .A2(n6049), .ZN(n5513) );
  NOR2_X1 U6163 ( .A1(n8514), .A2(n8513), .ZN(n5451) );
  NAND2_X1 U6164 ( .A1(n5452), .A2(n8518), .ZN(n7600) );
  AND2_X1 U6165 ( .A1(n9145), .A2(n7101), .ZN(n9148) );
  INV_X1 U6166 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9959) );
  INV_X1 U6167 ( .A(n9142), .ZN(n9125) );
  INV_X1 U6168 ( .A(n8689), .ZN(n9214) );
  INV_X1 U6169 ( .A(n8675), .ZN(n9217) );
  NAND2_X1 U6170 ( .A1(n9157), .A2(n5188), .ZN(n9218) );
  NAND2_X1 U6171 ( .A1(n9155), .A2(n9180), .ZN(n5456) );
  NAND2_X1 U6172 ( .A1(n9156), .A2(n9204), .ZN(n5457) );
  INV_X1 U6173 ( .A(n8806), .ZN(n9222) );
  NAND2_X1 U6174 ( .A1(n6178), .A2(n6177), .ZN(n9237) );
  INV_X1 U6175 ( .A(n8786), .ZN(n9242) );
  INV_X1 U6176 ( .A(n8758), .ZN(n9246) );
  INV_X1 U6177 ( .A(n8404), .ZN(n8824) );
  INV_X1 U6178 ( .A(n8162), .ZN(n8519) );
  NAND2_X1 U6179 ( .A1(n6495), .A2(n6494), .ZN(n6505) );
  INV_X1 U6180 ( .A(n5761), .ZN(n8699) );
  XNOR2_X1 U6181 ( .A(n6349), .B(n5694), .ZN(n8079) );
  INV_X1 U6182 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n7859) );
  INV_X1 U6183 ( .A(n8694), .ZN(n7857) );
  INV_X1 U6184 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n6295) );
  NAND2_X1 U6185 ( .A1(n6300), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6296) );
  INV_X1 U6186 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7695) );
  OR2_X1 U6187 ( .A1(n6298), .A2(n6297), .ZN(n6299) );
  INV_X1 U6188 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7655) );
  INV_X1 U6189 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7451) );
  INV_X1 U6190 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7140) );
  INV_X1 U6191 ( .A(n10879), .ZN(n8938) );
  INV_X1 U6192 ( .A(n10863), .ZN(n8933) );
  INV_X1 U6193 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6883) );
  INV_X1 U6194 ( .A(n10812), .ZN(n8927) );
  NAND2_X1 U6195 ( .A1(n5351), .A2(n5349), .ZN(n6613) );
  NAND2_X1 U6196 ( .A1(n5903), .A2(P2_IR_REG_2__SCAN_IN), .ZN(n5351) );
  NOR2_X1 U6197 ( .A1(n5924), .A2(n5350), .ZN(n5349) );
  NAND2_X1 U6198 ( .A1(n5615), .A2(n5880), .ZN(n6661) );
  AOI21_X1 U6199 ( .B1(n5206), .B2(P2_IR_REG_1__SCAN_IN), .A(n5616), .ZN(n5615) );
  NOR2_X1 U6200 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5616) );
  CLKBUF_X1 U6201 ( .A(P2_IR_REG_0__SCAN_IN), .Z(n10749) );
  NAND2_X1 U6202 ( .A1(n5658), .A2(n8249), .ZN(n9297) );
  NAND2_X1 U6203 ( .A1(n8086), .A2(n8085), .ZN(n9322) );
  NAND2_X1 U6204 ( .A1(n8134), .A2(n8133), .ZN(n10488) );
  INV_X1 U6205 ( .A(n5634), .ZN(n7827) );
  AOI21_X1 U6206 ( .B1(n7782), .B2(n5635), .A(n5639), .ZN(n5634) );
  INV_X1 U6207 ( .A(n5641), .ZN(n5635) );
  INV_X1 U6208 ( .A(n5656), .ZN(n5655) );
  AND2_X1 U6209 ( .A1(n8287), .A2(n5653), .ZN(n5652) );
  INV_X1 U6210 ( .A(n9391), .ZN(n9367) );
  AND4_X1 U6211 ( .A1(n7343), .A2(n7342), .A3(n7341), .A4(n7340), .ZN(n11110)
         );
  INV_X1 U6212 ( .A(n9402), .ZN(n9376) );
  AND4_X1 U6213 ( .A1(n6527), .A2(n6526), .A3(n6525), .A4(n6524), .ZN(n10378)
         );
  OR2_X1 U6214 ( .A1(n6966), .A2(n6897), .ZN(n6900) );
  OR2_X1 U6215 ( .A1(n6983), .A2(n6763), .ZN(n6764) );
  OR2_X1 U6216 ( .A1(n6966), .A2(n6761), .ZN(n6767) );
  NOR2_X1 U6217 ( .A1(n10669), .A2(n5226), .ZN(n6855) );
  AOI22_X1 U6218 ( .A1(n7356), .A2(n9676), .B1(P1_REG2_REG_10__SCAN_IN), .B2(
        n7525), .ZN(n10687) );
  NOR2_X1 U6219 ( .A1(n10687), .A2(n10686), .ZN(n10685) );
  NOR2_X1 U6220 ( .A1(n10685), .A2(n5386), .ZN(n7358) );
  AND2_X1 U6221 ( .A1(n10690), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n5386) );
  NAND2_X1 U6222 ( .A1(n7358), .A2(n7359), .ZN(n10121) );
  AND2_X1 U6223 ( .A1(n6540), .A2(n6858), .ZN(n10942) );
  XNOR2_X1 U6224 ( .A(n10125), .B(n5387), .ZN(n10715) );
  NAND2_X1 U6225 ( .A1(n6860), .A2(n6859), .ZN(n10958) );
  NAND2_X1 U6226 ( .A1(n5450), .A2(n5131), .ZN(n10392) );
  XNOR2_X1 U6227 ( .A(n10174), .B(n10393), .ZN(n5450) );
  NAND2_X1 U6228 ( .A1(n5598), .A2(n9447), .ZN(n10176) );
  NAND2_X1 U6229 ( .A1(n9446), .A2(n8029), .ZN(n5598) );
  AOI21_X1 U6230 ( .B1(n10218), .B2(n10220), .A(n10189), .ZN(n5334) );
  NAND2_X1 U6231 ( .A1(n10222), .A2(n10202), .ZN(n10205) );
  NAND2_X1 U6232 ( .A1(n8356), .A2(n8355), .ZN(n10244) );
  NOR2_X1 U6233 ( .A1(n5282), .A2(n5280), .ZN(n10250) );
  INV_X1 U6234 ( .A(n5335), .ZN(n5280) );
  NOR2_X1 U6235 ( .A1(n5337), .A2(n10305), .ZN(n5282) );
  INV_X1 U6236 ( .A(n10435), .ZN(n10271) );
  NAND2_X1 U6237 ( .A1(n10282), .A2(n10184), .ZN(n10263) );
  OAI21_X1 U6238 ( .B1(n10320), .B2(n5701), .A(n5699), .ZN(n10275) );
  INV_X1 U6239 ( .A(n10448), .ZN(n10299) );
  OAI21_X1 U6240 ( .B1(n10305), .B2(n10304), .A(n10180), .ZN(n10291) );
  NAND2_X1 U6241 ( .A1(n5704), .A2(n5702), .ZN(n10289) );
  INV_X1 U6242 ( .A(n5706), .ZN(n5702) );
  NAND2_X1 U6243 ( .A1(n10320), .A2(n5708), .ZN(n5704) );
  AOI21_X1 U6244 ( .B1(n10320), .B2(n10321), .A(n5705), .ZN(n10303) );
  INV_X1 U6245 ( .A(n5707), .ZN(n5705) );
  INV_X1 U6246 ( .A(n10466), .ZN(n10331) );
  AOI21_X1 U6247 ( .B1(n10361), .B2(n5546), .A(n9456), .ZN(n10322) );
  AND2_X1 U6248 ( .A1(n8235), .A2(n8234), .ZN(n10341) );
  NAND2_X1 U6249 ( .A1(n10361), .A2(n9455), .ZN(n10347) );
  AOI21_X1 U6250 ( .B1(n10353), .B2(n10193), .A(n5149), .ZN(n10338) );
  NAND2_X1 U6251 ( .A1(n8205), .A2(n8204), .ZN(n10483) );
  NAND2_X1 U6252 ( .A1(n9587), .A2(n8028), .ZN(n8033) );
  OAI21_X1 U6253 ( .B1(n7991), .B2(n5298), .A(n5297), .ZN(n8083) );
  INV_X1 U6254 ( .A(n5299), .ZN(n8037) );
  AOI21_X1 U6255 ( .B1(n7991), .B2(n5720), .A(n5301), .ZN(n5299) );
  NAND2_X1 U6256 ( .A1(n7795), .A2(n7794), .ZN(n7992) );
  NAND2_X1 U6257 ( .A1(n7756), .A2(n7755), .ZN(n7929) );
  OR2_X1 U6258 ( .A1(n7754), .A2(n6959), .ZN(n7756) );
  NAND2_X1 U6259 ( .A1(n5715), .A2(n5710), .ZN(n7768) );
  INV_X1 U6260 ( .A(n5714), .ZN(n5711) );
  OAI21_X1 U6261 ( .B1(n7610), .B2(n9569), .A(n5719), .ZN(n7633) );
  AND2_X1 U6262 ( .A1(n10367), .A2(n7189), .ZN(n11124) );
  INV_X1 U6263 ( .A(n11124), .ZN(n10387) );
  OR2_X1 U6264 ( .A1(n6968), .A2(n7022), .ZN(n7028) );
  INV_X1 U6265 ( .A(n11128), .ZN(n10333) );
  AND2_X1 U6266 ( .A1(n10367), .A2(n7174), .ZN(n11129) );
  AND2_X2 U6267 ( .A1(n7721), .A2(n7715), .ZN(n11202) );
  NAND2_X1 U6268 ( .A1(n10392), .A2(n5448), .ZN(n10491) );
  INV_X1 U6269 ( .A(n5449), .ZN(n5448) );
  OAI21_X1 U6270 ( .B1(n10393), .B2(n11195), .A(n10394), .ZN(n5449) );
  NAND2_X1 U6271 ( .A1(n5198), .A2(n5288), .ZN(n10494) );
  AND2_X2 U6272 ( .A1(n7722), .A2(n7721), .ZN(n11206) );
  AND2_X1 U6273 ( .A1(n6770), .A2(n6769), .ZN(n10507) );
  XNOR2_X1 U6274 ( .A(n8461), .B(n8460), .ZN(n9452) );
  NAND2_X1 U6275 ( .A1(n8467), .A2(n8457), .ZN(n8461) );
  XNOR2_X1 U6276 ( .A(n6406), .B(n6405), .ZN(n10519) );
  INV_X1 U6277 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n10013) );
  INV_X1 U6278 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n9801) );
  NAND2_X1 U6279 ( .A1(n6537), .A2(n6465), .ZN(n6466) );
  INV_X1 U6280 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n9805) );
  INV_X1 U6281 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10021) );
  INV_X1 U6282 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7657) );
  INV_X1 U6283 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n10025) );
  NAND2_X1 U6284 ( .A1(n5578), .A2(n5577), .ZN(n6037) );
  NAND2_X1 U6285 ( .A1(n5578), .A2(n5579), .ZN(n6035) );
  AND2_X1 U6286 ( .A1(n5134), .A2(P1_U3086), .ZN(n7489) );
  OAI21_X1 U6287 ( .B1(n5974), .B2(n5499), .A(n5498), .ZN(n5990) );
  NOR2_X1 U6288 ( .A1(n5989), .A2(n5499), .ZN(n5347) );
  INV_X1 U6289 ( .A(n5380), .ZN(n5379) );
  INV_X1 U6290 ( .A(n6481), .ZN(n5382) );
  OAI21_X1 U6291 ( .B1(P1_IR_REG_31__SCAN_IN), .B2(P1_IR_REG_1__SCAN_IN), .A(
        n5381), .ZN(n5380) );
  NAND2_X1 U6292 ( .A1(n5771), .A2(n5773), .ZN(n5876) );
  OAI211_X1 U6293 ( .C1(n8949), .C2(n8974), .A(n5373), .B(n5372), .ZN(P2_U3200) );
  OR2_X1 U6294 ( .A1(n8943), .A2(n10910), .ZN(n5372) );
  AOI21_X1 U6295 ( .B1(n8947), .B2(n8948), .A(n5374), .ZN(n5373) );
  OAI21_X1 U6296 ( .B1(n5332), .B2(n8974), .A(n5208), .ZN(P2_U3201) );
  XNOR2_X1 U6297 ( .A(n8952), .B(n8967), .ZN(n5332) );
  AOI21_X1 U6298 ( .B1(n8665), .B2(n6400), .A(n6399), .ZN(n6401) );
  NAND2_X1 U6299 ( .A1(n5404), .A2(n5403), .ZN(P2_U3486) );
  NAND2_X1 U6300 ( .A1(n9210), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n5403) );
  NAND2_X1 U6301 ( .A1(n9218), .A2(n9206), .ZN(n5404) );
  AOI21_X1 U6302 ( .B1(n6440), .B2(n6446), .A(n6445), .ZN(n6447) );
  NOR2_X1 U6303 ( .A1(n11186), .A2(n6444), .ZN(n6445) );
  INV_X1 U6304 ( .A(n5453), .ZN(P2_U3454) );
  AOI21_X1 U6305 ( .B1(n9218), .B2(n11186), .A(n5454), .ZN(n5453) );
  NOR2_X1 U6306 ( .A1(n11186), .A2(n5455), .ZN(n5454) );
  INV_X1 U6307 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n5455) );
  XNOR2_X1 U6308 ( .A(n5629), .B(n8394), .ZN(n8399) );
  AND2_X1 U6309 ( .A1(n7019), .A2(n7018), .ZN(n5624) );
  NAND2_X1 U6310 ( .A1(n5625), .A2(n6943), .ZN(n7054) );
  NAND2_X1 U6311 ( .A1(n5552), .A2(n5551), .ZN(P1_U3242) );
  OR2_X1 U6312 ( .A1(n9668), .A2(n9667), .ZN(n5551) );
  OR2_X1 U6313 ( .A1(n10729), .A2(n5248), .ZN(P1_U3261) );
  OR2_X1 U6314 ( .A1(n10728), .A2(n5249), .ZN(n5248) );
  INV_X1 U6315 ( .A(n5250), .ZN(n5249) );
  INV_X1 U6316 ( .A(n5445), .ZN(P1_U3521) );
  AOI21_X1 U6317 ( .B1(n10491), .B2(n11206), .A(n5446), .ZN(n5445) );
  NOR2_X1 U6318 ( .A1(n11206), .A2(n5447), .ZN(n5446) );
  INV_X1 U6319 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n5447) );
  INV_X1 U6320 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7162) );
  NOR2_X1 U6321 ( .A1(n6034), .A2(n5804), .ZN(n5577) );
  AND2_X1 U6322 ( .A1(n8429), .A2(n9065), .ZN(n5148) );
  INV_X1 U6323 ( .A(n5577), .ZN(n5576) );
  AND2_X1 U6324 ( .A1(n10355), .A2(n10349), .ZN(n5149) );
  AND2_X1 U6325 ( .A1(n9155), .A2(n8827), .ZN(n5150) );
  NAND2_X2 U6326 ( .A1(n5133), .A2(n6884), .ZN(n6959) );
  OR2_X1 U6327 ( .A1(n7854), .A2(n8835), .ZN(n5151) );
  AND2_X1 U6328 ( .A1(n5582), .A2(n6155), .ZN(n5152) );
  AND2_X1 U6329 ( .A1(n5496), .A2(n5420), .ZN(n5153) );
  NAND2_X1 U6330 ( .A1(n9048), .A2(n8651), .ZN(n5154) );
  AND4_X1 U6331 ( .A1(n6053), .A2(n6015), .A3(n6013), .A4(n6056), .ZN(n5155)
         );
  NOR2_X1 U6332 ( .A1(n7874), .A2(n11146), .ZN(n5156) );
  NOR2_X1 U6333 ( .A1(n6470), .A2(P1_IR_REG_25__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U6334 ( .A1(n9617), .A2(n10180), .ZN(n10304) );
  INV_X1 U6335 ( .A(n7698), .ZN(n5511) );
  NAND2_X1 U6336 ( .A1(n7628), .A2(n7570), .ZN(n8518) );
  INV_X1 U6337 ( .A(n9093), .ZN(n5463) );
  INV_X1 U6338 ( .A(n7238), .ZN(n7234) );
  AND2_X1 U6339 ( .A1(n5506), .A2(n5502), .ZN(n5158) );
  NAND2_X1 U6340 ( .A1(n10341), .A2(n10462), .ZN(n5159) );
  INV_X1 U6341 ( .A(n5339), .ZN(n5337) );
  NOR2_X1 U6342 ( .A1(n5537), .A2(n5187), .ZN(n5339) );
  AOI21_X1 U6343 ( .B1(n5429), .B2(n9080), .A(n8640), .ZN(n5428) );
  AND2_X1 U6344 ( .A1(n5493), .A2(n7385), .ZN(n5161) );
  AND2_X1 U6345 ( .A1(n8433), .A2(n9044), .ZN(n5162) );
  NAND2_X1 U6346 ( .A1(n5592), .A2(n5228), .ZN(n5163) );
  NOR2_X1 U6347 ( .A1(n5809), .A2(SI_11_), .ZN(n5164) );
  AND3_X1 U6348 ( .A1(n5691), .A2(n5870), .A3(n5868), .ZN(n5165) );
  NAND2_X1 U6349 ( .A1(n5756), .A2(n5694), .ZN(n5693) );
  INV_X1 U6350 ( .A(n5693), .ZN(n5691) );
  AND2_X1 U6351 ( .A1(n7576), .A2(n7572), .ZN(n5166) );
  NAND2_X1 U6352 ( .A1(n6910), .A2(n6909), .ZN(n6911) );
  INV_X1 U6353 ( .A(n10829), .ZN(n5366) );
  INV_X1 U6354 ( .A(n7215), .ZN(n5355) );
  INV_X1 U6355 ( .A(n6983), .ZN(n6836) );
  INV_X1 U6356 ( .A(n7077), .ZN(n5358) );
  NAND2_X1 U6357 ( .A1(n10363), .A2(n10362), .ZN(n10361) );
  AND2_X1 U6358 ( .A1(n6380), .A2(n5755), .ZN(n6345) );
  NAND2_X1 U6359 ( .A1(n6481), .A2(n6450), .ZN(n6482) );
  NAND2_X1 U6360 ( .A1(n5721), .A2(n5157), .ZN(n6515) );
  OR2_X1 U6361 ( .A1(n10265), .A2(n10257), .ZN(n5167) );
  INV_X1 U6362 ( .A(n6651), .ZN(n5602) );
  OR2_X1 U6363 ( .A1(n6011), .A2(n5418), .ZN(n5168) );
  NOR2_X1 U6364 ( .A1(n7664), .A2(n8837), .ZN(n5169) );
  AND2_X1 U6365 ( .A1(n11175), .A2(n5487), .ZN(n5170) );
  AND2_X1 U6366 ( .A1(n9375), .A2(n5723), .ZN(n5171) );
  AND2_X1 U6367 ( .A1(n9523), .A2(n9526), .ZN(n9569) );
  OR2_X1 U6368 ( .A1(n9179), .A2(n9064), .ZN(n5172) );
  AND4_X1 U6369 ( .A1(n6016), .A2(n5747), .A3(n5923), .A4(n6014), .ZN(n5173)
         );
  OAI21_X1 U6370 ( .B1(n8430), .B2(n5671), .A(n5670), .ZN(n8798) );
  OR2_X1 U6371 ( .A1(n5143), .A2(n7202), .ZN(n5174) );
  NAND2_X1 U6372 ( .A1(n5674), .A2(n5675), .ZN(n8731) );
  OR2_X1 U6373 ( .A1(n9400), .A2(n9671), .ZN(n5175) );
  AOI21_X1 U6374 ( .B1(n10248), .B2(n10249), .A(n10198), .ZN(n10234) );
  AND2_X1 U6375 ( .A1(n7990), .A2(n9575), .ZN(n5176) );
  OR2_X1 U6376 ( .A1(n10277), .A2(n10297), .ZN(n5177) );
  XNOR2_X1 U6377 ( .A(n8430), .B(n8429), .ZN(n8707) );
  NAND2_X1 U6378 ( .A1(n8217), .A2(n8216), .ZN(n10478) );
  OR2_X1 U6379 ( .A1(n10829), .A2(n8928), .ZN(n5178) );
  AND2_X1 U6380 ( .A1(n5649), .A2(n5648), .ZN(n5179) );
  AND2_X1 U6381 ( .A1(n9636), .A2(n10188), .ZN(n10220) );
  INV_X1 U6382 ( .A(n10220), .ZN(n5289) );
  NAND2_X1 U6383 ( .A1(n7636), .A2(n7635), .ZN(n7874) );
  INV_X1 U6384 ( .A(n8594), .ZN(n6110) );
  NAND2_X1 U6385 ( .A1(n5761), .A2(n9260), .ZN(n5915) );
  INV_X1 U6386 ( .A(n5915), .ZN(n5882) );
  NAND2_X1 U6387 ( .A1(n8334), .A2(n8333), .ZN(n10257) );
  INV_X1 U6388 ( .A(n10257), .ZN(n5490) );
  AND2_X1 U6389 ( .A1(n9621), .A2(n9640), .ZN(n5180) );
  NAND2_X1 U6390 ( .A1(n9009), .A2(n9015), .ZN(n5181) );
  AOI21_X1 U6391 ( .B1(n8798), .B2(n8799), .A(n8435), .ZN(n8700) );
  AND2_X1 U6392 ( .A1(n7854), .A2(n8835), .ZN(n5182) );
  AND2_X1 U6393 ( .A1(n5376), .A2(n5375), .ZN(n5183) );
  NAND2_X1 U6394 ( .A1(n8716), .A2(n8715), .ZN(n8714) );
  NAND2_X1 U6395 ( .A1(n6481), .A2(n5533), .ZN(n6489) );
  AND2_X1 U6396 ( .A1(n8646), .A2(n8645), .ZN(n9058) );
  NAND2_X1 U6397 ( .A1(n5666), .A2(n5749), .ZN(n6101) );
  INV_X1 U6398 ( .A(n9514), .ZN(n5542) );
  AND2_X1 U6399 ( .A1(n10220), .A2(n9634), .ZN(n5184) );
  NOR2_X1 U6400 ( .A1(n7826), .A2(n5639), .ZN(n5185) );
  NOR2_X1 U6401 ( .A1(n8115), .A2(n8817), .ZN(n5186) );
  AND2_X1 U6402 ( .A1(n5341), .A2(n5343), .ZN(n5187) );
  INV_X1 U6403 ( .A(n5258), .ZN(n5875) );
  OAI211_X1 U6404 ( .C1(n5134), .C2(P2_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n5259), .ZN(n5258) );
  AND2_X1 U6405 ( .A1(n5457), .A2(n5456), .ZN(n5188) );
  INV_X1 U6406 ( .A(n8514), .ZN(n6031) );
  NAND2_X1 U6407 ( .A1(n8516), .A2(n8522), .ZN(n8514) );
  OR2_X1 U6408 ( .A1(n7889), .A2(n7872), .ZN(n5189) );
  AND2_X1 U6409 ( .A1(n5698), .A2(n5709), .ZN(n5190) );
  AND2_X1 U6410 ( .A1(n11163), .A2(n7981), .ZN(n5191) );
  INV_X1 U6411 ( .A(n5677), .ZN(n5676) );
  NAND2_X1 U6412 ( .A1(n5682), .A2(n5680), .ZN(n5677) );
  AND2_X1 U6413 ( .A1(n6912), .A2(n6909), .ZN(n5192) );
  AND2_X1 U6414 ( .A1(n5289), .A2(n10200), .ZN(n5193) );
  AND2_X1 U6415 ( .A1(n10176), .A2(n9639), .ZN(n5194) );
  INV_X1 U6416 ( .A(n5430), .ZN(n5429) );
  NAND2_X1 U6417 ( .A1(n5431), .A2(n5434), .ZN(n5430) );
  OR2_X1 U6418 ( .A1(n5358), .A2(n7078), .ZN(n5195) );
  OR2_X1 U6419 ( .A1(n10442), .A2(n10297), .ZN(n10184) );
  INV_X1 U6420 ( .A(n10184), .ZN(n5539) );
  AND2_X1 U6421 ( .A1(n5170), .A2(n5486), .ZN(n5196) );
  AND2_X1 U6422 ( .A1(n10282), .A2(n5538), .ZN(n5197) );
  INV_X1 U6423 ( .A(n5799), .ZN(n5497) );
  NAND2_X1 U6424 ( .A1(n5796), .A2(SI_7_), .ZN(n5799) );
  AND2_X1 U6425 ( .A1(n10415), .A2(n10413), .ZN(n5198) );
  NAND2_X1 U6426 ( .A1(n7616), .A2(n5996), .ZN(n8560) );
  INV_X1 U6427 ( .A(n8560), .ZN(n5397) );
  INV_X1 U6428 ( .A(n8669), .ZN(n5509) );
  OR2_X1 U6429 ( .A1(n5358), .A2(n5357), .ZN(n5199) );
  INV_X1 U6430 ( .A(n5804), .ZN(n5579) );
  INV_X1 U6431 ( .A(n10319), .ZN(n10321) );
  AND2_X1 U6432 ( .A1(n5542), .A2(n9516), .ZN(n10319) );
  AND2_X1 U6433 ( .A1(n10179), .A2(n5281), .ZN(n5200) );
  OR2_X1 U6434 ( .A1(n5560), .A2(n5194), .ZN(n5201) );
  AND2_X1 U6435 ( .A1(n9523), .A2(n9535), .ZN(n5202) );
  NAND2_X1 U6436 ( .A1(n9039), .A2(n9054), .ZN(n5203) );
  OR2_X1 U6437 ( .A1(n6471), .A2(n6470), .ZN(n5204) );
  NAND2_X1 U6438 ( .A1(n5666), .A2(n5663), .ZN(n5205) );
  AND2_X1 U6439 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(n10749), .ZN(n5206) );
  NOR2_X1 U6440 ( .A1(n10473), .A2(n10462), .ZN(n5207) );
  AND2_X1 U6441 ( .A1(n5620), .A2(n5617), .ZN(n5208) );
  INV_X1 U6442 ( .A(n5669), .ZN(n5668) );
  NAND2_X1 U6443 ( .A1(n8419), .A2(n8770), .ZN(n5669) );
  AND2_X1 U6444 ( .A1(n9000), .A2(n8665), .ZN(n5209) );
  INV_X1 U6445 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n10083) );
  INV_X1 U6446 ( .A(n5465), .ZN(n5464) );
  NAND2_X1 U6447 ( .A1(n5435), .A2(n6335), .ZN(n5465) );
  AND2_X1 U6448 ( .A1(n5172), .A2(n6336), .ZN(n9080) );
  INV_X1 U6449 ( .A(n9080), .ZN(n5435) );
  INV_X1 U6450 ( .A(n8640), .ZN(n9067) );
  XNOR2_X1 U6451 ( .A(n7289), .B(n7288), .ZN(n7015) );
  INV_X1 U6452 ( .A(n7015), .ZN(n7016) );
  OR2_X1 U6453 ( .A1(n6338), .A2(n6337), .ZN(n5210) );
  INV_X1 U6454 ( .A(n7385), .ZN(n11048) );
  AND3_X1 U6455 ( .A1(n7287), .A2(n7286), .A3(n7285), .ZN(n7385) );
  OR2_X1 U6456 ( .A1(n8667), .A2(n5441), .ZN(n5211) );
  INV_X1 U6457 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6462) );
  AND2_X1 U6458 ( .A1(n9065), .A2(n5530), .ZN(n5212) );
  NOR2_X1 U6459 ( .A1(n10448), .A2(n10312), .ZN(n5213) );
  NAND2_X1 U6460 ( .A1(n10271), .A2(n10196), .ZN(n10185) );
  AND2_X1 U6461 ( .A1(n11046), .A2(n7394), .ZN(n5214) );
  INV_X1 U6462 ( .A(n5726), .ZN(n5648) );
  NAND2_X1 U6463 ( .A1(n6218), .A2(n5172), .ZN(n5215) );
  NAND2_X1 U6464 ( .A1(n9494), .A2(n5300), .ZN(n5216) );
  AND2_X1 U6465 ( .A1(n9179), .A2(n9091), .ZN(n5217) );
  XNOR2_X1 U6466 ( .A(n5803), .B(n9928), .ZN(n6011) );
  INV_X1 U6467 ( .A(n6011), .ZN(n5575) );
  AND2_X1 U6468 ( .A1(n5573), .A2(n5291), .ZN(n5218) );
  AND3_X1 U6469 ( .A1(n5496), .A2(n5420), .A3(n6011), .ZN(n5219) );
  AND2_X1 U6470 ( .A1(n5529), .A2(n5172), .ZN(n5220) );
  AND2_X1 U6471 ( .A1(n5699), .A2(n5177), .ZN(n5221) );
  NOR2_X1 U6472 ( .A1(n10889), .A2(n10888), .ZN(n5222) );
  AND2_X1 U6473 ( .A1(n9601), .A2(n9431), .ZN(n10191) );
  NOR2_X1 U6474 ( .A1(P1_IR_REG_28__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), .ZN(
        n5223) );
  AND2_X1 U6475 ( .A1(n5650), .A2(n5651), .ZN(n5224) );
  AND2_X1 U6476 ( .A1(n5608), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5225) );
  INV_X1 U6477 ( .A(n8036), .ZN(n5302) );
  AND2_X1 U6478 ( .A1(n8121), .A2(n11170), .ZN(n8036) );
  INV_X1 U6479 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5748) );
  INV_X1 U6480 ( .A(n8432), .ZN(n5682) );
  AND2_X1 U6481 ( .A1(n8431), .A2(n8709), .ZN(n8432) );
  INV_X1 U6482 ( .A(n5685), .ZN(n5684) );
  NAND2_X1 U6483 ( .A1(n7429), .A2(n7427), .ZN(n5685) );
  INV_X1 U6484 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5870) );
  BUF_X1 U6485 ( .A(n5916), .Z(n6149) );
  NAND2_X2 U6486 ( .A1(n6676), .A2(n8694), .ZN(n8676) );
  INV_X1 U6487 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n5597) );
  AND2_X1 U6488 ( .A1(n10677), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n5226) );
  INV_X1 U6489 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n5399) );
  AND2_X1 U6490 ( .A1(n7401), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n5227) );
  INV_X1 U6491 ( .A(n7219), .ZN(n7257) );
  NAND2_X1 U6492 ( .A1(n5843), .A2(SI_21_), .ZN(n5228) );
  NAND2_X1 U6493 ( .A1(n6082), .A2(n6081), .ZN(n7818) );
  NAND2_X1 U6494 ( .A1(n6333), .A2(n6332), .ZN(n9122) );
  INV_X1 U6495 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5694) );
  INV_X1 U6496 ( .A(n5795), .ZN(n5499) );
  NAND2_X1 U6497 ( .A1(n6258), .A2(n6257), .ZN(n8828) );
  INV_X1 U6498 ( .A(n8828), .ZN(n9044) );
  NAND2_X1 U6499 ( .A1(n5688), .A2(n5686), .ZN(n8740) );
  NAND2_X1 U6500 ( .A1(n5662), .A2(n7894), .ZN(n7895) );
  OR2_X1 U6501 ( .A1(n10379), .A2(n5483), .ZN(n5229) );
  NAND2_X1 U6502 ( .A1(n5392), .A2(n5395), .ZN(n7915) );
  AND2_X1 U6503 ( .A1(n8420), .A2(n9077), .ZN(n5230) );
  INV_X1 U6504 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9253) );
  NAND2_X1 U6505 ( .A1(n8376), .A2(n8375), .ZN(n10412) );
  AND2_X1 U6506 ( .A1(n5612), .A2(n5611), .ZN(n5231) );
  INV_X1 U6507 ( .A(n5546), .ZN(n5545) );
  AND2_X1 U6508 ( .A1(n5847), .A2(n5228), .ZN(n5232) );
  NAND2_X1 U6509 ( .A1(n8106), .A2(n8105), .ZN(n8403) );
  INV_X1 U6510 ( .A(n8665), .ZN(n8993) );
  NAND2_X1 U6511 ( .A1(n6283), .A2(n6282), .ZN(n8665) );
  AND2_X1 U6512 ( .A1(n5820), .A2(SI_15_), .ZN(n5233) );
  AND2_X1 U6513 ( .A1(n5831), .A2(SI_18_), .ZN(n5234) );
  INV_X1 U6514 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5749) );
  AND2_X1 U6515 ( .A1(n7986), .A2(n9575), .ZN(n5235) );
  OR2_X1 U6516 ( .A1(n7219), .A2(n5607), .ZN(n5236) );
  AND2_X1 U6517 ( .A1(n8927), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5237) );
  NAND2_X1 U6518 ( .A1(n7428), .A2(n5684), .ZN(n7503) );
  AND2_X1 U6519 ( .A1(n7637), .A2(n7889), .ZN(n5238) );
  NOR2_X1 U6520 ( .A1(n5139), .A2(n10013), .ZN(n5239) );
  INV_X1 U6521 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n5322) );
  OAI21_X1 U6522 ( .B1(n7135), .B2(n5948), .A(n5947), .ZN(n7441) );
  AND2_X1 U6523 ( .A1(n7459), .A2(n7458), .ZN(n5240) );
  INV_X1 U6524 ( .A(n10718), .ZN(n5387) );
  NAND2_X1 U6525 ( .A1(n6910), .A2(n5192), .ZN(n7035) );
  INV_X1 U6526 ( .A(n5720), .ZN(n5303) );
  OR2_X1 U6527 ( .A1(n7992), .A2(n9672), .ZN(n5720) );
  NAND2_X1 U6528 ( .A1(n7235), .A2(n7234), .ZN(n7428) );
  OR2_X1 U6529 ( .A1(n10981), .A2(n7198), .ZN(n7199) );
  INV_X1 U6530 ( .A(n7199), .ZN(n5492) );
  INV_X1 U6531 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n5607) );
  OR2_X1 U6532 ( .A1(n5237), .A2(n5366), .ZN(n5241) );
  INV_X1 U6533 ( .A(n8525), .ZN(n6676) );
  AND2_X1 U6534 ( .A1(n8938), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5242) );
  OAI22_X1 U6535 ( .A1(n10985), .A2(n10980), .B1(n9409), .B2(n11007), .ZN(
        n7197) );
  AND2_X1 U6536 ( .A1(n7501), .A2(n7500), .ZN(n5243) );
  AND2_X1 U6537 ( .A1(n5605), .A2(n5606), .ZN(n5244) );
  OR2_X1 U6538 ( .A1(n10625), .A2(n10626), .ZN(n5378) );
  AND2_X1 U6539 ( .A1(n5599), .A2(n5604), .ZN(n5245) );
  NAND2_X1 U6540 ( .A1(n7675), .A2(n10163), .ZN(n9666) );
  INV_X1 U6541 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n5357) );
  INV_X1 U6542 ( .A(n5989), .ZN(n5314) );
  NAND2_X1 U6543 ( .A1(n5974), .A2(n5498), .ZN(n5495) );
  NAND2_X1 U6544 ( .A1(n10374), .A2(n10373), .ZN(n10372) );
  OAI21_X1 U6545 ( .B1(n5335), .B2(n10249), .A(n5278), .ZN(n10237) );
  OAI21_X1 U6546 ( .B1(n7986), .B2(n5346), .A(n5344), .ZN(n8087) );
  OAI21_X1 U6547 ( .B1(n5176), .B2(n5346), .A(n9496), .ZN(n5345) );
  XNOR2_X1 U6548 ( .A(n5334), .B(n10203), .ZN(n10404) );
  INV_X2 U6549 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n5247) );
  NAND2_X2 U6550 ( .A1(n8232), .A2(n8231), .ZN(n9345) );
  NAND2_X2 U6551 ( .A1(n8291), .A2(n8290), .ZN(n9352) );
  INV_X1 U6552 ( .A(n7014), .ZN(n7017) );
  NAND2_X1 U6553 ( .A1(n7683), .A2(n7682), .ZN(n7782) );
  NAND2_X1 U6554 ( .A1(n7017), .A2(n7016), .ZN(n7018) );
  NAND2_X2 U6555 ( .A1(n9302), .A2(n9303), .ZN(n9301) );
  OR2_X1 U6556 ( .A1(n8330), .A2(n7394), .ZN(n7005) );
  NAND2_X1 U6557 ( .A1(n7019), .A2(n5623), .ZN(n7296) );
  NAND2_X1 U6558 ( .A1(n5944), .A2(n5253), .ZN(n6999) );
  NAND2_X1 U6559 ( .A1(n5943), .A2(n5942), .ZN(n5253) );
  NAND2_X1 U6560 ( .A1(n5976), .A2(n5347), .ZN(n5257) );
  NAND3_X1 U6561 ( .A1(n5773), .A2(n5771), .A3(n5875), .ZN(n5878) );
  NAND2_X1 U6562 ( .A1(n5260), .A2(n9940), .ZN(n5771) );
  NAND2_X1 U6563 ( .A1(n10237), .A2(n10236), .ZN(n10235) );
  MUX2_X1 U6564 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .S(n6884), .Z(n5803) );
  OR2_X1 U6565 ( .A1(n10353), .A2(n5307), .ZN(n5306) );
  NAND3_X1 U6566 ( .A1(n5306), .A2(n5221), .A3(n5304), .ZN(n5312) );
  AOI21_X1 U6567 ( .B1(n5318), .B2(n5795), .A(n5314), .ZN(n5498) );
  NAND3_X1 U6568 ( .A1(n5324), .A2(n5323), .A3(P2_DATAO_REG_6__SCAN_IN), .ZN(
        n5319) );
  INV_X1 U6569 ( .A(n5323), .ZN(n5321) );
  AND2_X2 U6570 ( .A1(n5353), .A2(n5352), .ZN(n5879) );
  INV_X1 U6571 ( .A(n10757), .ZN(n5359) );
  NAND2_X1 U6572 ( .A1(n10758), .A2(n10756), .ZN(n5360) );
  NOR2_X1 U6573 ( .A1(n10822), .A2(n5237), .ZN(n8928) );
  NAND2_X1 U6574 ( .A1(n5361), .A2(n5364), .ZN(n5367) );
  NAND3_X1 U6575 ( .A1(n5364), .A2(n5365), .A3(n5363), .ZN(n10839) );
  INV_X1 U6576 ( .A(n5367), .ZN(n10838) );
  AOI21_X1 U6577 ( .B1(n8935), .B2(n5371), .A(n5242), .ZN(n5369) );
  NAND2_X1 U6578 ( .A1(n10872), .A2(n5371), .ZN(n5370) );
  NAND3_X1 U6579 ( .A1(n8946), .A2(n8944), .A3(n8945), .ZN(n5374) );
  NAND3_X1 U6580 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_1__SCAN_IN), .A3(
        P1_IR_REG_0__SCAN_IN), .ZN(n5381) );
  NAND2_X1 U6581 ( .A1(n6082), .A2(n5393), .ZN(n5392) );
  NAND2_X1 U6582 ( .A1(n8515), .A2(n8518), .ZN(n6029) );
  NAND2_X1 U6583 ( .A1(n5495), .A2(n5219), .ZN(n5414) );
  NAND2_X1 U6584 ( .A1(n6541), .A2(n8468), .ZN(n6021) );
  NAND2_X1 U6585 ( .A1(n5421), .A2(n5422), .ZN(n8655) );
  NAND2_X1 U6586 ( .A1(n8638), .A2(n5423), .ZN(n5421) );
  NAND2_X1 U6587 ( .A1(n5595), .A2(n5438), .ZN(n5437) );
  NAND2_X1 U6588 ( .A1(n5452), .A2(n5451), .ZN(n7599) );
  NAND2_X1 U6589 ( .A1(n6333), .A2(n5460), .ZN(n5459) );
  NAND2_X1 U6590 ( .A1(n5459), .A2(n5458), .ZN(n9099) );
  OAI211_X2 U6591 ( .C1(n5138), .C2(n5597), .A(n5468), .B(n5467), .ZN(n9409)
         );
  OR2_X1 U6592 ( .A1(n6959), .A2(n6885), .ZN(n5468) );
  NOR2_X1 U6593 ( .A1(n9056), .A2(n5474), .ZN(n5473) );
  NAND2_X1 U6594 ( .A1(n6380), .A2(n5480), .ZN(n5482) );
  OR2_X1 U6595 ( .A1(n5926), .A2(n6486), .ZN(n5911) );
  AND4_X2 U6596 ( .A1(n5887), .A2(n5886), .A3(n5885), .A4(n5884), .ZN(n5897)
         );
  OR2_X1 U6597 ( .A1(n5912), .A2(n6661), .ZN(n5724) );
  INV_X1 U6598 ( .A(n8541), .ZN(n8529) );
  NAND2_X1 U6599 ( .A1(n8659), .A2(n8658), .ZN(n5595) );
  NAND2_X2 U6600 ( .A1(n6459), .A2(n6458), .ZN(n6471) );
  NAND2_X1 U6601 ( .A1(n9101), .A2(n8417), .ZN(n6186) );
  NAND2_X1 U6602 ( .A1(n9115), .A2(n6170), .ZN(n5494) );
  OR2_X1 U6603 ( .A1(n8999), .A2(n5505), .ZN(n5504) );
  OR2_X1 U6604 ( .A1(n8999), .A2(n5150), .ZN(n5508) );
  NAND3_X1 U6605 ( .A1(n5504), .A2(n5503), .A3(n5500), .ZN(n6415) );
  NAND3_X1 U6606 ( .A1(n8999), .A2(n5507), .A3(n5509), .ZN(n5503) );
  NAND2_X1 U6607 ( .A1(n5512), .A2(n5510), .ZN(n6082) );
  NAND2_X1 U6608 ( .A1(n7730), .A2(n5514), .ZN(n5512) );
  OAI21_X1 U6609 ( .B1(n7730), .B2(n5517), .A(n5514), .ZN(n7697) );
  AOI21_X1 U6610 ( .B1(n5518), .B2(n5520), .A(n5519), .ZN(n9024) );
  NAND2_X1 U6611 ( .A1(n5540), .A2(n5541), .ZN(n10179) );
  NAND2_X1 U6612 ( .A1(n5721), .A2(n5160), .ZN(n6532) );
  INV_X1 U6613 ( .A(n6517), .ZN(n6516) );
  NAND3_X1 U6614 ( .A1(n5721), .A2(n5223), .A3(n5160), .ZN(n6517) );
  XNOR2_X2 U6615 ( .A(n5550), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6522) );
  NAND3_X1 U6616 ( .A1(n5555), .A2(n9664), .A3(n5553), .ZN(n5552) );
  NAND4_X1 U6617 ( .A1(n9652), .A2(n9661), .A3(n5556), .A4(n9653), .ZN(n5555)
         );
  NAND3_X1 U6618 ( .A1(n9659), .A2(n9660), .A3(n9658), .ZN(n5556) );
  OR2_X1 U6619 ( .A1(n6222), .A2(n5568), .ZN(n5561) );
  NAND2_X1 U6620 ( .A1(n6222), .A2(n5565), .ZN(n5564) );
  NAND2_X1 U6621 ( .A1(n6012), .A2(n5218), .ZN(n5569) );
  NAND2_X1 U6622 ( .A1(n5569), .A2(n5570), .ZN(n6068) );
  OR2_X1 U6623 ( .A1(n6126), .A2(n6125), .ZN(n5586) );
  NAND2_X1 U6624 ( .A1(n5840), .A2(n5593), .ZN(n5592) );
  INV_X1 U6625 ( .A(n6615), .ZN(n5603) );
  NAND2_X1 U6626 ( .A1(n7071), .A2(n5225), .ZN(n5605) );
  INV_X1 U6627 ( .A(n7221), .ZN(n5608) );
  XNOR2_X1 U6628 ( .A(n8924), .B(n10797), .ZN(n10806) );
  NOR2_X1 U6629 ( .A1(n6809), .A2(n5622), .ZN(n10929) );
  AND2_X1 U6630 ( .A1(n7018), .A2(n7290), .ZN(n5623) );
  NAND2_X1 U6631 ( .A1(n7020), .A2(n5624), .ZN(n7031) );
  NAND3_X1 U6632 ( .A1(n5625), .A2(n6943), .A3(n6953), .ZN(n7012) );
  NAND2_X1 U6633 ( .A1(n6895), .A2(n6894), .ZN(n6943) );
  NAND2_X1 U6634 ( .A1(n9301), .A2(n8354), .ZN(n9375) );
  INV_X1 U6635 ( .A(n8354), .ZN(n5627) );
  NAND2_X1 U6636 ( .A1(n5633), .A2(n5636), .ZN(n7832) );
  NAND2_X1 U6637 ( .A1(n5644), .A2(n9326), .ZN(n8211) );
  NAND2_X1 U6638 ( .A1(n9364), .A2(n9365), .ZN(n8212) );
  NAND3_X1 U6639 ( .A1(n9351), .A2(n5224), .A3(n9352), .ZN(n5645) );
  NAND3_X1 U6640 ( .A1(n9351), .A2(n9352), .A3(n5650), .ZN(n5649) );
  NAND2_X1 U6641 ( .A1(n9351), .A2(n9352), .ZN(n9277) );
  INV_X1 U6642 ( .A(n5649), .ZN(n9278) );
  INV_X1 U6643 ( .A(n9279), .ZN(n5650) );
  OAI21_X1 U6644 ( .B1(n9345), .B2(n5655), .A(n5652), .ZN(n9356) );
  NAND3_X1 U6645 ( .A1(n7320), .A2(n7458), .A3(n7319), .ZN(n7460) );
  NAND2_X1 U6646 ( .A1(n7320), .A2(n7319), .ZN(n5659) );
  XNOR2_X1 U6647 ( .A(n5659), .B(n5240), .ZN(n7335) );
  NAND2_X1 U6648 ( .A1(n5662), .A2(n5660), .ZN(n7945) );
  AND2_X2 U6649 ( .A1(n5666), .A2(n5664), .ZN(n6380) );
  NAND2_X1 U6650 ( .A1(n7573), .A2(n5166), .ZN(n7705) );
  OAI21_X2 U6651 ( .B1(n8716), .B2(n5669), .A(n5667), .ZN(n8722) );
  AOI21_X1 U6652 ( .B1(n8430), .B2(n5680), .A(n5148), .ZN(n8761) );
  OAI21_X1 U6653 ( .B1(n7235), .B2(n5685), .A(n5683), .ZN(n7505) );
  NAND2_X1 U6654 ( .A1(n8106), .A2(n5689), .ZN(n5688) );
  NOR2_X1 U6655 ( .A1(n6348), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n6351) );
  NOR3_X1 U6656 ( .A1(n6348), .A2(P2_IR_REG_27__SCAN_IN), .A3(n5693), .ZN(
        n5867) );
  NAND2_X1 U6657 ( .A1(n5692), .A2(n5165), .ZN(n5758) );
  INV_X1 U6658 ( .A(n6348), .ZN(n5692) );
  AND2_X1 U6661 ( .A1(n11061), .A2(n11085), .ZN(n5696) );
  NAND3_X1 U6662 ( .A1(n5699), .A2(n5701), .A3(n5177), .ZN(n5698) );
  OR2_X1 U6663 ( .A1(n10442), .A2(n10445), .ZN(n5709) );
  NAND2_X1 U6664 ( .A1(n7610), .A2(n5711), .ZN(n5710) );
  NAND2_X1 U6665 ( .A1(n7610), .A2(n5713), .ZN(n5712) );
  NOR2_X1 U6666 ( .A1(n5156), .A2(n5714), .ZN(n5713) );
  NOR2_X2 U6667 ( .A1(n7792), .A2(n5191), .ZN(n7991) );
  INV_X2 U6668 ( .A(n6471), .ZN(n5721) );
  OAI21_X1 U6669 ( .B1(n6173), .B2(n6172), .A(n5835), .ZN(n6188) );
  NAND2_X1 U6670 ( .A1(n6517), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6518) );
  CLKBUF_X1 U6671 ( .A(n6929), .Z(n6934) );
  NAND2_X1 U6672 ( .A1(n9467), .A2(n9643), .ZN(n9506) );
  XNOR2_X1 U6673 ( .A(n6404), .B(n8496), .ZN(n6304) );
  NAND2_X1 U6674 ( .A1(n10407), .A2(n11199), .ZN(n10415) );
  NAND2_X1 U6675 ( .A1(n7013), .A2(n7012), .ZN(n7019) );
  OR2_X1 U6676 ( .A1(n5867), .A2(n9253), .ZN(n5869) );
  NAND2_X1 U6677 ( .A1(n6522), .A2(n6521), .ZN(n6983) );
  INV_X1 U6678 ( .A(n6522), .ZN(n10518) );
  OR2_X1 U6679 ( .A1(n8168), .A2(n6680), .ZN(n6935) );
  OR2_X1 U6680 ( .A1(n6535), .A2(n6534), .ZN(n6536) );
  CLKBUF_X1 U6681 ( .A(n8741), .Z(n8742) );
  OR2_X1 U6682 ( .A1(n5981), .A2(n5888), .ZN(n5895) );
  INV_X1 U6683 ( .A(n8526), .ZN(n6320) );
  NAND2_X1 U6684 ( .A1(n6533), .A2(n6536), .ZN(n10522) );
  AND2_X1 U6685 ( .A1(n9269), .A2(n9270), .ZN(n5723) );
  INV_X1 U6686 ( .A(n9669), .ZN(n10937) );
  NAND2_X1 U6687 ( .A1(n11186), .A2(n9180), .ZN(n9250) );
  INV_X1 U6688 ( .A(n9250), .ZN(n6446) );
  AND2_X1 U6689 ( .A1(n8299), .A2(n8298), .ZN(n5726) );
  OR2_X1 U6690 ( .A1(n8993), .A2(n9250), .ZN(n5727) );
  AND2_X1 U6691 ( .A1(n5813), .A2(n5812), .ZN(n5728) );
  AND2_X1 U6692 ( .A1(n5727), .A2(n6387), .ZN(n5730) );
  INV_X1 U6693 ( .A(n11186), .ZN(n6448) );
  INV_X1 U6694 ( .A(n8607), .ZN(n6330) );
  NAND2_X1 U6695 ( .A1(n5912), .A2(n5134), .ZN(n5909) );
  INV_X1 U6696 ( .A(n6440), .ZN(n8983) );
  INV_X1 U6697 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7912) );
  INV_X1 U6698 ( .A(n9609), .ZN(n9456) );
  INV_X1 U6699 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n5776) );
  INV_X1 U6700 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n5769) );
  NAND2_X1 U6701 ( .A1(n7170), .A2(n10968), .ZN(n10367) );
  INV_X1 U6702 ( .A(n10367), .ZN(n7171) );
  AND2_X1 U6703 ( .A1(n7186), .A2(n11010), .ZN(n5731) );
  NAND2_X2 U6704 ( .A1(n7098), .A2(n6397), .ZN(n9210) );
  INV_X1 U6705 ( .A(n9209), .ZN(n6400) );
  AND2_X1 U6706 ( .A1(n8508), .A2(n6676), .ZN(n5732) );
  INV_X1 U6707 ( .A(n9130), .ZN(n9116) );
  NAND2_X1 U6708 ( .A1(n6303), .A2(n6302), .ZN(n9130) );
  NAND2_X2 U6709 ( .A1(n7128), .A2(n9142), .ZN(n9145) );
  INV_X1 U6710 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n10061) );
  INV_X1 U6711 ( .A(n9561), .ZN(n7542) );
  NOR2_X1 U6712 ( .A1(n7543), .A2(n7542), .ZN(n7544) );
  INV_X1 U6713 ( .A(n6679), .ZN(n6680) );
  INV_X1 U6714 ( .A(n6914), .ZN(n6912) );
  OR2_X1 U6715 ( .A1(n6710), .A2(n7073), .ZN(n6711) );
  OAI21_X1 U6716 ( .B1(n9649), .B2(n10163), .A(n9648), .ZN(n9650) );
  INV_X1 U6717 ( .A(SI_26_), .ZN(n9693) );
  INV_X1 U6718 ( .A(n6251), .ZN(n5745) );
  NAND2_X1 U6719 ( .A1(n8957), .A2(n8956), .ZN(n8958) );
  INV_X1 U6720 ( .A(n6083), .ZN(n5739) );
  INV_X1 U6721 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7802) );
  NAND2_X1 U6722 ( .A1(n7006), .A2(n7005), .ZN(n7007) );
  INV_X1 U6723 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7531) );
  AND2_X1 U6724 ( .A1(n8321), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8336) );
  INV_X1 U6725 ( .A(n6246), .ZN(n5859) );
  INV_X1 U6726 ( .A(SI_19_), .ZN(n9907) );
  OR2_X1 U6727 ( .A1(n7087), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n7088) );
  INV_X1 U6728 ( .A(SI_9_), .ZN(n9928) );
  NAND2_X1 U6729 ( .A1(n5745), .A2(n9759), .ZN(n6253) );
  INV_X1 U6730 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n9979) );
  NAND2_X1 U6731 ( .A1(n5741), .A2(n9767), .ZN(n6164) );
  OR2_X1 U6732 ( .A1(n6061), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6075) );
  INV_X1 U6733 ( .A(n7586), .ZN(n7587) );
  INV_X1 U6734 ( .A(n6433), .ZN(n6434) );
  NOR2_X1 U6735 ( .A1(n7803), .A2(n7802), .ZN(n7994) );
  INV_X1 U6736 ( .A(n6734), .ZN(n8143) );
  AND2_X1 U6737 ( .A1(n9657), .A2(n10158), .ZN(n9658) );
  INV_X1 U6738 ( .A(n6520), .ZN(n6521) );
  INV_X1 U6739 ( .A(n9473), .ZN(n9510) );
  INV_X1 U6740 ( .A(n8218), .ZN(n8238) );
  OR2_X1 U6741 ( .A1(n7412), .A2(n7676), .ZN(n7532) );
  INV_X1 U6742 ( .A(n7322), .ZN(n8214) );
  AND2_X1 U6743 ( .A1(n6280), .A2(n6266), .ZN(n6267) );
  AND2_X1 U6744 ( .A1(n5852), .A2(n5851), .ZN(n6219) );
  INV_X1 U6745 ( .A(SI_15_), .ZN(n5819) );
  NOR2_X1 U6746 ( .A1(n6721), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6832) );
  AND2_X1 U6747 ( .A1(n6377), .A2(n6376), .ZN(n6378) );
  INV_X1 U6748 ( .A(n9054), .ZN(n8709) );
  NAND2_X1 U6749 ( .A1(n5742), .A2(n9752), .ZN(n6191) );
  OR2_X1 U6750 ( .A1(n6213), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6224) );
  NAND2_X2 U6751 ( .A1(n6305), .A2(n6580), .ZN(n5912) );
  INV_X1 U6752 ( .A(n8814), .ZN(n8803) );
  AOI211_X1 U6753 ( .C1(n8687), .C2(n8686), .A(n8685), .B(n8684), .ZN(n8688)
         );
  INV_X1 U6754 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10000) );
  OR2_X1 U6755 ( .A1(n6284), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n8978) );
  INV_X1 U6756 ( .A(n8998), .ZN(n9006) );
  INV_X1 U6757 ( .A(n9041), .ZN(n9048) );
  INV_X1 U6758 ( .A(n9058), .ZN(n9052) );
  OR2_X1 U6759 ( .A1(n6191), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6203) );
  INV_X1 U6760 ( .A(n8559), .ZN(n6323) );
  NAND2_X1 U6761 ( .A1(n6357), .A2(n6499), .ZN(n7095) );
  OR2_X1 U6762 ( .A1(n11186), .A2(n6386), .ZN(n6387) );
  INV_X1 U6763 ( .A(n8835), .ZN(n7892) );
  AND2_X1 U6764 ( .A1(n6371), .A2(n7129), .ZN(n6375) );
  INV_X1 U6765 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n6161) );
  INV_X1 U6766 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n5923) );
  OR2_X1 U6767 ( .A1(n5138), .A2(n10524), .ZN(n8355) );
  AND2_X1 U6768 ( .A1(n9377), .A2(n9374), .ZN(n8354) );
  INV_X1 U6769 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7336) );
  INV_X1 U6770 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7979) );
  INV_X1 U6771 ( .A(n9494), .ZN(n7990) );
  AND4_X1 U6772 ( .A1(n6564), .A2(n6563), .A3(n6562), .A4(n6561), .ZN(n7884)
         );
  AOI21_X1 U6773 ( .B1(n6780), .B2(n10097), .A(n6771), .ZN(n7713) );
  INV_X1 U6774 ( .A(n11195), .ZN(n11147) );
  INV_X1 U6775 ( .A(n7913), .ZN(n6817) );
  AND2_X1 U6776 ( .A1(n6244), .A2(n5856), .ZN(n6232) );
  OR2_X1 U6777 ( .A1(n6832), .A2(n6722), .ZN(n6743) );
  AND2_X1 U6778 ( .A1(n5799), .A2(n5798), .ZN(n5989) );
  AND2_X1 U6779 ( .A1(n5795), .A2(n5794), .ZN(n5973) );
  INV_X1 U6780 ( .A(n5904), .ZN(n5906) );
  NAND2_X1 U6781 ( .A1(n6379), .A2(n6378), .ZN(n6629) );
  AND3_X1 U6782 ( .A1(n6687), .A2(n8692), .A3(n6686), .ZN(n8814) );
  AND2_X1 U6783 ( .A1(n6291), .A2(n6290), .ZN(n8664) );
  AND4_X1 U6784 ( .A1(n6088), .A2(n6087), .A3(n6086), .A4(n6085), .ZN(n8110)
         );
  OR2_X1 U6785 ( .A1(n5891), .A2(n5890), .ZN(n5892) );
  NAND2_X1 U6786 ( .A1(n10752), .A2(n6307), .ZN(n10910) );
  OR3_X1 U6787 ( .A1(n7099), .A2(n7119), .A3(n9173), .ZN(n9142) );
  INV_X1 U6788 ( .A(n8417), .ZN(n9102) );
  AND2_X1 U6789 ( .A1(n8568), .A2(n8561), .ZN(n8480) );
  AND2_X1 U6790 ( .A1(n8547), .A2(n8555), .ZN(n8474) );
  OR2_X1 U6791 ( .A1(n8676), .A2(n6392), .ZN(n7129) );
  NOR2_X1 U6792 ( .A1(n6390), .A2(n6389), .ZN(n7098) );
  NAND2_X1 U6793 ( .A1(n7734), .A2(n7728), .ZN(n9204) );
  INV_X1 U6794 ( .A(P2_IR_REG_29__SCAN_IN), .ZN(n5759) );
  AND2_X1 U6795 ( .A1(n6071), .A2(n6058), .ZN(n10797) );
  AND2_X1 U6796 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n7024) );
  INV_X1 U6797 ( .A(n9397), .ZN(n9381) );
  AND4_X1 U6798 ( .A1(n8386), .A2(n8385), .A3(n8384), .A4(n8383), .ZN(n10401)
         );
  AND4_X1 U6799 ( .A1(n8223), .A2(n8222), .A3(n8221), .A4(n8220), .ZN(n10349)
         );
  AND4_X1 U6800 ( .A1(n7999), .A2(n7998), .A3(n7997), .A4(n7996), .ZN(n8178)
         );
  OR2_X1 U6801 ( .A1(n6968), .A2(n6865), .ZN(n6987) );
  INV_X1 U6802 ( .A(n10949), .ZN(n10744) );
  AND2_X1 U6803 ( .A1(n10184), .A2(n9622), .ZN(n10283) );
  INV_X1 U6804 ( .A(n10373), .ZN(n10370) );
  AND2_X1 U6805 ( .A1(n10367), .A2(n10163), .ZN(n11128) );
  INV_X1 U6806 ( .A(n10233), .ZN(n10335) );
  NOR2_X1 U6807 ( .A1(n10506), .A2(n7711), .ZN(n11123) );
  AND2_X1 U6808 ( .A1(n7714), .A2(n7713), .ZN(n7715) );
  NAND2_X1 U6809 ( .A1(n6814), .A2(n9666), .ZN(n11195) );
  INV_X1 U6810 ( .A(n11199), .ZN(n11176) );
  NAND2_X1 U6811 ( .A1(n10984), .A2(n11091), .ZN(n11199) );
  NOR2_X1 U6812 ( .A1(n10507), .A2(n7712), .ZN(n7721) );
  AND2_X1 U6813 ( .A1(n7141), .A2(n7089), .ZN(n10718) );
  NAND2_X1 U6814 ( .A1(n5904), .A2(n5774), .ZN(n5907) );
  OR2_X1 U6815 ( .A1(n6629), .A2(n6632), .ZN(n6593) );
  INV_X1 U6816 ( .A(n8819), .ZN(n8756) );
  NAND2_X1 U6817 ( .A1(n6639), .A2(n6638), .ZN(n8808) );
  AND2_X1 U6818 ( .A1(n7381), .A2(n7380), .ZN(n8977) );
  INV_X1 U6819 ( .A(n8110), .ZN(n8833) );
  OR2_X1 U6820 ( .A1(n7128), .A2(n9040), .ZN(n9141) );
  INV_X1 U6821 ( .A(n9148), .ZN(n9114) );
  INV_X1 U6822 ( .A(n6442), .ZN(n6443) );
  OR2_X1 U6823 ( .A1(n9210), .A2(n9173), .ZN(n9209) );
  INV_X1 U6824 ( .A(n9210), .ZN(n9206) );
  NOR2_X1 U6825 ( .A1(n8982), .A2(n6439), .ZN(n6449) );
  INV_X1 U6826 ( .A(n8768), .ZN(n9234) );
  AND2_X2 U6827 ( .A1(n6385), .A2(n6495), .ZN(n11186) );
  AND2_X1 U6828 ( .A1(n6477), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6500) );
  INV_X1 U6829 ( .A(n7929), .ZN(n11163) );
  OR2_X1 U6830 ( .A1(n6788), .A2(n6901), .ZN(n9391) );
  AND2_X1 U6831 ( .A1(n6826), .A2(n6825), .ZN(n9397) );
  AND4_X1 U6832 ( .A1(n6842), .A2(n6841), .A3(n6840), .A4(n6839), .ZN(n10408)
         );
  INV_X1 U6833 ( .A(n10297), .ZN(n10445) );
  INV_X1 U6834 ( .A(P1_U3973), .ZN(n9669) );
  INV_X1 U6835 ( .A(n10942), .ZN(n10733) );
  INV_X1 U6836 ( .A(n11129), .ZN(n10391) );
  INV_X1 U6837 ( .A(n11202), .ZN(n11201) );
  INV_X1 U6838 ( .A(n11206), .ZN(n11203) );
  NAND2_X1 U6839 ( .A1(n6575), .A2(n6786), .ZN(n10530) );
  INV_X1 U6840 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n10017) );
  INV_X1 U6841 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n7457) );
  NOR2_X2 U6842 ( .A1(n6593), .A2(P2_U3151), .ZN(P2_U3893) );
  OAI21_X1 U6843 ( .B1(n6402), .B2(n6448), .A(n5730), .ZN(P2_U3455) );
  AND2_X1 U6844 ( .A1(n6476), .A2(n6806), .ZN(P1_U3973) );
  NAND2_X1 U6845 ( .A1(n9959), .A2(n5733), .ZN(n5949) );
  INV_X1 U6846 ( .A(n5949), .ZN(n5734) );
  NAND2_X1 U6847 ( .A1(n5734), .A2(n9975), .ZN(n5965) );
  INV_X1 U6848 ( .A(n5982), .ZN(n5735) );
  NAND2_X1 U6849 ( .A1(n5735), .A2(n9951), .ZN(n6005) );
  OR2_X2 U6850 ( .A1(n6005), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6023) );
  INV_X1 U6851 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5738) );
  OR2_X2 U6852 ( .A1(n6104), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6117) );
  OR2_X2 U6853 ( .A1(n6164), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6179) );
  INV_X1 U6854 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n9759) );
  OR2_X2 U6855 ( .A1(n6253), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n6273) );
  NAND2_X1 U6856 ( .A1(n6253), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U6857 ( .A1(n6273), .A2(n5746), .ZN(n9018) );
  NOR2_X1 U6858 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), .ZN(
        n5752) );
  NOR2_X2 U6859 ( .A1(n5758), .A2(P2_IR_REG_29__SCAN_IN), .ZN(n9252) );
  XNOR2_X2 U6860 ( .A(n5757), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5761) );
  NAND2_X1 U6861 ( .A1(n5758), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5760) );
  NAND2_X1 U6862 ( .A1(n9018), .A2(n5137), .ZN(n5768) );
  INV_X1 U6863 ( .A(P2_REG2_REG_26__SCAN_IN), .ZN(n5765) );
  NAND2_X2 U6864 ( .A1(n8699), .A2(n9260), .ZN(n5981) );
  NAND2_X1 U6865 ( .A1(n7372), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n5764) );
  NAND2_X1 U6866 ( .A1(n5914), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n5763) );
  OAI211_X1 U6867 ( .C1(n5765), .C2(n7377), .A(n5764), .B(n5763), .ZN(n5766)
         );
  INV_X1 U6868 ( .A(n5766), .ZN(n5767) );
  INV_X1 U6869 ( .A(SI_1_), .ZN(n9940) );
  INV_X1 U6870 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n5772) );
  INV_X1 U6871 ( .A(SI_0_), .ZN(n6789) );
  INV_X1 U6872 ( .A(n5905), .ZN(n5774) );
  NAND2_X1 U6873 ( .A1(n5907), .A2(n5775), .ZN(n5928) );
  NAND2_X1 U6874 ( .A1(n6884), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n5777) );
  INV_X1 U6875 ( .A(n5780), .ZN(n5779) );
  INV_X1 U6876 ( .A(SI_3_), .ZN(n9936) );
  NAND2_X1 U6877 ( .A1(n5779), .A2(n9936), .ZN(n5781) );
  NAND2_X1 U6878 ( .A1(n5780), .A2(SI_3_), .ZN(n5782) );
  AND2_X1 U6879 ( .A1(n5781), .A2(n5782), .ZN(n5927) );
  NAND2_X1 U6880 ( .A1(n5928), .A2(n5927), .ZN(n5930) );
  NAND2_X1 U6881 ( .A1(n5930), .A2(n5782), .ZN(n5943) );
  MUX2_X1 U6882 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .S(n6884), .Z(n5783) );
  NAND2_X1 U6883 ( .A1(n5783), .A2(SI_4_), .ZN(n5786) );
  INV_X1 U6884 ( .A(n5783), .ZN(n5784) );
  INV_X1 U6885 ( .A(SI_4_), .ZN(n9941) );
  NAND2_X1 U6886 ( .A1(n5784), .A2(n9941), .ZN(n5785) );
  AND2_X1 U6887 ( .A1(n5786), .A2(n5785), .ZN(n5942) );
  MUX2_X1 U6888 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .S(n6884), .Z(n5787) );
  NAND2_X1 U6889 ( .A1(n5787), .A2(SI_5_), .ZN(n5791) );
  INV_X1 U6890 ( .A(n5787), .ZN(n5789) );
  INV_X1 U6891 ( .A(SI_5_), .ZN(n5788) );
  NAND2_X1 U6892 ( .A1(n5789), .A2(n5788), .ZN(n5790) );
  AND2_X1 U6893 ( .A1(n5791), .A2(n5790), .ZN(n5958) );
  NAND2_X1 U6894 ( .A1(n5792), .A2(SI_6_), .ZN(n5795) );
  INV_X1 U6895 ( .A(n5792), .ZN(n5793) );
  INV_X1 U6896 ( .A(SI_6_), .ZN(n9729) );
  NAND2_X1 U6897 ( .A1(n5793), .A2(n9729), .ZN(n5794) );
  MUX2_X1 U6898 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n6884), .Z(n5796) );
  INV_X1 U6899 ( .A(n5796), .ZN(n5797) );
  INV_X1 U6900 ( .A(SI_7_), .ZN(n9932) );
  NAND2_X1 U6901 ( .A1(n5797), .A2(n9932), .ZN(n5798) );
  MUX2_X1 U6902 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .S(n6884), .Z(n5800) );
  XNOR2_X1 U6903 ( .A(n5800), .B(SI_8_), .ZN(n5997) );
  INV_X1 U6904 ( .A(n5800), .ZN(n5801) );
  INV_X1 U6905 ( .A(SI_8_), .ZN(n9725) );
  NAND2_X1 U6906 ( .A1(n5801), .A2(n9725), .ZN(n5802) );
  NOR2_X1 U6907 ( .A1(n5803), .A2(SI_9_), .ZN(n5804) );
  MUX2_X1 U6908 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .S(n6884), .Z(n5805) );
  NAND2_X1 U6909 ( .A1(n5805), .A2(SI_10_), .ZN(n5808) );
  INV_X1 U6910 ( .A(n5805), .ZN(n5806) );
  NAND2_X1 U6911 ( .A1(n5806), .A2(n9923), .ZN(n5807) );
  NAND2_X1 U6912 ( .A1(n5808), .A2(n5807), .ZN(n6034) );
  MUX2_X1 U6913 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .S(n6884), .Z(n5809) );
  XNOR2_X1 U6914 ( .A(n5809), .B(SI_11_), .ZN(n6051) );
  MUX2_X1 U6915 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n6884), .Z(n5810) );
  NAND2_X1 U6916 ( .A1(n5810), .A2(SI_12_), .ZN(n6089) );
  OAI21_X1 U6917 ( .B1(n5810), .B2(SI_12_), .A(n6089), .ZN(n6067) );
  MUX2_X1 U6918 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n6884), .Z(n6091) );
  NAND2_X1 U6919 ( .A1(n6091), .A2(SI_13_), .ZN(n5811) );
  INV_X1 U6920 ( .A(n6091), .ZN(n5813) );
  INV_X1 U6921 ( .A(SI_13_), .ZN(n5812) );
  MUX2_X1 U6922 ( .A(n6883), .B(n10032), .S(n6884), .Z(n5815) );
  NAND2_X1 U6923 ( .A1(n5815), .A2(n9714), .ZN(n5818) );
  INV_X1 U6924 ( .A(n5815), .ZN(n5816) );
  NAND2_X1 U6925 ( .A1(n5816), .A2(SI_14_), .ZN(n5817) );
  NAND2_X1 U6926 ( .A1(n5818), .A2(n5817), .ZN(n6099) );
  MUX2_X1 U6927 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(P2_DATAO_REG_15__SCAN_IN), 
        .S(n6884), .Z(n5820) );
  XNOR2_X1 U6928 ( .A(n5820), .B(n5819), .ZN(n6111) );
  INV_X1 U6929 ( .A(n6111), .ZN(n5821) );
  MUX2_X1 U6930 ( .A(n7140), .B(n10025), .S(n6884), .Z(n5823) );
  NAND2_X1 U6931 ( .A1(n5823), .A2(n5822), .ZN(n5826) );
  INV_X1 U6932 ( .A(n5823), .ZN(n5824) );
  NAND2_X1 U6933 ( .A1(n5824), .A2(SI_16_), .ZN(n5825) );
  NAND2_X1 U6934 ( .A1(n5826), .A2(n5825), .ZN(n6125) );
  MUX2_X1 U6935 ( .A(n7451), .B(n7457), .S(n6884), .Z(n5827) );
  NAND2_X1 U6936 ( .A1(n5827), .A2(n9913), .ZN(n5830) );
  INV_X1 U6937 ( .A(n5827), .ZN(n5828) );
  NAND2_X1 U6938 ( .A1(n5828), .A2(SI_17_), .ZN(n5829) );
  MUX2_X1 U6939 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n6884), .Z(n5831) );
  XNOR2_X1 U6940 ( .A(n5831), .B(n9912), .ZN(n6155) );
  MUX2_X1 U6941 ( .A(n7655), .B(n7657), .S(n6884), .Z(n5832) );
  NAND2_X1 U6942 ( .A1(n5832), .A2(n9907), .ZN(n5835) );
  INV_X1 U6943 ( .A(n5832), .ZN(n5833) );
  NAND2_X1 U6944 ( .A1(n5833), .A2(SI_19_), .ZN(n5834) );
  NAND2_X1 U6945 ( .A1(n5835), .A2(n5834), .ZN(n6172) );
  MUX2_X1 U6946 ( .A(n7695), .B(n10021), .S(n6884), .Z(n5836) );
  INV_X1 U6947 ( .A(SI_20_), .ZN(n9706) );
  NAND2_X1 U6948 ( .A1(n5836), .A2(n9706), .ZN(n5839) );
  INV_X1 U6949 ( .A(n5836), .ZN(n5837) );
  NAND2_X1 U6950 ( .A1(n5837), .A2(SI_20_), .ZN(n5838) );
  NAND2_X1 U6951 ( .A1(n6188), .A2(n6187), .ZN(n5840) );
  MUX2_X1 U6952 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n6884), .Z(n5843) );
  XNOR2_X1 U6953 ( .A(n5843), .B(n5841), .ZN(n6199) );
  INV_X1 U6954 ( .A(n6199), .ZN(n5842) );
  MUX2_X1 U6955 ( .A(n7859), .B(n9805), .S(n6884), .Z(n5844) );
  INV_X1 U6956 ( .A(SI_22_), .ZN(n9702) );
  NAND2_X1 U6957 ( .A1(n5844), .A2(n9702), .ZN(n5848) );
  INV_X1 U6958 ( .A(n5844), .ZN(n5845) );
  NAND2_X1 U6959 ( .A1(n5845), .A2(SI_22_), .ZN(n5846) );
  NAND2_X1 U6960 ( .A1(n5848), .A2(n5846), .ZN(n6208) );
  INV_X1 U6961 ( .A(n6208), .ZN(n5847) );
  MUX2_X1 U6962 ( .A(n7912), .B(n10017), .S(n6884), .Z(n5849) );
  INV_X1 U6963 ( .A(SI_23_), .ZN(n9701) );
  NAND2_X1 U6964 ( .A1(n5849), .A2(n9701), .ZN(n5852) );
  INV_X1 U6965 ( .A(n5849), .ZN(n5850) );
  NAND2_X1 U6966 ( .A1(n5850), .A2(SI_23_), .ZN(n5851) );
  INV_X1 U6967 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n8082) );
  MUX2_X1 U6968 ( .A(n8082), .B(n9801), .S(n6884), .Z(n5854) );
  INV_X1 U6969 ( .A(SI_24_), .ZN(n5853) );
  NAND2_X1 U6970 ( .A1(n5854), .A2(n5853), .ZN(n6244) );
  INV_X1 U6971 ( .A(n5854), .ZN(n5855) );
  NAND2_X1 U6972 ( .A1(n5855), .A2(SI_24_), .ZN(n5856) );
  INV_X1 U6973 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n8080) );
  MUX2_X1 U6974 ( .A(n8080), .B(n10013), .S(n6884), .Z(n5857) );
  INV_X1 U6975 ( .A(SI_25_), .ZN(n9896) );
  NAND2_X1 U6976 ( .A1(n5857), .A2(n9896), .ZN(n6247) );
  AND2_X1 U6977 ( .A1(n6244), .A2(n6247), .ZN(n5860) );
  INV_X1 U6978 ( .A(n5857), .ZN(n5858) );
  NAND2_X1 U6979 ( .A1(n5858), .A2(SI_25_), .ZN(n6246) );
  INV_X1 U6980 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8157) );
  INV_X1 U6981 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n9797) );
  MUX2_X1 U6982 ( .A(n8157), .B(n9797), .S(n6884), .Z(n5861) );
  NAND2_X1 U6983 ( .A1(n5861), .A2(n9693), .ZN(n6262) );
  INV_X1 U6984 ( .A(n5861), .ZN(n5862) );
  NAND2_X1 U6985 ( .A1(n5862), .A2(SI_26_), .ZN(n5863) );
  OR2_X1 U6986 ( .A1(n5865), .A2(n5864), .ZN(n5866) );
  NAND2_X1 U6987 ( .A1(n6263), .A2(n5866), .ZN(n8332) );
  NAND2_X1 U6988 ( .A1(n8332), .A2(n8468), .ZN(n5874) );
  OR2_X1 U6989 ( .A1(n5926), .A2(n8157), .ZN(n5873) );
  NAND2_X1 U6990 ( .A1(n5876), .A2(n5258), .ZN(n5877) );
  NAND2_X1 U6991 ( .A1(n5878), .A2(n5877), .ZN(n6885) );
  OR2_X1 U6992 ( .A1(n5909), .A2(n6885), .ZN(n5881) );
  INV_X1 U6993 ( .A(n5879), .ZN(n5880) );
  INV_X1 U6994 ( .A(n6682), .ZN(n6932) );
  NAND2_X1 U6995 ( .A1(n5882), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5885) );
  INV_X1 U6996 ( .A(n5981), .ZN(n5883) );
  NAND2_X1 U6997 ( .A1(n5883), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n5886) );
  INV_X1 U6998 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6940) );
  OR2_X1 U6999 ( .A1(n5891), .A2(n6940), .ZN(n5884) );
  NAND2_X1 U7000 ( .A1(n8535), .A2(n8537), .ZN(n6929) );
  INV_X1 U7001 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n5888) );
  NAND2_X1 U7002 ( .A1(n5882), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5893) );
  INV_X1 U7003 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n5890) );
  NAND2_X1 U7004 ( .A1(n5134), .A2(SI_0_), .ZN(n5896) );
  XNOR2_X1 U7005 ( .A(n5896), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9268) );
  MUX2_X1 U7006 ( .A(n10749), .B(n9268), .S(n6479), .Z(n6679) );
  NAND2_X1 U7007 ( .A1(n6929), .A2(n6935), .ZN(n6933) );
  NAND2_X1 U7008 ( .A1(n5897), .A2(n6932), .ZN(n5898) );
  INV_X1 U7009 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n7116) );
  OR2_X1 U7010 ( .A1(n5916), .A2(n7116), .ZN(n5900) );
  INV_X1 U7011 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n7122) );
  OR2_X1 U7012 ( .A1(n5915), .A2(n7122), .ZN(n5899) );
  NAND4_X2 U7013 ( .A1(n5902), .A2(n5901), .A3(n5900), .A4(n5899), .ZN(n8844)
         );
  NOR2_X1 U7014 ( .A1(n5879), .A2(n9253), .ZN(n5903) );
  INV_X1 U7015 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n6486) );
  NAND2_X1 U7016 ( .A1(n5906), .A2(n5905), .ZN(n5908) );
  NAND2_X1 U7017 ( .A1(n5908), .A2(n5907), .ZN(n6944) );
  OR2_X1 U7018 ( .A1(n5909), .A2(n6944), .ZN(n5910) );
  NAND2_X1 U7019 ( .A1(n6923), .A2(n8541), .ZN(n6924) );
  INV_X1 U7020 ( .A(n8844), .ZN(n7046) );
  NAND2_X1 U7021 ( .A1(n7046), .A2(n8539), .ZN(n5913) );
  NAND2_X1 U7022 ( .A1(n6924), .A2(n5913), .ZN(n7044) );
  NAND2_X1 U7023 ( .A1(n6426), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5920) );
  INV_X1 U7024 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n7110) );
  OR2_X1 U7025 ( .A1(n5915), .A2(n7110), .ZN(n5918) );
  OR2_X1 U7026 ( .A1(n5916), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n5917) );
  NOR2_X1 U7027 ( .A1(n5924), .A2(n9253), .ZN(n5921) );
  MUX2_X1 U7028 ( .A(n9253), .B(n5921), .S(P2_IR_REG_3__SCAN_IN), .Z(n5922) );
  INV_X1 U7029 ( .A(n5922), .ZN(n5925) );
  NAND2_X1 U7030 ( .A1(n5924), .A2(n5923), .ZN(n6018) );
  NAND2_X1 U7031 ( .A1(n5925), .A2(n6018), .ZN(n6651) );
  OR2_X1 U7032 ( .A1(n5926), .A2(n5776), .ZN(n5932) );
  OR2_X1 U7033 ( .A1(n5928), .A2(n5927), .ZN(n5929) );
  NAND2_X1 U7034 ( .A1(n5930), .A2(n5929), .ZN(n6960) );
  OR2_X1 U7035 ( .A1(n5909), .A2(n6960), .ZN(n5931) );
  OAI211_X1 U7036 ( .C1(n6479), .C2(n6651), .A(n5932), .B(n5931), .ZN(n7111)
         );
  NAND2_X1 U7037 ( .A1(n8843), .A2(n7111), .ZN(n5933) );
  NAND2_X1 U7038 ( .A1(n7044), .A2(n5933), .ZN(n5935) );
  INV_X1 U7039 ( .A(n7111), .ZN(n7049) );
  NAND2_X1 U7040 ( .A1(n7137), .A2(n7049), .ZN(n5934) );
  NAND2_X1 U7041 ( .A1(n5935), .A2(n5934), .ZN(n7135) );
  NAND2_X1 U7042 ( .A1(n5914), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5941) );
  NAND2_X1 U7043 ( .A1(n6426), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5940) );
  NAND2_X1 U7044 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5936) );
  AND2_X1 U7045 ( .A1(n5949), .A2(n5936), .ZN(n7310) );
  OR2_X1 U7046 ( .A1(n6149), .A2(n7310), .ZN(n5939) );
  INV_X1 U7047 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n5937) );
  OR2_X1 U7048 ( .A1(n7377), .A2(n5937), .ZN(n5938) );
  NAND2_X1 U7049 ( .A1(n6018), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5956) );
  XNOR2_X1 U7050 ( .A(n5956), .B(n6015), .ZN(n6704) );
  INV_X1 U7051 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6488) );
  OR2_X1 U7052 ( .A1(n5926), .A2(n6488), .ZN(n5946) );
  OR2_X1 U7053 ( .A1(n5943), .A2(n5942), .ZN(n5944) );
  OR2_X1 U7054 ( .A1(n5909), .A2(n6999), .ZN(n5945) );
  OAI211_X1 U7055 ( .C1(n6479), .C2(n6704), .A(n5946), .B(n5945), .ZN(n6919)
         );
  NOR2_X1 U7056 ( .A1(n8842), .A2(n6919), .ZN(n5948) );
  NAND2_X1 U7057 ( .A1(n8842), .A2(n6919), .ZN(n5947) );
  NAND2_X1 U7058 ( .A1(n5914), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5955) );
  NAND2_X1 U7059 ( .A1(n5883), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5954) );
  NAND2_X1 U7060 ( .A1(n5949), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5950) );
  AND2_X1 U7061 ( .A1(n5965), .A2(n5950), .ZN(n7492) );
  OR2_X1 U7062 ( .A1(n6149), .A2(n7492), .ZN(n5953) );
  INV_X1 U7063 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n5951) );
  OR2_X1 U7064 ( .A1(n7377), .A2(n5951), .ZN(n5952) );
  NAND4_X1 U7065 ( .A1(n5955), .A2(n5954), .A3(n5953), .A4(n5952), .ZN(n8841)
         );
  NAND2_X1 U7066 ( .A1(n5956), .A2(n6015), .ZN(n5957) );
  NAND2_X1 U7067 ( .A1(n5957), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5971) );
  XNOR2_X1 U7068 ( .A(n5971), .B(n6013), .ZN(n7073) );
  OR2_X1 U7069 ( .A1(n5959), .A2(n5958), .ZN(n5960) );
  NAND2_X1 U7070 ( .A1(n5961), .A2(n5960), .ZN(n7283) );
  OR2_X1 U7071 ( .A1(n6070), .A2(n7283), .ZN(n5963) );
  INV_X1 U7072 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6491) );
  OR2_X1 U7073 ( .A1(n5926), .A2(n6491), .ZN(n5962) );
  OAI211_X1 U7074 ( .C1(n6479), .C2(n7073), .A(n5963), .B(n5962), .ZN(n7041)
         );
  AND2_X1 U7075 ( .A1(n8841), .A2(n7041), .ZN(n5964) );
  OAI22_X1 U7076 ( .A1(n7441), .A2(n5964), .B1(n8841), .B2(n7041), .ZN(n7347)
         );
  NAND2_X1 U7077 ( .A1(n6426), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5970) );
  NAND2_X1 U7078 ( .A1(n5882), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5969) );
  NAND2_X1 U7079 ( .A1(n5965), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n5966) );
  AND2_X1 U7080 ( .A1(n5982), .A2(n5966), .ZN(n7239) );
  OR2_X1 U7081 ( .A1(n6149), .A2(n7239), .ZN(n5968) );
  INV_X1 U7082 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n7078) );
  OR2_X1 U7083 ( .A1(n7374), .A2(n7078), .ZN(n5967) );
  NAND4_X1 U7084 ( .A1(n5970), .A2(n5969), .A3(n5968), .A4(n5967), .ZN(n8840)
         );
  NAND2_X1 U7085 ( .A1(n5971), .A2(n6013), .ZN(n5972) );
  NAND2_X1 U7086 ( .A1(n5972), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5992) );
  XNOR2_X1 U7087 ( .A(n5992), .B(n5991), .ZN(n7077) );
  OR2_X1 U7088 ( .A1(n5974), .A2(n5973), .ZN(n5975) );
  NAND2_X1 U7089 ( .A1(n5976), .A2(n5975), .ZN(n7321) );
  OR2_X1 U7090 ( .A1(n7321), .A2(n6070), .ZN(n5978) );
  OR2_X1 U7091 ( .A1(n5926), .A2(n5322), .ZN(n5977) );
  OAI211_X1 U7092 ( .C1(n6479), .C2(n7077), .A(n5978), .B(n5977), .ZN(n7518)
         );
  NOR2_X1 U7093 ( .A1(n8840), .A2(n7518), .ZN(n5980) );
  NAND2_X1 U7094 ( .A1(n8840), .A2(n7518), .ZN(n5979) );
  NAND2_X1 U7095 ( .A1(n6310), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5988) );
  INV_X2 U7096 ( .A(n5981), .ZN(n6426) );
  NAND2_X1 U7097 ( .A1(n6426), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5987) );
  NAND2_X1 U7098 ( .A1(n5982), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n5983) );
  AND2_X1 U7099 ( .A1(n6005), .A2(n5983), .ZN(n8160) );
  OR2_X1 U7100 ( .A1(n6149), .A2(n8160), .ZN(n5986) );
  INV_X1 U7101 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n5984) );
  OR2_X1 U7102 ( .A1(n7377), .A2(n5984), .ZN(n5985) );
  NAND4_X1 U7103 ( .A1(n5988), .A2(n5987), .A3(n5986), .A4(n5985), .ZN(n8839)
         );
  INV_X1 U7104 ( .A(n8839), .ZN(n7500) );
  OR2_X1 U7105 ( .A1(n7400), .A2(n6070), .ZN(n5995) );
  NAND2_X1 U7106 ( .A1(n5992), .A2(n5991), .ZN(n5993) );
  NAND2_X1 U7107 ( .A1(n5993), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5999) );
  XNOR2_X1 U7108 ( .A(n5999), .B(P2_IR_REG_7__SCAN_IN), .ZN(n7215) );
  AOI22_X1 U7109 ( .A1(n6176), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6175), .B2(
        n7215), .ZN(n5994) );
  NAND2_X1 U7110 ( .A1(n5995), .A2(n5994), .ZN(n8162) );
  NAND2_X1 U7111 ( .A1(n8839), .A2(n8162), .ZN(n5996) );
  NAND2_X1 U7112 ( .A1(n7539), .A2(n8468), .ZN(n6003) );
  INV_X1 U7113 ( .A(P2_IR_REG_7__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7114 ( .A1(n5999), .A2(n5998), .ZN(n6000) );
  NAND2_X1 U7115 ( .A1(n6000), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6001) );
  XNOR2_X1 U7116 ( .A(n6001), .B(P2_IR_REG_8__SCAN_IN), .ZN(n7219) );
  AOI22_X1 U7117 ( .A1(n6176), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6175), .B2(
        n7219), .ZN(n6002) );
  NAND2_X1 U7118 ( .A1(n6426), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n6010) );
  NAND2_X1 U7119 ( .A1(n5882), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n6009) );
  INV_X1 U7120 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n6004) );
  OR2_X1 U7121 ( .A1(n7374), .A2(n6004), .ZN(n6008) );
  NAND2_X1 U7122 ( .A1(n6005), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n6006) );
  AND2_X1 U7123 ( .A1(n6023), .A2(n6006), .ZN(n7508) );
  OR2_X1 U7124 ( .A1(n6149), .A2(n7508), .ZN(n6007) );
  NAND4_X1 U7125 ( .A1(n6016), .A2(n6015), .A3(n6014), .A4(n6013), .ZN(n6017)
         );
  NAND2_X1 U7126 ( .A1(n6038), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6019) );
  XNOR2_X1 U7127 ( .A(n6019), .B(P2_IR_REG_9__SCAN_IN), .ZN(n8920) );
  AOI22_X1 U7128 ( .A1(n6176), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6175), .B2(
        n8920), .ZN(n6020) );
  NAND2_X1 U7129 ( .A1(n6426), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n6028) );
  NAND2_X1 U7130 ( .A1(n5882), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n6027) );
  INV_X1 U7131 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n6022) );
  OR2_X1 U7132 ( .A1(n7374), .A2(n6022), .ZN(n6026) );
  NAND2_X1 U7133 ( .A1(n6023), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n6024) );
  AND2_X1 U7134 ( .A1(n6043), .A2(n6024), .ZN(n7597) );
  OR2_X1 U7135 ( .A1(n6149), .A2(n7597), .ZN(n6025) );
  NAND4_X1 U7136 ( .A1(n6028), .A2(n6027), .A3(n6026), .A4(n6025), .ZN(n8837)
         );
  NAND2_X1 U7137 ( .A1(n7664), .A2(n7510), .ZN(n8522) );
  OR2_X1 U7138 ( .A1(n7589), .A2(n6031), .ZN(n7585) );
  OR2_X1 U7139 ( .A1(n7628), .A2(n8838), .ZN(n7593) );
  INV_X1 U7140 ( .A(n6029), .ZN(n6030) );
  OR2_X1 U7141 ( .A1(n6030), .A2(n7616), .ZN(n7591) );
  NAND2_X1 U7142 ( .A1(n6035), .A2(n6034), .ZN(n6036) );
  NAND2_X1 U7143 ( .A1(n6037), .A2(n6036), .ZN(n7524) );
  OR2_X1 U7144 ( .A1(n7524), .A2(n6070), .ZN(n6041) );
  NOR2_X1 U7145 ( .A1(n6038), .A2(P2_IR_REG_9__SCAN_IN), .ZN(n6054) );
  OR2_X1 U7146 ( .A1(n6054), .A2(n9253), .ZN(n6039) );
  XNOR2_X1 U7147 ( .A(n6039), .B(P2_IR_REG_10__SCAN_IN), .ZN(n10777) );
  AOI22_X1 U7148 ( .A1(n6176), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6175), .B2(
        n10777), .ZN(n6040) );
  NAND2_X1 U7149 ( .A1(n5914), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n6048) );
  INV_X1 U7150 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n6042) );
  OR2_X1 U7151 ( .A1(n5981), .A2(n6042), .ZN(n6047) );
  NAND2_X1 U7152 ( .A1(n6043), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n6044) );
  AND2_X1 U7153 ( .A1(n6061), .A2(n6044), .ZN(n7739) );
  OR2_X1 U7154 ( .A1(n6149), .A2(n7739), .ZN(n6046) );
  INV_X1 U7155 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n8894) );
  OR2_X1 U7156 ( .A1(n7377), .A2(n8894), .ZN(n6045) );
  NAND2_X1 U7157 ( .A1(n7741), .A2(n8836), .ZN(n6049) );
  OR2_X1 U7158 ( .A1(n7741), .A2(n8836), .ZN(n6050) );
  XNOR2_X1 U7159 ( .A(n6052), .B(n6051), .ZN(n7634) );
  NAND2_X1 U7160 ( .A1(n7634), .A2(n8468), .ZN(n6060) );
  NAND2_X1 U7161 ( .A1(n6054), .A2(n6053), .ZN(n6055) );
  NAND2_X1 U7162 ( .A1(n6055), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6057) );
  NAND2_X1 U7163 ( .A1(n6057), .A2(n6056), .ZN(n6071) );
  OR2_X1 U7164 ( .A1(n6057), .A2(n6056), .ZN(n6058) );
  AOI22_X1 U7165 ( .A1(n6176), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6175), .B2(
        n10797), .ZN(n6059) );
  NAND2_X1 U7166 ( .A1(n6060), .A2(n6059), .ZN(n7854) );
  NAND2_X1 U7167 ( .A1(n6426), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n6066) );
  INV_X1 U7168 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n8890) );
  OR2_X1 U7169 ( .A1(n7377), .A2(n8890), .ZN(n6065) );
  NAND2_X1 U7170 ( .A1(n6061), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6062) );
  AND2_X1 U7171 ( .A1(n6075), .A2(n6062), .ZN(n7852) );
  OR2_X1 U7172 ( .A1(n6149), .A2(n7852), .ZN(n6064) );
  INV_X1 U7173 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n8889) );
  OR2_X1 U7174 ( .A1(n7374), .A2(n8889), .ZN(n6063) );
  NAND4_X1 U7175 ( .A1(n6066), .A2(n6065), .A3(n6064), .A4(n6063), .ZN(n8835)
         );
  NAND2_X1 U7176 ( .A1(n6068), .A2(n6067), .ZN(n6069) );
  NAND2_X1 U7177 ( .A1(n6069), .A2(n6090), .ZN(n7754) );
  OR2_X1 U7178 ( .A1(n7754), .A2(n6070), .ZN(n6074) );
  NAND2_X1 U7179 ( .A1(n6071), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6072) );
  XNOR2_X1 U7180 ( .A(n6072), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10812) );
  AOI22_X1 U7181 ( .A1(n6176), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6175), .B2(
        n10812), .ZN(n6073) );
  INV_X1 U7182 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n8886) );
  OR2_X1 U7183 ( .A1(n7374), .A2(n8886), .ZN(n6080) );
  NAND2_X1 U7184 ( .A1(n6426), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U7185 ( .A1(n6075), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n6076) );
  AND2_X1 U7186 ( .A1(n6083), .A2(n6076), .ZN(n7898) );
  OR2_X1 U7187 ( .A1(n6149), .A2(n7898), .ZN(n6078) );
  INV_X1 U7188 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n8887) );
  OR2_X1 U7189 ( .A1(n7377), .A2(n8887), .ZN(n6077) );
  NAND4_X1 U7190 ( .A1(n6080), .A2(n6079), .A3(n6078), .A4(n6077), .ZN(n8834)
         );
  OR2_X1 U7191 ( .A1(n7908), .A2(n7947), .ZN(n8586) );
  NAND2_X1 U7192 ( .A1(n7908), .A2(n7947), .ZN(n8585) );
  NAND2_X1 U7193 ( .A1(n8586), .A2(n8585), .ZN(n7698) );
  NAND2_X1 U7194 ( .A1(n7908), .A2(n8834), .ZN(n6081) );
  NAND2_X1 U7195 ( .A1(n6426), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n6088) );
  INV_X1 U7196 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n8883) );
  OR2_X1 U7197 ( .A1(n7374), .A2(n8883), .ZN(n6087) );
  NAND2_X1 U7198 ( .A1(n6083), .A2(P2_REG3_REG_13__SCAN_IN), .ZN(n6084) );
  AND2_X1 U7199 ( .A1(n6104), .A2(n6084), .ZN(n7950) );
  OR2_X1 U7200 ( .A1(n6149), .A2(n7950), .ZN(n6086) );
  INV_X1 U7201 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n8884) );
  OR2_X1 U7202 ( .A1(n7377), .A2(n8884), .ZN(n6085) );
  NAND2_X1 U7203 ( .A1(n6090), .A2(n6089), .ZN(n6093) );
  XNOR2_X1 U7204 ( .A(n6091), .B(SI_13_), .ZN(n6092) );
  XNOR2_X1 U7205 ( .A(n6093), .B(n6092), .ZN(n7793) );
  NAND2_X1 U7206 ( .A1(n7793), .A2(n8468), .ZN(n6098) );
  NAND2_X1 U7207 ( .A1(n6095), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6096) );
  XNOR2_X1 U7208 ( .A(n6096), .B(P2_IR_REG_13__SCAN_IN), .ZN(n10829) );
  AOI22_X1 U7209 ( .A1(n6176), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6175), .B2(
        n10829), .ZN(n6097) );
  NAND2_X1 U7210 ( .A1(n6098), .A2(n6097), .ZN(n7952) );
  INV_X1 U7211 ( .A(n7952), .ZN(n7860) );
  XNOR2_X1 U7212 ( .A(n6100), .B(n6099), .ZN(n7987) );
  NAND2_X1 U7213 ( .A1(n7987), .A2(n8468), .ZN(n6103) );
  NAND2_X1 U7214 ( .A1(n6101), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6160) );
  XNOR2_X1 U7215 ( .A(n6160), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U7216 ( .A1(n6176), .A2(P1_DATAO_REG_14__SCAN_IN), .B1(n6175), .B2(
        n10845), .ZN(n6102) );
  NAND2_X1 U7217 ( .A1(n6310), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n6109) );
  NAND2_X1 U7218 ( .A1(n6426), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n6108) );
  NAND2_X1 U7219 ( .A1(n6104), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n6105) );
  AND2_X1 U7220 ( .A1(n6117), .A2(n6105), .ZN(n8113) );
  OR2_X1 U7221 ( .A1(n6149), .A2(n8113), .ZN(n6107) );
  INV_X1 U7222 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n8929) );
  OR2_X1 U7223 ( .A1(n7377), .A2(n8929), .ZN(n6106) );
  NAND4_X1 U7224 ( .A1(n6109), .A2(n6108), .A3(n6107), .A4(n6106), .ZN(n8832)
         );
  XNOR2_X1 U7225 ( .A(n8115), .B(n8832), .ZN(n8594) );
  NAND2_X1 U7226 ( .A1(n8115), .A2(n8832), .ZN(n8606) );
  NAND2_X1 U7227 ( .A1(n7917), .A2(n8606), .ZN(n7956) );
  XNOR2_X1 U7228 ( .A(n6112), .B(n6111), .ZN(n8030) );
  NAND2_X1 U7229 ( .A1(n8030), .A2(n8468), .ZN(n6116) );
  INV_X1 U7230 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n6113) );
  NAND2_X1 U7231 ( .A1(n6160), .A2(n6113), .ZN(n6114) );
  NAND2_X1 U7232 ( .A1(n6114), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6128) );
  XNOR2_X1 U7233 ( .A(n6128), .B(P2_IR_REG_15__SCAN_IN), .ZN(n10863) );
  AOI22_X1 U7234 ( .A1(n6176), .A2(P1_DATAO_REG_15__SCAN_IN), .B1(n6175), .B2(
        n10863), .ZN(n6115) );
  INV_X1 U7235 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n8879) );
  OR2_X1 U7236 ( .A1(n7374), .A2(n8879), .ZN(n6122) );
  NAND2_X1 U7237 ( .A1(n6426), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n6121) );
  NAND2_X1 U7238 ( .A1(n6117), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n6118) );
  AND2_X1 U7239 ( .A1(n6132), .A2(n6118), .ZN(n7961) );
  OR2_X1 U7240 ( .A1(n6149), .A2(n7961), .ZN(n6120) );
  INV_X1 U7241 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n8880) );
  OR2_X1 U7242 ( .A1(n7377), .A2(n8880), .ZN(n6119) );
  NAND4_X1 U7243 ( .A1(n6122), .A2(n6121), .A3(n6120), .A4(n6119), .ZN(n8831)
         );
  INV_X1 U7244 ( .A(n8831), .ZN(n6123) );
  OR2_X1 U7245 ( .A1(n8404), .A2(n6123), .ZN(n8598) );
  NAND2_X1 U7246 ( .A1(n8404), .A2(n6123), .ZN(n8599) );
  NAND2_X1 U7247 ( .A1(n8598), .A2(n8599), .ZN(n8607) );
  NAND2_X1 U7248 ( .A1(n7956), .A2(n8607), .ZN(n7955) );
  NAND2_X1 U7249 ( .A1(n8404), .A2(n8831), .ZN(n6124) );
  NAND2_X1 U7250 ( .A1(n7955), .A2(n6124), .ZN(n8013) );
  XNOR2_X1 U7251 ( .A(n6126), .B(n6125), .ZN(n8084) );
  NAND2_X1 U7252 ( .A1(n8084), .A2(n8468), .ZN(n6131) );
  INV_X1 U7253 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n6127) );
  NAND2_X1 U7254 ( .A1(n6128), .A2(n6127), .ZN(n6129) );
  NAND2_X1 U7255 ( .A1(n6129), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6142) );
  XNOR2_X1 U7256 ( .A(n6142), .B(P2_IR_REG_16__SCAN_IN), .ZN(n10879) );
  AOI22_X1 U7257 ( .A1(n6176), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6175), .B2(
        n10879), .ZN(n6130) );
  INV_X1 U7258 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n9207) );
  OR2_X1 U7259 ( .A1(n7374), .A2(n9207), .ZN(n6137) );
  NAND2_X1 U7260 ( .A1(n6426), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n6136) );
  NAND2_X1 U7261 ( .A1(n6132), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n6133) );
  AND2_X1 U7262 ( .A1(n6147), .A2(n6133), .ZN(n8745) );
  OR2_X1 U7263 ( .A1(n6149), .A2(n8745), .ZN(n6135) );
  INV_X1 U7264 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n8936) );
  OR2_X1 U7265 ( .A1(n7377), .A2(n8936), .ZN(n6134) );
  NAND4_X1 U7266 ( .A1(n6137), .A2(n6136), .A3(n6135), .A4(n6134), .ZN(n9135)
         );
  INV_X1 U7267 ( .A(n9135), .ZN(n8408) );
  OR2_X1 U7268 ( .A1(n8739), .A2(n8408), .ZN(n8611) );
  NAND2_X1 U7269 ( .A1(n8739), .A2(n8408), .ZN(n8612) );
  NAND2_X1 U7270 ( .A1(n8611), .A2(n8612), .ZN(n8608) );
  NAND2_X1 U7271 ( .A1(n8013), .A2(n8608), .ZN(n8012) );
  NAND2_X1 U7272 ( .A1(n8739), .A2(n9135), .ZN(n6138) );
  NAND2_X1 U7273 ( .A1(n8012), .A2(n6138), .ZN(n9132) );
  XNOR2_X1 U7274 ( .A(n6140), .B(n6139), .ZN(n8132) );
  NAND2_X1 U7275 ( .A1(n8132), .A2(n8468), .ZN(n6146) );
  INV_X1 U7276 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7277 ( .A1(n6142), .A2(n6141), .ZN(n6143) );
  NAND2_X1 U7278 ( .A1(n6143), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6144) );
  XNOR2_X1 U7279 ( .A(n6144), .B(P2_IR_REG_17__SCAN_IN), .ZN(n10897) );
  AOI22_X1 U7280 ( .A1(n6176), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6175), .B2(
        n10897), .ZN(n6145) );
  INV_X1 U7281 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9200) );
  OR2_X1 U7282 ( .A1(n7374), .A2(n9200), .ZN(n6153) );
  NAND2_X1 U7283 ( .A1(n6426), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n6152) );
  NAND2_X1 U7284 ( .A1(n6147), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n6148) );
  AND2_X1 U7285 ( .A1(n6164), .A2(n6148), .ZN(n9143) );
  OR2_X1 U7286 ( .A1(n6149), .A2(n9143), .ZN(n6151) );
  INV_X1 U7287 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n9144) );
  OR2_X1 U7288 ( .A1(n7377), .A2(n9144), .ZN(n6150) );
  NAND4_X1 U7289 ( .A1(n6153), .A2(n6152), .A3(n6151), .A4(n6150), .ZN(n8830)
         );
  XNOR2_X1 U7290 ( .A(n8758), .B(n9118), .ZN(n9140) );
  NAND2_X1 U7291 ( .A1(n9132), .A2(n9140), .ZN(n9131) );
  NAND2_X1 U7292 ( .A1(n8758), .A2(n8830), .ZN(n6154) );
  XNOR2_X1 U7293 ( .A(n6156), .B(n6155), .ZN(n8203) );
  NAND2_X1 U7294 ( .A1(n8203), .A2(n8468), .ZN(n6163) );
  INV_X1 U7295 ( .A(n6157), .ZN(n6158) );
  NAND2_X1 U7296 ( .A1(n6158), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6159) );
  NAND2_X1 U7297 ( .A1(n6160), .A2(n6159), .ZN(n6174) );
  XNOR2_X1 U7298 ( .A(n6174), .B(n6161), .ZN(n8948) );
  AOI22_X1 U7299 ( .A1(n6176), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6175), .B2(
        n8948), .ZN(n6162) );
  NAND2_X1 U7300 ( .A1(n5914), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n6169) );
  NAND2_X1 U7301 ( .A1(n6164), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n6165) );
  NAND2_X1 U7302 ( .A1(n6179), .A2(n6165), .ZN(n9124) );
  NAND2_X1 U7303 ( .A1(n5137), .A2(n9124), .ZN(n6168) );
  INV_X1 U7304 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n9240) );
  OR2_X1 U7305 ( .A1(n5981), .A2(n9240), .ZN(n6167) );
  INV_X1 U7306 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n8916) );
  OR2_X1 U7307 ( .A1(n7377), .A2(n8916), .ZN(n6166) );
  NAND4_X1 U7308 ( .A1(n6169), .A2(n6168), .A3(n6167), .A4(n6166), .ZN(n9134)
         );
  OR2_X1 U7309 ( .A1(n8786), .A2(n9134), .ZN(n6170) );
  NAND2_X1 U7310 ( .A1(n8786), .A2(n9134), .ZN(n6171) );
  XNOR2_X1 U7311 ( .A(n6173), .B(n6172), .ZN(n8213) );
  NAND2_X1 U7312 ( .A1(n8213), .A2(n8468), .ZN(n6178) );
  XNOR2_X2 U7313 ( .A(n6293), .B(P2_IR_REG_19__SCAN_IN), .ZN(n8962) );
  AOI22_X1 U7314 ( .A1(n6176), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n6175), .B2(
        n8962), .ZN(n6177) );
  NAND2_X1 U7315 ( .A1(n6179), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n6180) );
  NAND2_X1 U7316 ( .A1(n6191), .A2(n6180), .ZN(n9107) );
  NAND2_X1 U7317 ( .A1(n9107), .A2(n5136), .ZN(n6184) );
  NAND2_X1 U7318 ( .A1(n5914), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n6183) );
  NAND2_X1 U7319 ( .A1(n6426), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n6182) );
  INV_X1 U7320 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9109) );
  OR2_X1 U7321 ( .A1(n7377), .A2(n9109), .ZN(n6181) );
  NAND2_X1 U7322 ( .A1(n9237), .A2(n9120), .ZN(n8630) );
  NAND2_X1 U7323 ( .A1(n8631), .A2(n8630), .ZN(n8417) );
  INV_X1 U7324 ( .A(n9120), .ZN(n8829) );
  NAND2_X1 U7325 ( .A1(n9237), .A2(n8829), .ZN(n6185) );
  NAND2_X1 U7326 ( .A1(n6186), .A2(n6185), .ZN(n9089) );
  XNOR2_X1 U7327 ( .A(n6188), .B(n6187), .ZN(n8233) );
  NAND2_X1 U7328 ( .A1(n8233), .A2(n8468), .ZN(n6190) );
  OR2_X1 U7329 ( .A1(n5926), .A2(n7695), .ZN(n6189) );
  INV_X1 U7330 ( .A(P2_REG2_REG_20__SCAN_IN), .ZN(n9095) );
  NAND2_X1 U7331 ( .A1(n6191), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7332 ( .A1(n6203), .A2(n6192), .ZN(n9092) );
  NAND2_X1 U7333 ( .A1(n9092), .A2(n5137), .ZN(n6196) );
  NAND2_X1 U7334 ( .A1(n6310), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n6194) );
  NAND2_X1 U7335 ( .A1(n7372), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n6193) );
  AND2_X1 U7336 ( .A1(n6194), .A2(n6193), .ZN(n6195) );
  OAI211_X1 U7337 ( .C1(n7377), .C2(n9095), .A(n6196), .B(n6195), .ZN(n9104)
         );
  OR2_X1 U7338 ( .A1(n8768), .A2(n9104), .ZN(n6198) );
  NAND2_X1 U7339 ( .A1(n8768), .A2(n9104), .ZN(n6197) );
  NAND2_X1 U7340 ( .A1(n6198), .A2(n6197), .ZN(n9093) );
  XNOR2_X1 U7341 ( .A(n6200), .B(n6199), .ZN(n8250) );
  NAND2_X1 U7342 ( .A1(n8250), .A2(n8468), .ZN(n6202) );
  INV_X1 U7343 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7751) );
  OR2_X1 U7344 ( .A1(n5926), .A2(n7751), .ZN(n6201) );
  INV_X1 U7345 ( .A(P2_REG2_REG_21__SCAN_IN), .ZN(n6207) );
  NAND2_X1 U7346 ( .A1(n6203), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n6204) );
  NAND2_X1 U7347 ( .A1(n6213), .A2(n6204), .ZN(n9084) );
  NAND2_X1 U7348 ( .A1(n9084), .A2(n5136), .ZN(n6206) );
  AOI22_X1 U7349 ( .A1(n7372), .A2(P2_REG0_REG_21__SCAN_IN), .B1(n6310), .B2(
        P2_REG1_REG_21__SCAN_IN), .ZN(n6205) );
  OAI211_X1 U7350 ( .C1(n7377), .C2(n6207), .A(n6206), .B(n6205), .ZN(n9064)
         );
  NAND2_X1 U7351 ( .A1(n9179), .A2(n9064), .ZN(n6336) );
  NAND2_X1 U7352 ( .A1(n5163), .A2(n6208), .ZN(n6209) );
  NAND2_X1 U7353 ( .A1(n6210), .A2(n6209), .ZN(n8272) );
  NAND2_X1 U7354 ( .A1(n8272), .A2(n8468), .ZN(n6212) );
  OR2_X1 U7355 ( .A1(n5926), .A2(n7859), .ZN(n6211) );
  INV_X1 U7356 ( .A(n9175), .ZN(n8785) );
  INV_X1 U7357 ( .A(P2_REG2_REG_22__SCAN_IN), .ZN(n6217) );
  NAND2_X1 U7358 ( .A1(n6213), .A2(P2_REG3_REG_22__SCAN_IN), .ZN(n6214) );
  NAND2_X1 U7359 ( .A1(n6224), .A2(n6214), .ZN(n9069) );
  NAND2_X1 U7360 ( .A1(n9069), .A2(n5137), .ZN(n6216) );
  AOI22_X1 U7361 ( .A1(n7372), .A2(P2_REG0_REG_22__SCAN_IN), .B1(n5914), .B2(
        P2_REG1_REG_22__SCAN_IN), .ZN(n6215) );
  OAI211_X1 U7362 ( .C1(n7377), .C2(n6217), .A(n6216), .B(n6215), .ZN(n9075)
         );
  INV_X1 U7363 ( .A(n9075), .ZN(n8727) );
  NAND2_X1 U7364 ( .A1(n8785), .A2(n8727), .ZN(n6218) );
  OR2_X1 U7365 ( .A1(n6220), .A2(n6219), .ZN(n6221) );
  NAND2_X1 U7366 ( .A1(n6222), .A2(n6221), .ZN(n8292) );
  NOR2_X1 U7367 ( .A1(n5926), .A2(n7912), .ZN(n6223) );
  NAND2_X1 U7368 ( .A1(n6224), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6225) );
  NAND2_X1 U7369 ( .A1(n6236), .A2(n6225), .ZN(n9060) );
  NAND2_X1 U7370 ( .A1(n9060), .A2(n5136), .ZN(n6231) );
  INV_X1 U7371 ( .A(P2_REG2_REG_23__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U7372 ( .A1(n7372), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n6227) );
  NAND2_X1 U7373 ( .A1(n6310), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6226) );
  OAI211_X1 U7374 ( .C1(n6228), .C2(n7377), .A(n6227), .B(n6226), .ZN(n6229)
         );
  INV_X1 U7375 ( .A(n6229), .ZN(n6230) );
  NAND2_X1 U7376 ( .A1(n6231), .A2(n6230), .ZN(n9065) );
  OR2_X1 U7377 ( .A1(n9174), .A2(n9065), .ZN(n8646) );
  NAND2_X1 U7378 ( .A1(n9174), .A2(n9065), .ZN(n8645) );
  INV_X1 U7379 ( .A(n9065), .ZN(n9045) );
  XNOR2_X1 U7380 ( .A(n6233), .B(n6232), .ZN(n8300) );
  NAND2_X1 U7381 ( .A1(n8300), .A2(n8468), .ZN(n6235) );
  OR2_X1 U7382 ( .A1(n5926), .A2(n8082), .ZN(n6234) );
  NAND2_X1 U7383 ( .A1(n6236), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6237) );
  NAND2_X1 U7384 ( .A1(n6251), .A2(n6237), .ZN(n9047) );
  NAND2_X1 U7385 ( .A1(n9047), .A2(n5137), .ZN(n6243) );
  INV_X1 U7386 ( .A(P2_REG2_REG_24__SCAN_IN), .ZN(n6240) );
  NAND2_X1 U7387 ( .A1(n7372), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n6239) );
  NAND2_X1 U7388 ( .A1(n5914), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6238) );
  OAI211_X1 U7389 ( .C1(n6240), .C2(n7377), .A(n6239), .B(n6238), .ZN(n6241)
         );
  INV_X1 U7390 ( .A(n6241), .ZN(n6242) );
  XNOR2_X1 U7391 ( .A(n9039), .B(n8709), .ZN(n9041) );
  AND2_X1 U7392 ( .A1(n6247), .A2(n6246), .ZN(n6248) );
  NAND2_X1 U7393 ( .A1(n8319), .A2(n8468), .ZN(n6250) );
  OR2_X1 U7394 ( .A1(n5926), .A2(n8080), .ZN(n6249) );
  NAND2_X1 U7395 ( .A1(n6251), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n6252) );
  NAND2_X1 U7396 ( .A1(n6253), .A2(n6252), .ZN(n9027) );
  NAND2_X1 U7397 ( .A1(n9027), .A2(n5136), .ZN(n6258) );
  INV_X1 U7398 ( .A(P2_REG2_REG_25__SCAN_IN), .ZN(n9038) );
  NAND2_X1 U7399 ( .A1(n6310), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6255) );
  NAND2_X1 U7400 ( .A1(n7372), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n6254) );
  OAI211_X1 U7401 ( .C1(n9038), .C2(n7377), .A(n6255), .B(n6254), .ZN(n6256)
         );
  INV_X1 U7402 ( .A(n6256), .ZN(n6257) );
  NAND2_X1 U7403 ( .A1(n9162), .A2(n8828), .ZN(n6259) );
  INV_X1 U7404 ( .A(n9162), .ZN(n9029) );
  AOI22_X1 U7405 ( .A1(n9024), .A2(n6259), .B1(n9044), .B2(n9029), .ZN(n9013)
         );
  NAND2_X1 U7406 ( .A1(n9013), .A2(n6260), .ZN(n6261) );
  OAI21_X1 U7407 ( .B1(n8735), .B2(n9222), .A(n6261), .ZN(n8999) );
  NAND2_X1 U7408 ( .A1(n6263), .A2(n6262), .ZN(n6268) );
  INV_X1 U7409 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8449) );
  INV_X1 U7410 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n10524) );
  MUX2_X1 U7411 ( .A(n8449), .B(n10524), .S(n6884), .Z(n6264) );
  INV_X1 U7412 ( .A(SI_27_), .ZN(n9893) );
  NAND2_X1 U7413 ( .A1(n6264), .A2(n9893), .ZN(n6280) );
  INV_X1 U7414 ( .A(n6264), .ZN(n6265) );
  NAND2_X1 U7415 ( .A1(n6265), .A2(SI_27_), .ZN(n6266) );
  NAND2_X1 U7416 ( .A1(n6268), .A2(n6267), .ZN(n6281) );
  OR2_X1 U7417 ( .A1(n6268), .A2(n6267), .ZN(n6269) );
  NAND2_X1 U7418 ( .A1(n6281), .A2(n6269), .ZN(n8448) );
  OR2_X1 U7419 ( .A1(n5926), .A2(n8449), .ZN(n6270) );
  INV_X1 U7420 ( .A(n6273), .ZN(n6272) );
  INV_X1 U7421 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n6271) );
  NAND2_X1 U7422 ( .A1(n6272), .A2(n6271), .ZN(n6284) );
  NAND2_X1 U7423 ( .A1(n6273), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n6274) );
  NAND2_X1 U7424 ( .A1(n6284), .A2(n6274), .ZN(n9003) );
  NAND2_X1 U7425 ( .A1(n9003), .A2(n5136), .ZN(n6279) );
  INV_X1 U7426 ( .A(P2_REG2_REG_27__SCAN_IN), .ZN(n9008) );
  NAND2_X1 U7427 ( .A1(n7372), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n6276) );
  NAND2_X1 U7428 ( .A1(n6310), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6275) );
  OAI211_X1 U7429 ( .C1(n9008), .C2(n7377), .A(n6276), .B(n6275), .ZN(n6277)
         );
  INV_X1 U7430 ( .A(n6277), .ZN(n6278) );
  INV_X1 U7431 ( .A(n9015), .ZN(n8827) );
  INV_X1 U7432 ( .A(n9155), .ZN(n9009) );
  MUX2_X1 U7433 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n6884), .Z(n6407) );
  INV_X1 U7434 ( .A(SI_28_), .ZN(n6408) );
  XNOR2_X1 U7435 ( .A(n6407), .B(n6408), .ZN(n6405) );
  NAND2_X1 U7436 ( .A1(n10519), .A2(n8468), .ZN(n6283) );
  INV_X1 U7437 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n9266) );
  OR2_X1 U7438 ( .A1(n5926), .A2(n9266), .ZN(n6282) );
  NAND2_X1 U7439 ( .A1(n6284), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n6285) );
  NAND2_X1 U7440 ( .A1(n8978), .A2(n6285), .ZN(n8991) );
  NAND2_X1 U7441 ( .A1(n8991), .A2(n5137), .ZN(n6291) );
  INV_X1 U7442 ( .A(P2_REG2_REG_28__SCAN_IN), .ZN(n6288) );
  NAND2_X1 U7443 ( .A1(n7372), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n6287) );
  NAND2_X1 U7444 ( .A1(n6310), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6286) );
  OAI211_X1 U7445 ( .C1(n6288), .C2(n7377), .A(n6287), .B(n6286), .ZN(n6289)
         );
  INV_X1 U7446 ( .A(n6289), .ZN(n6290) );
  NAND2_X1 U7447 ( .A1(n8665), .A2(n8664), .ZN(n8499) );
  NAND2_X1 U7448 ( .A1(n6417), .A2(n8499), .ZN(n8439) );
  NAND2_X1 U7449 ( .A1(n6293), .A2(n6292), .ZN(n6294) );
  NAND2_X2 U7450 ( .A1(n6300), .A2(n6299), .ZN(n8673) );
  OR2_X1 U7451 ( .A1(n5140), .A2(n8673), .ZN(n6303) );
  NAND2_X1 U7452 ( .A1(n5205), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6301) );
  NAND2_X1 U7453 ( .A1(n8962), .A2(n8694), .ZN(n6302) );
  INV_X1 U7454 ( .A(n6306), .ZN(n8691) );
  INV_X1 U7455 ( .A(n6580), .ZN(n6307) );
  INV_X2 U7456 ( .A(n6307), .ZN(n6588) );
  NAND2_X1 U7457 ( .A1(n8691), .A2(n6307), .ZN(n6308) );
  NAND2_X1 U7458 ( .A1(n6479), .A2(n6308), .ZN(n6686) );
  NOR2_X1 U7459 ( .A1(n9015), .A2(n9119), .ZN(n6317) );
  INV_X1 U7460 ( .A(n8978), .ZN(n6309) );
  NAND2_X1 U7461 ( .A1(n6309), .A2(n5136), .ZN(n7381) );
  INV_X1 U7462 ( .A(P2_REG2_REG_29__SCAN_IN), .ZN(n6313) );
  NAND2_X1 U7463 ( .A1(n7372), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n6312) );
  NAND2_X1 U7464 ( .A1(n6310), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6311) );
  OAI211_X1 U7465 ( .C1(n7377), .C2(n6313), .A(n6312), .B(n6311), .ZN(n6314)
         );
  INV_X1 U7466 ( .A(n6314), .ZN(n6315) );
  NAND2_X1 U7467 ( .A1(n7381), .A2(n6315), .ZN(n8826) );
  INV_X1 U7468 ( .A(n8826), .ZN(n6414) );
  NOR2_X1 U7469 ( .A1(n6414), .A2(n9121), .ZN(n6316) );
  INV_X1 U7470 ( .A(n6929), .ZN(n8477) );
  NAND2_X1 U7471 ( .A1(n8477), .A2(n6320), .ZN(n6931) );
  NAND2_X1 U7472 ( .A1(n6931), .A2(n8537), .ZN(n6922) );
  NAND2_X1 U7473 ( .A1(n6922), .A2(n8529), .ZN(n6321) );
  NAND2_X1 U7474 ( .A1(n7046), .A2(n6730), .ZN(n8531) );
  NAND2_X1 U7475 ( .A1(n6321), .A2(n8531), .ZN(n7048) );
  NAND2_X1 U7476 ( .A1(n7137), .A2(n7111), .ZN(n8547) );
  NAND2_X1 U7477 ( .A1(n8843), .A2(n7049), .ZN(n8555) );
  NAND2_X1 U7478 ( .A1(n7048), .A2(n8474), .ZN(n6322) );
  NAND2_X1 U7479 ( .A1(n6322), .A2(n8547), .ZN(n7134) );
  NAND2_X1 U7480 ( .A1(n7047), .A2(n6919), .ZN(n8552) );
  INV_X1 U7481 ( .A(n6919), .ZN(n7311) );
  NAND2_X1 U7482 ( .A1(n8842), .A2(n7311), .ZN(n8548) );
  NAND2_X1 U7483 ( .A1(n7349), .A2(n7041), .ZN(n8553) );
  AND2_X1 U7484 ( .A1(n8552), .A2(n8553), .ZN(n6324) );
  INV_X1 U7485 ( .A(n7041), .ZN(n7493) );
  NAND2_X1 U7486 ( .A1(n8841), .A2(n7493), .ZN(n8559) );
  INV_X1 U7487 ( .A(n8840), .ZN(n6325) );
  NAND2_X1 U7488 ( .A1(n6325), .A2(n7518), .ZN(n8568) );
  INV_X1 U7489 ( .A(n7518), .ZN(n7351) );
  NAND2_X1 U7490 ( .A1(n8840), .A2(n7351), .ZN(n8561) );
  NAND2_X1 U7491 ( .A1(n7350), .A2(n8480), .ZN(n6326) );
  NAND2_X1 U7492 ( .A1(n6326), .A2(n8568), .ZN(n7478) );
  INV_X1 U7493 ( .A(n7478), .ZN(n6327) );
  NAND2_X1 U7494 ( .A1(n6327), .A2(n8560), .ZN(n7477) );
  NAND2_X1 U7495 ( .A1(n8519), .A2(n8839), .ZN(n7614) );
  AND2_X1 U7496 ( .A1(n8515), .A2(n7614), .ZN(n8573) );
  OR2_X1 U7497 ( .A1(n7741), .A2(n7849), .ZN(n8578) );
  AND2_X1 U7498 ( .A1(n8578), .A2(n8516), .ZN(n8571) );
  NAND2_X1 U7499 ( .A1(n7599), .A2(n8571), .ZN(n6328) );
  NAND2_X1 U7500 ( .A1(n7741), .A2(n7849), .ZN(n8574) );
  NAND2_X1 U7501 ( .A1(n6328), .A2(n8574), .ZN(n7670) );
  OR2_X1 U7502 ( .A1(n7854), .A2(n7892), .ZN(n8579) );
  NAND2_X1 U7503 ( .A1(n7854), .A2(n7892), .ZN(n8580) );
  NAND2_X1 U7504 ( .A1(n7670), .A2(n8486), .ZN(n7669) );
  NAND2_X1 U7505 ( .A1(n7669), .A2(n8580), .ZN(n7696) );
  NAND2_X1 U7506 ( .A1(n7696), .A2(n5511), .ZN(n6329) );
  AND2_X1 U7507 ( .A1(n7952), .A2(n8110), .ZN(n8591) );
  OR2_X1 U7508 ( .A1(n7952), .A2(n8110), .ZN(n7816) );
  INV_X1 U7509 ( .A(n8832), .ZN(n8817) );
  INV_X1 U7510 ( .A(n8608), .ZN(n8489) );
  INV_X1 U7511 ( .A(n9140), .ZN(n6331) );
  NAND2_X1 U7512 ( .A1(n9139), .A2(n6331), .ZN(n6333) );
  OR2_X1 U7513 ( .A1(n8758), .A2(n9118), .ZN(n6332) );
  INV_X1 U7514 ( .A(n9134), .ZN(n8753) );
  OR2_X1 U7515 ( .A1(n8786), .A2(n8753), .ZN(n8620) );
  NAND2_X1 U7516 ( .A1(n8786), .A2(n8753), .ZN(n8618) );
  NAND2_X1 U7517 ( .A1(n8620), .A2(n8618), .ZN(n9123) );
  INV_X1 U7518 ( .A(n8618), .ZN(n6334) );
  INV_X1 U7519 ( .A(n9104), .ZN(n9077) );
  OR2_X1 U7520 ( .A1(n8768), .A2(n9077), .ZN(n6335) );
  INV_X1 U7521 ( .A(n9064), .ZN(n9091) );
  AND2_X1 U7522 ( .A1(n9175), .A2(n8727), .ZN(n8472) );
  INV_X1 U7523 ( .A(n8651), .ZN(n6338) );
  NAND2_X1 U7524 ( .A1(n9039), .A2(n8709), .ZN(n9032) );
  NAND2_X1 U7525 ( .A1(n9162), .A2(n9044), .ZN(n8652) );
  AND2_X1 U7526 ( .A1(n9032), .A2(n8652), .ZN(n6337) );
  NOR2_X1 U7527 ( .A1(n8806), .A2(n8735), .ZN(n8656) );
  NAND2_X1 U7528 ( .A1(n9155), .A2(n9015), .ZN(n8661) );
  NAND2_X1 U7529 ( .A1(n8806), .A2(n8735), .ZN(n8471) );
  NAND2_X1 U7530 ( .A1(n8661), .A2(n8471), .ZN(n6416) );
  NOR2_X1 U7531 ( .A1(n9005), .A2(n6416), .ZN(n6340) );
  INV_X1 U7532 ( .A(n8660), .ZN(n6339) );
  NOR2_X1 U7533 ( .A1(n6340), .A2(n6339), .ZN(n6341) );
  INV_X1 U7534 ( .A(n8439), .ZN(n8496) );
  XNOR2_X1 U7535 ( .A(n6341), .B(n8496), .ZN(n8995) );
  INV_X1 U7536 ( .A(n8962), .ZN(n7654) );
  NAND2_X1 U7537 ( .A1(n8673), .A2(n7654), .ZN(n6392) );
  OR2_X1 U7538 ( .A1(n8962), .A2(n7857), .ZN(n6394) );
  NAND2_X1 U7539 ( .A1(n6392), .A2(n6394), .ZN(n6342) );
  AND2_X1 U7540 ( .A1(n9173), .A2(n6342), .ZN(n6343) );
  NAND2_X1 U7541 ( .A1(n6343), .A2(n7129), .ZN(n7734) );
  NOR2_X1 U7542 ( .A1(n7119), .A2(n8694), .ZN(n7448) );
  INV_X1 U7543 ( .A(n7448), .ZN(n7728) );
  NOR2_X1 U7544 ( .A1(n8990), .A2(n6344), .ZN(n6402) );
  XNOR2_X1 U7545 ( .A(n6354), .B(P2_B_REG_SCAN_IN), .ZN(n6350) );
  NAND2_X1 U7546 ( .A1(n6348), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6349) );
  NAND2_X1 U7547 ( .A1(n6350), .A2(n8079), .ZN(n6353) );
  INV_X1 U7548 ( .A(n6379), .ZN(n6356) );
  NAND2_X1 U7549 ( .A1(n6356), .A2(n6354), .ZN(n6496) );
  OAI21_X1 U7550 ( .B1(n6494), .B2(P2_D_REG_0__SCAN_IN), .A(n6496), .ZN(n6355)
         );
  INV_X1 U7551 ( .A(n6355), .ZN(n6675) );
  NAND2_X1 U7552 ( .A1(n6356), .A2(n8079), .ZN(n6499) );
  INV_X1 U7553 ( .A(n7095), .ZN(n6358) );
  AND2_X1 U7554 ( .A1(n6675), .A2(n6358), .ZN(n6390) );
  NOR2_X1 U7555 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .ZN(
        n6362) );
  NOR4_X1 U7556 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6361) );
  NOR4_X1 U7557 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6360) );
  NOR4_X1 U7558 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6359) );
  NAND4_X1 U7559 ( .A1(n6362), .A2(n6361), .A3(n6360), .A4(n6359), .ZN(n6368)
         );
  NOR4_X1 U7560 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6366) );
  NOR4_X1 U7561 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6365) );
  NOR4_X1 U7562 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6364) );
  NOR4_X1 U7563 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6363) );
  NAND4_X1 U7564 ( .A1(n6366), .A2(n6365), .A3(n6364), .A4(n6363), .ZN(n6367)
         );
  NOR2_X1 U7565 ( .A1(n6368), .A2(n6367), .ZN(n6369) );
  NAND2_X1 U7566 ( .A1(n6390), .A2(n6388), .ZN(n6640) );
  NOR3_X1 U7567 ( .A1(n8673), .A2(n7654), .A3(n7857), .ZN(n6370) );
  AND2_X1 U7568 ( .A1(n5140), .A2(n6370), .ZN(n6626) );
  INV_X1 U7569 ( .A(n6626), .ZN(n6371) );
  NAND2_X1 U7570 ( .A1(n8676), .A2(n9173), .ZN(n6637) );
  OR2_X1 U7571 ( .A1(n6637), .A2(n6626), .ZN(n6373) );
  INV_X1 U7572 ( .A(n7119), .ZN(n6372) );
  NAND2_X1 U7573 ( .A1(n6373), .A2(n9040), .ZN(n6625) );
  NAND2_X1 U7574 ( .A1(n6687), .A2(n6625), .ZN(n6374) );
  OAI21_X1 U7575 ( .B1(n6640), .B2(n6375), .A(n6374), .ZN(n6385) );
  INV_X1 U7576 ( .A(n8079), .ZN(n6377) );
  INV_X1 U7577 ( .A(n6354), .ZN(n6376) );
  INV_X1 U7578 ( .A(n6380), .ZN(n6381) );
  NAND2_X1 U7579 ( .A1(n6381), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6382) );
  MUX2_X1 U7580 ( .A(P2_IR_REG_31__SCAN_IN), .B(n6382), .S(
        P2_IR_REG_23__SCAN_IN), .Z(n6384) );
  INV_X1 U7581 ( .A(n6345), .ZN(n6383) );
  NAND2_X1 U7582 ( .A1(n6384), .A2(n6383), .ZN(n6477) );
  INV_X1 U7583 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6386) );
  NAND2_X1 U7584 ( .A1(n6495), .A2(n6388), .ZN(n6389) );
  NAND2_X1 U7585 ( .A1(n7448), .A2(n5140), .ZN(n6391) );
  NAND2_X1 U7586 ( .A1(n6675), .A2(n6391), .ZN(n6396) );
  INV_X1 U7587 ( .A(n6392), .ZN(n6393) );
  OR2_X1 U7588 ( .A1(n8676), .A2(n6393), .ZN(n6630) );
  OR2_X1 U7589 ( .A1(n6394), .A2(n8673), .ZN(n6395) );
  NAND2_X1 U7590 ( .A1(n8676), .A2(n6395), .ZN(n7096) );
  NAND2_X1 U7591 ( .A1(n6630), .A2(n7096), .ZN(n7092) );
  AOI22_X1 U7592 ( .A1(n6396), .A2(n7092), .B1(n7095), .B2(n7096), .ZN(n6397)
         );
  INV_X1 U7593 ( .A(P2_REG1_REG_28__SCAN_IN), .ZN(n6398) );
  NOR2_X1 U7594 ( .A1(n9206), .A2(n6398), .ZN(n6399) );
  OAI21_X1 U7595 ( .B1(n6402), .B2(n9210), .A(n6401), .ZN(P2_U3487) );
  NAND2_X1 U7596 ( .A1(n8993), .A2(n8664), .ZN(n6403) );
  NAND2_X1 U7597 ( .A1(n6406), .A2(n6405), .ZN(n6411) );
  INV_X1 U7598 ( .A(n6407), .ZN(n6409) );
  NAND2_X1 U7599 ( .A1(n6409), .A2(n6408), .ZN(n6410) );
  INV_X1 U7600 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n9406) );
  INV_X1 U7601 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9259) );
  MUX2_X1 U7602 ( .A(n9406), .B(n9259), .S(n5134), .Z(n8450) );
  NAND2_X1 U7603 ( .A1(n9405), .A2(n8468), .ZN(n6413) );
  OR2_X1 U7604 ( .A1(n5926), .A2(n9259), .ZN(n6412) );
  NAND2_X1 U7605 ( .A1(n6413), .A2(n6412), .ZN(n6440) );
  OR2_X1 U7606 ( .A1(n6440), .A2(n6414), .ZN(n8679) );
  NAND2_X1 U7607 ( .A1(n6440), .A2(n6414), .ZN(n8671) );
  NAND2_X1 U7608 ( .A1(n8679), .A2(n8671), .ZN(n8669) );
  NAND2_X1 U7609 ( .A1(n6415), .A2(n9130), .ZN(n6437) );
  INV_X1 U7610 ( .A(n9017), .ZN(n6422) );
  INV_X1 U7611 ( .A(n6416), .ZN(n8500) );
  NAND2_X1 U7612 ( .A1(n8496), .A2(n8500), .ZN(n6421) );
  NAND2_X1 U7613 ( .A1(n6417), .A2(n8660), .ZN(n6419) );
  AND2_X1 U7614 ( .A1(n8661), .A2(n8656), .ZN(n6418) );
  OR2_X1 U7615 ( .A1(n6419), .A2(n6418), .ZN(n6420) );
  NAND2_X1 U7616 ( .A1(n6420), .A2(n8499), .ZN(n8501) );
  OAI21_X1 U7617 ( .B1(n6422), .B2(n6421), .A(n8501), .ZN(n6424) );
  INV_X1 U7618 ( .A(n6424), .ZN(n6423) );
  NOR2_X1 U7619 ( .A1(n8989), .A2(n7734), .ZN(n6435) );
  AND2_X1 U7620 ( .A1(n6479), .A2(P2_B_REG_SCAN_IN), .ZN(n6425) );
  NOR2_X1 U7621 ( .A1(n9121), .A2(n6425), .ZN(n8975) );
  INV_X1 U7622 ( .A(P2_REG2_REG_30__SCAN_IN), .ZN(n6430) );
  NAND2_X1 U7623 ( .A1(n6426), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n6429) );
  INV_X1 U7624 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n6427) );
  OR2_X1 U7625 ( .A1(n7374), .A2(n6427), .ZN(n6428) );
  OAI211_X1 U7626 ( .C1(n6430), .C2(n7377), .A(n6429), .B(n6428), .ZN(n6431)
         );
  INV_X1 U7627 ( .A(n6431), .ZN(n6432) );
  NAND2_X1 U7628 ( .A1(n7381), .A2(n6432), .ZN(n8825) );
  AOI22_X1 U7629 ( .A1(n9000), .A2(n9136), .B1(n8975), .B2(n8825), .ZN(n6433)
         );
  NOR2_X1 U7630 ( .A1(n6435), .A2(n6434), .ZN(n6436) );
  NAND2_X1 U7631 ( .A1(n6437), .A2(n6436), .ZN(n8982) );
  INV_X1 U7632 ( .A(n8989), .ZN(n6438) );
  NAND2_X1 U7633 ( .A1(n9210), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6441) );
  OAI21_X1 U7634 ( .B1(n8983), .B2(n9209), .A(n6441), .ZN(n6442) );
  OAI21_X1 U7635 ( .B1(n6449), .B2(n9210), .A(n6443), .ZN(P2_U3488) );
  INV_X1 U7636 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6444) );
  OAI21_X1 U7637 ( .B1(n6449), .B2(n6448), .A(n6447), .ZN(P2_U3456) );
  NAND4_X1 U7638 ( .A1(n6544), .A2(n10062), .A3(n10061), .A4(n9846), .ZN(n6456) );
  NOR2_X1 U7639 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6454) );
  NAND4_X1 U7640 ( .A1(n6454), .A2(n6453), .A3(n6452), .A4(n6451), .ZN(n6455)
         );
  NOR2_X1 U7641 ( .A1(n6456), .A2(n6455), .ZN(n6457) );
  NAND2_X1 U7642 ( .A1(n6492), .A2(n6457), .ZN(n7487) );
  INV_X1 U7643 ( .A(n7487), .ZN(n6459) );
  NAND2_X1 U7644 ( .A1(n6537), .A2(n10069), .ZN(n6463) );
  NAND2_X1 U7645 ( .A1(n6463), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6464) );
  NAND2_X1 U7646 ( .A1(n6817), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6574) );
  INV_X1 U7647 ( .A(n6574), .ZN(n6476) );
  OAI21_X1 U7648 ( .B1(P1_IR_REG_22__SCAN_IN), .B2(P1_IR_REG_23__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6465) );
  XNOR2_X2 U7649 ( .A(n6466), .B(n10082), .ZN(n6571) );
  NOR2_X1 U7650 ( .A1(P1_IR_REG_24__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n6469) );
  NOR2_X1 U7651 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_20__SCAN_IN), .ZN(
        n6468) );
  NAND4_X1 U7652 ( .A1(n6469), .A2(n6468), .A3(n10069), .A4(n6467), .ZN(n6470)
         );
  NAND2_X1 U7653 ( .A1(n6515), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6472) );
  NAND2_X1 U7654 ( .A1(n5204), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6473) );
  MUX2_X1 U7655 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6473), .S(
        P1_IR_REG_25__SCAN_IN), .Z(n6474) );
  NAND2_X1 U7656 ( .A1(n6474), .A2(n6515), .ZN(n8071) );
  NOR2_X1 U7657 ( .A1(n8155), .A2(n8071), .ZN(n6475) );
  INV_X1 U7658 ( .A(n6477), .ZN(n6632) );
  OR2_X1 U7659 ( .A1(n8676), .A2(n6632), .ZN(n6478) );
  NAND2_X1 U7660 ( .A1(n6594), .A2(n6479), .ZN(n6480) );
  NAND2_X1 U7661 ( .A1(n6480), .A2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3150) );
  NOR2_X1 U7662 ( .A1(n5134), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10513) );
  INV_X2 U7663 ( .A(n10513), .ZN(n10517) );
  OAI222_X1 U7664 ( .A1(P1_U3086), .A2(n10600), .B1(n10517), .B2(n6885), .C1(
        n5597), .C2(n5141), .ZN(P1_U3354) );
  NOR2_X1 U7665 ( .A1(n6481), .A2(n6722), .ZN(n6483) );
  INV_X1 U7666 ( .A(n6484), .ZN(n6485) );
  INV_X1 U7667 ( .A(n6863), .ZN(n10920) );
  OAI222_X1 U7668 ( .A1(P1_U3086), .A2(n10920), .B1(n10517), .B2(n6944), .C1(
        n5399), .C2(n5141), .ZN(P1_U3353) );
  AND2_X1 U7669 ( .A1(n5134), .A2(P2_U3151), .ZN(n9263) );
  INV_X2 U7670 ( .A(n9263), .ZN(n9262) );
  NOR2_X1 U7671 ( .A1(n5134), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9256) );
  INV_X2 U7672 ( .A(n9256), .ZN(n9267) );
  OAI222_X1 U7673 ( .A1(n9262), .A2(n6944), .B1(n9267), .B2(n6486), .C1(
        P2_U3151), .C2(n6613), .ZN(P2_U3293) );
  OAI222_X1 U7674 ( .A1(n9262), .A2(n6885), .B1(n9267), .B2(n5769), .C1(
        P2_U3151), .C2(n6661), .ZN(P2_U3294) );
  OAI222_X1 U7675 ( .A1(n9262), .A2(n6960), .B1(n9267), .B2(n5776), .C1(
        P2_U3151), .C2(n6651), .ZN(P2_U3292) );
  NAND2_X1 U7676 ( .A1(n6482), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6487) );
  XNOR2_X1 U7677 ( .A(n6487), .B(P1_IR_REG_3__SCAN_IN), .ZN(n10620) );
  INV_X1 U7678 ( .A(n10620), .ZN(n6961) );
  INV_X1 U7679 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n6958) );
  OAI222_X1 U7680 ( .A1(P1_U3086), .A2(n6961), .B1(n10517), .B2(n6960), .C1(
        n6958), .C2(n5141), .ZN(P1_U3352) );
  OAI222_X1 U7681 ( .A1(n9262), .A2(n6999), .B1(n9267), .B2(n6488), .C1(
        P2_U3151), .C2(n6704), .ZN(P2_U3291) );
  INV_X1 U7682 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n7000) );
  NAND2_X1 U7683 ( .A1(n6489), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6490) );
  XNOR2_X1 U7684 ( .A(n6490), .B(P1_IR_REG_4__SCAN_IN), .ZN(n6866) );
  INV_X1 U7685 ( .A(n6866), .ZN(n10948) );
  OAI222_X1 U7686 ( .A1(n5141), .A2(n7000), .B1(n10517), .B2(n6999), .C1(
        n10948), .C2(P1_U3086), .ZN(P1_U3351) );
  OAI222_X1 U7687 ( .A1(n9267), .A2(n6491), .B1(n9262), .B2(n7283), .C1(n7073), 
        .C2(P2_U3151), .ZN(P2_U3290) );
  INV_X1 U7688 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n7284) );
  OR2_X1 U7689 ( .A1(n6492), .A2(n6722), .ZN(n6493) );
  XNOR2_X1 U7690 ( .A(n6493), .B(P1_IR_REG_5__SCAN_IN), .ZN(n6869) );
  INV_X1 U7691 ( .A(n6869), .ZN(n10628) );
  OAI222_X1 U7692 ( .A1(n5141), .A2(n7284), .B1(n10517), .B2(n7283), .C1(
        n10628), .C2(P1_U3086), .ZN(P1_U3350) );
  INV_X1 U7693 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n6498) );
  INV_X1 U7694 ( .A(n6496), .ZN(n6497) );
  AOI22_X1 U7695 ( .A1(n6505), .A2(n6498), .B1(n6497), .B2(n6500), .ZN(
        P2_U3376) );
  INV_X1 U7696 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n6502) );
  INV_X1 U7697 ( .A(n6499), .ZN(n6501) );
  AOI22_X1 U7698 ( .A1(n6505), .A2(n6502), .B1(n6501), .B2(n6500), .ZN(
        P2_U3377) );
  INV_X1 U7699 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6504) );
  INV_X1 U7700 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n6503) );
  AND2_X1 U7701 ( .A1(n6492), .A2(n6503), .ZN(n6546) );
  OR2_X1 U7702 ( .A1(n6546), .A2(n6722), .ZN(n6512) );
  XNOR2_X1 U7703 ( .A(n6512), .B(P1_IR_REG_6__SCAN_IN), .ZN(n10648) );
  INV_X1 U7704 ( .A(n10648), .ZN(n6852) );
  OAI222_X1 U7705 ( .A1(n5141), .A2(n6504), .B1(n10517), .B2(n7321), .C1(n6852), .C2(P1_U3086), .ZN(P1_U3349) );
  OAI222_X1 U7706 ( .A1(n9267), .A2(n5322), .B1(n9262), .B2(n7321), .C1(n7077), 
        .C2(P2_U3151), .ZN(P2_U3289) );
  AND2_X1 U7707 ( .A1(n6505), .A2(P2_D_REG_27__SCAN_IN), .ZN(P2_U3238) );
  AND2_X1 U7708 ( .A1(n6505), .A2(P2_D_REG_26__SCAN_IN), .ZN(P2_U3239) );
  AND2_X1 U7709 ( .A1(n6505), .A2(P2_D_REG_23__SCAN_IN), .ZN(P2_U3242) );
  AND2_X1 U7710 ( .A1(n6505), .A2(P2_D_REG_25__SCAN_IN), .ZN(P2_U3240) );
  AND2_X1 U7711 ( .A1(n6505), .A2(P2_D_REG_15__SCAN_IN), .ZN(P2_U3250) );
  AND2_X1 U7712 ( .A1(n6505), .A2(P2_D_REG_14__SCAN_IN), .ZN(P2_U3251) );
  AND2_X1 U7713 ( .A1(n6505), .A2(P2_D_REG_31__SCAN_IN), .ZN(P2_U3234) );
  AND2_X1 U7714 ( .A1(n6505), .A2(P2_D_REG_17__SCAN_IN), .ZN(P2_U3248) );
  AND2_X1 U7715 ( .A1(n6505), .A2(P2_D_REG_16__SCAN_IN), .ZN(P2_U3249) );
  AND2_X1 U7716 ( .A1(n6505), .A2(P2_D_REG_10__SCAN_IN), .ZN(P2_U3255) );
  AND2_X1 U7717 ( .A1(n6505), .A2(P2_D_REG_24__SCAN_IN), .ZN(P2_U3241) );
  AND2_X1 U7718 ( .A1(n6505), .A2(P2_D_REG_21__SCAN_IN), .ZN(P2_U3244) );
  AND2_X1 U7719 ( .A1(n6505), .A2(P2_D_REG_22__SCAN_IN), .ZN(P2_U3243) );
  AND2_X1 U7720 ( .A1(n6505), .A2(P2_D_REG_6__SCAN_IN), .ZN(P2_U3259) );
  AND2_X1 U7721 ( .A1(n6505), .A2(P2_D_REG_5__SCAN_IN), .ZN(P2_U3260) );
  AND2_X1 U7722 ( .A1(n6505), .A2(P2_D_REG_4__SCAN_IN), .ZN(P2_U3261) );
  AND2_X1 U7723 ( .A1(n6505), .A2(P2_D_REG_3__SCAN_IN), .ZN(P2_U3262) );
  AND2_X1 U7724 ( .A1(n6505), .A2(P2_D_REG_2__SCAN_IN), .ZN(P2_U3263) );
  AND2_X1 U7725 ( .A1(n6505), .A2(P2_D_REG_13__SCAN_IN), .ZN(P2_U3252) );
  AND2_X1 U7726 ( .A1(n6505), .A2(P2_D_REG_12__SCAN_IN), .ZN(P2_U3253) );
  AND2_X1 U7727 ( .A1(n6505), .A2(P2_D_REG_11__SCAN_IN), .ZN(P2_U3254) );
  AND2_X1 U7728 ( .A1(n6505), .A2(P2_D_REG_28__SCAN_IN), .ZN(P2_U3237) );
  AND2_X1 U7729 ( .A1(n6505), .A2(P2_D_REG_9__SCAN_IN), .ZN(P2_U3256) );
  AND2_X1 U7730 ( .A1(n6505), .A2(P2_D_REG_8__SCAN_IN), .ZN(P2_U3257) );
  AND2_X1 U7731 ( .A1(n6505), .A2(P2_D_REG_7__SCAN_IN), .ZN(P2_U3258) );
  AND2_X1 U7732 ( .A1(n6505), .A2(P2_D_REG_19__SCAN_IN), .ZN(P2_U3246) );
  AND2_X1 U7733 ( .A1(n6505), .A2(P2_D_REG_20__SCAN_IN), .ZN(P2_U3245) );
  AND2_X1 U7734 ( .A1(n6505), .A2(P2_D_REG_29__SCAN_IN), .ZN(P2_U3236) );
  AND2_X1 U7735 ( .A1(n6505), .A2(P2_D_REG_30__SCAN_IN), .ZN(P2_U3235) );
  AND2_X1 U7736 ( .A1(n6505), .A2(P2_D_REG_18__SCAN_IN), .ZN(P2_U3247) );
  INV_X1 U7737 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6506) );
  OAI222_X1 U7738 ( .A1(n9267), .A2(n6506), .B1(n9262), .B2(n7400), .C1(n5355), 
        .C2(P2_U3151), .ZN(P2_U3288) );
  INV_X1 U7739 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n6510) );
  INV_X1 U7740 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6507) );
  NAND2_X1 U7741 ( .A1(n6512), .A2(n6507), .ZN(n6508) );
  NAND2_X1 U7742 ( .A1(n6508), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6509) );
  XNOR2_X1 U7743 ( .A(n6509), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7401) );
  INV_X1 U7744 ( .A(n7401), .ZN(n10657) );
  OAI222_X1 U7745 ( .A1(n5141), .A2(n6510), .B1(n10517), .B2(n7400), .C1(
        n10657), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U7746 ( .A(n7539), .ZN(n6529) );
  OAI21_X1 U7747 ( .B1(P1_IR_REG_7__SCAN_IN), .B2(P1_IR_REG_6__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6511) );
  NAND2_X1 U7748 ( .A1(n6512), .A2(n6511), .ZN(n6567) );
  INV_X1 U7749 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6513) );
  XNOR2_X1 U7750 ( .A(n6567), .B(n6513), .ZN(n10677) );
  AOI22_X1 U7751 ( .A1(n10677), .A2(P1_STATE_REG_SCAN_IN), .B1(n7489), .B2(
        P2_DATAO_REG_8__SCAN_IN), .ZN(n6514) );
  OAI21_X1 U7752 ( .B1(n6529), .B2(n10517), .A(n6514), .ZN(P1_U3347) );
  NAND2_X1 U7753 ( .A1(n6516), .A2(n10093), .ZN(n10508) );
  NAND2_X2 U7754 ( .A1(n10518), .A2(n6520), .ZN(n6966) );
  NAND2_X1 U7755 ( .A1(n8377), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n6527) );
  INV_X1 U7756 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n8138) );
  OR2_X1 U7757 ( .A1(n5143), .A2(n8138), .ZN(n6526) );
  INV_X1 U7758 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n6519) );
  OR2_X1 U7759 ( .A1(n6968), .A2(n6519), .ZN(n6525) );
  NAND2_X1 U7760 ( .A1(n7024), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7300) );
  NOR2_X1 U7761 ( .A1(n7300), .A2(n7336), .ZN(n7338) );
  NAND2_X1 U7762 ( .A1(n7338), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7412) );
  AND2_X1 U7763 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_REG3_REG_12__SCAN_IN), 
        .ZN(n6523) );
  NAND2_X1 U7764 ( .A1(n7642), .A2(n6523), .ZN(n7760) );
  NAND2_X1 U7765 ( .A1(n7994), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8020) );
  NAND2_X1 U7766 ( .A1(n8021), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n6734) );
  OAI21_X1 U7767 ( .B1(n8021), .B2(P1_REG3_REG_17__SCAN_IN), .A(n6734), .ZN(
        n9331) );
  OR2_X1 U7768 ( .A1(n8382), .A2(n9331), .ZN(n6524) );
  NAND2_X1 U7769 ( .A1(n9669), .A2(P1_DATAO_REG_17__SCAN_IN), .ZN(n6528) );
  OAI21_X1 U7770 ( .B1(n10378), .B2(n9669), .A(n6528), .ZN(P1_U3571) );
  INV_X1 U7771 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6530) );
  OAI222_X1 U7772 ( .A1(n9267), .A2(n6530), .B1(n9262), .B2(n6529), .C1(
        P2_U3151), .C2(n7257), .ZN(P2_U3287) );
  NAND2_X1 U7773 ( .A1(n6817), .A2(n6806), .ZN(n6531) );
  NAND2_X1 U7774 ( .A1(n6531), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6857) );
  INV_X1 U7775 ( .A(n6857), .ZN(n6540) );
  NAND2_X1 U7776 ( .A1(n6535), .A2(n6534), .ZN(n6533) );
  XNOR2_X2 U7777 ( .A(n6537), .B(P1_IR_REG_22__SCAN_IN), .ZN(n6792) );
  XNOR2_X2 U7778 ( .A(n6538), .B(P1_IR_REG_21__SCAN_IN), .ZN(n9655) );
  NAND2_X1 U7779 ( .A1(n6792), .A2(n9655), .ZN(n9469) );
  OR2_X1 U7780 ( .A1(n7913), .A2(n9469), .ZN(n6539) );
  NAND2_X1 U7781 ( .A1(n7322), .A2(n6539), .ZN(n6858) );
  NOR2_X1 U7782 ( .A1(n10942), .A2(n10937), .ZN(P1_U3085) );
  INV_X1 U7783 ( .A(n6541), .ZN(n6569) );
  AOI22_X1 U7784 ( .A1(n8920), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n9256), .ZN(n6542) );
  OAI21_X1 U7785 ( .B1(n6569), .B2(n9262), .A(n6542), .ZN(P2_U3286) );
  INV_X1 U7786 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n6548) );
  NOR2_X1 U7787 ( .A1(P1_IR_REG_9__SCAN_IN), .A2(P1_IR_REG_6__SCAN_IN), .ZN(
        n6543) );
  AND2_X1 U7788 ( .A1(n6544), .A2(n6543), .ZN(n6545) );
  NAND2_X1 U7789 ( .A1(n6546), .A2(n6545), .ZN(n6645) );
  NAND2_X1 U7790 ( .A1(n6645), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6547) );
  XNOR2_X1 U7791 ( .A(n6547), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7525) );
  INV_X1 U7792 ( .A(n7525), .ZN(n9683) );
  OAI222_X1 U7793 ( .A1(n5141), .A2(n6548), .B1(n10517), .B2(n7524), .C1(n9683), .C2(P1_U3086), .ZN(P1_U3345) );
  INV_X1 U7794 ( .A(n10777), .ZN(n8923) );
  INV_X1 U7795 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n6566) );
  OAI222_X1 U7796 ( .A1(P2_U3151), .A2(n8923), .B1(n9267), .B2(n6566), .C1(
        n7524), .C2(n9262), .ZN(P2_U3285) );
  INV_X1 U7797 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6553) );
  INV_X1 U7798 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6551) );
  NAND2_X1 U7799 ( .A1(n6762), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6550) );
  NAND2_X1 U7800 ( .A1(n8377), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6549) );
  OAI211_X1 U7801 ( .C1(n6968), .C2(n6551), .A(n6550), .B(n6549), .ZN(n10170)
         );
  NAND2_X1 U7802 ( .A1(n10170), .A2(n10937), .ZN(n6552) );
  OAI21_X1 U7803 ( .B1(n10937), .B2(n6553), .A(n6552), .ZN(P1_U3585) );
  INV_X1 U7804 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8698) );
  INV_X1 U7805 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n6556) );
  NAND2_X1 U7806 ( .A1(n6762), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n6555) );
  NAND2_X1 U7807 ( .A1(n8377), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n6554) );
  OAI211_X1 U7808 ( .C1(n6968), .C2(n6556), .A(n6555), .B(n6554), .ZN(n10208)
         );
  NAND2_X1 U7809 ( .A1(n10208), .A2(n10937), .ZN(n6557) );
  OAI21_X1 U7810 ( .B1(n8698), .B2(n10937), .A(n6557), .ZN(P1_U3584) );
  NAND2_X1 U7811 ( .A1(n8357), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n6564) );
  INV_X1 U7812 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n6558) );
  OR2_X1 U7813 ( .A1(n6966), .A2(n6558), .ZN(n6563) );
  NOR2_X1 U7814 ( .A1(n7533), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n6559) );
  OR2_X1 U7815 ( .A1(n7642), .A2(n6559), .ZN(n7839) );
  OR2_X1 U7816 ( .A1(n8382), .A2(n7839), .ZN(n6562) );
  INV_X1 U7817 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6560) );
  OR2_X1 U7818 ( .A1(n5143), .A2(n6560), .ZN(n6561) );
  INV_X1 U7819 ( .A(n7884), .ZN(n7776) );
  NAND2_X1 U7820 ( .A1(n7776), .A2(n10937), .ZN(n6565) );
  OAI21_X1 U7821 ( .B1(n6566), .B2(n10937), .A(n6565), .ZN(P1_U3564) );
  INV_X1 U7822 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6570) );
  OAI21_X1 U7823 ( .B1(n6567), .B2(P1_IR_REG_8__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n6568) );
  XNOR2_X1 U7824 ( .A(n6568), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7528) );
  INV_X1 U7825 ( .A(n7528), .ZN(n7362) );
  OAI222_X1 U7826 ( .A1(n5141), .A2(n6570), .B1(n10517), .B2(n6569), .C1(n7362), .C2(P1_U3086), .ZN(P1_U3346) );
  NAND2_X1 U7827 ( .A1(n8071), .A2(P1_B_REG_SCAN_IN), .ZN(n6572) );
  MUX2_X1 U7828 ( .A(n6572), .B(P1_B_REG_SCAN_IN), .S(n6571), .Z(n6573) );
  INV_X1 U7829 ( .A(n8155), .ZN(n6576) );
  INV_X1 U7830 ( .A(n6780), .ZN(n6575) );
  INV_X1 U7831 ( .A(n10506), .ZN(n6786) );
  INV_X1 U7832 ( .A(n10530), .ZN(n10529) );
  NOR2_X1 U7833 ( .A1(n10529), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6577) );
  NOR2_X1 U7834 ( .A1(n6571), .A2(n6576), .ZN(n6771) );
  INV_X1 U7835 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n10097) );
  OAI22_X1 U7836 ( .A1(n6577), .A2(n6771), .B1(n6786), .B2(n10097), .ZN(
        P1_U3439) );
  INV_X1 U7837 ( .A(P2_ADDR_REG_4__SCAN_IN), .ZN(n6624) );
  INV_X1 U7838 ( .A(n6593), .ZN(n6578) );
  NOR2_X2 U7839 ( .A1(P2_U3150), .A2(n6578), .ZN(n10895) );
  INV_X1 U7840 ( .A(n10895), .ZN(n7260) );
  MUX2_X1 U7841 ( .A(P2_REG2_REG_3__SCAN_IN), .B(P2_REG1_REG_3__SCAN_IN), .S(
        n6588), .Z(n6586) );
  INV_X1 U7842 ( .A(n6586), .ZN(n6587) );
  INV_X1 U7843 ( .A(n6613), .ZN(n8848) );
  MUX2_X1 U7844 ( .A(P2_REG2_REG_2__SCAN_IN), .B(P2_REG1_REG_2__SCAN_IN), .S(
        n6580), .Z(n6584) );
  INV_X1 U7845 ( .A(n6584), .ZN(n6585) );
  INV_X1 U7846 ( .A(n6661), .ZN(n6583) );
  MUX2_X1 U7847 ( .A(P2_REG2_REG_1__SCAN_IN), .B(P2_REG1_REG_1__SCAN_IN), .S(
        n6580), .Z(n6579) );
  INV_X1 U7848 ( .A(n6579), .ZN(n6582) );
  XOR2_X1 U7849 ( .A(n6661), .B(n6579), .Z(n6671) );
  INV_X1 U7850 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n6581) );
  MUX2_X1 U7851 ( .A(n6581), .B(n5890), .S(n6580), .Z(n10750) );
  NAND2_X1 U7852 ( .A1(n10750), .A2(n10749), .ZN(n6670) );
  NAND2_X1 U7853 ( .A1(n6671), .A2(n6670), .ZN(n6669) );
  OAI21_X1 U7854 ( .B1(n6583), .B2(n6582), .A(n6669), .ZN(n8847) );
  XOR2_X1 U7855 ( .A(n6613), .B(n6584), .Z(n8846) );
  NAND2_X1 U7856 ( .A1(n8847), .A2(n8846), .ZN(n8845) );
  OAI21_X1 U7857 ( .B1(n8848), .B2(n6585), .A(n8845), .ZN(n6649) );
  XNOR2_X1 U7858 ( .A(n6586), .B(n6651), .ZN(n6650) );
  NOR2_X1 U7859 ( .A1(n6649), .A2(n6650), .ZN(n6648) );
  AOI21_X1 U7860 ( .B1(n5602), .B2(n6587), .A(n6648), .ZN(n6590) );
  MUX2_X1 U7861 ( .A(P2_REG2_REG_4__SCAN_IN), .B(P2_REG1_REG_4__SCAN_IN), .S(
        n6588), .Z(n6698) );
  XOR2_X1 U7862 ( .A(n6704), .B(n6698), .Z(n6589) );
  NAND2_X1 U7863 ( .A1(n6590), .A2(n6589), .ZN(n6699) );
  NAND2_X1 U7864 ( .A1(P2_U3893), .A2(n6306), .ZN(n10772) );
  OAI211_X1 U7865 ( .C1(n6590), .C2(n6589), .A(n6699), .B(n10904), .ZN(n6623)
         );
  OR2_X1 U7866 ( .A1(n6306), .A2(P2_U3151), .ZN(n9264) );
  NOR2_X1 U7867 ( .A1(n6588), .A2(P2_U3151), .ZN(n6591) );
  NAND3_X1 U7868 ( .A1(n6594), .A2(n6591), .A3(n6306), .ZN(n6592) );
  OAI21_X2 U7869 ( .B1(n9264), .B2(n6593), .A(n6592), .ZN(n10896) );
  INV_X1 U7870 ( .A(n10896), .ZN(n8912) );
  INV_X1 U7871 ( .A(n6594), .ZN(n6595) );
  NOR2_X1 U7872 ( .A1(n9264), .A2(n6595), .ZN(n10752) );
  NAND2_X1 U7873 ( .A1(n10752), .A2(n6588), .ZN(n8974) );
  INV_X1 U7874 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n6596) );
  MUX2_X1 U7875 ( .A(P2_REG1_REG_4__SCAN_IN), .B(n6596), .S(n6704), .Z(n6609)
         );
  INV_X1 U7876 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n6597) );
  MUX2_X1 U7877 ( .A(P2_REG1_REG_2__SCAN_IN), .B(n6597), .S(n6613), .Z(n8851)
         );
  NAND2_X1 U7878 ( .A1(n5879), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6602) );
  NAND2_X1 U7879 ( .A1(n6661), .A2(n6602), .ZN(n6601) );
  INV_X1 U7880 ( .A(n10749), .ZN(n6598) );
  NAND2_X1 U7881 ( .A1(n6598), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n6599) );
  OR2_X1 U7882 ( .A1(n6599), .A2(n5879), .ZN(n6600) );
  NAND2_X1 U7883 ( .A1(n6601), .A2(n6600), .ZN(n6660) );
  NAND2_X1 U7884 ( .A1(n6660), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6603) );
  NAND2_X1 U7885 ( .A1(n6603), .A2(n6602), .ZN(n8850) );
  NAND2_X1 U7886 ( .A1(n8851), .A2(n8850), .ZN(n8849) );
  NAND2_X1 U7887 ( .A1(n6613), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6604) );
  NAND2_X1 U7888 ( .A1(n8849), .A2(n6604), .ZN(n6605) );
  XNOR2_X1 U7889 ( .A(n6605), .B(n5602), .ZN(n6652) );
  NAND2_X1 U7890 ( .A1(n6652), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n6607) );
  NAND2_X1 U7891 ( .A1(n6605), .A2(n6651), .ZN(n6606) );
  NAND2_X1 U7892 ( .A1(n6607), .A2(n6606), .ZN(n6608) );
  NAND2_X1 U7893 ( .A1(n6608), .A2(n6609), .ZN(n6706) );
  OAI21_X1 U7894 ( .B1(n6609), .B2(n6608), .A(n6706), .ZN(n6619) );
  INV_X1 U7895 ( .A(n10910), .ZN(n10790) );
  NAND2_X1 U7896 ( .A1(n6704), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6708) );
  OR2_X1 U7897 ( .A1(n6704), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n6610) );
  AND2_X1 U7898 ( .A1(n6708), .A2(n6610), .ZN(n6617) );
  NOR2_X1 U7899 ( .A1(n6581), .A2(n10749), .ZN(n6611) );
  NAND2_X1 U7900 ( .A1(n5879), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n6612) );
  INV_X1 U7901 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6662) );
  NAND2_X1 U7902 ( .A1(n6665), .A2(n6612), .ZN(n8853) );
  NAND2_X1 U7903 ( .A1(n8854), .A2(n8853), .ZN(n8852) );
  NAND2_X1 U7904 ( .A1(n6613), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n6614) );
  NAND2_X1 U7905 ( .A1(n8852), .A2(n6614), .ZN(n6615) );
  OAI21_X1 U7906 ( .B1(n6617), .B2(n6616), .A(n6709), .ZN(n6618) );
  AOI22_X1 U7907 ( .A1(n10905), .A2(n6619), .B1(n10790), .B2(n6618), .ZN(n6620) );
  NAND2_X1 U7908 ( .A1(P2_U3151), .A2(P2_REG3_REG_4__SCAN_IN), .ZN(n6915) );
  OAI211_X1 U7909 ( .C1(n8912), .C2(n6704), .A(n6620), .B(n6915), .ZN(n6621)
         );
  INV_X1 U7910 ( .A(n6621), .ZN(n6622) );
  OAI211_X1 U7911 ( .C1(n6624), .C2(n7260), .A(n6623), .B(n6622), .ZN(P2_U3186) );
  NAND2_X1 U7912 ( .A1(n6640), .A2(n6625), .ZN(n6628) );
  INV_X1 U7913 ( .A(n6687), .ZN(n6633) );
  NAND2_X1 U7914 ( .A1(n6633), .A2(n6626), .ZN(n6627) );
  NAND2_X1 U7915 ( .A1(n6628), .A2(n6627), .ZN(n6636) );
  NAND2_X1 U7916 ( .A1(n6630), .A2(n6629), .ZN(n6631) );
  OAI21_X1 U7917 ( .B1(n6636), .B2(n6631), .A(P2_STATE_REG_SCAN_IN), .ZN(n6635) );
  NOR2_X1 U7918 ( .A1(n7099), .A2(n7129), .ZN(n8692) );
  AND2_X1 U7919 ( .A1(n6632), .A2(P2_STATE_REG_SCAN_IN), .ZN(n7910) );
  AOI21_X1 U7920 ( .B1(n6633), .B2(n8692), .A(n7910), .ZN(n6634) );
  NOR2_X1 U7921 ( .A1(n8819), .A2(P2_U3151), .ZN(n6727) );
  INV_X1 U7922 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10755) );
  NAND2_X1 U7923 ( .A1(n8534), .A2(n8526), .ZN(n8473) );
  INV_X1 U7924 ( .A(n6636), .ZN(n6639) );
  NOR2_X1 U7925 ( .A1(n7099), .A2(n6637), .ZN(n6638) );
  NAND2_X1 U7926 ( .A1(n6640), .A2(n7119), .ZN(n6642) );
  NOR2_X1 U7927 ( .A1(n7099), .A2(n9173), .ZN(n6641) );
  INV_X1 U7928 ( .A(n8805), .ZN(n8823) );
  OAI22_X1 U7929 ( .A1(n5897), .A2(n8803), .B1(n8823), .B2(n6680), .ZN(n6643)
         );
  AOI21_X1 U7930 ( .B1(n8473), .B2(n8810), .A(n6643), .ZN(n6644) );
  OAI21_X1 U7931 ( .B1(n6727), .B2(n10755), .A(n6644), .ZN(P2_U3172) );
  INV_X1 U7932 ( .A(n7634), .ZN(n6693) );
  NAND2_X1 U7933 ( .A1(n6721), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6646) );
  XNOR2_X1 U7934 ( .A(n6646), .B(P1_IR_REG_11__SCAN_IN), .ZN(n10690) );
  AOI22_X1 U7935 ( .A1(n10690), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n7489), .ZN(n6647) );
  OAI21_X1 U7936 ( .B1(n6693), .B2(n10517), .A(n6647), .ZN(P1_U3344) );
  AOI21_X1 U7937 ( .B1(n6650), .B2(n6649), .A(n6648), .ZN(n6659) );
  NAND2_X1 U7938 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_U3151), .ZN(n6757) );
  OAI21_X1 U7939 ( .B1(n8912), .B2(n6651), .A(n6757), .ZN(n6657) );
  XOR2_X1 U7940 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6652), .Z(n6655) );
  AOI21_X1 U7941 ( .B1(n7110), .B2(n6653), .A(n5245), .ZN(n6654) );
  OAI22_X1 U7942 ( .A1(n6655), .A2(n8974), .B1(n10910), .B2(n6654), .ZN(n6656)
         );
  AOI211_X1 U7943 ( .C1(n10895), .C2(P2_ADDR_REG_3__SCAN_IN), .A(n6657), .B(
        n6656), .ZN(n6658) );
  OAI21_X1 U7944 ( .B1(n6659), .B2(n10772), .A(n6658), .ZN(P2_U3185) );
  INV_X1 U7945 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10535) );
  XNOR2_X1 U7946 ( .A(n6660), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n6668) );
  INV_X1 U7947 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n6692) );
  OAI22_X1 U7948 ( .A1(n8912), .A2(n6661), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n6692), .ZN(n6667) );
  NAND2_X1 U7949 ( .A1(n6663), .A2(n6662), .ZN(n6664) );
  AOI21_X1 U7950 ( .B1(n6665), .B2(n6664), .A(n10910), .ZN(n6666) );
  AOI211_X1 U7951 ( .C1(n10905), .C2(n6668), .A(n6667), .B(n6666), .ZN(n6673)
         );
  OAI211_X1 U7952 ( .C1(n6671), .C2(n6670), .A(n6669), .B(n10904), .ZN(n6672)
         );
  OAI211_X1 U7953 ( .C1(n10535), .C2(n7260), .A(n6673), .B(n6672), .ZN(
        P2_U3183) );
  NAND2_X1 U7954 ( .A1(n6675), .A2(n6674), .ZN(n6678) );
  NAND2_X1 U7955 ( .A1(n6676), .A2(n8673), .ZN(n6677) );
  INV_X2 U7956 ( .A(n6752), .ZN(n8424) );
  NAND2_X1 U7957 ( .A1(n8526), .A2(n6681), .ZN(n6684) );
  XNOR2_X1 U7958 ( .A(n6724), .B(n6695), .ZN(n6683) );
  NAND2_X1 U7959 ( .A1(n6684), .A2(n6683), .ZN(n6726) );
  OAI21_X1 U7960 ( .B1(n6684), .B2(n6683), .A(n6726), .ZN(n6685) );
  NAND2_X1 U7961 ( .A1(n6685), .A2(n8810), .ZN(n6691) );
  INV_X1 U7962 ( .A(n6686), .ZN(n6688) );
  NAND3_X1 U7963 ( .A1(n6688), .A2(n6687), .A3(n8692), .ZN(n8816) );
  OAI22_X1 U7964 ( .A1(n7046), .A2(n8803), .B1(n8168), .B2(n8816), .ZN(n6689)
         );
  AOI21_X1 U7965 ( .B1(n8805), .B2(n6682), .A(n6689), .ZN(n6690) );
  OAI211_X1 U7966 ( .C1(n6727), .C2(n6692), .A(n6691), .B(n6690), .ZN(P2_U3162) );
  INV_X1 U7967 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n6694) );
  INV_X1 U7968 ( .A(n10797), .ZN(n8898) );
  OAI222_X1 U7969 ( .A1(n9267), .A2(n6694), .B1(n9262), .B2(n6693), .C1(
        P2_U3151), .C2(n8898), .ZN(P2_U3284) );
  OAI21_X1 U7970 ( .B1(n9130), .B2(n9204), .A(n8473), .ZN(n6696) );
  NAND2_X1 U7971 ( .A1(n6695), .A2(n9133), .ZN(n7125) );
  OAI211_X1 U7972 ( .C1(n9173), .C2(n6680), .A(n6696), .B(n7125), .ZN(n9211)
         );
  NAND2_X1 U7973 ( .A1(n9211), .A2(n11186), .ZN(n6697) );
  OAI21_X1 U7974 ( .B1(n11186), .B2(n5888), .A(n6697), .ZN(P2_U3390) );
  INV_X1 U7975 ( .A(n6704), .ZN(n6701) );
  INV_X1 U7976 ( .A(n6698), .ZN(n6700) );
  OAI21_X1 U7977 ( .B1(n6701), .B2(n6700), .A(n6699), .ZN(n6703) );
  MUX2_X1 U7978 ( .A(P2_REG2_REG_5__SCAN_IN), .B(P2_REG1_REG_5__SCAN_IN), .S(
        n6588), .Z(n7061) );
  XOR2_X1 U7979 ( .A(n7073), .B(n7061), .Z(n6702) );
  NAND2_X1 U7980 ( .A1(n6703), .A2(n6702), .ZN(n7062) );
  OAI211_X1 U7981 ( .C1(n6703), .C2(n6702), .A(n7062), .B(n10904), .ZN(n6719)
         );
  NAND2_X1 U7982 ( .A1(n6704), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n6705) );
  NAND2_X1 U7983 ( .A1(n6706), .A2(n6705), .ZN(n7074) );
  INV_X1 U7984 ( .A(n7073), .ZN(n7064) );
  XNOR2_X1 U7985 ( .A(n7074), .B(n7064), .ZN(n7072) );
  INV_X1 U7986 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n7450) );
  XNOR2_X1 U7987 ( .A(n7072), .B(n7450), .ZN(n6707) );
  NOR2_X1 U7988 ( .A1(n8974), .A2(n6707), .ZN(n6717) );
  NAND2_X1 U7989 ( .A1(n6709), .A2(n6708), .ZN(n6710) );
  NAND2_X1 U7990 ( .A1(n6710), .A2(n7073), .ZN(n10756) );
  AND2_X1 U7991 ( .A1(n6711), .A2(n10756), .ZN(n6712) );
  OAI21_X1 U7992 ( .B1(n6712), .B2(P2_REG2_REG_5__SCAN_IN), .A(n10758), .ZN(
        n6713) );
  INV_X1 U7993 ( .A(n6713), .ZN(n6715) );
  NAND2_X1 U7994 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3151), .ZN(n7036) );
  NAND2_X1 U7995 ( .A1(n10896), .A2(n7064), .ZN(n6714) );
  OAI211_X1 U7996 ( .C1(n10910), .C2(n6715), .A(n7036), .B(n6714), .ZN(n6716)
         );
  AOI211_X1 U7997 ( .C1(n10895), .C2(P2_ADDR_REG_5__SCAN_IN), .A(n6717), .B(
        n6716), .ZN(n6718) );
  NAND2_X1 U7998 ( .A1(n6719), .A2(n6718), .ZN(P2_U3187) );
  INV_X1 U7999 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n6720) );
  OAI222_X1 U8000 ( .A1(n9267), .A2(n6720), .B1(n9262), .B2(n7754), .C1(n8927), 
        .C2(P2_U3151), .ZN(P2_U3283) );
  INV_X1 U8001 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n6723) );
  XNOR2_X1 U8002 ( .A(n6743), .B(P1_IR_REG_12__SCAN_IN), .ZN(n10122) );
  INV_X1 U8003 ( .A(n10122), .ZN(n7368) );
  OAI222_X1 U8004 ( .A1(n5141), .A2(n6723), .B1(n10517), .B2(n7754), .C1(n7368), .C2(P1_U3086), .ZN(P1_U3343) );
  NAND2_X1 U8005 ( .A1(n5897), .A2(n6724), .ZN(n6725) );
  NAND2_X1 U8006 ( .A1(n6726), .A2(n6725), .ZN(n6751) );
  XNOR2_X1 U8007 ( .A(n6730), .B(n6752), .ZN(n6747) );
  XNOR2_X1 U8008 ( .A(n6747), .B(n8844), .ZN(n6750) );
  XOR2_X1 U8009 ( .A(n6751), .B(n6750), .Z(n6732) );
  OAI22_X1 U8010 ( .A1(n5897), .A2(n8816), .B1(n7137), .B2(n8803), .ZN(n6729)
         );
  NOR2_X1 U8011 ( .A1(n6727), .A2(n7116), .ZN(n6728) );
  AOI211_X1 U8012 ( .C1(n8805), .C2(n6730), .A(n6729), .B(n6728), .ZN(n6731)
         );
  OAI21_X1 U8013 ( .B1(n6732), .B2(n8808), .A(n6731), .ZN(P2_U3177) );
  NAND2_X1 U8014 ( .A1(n8357), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6741) );
  INV_X1 U8015 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n6733) );
  OR2_X1 U8016 ( .A1(n6966), .A2(n6733), .ZN(n6740) );
  INV_X2 U8017 ( .A(n6836), .ZN(n8382) );
  NAND2_X1 U8018 ( .A1(n8143), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8142) );
  NAND2_X1 U8019 ( .A1(n8219), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n8218) );
  INV_X1 U8020 ( .A(n6837), .ZN(n8306) );
  INV_X1 U8021 ( .A(n6735), .ZN(n8279) );
  INV_X1 U8022 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6736) );
  NAND2_X1 U8023 ( .A1(n8279), .A2(n6736), .ZN(n6737) );
  NAND2_X1 U8024 ( .A1(n8306), .A2(n6737), .ZN(n10293) );
  OR2_X1 U8025 ( .A1(n8382), .A2(n10293), .ZN(n6739) );
  INV_X1 U8026 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n10294) );
  OR2_X1 U8027 ( .A1(n5143), .A2(n10294), .ZN(n6738) );
  NAND4_X1 U8028 ( .A1(n6741), .A2(n6740), .A3(n6739), .A4(n6738), .ZN(n10453)
         );
  NAND2_X1 U8029 ( .A1(n10453), .A2(n10937), .ZN(n6742) );
  OAI21_X1 U8030 ( .B1(n10937), .B2(n7912), .A(n6742), .ZN(P1_U3577) );
  INV_X1 U8031 ( .A(n7793), .ZN(n6829) );
  NAND2_X1 U8032 ( .A1(n6743), .A2(n9846), .ZN(n6744) );
  NAND2_X1 U8033 ( .A1(n6744), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6745) );
  XNOR2_X1 U8034 ( .A(n6745), .B(P1_IR_REG_13__SCAN_IN), .ZN(n10743) );
  AOI22_X1 U8035 ( .A1(n10743), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7489), .ZN(n6746) );
  OAI21_X1 U8036 ( .B1(n6829), .B2(n10517), .A(n6746), .ZN(P1_U3342) );
  INV_X1 U8037 ( .A(n6747), .ZN(n6748) );
  NOR2_X1 U8038 ( .A1(n6748), .A2(n8844), .ZN(n6749) );
  AOI21_X1 U8039 ( .B1(n6751), .B2(n6750), .A(n6749), .ZN(n6753) );
  XNOR2_X1 U8040 ( .A(n7111), .B(n8440), .ZN(n6907) );
  XNOR2_X1 U8041 ( .A(n6907), .B(n8843), .ZN(n6755) );
  OAI211_X1 U8042 ( .C1(n6753), .C2(n6755), .A(n6754), .B(n8810), .ZN(n6760)
         );
  NAND2_X1 U8043 ( .A1(n8844), .A2(n8800), .ZN(n6756) );
  OAI211_X1 U8044 ( .C1(n7047), .C2(n8803), .A(n6757), .B(n6756), .ZN(n6758)
         );
  AOI21_X1 U8045 ( .B1(n8805), .B2(n7111), .A(n6758), .ZN(n6759) );
  OAI211_X1 U8046 ( .C1(P2_REG3_REG_3__SCAN_IN), .C2(n8756), .A(n6760), .B(
        n6759), .ZN(P2_U3158) );
  INV_X1 U8047 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n6761) );
  NAND2_X1 U8048 ( .A1(n6762), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6766) );
  INV_X1 U8049 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10992) );
  INV_X1 U8050 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n6763) );
  INV_X1 U8051 ( .A(n11007), .ZN(n10963) );
  INV_X1 U8052 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6768) );
  NAND2_X1 U8053 ( .A1(n6780), .A2(n6768), .ZN(n6770) );
  NAND2_X1 U8054 ( .A1(n8155), .A2(n8071), .ZN(n6769) );
  NOR4_X1 U8055 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_16__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_14__SCAN_IN), .ZN(n6775) );
  NOR4_X1 U8056 ( .A1(P1_D_REG_19__SCAN_IN), .A2(P1_D_REG_21__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_18__SCAN_IN), .ZN(n6774) );
  NOR4_X1 U8057 ( .A1(P1_D_REG_9__SCAN_IN), .A2(P1_D_REG_8__SCAN_IN), .A3(
        P1_D_REG_7__SCAN_IN), .A4(P1_D_REG_4__SCAN_IN), .ZN(n6773) );
  NOR4_X1 U8058 ( .A1(P1_D_REG_13__SCAN_IN), .A2(P1_D_REG_12__SCAN_IN), .A3(
        P1_D_REG_11__SCAN_IN), .A4(P1_D_REG_10__SCAN_IN), .ZN(n6772) );
  NAND4_X1 U8059 ( .A1(n6775), .A2(n6774), .A3(n6773), .A4(n6772), .ZN(n6782)
         );
  NOR2_X1 U8060 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n6779) );
  NOR4_X1 U8061 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_5__SCAN_IN), .A3(
        P1_D_REG_31__SCAN_IN), .A4(P1_D_REG_30__SCAN_IN), .ZN(n6778) );
  NOR4_X1 U8062 ( .A1(P1_D_REG_25__SCAN_IN), .A2(P1_D_REG_24__SCAN_IN), .A3(
        P1_D_REG_23__SCAN_IN), .A4(P1_D_REG_22__SCAN_IN), .ZN(n6777) );
  NOR4_X1 U8063 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_28__SCAN_IN), .A3(
        P1_D_REG_27__SCAN_IN), .A4(P1_D_REG_26__SCAN_IN), .ZN(n6776) );
  NAND4_X1 U8064 ( .A1(n6779), .A2(n6778), .A3(n6777), .A4(n6776), .ZN(n6781)
         );
  OAI21_X1 U8065 ( .B1(n6782), .B2(n6781), .A(n6780), .ZN(n7168) );
  NAND3_X1 U8066 ( .A1(n10507), .A2(n7713), .A3(n7168), .ZN(n6824) );
  XNOR2_X2 U8067 ( .A(n6783), .B(P1_IR_REG_20__SCAN_IN), .ZN(n9652) );
  OR2_X1 U8068 ( .A1(n9469), .A2(n9666), .ZN(n9404) );
  INV_X1 U8069 ( .A(n9404), .ZN(n6785) );
  NAND2_X1 U8070 ( .A1(n6786), .A2(n6785), .ZN(n6822) );
  NOR2_X1 U8071 ( .A1(n6824), .A2(n6822), .ZN(n6902) );
  INV_X1 U8072 ( .A(n6902), .ZN(n6788) );
  INV_X1 U8073 ( .A(n5145), .ZN(n6901) );
  NOR2_X1 U8074 ( .A1(n5134), .A2(n6789), .ZN(n6790) );
  XNOR2_X1 U8075 ( .A(n6790), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n10525) );
  MUX2_X1 U8076 ( .A(n5247), .B(n10525), .S(n5133), .Z(n10982) );
  NAND2_X1 U8077 ( .A1(n6792), .A2(n10163), .ZN(n7172) );
  NAND2_X1 U8078 ( .A1(n9655), .A2(n7675), .ZN(n6799) );
  NAND2_X1 U8079 ( .A1(n7172), .A2(n6799), .ZN(n6791) );
  OAI21_X1 U8080 ( .B1(n6792), .B2(n9666), .A(n10995), .ZN(n6793) );
  AND2_X4 U8081 ( .A1(n6949), .A2(n5146), .ZN(n8330) );
  NAND2_X1 U8082 ( .A1(n6836), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6798) );
  INV_X1 U8083 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6794) );
  OR2_X1 U8084 ( .A1(n6966), .A2(n6794), .ZN(n6797) );
  INV_X1 U8085 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10588) );
  OR2_X1 U8086 ( .A1(n5143), .A2(n10588), .ZN(n6796) );
  INV_X1 U8087 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10590) );
  OR2_X1 U8088 ( .A1(n6968), .A2(n10590), .ZN(n6795) );
  NAND2_X1 U8089 ( .A1(n7175), .A2(n8387), .ZN(n6801) );
  NAND2_X1 U8090 ( .A1(n7175), .A2(n8264), .ZN(n6803) );
  OR2_X1 U8091 ( .A1(n10982), .A2(n7325), .ZN(n6802) );
  NAND2_X1 U8092 ( .A1(n6803), .A2(n6802), .ZN(n6805) );
  INV_X1 U8093 ( .A(n6806), .ZN(n6818) );
  AOI21_X1 U8094 ( .B1(n5247), .B2(n10590), .A(n6818), .ZN(n6804) );
  NOR3_X1 U8095 ( .A1(n6888), .A2(n6805), .A3(n6804), .ZN(n6809) );
  NAND2_X1 U8096 ( .A1(n6888), .A2(n6805), .ZN(n6808) );
  NAND3_X1 U8097 ( .A1(n6806), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG1_REG_0__SCAN_IN), .ZN(n6807) );
  INV_X1 U8098 ( .A(n6824), .ZN(n6813) );
  AND2_X1 U8099 ( .A1(n11195), .A2(n9469), .ZN(n6820) );
  INV_X1 U8100 ( .A(n6820), .ZN(n6810) );
  NOR2_X1 U8101 ( .A1(n6810), .A2(n10506), .ZN(n6811) );
  INV_X1 U8102 ( .A(n10982), .ZN(n7176) );
  NAND2_X1 U8103 ( .A1(n6814), .A2(n9652), .ZN(n7188) );
  NOR2_X1 U8104 ( .A1(n10506), .A2(n7188), .ZN(n6812) );
  NAND2_X1 U8105 ( .A1(n6813), .A2(n6812), .ZN(n6815) );
  AOI22_X1 U8106 ( .A1(n10929), .A2(n9376), .B1(n7176), .B2(n9399), .ZN(n6828)
         );
  INV_X1 U8107 ( .A(n9666), .ZN(n6816) );
  OR2_X1 U8108 ( .A1(n9469), .A2(n6816), .ZN(n7165) );
  NAND3_X1 U8109 ( .A1(n6818), .A2(n6817), .A3(n7165), .ZN(n6819) );
  AOI21_X1 U8110 ( .B1(n6824), .B2(n6820), .A(n6819), .ZN(n6821) );
  OR2_X1 U8111 ( .A1(n6821), .A2(P1_U3086), .ZN(n6826) );
  OAI21_X1 U8112 ( .B1(n7188), .B2(P1_U3086), .A(n6822), .ZN(n6823) );
  NAND2_X1 U8113 ( .A1(n6824), .A2(n6823), .ZN(n6825) );
  NAND2_X1 U8114 ( .A1(n9397), .A2(P1_STATE_REG_SCAN_IN), .ZN(n7058) );
  NAND2_X1 U8115 ( .A1(n7058), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6827) );
  OAI211_X1 U8116 ( .C1(n10963), .C2(n9391), .A(n6828), .B(n6827), .ZN(
        P1_U3232) );
  INV_X1 U8117 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6830) );
  OAI222_X1 U8118 ( .A1(n9267), .A2(n6830), .B1(n9262), .B2(n6829), .C1(
        P2_U3151), .C2(n5366), .ZN(P2_U3282) );
  INV_X1 U8119 ( .A(n7987), .ZN(n6882) );
  NOR2_X1 U8120 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6831) );
  NAND2_X1 U8121 ( .A1(n6832), .A2(n6831), .ZN(n7087) );
  NAND2_X1 U8122 ( .A1(n7087), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6833) );
  XNOR2_X1 U8123 ( .A(n6833), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10699) );
  AOI22_X1 U8124 ( .A1(n10699), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n7489), .ZN(n6834) );
  OAI21_X1 U8125 ( .B1(n6882), .B2(n10517), .A(n6834), .ZN(P1_U3341) );
  NAND2_X1 U8126 ( .A1(n8357), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n6842) );
  INV_X1 U8127 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n6835) );
  OR2_X1 U8128 ( .A1(n6966), .A2(n6835), .ZN(n6841) );
  NAND2_X1 U8129 ( .A1(n8359), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n10209) );
  OR2_X1 U8130 ( .A1(n8382), .A2(n10209), .ZN(n6840) );
  INV_X1 U8131 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n6838) );
  OR2_X1 U8132 ( .A1(n5143), .A2(n6838), .ZN(n6839) );
  NAND2_X1 U8133 ( .A1(n9669), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n6843) );
  OAI21_X1 U8134 ( .B1(n10408), .B2(n9669), .A(n6843), .ZN(P1_U3583) );
  NOR2_X1 U8135 ( .A1(P1_REG2_REG_9__SCAN_IN), .A2(n7528), .ZN(n6844) );
  AOI21_X1 U8136 ( .B1(n7528), .B2(P1_REG2_REG_9__SCAN_IN), .A(n6844), .ZN(
        n6856) );
  NAND2_X1 U8137 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n10933) );
  NAND2_X1 U8138 ( .A1(n6846), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6845) );
  OAI21_X1 U8139 ( .B1(n6846), .B2(P1_REG2_REG_1__SCAN_IN), .A(n6845), .ZN(
        n10596) );
  NOR2_X1 U8140 ( .A1(n10933), .A2(n10596), .ZN(n10597) );
  AOI21_X1 U8141 ( .B1(P1_REG2_REG_1__SCAN_IN), .B2(n6846), .A(n10597), .ZN(
        n10915) );
  NAND2_X1 U8142 ( .A1(n6863), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6847) );
  OAI21_X1 U8143 ( .B1(n6863), .B2(P1_REG2_REG_2__SCAN_IN), .A(n6847), .ZN(
        n10916) );
  NOR2_X1 U8144 ( .A1(n10915), .A2(n10916), .ZN(n10917) );
  NAND2_X1 U8145 ( .A1(n10620), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6848) );
  OAI21_X1 U8146 ( .B1(n10620), .B2(P1_REG2_REG_3__SCAN_IN), .A(n6848), .ZN(
        n10613) );
  INV_X1 U8147 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6849) );
  AOI22_X1 U8148 ( .A1(P1_REG2_REG_4__SCAN_IN), .A2(n10948), .B1(n6866), .B2(
        n6849), .ZN(n10944) );
  AOI21_X1 U8149 ( .B1(n6866), .B2(P1_REG2_REG_4__SCAN_IN), .A(n10945), .ZN(
        n10625) );
  NAND2_X1 U8150 ( .A1(P1_REG2_REG_5__SCAN_IN), .A2(n6869), .ZN(n6850) );
  OAI21_X1 U8151 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n6869), .A(n6850), .ZN(
        n10626) );
  INV_X1 U8152 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n6851) );
  AOI22_X1 U8153 ( .A1(P1_REG2_REG_6__SCAN_IN), .A2(n6852), .B1(n10648), .B2(
        n6851), .ZN(n10641) );
  NAND2_X1 U8154 ( .A1(P1_REG2_REG_7__SCAN_IN), .A2(n7401), .ZN(n6853) );
  OAI21_X1 U8155 ( .B1(P1_REG2_REG_7__SCAN_IN), .B2(n7401), .A(n6853), .ZN(
        n10653) );
  NOR2_X1 U8156 ( .A1(n5183), .A2(n10653), .ZN(n10654) );
  NAND2_X1 U8157 ( .A1(n10677), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n6854) );
  OAI21_X1 U8158 ( .B1(n10677), .B2(P1_REG2_REG_8__SCAN_IN), .A(n6854), .ZN(
        n10670) );
  OAI21_X1 U8159 ( .B1(n6856), .B2(n6855), .A(n7355), .ZN(n6880) );
  OR2_X1 U8160 ( .A1(n6858), .A2(n6857), .ZN(n10594) );
  INV_X1 U8161 ( .A(n10594), .ZN(n6860) );
  INV_X1 U8162 ( .A(n10522), .ZN(n10587) );
  NAND2_X1 U8163 ( .A1(n6901), .A2(n10587), .ZN(n10930) );
  INV_X1 U8164 ( .A(n10930), .ZN(n6859) );
  INV_X1 U8165 ( .A(n10958), .ZN(n9685) );
  NAND2_X1 U8166 ( .A1(n6860), .A2(n5145), .ZN(n10949) );
  NOR2_X1 U8167 ( .A1(P1_REG1_REG_9__SCAN_IN), .A2(n7528), .ZN(n6861) );
  AOI21_X1 U8168 ( .B1(n7528), .B2(P1_REG1_REG_9__SCAN_IN), .A(n6861), .ZN(
        n6875) );
  XNOR2_X1 U8169 ( .A(n10600), .B(n10992), .ZN(n10603) );
  NOR3_X1 U8170 ( .A1(n5247), .A2(n10590), .A3(n10603), .ZN(n10601) );
  NOR2_X1 U8171 ( .A1(n10600), .A2(n10992), .ZN(n6862) );
  NOR2_X1 U8172 ( .A1(n10601), .A2(n6862), .ZN(n10923) );
  XNOR2_X1 U8173 ( .A(n6863), .B(P1_REG1_REG_2__SCAN_IN), .ZN(n10922) );
  NOR2_X1 U8174 ( .A1(n10923), .A2(n10922), .ZN(n10921) );
  AOI21_X1 U8175 ( .B1(n6863), .B2(P1_REG1_REG_2__SCAN_IN), .A(n10921), .ZN(
        n10617) );
  NAND2_X1 U8176 ( .A1(n10620), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6864) );
  OAI21_X1 U8177 ( .B1(n10620), .B2(P1_REG1_REG_3__SCAN_IN), .A(n6864), .ZN(
        n10616) );
  NOR2_X1 U8178 ( .A1(n10617), .A2(n10616), .ZN(n10615) );
  INV_X1 U8179 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6865) );
  MUX2_X1 U8180 ( .A(n6865), .B(P1_REG1_REG_4__SCAN_IN), .S(n6866), .Z(n10952)
         );
  NOR2_X1 U8181 ( .A1(n10951), .A2(n10952), .ZN(n10950) );
  AOI21_X1 U8182 ( .B1(n6866), .B2(P1_REG1_REG_4__SCAN_IN), .A(n10950), .ZN(
        n10630) );
  OR2_X1 U8183 ( .A1(n6869), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6868) );
  NAND2_X1 U8184 ( .A1(P1_REG1_REG_5__SCAN_IN), .A2(n6869), .ZN(n6867) );
  NAND2_X1 U8185 ( .A1(n6868), .A2(n6867), .ZN(n10631) );
  NOR2_X1 U8186 ( .A1(n10630), .A2(n10631), .ZN(n10629) );
  INV_X1 U8187 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n6870) );
  MUX2_X1 U8188 ( .A(n6870), .B(P1_REG1_REG_6__SCAN_IN), .S(n10648), .Z(n10644) );
  NOR2_X1 U8189 ( .A1(n10645), .A2(n10644), .ZN(n10643) );
  OR2_X1 U8190 ( .A1(n7401), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6872) );
  NAND2_X1 U8191 ( .A1(P1_REG1_REG_7__SCAN_IN), .A2(n7401), .ZN(n6871) );
  NAND2_X1 U8192 ( .A1(n6872), .A2(n6871), .ZN(n10660) );
  NOR2_X1 U8193 ( .A1(n10659), .A2(n10660), .ZN(n10658) );
  AOI21_X1 U8194 ( .B1(n7401), .B2(P1_REG1_REG_7__SCAN_IN), .A(n10658), .ZN(
        n10674) );
  NAND2_X1 U8195 ( .A1(n10677), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n6873) );
  OAI21_X1 U8196 ( .B1(n10677), .B2(P1_REG1_REG_8__SCAN_IN), .A(n6873), .ZN(
        n10673) );
  NOR2_X1 U8197 ( .A1(n10674), .A2(n10673), .ZN(n10672) );
  NAND2_X1 U8198 ( .A1(n6875), .A2(n6874), .ZN(n7360) );
  OAI21_X1 U8199 ( .B1(n6875), .B2(n6874), .A(n7360), .ZN(n6876) );
  NOR2_X2 U8200 ( .A1(n10594), .A2(n10587), .ZN(n10954) );
  NAND2_X1 U8201 ( .A1(n6876), .A2(n10954), .ZN(n6878) );
  AND2_X1 U8202 ( .A1(P1_U3086), .A2(P1_REG3_REG_9__SCAN_IN), .ZN(n7775) );
  AOI21_X1 U8203 ( .B1(n10942), .B2(P1_ADDR_REG_9__SCAN_IN), .A(n7775), .ZN(
        n6877) );
  OAI211_X1 U8204 ( .C1(n10949), .C2(n7362), .A(n6878), .B(n6877), .ZN(n6879)
         );
  AOI21_X1 U8205 ( .B1(n6880), .B2(n9685), .A(n6879), .ZN(n6881) );
  INV_X1 U8206 ( .A(n6881), .ZN(P1_U3252) );
  INV_X1 U8207 ( .A(n10845), .ZN(n8930) );
  OAI222_X1 U8208 ( .A1(n9267), .A2(n6883), .B1(n9262), .B2(n6882), .C1(
        P2_U3151), .C2(n8930), .ZN(P2_U3281) );
  NAND2_X1 U8209 ( .A1(n11007), .A2(n8264), .ZN(n6887) );
  NAND2_X1 U8210 ( .A1(n9409), .A2(n8387), .ZN(n6886) );
  NAND2_X1 U8211 ( .A1(n6887), .A2(n6886), .ZN(n6941) );
  NOR2_X1 U8212 ( .A1(n6888), .A2(n8346), .ZN(n6889) );
  NAND2_X1 U8213 ( .A1(n11007), .A2(n8387), .ZN(n6890) );
  XNOR2_X1 U8214 ( .A(n6891), .B(n8314), .ZN(n6893) );
  NAND2_X1 U8215 ( .A1(n6892), .A2(n6893), .ZN(n6942) );
  INV_X1 U8216 ( .A(n6892), .ZN(n6895) );
  INV_X1 U8217 ( .A(n6893), .ZN(n6894) );
  NAND2_X1 U8218 ( .A1(n6942), .A2(n6943), .ZN(n6896) );
  XOR2_X1 U8219 ( .A(n6941), .B(n6896), .Z(n6906) );
  INV_X1 U8220 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n7202) );
  INV_X1 U8221 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n6897) );
  INV_X1 U8222 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n11015) );
  OR2_X1 U8223 ( .A1(n6968), .A2(n11015), .ZN(n6899) );
  INV_X1 U8224 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n7201) );
  OR2_X1 U8225 ( .A1(n6983), .A2(n7201), .ZN(n6898) );
  INV_X1 U8226 ( .A(n11020), .ZN(n7186) );
  AOI22_X1 U8227 ( .A1(n9394), .A2(n7175), .B1(n9409), .B2(n9399), .ZN(n6903)
         );
  OAI21_X1 U8228 ( .B1(n7186), .B2(n9391), .A(n6903), .ZN(n6904) );
  AOI21_X1 U8229 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n7058), .A(n6904), .ZN(
        n6905) );
  OAI21_X1 U8230 ( .B1(n6906), .B2(n9402), .A(n6905), .ZN(P1_U3222) );
  XNOR2_X1 U8231 ( .A(n6919), .B(n8424), .ZN(n7032) );
  XNOR2_X1 U8232 ( .A(n7032), .B(n8842), .ZN(n6914) );
  INV_X1 U8233 ( .A(n6907), .ZN(n6908) );
  NAND2_X1 U8234 ( .A1(n6908), .A2(n8843), .ZN(n6909) );
  INV_X1 U8235 ( .A(n7035), .ZN(n6913) );
  AOI21_X1 U8236 ( .B1(n6914), .B2(n6911), .A(n6913), .ZN(n6921) );
  NAND2_X1 U8237 ( .A1(n8841), .A2(n8814), .ZN(n6916) );
  OAI211_X1 U8238 ( .C1(n7137), .C2(n8816), .A(n6916), .B(n6915), .ZN(n6918)
         );
  NOR2_X1 U8239 ( .A1(n8756), .A2(n7310), .ZN(n6917) );
  AOI211_X1 U8240 ( .C1(n8805), .C2(n6919), .A(n6918), .B(n6917), .ZN(n6920)
         );
  OAI21_X1 U8241 ( .B1(n6921), .B2(n8808), .A(n6920), .ZN(P2_U3170) );
  XNOR2_X1 U8242 ( .A(n6922), .B(n8529), .ZN(n7115) );
  NOR2_X1 U8243 ( .A1(n8539), .A2(n9173), .ZN(n7120) );
  OAI21_X1 U8244 ( .B1(n8541), .B2(n6923), .A(n6924), .ZN(n6925) );
  NAND2_X1 U8245 ( .A1(n6925), .A2(n9130), .ZN(n6927) );
  AOI22_X1 U8246 ( .A1(n9136), .A2(n6695), .B1(n8843), .B2(n9133), .ZN(n6926)
         );
  NAND2_X1 U8247 ( .A1(n6927), .A2(n6926), .ZN(n7117) );
  AOI211_X1 U8248 ( .C1(n9204), .C2(n7115), .A(n7120), .B(n7117), .ZN(n11018)
         );
  NAND2_X1 U8249 ( .A1(n9210), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n6928) );
  OAI21_X1 U8250 ( .B1(n11018), .B2(n9210), .A(n6928), .ZN(P2_U3461) );
  NAND2_X1 U8251 ( .A1(n6934), .A2(n8526), .ZN(n6930) );
  NAND2_X1 U8252 ( .A1(n6931), .A2(n6930), .ZN(n7102) );
  NOR2_X1 U8253 ( .A1(n6932), .A2(n9173), .ZN(n6938) );
  OAI21_X1 U8254 ( .B1(n6935), .B2(n6934), .A(n6933), .ZN(n6936) );
  INV_X1 U8255 ( .A(n6936), .ZN(n6937) );
  OAI222_X1 U8256 ( .A1(n9119), .A2(n8168), .B1(n9121), .B2(n7046), .C1(n9116), 
        .C2(n6937), .ZN(n7103) );
  AOI211_X1 U8257 ( .C1(n9204), .C2(n7102), .A(n6938), .B(n7103), .ZN(n10979)
         );
  OR2_X1 U8258 ( .A1(n10979), .A2(n9210), .ZN(n6939) );
  OAI21_X1 U8259 ( .B1(n9206), .B2(n6940), .A(n6939), .ZN(P2_U3460) );
  OR2_X1 U8260 ( .A1(n5139), .A2(n5399), .ZN(n6947) );
  OR2_X1 U8261 ( .A1(n6959), .A2(n6944), .ZN(n6946) );
  OR2_X1 U8262 ( .A1(n7322), .A2(n10920), .ZN(n6945) );
  NAND2_X1 U8263 ( .A1(n11020), .A2(n8387), .ZN(n6948) );
  OAI21_X1 U8264 ( .B1(n11010), .B2(n8330), .A(n6948), .ZN(n6950) );
  XNOR2_X1 U8265 ( .A(n6950), .B(n8346), .ZN(n6954) );
  OR2_X1 U8266 ( .A1(n11010), .A2(n7325), .ZN(n6952) );
  NAND2_X1 U8267 ( .A1(n11020), .A2(n8264), .ZN(n6951) );
  NAND2_X1 U8268 ( .A1(n6952), .A2(n6951), .ZN(n6955) );
  XNOR2_X1 U8269 ( .A(n6954), .B(n6955), .ZN(n7055) );
  INV_X1 U8270 ( .A(n6954), .ZN(n6957) );
  INV_X1 U8271 ( .A(n6955), .ZN(n6956) );
  NAND2_X1 U8272 ( .A1(n6957), .A2(n6956), .ZN(n6994) );
  NAND2_X1 U8273 ( .A1(n7012), .A2(n6994), .ZN(n6977) );
  OR2_X1 U8274 ( .A1(n5139), .A2(n6958), .ZN(n6964) );
  OR2_X1 U8275 ( .A1(n6959), .A2(n6960), .ZN(n6963) );
  OR2_X1 U8276 ( .A1(n7322), .A2(n6961), .ZN(n6962) );
  INV_X1 U8277 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6965) );
  OR2_X1 U8278 ( .A1(n6966), .A2(n6965), .ZN(n6972) );
  INV_X1 U8279 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n7190) );
  OR2_X1 U8280 ( .A1(n5143), .A2(n7190), .ZN(n6971) );
  INV_X1 U8281 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6967) );
  OR2_X1 U8282 ( .A1(n6968), .A2(n6967), .ZN(n6970) );
  OR2_X1 U8283 ( .A1(n6983), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n6969) );
  NAND2_X1 U8284 ( .A1(n11006), .A2(n8387), .ZN(n6973) );
  XNOR2_X1 U8285 ( .A(n6974), .B(n8314), .ZN(n6993) );
  OR2_X1 U8286 ( .A1(n11023), .A2(n7325), .ZN(n6976) );
  NAND2_X1 U8287 ( .A1(n5142), .A2(n8264), .ZN(n6975) );
  NAND2_X1 U8288 ( .A1(n6976), .A2(n6975), .ZN(n6991) );
  XNOR2_X1 U8289 ( .A(n6993), .B(n6991), .ZN(n6996) );
  XNOR2_X1 U8290 ( .A(n6977), .B(n6996), .ZN(n6978) );
  NAND2_X1 U8291 ( .A1(n6978), .A2(n9376), .ZN(n6990) );
  INV_X1 U8292 ( .A(n11023), .ZN(n7268) );
  INV_X1 U8293 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6980) );
  NOR2_X1 U8294 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6980), .ZN(n10622) );
  INV_X1 U8295 ( .A(n9394), .ZN(n9369) );
  INV_X1 U8296 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n6979) );
  OR2_X1 U8297 ( .A1(n6966), .A2(n6979), .ZN(n6986) );
  INV_X1 U8298 ( .A(n7024), .ZN(n6982) );
  INV_X1 U8299 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n7021) );
  NAND2_X1 U8300 ( .A1(n6980), .A2(n7021), .ZN(n6981) );
  NAND2_X1 U8301 ( .A1(n6982), .A2(n6981), .ZN(n7274) );
  OR2_X1 U8302 ( .A1(n6983), .A2(n7274), .ZN(n6985) );
  OR2_X1 U8303 ( .A1(n5143), .A2(n6849), .ZN(n6984) );
  INV_X1 U8304 ( .A(n11019), .ZN(n11046) );
  OAI22_X1 U8305 ( .A1(n9369), .A2(n7186), .B1(n11046), .B2(n9391), .ZN(n6988)
         );
  AOI211_X1 U8306 ( .C1(n7268), .C2(n9399), .A(n10622), .B(n6988), .ZN(n6989)
         );
  OAI211_X1 U8307 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9397), .A(n6990), .B(
        n6989), .ZN(P1_U3218) );
  INV_X1 U8308 ( .A(n6991), .ZN(n6992) );
  NAND2_X1 U8309 ( .A1(n6993), .A2(n6992), .ZN(n6995) );
  AND2_X1 U8310 ( .A1(n6994), .A2(n6995), .ZN(n7011) );
  NAND2_X1 U8311 ( .A1(n7012), .A2(n7011), .ZN(n6998) );
  INV_X1 U8312 ( .A(n6995), .ZN(n6997) );
  AND2_X1 U8313 ( .A1(n6998), .A2(n7014), .ZN(n7010) );
  NAND2_X1 U8314 ( .A1(n11019), .A2(n8387), .ZN(n7006) );
  OR2_X1 U8315 ( .A1(n6959), .A2(n6999), .ZN(n7003) );
  OR2_X1 U8316 ( .A1(n5138), .A2(n7000), .ZN(n7002) );
  OR2_X1 U8317 ( .A1(n5133), .A2(n10948), .ZN(n7001) );
  XNOR2_X1 U8318 ( .A(n7007), .B(n8346), .ZN(n7289) );
  OR2_X1 U8319 ( .A1(n7394), .A2(n7325), .ZN(n7009) );
  NAND2_X1 U8320 ( .A1(n11019), .A2(n8264), .ZN(n7008) );
  NAND2_X1 U8321 ( .A1(n7009), .A2(n7008), .ZN(n7288) );
  AOI21_X1 U8322 ( .B1(n7010), .B2(n7015), .A(n9402), .ZN(n7020) );
  AND2_X1 U8323 ( .A1(n7011), .A2(n7016), .ZN(n7013) );
  NOR2_X1 U8324 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7021), .ZN(n10941) );
  INV_X1 U8325 ( .A(n5142), .ZN(n11036) );
  INV_X1 U8326 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7022) );
  INV_X1 U8327 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7023) );
  OR2_X1 U8328 ( .A1(n6966), .A2(n7023), .ZN(n7027) );
  OAI21_X1 U8329 ( .B1(n7024), .B2(P1_REG3_REG_5__SCAN_IN), .A(n7300), .ZN(
        n7387) );
  OR2_X1 U8330 ( .A1(n8382), .A2(n7387), .ZN(n7026) );
  INV_X1 U8331 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7388) );
  OR2_X1 U8332 ( .A1(n5143), .A2(n7388), .ZN(n7025) );
  NAND4_X1 U8333 ( .A1(n7028), .A2(n7027), .A3(n7026), .A4(n7025), .ZN(n11064)
         );
  OAI22_X1 U8334 ( .A1(n9369), .A2(n11036), .B1(n11035), .B2(n9391), .ZN(n7029) );
  AOI211_X1 U8335 ( .C1(n7004), .C2(n9399), .A(n10941), .B(n7029), .ZN(n7030)
         );
  OAI211_X1 U8336 ( .C1(n9397), .C2(n7274), .A(n7031), .B(n7030), .ZN(P1_U3230) );
  INV_X1 U8337 ( .A(n7032), .ZN(n7033) );
  NAND2_X1 U8338 ( .A1(n7047), .A2(n7033), .ZN(n7034) );
  NAND2_X1 U8339 ( .A1(n7035), .A2(n7034), .ZN(n7230) );
  XNOR2_X1 U8340 ( .A(n7041), .B(n8440), .ZN(n7231) );
  XNOR2_X1 U8341 ( .A(n7231), .B(n8841), .ZN(n7229) );
  XOR2_X1 U8342 ( .A(n7230), .B(n7229), .Z(n7043) );
  NAND2_X1 U8343 ( .A1(n8840), .A2(n8814), .ZN(n7038) );
  NAND2_X1 U8344 ( .A1(n8842), .A2(n8800), .ZN(n7037) );
  NAND3_X1 U8345 ( .A1(n7038), .A2(n7037), .A3(n7036), .ZN(n7040) );
  NOR2_X1 U8346 ( .A1(n8756), .A2(n7492), .ZN(n7039) );
  AOI211_X1 U8347 ( .C1(n8805), .C2(n7041), .A(n7040), .B(n7039), .ZN(n7042)
         );
  OAI21_X1 U8348 ( .B1(n7043), .B2(n8808), .A(n7042), .ZN(P2_U3167) );
  XNOR2_X1 U8349 ( .A(n7044), .B(n8474), .ZN(n7045) );
  OAI222_X1 U8350 ( .A1(n9121), .A2(n7047), .B1(n9119), .B2(n7046), .C1(n9116), 
        .C2(n7045), .ZN(n7108) );
  XOR2_X1 U8351 ( .A(n7048), .B(n8474), .Z(n7114) );
  INV_X1 U8352 ( .A(n9204), .ZN(n9188) );
  OAI22_X1 U8353 ( .A1(n7114), .A2(n9188), .B1(n7049), .B2(n9173), .ZN(n7050)
         );
  NOR2_X1 U8354 ( .A1(n7108), .A2(n7050), .ZN(n11032) );
  INV_X1 U8355 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n7051) );
  OR2_X1 U8356 ( .A1(n9206), .A2(n7051), .ZN(n7052) );
  OAI21_X1 U8357 ( .B1(n11032), .B2(n9210), .A(n7052), .ZN(P2_U3462) );
  INV_X1 U8358 ( .A(n7012), .ZN(n7053) );
  AOI21_X1 U8359 ( .B1(n7055), .B2(n7054), .A(n7053), .ZN(n7060) );
  INV_X1 U8360 ( .A(n11010), .ZN(n7198) );
  AOI22_X1 U8361 ( .A1(n9394), .A2(n11007), .B1(n7198), .B2(n9399), .ZN(n7056)
         );
  OAI21_X1 U8362 ( .B1(n11036), .B2(n9391), .A(n7056), .ZN(n7057) );
  AOI21_X1 U8363 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n7058), .A(n7057), .ZN(
        n7059) );
  OAI21_X1 U8364 ( .B1(n7060), .B2(n9402), .A(n7059), .ZN(P1_U3237) );
  MUX2_X1 U8365 ( .A(P2_REG2_REG_6__SCAN_IN), .B(P2_REG1_REG_6__SCAN_IN), .S(
        n6588), .Z(n7065) );
  INV_X1 U8366 ( .A(n7065), .ZN(n7066) );
  INV_X1 U8367 ( .A(n7061), .ZN(n7063) );
  OAI21_X1 U8368 ( .B1(n7064), .B2(n7063), .A(n7062), .ZN(n10770) );
  XNOR2_X1 U8369 ( .A(n7065), .B(n7077), .ZN(n10771) );
  NOR2_X1 U8370 ( .A1(n10770), .A2(n10771), .ZN(n10769) );
  AOI21_X1 U8371 ( .B1(n5358), .B2(n7066), .A(n10769), .ZN(n7068) );
  MUX2_X1 U8372 ( .A(P2_REG2_REG_7__SCAN_IN), .B(P2_REG1_REG_7__SCAN_IN), .S(
        n6588), .Z(n7212) );
  XOR2_X1 U8373 ( .A(n7215), .B(n7212), .Z(n7067) );
  NOR2_X1 U8374 ( .A1(n7068), .A2(n7067), .ZN(n7213) );
  AOI21_X1 U8375 ( .B1(n7068), .B2(n7067), .A(n7213), .ZN(n7085) );
  XNOR2_X1 U8376 ( .A(n7077), .B(P2_REG2_REG_6__SCAN_IN), .ZN(n10757) );
  OAI21_X1 U8377 ( .B1(n7071), .B2(P2_REG2_REG_7__SCAN_IN), .A(n7222), .ZN(
        n7083) );
  NAND2_X1 U8378 ( .A1(n7072), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n7076) );
  NAND2_X1 U8379 ( .A1(n7074), .A2(n7073), .ZN(n7075) );
  NAND2_X1 U8380 ( .A1(n7076), .A2(n7075), .ZN(n10762) );
  MUX2_X1 U8381 ( .A(P2_REG1_REG_6__SCAN_IN), .B(n7078), .S(n7077), .Z(n10763)
         );
  XOR2_X1 U8382 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n7209), .Z(n7079) );
  NOR2_X1 U8383 ( .A1(n7079), .A2(n8974), .ZN(n7082) );
  NAND2_X1 U8384 ( .A1(n10895), .A2(P2_ADDR_REG_7__SCAN_IN), .ZN(n7080) );
  NAND2_X1 U8385 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_U3151), .ZN(n7432) );
  OAI211_X1 U8386 ( .C1(n8912), .C2(n5355), .A(n7080), .B(n7432), .ZN(n7081)
         );
  AOI211_X1 U8387 ( .C1(n7083), .C2(n10790), .A(n7082), .B(n7081), .ZN(n7084)
         );
  OAI21_X1 U8388 ( .B1(n7085), .B2(n10772), .A(n7084), .ZN(P2_U3189) );
  INV_X1 U8389 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n7086) );
  INV_X1 U8390 ( .A(n8030), .ZN(n7090) );
  OAI222_X1 U8391 ( .A1(n9267), .A2(n7086), .B1(n9262), .B2(n7090), .C1(n8933), 
        .C2(P2_U3151), .ZN(P2_U3280) );
  INV_X1 U8392 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7091) );
  NAND2_X1 U8393 ( .A1(n7088), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7453) );
  INV_X1 U8394 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9853) );
  NAND2_X1 U8395 ( .A1(n7453), .A2(n9853), .ZN(n7141) );
  OR2_X1 U8396 ( .A1(n7453), .A2(n9853), .ZN(n7089) );
  OAI222_X1 U8397 ( .A1(n5141), .A2(n7091), .B1(n10517), .B2(n7090), .C1(n5387), .C2(P1_U3086), .ZN(P1_U3340) );
  INV_X1 U8398 ( .A(n7092), .ZN(n7093) );
  NAND2_X1 U8399 ( .A1(n7093), .A2(n6675), .ZN(n7094) );
  OAI21_X1 U8400 ( .B1(n7096), .B2(n7095), .A(n7094), .ZN(n7097) );
  NAND2_X1 U8401 ( .A1(n7098), .A2(n7097), .ZN(n7128) );
  NOR2_X1 U8402 ( .A1(n5140), .A2(n7119), .ZN(n7491) );
  INV_X1 U8403 ( .A(n7491), .ZN(n7100) );
  NAND2_X1 U8404 ( .A1(n7734), .A2(n7100), .ZN(n7101) );
  INV_X1 U8405 ( .A(n7102), .ZN(n7107) );
  INV_X1 U8406 ( .A(n7103), .ZN(n7104) );
  MUX2_X1 U8407 ( .A(n6662), .B(n7104), .S(n9145), .Z(n7106) );
  INV_X1 U8408 ( .A(n9141), .ZN(n9111) );
  AOI22_X1 U8409 ( .A1(n9111), .A2(n6682), .B1(P2_REG3_REG_1__SCAN_IN), .B2(
        n9125), .ZN(n7105) );
  OAI211_X1 U8410 ( .C1(n9114), .C2(n7107), .A(n7106), .B(n7105), .ZN(P2_U3232) );
  INV_X1 U8411 ( .A(n7108), .ZN(n7109) );
  MUX2_X1 U8412 ( .A(n7110), .B(n7109), .S(n9145), .Z(n7113) );
  AOI22_X1 U8413 ( .A1(n9111), .A2(n7111), .B1(n9125), .B2(n9959), .ZN(n7112)
         );
  OAI211_X1 U8414 ( .C1(n9114), .C2(n7114), .A(n7113), .B(n7112), .ZN(P2_U3230) );
  INV_X1 U8415 ( .A(n7115), .ZN(n7124) );
  NOR2_X1 U8416 ( .A1(n9142), .A2(n7116), .ZN(n7118) );
  AOI211_X1 U8417 ( .C1(n7120), .C2(n7119), .A(n7118), .B(n7117), .ZN(n7121)
         );
  MUX2_X1 U8418 ( .A(n7122), .B(n7121), .S(n9145), .Z(n7123) );
  OAI21_X1 U8419 ( .B1(n7124), .B2(n9114), .A(n7123), .ZN(P2_U3231) );
  OAI22_X1 U8420 ( .A1(n9141), .A2(n6680), .B1(n10755), .B2(n9142), .ZN(n7127)
         );
  NOR2_X1 U8421 ( .A1(n7125), .A2(n9150), .ZN(n7126) );
  AOI211_X1 U8422 ( .C1(n9150), .C2(P2_REG2_REG_0__SCAN_IN), .A(n7127), .B(
        n7126), .ZN(n7132) );
  INV_X1 U8423 ( .A(n7128), .ZN(n7130) );
  NAND4_X1 U8424 ( .A1(n8473), .A2(n7130), .A3(n9173), .A4(n7129), .ZN(n7131)
         );
  NAND2_X1 U8425 ( .A1(n7132), .A2(n7131), .ZN(P2_U3233) );
  OAI21_X1 U8426 ( .B1(n7134), .B2(n8545), .A(n7133), .ZN(n7315) );
  NOR2_X1 U8427 ( .A1(n7311), .A2(n9173), .ZN(n7138) );
  XNOR2_X1 U8428 ( .A(n7135), .B(n8545), .ZN(n7136) );
  OAI222_X1 U8429 ( .A1(n9119), .A2(n7137), .B1(n9121), .B2(n7349), .C1(n9116), 
        .C2(n7136), .ZN(n7312) );
  AOI211_X1 U8430 ( .C1(n9204), .C2(n7315), .A(n7138), .B(n7312), .ZN(n11034)
         );
  NAND2_X1 U8431 ( .A1(n9210), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n7139) );
  OAI21_X1 U8432 ( .B1(n11034), .B2(n9210), .A(n7139), .ZN(P2_U3463) );
  INV_X1 U8433 ( .A(n8084), .ZN(n7143) );
  OAI222_X1 U8434 ( .A1(n9267), .A2(n7140), .B1(n9262), .B2(n7143), .C1(
        P2_U3151), .C2(n8938), .ZN(P2_U3279) );
  NAND2_X1 U8435 ( .A1(n7141), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7142) );
  XNOR2_X1 U8436 ( .A(n7142), .B(P1_IR_REG_16__SCAN_IN), .ZN(n10140) );
  INV_X1 U8437 ( .A(n10140), .ZN(n10120) );
  OAI222_X1 U8438 ( .A1(n5141), .A2(n10025), .B1(n10517), .B2(n7143), .C1(
        P1_U3086), .C2(n10120), .ZN(P1_U3339) );
  NOR2_X1 U8439 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(P1_ADDR_REG_18__SCAN_IN), 
        .ZN(n7144) );
  AOI21_X1 U8440 ( .B1(P1_ADDR_REG_18__SCAN_IN), .B2(P2_ADDR_REG_18__SCAN_IN), 
        .A(n7144), .ZN(n10586) );
  NOR2_X1 U8441 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n7145) );
  AOI21_X1 U8442 ( .B1(P1_ADDR_REG_17__SCAN_IN), .B2(P2_ADDR_REG_17__SCAN_IN), 
        .A(n7145), .ZN(n10583) );
  NOR2_X1 U8443 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n7146) );
  AOI21_X1 U8444 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(P2_ADDR_REG_16__SCAN_IN), 
        .A(n7146), .ZN(n10580) );
  NOR2_X1 U8445 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n7147) );
  AOI21_X1 U8446 ( .B1(P1_ADDR_REG_15__SCAN_IN), .B2(P2_ADDR_REG_15__SCAN_IN), 
        .A(n7147), .ZN(n10577) );
  NOR2_X1 U8447 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n7148) );
  AOI21_X1 U8448 ( .B1(P1_ADDR_REG_14__SCAN_IN), .B2(P2_ADDR_REG_14__SCAN_IN), 
        .A(n7148), .ZN(n10574) );
  NOR2_X1 U8449 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n7149) );
  AOI21_X1 U8450 ( .B1(P1_ADDR_REG_13__SCAN_IN), .B2(P2_ADDR_REG_13__SCAN_IN), 
        .A(n7149), .ZN(n10571) );
  NOR2_X1 U8451 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n7150) );
  AOI21_X1 U8452 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(P2_ADDR_REG_12__SCAN_IN), 
        .A(n7150), .ZN(n10568) );
  NOR2_X1 U8453 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n7151) );
  AOI21_X1 U8454 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(P2_ADDR_REG_11__SCAN_IN), 
        .A(n7151), .ZN(n10565) );
  NOR2_X1 U8455 ( .A1(P1_ADDR_REG_10__SCAN_IN), .A2(P2_ADDR_REG_10__SCAN_IN), 
        .ZN(n7152) );
  AOI21_X1 U8456 ( .B1(P2_ADDR_REG_10__SCAN_IN), .B2(P1_ADDR_REG_10__SCAN_IN), 
        .A(n7152), .ZN(n10562) );
  NOR2_X1 U8457 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(P1_ADDR_REG_9__SCAN_IN), 
        .ZN(n7153) );
  AOI21_X1 U8458 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(P2_ADDR_REG_9__SCAN_IN), 
        .A(n7153), .ZN(n10559) );
  NOR2_X1 U8459 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(P1_ADDR_REG_8__SCAN_IN), 
        .ZN(n7154) );
  AOI21_X1 U8460 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(P2_ADDR_REG_8__SCAN_IN), 
        .A(n7154), .ZN(n10556) );
  NOR2_X1 U8461 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(P1_ADDR_REG_7__SCAN_IN), 
        .ZN(n7155) );
  AOI21_X1 U8462 ( .B1(P1_ADDR_REG_7__SCAN_IN), .B2(P2_ADDR_REG_7__SCAN_IN), 
        .A(n7155), .ZN(n10553) );
  NOR2_X1 U8463 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(P1_ADDR_REG_6__SCAN_IN), 
        .ZN(n7156) );
  AOI21_X1 U8464 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(P2_ADDR_REG_6__SCAN_IN), 
        .A(n7156), .ZN(n10550) );
  NOR2_X1 U8465 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(P1_ADDR_REG_5__SCAN_IN), 
        .ZN(n7157) );
  AOI21_X1 U8466 ( .B1(P1_ADDR_REG_5__SCAN_IN), .B2(P2_ADDR_REG_5__SCAN_IN), 
        .A(n7157), .ZN(n10547) );
  AND2_X1 U8467 ( .A1(P2_ADDR_REG_0__SCAN_IN), .A2(P1_ADDR_REG_0__SCAN_IN), 
        .ZN(n7158) );
  NOR2_X1 U8468 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n7158), .ZN(n10532) );
  INV_X1 U8469 ( .A(n10532), .ZN(n10533) );
  NAND3_X1 U8470 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10534) );
  NAND2_X1 U8471 ( .A1(n10535), .A2(n10534), .ZN(n10531) );
  NAND2_X1 U8472 ( .A1(n10533), .A2(n10531), .ZN(n10538) );
  NAND2_X1 U8473 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n7159) );
  OAI21_X1 U8474 ( .B1(P1_ADDR_REG_2__SCAN_IN), .B2(P2_ADDR_REG_2__SCAN_IN), 
        .A(n7159), .ZN(n10537) );
  NOR2_X1 U8475 ( .A1(n10538), .A2(n10537), .ZN(n10536) );
  AOI21_X1 U8476 ( .B1(P2_ADDR_REG_2__SCAN_IN), .B2(P1_ADDR_REG_2__SCAN_IN), 
        .A(n10536), .ZN(n10541) );
  NAND2_X1 U8477 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n7160) );
  OAI21_X1 U8478 ( .B1(P2_ADDR_REG_3__SCAN_IN), .B2(P1_ADDR_REG_3__SCAN_IN), 
        .A(n7160), .ZN(n10540) );
  NOR2_X1 U8479 ( .A1(n10541), .A2(n10540), .ZN(n10539) );
  AOI21_X1 U8480 ( .B1(P1_ADDR_REG_3__SCAN_IN), .B2(P2_ADDR_REG_3__SCAN_IN), 
        .A(n10539), .ZN(n10544) );
  NOR2_X1 U8481 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n7161) );
  AOI21_X1 U8482 ( .B1(P2_ADDR_REG_4__SCAN_IN), .B2(P1_ADDR_REG_4__SCAN_IN), 
        .A(n7161), .ZN(n10543) );
  NAND2_X1 U8483 ( .A1(n10544), .A2(n10543), .ZN(n10542) );
  OAI21_X1 U8484 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(P2_ADDR_REG_4__SCAN_IN), 
        .A(n10542), .ZN(n10546) );
  NAND2_X1 U8485 ( .A1(n10547), .A2(n10546), .ZN(n10545) );
  OAI21_X1 U8486 ( .B1(P2_ADDR_REG_5__SCAN_IN), .B2(P1_ADDR_REG_5__SCAN_IN), 
        .A(n10545), .ZN(n10549) );
  NAND2_X1 U8487 ( .A1(n10550), .A2(n10549), .ZN(n10548) );
  OAI21_X1 U8488 ( .B1(P2_ADDR_REG_6__SCAN_IN), .B2(P1_ADDR_REG_6__SCAN_IN), 
        .A(n10548), .ZN(n10552) );
  NAND2_X1 U8489 ( .A1(n10553), .A2(n10552), .ZN(n10551) );
  OAI21_X1 U8490 ( .B1(P2_ADDR_REG_7__SCAN_IN), .B2(P1_ADDR_REG_7__SCAN_IN), 
        .A(n10551), .ZN(n10555) );
  NAND2_X1 U8491 ( .A1(n10556), .A2(n10555), .ZN(n10554) );
  OAI21_X1 U8492 ( .B1(P2_ADDR_REG_8__SCAN_IN), .B2(P1_ADDR_REG_8__SCAN_IN), 
        .A(n10554), .ZN(n10558) );
  NAND2_X1 U8493 ( .A1(n10559), .A2(n10558), .ZN(n10557) );
  OAI21_X1 U8494 ( .B1(P2_ADDR_REG_9__SCAN_IN), .B2(P1_ADDR_REG_9__SCAN_IN), 
        .A(n10557), .ZN(n10561) );
  NAND2_X1 U8495 ( .A1(n10562), .A2(n10561), .ZN(n10560) );
  OAI21_X1 U8496 ( .B1(P1_ADDR_REG_10__SCAN_IN), .B2(P2_ADDR_REG_10__SCAN_IN), 
        .A(n10560), .ZN(n10564) );
  NAND2_X1 U8497 ( .A1(n10565), .A2(n10564), .ZN(n10563) );
  OAI21_X1 U8498 ( .B1(P2_ADDR_REG_11__SCAN_IN), .B2(P1_ADDR_REG_11__SCAN_IN), 
        .A(n10563), .ZN(n10567) );
  NAND2_X1 U8499 ( .A1(n10568), .A2(n10567), .ZN(n10566) );
  OAI21_X1 U8500 ( .B1(P2_ADDR_REG_12__SCAN_IN), .B2(P1_ADDR_REG_12__SCAN_IN), 
        .A(n10566), .ZN(n10570) );
  NAND2_X1 U8501 ( .A1(n10571), .A2(n10570), .ZN(n10569) );
  OAI21_X1 U8502 ( .B1(P2_ADDR_REG_13__SCAN_IN), .B2(P1_ADDR_REG_13__SCAN_IN), 
        .A(n10569), .ZN(n10573) );
  NAND2_X1 U8503 ( .A1(n10574), .A2(n10573), .ZN(n10572) );
  OAI21_X1 U8504 ( .B1(P2_ADDR_REG_14__SCAN_IN), .B2(P1_ADDR_REG_14__SCAN_IN), 
        .A(n10572), .ZN(n10576) );
  NAND2_X1 U8505 ( .A1(n10577), .A2(n10576), .ZN(n10575) );
  OAI21_X1 U8506 ( .B1(P2_ADDR_REG_15__SCAN_IN), .B2(P1_ADDR_REG_15__SCAN_IN), 
        .A(n10575), .ZN(n10579) );
  NAND2_X1 U8507 ( .A1(n10580), .A2(n10579), .ZN(n10578) );
  OAI21_X1 U8508 ( .B1(P2_ADDR_REG_16__SCAN_IN), .B2(P1_ADDR_REG_16__SCAN_IN), 
        .A(n10578), .ZN(n10582) );
  NAND2_X1 U8509 ( .A1(n10583), .A2(n10582), .ZN(n10581) );
  OAI21_X1 U8510 ( .B1(P2_ADDR_REG_17__SCAN_IN), .B2(P1_ADDR_REG_17__SCAN_IN), 
        .A(n10581), .ZN(n10585) );
  NAND2_X1 U8511 ( .A1(n10586), .A2(n10585), .ZN(n10584) );
  OAI21_X1 U8512 ( .B1(P2_ADDR_REG_18__SCAN_IN), .B2(P1_ADDR_REG_18__SCAN_IN), 
        .A(n10584), .ZN(n7164) );
  XNOR2_X1 U8513 ( .A(n7162), .B(P1_ADDR_REG_19__SCAN_IN), .ZN(n7163) );
  XNOR2_X1 U8514 ( .A(n7164), .B(n7163), .ZN(ADD_1068_U4) );
  INV_X1 U8515 ( .A(n7713), .ZN(n7169) );
  INV_X1 U8516 ( .A(n7165), .ZN(n7166) );
  NOR2_X1 U8517 ( .A1(n10506), .A2(n7166), .ZN(n7167) );
  NAND2_X1 U8518 ( .A1(n7722), .A2(n10507), .ZN(n7170) );
  AND2_X1 U8519 ( .A1(n9404), .A2(n10964), .ZN(n10971) );
  NAND2_X1 U8520 ( .A1(n7172), .A2(n9666), .ZN(n7173) );
  NAND2_X1 U8521 ( .A1(n10971), .A2(n7173), .ZN(n10984) );
  NAND2_X1 U8522 ( .A1(n10984), .A2(n10995), .ZN(n7174) );
  XNOR2_X2 U8523 ( .A(n11007), .B(n9409), .ZN(n10985) );
  AND2_X1 U8524 ( .A1(n7176), .A2(n7175), .ZN(n10980) );
  OR2_X1 U8525 ( .A1(n11020), .A2(n11010), .ZN(n9536) );
  NAND2_X1 U8526 ( .A1(n11010), .A2(n11020), .ZN(n9540) );
  NAND2_X1 U8527 ( .A1(n9536), .A2(n9540), .ZN(n7179) );
  NAND2_X1 U8528 ( .A1(n11023), .A2(n5142), .ZN(n9541) );
  INV_X1 U8529 ( .A(n7269), .ZN(n9480) );
  XNOR2_X1 U8530 ( .A(n7270), .B(n9480), .ZN(n11027) );
  NOR2_X1 U8531 ( .A1(n7175), .A2(n10982), .ZN(n9477) );
  NAND2_X1 U8532 ( .A1(n10985), .A2(n9477), .ZN(n7178) );
  NAND2_X1 U8533 ( .A1(n10963), .A2(n9409), .ZN(n7177) );
  NAND2_X1 U8534 ( .A1(n7178), .A2(n7177), .ZN(n9542) );
  NAND2_X1 U8535 ( .A1(n9542), .A2(n7180), .ZN(n9539) );
  NAND2_X1 U8536 ( .A1(n9539), .A2(n9536), .ZN(n7181) );
  NAND2_X1 U8537 ( .A1(n7181), .A2(n7269), .ZN(n7280) );
  OAI21_X1 U8538 ( .B1(n7269), .B2(n7181), .A(n7280), .ZN(n7184) );
  NAND2_X1 U8539 ( .A1(n6792), .A2(n10158), .ZN(n7183) );
  NAND2_X1 U8540 ( .A1(n9655), .A2(n9652), .ZN(n7182) );
  NAND2_X1 U8541 ( .A1(n7184), .A2(n11181), .ZN(n11025) );
  INV_X1 U8542 ( .A(n11025), .ZN(n7195) );
  NAND2_X1 U8543 ( .A1(n10983), .A2(n10982), .ZN(n10981) );
  AOI21_X1 U8544 ( .B1(n7199), .B2(n7268), .A(n11212), .ZN(n7185) );
  NAND2_X1 U8545 ( .A1(n7185), .A2(n7271), .ZN(n11022) );
  NAND2_X1 U8546 ( .A1(n10367), .A2(n11172), .ZN(n10213) );
  OAI22_X1 U8547 ( .A1(n10333), .A2(n11022), .B1(n7186), .B2(n10213), .ZN(
        n7194) );
  INV_X1 U8548 ( .A(n9469), .ZN(n7187) );
  NAND2_X1 U8549 ( .A1(n10367), .A2(n11169), .ZN(n10328) );
  INV_X1 U8550 ( .A(n7188), .ZN(n7189) );
  INV_X1 U8551 ( .A(n7171), .ZN(n10358) );
  OAI22_X1 U8552 ( .A1(n10358), .A2(n7190), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n10968), .ZN(n7191) );
  AOI21_X1 U8553 ( .B1(n11124), .B2(n7268), .A(n7191), .ZN(n7192) );
  OAI21_X1 U8554 ( .B1(n11046), .B2(n10328), .A(n7192), .ZN(n7193) );
  AOI211_X1 U8555 ( .C1(n7195), .C2(n10367), .A(n7194), .B(n7193), .ZN(n7196)
         );
  OAI21_X1 U8556 ( .B1(n10391), .B2(n11027), .A(n7196), .ZN(P1_U3290) );
  NAND2_X1 U8557 ( .A1(n10367), .A2(n11181), .ZN(n10233) );
  XNOR2_X1 U8558 ( .A(n9542), .B(n7179), .ZN(n11011) );
  XNOR2_X1 U8559 ( .A(n7197), .B(n7179), .ZN(n11014) );
  INV_X1 U8560 ( .A(n10213), .ZN(n10326) );
  AOI22_X1 U8561 ( .A1(n10326), .A2(n11007), .B1(n11124), .B2(n7198), .ZN(
        n7206) );
  AOI21_X1 U8562 ( .B1(n10981), .B2(n7198), .A(n11212), .ZN(n7200) );
  NAND2_X1 U8563 ( .A1(n7200), .A2(n7199), .ZN(n11009) );
  INV_X1 U8564 ( .A(n11009), .ZN(n7204) );
  OAI22_X1 U8565 ( .A1(n10367), .A2(n7202), .B1(n7201), .B2(n10968), .ZN(n7203) );
  AOI21_X1 U8566 ( .B1(n11128), .B2(n7204), .A(n7203), .ZN(n7205) );
  OAI211_X1 U8567 ( .C1(n11036), .C2(n10328), .A(n7206), .B(n7205), .ZN(n7207)
         );
  AOI21_X1 U8568 ( .B1(n11129), .B2(n11014), .A(n7207), .ZN(n7208) );
  OAI21_X1 U8569 ( .B1(n10233), .B2(n11011), .A(n7208), .ZN(P1_U3291) );
  MUX2_X1 U8570 ( .A(P2_REG1_REG_8__SCAN_IN), .B(n6004), .S(n7219), .Z(n7211)
         );
  NOR2_X1 U8571 ( .A1(n7210), .A2(n7211), .ZN(n7255) );
  AOI21_X1 U8572 ( .B1(n7211), .B2(n7210), .A(n7255), .ZN(n7228) );
  INV_X1 U8573 ( .A(n7212), .ZN(n7214) );
  AOI21_X1 U8574 ( .B1(n7215), .B2(n7214), .A(n7213), .ZN(n7249) );
  MUX2_X1 U8575 ( .A(P2_REG2_REG_8__SCAN_IN), .B(P2_REG1_REG_8__SCAN_IN), .S(
        n6588), .Z(n7247) );
  XOR2_X1 U8576 ( .A(n7219), .B(n7247), .Z(n7248) );
  XNOR2_X1 U8577 ( .A(n7249), .B(n7248), .ZN(n7216) );
  NAND2_X1 U8578 ( .A1(n7216), .A2(n10904), .ZN(n7227) );
  NAND2_X1 U8579 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3151), .ZN(n7217) );
  OAI21_X1 U8580 ( .B1(n8912), .B2(n7257), .A(n7217), .ZN(n7225) );
  MUX2_X1 U8581 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n5607), .S(n7219), .Z(n7221)
         );
  NAND3_X1 U8582 ( .A1(n7222), .A2(n7221), .A3(n7220), .ZN(n7223) );
  AOI21_X1 U8583 ( .B1(n5244), .B2(n7223), .A(n10910), .ZN(n7224) );
  AOI211_X1 U8584 ( .C1(n10895), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n7225), .B(
        n7224), .ZN(n7226) );
  OAI211_X1 U8585 ( .C1(n7228), .C2(n8974), .A(n7227), .B(n7226), .ZN(P2_U3190) );
  XNOR2_X1 U8586 ( .A(n7518), .B(n8424), .ZN(n7426) );
  XNOR2_X1 U8587 ( .A(n7426), .B(n8840), .ZN(n7238) );
  NAND2_X1 U8588 ( .A1(n7230), .A2(n7229), .ZN(n7233) );
  NAND2_X1 U8589 ( .A1(n7349), .A2(n7231), .ZN(n7232) );
  NAND2_X1 U8590 ( .A1(n7233), .A2(n7232), .ZN(n7237) );
  INV_X1 U8591 ( .A(n7237), .ZN(n7235) );
  INV_X1 U8592 ( .A(n7428), .ZN(n7236) );
  AOI211_X1 U8593 ( .C1(n7238), .C2(n7237), .A(n8808), .B(n7236), .ZN(n7246)
         );
  INV_X1 U8594 ( .A(n7239), .ZN(n7517) );
  NAND2_X1 U8595 ( .A1(n8819), .A2(n7517), .ZN(n7244) );
  INV_X1 U8596 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n7240) );
  NOR2_X1 U8597 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7240), .ZN(n10765) );
  AOI21_X1 U8598 ( .B1(n8841), .B2(n8800), .A(n10765), .ZN(n7243) );
  NAND2_X1 U8599 ( .A1(n8805), .A2(n7518), .ZN(n7242) );
  NAND2_X1 U8600 ( .A1(n8839), .A2(n8814), .ZN(n7241) );
  NAND4_X1 U8601 ( .A1(n7244), .A2(n7243), .A3(n7242), .A4(n7241), .ZN(n7245)
         );
  OR2_X1 U8602 ( .A1(n7246), .A2(n7245), .ZN(P2_U3179) );
  OAI22_X1 U8603 ( .A1(n7249), .A2(n7248), .B1(n7247), .B2(n7257), .ZN(n8892)
         );
  INV_X1 U8604 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8921) );
  OR2_X1 U8605 ( .A1(n6588), .A2(n8921), .ZN(n7251) );
  NAND2_X1 U8606 ( .A1(n6588), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n7250) );
  AND3_X1 U8607 ( .A1(n7251), .A2(n7250), .A3(n8920), .ZN(n8891) );
  INV_X1 U8608 ( .A(n8891), .ZN(n7253) );
  AOI21_X1 U8609 ( .B1(n6588), .B2(n6022), .A(n8920), .ZN(n7252) );
  OAI21_X1 U8610 ( .B1(n6588), .B2(P2_REG2_REG_9__SCAN_IN), .A(n7252), .ZN(
        n8893) );
  NAND2_X1 U8611 ( .A1(n7253), .A2(n8893), .ZN(n7254) );
  XNOR2_X1 U8612 ( .A(n8892), .B(n7254), .ZN(n7267) );
  OAI21_X1 U8613 ( .B1(n7256), .B2(P2_REG1_REG_9__SCAN_IN), .A(n8862), .ZN(
        n7265) );
  XOR2_X1 U8614 ( .A(n8921), .B(n8922), .Z(n7263) );
  NOR2_X1 U8615 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n7258), .ZN(n7578) );
  INV_X1 U8616 ( .A(P2_ADDR_REG_9__SCAN_IN), .ZN(n7259) );
  NOR2_X1 U8617 ( .A1(n7260), .A2(n7259), .ZN(n7261) );
  AOI211_X1 U8618 ( .C1(n8920), .C2(n10896), .A(n7578), .B(n7261), .ZN(n7262)
         );
  OAI21_X1 U8619 ( .B1(n7263), .B2(n10910), .A(n7262), .ZN(n7264) );
  AOI21_X1 U8620 ( .B1(n10905), .B2(n7265), .A(n7264), .ZN(n7266) );
  OAI21_X1 U8621 ( .B1(n7267), .B2(n10772), .A(n7266), .ZN(P2_U3191) );
  NAND2_X1 U8622 ( .A1(n7394), .A2(n11019), .ZN(n9546) );
  XNOR2_X1 U8623 ( .A(n7393), .B(n7395), .ZN(n11040) );
  INV_X1 U8624 ( .A(n10328), .ZN(n7564) );
  OAI22_X1 U8625 ( .A1(n10387), .A2(n7394), .B1(n11036), .B2(n10213), .ZN(
        n7279) );
  NAND2_X1 U8626 ( .A1(n7271), .A2(n7004), .ZN(n7272) );
  NAND2_X1 U8627 ( .A1(n7272), .A2(n5131), .ZN(n7273) );
  NOR2_X1 U8628 ( .A1(n7386), .A2(n7273), .ZN(n11037) );
  INV_X1 U8629 ( .A(n11037), .ZN(n7277) );
  INV_X1 U8630 ( .A(n7274), .ZN(n7275) );
  AOI22_X1 U8631 ( .A1(n7171), .A2(P1_REG2_REG_4__SCAN_IN), .B1(n7275), .B2(
        n11123), .ZN(n7276) );
  OAI21_X1 U8632 ( .B1(n7277), .B2(n10333), .A(n7276), .ZN(n7278) );
  AOI211_X1 U8633 ( .C1(n7564), .C2(n11064), .A(n7279), .B(n7278), .ZN(n7282)
         );
  NAND2_X1 U8634 ( .A1(n7280), .A2(n9543), .ZN(n7383) );
  XNOR2_X1 U8635 ( .A(n7393), .B(n7383), .ZN(n11042) );
  NAND2_X1 U8636 ( .A1(n11042), .A2(n10335), .ZN(n7281) );
  OAI211_X1 U8637 ( .C1(n11040), .C2(n10391), .A(n7282), .B(n7281), .ZN(
        P1_U3289) );
  OR2_X1 U8638 ( .A1(n7283), .A2(n6959), .ZN(n7287) );
  OR2_X1 U8639 ( .A1(n7322), .A2(n10628), .ZN(n7286) );
  OR2_X1 U8640 ( .A1(n5138), .A2(n7284), .ZN(n7285) );
  AOI22_X1 U8641 ( .A1(n11048), .A2(n8349), .B1(n8264), .B2(n11064), .ZN(n7317) );
  NAND2_X1 U8642 ( .A1(n7289), .A2(n7288), .ZN(n7290) );
  INV_X1 U8643 ( .A(n7296), .ZN(n7294) );
  NAND2_X1 U8644 ( .A1(n11064), .A2(n8387), .ZN(n7291) );
  OAI21_X1 U8645 ( .B1(n7385), .B2(n8330), .A(n7291), .ZN(n7292) );
  XNOR2_X1 U8646 ( .A(n7292), .B(n8346), .ZN(n7295) );
  INV_X1 U8647 ( .A(n7295), .ZN(n7293) );
  NAND2_X1 U8648 ( .A1(n7294), .A2(n7293), .ZN(n7319) );
  NAND2_X1 U8649 ( .A1(n7296), .A2(n7295), .ZN(n7318) );
  NAND2_X1 U8650 ( .A1(n7319), .A2(n7318), .ZN(n7297) );
  XOR2_X1 U8651 ( .A(n7317), .B(n7297), .Z(n7298) );
  NAND2_X1 U8652 ( .A1(n7298), .A2(n9376), .ZN(n7309) );
  NAND2_X1 U8653 ( .A1(P1_U3086), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n10637) );
  INV_X1 U8654 ( .A(n10637), .ZN(n7307) );
  NAND2_X1 U8655 ( .A1(n8357), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7305) );
  INV_X1 U8656 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7299) );
  OR2_X1 U8657 ( .A1(n6966), .A2(n7299), .ZN(n7304) );
  AND2_X1 U8658 ( .A1(n7300), .A2(n7336), .ZN(n7301) );
  OR2_X1 U8659 ( .A1(n7301), .A2(n7338), .ZN(n11073) );
  OR2_X1 U8660 ( .A1(n8382), .A2(n11073), .ZN(n7303) );
  OR2_X1 U8661 ( .A1(n5143), .A2(n6851), .ZN(n7302) );
  OAI22_X1 U8662 ( .A1(n9369), .A2(n11046), .B1(n11085), .B2(n9391), .ZN(n7306) );
  AOI211_X1 U8663 ( .C1(n11048), .C2(n9399), .A(n7307), .B(n7306), .ZN(n7308)
         );
  OAI211_X1 U8664 ( .C1(n9397), .C2(n7387), .A(n7309), .B(n7308), .ZN(P1_U3227) );
  OAI22_X1 U8665 ( .A1(n9141), .A2(n7311), .B1(n7310), .B2(n9142), .ZN(n7314)
         );
  MUX2_X1 U8666 ( .A(P2_REG2_REG_4__SCAN_IN), .B(n7312), .S(n9145), .Z(n7313)
         );
  AOI211_X1 U8667 ( .C1(n9148), .C2(n7315), .A(n7314), .B(n7313), .ZN(n7316)
         );
  INV_X1 U8668 ( .A(n7316), .ZN(P2_U3229) );
  NAND2_X1 U8669 ( .A1(n7318), .A2(n7317), .ZN(n7320) );
  OR2_X1 U8670 ( .A1(n7321), .A2(n6959), .ZN(n7324) );
  AOI22_X1 U8671 ( .A1(n8215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n8214), .B2(
        n10648), .ZN(n7323) );
  NAND2_X1 U8672 ( .A1(n7324), .A2(n7323), .ZN(n11075) );
  NAND2_X1 U8673 ( .A1(n11075), .A2(n8388), .ZN(n7327) );
  OR2_X1 U8674 ( .A1(n11085), .A2(n8390), .ZN(n7326) );
  NAND2_X1 U8675 ( .A1(n7327), .A2(n7326), .ZN(n7328) );
  XNOR2_X1 U8676 ( .A(n7328), .B(n8314), .ZN(n7334) );
  INV_X1 U8677 ( .A(n7334), .ZN(n7332) );
  NAND2_X1 U8678 ( .A1(n11075), .A2(n8349), .ZN(n7330) );
  OR2_X1 U8679 ( .A1(n11085), .A2(n5144), .ZN(n7329) );
  AND2_X1 U8680 ( .A1(n7330), .A2(n7329), .ZN(n7333) );
  INV_X1 U8681 ( .A(n7333), .ZN(n7331) );
  NAND2_X1 U8682 ( .A1(n7332), .A2(n7331), .ZN(n7459) );
  NAND2_X1 U8683 ( .A1(n7334), .A2(n7333), .ZN(n7458) );
  NAND2_X1 U8684 ( .A1(n7335), .A2(n9376), .ZN(n7346) );
  NOR2_X1 U8685 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7336), .ZN(n10650) );
  NAND2_X1 U8686 ( .A1(n8357), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7343) );
  INV_X1 U8687 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7337) );
  OR2_X1 U8688 ( .A1(n6966), .A2(n7337), .ZN(n7342) );
  OR2_X1 U8689 ( .A1(n7338), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7339) );
  NAND2_X1 U8690 ( .A1(n7412), .A2(n7339), .ZN(n7472) );
  OR2_X1 U8691 ( .A1(n8382), .A2(n7472), .ZN(n7341) );
  INV_X1 U8692 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7409) );
  OR2_X1 U8693 ( .A1(n5143), .A2(n7409), .ZN(n7340) );
  OAI22_X1 U8694 ( .A1(n9369), .A2(n11035), .B1(n11110), .B2(n9391), .ZN(n7344) );
  AOI211_X1 U8695 ( .C1(n11075), .C2(n9399), .A(n10650), .B(n7344), .ZN(n7345)
         );
  OAI211_X1 U8696 ( .C1(n9397), .C2(n11073), .A(n7346), .B(n7345), .ZN(
        P1_U3239) );
  XNOR2_X1 U8697 ( .A(n7347), .B(n8480), .ZN(n7348) );
  OAI222_X1 U8698 ( .A1(n9121), .A2(n7500), .B1(n9119), .B2(n7349), .C1(n9116), 
        .C2(n7348), .ZN(n7515) );
  XOR2_X1 U8699 ( .A(n7350), .B(n8480), .Z(n7521) );
  OAI22_X1 U8700 ( .A1(n7521), .A2(n9188), .B1(n7351), .B2(n9173), .ZN(n7352)
         );
  NOR2_X1 U8701 ( .A1(n7515), .A2(n7352), .ZN(n11056) );
  OR2_X1 U8702 ( .A1(n9206), .A2(n7078), .ZN(n7353) );
  OAI21_X1 U8703 ( .B1(n11056), .B2(n9210), .A(n7353), .ZN(P2_U3465) );
  NOR2_X1 U8704 ( .A1(n10122), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n7354) );
  AOI21_X1 U8705 ( .B1(P1_REG2_REG_12__SCAN_IN), .B2(n10122), .A(n7354), .ZN(
        n7359) );
  AOI22_X1 U8706 ( .A1(n7525), .A2(P1_REG2_REG_10__SCAN_IN), .B1(n6560), .B2(
        n9683), .ZN(n9676) );
  OAI21_X1 U8707 ( .B1(P1_REG2_REG_9__SCAN_IN), .B2(n7528), .A(n7355), .ZN(
        n9675) );
  INV_X1 U8708 ( .A(n9675), .ZN(n7356) );
  NAND2_X1 U8709 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n10690), .ZN(n7357) );
  OAI21_X1 U8710 ( .B1(P1_REG2_REG_11__SCAN_IN), .B2(n10690), .A(n7357), .ZN(
        n10686) );
  OAI21_X1 U8711 ( .B1(n7359), .B2(n7358), .A(n10121), .ZN(n7370) );
  INV_X1 U8712 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n11166) );
  AOI22_X1 U8713 ( .A1(n10122), .A2(P1_REG1_REG_12__SCAN_IN), .B1(n11166), 
        .B2(n7368), .ZN(n7364) );
  INV_X1 U8714 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n11143) );
  INV_X1 U8715 ( .A(n7360), .ZN(n7361) );
  AOI21_X1 U8716 ( .B1(n11143), .B2(n7362), .A(n7361), .ZN(n9678) );
  INV_X1 U8717 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n11154) );
  AOI22_X1 U8718 ( .A1(n7525), .A2(P1_REG1_REG_10__SCAN_IN), .B1(n11154), .B2(
        n9683), .ZN(n9679) );
  INV_X1 U8719 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n7557) );
  MUX2_X1 U8720 ( .A(n7557), .B(P1_REG1_REG_11__SCAN_IN), .S(n10690), .Z(
        n10683) );
  NOR2_X1 U8721 ( .A1(n10684), .A2(n10683), .ZN(n10682) );
  NAND2_X1 U8722 ( .A1(n7364), .A2(n7363), .ZN(n10112) );
  OAI21_X1 U8723 ( .B1(n7364), .B2(n7363), .A(n10112), .ZN(n7365) );
  NAND2_X1 U8724 ( .A1(n7365), .A2(n10954), .ZN(n7367) );
  AND2_X1 U8725 ( .A1(P1_U3086), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7937) );
  AOI21_X1 U8726 ( .B1(n10942), .B2(P1_ADDR_REG_12__SCAN_IN), .A(n7937), .ZN(
        n7366) );
  OAI211_X1 U8727 ( .C1(n10949), .C2(n7368), .A(n7367), .B(n7366), .ZN(n7369)
         );
  AOI21_X1 U8728 ( .B1(n7370), .B2(n9685), .A(n7369), .ZN(n7371) );
  INV_X1 U8729 ( .A(n7371), .ZN(P1_U3255) );
  INV_X1 U8730 ( .A(P2_REG2_REG_31__SCAN_IN), .ZN(n7378) );
  NAND2_X1 U8731 ( .A1(n7372), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n7376) );
  INV_X1 U8732 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n7373) );
  OR2_X1 U8733 ( .A1(n7374), .A2(n7373), .ZN(n7375) );
  OAI211_X1 U8734 ( .C1(n7378), .C2(n7377), .A(n7376), .B(n7375), .ZN(n7379)
         );
  INV_X1 U8735 ( .A(n7379), .ZN(n7380) );
  NAND2_X1 U8736 ( .A1(n8913), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n7382) );
  OAI21_X1 U8737 ( .B1(n8977), .B2(n8913), .A(n7382), .ZN(P2_U3522) );
  NAND2_X1 U8738 ( .A1(n7383), .A2(n7393), .ZN(n7384) );
  NAND2_X1 U8739 ( .A1(n7384), .A2(n9544), .ZN(n7404) );
  NAND2_X1 U8740 ( .A1(n11035), .A2(n11048), .ZN(n9415) );
  NAND2_X1 U8741 ( .A1(n7385), .A2(n11064), .ZN(n9552) );
  NAND2_X1 U8742 ( .A1(n9415), .A2(n9552), .ZN(n9482) );
  INV_X1 U8743 ( .A(n9482), .ZN(n9557) );
  XNOR2_X1 U8744 ( .A(n7404), .B(n9557), .ZN(n11053) );
  OAI211_X1 U8745 ( .C1(n7386), .C2(n7385), .A(n5131), .B(n11058), .ZN(n11049)
         );
  OAI22_X1 U8746 ( .A1(n10367), .A2(n7388), .B1(n7387), .B2(n10968), .ZN(n7389) );
  AOI21_X1 U8747 ( .B1(n11124), .B2(n11048), .A(n7389), .ZN(n7392) );
  OAI22_X1 U8748 ( .A1(n11046), .A2(n10213), .B1(n10328), .B2(n11085), .ZN(
        n7390) );
  INV_X1 U8749 ( .A(n7390), .ZN(n7391) );
  OAI211_X1 U8750 ( .C1(n11049), .C2(n10333), .A(n7392), .B(n7391), .ZN(n7397)
         );
  INV_X1 U8751 ( .A(n7393), .ZN(n9481) );
  XNOR2_X1 U8752 ( .A(n7399), .B(n9482), .ZN(n11051) );
  NOR2_X1 U8753 ( .A1(n11051), .A2(n10391), .ZN(n7396) );
  AOI211_X1 U8754 ( .C1(n11053), .C2(n10335), .A(n7397), .B(n7396), .ZN(n7398)
         );
  INV_X1 U8755 ( .A(n7398), .ZN(P1_U3288) );
  AND2_X1 U8756 ( .A1(n11075), .A2(n11085), .ZN(n9483) );
  INV_X1 U8757 ( .A(n9483), .ZN(n9559) );
  INV_X1 U8758 ( .A(n11075), .ZN(n11061) );
  INV_X1 U8759 ( .A(n11085), .ZN(n9674) );
  AOI22_X1 U8760 ( .A1(n8215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n8214), .B2(
        n7401), .ZN(n7402) );
  XNOR2_X1 U8761 ( .A(n7552), .B(n9562), .ZN(n11092) );
  AND2_X1 U8762 ( .A1(n7546), .A2(n9561), .ZN(n7405) );
  NAND2_X1 U8763 ( .A1(n7405), .A2(n9553), .ZN(n11103) );
  OAI21_X1 U8764 ( .B1(n9553), .B2(n7405), .A(n11103), .ZN(n7406) );
  NAND2_X1 U8765 ( .A1(n7406), .A2(n11181), .ZN(n11089) );
  INV_X1 U8766 ( .A(n11089), .ZN(n7424) );
  NAND2_X1 U8767 ( .A1(n11059), .A2(n11088), .ZN(n7407) );
  NAND2_X1 U8768 ( .A1(n7407), .A2(n5131), .ZN(n7408) );
  NOR2_X1 U8769 ( .A1(n11116), .A2(n7408), .ZN(n11086) );
  NAND2_X1 U8770 ( .A1(n11086), .A2(n11128), .ZN(n7422) );
  OAI22_X1 U8771 ( .A1(n10367), .A2(n7409), .B1(n7472), .B2(n10968), .ZN(n7410) );
  AOI21_X1 U8772 ( .B1(n11124), .B2(n11088), .A(n7410), .ZN(n7421) );
  NAND2_X1 U8773 ( .A1(n8377), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n7418) );
  INV_X1 U8774 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n7411) );
  OR2_X1 U8775 ( .A1(n6968), .A2(n7411), .ZN(n7417) );
  NAND2_X1 U8776 ( .A1(n7412), .A2(n7676), .ZN(n7413) );
  NAND2_X1 U8777 ( .A1(n7532), .A2(n7413), .ZN(n11121) );
  OR2_X1 U8778 ( .A1(n8382), .A2(n11121), .ZN(n7416) );
  INV_X1 U8779 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n7414) );
  OR2_X1 U8780 ( .A1(n5143), .A2(n7414), .ZN(n7415) );
  OAI22_X1 U8781 ( .A1(n11085), .A2(n10213), .B1(n10328), .B2(n11084), .ZN(
        n7419) );
  INV_X1 U8782 ( .A(n7419), .ZN(n7420) );
  NAND3_X1 U8783 ( .A1(n7422), .A2(n7421), .A3(n7420), .ZN(n7423) );
  AOI21_X1 U8784 ( .B1(n7424), .B2(n10358), .A(n7423), .ZN(n7425) );
  OAI21_X1 U8785 ( .B1(n11092), .B2(n10391), .A(n7425), .ZN(P1_U3286) );
  NAND2_X1 U8786 ( .A1(n7426), .A2(n8840), .ZN(n7427) );
  XNOR2_X1 U8787 ( .A(n8162), .B(n8440), .ZN(n7501) );
  XNOR2_X1 U8788 ( .A(n7501), .B(n8839), .ZN(n7429) );
  OAI21_X1 U8789 ( .B1(n7430), .B2(n7429), .A(n7503), .ZN(n7438) );
  NOR2_X1 U8790 ( .A1(n8519), .A2(n8823), .ZN(n7437) );
  INV_X1 U8791 ( .A(n8160), .ZN(n7431) );
  NAND2_X1 U8792 ( .A1(n8819), .A2(n7431), .ZN(n7435) );
  INV_X1 U8793 ( .A(n7432), .ZN(n7433) );
  AOI21_X1 U8794 ( .B1(n8840), .B2(n8800), .A(n7433), .ZN(n7434) );
  OAI211_X1 U8795 ( .C1(n7570), .C2(n8803), .A(n7435), .B(n7434), .ZN(n7436)
         );
  AOI211_X1 U8796 ( .C1(n7438), .C2(n8810), .A(n7437), .B(n7436), .ZN(n7439)
         );
  INV_X1 U8797 ( .A(n7439), .ZN(P2_U3153) );
  NAND2_X1 U8798 ( .A1(n7133), .A2(n8552), .ZN(n7440) );
  AND2_X1 U8799 ( .A1(n8553), .A2(n8559), .ZN(n8476) );
  XNOR2_X1 U8800 ( .A(n7440), .B(n8476), .ZN(n7498) );
  NOR2_X1 U8801 ( .A1(n7493), .A2(n9173), .ZN(n7447) );
  INV_X1 U8802 ( .A(n8476), .ZN(n7442) );
  XNOR2_X1 U8803 ( .A(n7441), .B(n7442), .ZN(n7446) );
  INV_X1 U8804 ( .A(n7734), .ZN(n7443) );
  NAND2_X1 U8805 ( .A1(n7498), .A2(n7443), .ZN(n7445) );
  AOI22_X1 U8806 ( .A1(n9136), .A2(n8842), .B1(n8840), .B2(n9133), .ZN(n7444)
         );
  OAI211_X1 U8807 ( .C1(n9116), .C2(n7446), .A(n7445), .B(n7444), .ZN(n7494)
         );
  AOI211_X1 U8808 ( .C1(n7498), .C2(n7448), .A(n7447), .B(n7494), .ZN(n11045)
         );
  OR2_X1 U8809 ( .A1(n11045), .A2(n9210), .ZN(n7449) );
  OAI21_X1 U8810 ( .B1(n9206), .B2(n7450), .A(n7449), .ZN(P2_U3464) );
  INV_X1 U8811 ( .A(n8132), .ZN(n7456) );
  INV_X1 U8812 ( .A(n10897), .ZN(n8941) );
  OAI222_X1 U8813 ( .A1(n9267), .A2(n7451), .B1(n9262), .B2(n7456), .C1(n8941), 
        .C2(P2_U3151), .ZN(P2_U3278) );
  OAI21_X1 U8814 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(P1_IR_REG_15__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n7452) );
  NAND2_X1 U8815 ( .A1(n7453), .A2(n7452), .ZN(n7455) );
  INV_X1 U8816 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n7454) );
  XNOR2_X1 U8817 ( .A(n7455), .B(n7454), .ZN(n10154) );
  INV_X1 U8818 ( .A(n10154), .ZN(n10145) );
  OAI222_X1 U8819 ( .A1(n5141), .A2(n7457), .B1(P1_U3086), .B2(n10145), .C1(
        n7456), .C2(n10517), .ZN(P1_U3338) );
  NAND2_X1 U8820 ( .A1(n11088), .A2(n8388), .ZN(n7462) );
  OR2_X1 U8821 ( .A1(n11110), .A2(n8390), .ZN(n7461) );
  NAND2_X1 U8822 ( .A1(n7462), .A2(n7461), .ZN(n7463) );
  XNOR2_X1 U8823 ( .A(n7463), .B(n8346), .ZN(n7679) );
  NAND2_X1 U8824 ( .A1(n11088), .A2(n8349), .ZN(n7465) );
  OR2_X1 U8825 ( .A1(n11110), .A2(n5144), .ZN(n7464) );
  NAND2_X1 U8826 ( .A1(n7465), .A2(n7464), .ZN(n7680) );
  XNOR2_X1 U8827 ( .A(n7679), .B(n7680), .ZN(n7466) );
  XNOR2_X1 U8828 ( .A(n7681), .B(n7466), .ZN(n7467) );
  NAND2_X1 U8829 ( .A1(n7467), .A2(n9376), .ZN(n7471) );
  NAND2_X1 U8830 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10666) );
  INV_X1 U8831 ( .A(n10666), .ZN(n7469) );
  OAI22_X1 U8832 ( .A1(n9369), .A2(n11085), .B1(n11084), .B2(n9391), .ZN(n7468) );
  AOI211_X1 U8833 ( .C1(n11088), .C2(n9399), .A(n7469), .B(n7468), .ZN(n7470)
         );
  OAI211_X1 U8834 ( .C1(n9397), .C2(n7472), .A(n7471), .B(n7470), .ZN(P1_U3213) );
  OR2_X1 U8835 ( .A1(n7590), .A2(n8560), .ZN(n7617) );
  NAND2_X1 U8836 ( .A1(n7590), .A2(n8560), .ZN(n7473) );
  NAND2_X1 U8837 ( .A1(n7617), .A2(n7473), .ZN(n7474) );
  NAND2_X1 U8838 ( .A1(n7474), .A2(n9130), .ZN(n7476) );
  AOI22_X1 U8839 ( .A1(n9136), .A2(n8840), .B1(n8838), .B2(n9133), .ZN(n7475)
         );
  NAND2_X1 U8840 ( .A1(n7476), .A2(n7475), .ZN(n8158) );
  NAND2_X1 U8841 ( .A1(n7478), .A2(n5397), .ZN(n8159) );
  AND3_X1 U8842 ( .A1(n7477), .A2(n9204), .A3(n8159), .ZN(n7479) );
  NOR2_X1 U8843 ( .A1(n8158), .A2(n7479), .ZN(n7486) );
  INV_X1 U8844 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n7480) );
  OAI22_X1 U8845 ( .A1(n8519), .A2(n9250), .B1(n11186), .B2(n7480), .ZN(n7481)
         );
  INV_X1 U8846 ( .A(n7481), .ZN(n7482) );
  OAI21_X1 U8847 ( .B1(n7486), .B2(n6448), .A(n7482), .ZN(P2_U3411) );
  INV_X1 U8848 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n7483) );
  OAI22_X1 U8849 ( .A1(n8519), .A2(n9209), .B1(n9206), .B2(n7483), .ZN(n7484)
         );
  INV_X1 U8850 ( .A(n7484), .ZN(n7485) );
  OAI21_X1 U8851 ( .B1(n7486), .B2(n9210), .A(n7485), .ZN(P2_U3466) );
  INV_X1 U8852 ( .A(n8203), .ZN(n7522) );
  NAND2_X1 U8853 ( .A1(n7487), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7488) );
  XNOR2_X1 U8854 ( .A(n7488), .B(P1_IR_REG_18__SCAN_IN), .ZN(n10730) );
  AOI22_X1 U8855 ( .A1(n10730), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n7489), .ZN(n7490) );
  OAI21_X1 U8856 ( .B1(n7522), .B2(n10517), .A(n7490), .ZN(P1_U3337) );
  NAND2_X1 U8857 ( .A1(n9145), .A2(n7491), .ZN(n8988) );
  INV_X1 U8858 ( .A(n8988), .ZN(n7497) );
  OAI22_X1 U8859 ( .A1(n9141), .A2(n7493), .B1(n7492), .B2(n9142), .ZN(n7496)
         );
  MUX2_X1 U8860 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7494), .S(n9145), .Z(n7495)
         );
  AOI211_X1 U8861 ( .C1(n7498), .C2(n7497), .A(n7496), .B(n7495), .ZN(n7499)
         );
  INV_X1 U8862 ( .A(n7499), .ZN(P2_U3228) );
  INV_X1 U8863 ( .A(n7628), .ZN(n7514) );
  INV_X1 U8864 ( .A(n7503), .ZN(n7502) );
  XNOR2_X1 U8865 ( .A(n7628), .B(n8440), .ZN(n7571) );
  XNOR2_X1 U8866 ( .A(n7571), .B(n8838), .ZN(n7504) );
  NOR3_X1 U8867 ( .A1(n7502), .A2(n5243), .A3(n7504), .ZN(n7507) );
  NAND2_X1 U8868 ( .A1(n7505), .A2(n7504), .ZN(n7573) );
  INV_X1 U8869 ( .A(n7573), .ZN(n7506) );
  OAI21_X1 U8870 ( .B1(n7507), .B2(n7506), .A(n8810), .ZN(n7513) );
  INV_X1 U8871 ( .A(n7508), .ZN(n7627) );
  AOI22_X1 U8872 ( .A1(n8839), .A2(n8800), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3151), .ZN(n7509) );
  OAI21_X1 U8873 ( .B1(n7510), .B2(n8803), .A(n7509), .ZN(n7511) );
  AOI21_X1 U8874 ( .B1(n7627), .B2(n8819), .A(n7511), .ZN(n7512) );
  OAI211_X1 U8875 ( .C1(n7514), .C2(n8823), .A(n7513), .B(n7512), .ZN(P2_U3161) );
  INV_X1 U8876 ( .A(n7515), .ZN(n7516) );
  MUX2_X1 U8877 ( .A(n5357), .B(n7516), .S(n9145), .Z(n7520) );
  AOI22_X1 U8878 ( .A1(n9111), .A2(n7518), .B1(n9125), .B2(n7517), .ZN(n7519)
         );
  OAI211_X1 U8879 ( .C1(n9114), .C2(n7521), .A(n7520), .B(n7519), .ZN(P2_U3227) );
  INV_X1 U8880 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n7523) );
  INV_X1 U8881 ( .A(n8948), .ZN(n8965) );
  OAI222_X1 U8882 ( .A1(n9267), .A2(n7523), .B1(P2_U3151), .B2(n8965), .C1(
        n7522), .C2(n9262), .ZN(P2_U3277) );
  OR2_X1 U8883 ( .A1(n7524), .A2(n6959), .ZN(n7527) );
  AOI22_X1 U8884 ( .A1(n8215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n8214), .B2(
        n7525), .ZN(n7526) );
  NAND2_X1 U8885 ( .A1(n11148), .A2(n7884), .ZN(n9533) );
  NAND2_X1 U8886 ( .A1(n6541), .A2(n8029), .ZN(n7530) );
  AOI22_X1 U8887 ( .A1(n8215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n8214), .B2(
        n7528), .ZN(n7529) );
  NAND2_X1 U8888 ( .A1(n8377), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7538) );
  OR2_X1 U8889 ( .A1(n6968), .A2(n11143), .ZN(n7537) );
  AND2_X1 U8890 ( .A1(n7532), .A2(n7531), .ZN(n7534) );
  OR2_X1 U8891 ( .A1(n7534), .A2(n7533), .ZN(n7779) );
  OR2_X1 U8892 ( .A1(n8382), .A2(n7779), .ZN(n7536) );
  INV_X1 U8893 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n7606) );
  OR2_X1 U8894 ( .A1(n5143), .A2(n7606), .ZN(n7535) );
  NAND2_X1 U8895 ( .A1(n7539), .A2(n8029), .ZN(n7541) );
  AOI22_X1 U8896 ( .A1(n8215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n8214), .B2(
        n10677), .ZN(n7540) );
  NAND2_X1 U8897 ( .A1(n7541), .A2(n7540), .ZN(n11125) );
  OR2_X1 U8898 ( .A1(n11125), .A2(n11084), .ZN(n9535) );
  NAND2_X1 U8899 ( .A1(n5202), .A2(n7544), .ZN(n9488) );
  INV_X1 U8900 ( .A(n9488), .ZN(n7545) );
  NAND2_X1 U8901 ( .A1(n11125), .A2(n11084), .ZN(n9532) );
  NAND2_X1 U8902 ( .A1(n11137), .A2(n11108), .ZN(n9526) );
  AND2_X1 U8903 ( .A1(n7547), .A2(n9526), .ZN(n9418) );
  NAND2_X1 U8904 ( .A1(n7548), .A2(n9418), .ZN(n7549) );
  NAND2_X1 U8905 ( .A1(n7549), .A2(n7553), .ZN(n7650) );
  OAI21_X1 U8906 ( .B1(n7553), .B2(n7549), .A(n7650), .ZN(n7551) );
  NOR2_X1 U8907 ( .A1(n11108), .A2(n11109), .ZN(n7550) );
  AOI21_X1 U8908 ( .B1(n7551), .B2(n11181), .A(n7550), .ZN(n11151) );
  INV_X1 U8909 ( .A(n11110), .ZN(n11065) );
  OAI22_X1 U8910 ( .A1(n7552), .A2(n9553), .B1(n11088), .B2(n11065), .ZN(
        n11099) );
  INV_X1 U8911 ( .A(n11101), .ZN(n11098) );
  INV_X1 U8912 ( .A(n11125), .ZN(n11117) );
  AOI22_X2 U8913 ( .A1(n11099), .A2(n11098), .B1(n11117), .B2(n11084), .ZN(
        n7610) );
  INV_X1 U8914 ( .A(n11108), .ZN(n9673) );
  XNOR2_X1 U8915 ( .A(n7633), .B(n9489), .ZN(n11153) );
  NAND2_X1 U8916 ( .A1(n11153), .A2(n11129), .ZN(n7569) );
  INV_X1 U8917 ( .A(n11137), .ZN(n7554) );
  INV_X1 U8918 ( .A(n7555), .ZN(n7556) );
  INV_X1 U8919 ( .A(n11148), .ZN(n7632) );
  OAI211_X1 U8920 ( .C1(n7556), .C2(n7632), .A(n5131), .B(n7638), .ZN(n11149)
         );
  INV_X1 U8921 ( .A(n11149), .ZN(n7567) );
  NAND2_X1 U8922 ( .A1(n8377), .A2(P1_REG0_REG_11__SCAN_IN), .ZN(n7562) );
  OR2_X1 U8923 ( .A1(n6968), .A2(n7557), .ZN(n7561) );
  XNOR2_X1 U8924 ( .A(n7642), .B(P1_REG3_REG_11__SCAN_IN), .ZN(n7883) );
  OR2_X1 U8925 ( .A1(n8382), .A2(n7883), .ZN(n7560) );
  INV_X1 U8926 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7639) );
  OR2_X1 U8927 ( .A1(n5143), .A2(n7639), .ZN(n7559) );
  INV_X1 U8928 ( .A(n7872), .ZN(n11146) );
  OAI22_X1 U8929 ( .A1(n10358), .A2(n6560), .B1(n7839), .B2(n10968), .ZN(n7563) );
  AOI21_X1 U8930 ( .B1(n7564), .B2(n11146), .A(n7563), .ZN(n7565) );
  OAI21_X1 U8931 ( .B1(n7632), .B2(n10387), .A(n7565), .ZN(n7566) );
  AOI21_X1 U8932 ( .B1(n7567), .B2(n11128), .A(n7566), .ZN(n7568) );
  OAI211_X1 U8933 ( .C1(n7171), .C2(n11151), .A(n7569), .B(n7568), .ZN(
        P1_U3283) );
  INV_X1 U8934 ( .A(n7664), .ZN(n7584) );
  NAND2_X1 U8935 ( .A1(n7571), .A2(n7570), .ZN(n7572) );
  XNOR2_X1 U8936 ( .A(n7664), .B(n8424), .ZN(n7703) );
  XNOR2_X1 U8937 ( .A(n7703), .B(n8837), .ZN(n7575) );
  AOI21_X1 U8938 ( .B1(n7574), .B2(n7575), .A(n8808), .ZN(n7577) );
  INV_X1 U8939 ( .A(n7575), .ZN(n7576) );
  NAND2_X1 U8940 ( .A1(n7577), .A2(n7705), .ZN(n7583) );
  INV_X1 U8941 ( .A(n7597), .ZN(n7581) );
  AOI21_X1 U8942 ( .B1(n8838), .B2(n8800), .A(n7578), .ZN(n7579) );
  OAI21_X1 U8943 ( .B1(n7849), .B2(n8803), .A(n7579), .ZN(n7580) );
  AOI21_X1 U8944 ( .B1(n7581), .B2(n8819), .A(n7580), .ZN(n7582) );
  OAI211_X1 U8945 ( .C1(n7584), .C2(n8823), .A(n7583), .B(n7582), .ZN(P2_U3171) );
  OR2_X1 U8946 ( .A1(n7590), .A2(n7585), .ZN(n7588) );
  AND2_X1 U8947 ( .A1(n7588), .A2(n7587), .ZN(n7595) );
  OR2_X1 U8948 ( .A1(n7590), .A2(n7589), .ZN(n7592) );
  AND2_X1 U8949 ( .A1(n7592), .A2(n7591), .ZN(n7619) );
  NAND3_X1 U8950 ( .A1(n7619), .A2(n6031), .A3(n7593), .ZN(n7594) );
  NAND2_X1 U8951 ( .A1(n7595), .A2(n7594), .ZN(n7596) );
  AOI222_X1 U8952 ( .A1(n9130), .A2(n7596), .B1(n8836), .B2(n9133), .C1(n8838), 
        .C2(n9136), .ZN(n7660) );
  OAI22_X1 U8953 ( .A1(n9145), .A2(n8921), .B1(n7597), .B2(n9142), .ZN(n7598)
         );
  AOI21_X1 U8954 ( .B1(n7664), .B2(n9111), .A(n7598), .ZN(n7602) );
  NAND2_X1 U8955 ( .A1(n7600), .A2(n8514), .ZN(n7658) );
  NAND3_X1 U8956 ( .A1(n7599), .A2(n9148), .A3(n7658), .ZN(n7601) );
  OAI211_X1 U8957 ( .C1(n7660), .C2(n9150), .A(n7602), .B(n7601), .ZN(P2_U3224) );
  NAND3_X1 U8958 ( .A1(n11103), .A2(n11101), .A3(n11102), .ZN(n11100) );
  NAND2_X1 U8959 ( .A1(n11100), .A2(n9535), .ZN(n7603) );
  XOR2_X1 U8960 ( .A(n9569), .B(n7603), .Z(n11142) );
  XNOR2_X1 U8961 ( .A(n11113), .B(n11137), .ZN(n7605) );
  NOR2_X1 U8962 ( .A1(n7884), .A2(n11107), .ZN(n7604) );
  AOI21_X1 U8963 ( .B1(n7605), .B2(n5131), .A(n7604), .ZN(n11139) );
  INV_X1 U8964 ( .A(n11084), .ZN(n11136) );
  OAI22_X1 U8965 ( .A1(n10367), .A2(n7606), .B1(n7779), .B2(n10968), .ZN(n7607) );
  AOI21_X1 U8966 ( .B1(n10326), .B2(n11136), .A(n7607), .ZN(n7609) );
  NAND2_X1 U8967 ( .A1(n11137), .A2(n11124), .ZN(n7608) );
  OAI211_X1 U8968 ( .C1(n11139), .C2(n10333), .A(n7609), .B(n7608), .ZN(n7612)
         );
  XOR2_X1 U8969 ( .A(n9569), .B(n7610), .Z(n11140) );
  NOR2_X1 U8970 ( .A1(n11140), .A2(n10391), .ZN(n7611) );
  AOI211_X1 U8971 ( .C1(n10335), .C2(n11142), .A(n7612), .B(n7611), .ZN(n7613)
         );
  INV_X1 U8972 ( .A(n7613), .ZN(P1_U3284) );
  NAND2_X1 U8973 ( .A1(n7477), .A2(n7614), .ZN(n7615) );
  XNOR2_X1 U8974 ( .A(n7615), .B(n6030), .ZN(n7631) );
  NOR2_X1 U8975 ( .A1(n7631), .A2(n9188), .ZN(n7623) );
  NAND3_X1 U8976 ( .A1(n7617), .A2(n6030), .A3(n7616), .ZN(n7618) );
  NAND2_X1 U8977 ( .A1(n7619), .A2(n7618), .ZN(n7620) );
  NAND2_X1 U8978 ( .A1(n7620), .A2(n9130), .ZN(n7622) );
  AOI22_X1 U8979 ( .A1(n9136), .A2(n8839), .B1(n8837), .B2(n9133), .ZN(n7621)
         );
  NAND2_X1 U8980 ( .A1(n7622), .A2(n7621), .ZN(n7625) );
  AOI211_X1 U8981 ( .C1(n9180), .C2(n7628), .A(n7623), .B(n7625), .ZN(n11135)
         );
  NAND2_X1 U8982 ( .A1(n9210), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n7624) );
  OAI21_X1 U8983 ( .B1(n11135), .B2(n9210), .A(n7624), .ZN(P2_U3467) );
  MUX2_X1 U8984 ( .A(n7625), .B(P2_REG2_REG_8__SCAN_IN), .S(n9150), .Z(n7626)
         );
  INV_X1 U8985 ( .A(n7626), .ZN(n7630) );
  AOI22_X1 U8986 ( .A1(n7628), .A2(n9111), .B1(n9125), .B2(n7627), .ZN(n7629)
         );
  OAI211_X1 U8987 ( .C1(n7631), .C2(n9114), .A(n7630), .B(n7629), .ZN(P2_U3225) );
  NAND2_X1 U8988 ( .A1(n7634), .A2(n8029), .ZN(n7636) );
  AOI22_X1 U8989 ( .A1(n8215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n8214), .B2(
        n10690), .ZN(n7635) );
  OR2_X1 U8990 ( .A1(n7874), .A2(n7872), .ZN(n9522) );
  NAND2_X1 U8991 ( .A1(n7874), .A2(n7872), .ZN(n9517) );
  NAND2_X1 U8992 ( .A1(n9522), .A2(n9517), .ZN(n9492) );
  XNOR2_X1 U8993 ( .A(n7768), .B(n9492), .ZN(n7719) );
  AOI211_X1 U8994 ( .C1(n7874), .C2(n7638), .A(n11212), .B(n5238), .ZN(n7717)
         );
  INV_X1 U8995 ( .A(n7874), .ZN(n7889) );
  NOR2_X1 U8996 ( .A1(n7889), .A2(n10387), .ZN(n7641) );
  OAI22_X1 U8997 ( .A1(n10367), .A2(n7639), .B1(n7883), .B2(n10968), .ZN(n7640) );
  AOI211_X1 U8998 ( .C1(n7717), .C2(n11128), .A(n7641), .B(n7640), .ZN(n7653)
         );
  NAND2_X1 U8999 ( .A1(n8377), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n7649) );
  OR2_X1 U9000 ( .A1(n6968), .A2(n11166), .ZN(n7648) );
  NAND2_X1 U9001 ( .A1(n7642), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7644) );
  INV_X1 U9002 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7643) );
  NAND2_X1 U9003 ( .A1(n7644), .A2(n7643), .ZN(n7645) );
  NAND2_X1 U9004 ( .A1(n7645), .A2(n7760), .ZN(n7936) );
  OR2_X1 U9005 ( .A1(n8382), .A2(n7936), .ZN(n7647) );
  INV_X1 U9006 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n7769) );
  OR2_X1 U9007 ( .A1(n5143), .A2(n7769), .ZN(n7646) );
  NAND2_X1 U9008 ( .A1(n7650), .A2(n9533), .ZN(n7752) );
  XNOR2_X1 U9009 ( .A(n7752), .B(n9492), .ZN(n7651) );
  OAI222_X1 U9010 ( .A1(n11107), .A2(n7981), .B1(n11109), .B2(n7884), .C1(
        n7651), .C2(n11104), .ZN(n7716) );
  NAND2_X1 U9011 ( .A1(n7716), .A2(n10358), .ZN(n7652) );
  OAI211_X1 U9012 ( .C1(n7719), .C2(n10391), .A(n7653), .B(n7652), .ZN(
        P1_U3282) );
  INV_X1 U9013 ( .A(n8213), .ZN(n7656) );
  OAI222_X1 U9014 ( .A1(n9267), .A2(n7655), .B1(n9262), .B2(n7656), .C1(n7654), 
        .C2(P2_U3151), .ZN(P2_U3276) );
  OAI222_X1 U9015 ( .A1(n5141), .A2(n7657), .B1(n10517), .B2(n7656), .C1(
        P1_U3086), .C2(n10163), .ZN(P1_U3336) );
  NAND3_X1 U9016 ( .A1(n7599), .A2(n9204), .A3(n7658), .ZN(n7659) );
  AND2_X1 U9017 ( .A1(n7660), .A2(n7659), .ZN(n7666) );
  INV_X1 U9018 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n7661) );
  NOR2_X1 U9019 ( .A1(n11186), .A2(n7661), .ZN(n7662) );
  AOI21_X1 U9020 ( .B1(n7664), .B2(n6446), .A(n7662), .ZN(n7663) );
  OAI21_X1 U9021 ( .B1(n7666), .B2(n6448), .A(n7663), .ZN(P2_U3417) );
  AOI22_X1 U9022 ( .A1(n7664), .A2(n6400), .B1(n9210), .B2(
        P2_REG1_REG_9__SCAN_IN), .ZN(n7665) );
  OAI21_X1 U9023 ( .B1(n7666), .B2(n9210), .A(n7665), .ZN(P2_U3468) );
  XNOR2_X1 U9024 ( .A(n7667), .B(n8486), .ZN(n7668) );
  OAI222_X1 U9025 ( .A1(n9121), .A2(n7947), .B1(n9119), .B2(n7849), .C1(n9116), 
        .C2(n7668), .ZN(n7746) );
  INV_X1 U9026 ( .A(n7746), .ZN(n7674) );
  OAI21_X1 U9027 ( .B1(n7670), .B2(n8486), .A(n7669), .ZN(n7748) );
  INV_X1 U9028 ( .A(n7854), .ZN(n7745) );
  NOR2_X1 U9029 ( .A1(n7745), .A2(n9141), .ZN(n7672) );
  OAI22_X1 U9030 ( .A1(n9145), .A2(n8890), .B1(n7852), .B2(n9142), .ZN(n7671)
         );
  AOI211_X1 U9031 ( .C1(n7748), .C2(n9148), .A(n7672), .B(n7671), .ZN(n7673)
         );
  OAI21_X1 U9032 ( .B1(n7674), .B2(n9150), .A(n7673), .ZN(P2_U3222) );
  INV_X1 U9033 ( .A(n8233), .ZN(n7694) );
  OAI222_X1 U9034 ( .A1(n5141), .A2(n10021), .B1(n10517), .B2(n7694), .C1(
        n7675), .C2(P1_U3086), .ZN(P1_U3335) );
  NOR2_X1 U9035 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7676), .ZN(n10679) );
  AOI21_X1 U9036 ( .B1(n9367), .B2(n9673), .A(n10679), .ZN(n7678) );
  NAND2_X1 U9037 ( .A1(n9394), .A2(n11065), .ZN(n7677) );
  OAI211_X1 U9038 ( .C1(n9397), .C2(n11121), .A(n7678), .B(n7677), .ZN(n7692)
         );
  OAI21_X1 U9039 ( .B1(n7681), .B2(n7680), .A(n7679), .ZN(n7683) );
  NAND2_X1 U9040 ( .A1(n7681), .A2(n7680), .ZN(n7682) );
  NAND2_X1 U9041 ( .A1(n11125), .A2(n8349), .ZN(n7685) );
  OR2_X1 U9042 ( .A1(n11084), .A2(n5144), .ZN(n7684) );
  NAND2_X1 U9043 ( .A1(n7685), .A2(n7684), .ZN(n7780) );
  NAND2_X1 U9044 ( .A1(n11125), .A2(n8388), .ZN(n7687) );
  OR2_X1 U9045 ( .A1(n11084), .A2(n8390), .ZN(n7686) );
  NAND2_X1 U9046 ( .A1(n7687), .A2(n7686), .ZN(n7688) );
  XNOR2_X1 U9047 ( .A(n7688), .B(n8346), .ZN(n7781) );
  XOR2_X1 U9048 ( .A(n7780), .B(n7781), .Z(n7689) );
  XNOR2_X1 U9049 ( .A(n7782), .B(n7689), .ZN(n7690) );
  NOR2_X1 U9050 ( .A1(n7690), .A2(n9402), .ZN(n7691) );
  AOI211_X1 U9051 ( .C1(n11125), .C2(n9399), .A(n7692), .B(n7691), .ZN(n7693)
         );
  INV_X1 U9052 ( .A(n7693), .ZN(P1_U3221) );
  OAI222_X1 U9053 ( .A1(n9267), .A2(n7695), .B1(P2_U3151), .B2(n8673), .C1(
        n9262), .C2(n7694), .ZN(P2_U3275) );
  XNOR2_X1 U9054 ( .A(n7696), .B(n7698), .ZN(n7905) );
  XNOR2_X1 U9055 ( .A(n7697), .B(n7698), .ZN(n7699) );
  OAI222_X1 U9056 ( .A1(n9119), .A2(n7892), .B1(n9121), .B2(n8110), .C1(n7699), 
        .C2(n9116), .ZN(n7906) );
  NAND2_X1 U9057 ( .A1(n7906), .A2(n9145), .ZN(n7702) );
  OAI22_X1 U9058 ( .A1(n9145), .A2(n8887), .B1(n7898), .B2(n9142), .ZN(n7700)
         );
  AOI21_X1 U9059 ( .B1(n7908), .B2(n9111), .A(n7700), .ZN(n7701) );
  OAI211_X1 U9060 ( .C1(n7905), .C2(n9114), .A(n7702), .B(n7701), .ZN(P2_U3221) );
  NAND2_X1 U9061 ( .A1(n7703), .A2(n8837), .ZN(n7704) );
  XNOR2_X1 U9062 ( .A(n7741), .B(n8440), .ZN(n7845) );
  XNOR2_X1 U9063 ( .A(n7844), .B(n7845), .ZN(n7843) );
  XNOR2_X1 U9064 ( .A(n7843), .B(n8836), .ZN(n7710) );
  AOI22_X1 U9065 ( .A1(n8837), .A2(n8800), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3151), .ZN(n7707) );
  NAND2_X1 U9066 ( .A1(n8835), .A2(n8814), .ZN(n7706) );
  OAI211_X1 U9067 ( .C1(n8756), .C2(n7739), .A(n7707), .B(n7706), .ZN(n7708)
         );
  AOI21_X1 U9068 ( .B1(n7741), .B2(n8805), .A(n7708), .ZN(n7709) );
  OAI21_X1 U9069 ( .B1(n7710), .B2(n8808), .A(n7709), .ZN(P2_U3157) );
  INV_X1 U9070 ( .A(n7711), .ZN(n7712) );
  INV_X1 U9071 ( .A(n9663), .ZN(n10965) );
  OR2_X1 U9072 ( .A1(n6792), .A2(n10965), .ZN(n11091) );
  AOI211_X1 U9073 ( .C1(n11147), .C2(n7874), .A(n7717), .B(n7716), .ZN(n7718)
         );
  OAI21_X1 U9074 ( .B1(n7719), .B2(n11176), .A(n7718), .ZN(n7723) );
  NAND2_X1 U9075 ( .A1(n7723), .A2(n11202), .ZN(n7720) );
  OAI21_X1 U9076 ( .B1(n11202), .B2(n7557), .A(n7720), .ZN(P1_U3533) );
  INV_X1 U9077 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7725) );
  NAND2_X1 U9078 ( .A1(n7723), .A2(n11206), .ZN(n7724) );
  OAI21_X1 U9079 ( .B1(n11206), .B2(n7725), .A(n7724), .ZN(P1_U3486) );
  INV_X1 U9080 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8251) );
  INV_X1 U9081 ( .A(n8250), .ZN(n7750) );
  INV_X1 U9082 ( .A(n9655), .ZN(n7726) );
  OAI222_X1 U9083 ( .A1(n5141), .A2(n8251), .B1(n10517), .B2(n7750), .C1(n7726), .C2(P1_U3086), .ZN(P1_U3334) );
  NAND2_X1 U9084 ( .A1(n7599), .A2(n8516), .ZN(n7727) );
  XNOR2_X1 U9085 ( .A(n7741), .B(n8836), .ZN(n8484) );
  XNOR2_X1 U9086 ( .A(n7727), .B(n8484), .ZN(n7744) );
  NOR2_X1 U9087 ( .A1(n7744), .A2(n7728), .ZN(n7735) );
  INV_X1 U9088 ( .A(n8484), .ZN(n7729) );
  XNOR2_X1 U9089 ( .A(n7730), .B(n7729), .ZN(n7731) );
  NAND2_X1 U9090 ( .A1(n7731), .A2(n9130), .ZN(n7733) );
  AOI22_X1 U9091 ( .A1(n9136), .A2(n8837), .B1(n8835), .B2(n9133), .ZN(n7732)
         );
  OAI211_X1 U9092 ( .C1(n7744), .C2(n7734), .A(n7733), .B(n7732), .ZN(n7737)
         );
  AOI211_X1 U9093 ( .C1(n9180), .C2(n7741), .A(n7735), .B(n7737), .ZN(n11156)
         );
  NAND2_X1 U9094 ( .A1(n9210), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n7736) );
  OAI21_X1 U9095 ( .B1(n11156), .B2(n9210), .A(n7736), .ZN(P2_U3469) );
  MUX2_X1 U9096 ( .A(n7737), .B(P2_REG2_REG_10__SCAN_IN), .S(n9150), .Z(n7738)
         );
  INV_X1 U9097 ( .A(n7738), .ZN(n7743) );
  INV_X1 U9098 ( .A(n7739), .ZN(n7740) );
  AOI22_X1 U9099 ( .A1(n7741), .A2(n9111), .B1(n9125), .B2(n7740), .ZN(n7742)
         );
  OAI211_X1 U9100 ( .C1(n7744), .C2(n8988), .A(n7743), .B(n7742), .ZN(P2_U3223) );
  NOR2_X1 U9101 ( .A1(n7745), .A2(n9173), .ZN(n7747) );
  AOI211_X1 U9102 ( .C1(n9204), .C2(n7748), .A(n7747), .B(n7746), .ZN(n11158)
         );
  OR2_X1 U9103 ( .A1(n11158), .A2(n9210), .ZN(n7749) );
  OAI21_X1 U9104 ( .B1(n9206), .B2(n8889), .A(n7749), .ZN(P2_U3470) );
  OAI222_X1 U9105 ( .A1(n9267), .A2(n7751), .B1(P2_U3151), .B2(n5140), .C1(
        n9262), .C2(n7750), .ZN(P2_U3274) );
  NAND2_X1 U9106 ( .A1(n7752), .A2(n9522), .ZN(n7753) );
  AOI22_X1 U9107 ( .A1(n8215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n8214), .B2(
        n10122), .ZN(n7755) );
  NAND2_X1 U9108 ( .A1(n7929), .A2(n7981), .ZN(n9518) );
  NAND2_X1 U9109 ( .A1(n9577), .A2(n9518), .ZN(n9490) );
  INV_X1 U9110 ( .A(n7759), .ZN(n7758) );
  INV_X1 U9111 ( .A(n9490), .ZN(n7757) );
  INV_X1 U9112 ( .A(n7799), .ZN(n7796) );
  AOI211_X1 U9113 ( .C1(n7759), .C2(n9490), .A(n11104), .B(n7796), .ZN(n7767)
         );
  NAND2_X1 U9114 ( .A1(n8377), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n7765) );
  INV_X1 U9115 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7809) );
  OR2_X1 U9116 ( .A1(n5143), .A2(n7809), .ZN(n7764) );
  NAND2_X1 U9117 ( .A1(n7760), .A2(n7979), .ZN(n7761) );
  NAND2_X1 U9118 ( .A1(n7803), .A2(n7761), .ZN(n7978) );
  OR2_X1 U9119 ( .A1(n8382), .A2(n7978), .ZN(n7763) );
  INV_X1 U9120 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n10111) );
  OR2_X1 U9121 ( .A1(n6968), .A2(n10111), .ZN(n7762) );
  OAI22_X1 U9122 ( .A1(n7872), .A2(n11109), .B1(n8119), .B2(n11107), .ZN(n7766) );
  NOR2_X1 U9123 ( .A1(n7767), .A2(n7766), .ZN(n11162) );
  XOR2_X1 U9124 ( .A(n9490), .B(n7791), .Z(n11165) );
  NAND2_X1 U9125 ( .A1(n11165), .A2(n11129), .ZN(n7774) );
  OAI22_X1 U9126 ( .A1(n10367), .A2(n7769), .B1(n7936), .B2(n10968), .ZN(n7772) );
  INV_X1 U9127 ( .A(n7801), .ZN(n7770) );
  OAI211_X1 U9128 ( .C1(n11163), .C2(n5238), .A(n7770), .B(n5131), .ZN(n11161)
         );
  NOR2_X1 U9129 ( .A1(n11161), .A2(n10333), .ZN(n7771) );
  AOI211_X1 U9130 ( .C1(n11124), .C2(n7929), .A(n7772), .B(n7771), .ZN(n7773)
         );
  OAI211_X1 U9131 ( .C1(n7171), .C2(n11162), .A(n7774), .B(n7773), .ZN(
        P1_U3281) );
  AOI21_X1 U9132 ( .B1(n9394), .B2(n11136), .A(n7775), .ZN(n7778) );
  NAND2_X1 U9133 ( .A1(n9367), .A2(n7776), .ZN(n7777) );
  OAI211_X1 U9134 ( .C1(n9397), .C2(n7779), .A(n7778), .B(n7777), .ZN(n7789)
         );
  NAND2_X1 U9135 ( .A1(n11137), .A2(n8388), .ZN(n7784) );
  OR2_X1 U9136 ( .A1(n11108), .A2(n8390), .ZN(n7783) );
  NAND2_X1 U9137 ( .A1(n7784), .A2(n7783), .ZN(n7785) );
  XNOR2_X1 U9138 ( .A(n7785), .B(n8314), .ZN(n7824) );
  NOR2_X1 U9139 ( .A1(n11108), .A2(n5144), .ZN(n7786) );
  AOI21_X1 U9140 ( .B1(n11137), .B2(n8349), .A(n7786), .ZN(n7823) );
  XNOR2_X1 U9141 ( .A(n7824), .B(n7823), .ZN(n7826) );
  XOR2_X1 U9142 ( .A(n7827), .B(n7826), .Z(n7787) );
  NOR2_X1 U9143 ( .A1(n7787), .A2(n9402), .ZN(n7788) );
  AOI211_X1 U9144 ( .C1(n11137), .C2(n9399), .A(n7789), .B(n7788), .ZN(n7790)
         );
  INV_X1 U9145 ( .A(n7790), .ZN(P1_U3231) );
  INV_X1 U9146 ( .A(n7981), .ZN(n11171) );
  NAND2_X1 U9147 ( .A1(n7793), .A2(n8029), .ZN(n7795) );
  AOI22_X1 U9148 ( .A1(n8215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n8214), .B2(
        n10743), .ZN(n7794) );
  OR2_X1 U9149 ( .A1(n7992), .A2(n8119), .ZN(n9583) );
  NAND2_X1 U9150 ( .A1(n7992), .A2(n8119), .ZN(n9575) );
  NAND2_X1 U9151 ( .A1(n9583), .A2(n9575), .ZN(n9493) );
  XNOR2_X1 U9152 ( .A(n7991), .B(n9493), .ZN(n11177) );
  INV_X1 U9153 ( .A(n9577), .ZN(n7797) );
  OAI21_X1 U9154 ( .B1(n7796), .B2(n7797), .A(n9493), .ZN(n7800) );
  NOR2_X1 U9155 ( .A1(n9493), .A2(n7797), .ZN(n7798) );
  NAND2_X1 U9156 ( .A1(n7800), .A2(n7986), .ZN(n11180) );
  OAI211_X1 U9157 ( .C1(n7801), .C2(n11175), .A(n8003), .B(n5131), .ZN(n11174)
         );
  NAND2_X1 U9158 ( .A1(n8377), .A2(P1_REG0_REG_14__SCAN_IN), .ZN(n7808) );
  INV_X1 U9159 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n8000) );
  OR2_X1 U9160 ( .A1(n5143), .A2(n8000), .ZN(n7807) );
  AND2_X1 U9161 ( .A1(n7803), .A2(n7802), .ZN(n7804) );
  OR2_X1 U9162 ( .A1(n7994), .A2(n7804), .ZN(n8067) );
  OR2_X1 U9163 ( .A1(n8382), .A2(n8067), .ZN(n7806) );
  INV_X1 U9164 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10113) );
  OR2_X1 U9165 ( .A1(n6968), .A2(n10113), .ZN(n7805) );
  OAI22_X1 U9166 ( .A1(n10367), .A2(n7809), .B1(n7978), .B2(n10968), .ZN(n7810) );
  AOI21_X1 U9167 ( .B1(n10326), .B2(n11171), .A(n7810), .ZN(n7811) );
  OAI21_X1 U9168 ( .B1(n8062), .B2(n10328), .A(n7811), .ZN(n7812) );
  AOI21_X1 U9169 ( .B1(n7992), .B2(n11124), .A(n7812), .ZN(n7813) );
  OAI21_X1 U9170 ( .B1(n11174), .B2(n10333), .A(n7813), .ZN(n7814) );
  AOI21_X1 U9171 ( .B1(n11180), .B2(n10335), .A(n7814), .ZN(n7815) );
  OAI21_X1 U9172 ( .B1(n11177), .B2(n10391), .A(n7815), .ZN(P1_U3280) );
  INV_X1 U9173 ( .A(n7816), .ZN(n8590) );
  XNOR2_X1 U9174 ( .A(n7817), .B(n8589), .ZN(n7861) );
  XNOR2_X1 U9175 ( .A(n7818), .B(n8589), .ZN(n7819) );
  OAI222_X1 U9176 ( .A1(n9121), .A2(n8817), .B1(n9119), .B2(n7947), .C1(n7819), 
        .C2(n9116), .ZN(n7863) );
  OAI22_X1 U9177 ( .A1(n7860), .A2(n9040), .B1(n7950), .B2(n9142), .ZN(n7820)
         );
  OAI21_X1 U9178 ( .B1(n7863), .B2(n7820), .A(n9145), .ZN(n7822) );
  NAND2_X1 U9179 ( .A1(n9150), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n7821) );
  OAI211_X1 U9180 ( .C1(n7861), .C2(n9114), .A(n7822), .B(n7821), .ZN(P2_U3220) );
  NAND2_X1 U9181 ( .A1(n7824), .A2(n7823), .ZN(n7825) );
  NAND2_X1 U9182 ( .A1(n11148), .A2(n8388), .ZN(n7829) );
  OR2_X1 U9183 ( .A1(n7884), .A2(n8390), .ZN(n7828) );
  NAND2_X1 U9184 ( .A1(n7829), .A2(n7828), .ZN(n7830) );
  XNOR2_X1 U9185 ( .A(n7830), .B(n8314), .ZN(n7831) );
  NAND2_X1 U9186 ( .A1(n7832), .A2(n7831), .ZN(n7867) );
  NAND2_X1 U9187 ( .A1(n7866), .A2(n7867), .ZN(n7834) );
  NOR2_X1 U9188 ( .A1(n7884), .A2(n5144), .ZN(n7833) );
  AOI21_X1 U9189 ( .B1(n11148), .B2(n8349), .A(n7833), .ZN(n7865) );
  XNOR2_X1 U9190 ( .A(n7834), .B(n7865), .ZN(n7842) );
  INV_X1 U9191 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7835) );
  NOR2_X1 U9192 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7835), .ZN(n7837) );
  NOR2_X1 U9193 ( .A1(n9391), .A2(n7872), .ZN(n7836) );
  AOI211_X1 U9194 ( .C1(n9394), .C2(n9673), .A(n7837), .B(n7836), .ZN(n7838)
         );
  OAI21_X1 U9195 ( .B1(n9397), .B2(n7839), .A(n7838), .ZN(n7840) );
  AOI21_X1 U9196 ( .B1(n11148), .B2(n9399), .A(n7840), .ZN(n7841) );
  OAI21_X1 U9197 ( .B1(n7842), .B2(n9402), .A(n7841), .ZN(P1_U3217) );
  NAND2_X1 U9198 ( .A1(n7843), .A2(n7849), .ZN(n7848) );
  INV_X1 U9199 ( .A(n7844), .ZN(n7846) );
  NAND2_X1 U9200 ( .A1(n7846), .A2(n7845), .ZN(n7847) );
  NAND2_X1 U9201 ( .A1(n7848), .A2(n7847), .ZN(n7891) );
  XNOR2_X1 U9202 ( .A(n7854), .B(n8440), .ZN(n7893) );
  XNOR2_X1 U9203 ( .A(n7893), .B(n8835), .ZN(n7890) );
  XOR2_X1 U9204 ( .A(n7891), .B(n7890), .Z(n7856) );
  INV_X1 U9205 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9984) );
  OAI22_X1 U9206 ( .A1(n7849), .A2(n8816), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n9984), .ZN(n7850) );
  AOI21_X1 U9207 ( .B1(n8814), .B2(n8834), .A(n7850), .ZN(n7851) );
  OAI21_X1 U9208 ( .B1(n7852), .B2(n8756), .A(n7851), .ZN(n7853) );
  AOI21_X1 U9209 ( .B1(n7854), .B2(n8805), .A(n7853), .ZN(n7855) );
  OAI21_X1 U9210 ( .B1(n7856), .B2(n8808), .A(n7855), .ZN(P2_U3176) );
  INV_X1 U9211 ( .A(n8272), .ZN(n7858) );
  INV_X1 U9212 ( .A(n6792), .ZN(n9647) );
  OAI222_X1 U9213 ( .A1(n5141), .A2(n9805), .B1(n10517), .B2(n7858), .C1(
        P1_U3086), .C2(n9647), .ZN(P1_U3333) );
  OAI222_X1 U9214 ( .A1(n9267), .A2(n7859), .B1(n9262), .B2(n7858), .C1(
        P2_U3151), .C2(n7857), .ZN(P2_U3273) );
  OAI22_X1 U9215 ( .A1(n7861), .A2(n9188), .B1(n7860), .B2(n9173), .ZN(n7862)
         );
  NOR2_X1 U9216 ( .A1(n7863), .A2(n7862), .ZN(n11185) );
  OR2_X1 U9217 ( .A1(n9206), .A2(n8883), .ZN(n7864) );
  OAI21_X1 U9218 ( .B1(n11185), .B2(n9210), .A(n7864), .ZN(P2_U3472) );
  INV_X1 U9219 ( .A(n9399), .ZN(n9385) );
  NAND2_X1 U9220 ( .A1(n7866), .A2(n7865), .ZN(n7868) );
  NAND2_X1 U9221 ( .A1(n7868), .A2(n7867), .ZN(n7879) );
  NAND2_X1 U9222 ( .A1(n7874), .A2(n8388), .ZN(n7870) );
  OR2_X1 U9223 ( .A1(n7872), .A2(n8390), .ZN(n7869) );
  NAND2_X1 U9224 ( .A1(n7870), .A2(n7869), .ZN(n7871) );
  XNOR2_X1 U9225 ( .A(n7871), .B(n8314), .ZN(n7875) );
  NOR2_X1 U9226 ( .A1(n7872), .A2(n5144), .ZN(n7873) );
  AOI21_X1 U9227 ( .B1(n7874), .B2(n8349), .A(n7873), .ZN(n7876) );
  AND2_X1 U9228 ( .A1(n7875), .A2(n7876), .ZN(n7880) );
  INV_X1 U9229 ( .A(n7875), .ZN(n7878) );
  INV_X1 U9230 ( .A(n7876), .ZN(n7877) );
  NAND2_X1 U9231 ( .A1(n7878), .A2(n7877), .ZN(n7933) );
  INV_X1 U9232 ( .A(n7933), .ZN(n7882) );
  OAI21_X1 U9233 ( .B1(n7880), .B2(n7882), .A(n7879), .ZN(n7881) );
  OAI211_X1 U9234 ( .C1(n7931), .C2(n7882), .A(n9376), .B(n7881), .ZN(n7888)
         );
  NOR2_X1 U9235 ( .A1(n9397), .A2(n7883), .ZN(n7886) );
  NAND2_X1 U9236 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n10691) );
  OAI21_X1 U9237 ( .B1(n9369), .B2(n7884), .A(n10691), .ZN(n7885) );
  AOI211_X1 U9238 ( .C1(n9367), .C2(n11171), .A(n7886), .B(n7885), .ZN(n7887)
         );
  OAI211_X1 U9239 ( .C1(n7889), .C2(n9385), .A(n7888), .B(n7887), .ZN(P1_U3236) );
  INV_X1 U9240 ( .A(n7908), .ZN(n7904) );
  NAND2_X1 U9241 ( .A1(n7893), .A2(n7892), .ZN(n7894) );
  XNOR2_X1 U9242 ( .A(n7908), .B(n8424), .ZN(n7943) );
  XNOR2_X1 U9243 ( .A(n7943), .B(n8834), .ZN(n7896) );
  AOI21_X1 U9244 ( .B1(n7895), .B2(n7896), .A(n8808), .ZN(n7897) );
  NAND2_X1 U9245 ( .A1(n7897), .A2(n7945), .ZN(n7903) );
  INV_X1 U9246 ( .A(n7898), .ZN(n7901) );
  NOR2_X1 U9247 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9967), .ZN(n10821) );
  AOI21_X1 U9248 ( .B1(n8835), .B2(n8800), .A(n10821), .ZN(n7899) );
  OAI21_X1 U9249 ( .B1(n8110), .B2(n8803), .A(n7899), .ZN(n7900) );
  AOI21_X1 U9250 ( .B1(n7901), .B2(n8819), .A(n7900), .ZN(n7902) );
  OAI211_X1 U9251 ( .C1(n7904), .C2(n8823), .A(n7903), .B(n7902), .ZN(P2_U3164) );
  NOR2_X1 U9252 ( .A1(n7905), .A2(n9188), .ZN(n7907) );
  AOI211_X1 U9253 ( .C1(n9180), .C2(n7908), .A(n7907), .B(n7906), .ZN(n11160)
         );
  OR2_X1 U9254 ( .A1(n11160), .A2(n9210), .ZN(n7909) );
  OAI21_X1 U9255 ( .B1(n9206), .B2(n8886), .A(n7909), .ZN(P2_U3471) );
  NAND2_X1 U9256 ( .A1(n8292), .A2(n9263), .ZN(n7911) );
  INV_X1 U9257 ( .A(n7910), .ZN(n8696) );
  OAI211_X1 U9258 ( .C1(n7912), .C2(n9267), .A(n7911), .B(n8696), .ZN(P2_U3272) );
  NAND2_X1 U9259 ( .A1(n8292), .A2(n10513), .ZN(n7914) );
  NAND2_X1 U9260 ( .A1(n7913), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9662) );
  OAI211_X1 U9261 ( .C1(n10017), .C2(n5141), .A(n7914), .B(n9662), .ZN(
        P1_U3332) );
  NAND2_X1 U9262 ( .A1(n7915), .A2(n8594), .ZN(n7916) );
  NAND3_X1 U9263 ( .A1(n7917), .A2(n9130), .A3(n7916), .ZN(n7919) );
  AOI22_X1 U9264 ( .A1(n8833), .A2(n9136), .B1(n9133), .B2(n8831), .ZN(n7918)
         );
  AND2_X1 U9265 ( .A1(n7919), .A2(n7918), .ZN(n8049) );
  INV_X1 U9266 ( .A(n8049), .ZN(n7921) );
  INV_X1 U9267 ( .A(n8115), .ZN(n8595) );
  OAI22_X1 U9268 ( .A1(n8595), .A2(n9040), .B1(n8113), .B2(n9142), .ZN(n7920)
         );
  OAI21_X1 U9269 ( .B1(n7921), .B2(n7920), .A(n9145), .ZN(n7924) );
  XNOR2_X1 U9270 ( .A(n7922), .B(n6110), .ZN(n8047) );
  AOI22_X1 U9271 ( .A1(n8047), .A2(n9148), .B1(P2_REG2_REG_14__SCAN_IN), .B2(
        n9150), .ZN(n7923) );
  NAND2_X1 U9272 ( .A1(n7924), .A2(n7923), .ZN(P2_U3219) );
  NAND2_X1 U9273 ( .A1(n7929), .A2(n8388), .ZN(n7926) );
  OR2_X1 U9274 ( .A1(n7981), .A2(n8390), .ZN(n7925) );
  NAND2_X1 U9275 ( .A1(n7926), .A2(n7925), .ZN(n7927) );
  XNOR2_X1 U9276 ( .A(n7927), .B(n8346), .ZN(n7966) );
  NOR2_X1 U9277 ( .A1(n7981), .A2(n5144), .ZN(n7928) );
  AOI21_X1 U9278 ( .B1(n7929), .B2(n8349), .A(n7928), .ZN(n7967) );
  XNOR2_X1 U9279 ( .A(n7966), .B(n7967), .ZN(n7932) );
  AND2_X1 U9280 ( .A1(n7932), .A2(n7933), .ZN(n7930) );
  NAND2_X2 U9281 ( .A1(n7931), .A2(n7930), .ZN(n7975) );
  INV_X1 U9282 ( .A(n7975), .ZN(n7935) );
  AOI21_X1 U9283 ( .B1(n7931), .B2(n7933), .A(n7932), .ZN(n7934) );
  OAI21_X1 U9284 ( .B1(n7935), .B2(n7934), .A(n9376), .ZN(n7942) );
  INV_X1 U9285 ( .A(n7936), .ZN(n7940) );
  AOI21_X1 U9286 ( .B1(n9394), .B2(n11146), .A(n7937), .ZN(n7938) );
  OAI21_X1 U9287 ( .B1(n8119), .B2(n9391), .A(n7938), .ZN(n7939) );
  AOI21_X1 U9288 ( .B1(n7940), .B2(n9381), .A(n7939), .ZN(n7941) );
  OAI211_X1 U9289 ( .C1(n11163), .C2(n9385), .A(n7942), .B(n7941), .ZN(
        P1_U3224) );
  NAND2_X1 U9290 ( .A1(n7943), .A2(n8834), .ZN(n7944) );
  NAND2_X1 U9291 ( .A1(n7945), .A2(n7944), .ZN(n8099) );
  XNOR2_X1 U9292 ( .A(n7952), .B(n8440), .ZN(n8100) );
  XNOR2_X1 U9293 ( .A(n8100), .B(n8833), .ZN(n7946) );
  XNOR2_X1 U9294 ( .A(n8099), .B(n7946), .ZN(n7954) );
  NOR2_X1 U9295 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5738), .ZN(n10837) );
  NOR2_X1 U9296 ( .A1(n7947), .A2(n8816), .ZN(n7948) );
  AOI211_X1 U9297 ( .C1(n8814), .C2(n8832), .A(n10837), .B(n7948), .ZN(n7949)
         );
  OAI21_X1 U9298 ( .B1(n7950), .B2(n8756), .A(n7949), .ZN(n7951) );
  AOI21_X1 U9299 ( .B1(n7952), .B2(n8805), .A(n7951), .ZN(n7953) );
  OAI21_X1 U9300 ( .B1(n7954), .B2(n8808), .A(n7953), .ZN(P2_U3174) );
  OAI211_X1 U9301 ( .C1(n7956), .C2(n8607), .A(n7955), .B(n9130), .ZN(n7958)
         );
  AOI22_X1 U9302 ( .A1(n9136), .A2(n8832), .B1(n9135), .B2(n9133), .ZN(n7957)
         );
  NAND2_X1 U9303 ( .A1(n7958), .A2(n7957), .ZN(n8072) );
  INV_X1 U9304 ( .A(n8072), .ZN(n7965) );
  OAI21_X1 U9305 ( .B1(n7960), .B2(n6330), .A(n7959), .ZN(n8073) );
  INV_X1 U9306 ( .A(n7961), .ZN(n8820) );
  AOI22_X1 U9307 ( .A1(n9150), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n9125), .B2(
        n8820), .ZN(n7962) );
  OAI21_X1 U9308 ( .B1(n8824), .B2(n9141), .A(n7962), .ZN(n7963) );
  AOI21_X1 U9309 ( .B1(n8073), .B2(n9148), .A(n7963), .ZN(n7964) );
  OAI21_X1 U9310 ( .B1(n7965), .B2(n9150), .A(n7964), .ZN(P2_U3218) );
  INV_X1 U9311 ( .A(n7966), .ZN(n7968) );
  NAND2_X1 U9312 ( .A1(n7968), .A2(n7967), .ZN(n7973) );
  AND2_X1 U9313 ( .A1(n7975), .A2(n7973), .ZN(n7977) );
  NAND2_X1 U9314 ( .A1(n7992), .A2(n8388), .ZN(n7970) );
  OR2_X1 U9315 ( .A1(n8119), .A2(n8390), .ZN(n7969) );
  NAND2_X1 U9316 ( .A1(n7970), .A2(n7969), .ZN(n7971) );
  XNOR2_X1 U9317 ( .A(n7971), .B(n8346), .ZN(n8055) );
  NOR2_X1 U9318 ( .A1(n8119), .A2(n5144), .ZN(n7972) );
  AOI21_X1 U9319 ( .B1(n7992), .B2(n8349), .A(n7972), .ZN(n8056) );
  XNOR2_X1 U9320 ( .A(n8055), .B(n8056), .ZN(n7976) );
  AND2_X1 U9321 ( .A1(n7976), .A2(n7973), .ZN(n7974) );
  OAI211_X1 U9322 ( .C1(n7977), .C2(n7976), .A(n9376), .B(n8058), .ZN(n7985)
         );
  INV_X1 U9323 ( .A(n7978), .ZN(n7983) );
  INV_X1 U9324 ( .A(n8062), .ZN(n11170) );
  NOR2_X1 U9325 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7979), .ZN(n10746) );
  AOI21_X1 U9326 ( .B1(n9367), .B2(n11170), .A(n10746), .ZN(n7980) );
  OAI21_X1 U9327 ( .B1(n9369), .B2(n7981), .A(n7980), .ZN(n7982) );
  AOI21_X1 U9328 ( .B1(n7983), .B2(n9381), .A(n7982), .ZN(n7984) );
  OAI211_X1 U9329 ( .C1(n11175), .C2(n9385), .A(n7985), .B(n7984), .ZN(
        P1_U3234) );
  NAND2_X1 U9330 ( .A1(n7987), .A2(n8029), .ZN(n7989) );
  AOI22_X1 U9331 ( .A1(n8215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n8214), .B2(
        n10699), .ZN(n7988) );
  NAND2_X1 U9332 ( .A1(n8121), .A2(n8062), .ZN(n9585) );
  NAND2_X1 U9333 ( .A1(n9587), .A2(n9585), .ZN(n9494) );
  OAI211_X1 U9334 ( .C1(n5235), .C2(n7990), .A(n8028), .B(n11181), .ZN(n8123)
         );
  INV_X1 U9335 ( .A(n8119), .ZN(n9672) );
  XOR2_X1 U9336 ( .A(n9494), .B(n8037), .Z(n8118) );
  NAND2_X1 U9337 ( .A1(n8118), .A2(n11129), .ZN(n8008) );
  NAND2_X1 U9338 ( .A1(n8377), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7999) );
  INV_X1 U9339 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7993) );
  OR2_X1 U9340 ( .A1(n6968), .A2(n7993), .ZN(n7998) );
  OR2_X1 U9341 ( .A1(n7994), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7995) );
  NAND2_X1 U9342 ( .A1(n8020), .A2(n7995), .ZN(n9396) );
  OR2_X1 U9343 ( .A1(n8382), .A2(n9396), .ZN(n7997) );
  INV_X1 U9344 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n8038) );
  OR2_X1 U9345 ( .A1(n5143), .A2(n8038), .ZN(n7996) );
  OAI22_X1 U9346 ( .A1(n10358), .A2(n8000), .B1(n8067), .B2(n10968), .ZN(n8001) );
  AOI21_X1 U9347 ( .B1(n10326), .B2(n9672), .A(n8001), .ZN(n8002) );
  OAI21_X1 U9348 ( .B1(n8178), .B2(n10328), .A(n8002), .ZN(n8006) );
  AOI21_X1 U9349 ( .B1(n8003), .B2(n8121), .A(n11212), .ZN(n8004) );
  NAND2_X1 U9350 ( .A1(n8004), .A2(n8039), .ZN(n8122) );
  NOR2_X1 U9351 ( .A1(n8122), .A2(n10333), .ZN(n8005) );
  AOI211_X1 U9352 ( .C1(n11124), .C2(n8121), .A(n8006), .B(n8005), .ZN(n8007)
         );
  OAI211_X1 U9353 ( .C1(n7171), .C2(n8123), .A(n8008), .B(n8007), .ZN(P1_U3279) );
  INV_X1 U9354 ( .A(n6571), .ZN(n8009) );
  INV_X1 U9355 ( .A(n8300), .ZN(n8081) );
  OAI222_X1 U9356 ( .A1(n5141), .A2(n9801), .B1(P1_U3086), .B2(n8009), .C1(
        n8081), .C2(n10517), .ZN(P1_U3331) );
  OAI21_X1 U9357 ( .B1(n8011), .B2(n8489), .A(n8010), .ZN(n9202) );
  OAI211_X1 U9358 ( .C1(n8013), .C2(n8608), .A(n8012), .B(n9130), .ZN(n8015)
         );
  AOI22_X1 U9359 ( .A1(n9133), .A2(n8830), .B1(n8831), .B2(n9136), .ZN(n8014)
         );
  NAND2_X1 U9360 ( .A1(n8015), .A2(n8014), .ZN(n9203) );
  NAND2_X1 U9361 ( .A1(n9203), .A2(n9145), .ZN(n8018) );
  OAI22_X1 U9362 ( .A1(n9145), .A2(n8936), .B1(n8745), .B2(n9142), .ZN(n8016)
         );
  AOI21_X1 U9363 ( .B1(n8739), .B2(n9111), .A(n8016), .ZN(n8017) );
  OAI211_X1 U9364 ( .C1(n9202), .C2(n9114), .A(n8018), .B(n8017), .ZN(P2_U3217) );
  NAND2_X1 U9365 ( .A1(n8377), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8027) );
  INV_X1 U9366 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n8019) );
  OR2_X1 U9367 ( .A1(n6968), .A2(n8019), .ZN(n8026) );
  NAND2_X1 U9368 ( .A1(n8020), .A2(n9317), .ZN(n8023) );
  INV_X1 U9369 ( .A(n8021), .ZN(n8022) );
  NAND2_X1 U9370 ( .A1(n8023), .A2(n8022), .ZN(n9320) );
  OR2_X1 U9371 ( .A1(n8382), .A2(n9320), .ZN(n8025) );
  INV_X1 U9372 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n8092) );
  OR2_X1 U9373 ( .A1(n5143), .A2(n8092), .ZN(n8024) );
  NAND2_X1 U9374 ( .A1(n8030), .A2(n8029), .ZN(n8032) );
  AOI22_X1 U9375 ( .A1(n8215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8214), .B2(
        n10718), .ZN(n8031) );
  NAND2_X1 U9376 ( .A1(n9400), .A2(n8178), .ZN(n9593) );
  OAI211_X1 U9377 ( .C1(n8033), .C2(n9496), .A(n8087), .B(n11181), .ZN(n8035)
         );
  OR2_X1 U9378 ( .A1(n8062), .A2(n11109), .ZN(n8034) );
  OAI211_X1 U9379 ( .C1(n9390), .C2(n11107), .A(n8035), .B(n8034), .ZN(n11190)
         );
  INV_X1 U9380 ( .A(n11190), .ZN(n8046) );
  XOR2_X1 U9381 ( .A(n8083), .B(n9496), .Z(n11191) );
  NAND2_X1 U9382 ( .A1(n11191), .A2(n11129), .ZN(n8045) );
  OAI22_X1 U9383 ( .A1(n10358), .A2(n8038), .B1(n9396), .B2(n10968), .ZN(n8043) );
  INV_X1 U9384 ( .A(n9400), .ZN(n11188) );
  INV_X1 U9385 ( .A(n8039), .ZN(n8041) );
  INV_X1 U9386 ( .A(n8091), .ZN(n8040) );
  OAI211_X1 U9387 ( .C1(n11188), .C2(n8041), .A(n8040), .B(n5131), .ZN(n11187)
         );
  NOR2_X1 U9388 ( .A1(n11187), .A2(n10333), .ZN(n8042) );
  AOI211_X1 U9389 ( .C1(n11124), .C2(n9400), .A(n8043), .B(n8042), .ZN(n8044)
         );
  OAI211_X1 U9390 ( .C1(n7171), .C2(n8046), .A(n8045), .B(n8044), .ZN(P1_U3278) );
  NAND2_X1 U9391 ( .A1(n8047), .A2(n9204), .ZN(n8048) );
  NAND2_X1 U9392 ( .A1(n8049), .A2(n8048), .ZN(n8052) );
  MUX2_X1 U9393 ( .A(P2_REG0_REG_14__SCAN_IN), .B(n8052), .S(n11186), .Z(n8050) );
  AOI21_X1 U9394 ( .B1(n6446), .B2(n8115), .A(n8050), .ZN(n8051) );
  INV_X1 U9395 ( .A(n8051), .ZN(P2_U3432) );
  MUX2_X1 U9396 ( .A(n8052), .B(P2_REG1_REG_14__SCAN_IN), .S(n9210), .Z(n8053)
         );
  AOI21_X1 U9397 ( .B1(n6400), .B2(n8115), .A(n8053), .ZN(n8054) );
  INV_X1 U9398 ( .A(n8054), .ZN(P2_U3473) );
  INV_X1 U9399 ( .A(n8055), .ZN(n8057) );
  NAND2_X1 U9400 ( .A1(n8121), .A2(n8388), .ZN(n8060) );
  OR2_X1 U9401 ( .A1(n8062), .A2(n8390), .ZN(n8059) );
  NAND2_X1 U9402 ( .A1(n8060), .A2(n8059), .ZN(n8061) );
  XNOR2_X1 U9403 ( .A(n8061), .B(n8314), .ZN(n8172) );
  NOR2_X1 U9404 ( .A1(n8062), .A2(n5144), .ZN(n8063) );
  AOI21_X1 U9405 ( .B1(n8121), .B2(n8349), .A(n8063), .ZN(n8169) );
  INV_X1 U9406 ( .A(n8169), .ZN(n8173) );
  XNOR2_X1 U9407 ( .A(n8172), .B(n8173), .ZN(n8064) );
  XNOR2_X1 U9408 ( .A(n8171), .B(n8064), .ZN(n8070) );
  INV_X1 U9409 ( .A(n8178), .ZN(n9671) );
  NAND2_X1 U9410 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n10709) );
  OAI21_X1 U9411 ( .B1(n9369), .B2(n8119), .A(n10709), .ZN(n8065) );
  AOI21_X1 U9412 ( .B1(n9367), .B2(n9671), .A(n8065), .ZN(n8066) );
  OAI21_X1 U9413 ( .B1(n9397), .B2(n8067), .A(n8066), .ZN(n8068) );
  AOI21_X1 U9414 ( .B1(n8121), .B2(n9399), .A(n8068), .ZN(n8069) );
  OAI21_X1 U9415 ( .B1(n8070), .B2(n9402), .A(n8069), .ZN(P1_U3215) );
  INV_X1 U9416 ( .A(n8319), .ZN(n8078) );
  OAI222_X1 U9417 ( .A1(P1_U3086), .A2(n8071), .B1(n10517), .B2(n8078), .C1(
        n10013), .C2(n5141), .ZN(P1_U3330) );
  INV_X1 U9418 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n8074) );
  AOI21_X1 U9419 ( .B1(n9204), .B2(n8073), .A(n8072), .ZN(n8076) );
  MUX2_X1 U9420 ( .A(n8074), .B(n8076), .S(n11186), .Z(n8075) );
  OAI21_X1 U9421 ( .B1(n8824), .B2(n9250), .A(n8075), .ZN(P2_U3435) );
  MUX2_X1 U9422 ( .A(n8879), .B(n8076), .S(n9206), .Z(n8077) );
  OAI21_X1 U9423 ( .B1(n8824), .B2(n9209), .A(n8077), .ZN(P2_U3474) );
  OAI222_X1 U9424 ( .A1(n9267), .A2(n8080), .B1(P2_U3151), .B2(n8079), .C1(
        n9262), .C2(n8078), .ZN(P2_U3270) );
  OAI222_X1 U9425 ( .A1(n9267), .A2(n8082), .B1(P2_U3151), .B2(n6354), .C1(
        n9262), .C2(n8081), .ZN(P2_U3271) );
  NAND2_X1 U9426 ( .A1(n8084), .A2(n8029), .ZN(n8086) );
  AOI22_X1 U9427 ( .A1(n8215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n8214), .B2(
        n10140), .ZN(n8085) );
  NAND2_X1 U9428 ( .A1(n9322), .A2(n9390), .ZN(n9594) );
  XNOR2_X1 U9429 ( .A(n8131), .B(n9497), .ZN(n11200) );
  INV_X1 U9430 ( .A(n11200), .ZN(n8097) );
  NAND2_X1 U9431 ( .A1(n8087), .A2(n9591), .ZN(n8088) );
  NAND2_X1 U9432 ( .A1(n8088), .A2(n9497), .ZN(n8149) );
  OAI211_X1 U9433 ( .C1(n8088), .C2(n9497), .A(n8149), .B(n11181), .ZN(n8090)
         );
  NAND2_X1 U9434 ( .A1(n9671), .A2(n11172), .ZN(n8089) );
  OAI211_X1 U9435 ( .C1(n10378), .C2(n11107), .A(n8090), .B(n8089), .ZN(n11198) );
  INV_X1 U9436 ( .A(n9322), .ZN(n11196) );
  INV_X1 U9437 ( .A(n8135), .ZN(n8137) );
  OAI211_X1 U9438 ( .C1(n11196), .C2(n8091), .A(n8137), .B(n5131), .ZN(n11194)
         );
  OAI22_X1 U9439 ( .A1(n10358), .A2(n8092), .B1(n9320), .B2(n10968), .ZN(n8093) );
  AOI21_X1 U9440 ( .B1(n9322), .B2(n11124), .A(n8093), .ZN(n8094) );
  OAI21_X1 U9441 ( .B1(n11194), .B2(n10333), .A(n8094), .ZN(n8095) );
  AOI21_X1 U9442 ( .B1(n11198), .B2(n10358), .A(n8095), .ZN(n8096) );
  OAI21_X1 U9443 ( .B1(n8097), .B2(n10391), .A(n8096), .ZN(P1_U3277) );
  XNOR2_X1 U9444 ( .A(n8115), .B(n8424), .ZN(n8400) );
  XNOR2_X1 U9445 ( .A(n8400), .B(n8832), .ZN(n8108) );
  NAND2_X1 U9446 ( .A1(n8100), .A2(n8110), .ZN(n8098) );
  NAND2_X1 U9447 ( .A1(n8099), .A2(n8098), .ZN(n8103) );
  INV_X1 U9448 ( .A(n8100), .ZN(n8101) );
  NAND2_X1 U9449 ( .A1(n8101), .A2(n8833), .ZN(n8102) );
  NAND2_X1 U9450 ( .A1(n8103), .A2(n8102), .ZN(n8104) );
  INV_X1 U9451 ( .A(n8104), .ZN(n8106) );
  INV_X1 U9452 ( .A(n8108), .ZN(n8105) );
  INV_X1 U9453 ( .A(n8403), .ZN(n8107) );
  AOI21_X1 U9454 ( .B1(n8108), .B2(n8104), .A(n8107), .ZN(n8117) );
  INV_X1 U9455 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n8109) );
  NOR2_X1 U9456 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8109), .ZN(n10853) );
  NOR2_X1 U9457 ( .A1(n8110), .A2(n8816), .ZN(n8111) );
  AOI211_X1 U9458 ( .C1(n8814), .C2(n8831), .A(n10853), .B(n8111), .ZN(n8112)
         );
  OAI21_X1 U9459 ( .B1(n8113), .B2(n8756), .A(n8112), .ZN(n8114) );
  AOI21_X1 U9460 ( .B1(n8115), .B2(n8805), .A(n8114), .ZN(n8116) );
  OAI21_X1 U9461 ( .B1(n8117), .B2(n8808), .A(n8116), .ZN(P2_U3155) );
  INV_X1 U9462 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n8127) );
  NAND2_X1 U9463 ( .A1(n8118), .A2(n11199), .ZN(n8125) );
  OAI22_X1 U9464 ( .A1(n8178), .A2(n11107), .B1(n8119), .B2(n11109), .ZN(n8120) );
  AOI21_X1 U9465 ( .B1(n8121), .B2(n11147), .A(n8120), .ZN(n8124) );
  NAND4_X1 U9466 ( .A1(n8125), .A2(n8124), .A3(n8123), .A4(n8122), .ZN(n8128)
         );
  NAND2_X1 U9467 ( .A1(n8128), .A2(n11206), .ZN(n8126) );
  OAI21_X1 U9468 ( .B1(n11206), .B2(n8127), .A(n8126), .ZN(P1_U3495) );
  NAND2_X1 U9469 ( .A1(n8128), .A2(n11202), .ZN(n8129) );
  OAI21_X1 U9470 ( .B1(n11202), .B2(n10113), .A(n8129), .ZN(P1_U3536) );
  INV_X1 U9471 ( .A(n9497), .ZN(n8130) );
  INV_X1 U9472 ( .A(n9390), .ZN(n9670) );
  AOI22_X1 U9473 ( .A1(n8131), .A2(n8130), .B1(n9322), .B2(n9670), .ZN(n10192)
         );
  NAND2_X1 U9474 ( .A1(n8132), .A2(n8029), .ZN(n8134) );
  AOI22_X1 U9475 ( .A1(n8215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n8214), .B2(
        n10154), .ZN(n8133) );
  NAND2_X1 U9476 ( .A1(n10488), .A2(n10378), .ZN(n9431) );
  XNOR2_X1 U9477 ( .A(n10192), .B(n10191), .ZN(n10490) );
  INV_X1 U9478 ( .A(n10488), .ZN(n10190) );
  NAND2_X1 U9479 ( .A1(n10190), .A2(n8135), .ZN(n10382) );
  INV_X1 U9480 ( .A(n10382), .ZN(n8136) );
  AOI211_X1 U9481 ( .C1(n10488), .C2(n8137), .A(n11212), .B(n8136), .ZN(n10486) );
  NOR2_X1 U9482 ( .A1(n10190), .A2(n10387), .ZN(n8140) );
  OAI22_X1 U9483 ( .A1(n10358), .A2(n8138), .B1(n9331), .B2(n10968), .ZN(n8139) );
  AOI211_X1 U9484 ( .C1(n10486), .C2(n11128), .A(n8140), .B(n8139), .ZN(n8154)
         );
  NAND2_X1 U9485 ( .A1(n8377), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8148) );
  INV_X1 U9486 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n8141) );
  OR2_X1 U9487 ( .A1(n5143), .A2(n8141), .ZN(n8147) );
  OAI21_X1 U9488 ( .B1(P1_REG3_REG_18__SCAN_IN), .B2(n8143), .A(n8142), .ZN(
        n10383) );
  OR2_X1 U9489 ( .A1(n8382), .A2(n10383), .ZN(n8146) );
  INV_X1 U9490 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n8144) );
  OR2_X1 U9491 ( .A1(n6968), .A2(n8144), .ZN(n8145) );
  NAND2_X1 U9492 ( .A1(n8150), .A2(n10191), .ZN(n9454) );
  OAI211_X1 U9493 ( .C1(n8150), .C2(n10191), .A(n9454), .B(n11181), .ZN(n8152)
         );
  OR2_X1 U9494 ( .A1(n9390), .A2(n11109), .ZN(n8151) );
  OAI211_X1 U9495 ( .C1(n9432), .C2(n11107), .A(n8152), .B(n8151), .ZN(n10487)
         );
  NAND2_X1 U9496 ( .A1(n10487), .A2(n10367), .ZN(n8153) );
  OAI211_X1 U9497 ( .C1(n10490), .C2(n10391), .A(n8154), .B(n8153), .ZN(
        P1_U3276) );
  INV_X1 U9498 ( .A(n8332), .ZN(n8156) );
  OAI222_X1 U9499 ( .A1(n5141), .A2(n9797), .B1(n10517), .B2(n8156), .C1(
        P1_U3086), .C2(n8155), .ZN(P1_U3329) );
  OAI222_X1 U9500 ( .A1(n9267), .A2(n8157), .B1(n9262), .B2(n8156), .C1(n6356), 
        .C2(P2_U3151), .ZN(P2_U3269) );
  MUX2_X1 U9501 ( .A(n8158), .B(P2_REG2_REG_7__SCAN_IN), .S(n9150), .Z(n8166)
         );
  NAND3_X1 U9502 ( .A1(n7477), .A2(n9148), .A3(n8159), .ZN(n8164) );
  NOR2_X1 U9503 ( .A1(n9142), .A2(n8160), .ZN(n8161) );
  AOI21_X1 U9504 ( .B1(n9111), .B2(n8162), .A(n8161), .ZN(n8163) );
  NAND2_X1 U9505 ( .A1(n8164), .A2(n8163), .ZN(n8165) );
  OR2_X1 U9506 ( .A1(n8166), .A2(n8165), .ZN(P2_U3226) );
  INV_X1 U9507 ( .A(n9405), .ZN(n9261) );
  OAI222_X1 U9508 ( .A1(n5141), .A2(n9406), .B1(n10517), .B2(n9261), .C1(n6520), .C2(P1_U3086), .ZN(P1_U3326) );
  NAND2_X1 U9509 ( .A1(n8913), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n8167) );
  OAI21_X1 U9510 ( .B1(n8168), .B2(n8913), .A(n8167), .ZN(P2_U3491) );
  NAND2_X1 U9511 ( .A1(n8172), .A2(n8169), .ZN(n8170) );
  NAND2_X1 U9512 ( .A1(n8171), .A2(n8170), .ZN(n8176) );
  INV_X1 U9513 ( .A(n8172), .ZN(n8174) );
  NAND2_X1 U9514 ( .A1(n8174), .A2(n8173), .ZN(n8175) );
  NOR2_X1 U9515 ( .A1(n8178), .A2(n5144), .ZN(n8177) );
  AOI21_X1 U9516 ( .B1(n9400), .B2(n8349), .A(n8177), .ZN(n9386) );
  NAND2_X1 U9517 ( .A1(n9400), .A2(n8388), .ZN(n8180) );
  OR2_X1 U9518 ( .A1(n8178), .A2(n8390), .ZN(n8179) );
  NAND2_X1 U9519 ( .A1(n8180), .A2(n8179), .ZN(n8181) );
  XNOR2_X1 U9520 ( .A(n8181), .B(n8314), .ZN(n9312) );
  NAND2_X1 U9521 ( .A1(n9322), .A2(n8388), .ZN(n8183) );
  OR2_X1 U9522 ( .A1(n9390), .A2(n8390), .ZN(n8182) );
  NAND2_X1 U9523 ( .A1(n8183), .A2(n8182), .ZN(n8184) );
  XNOR2_X1 U9524 ( .A(n8184), .B(n8346), .ZN(n8187) );
  NAND2_X1 U9525 ( .A1(n9322), .A2(n8349), .ZN(n8186) );
  OR2_X1 U9526 ( .A1(n9390), .A2(n5144), .ZN(n8185) );
  NAND2_X1 U9527 ( .A1(n8186), .A2(n8185), .ZN(n8188) );
  NAND2_X1 U9528 ( .A1(n8187), .A2(n8188), .ZN(n9311) );
  OAI21_X1 U9529 ( .B1(n9386), .B2(n9312), .A(n9311), .ZN(n8193) );
  NAND3_X1 U9530 ( .A1(n9311), .A2(n9386), .A3(n9312), .ZN(n8191) );
  INV_X1 U9531 ( .A(n8187), .ZN(n8190) );
  INV_X1 U9532 ( .A(n8188), .ZN(n8189) );
  NAND2_X1 U9533 ( .A1(n8190), .A2(n8189), .ZN(n9310) );
  AND2_X1 U9534 ( .A1(n8191), .A2(n9310), .ZN(n8192) );
  NAND2_X1 U9535 ( .A1(n10488), .A2(n8388), .ZN(n8195) );
  OR2_X1 U9536 ( .A1(n10378), .A2(n8390), .ZN(n8194) );
  NAND2_X1 U9537 ( .A1(n8195), .A2(n8194), .ZN(n8196) );
  XNOR2_X1 U9538 ( .A(n8196), .B(n8346), .ZN(n8199) );
  NAND2_X1 U9539 ( .A1(n10488), .A2(n8349), .ZN(n8198) );
  OR2_X1 U9540 ( .A1(n10378), .A2(n5144), .ZN(n8197) );
  NAND2_X1 U9541 ( .A1(n8198), .A2(n8197), .ZN(n8200) );
  NAND2_X1 U9542 ( .A1(n8199), .A2(n8200), .ZN(n9327) );
  INV_X1 U9543 ( .A(n8199), .ZN(n8202) );
  INV_X1 U9544 ( .A(n8200), .ZN(n8201) );
  NAND2_X1 U9545 ( .A1(n8202), .A2(n8201), .ZN(n9326) );
  NAND2_X1 U9546 ( .A1(n8203), .A2(n8029), .ZN(n8205) );
  AOI22_X1 U9547 ( .A1(n8215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n8214), .B2(
        n10730), .ZN(n8204) );
  NAND2_X1 U9548 ( .A1(n10483), .A2(n8388), .ZN(n8207) );
  OR2_X1 U9549 ( .A1(n9432), .A2(n8390), .ZN(n8206) );
  NAND2_X1 U9550 ( .A1(n8207), .A2(n8206), .ZN(n8208) );
  XNOR2_X1 U9551 ( .A(n8208), .B(n8314), .ZN(n8210) );
  NOR2_X1 U9552 ( .A1(n9432), .A2(n5144), .ZN(n8209) );
  AOI21_X1 U9553 ( .B1(n10483), .B2(n8349), .A(n8209), .ZN(n9365) );
  NAND2_X1 U9554 ( .A1(n8211), .A2(n8210), .ZN(n9363) );
  NAND2_X1 U9555 ( .A1(n8212), .A2(n9363), .ZN(n9285) );
  NAND2_X1 U9556 ( .A1(n8213), .A2(n8029), .ZN(n8217) );
  AOI22_X1 U9557 ( .A1(n8215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n10158), 
        .B2(n8214), .ZN(n8216) );
  NAND2_X1 U9558 ( .A1(n10478), .A2(n8388), .ZN(n8225) );
  NAND2_X1 U9559 ( .A1(n8377), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8223) );
  INV_X1 U9560 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n10157) );
  OR2_X1 U9561 ( .A1(n6968), .A2(n10157), .ZN(n8222) );
  OAI21_X1 U9562 ( .B1(P1_REG3_REG_19__SCAN_IN), .B2(n8219), .A(n8218), .ZN(
        n10356) );
  OR2_X1 U9563 ( .A1(n8382), .A2(n10356), .ZN(n8221) );
  INV_X1 U9564 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n10357) );
  OR2_X1 U9565 ( .A1(n5143), .A2(n10357), .ZN(n8220) );
  OR2_X1 U9566 ( .A1(n10349), .A2(n8390), .ZN(n8224) );
  NAND2_X1 U9567 ( .A1(n8225), .A2(n8224), .ZN(n8226) );
  XNOR2_X1 U9568 ( .A(n8226), .B(n8346), .ZN(n8228) );
  NOR2_X1 U9569 ( .A1(n10349), .A2(n5144), .ZN(n8227) );
  AOI21_X1 U9570 ( .B1(n10478), .B2(n8349), .A(n8227), .ZN(n8229) );
  XNOR2_X1 U9571 ( .A(n8228), .B(n8229), .ZN(n9286) );
  NAND2_X1 U9572 ( .A1(n9285), .A2(n9286), .ZN(n8232) );
  INV_X1 U9573 ( .A(n8228), .ZN(n8230) );
  NAND2_X1 U9574 ( .A1(n8230), .A2(n8229), .ZN(n8231) );
  NAND2_X1 U9575 ( .A1(n8233), .A2(n8029), .ZN(n8235) );
  OR2_X1 U9576 ( .A1(n5138), .A2(n10021), .ZN(n8234) );
  NAND2_X1 U9577 ( .A1(n8377), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8242) );
  INV_X1 U9578 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8236) );
  OR2_X1 U9579 ( .A1(n6968), .A2(n8236), .ZN(n8241) );
  INV_X1 U9580 ( .A(n8237), .ZN(n8257) );
  OAI21_X1 U9581 ( .B1(P1_REG3_REG_20__SCAN_IN), .B2(n8238), .A(n8257), .ZN(
        n10342) );
  OR2_X1 U9582 ( .A1(n8382), .A2(n10342), .ZN(n8240) );
  INV_X1 U9583 ( .A(P1_REG2_REG_20__SCAN_IN), .ZN(n10343) );
  OR2_X1 U9584 ( .A1(n5143), .A2(n10343), .ZN(n8239) );
  NAND4_X1 U9585 ( .A1(n8242), .A2(n8241), .A3(n8240), .A4(n8239), .ZN(n10462)
         );
  INV_X1 U9586 ( .A(n10462), .ZN(n9435) );
  OAI22_X1 U9587 ( .A1(n10341), .A2(n8330), .B1(n9435), .B2(n8390), .ZN(n8243)
         );
  XNOR2_X1 U9588 ( .A(n8243), .B(n8314), .ZN(n8248) );
  OR2_X1 U9589 ( .A1(n10341), .A2(n8390), .ZN(n8245) );
  NAND2_X1 U9590 ( .A1(n10462), .A2(n8264), .ZN(n8244) );
  NAND2_X1 U9591 ( .A1(n8245), .A2(n8244), .ZN(n8246) );
  XNOR2_X1 U9592 ( .A(n8248), .B(n8246), .ZN(n9344) );
  INV_X1 U9593 ( .A(n8246), .ZN(n8247) );
  NAND2_X1 U9594 ( .A1(n8248), .A2(n8247), .ZN(n8249) );
  NAND2_X1 U9595 ( .A1(n8250), .A2(n8029), .ZN(n8253) );
  OR2_X1 U9596 ( .A1(n5139), .A2(n8251), .ZN(n8252) );
  NAND2_X1 U9597 ( .A1(n8357), .A2(P1_REG1_REG_21__SCAN_IN), .ZN(n8262) );
  INV_X1 U9598 ( .A(P1_REG0_REG_21__SCAN_IN), .ZN(n8254) );
  OR2_X1 U9599 ( .A1(n6966), .A2(n8254), .ZN(n8261) );
  INV_X1 U9600 ( .A(n8255), .ZN(n8277) );
  INV_X1 U9601 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n8256) );
  NAND2_X1 U9602 ( .A1(n8257), .A2(n8256), .ZN(n8258) );
  NAND2_X1 U9603 ( .A1(n8277), .A2(n8258), .ZN(n10323) );
  OR2_X1 U9604 ( .A1(n8382), .A2(n10323), .ZN(n8260) );
  INV_X1 U9605 ( .A(P1_REG2_REG_21__SCAN_IN), .ZN(n10324) );
  OR2_X1 U9606 ( .A1(n5143), .A2(n10324), .ZN(n8259) );
  NAND4_X1 U9607 ( .A1(n8262), .A2(n8261), .A3(n8260), .A4(n8259), .ZN(n10454)
         );
  OAI22_X1 U9608 ( .A1(n10466), .A2(n8330), .B1(n10350), .B2(n8390), .ZN(n8263) );
  XNOR2_X1 U9609 ( .A(n8263), .B(n8346), .ZN(n8267) );
  OR2_X1 U9610 ( .A1(n10466), .A2(n8390), .ZN(n8266) );
  NAND2_X1 U9611 ( .A1(n10454), .A2(n8264), .ZN(n8265) );
  NAND2_X1 U9612 ( .A1(n8266), .A2(n8265), .ZN(n8268) );
  NAND2_X1 U9613 ( .A1(n8267), .A2(n8268), .ZN(n8288) );
  INV_X1 U9614 ( .A(n8267), .ZN(n8270) );
  INV_X1 U9615 ( .A(n8268), .ZN(n8269) );
  NAND2_X1 U9616 ( .A1(n8270), .A2(n8269), .ZN(n8271) );
  NAND2_X1 U9617 ( .A1(n8288), .A2(n8271), .ZN(n9296) );
  NAND2_X1 U9618 ( .A1(n8272), .A2(n8029), .ZN(n8274) );
  OR2_X1 U9619 ( .A1(n5138), .A2(n9805), .ZN(n8273) );
  NAND2_X1 U9620 ( .A1(n10306), .A2(n8388), .ZN(n8285) );
  NAND2_X1 U9621 ( .A1(n8377), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n8283) );
  INV_X1 U9622 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n8275) );
  OR2_X1 U9623 ( .A1(n6968), .A2(n8275), .ZN(n8282) );
  INV_X1 U9624 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8276) );
  NAND2_X1 U9625 ( .A1(n8277), .A2(n8276), .ZN(n8278) );
  NAND2_X1 U9626 ( .A1(n8279), .A2(n8278), .ZN(n10310) );
  OR2_X1 U9627 ( .A1(n8382), .A2(n10310), .ZN(n8281) );
  INV_X1 U9628 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n10311) );
  OR2_X1 U9629 ( .A1(n5143), .A2(n10311), .ZN(n8280) );
  OR2_X1 U9630 ( .A1(n10329), .A2(n8390), .ZN(n8284) );
  NAND2_X1 U9631 ( .A1(n8285), .A2(n8284), .ZN(n8286) );
  XNOR2_X1 U9632 ( .A(n8286), .B(n8314), .ZN(n8289) );
  AND2_X1 U9633 ( .A1(n8288), .A2(n8289), .ZN(n8287) );
  INV_X1 U9634 ( .A(n10306), .ZN(n10456) );
  OAI22_X1 U9635 ( .A1(n10456), .A2(n8390), .B1(n10329), .B2(n5144), .ZN(n9354) );
  NAND2_X1 U9636 ( .A1(n9356), .A2(n9354), .ZN(n9351) );
  NAND2_X1 U9637 ( .A1(n9294), .A2(n8288), .ZN(n8291) );
  INV_X1 U9638 ( .A(n8289), .ZN(n8290) );
  NAND2_X1 U9639 ( .A1(n8292), .A2(n8029), .ZN(n8294) );
  OR2_X1 U9640 ( .A1(n5138), .A2(n10017), .ZN(n8293) );
  OAI22_X1 U9641 ( .A1(n10448), .A2(n8330), .B1(n10312), .B2(n8390), .ZN(n8295) );
  XNOR2_X1 U9642 ( .A(n8295), .B(n8346), .ZN(n8296) );
  OAI22_X1 U9643 ( .A1(n10448), .A2(n8390), .B1(n10312), .B2(n5144), .ZN(n8297) );
  XNOR2_X1 U9644 ( .A(n8296), .B(n8297), .ZN(n9279) );
  INV_X1 U9645 ( .A(n8296), .ZN(n8299) );
  INV_X1 U9646 ( .A(n8297), .ZN(n8298) );
  NAND2_X1 U9647 ( .A1(n8300), .A2(n8029), .ZN(n8302) );
  OR2_X1 U9648 ( .A1(n5139), .A2(n9801), .ZN(n8301) );
  NAND2_X1 U9649 ( .A1(n10442), .A2(n8388), .ZN(n8313) );
  NAND2_X1 U9650 ( .A1(n8357), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8311) );
  INV_X1 U9651 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n8303) );
  OR2_X1 U9652 ( .A1(n6966), .A2(n8303), .ZN(n8310) );
  INV_X1 U9653 ( .A(n8304), .ZN(n8323) );
  INV_X1 U9654 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8305) );
  NAND2_X1 U9655 ( .A1(n8306), .A2(n8305), .ZN(n8307) );
  NAND2_X1 U9656 ( .A1(n8323), .A2(n8307), .ZN(n10278) );
  OR2_X1 U9657 ( .A1(n8382), .A2(n10278), .ZN(n8309) );
  INV_X1 U9658 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n10279) );
  OR2_X1 U9659 ( .A1(n5143), .A2(n10279), .ZN(n8308) );
  OR2_X1 U9660 ( .A1(n10297), .A2(n8390), .ZN(n8312) );
  NAND2_X1 U9661 ( .A1(n8313), .A2(n8312), .ZN(n8315) );
  XNOR2_X1 U9662 ( .A(n8315), .B(n8314), .ZN(n8318) );
  NOR2_X1 U9663 ( .A1(n10297), .A2(n5144), .ZN(n8316) );
  AOI21_X1 U9664 ( .B1(n10442), .B2(n8349), .A(n8316), .ZN(n8317) );
  NOR2_X1 U9665 ( .A1(n8318), .A2(n8317), .ZN(n9337) );
  NAND2_X1 U9666 ( .A1(n8318), .A2(n8317), .ZN(n9335) );
  NAND2_X1 U9667 ( .A1(n8377), .A2(P1_REG0_REG_25__SCAN_IN), .ZN(n8329) );
  INV_X1 U9668 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n8320) );
  OR2_X1 U9669 ( .A1(n6968), .A2(n8320), .ZN(n8328) );
  INV_X1 U9670 ( .A(n8321), .ZN(n8338) );
  INV_X1 U9671 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8322) );
  NAND2_X1 U9672 ( .A1(n8323), .A2(n8322), .ZN(n8324) );
  NAND2_X1 U9673 ( .A1(n8338), .A2(n8324), .ZN(n9305) );
  OR2_X1 U9674 ( .A1(n8382), .A2(n9305), .ZN(n8327) );
  INV_X1 U9675 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n8325) );
  OR2_X1 U9676 ( .A1(n5143), .A2(n8325), .ZN(n8326) );
  NAND4_X1 U9677 ( .A1(n8329), .A2(n8328), .A3(n8327), .A4(n8326), .ZN(n10424)
         );
  OAI22_X1 U9678 ( .A1(n10435), .A2(n8390), .B1(n10196), .B2(n5144), .ZN(n8351) );
  OAI22_X1 U9679 ( .A1(n10435), .A2(n8330), .B1(n10196), .B2(n8390), .ZN(n8331) );
  XNOR2_X1 U9680 ( .A(n8331), .B(n8346), .ZN(n8350) );
  XOR2_X1 U9681 ( .A(n8351), .B(n8350), .Z(n9303) );
  NAND2_X1 U9682 ( .A1(n8332), .A2(n8029), .ZN(n8334) );
  OR2_X1 U9683 ( .A1(n5139), .A2(n9797), .ZN(n8333) );
  NAND2_X1 U9684 ( .A1(n10257), .A2(n8388), .ZN(n8345) );
  NAND2_X1 U9685 ( .A1(n8377), .A2(P1_REG0_REG_26__SCAN_IN), .ZN(n8343) );
  INV_X1 U9686 ( .A(P1_REG1_REG_26__SCAN_IN), .ZN(n8335) );
  OR2_X1 U9687 ( .A1(n6968), .A2(n8335), .ZN(n8342) );
  INV_X1 U9688 ( .A(n8336), .ZN(n8361) );
  INV_X1 U9689 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8337) );
  NAND2_X1 U9690 ( .A1(n8338), .A2(n8337), .ZN(n8339) );
  NAND2_X1 U9691 ( .A1(n8361), .A2(n8339), .ZN(n10252) );
  OR2_X1 U9692 ( .A1(n8382), .A2(n10252), .ZN(n8341) );
  INV_X1 U9693 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n10253) );
  OR2_X1 U9694 ( .A1(n5143), .A2(n10253), .ZN(n8340) );
  OR2_X1 U9695 ( .A1(n10269), .A2(n8390), .ZN(n8344) );
  NAND2_X1 U9696 ( .A1(n8345), .A2(n8344), .ZN(n8347) );
  XNOR2_X1 U9697 ( .A(n8347), .B(n8346), .ZN(n8371) );
  NOR2_X1 U9698 ( .A1(n10269), .A2(n5144), .ZN(n8348) );
  AOI21_X1 U9699 ( .B1(n10257), .B2(n8349), .A(n8348), .ZN(n8372) );
  XNOR2_X1 U9700 ( .A(n8371), .B(n8372), .ZN(n9377) );
  INV_X1 U9701 ( .A(n8350), .ZN(n8353) );
  INV_X1 U9702 ( .A(n8351), .ZN(n8352) );
  NAND2_X1 U9703 ( .A1(n8353), .A2(n8352), .ZN(n9374) );
  NAND2_X1 U9704 ( .A1(n8448), .A2(n8029), .ZN(n8356) );
  NAND2_X1 U9705 ( .A1(n8357), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8367) );
  INV_X1 U9706 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n8358) );
  OR2_X1 U9707 ( .A1(n6966), .A2(n8358), .ZN(n8366) );
  INV_X1 U9708 ( .A(n8359), .ZN(n8380) );
  INV_X1 U9709 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8360) );
  NAND2_X1 U9710 ( .A1(n8361), .A2(n8360), .ZN(n8362) );
  NAND2_X1 U9711 ( .A1(n8380), .A2(n8362), .ZN(n9272) );
  OR2_X1 U9712 ( .A1(n8382), .A2(n9272), .ZN(n8365) );
  INV_X1 U9713 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n8363) );
  OR2_X1 U9714 ( .A1(n5143), .A2(n8363), .ZN(n8364) );
  INV_X1 U9715 ( .A(n10409), .ZN(n10425) );
  AOI22_X1 U9716 ( .A1(n10244), .A2(n8388), .B1(n8349), .B2(n10425), .ZN(n8368) );
  XOR2_X1 U9717 ( .A(n8346), .B(n8368), .Z(n8370) );
  OAI22_X1 U9718 ( .A1(n10419), .A2(n8390), .B1(n10409), .B2(n5144), .ZN(n8369) );
  NOR2_X1 U9719 ( .A1(n8370), .A2(n8369), .ZN(n8374) );
  AOI21_X1 U9720 ( .B1(n8370), .B2(n8369), .A(n8374), .ZN(n9269) );
  INV_X1 U9721 ( .A(n8371), .ZN(n8373) );
  OR2_X1 U9722 ( .A1(n8373), .A2(n8372), .ZN(n9270) );
  NAND2_X1 U9723 ( .A1(n10519), .A2(n8029), .ZN(n8376) );
  INV_X1 U9724 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n10521) );
  OR2_X1 U9725 ( .A1(n5139), .A2(n10521), .ZN(n8375) );
  NAND2_X1 U9726 ( .A1(n8377), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n8386) );
  INV_X1 U9727 ( .A(P1_REG1_REG_28__SCAN_IN), .ZN(n8378) );
  OR2_X1 U9728 ( .A1(n6968), .A2(n8378), .ZN(n8385) );
  INV_X1 U9729 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n8379) );
  NAND2_X1 U9730 ( .A1(n8380), .A2(n8379), .ZN(n8381) );
  NAND2_X1 U9731 ( .A1(n10209), .A2(n8381), .ZN(n10225) );
  OR2_X1 U9732 ( .A1(n8382), .A2(n10225), .ZN(n8384) );
  INV_X1 U9733 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n10226) );
  OR2_X1 U9734 ( .A1(n5143), .A2(n10226), .ZN(n8383) );
  INV_X1 U9735 ( .A(n10401), .ZN(n10416) );
  AOI22_X1 U9736 ( .A1(n10412), .A2(n8388), .B1(n8349), .B2(n10416), .ZN(n8393) );
  INV_X1 U9737 ( .A(n10412), .ZN(n10201) );
  OAI22_X1 U9738 ( .A1(n10201), .A2(n8390), .B1(n10401), .B2(n5144), .ZN(n8391) );
  XNOR2_X1 U9739 ( .A(n8391), .B(n8346), .ZN(n8392) );
  XOR2_X1 U9740 ( .A(n8393), .B(n8392), .Z(n8394) );
  NOR2_X1 U9741 ( .A1(n9397), .A2(n10225), .ZN(n8397) );
  AOI22_X1 U9742 ( .A1(n9394), .A2(n10425), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3086), .ZN(n8395) );
  OAI21_X1 U9743 ( .B1(n10408), .B2(n9391), .A(n8395), .ZN(n8396) );
  AOI211_X1 U9744 ( .C1(n10412), .C2(n9399), .A(n8397), .B(n8396), .ZN(n8398)
         );
  OAI21_X1 U9745 ( .B1(n8399), .B2(n9402), .A(n8398), .ZN(P1_U3220) );
  INV_X1 U9746 ( .A(n8400), .ZN(n8401) );
  NAND2_X1 U9747 ( .A1(n8401), .A2(n8817), .ZN(n8402) );
  XNOR2_X1 U9748 ( .A(n8404), .B(n8440), .ZN(n8405) );
  XNOR2_X1 U9749 ( .A(n8405), .B(n8831), .ZN(n8812) );
  INV_X1 U9750 ( .A(n8405), .ZN(n8406) );
  NAND2_X1 U9751 ( .A1(n8406), .A2(n8831), .ZN(n8407) );
  XNOR2_X1 U9752 ( .A(n8739), .B(n8440), .ZN(n8409) );
  XNOR2_X1 U9753 ( .A(n8409), .B(n9135), .ZN(n8743) );
  NAND2_X1 U9754 ( .A1(n8740), .A2(n8743), .ZN(n8741) );
  NAND2_X1 U9755 ( .A1(n8409), .A2(n8408), .ZN(n8410) );
  NAND2_X1 U9756 ( .A1(n8741), .A2(n8410), .ZN(n8750) );
  XNOR2_X1 U9757 ( .A(n8758), .B(n8424), .ZN(n8751) );
  NAND2_X1 U9758 ( .A1(n8751), .A2(n8830), .ZN(n8411) );
  NAND2_X1 U9759 ( .A1(n8750), .A2(n8411), .ZN(n8788) );
  XNOR2_X1 U9760 ( .A(n8786), .B(n8424), .ZN(n8415) );
  XNOR2_X1 U9761 ( .A(n8415), .B(n9134), .ZN(n8789) );
  INV_X1 U9762 ( .A(n8789), .ZN(n8413) );
  INV_X1 U9763 ( .A(n8751), .ZN(n8412) );
  NAND2_X1 U9764 ( .A1(n8412), .A2(n9118), .ZN(n8787) );
  AND2_X1 U9765 ( .A1(n8413), .A2(n8787), .ZN(n8414) );
  NAND2_X1 U9766 ( .A1(n8788), .A2(n8414), .ZN(n8791) );
  NAND2_X1 U9767 ( .A1(n8415), .A2(n9134), .ZN(n8416) );
  NAND2_X1 U9768 ( .A1(n8791), .A2(n8416), .ZN(n8716) );
  XNOR2_X1 U9769 ( .A(n8417), .B(n8424), .ZN(n8715) );
  INV_X1 U9770 ( .A(n8715), .ZN(n8418) );
  NAND2_X1 U9771 ( .A1(n8418), .A2(n8829), .ZN(n8419) );
  XNOR2_X1 U9772 ( .A(n8768), .B(n8440), .ZN(n8420) );
  XNOR2_X1 U9773 ( .A(n8420), .B(n9104), .ZN(n8770) );
  XNOR2_X1 U9774 ( .A(n9179), .B(n8440), .ZN(n8421) );
  XNOR2_X1 U9775 ( .A(n8421), .B(n9064), .ZN(n8724) );
  NAND2_X1 U9776 ( .A1(n8722), .A2(n8724), .ZN(n8423) );
  NAND2_X1 U9777 ( .A1(n8421), .A2(n9091), .ZN(n8422) );
  NAND2_X1 U9778 ( .A1(n8423), .A2(n8422), .ZN(n8777) );
  INV_X1 U9779 ( .A(n8777), .ZN(n8426) );
  XNOR2_X1 U9780 ( .A(n9175), .B(n8424), .ZN(n8427) );
  XNOR2_X1 U9781 ( .A(n8427), .B(n9075), .ZN(n8778) );
  INV_X1 U9782 ( .A(n8778), .ZN(n8425) );
  NAND2_X1 U9783 ( .A1(n8427), .A2(n9075), .ZN(n8428) );
  XNOR2_X1 U9784 ( .A(n9174), .B(n8440), .ZN(n8429) );
  XNOR2_X1 U9785 ( .A(n9039), .B(n8440), .ZN(n8431) );
  XNOR2_X1 U9786 ( .A(n8431), .B(n9054), .ZN(n8762) );
  XNOR2_X1 U9787 ( .A(n9162), .B(n8440), .ZN(n8433) );
  XNOR2_X1 U9788 ( .A(n8806), .B(n8440), .ZN(n8434) );
  XNOR2_X1 U9789 ( .A(n8434), .B(n9025), .ZN(n8799) );
  XNOR2_X1 U9790 ( .A(n9155), .B(n8440), .ZN(n8436) );
  NOR2_X1 U9791 ( .A1(n8436), .A2(n9015), .ZN(n8437) );
  AOI21_X1 U9792 ( .B1(n9015), .B2(n8436), .A(n8437), .ZN(n8702) );
  INV_X1 U9793 ( .A(n8437), .ZN(n8438) );
  NAND2_X1 U9794 ( .A1(n8701), .A2(n8438), .ZN(n8442) );
  XOR2_X1 U9795 ( .A(n8440), .B(n8439), .Z(n8441) );
  XNOR2_X1 U9796 ( .A(n8442), .B(n8441), .ZN(n8447) );
  NAND2_X1 U9797 ( .A1(n8826), .A2(n8814), .ZN(n8444) );
  AOI22_X1 U9798 ( .A1(n8991), .A2(n8819), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3151), .ZN(n8443) );
  OAI211_X1 U9799 ( .C1(n9015), .C2(n8816), .A(n8444), .B(n8443), .ZN(n8445)
         );
  AOI21_X1 U9800 ( .B1(n8665), .B2(n8805), .A(n8445), .ZN(n8446) );
  OAI21_X1 U9801 ( .B1(n8447), .B2(n8808), .A(n8446), .ZN(P2_U3160) );
  INV_X1 U9802 ( .A(n8448), .ZN(n10523) );
  OAI222_X1 U9803 ( .A1(n9267), .A2(n8449), .B1(n9262), .B2(n10523), .C1(n6588), .C2(P2_U3151), .ZN(P2_U3268) );
  INV_X1 U9804 ( .A(SI_29_), .ZN(n9687) );
  INV_X1 U9805 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10515) );
  MUX2_X1 U9806 ( .A(n10515), .B(n8698), .S(n5134), .Z(n8454) );
  INV_X1 U9807 ( .A(SI_30_), .ZN(n9889) );
  NAND2_X1 U9808 ( .A1(n8454), .A2(n9889), .ZN(n8457) );
  INV_X1 U9809 ( .A(n8454), .ZN(n8455) );
  NAND2_X1 U9810 ( .A1(n8455), .A2(SI_30_), .ZN(n8456) );
  NAND2_X1 U9811 ( .A1(n8457), .A2(n8456), .ZN(n8464) );
  MUX2_X1 U9812 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n5134), .Z(n8459) );
  INV_X1 U9813 ( .A(SI_31_), .ZN(n8458) );
  XNOR2_X1 U9814 ( .A(n8459), .B(n8458), .ZN(n8460) );
  NAND2_X1 U9815 ( .A1(n9452), .A2(n8468), .ZN(n8463) );
  OR2_X1 U9816 ( .A1(n5926), .A2(n6553), .ZN(n8462) );
  NOR2_X1 U9817 ( .A1(n8689), .A2(n8977), .ZN(n8672) );
  NAND2_X1 U9818 ( .A1(n8465), .A2(n8464), .ZN(n8466) );
  NAND2_X1 U9819 ( .A1(n9446), .A2(n8468), .ZN(n8470) );
  OR2_X1 U9820 ( .A1(n5926), .A2(n8698), .ZN(n8469) );
  INV_X1 U9821 ( .A(n8825), .ZN(n8674) );
  NAND2_X1 U9822 ( .A1(n8675), .A2(n8674), .ZN(n8504) );
  INV_X1 U9823 ( .A(n8471), .ZN(n9004) );
  NAND2_X1 U9824 ( .A1(n8651), .A2(n8652), .ZN(n9023) );
  INV_X1 U9825 ( .A(n8472), .ZN(n8643) );
  NAND2_X1 U9826 ( .A1(n8643), .A2(n8642), .ZN(n8640) );
  INV_X1 U9827 ( .A(n8473), .ZN(n8475) );
  NAND3_X1 U9828 ( .A1(n8475), .A2(n8474), .A3(n8545), .ZN(n8479) );
  NAND2_X1 U9829 ( .A1(n8477), .A2(n8476), .ZN(n8478) );
  NOR2_X1 U9830 ( .A1(n8479), .A2(n8478), .ZN(n8482) );
  AND2_X1 U9831 ( .A1(n8480), .A2(n8529), .ZN(n8481) );
  NAND4_X1 U9832 ( .A1(n8482), .A2(n6030), .A3(n8481), .A4(n8560), .ZN(n8483)
         );
  NOR2_X1 U9833 ( .A1(n8483), .A2(n8514), .ZN(n8485) );
  NAND4_X1 U9834 ( .A1(n5511), .A2(n8486), .A3(n8485), .A4(n8484), .ZN(n8487)
         );
  NOR2_X1 U9835 ( .A1(n8589), .A2(n8487), .ZN(n8488) );
  NAND4_X1 U9836 ( .A1(n8489), .A2(n6330), .A3(n8488), .A4(n8594), .ZN(n8490)
         );
  NOR3_X1 U9837 ( .A1(n9123), .A2(n9140), .A3(n8490), .ZN(n8491) );
  NAND3_X1 U9838 ( .A1(n9093), .A2(n9102), .A3(n8491), .ZN(n8492) );
  NOR2_X1 U9839 ( .A1(n8640), .A2(n8492), .ZN(n8493) );
  NAND3_X1 U9840 ( .A1(n9058), .A2(n8493), .A3(n5435), .ZN(n8494) );
  NOR4_X1 U9841 ( .A1(n9016), .A2(n9041), .A3(n9023), .A4(n8494), .ZN(n8495)
         );
  NAND4_X1 U9842 ( .A1(n8504), .A2(n8496), .A3(n8998), .A4(n8495), .ZN(n8497)
         );
  NOR4_X2 U9843 ( .A1(n8672), .A2(n8677), .A3(n8497), .A4(n8669), .ZN(n8498)
         );
  NAND2_X1 U9844 ( .A1(n8498), .A2(n5140), .ZN(n8512) );
  NAND3_X1 U9845 ( .A1(n9017), .A2(n8500), .A3(n8499), .ZN(n8503) );
  AND2_X1 U9846 ( .A1(n8501), .A2(n8679), .ZN(n8502) );
  NAND2_X1 U9847 ( .A1(n8503), .A2(n8502), .ZN(n8505) );
  NAND3_X1 U9848 ( .A1(n8505), .A2(n8671), .A3(n8504), .ZN(n8510) );
  NAND2_X1 U9849 ( .A1(n8512), .A2(n8511), .ZN(n8687) );
  INV_X1 U9850 ( .A(n8673), .ZN(n8686) );
  INV_X1 U9851 ( .A(n8518), .ZN(n8513) );
  NAND2_X1 U9852 ( .A1(n8516), .A2(n8515), .ZN(n8517) );
  OAI21_X1 U9853 ( .B1(n8519), .B2(n8839), .A(n8518), .ZN(n8520) );
  NAND2_X1 U9854 ( .A1(n8521), .A2(n8520), .ZN(n8523) );
  NAND3_X1 U9855 ( .A1(n8523), .A2(n8522), .A3(n8574), .ZN(n8524) );
  NAND2_X1 U9856 ( .A1(n8524), .A2(n8663), .ZN(n8567) );
  NAND2_X1 U9857 ( .A1(n8526), .A2(n5140), .ZN(n8527) );
  NAND3_X1 U9858 ( .A1(n8527), .A2(n8534), .A3(n8535), .ZN(n8528) );
  NAND2_X1 U9859 ( .A1(n8528), .A2(n8537), .ZN(n8530) );
  NAND2_X1 U9860 ( .A1(n8530), .A2(n8529), .ZN(n8533) );
  AND2_X1 U9861 ( .A1(n8547), .A2(n8531), .ZN(n8532) );
  NAND2_X1 U9862 ( .A1(n8533), .A2(n8532), .ZN(n8544) );
  INV_X1 U9863 ( .A(n8534), .ZN(n8538) );
  INV_X1 U9864 ( .A(n8535), .ZN(n8536) );
  AOI21_X1 U9865 ( .B1(n8538), .B2(n8537), .A(n8536), .ZN(n8542) );
  NAND2_X1 U9866 ( .A1(n8844), .A2(n8539), .ZN(n8540) );
  OAI211_X1 U9867 ( .C1(n8542), .C2(n8541), .A(n8555), .B(n8540), .ZN(n8543)
         );
  MUX2_X1 U9868 ( .A(n8544), .B(n8543), .S(n8663), .Z(n8546) );
  NAND2_X1 U9869 ( .A1(n8546), .A2(n8545), .ZN(n8551) );
  INV_X1 U9870 ( .A(n8547), .ZN(n8549) );
  OAI211_X1 U9871 ( .C1(n8551), .C2(n8549), .A(n8559), .B(n8548), .ZN(n8550)
         );
  NAND3_X1 U9872 ( .A1(n8550), .A2(n8553), .A3(n8568), .ZN(n8558) );
  INV_X1 U9873 ( .A(n8551), .ZN(n8556) );
  NAND2_X1 U9874 ( .A1(n8553), .A2(n8552), .ZN(n8554) );
  AOI21_X1 U9875 ( .B1(n8556), .B2(n8555), .A(n8554), .ZN(n8557) );
  MUX2_X1 U9876 ( .A(n8558), .B(n8557), .S(n8676), .Z(n8565) );
  AOI21_X1 U9877 ( .B1(n8559), .B2(n8561), .A(n8663), .ZN(n8564) );
  OAI21_X1 U9878 ( .B1(n8676), .B2(n8561), .A(n8560), .ZN(n8562) );
  NOR2_X1 U9879 ( .A1(n8572), .A2(n8562), .ZN(n8563) );
  OAI21_X1 U9880 ( .B1(n8565), .B2(n8564), .A(n8563), .ZN(n8566) );
  NAND2_X1 U9881 ( .A1(n8567), .A2(n8566), .ZN(n8570) );
  OR2_X1 U9882 ( .A1(n8568), .A2(n8663), .ZN(n8569) );
  NAND2_X1 U9883 ( .A1(n8570), .A2(n8569), .ZN(n8577) );
  OAI211_X1 U9884 ( .C1(n8573), .C2(n8572), .A(n8577), .B(n8571), .ZN(n8576)
         );
  AND2_X1 U9885 ( .A1(n8580), .A2(n8574), .ZN(n8575) );
  INV_X1 U9886 ( .A(n8577), .ZN(n8583) );
  AND2_X1 U9887 ( .A1(n8579), .A2(n8578), .ZN(n8582) );
  INV_X1 U9888 ( .A(n8580), .ZN(n8581) );
  AOI21_X1 U9889 ( .B1(n8583), .B2(n8582), .A(n8581), .ZN(n8584) );
  MUX2_X1 U9890 ( .A(n8586), .B(n8585), .S(n8676), .Z(n8587) );
  INV_X1 U9891 ( .A(n8587), .ZN(n8588) );
  NOR2_X1 U9892 ( .A1(n8589), .A2(n8588), .ZN(n8593) );
  MUX2_X1 U9893 ( .A(n8591), .B(n8590), .S(n8676), .Z(n8592) );
  NAND2_X1 U9894 ( .A1(n8605), .A2(n8594), .ZN(n8602) );
  AND2_X1 U9895 ( .A1(n8599), .A2(n8595), .ZN(n8597) );
  INV_X1 U9896 ( .A(n8598), .ZN(n8596) );
  AOI21_X1 U9897 ( .B1(n8602), .B2(n8597), .A(n8596), .ZN(n8604) );
  AND2_X1 U9898 ( .A1(n8598), .A2(n8817), .ZN(n8601) );
  INV_X1 U9899 ( .A(n8599), .ZN(n8600) );
  AOI21_X1 U9900 ( .B1(n8602), .B2(n8601), .A(n8600), .ZN(n8603) );
  INV_X1 U9901 ( .A(n8605), .ZN(n8610) );
  NOR2_X1 U9902 ( .A1(n8607), .A2(n8606), .ZN(n8609) );
  AOI21_X1 U9903 ( .B1(n8610), .B2(n8609), .A(n8608), .ZN(n8615) );
  MUX2_X1 U9904 ( .A(n8612), .B(n8611), .S(n8663), .Z(n8613) );
  INV_X1 U9905 ( .A(n8613), .ZN(n8614) );
  MUX2_X1 U9906 ( .A(n9118), .B(n9246), .S(n8676), .Z(n8625) );
  NAND2_X1 U9907 ( .A1(n8624), .A2(n8625), .ZN(n8619) );
  NAND3_X1 U9908 ( .A1(n8619), .A2(n9118), .A3(n8620), .ZN(n8617) );
  NAND2_X1 U9909 ( .A1(n8617), .A2(n8618), .ZN(n8623) );
  NAND3_X1 U9910 ( .A1(n8619), .A2(n9246), .A3(n8618), .ZN(n8621) );
  NAND2_X1 U9911 ( .A1(n8621), .A2(n8620), .ZN(n8622) );
  INV_X1 U9912 ( .A(n8624), .ZN(n8628) );
  INV_X1 U9913 ( .A(n9123), .ZN(n8627) );
  INV_X1 U9914 ( .A(n8625), .ZN(n8626) );
  NAND3_X1 U9915 ( .A1(n8628), .A2(n8627), .A3(n8626), .ZN(n8629) );
  NAND2_X1 U9916 ( .A1(n8629), .A2(n9102), .ZN(n8633) );
  MUX2_X1 U9917 ( .A(n8631), .B(n8630), .S(n8663), .Z(n8632) );
  OR2_X1 U9918 ( .A1(n8768), .A2(n8676), .ZN(n8636) );
  NAND2_X1 U9919 ( .A1(n8768), .A2(n8676), .ZN(n8635) );
  MUX2_X1 U9920 ( .A(n8636), .B(n8635), .S(n9077), .Z(n8637) );
  NOR2_X1 U9921 ( .A1(n9179), .A2(n9091), .ZN(n8639) );
  MUX2_X1 U9922 ( .A(n8639), .B(n5217), .S(n8676), .Z(n8641) );
  MUX2_X1 U9923 ( .A(n8643), .B(n8642), .S(n8663), .Z(n8644) );
  MUX2_X1 U9924 ( .A(n8646), .B(n8645), .S(n8663), .Z(n8647) );
  NAND2_X1 U9925 ( .A1(n9048), .A2(n8647), .ZN(n8650) );
  INV_X1 U9926 ( .A(n9023), .ZN(n9034) );
  OR2_X1 U9927 ( .A1(n9039), .A2(n8709), .ZN(n8648) );
  MUX2_X1 U9928 ( .A(n8648), .B(n9032), .S(n8663), .Z(n8649) );
  INV_X1 U9929 ( .A(n9016), .ZN(n8654) );
  MUX2_X1 U9930 ( .A(n8652), .B(n8651), .S(n8663), .Z(n8653) );
  NAND3_X1 U9931 ( .A1(n8655), .A2(n8654), .A3(n8653), .ZN(n8659) );
  MUX2_X1 U9932 ( .A(n8656), .B(n9004), .S(n8663), .Z(n8657) );
  NOR2_X1 U9933 ( .A1(n9006), .A2(n8657), .ZN(n8658) );
  MUX2_X1 U9934 ( .A(n8661), .B(n8660), .S(n8663), .Z(n8662) );
  MUX2_X1 U9935 ( .A(n8664), .B(n8993), .S(n8663), .Z(n8667) );
  MUX2_X1 U9936 ( .A(n9000), .B(n8665), .S(n8676), .Z(n8666) );
  INV_X1 U9937 ( .A(n8667), .ZN(n8668) );
  NAND2_X1 U9938 ( .A1(n8676), .A2(n8673), .ZN(n8670) );
  AOI211_X1 U9939 ( .C1(n8671), .C2(n8681), .A(n8670), .B(n8677), .ZN(n8685)
         );
  NAND3_X1 U9940 ( .A1(n8675), .A2(n8674), .A3(n8673), .ZN(n8683) );
  NOR2_X1 U9941 ( .A1(n8676), .A2(n8686), .ZN(n8680) );
  INV_X1 U9942 ( .A(n8677), .ZN(n8678) );
  NAND4_X1 U9943 ( .A1(n8681), .A2(n8680), .A3(n8679), .A4(n8678), .ZN(n8682)
         );
  OAI211_X1 U9944 ( .C1(n8507), .C2(n8686), .A(n8683), .B(n8682), .ZN(n8684)
         );
  AOI21_X1 U9945 ( .B1(n8977), .B2(n8689), .A(n8688), .ZN(n8690) );
  XNOR2_X1 U9946 ( .A(n8690), .B(n8962), .ZN(n8697) );
  NAND3_X1 U9947 ( .A1(n8692), .A2(n8691), .A3(n6588), .ZN(n8693) );
  OAI211_X1 U9948 ( .C1(n8694), .C2(n8696), .A(n8693), .B(P2_B_REG_SCAN_IN), 
        .ZN(n8695) );
  OAI21_X1 U9949 ( .B1(n8697), .B2(n8696), .A(n8695), .ZN(P2_U3296) );
  INV_X1 U9950 ( .A(n9446), .ZN(n10516) );
  OAI222_X1 U9951 ( .A1(P2_U3151), .A2(n8699), .B1(n9262), .B2(n10516), .C1(
        n9267), .C2(n8698), .ZN(P2_U3265) );
  OAI211_X1 U9952 ( .C1(n8700), .C2(n8702), .A(n8701), .B(n8810), .ZN(n8706)
         );
  AOI22_X1 U9953 ( .A1(n9003), .A2(n8819), .B1(P2_REG3_REG_27__SCAN_IN), .B2(
        P2_U3151), .ZN(n8703) );
  OAI21_X1 U9954 ( .B1(n8735), .B2(n8816), .A(n8703), .ZN(n8704) );
  AOI21_X1 U9955 ( .B1(n9000), .B2(n8814), .A(n8704), .ZN(n8705) );
  OAI211_X1 U9956 ( .C1(n9009), .C2(n8823), .A(n8706), .B(n8705), .ZN(P2_U3154) );
  XNOR2_X1 U9957 ( .A(n8707), .B(n9045), .ZN(n8713) );
  AOI22_X1 U9958 ( .A1(n9075), .A2(n8800), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3151), .ZN(n8708) );
  OAI21_X1 U9959 ( .B1(n8709), .B2(n8803), .A(n8708), .ZN(n8711) );
  NOR2_X1 U9960 ( .A1(n9174), .A2(n8823), .ZN(n8710) );
  AOI211_X1 U9961 ( .C1(n9060), .C2(n8819), .A(n8711), .B(n8710), .ZN(n8712)
         );
  OAI21_X1 U9962 ( .B1(n8713), .B2(n8808), .A(n8712), .ZN(P2_U3156) );
  INV_X1 U9963 ( .A(n9237), .ZN(n8721) );
  OAI211_X1 U9964 ( .C1(n8716), .C2(n8715), .A(n8714), .B(n8810), .ZN(n8720)
         );
  NOR2_X1 U9965 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9752), .ZN(n8961) );
  AOI21_X1 U9966 ( .B1(n9104), .B2(n8814), .A(n8961), .ZN(n8717) );
  OAI21_X1 U9967 ( .B1(n8753), .B2(n8816), .A(n8717), .ZN(n8718) );
  AOI21_X1 U9968 ( .B1(n9107), .B2(n8819), .A(n8718), .ZN(n8719) );
  OAI211_X1 U9969 ( .C1(n8721), .C2(n8823), .A(n8720), .B(n8719), .ZN(P2_U3159) );
  XOR2_X1 U9970 ( .A(n8723), .B(n8724), .Z(n8730) );
  AOI22_X1 U9971 ( .A1(n9104), .A2(n8800), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3151), .ZN(n8726) );
  NAND2_X1 U9972 ( .A1(n8819), .A2(n9084), .ZN(n8725) );
  OAI211_X1 U9973 ( .C1(n8727), .C2(n8803), .A(n8726), .B(n8725), .ZN(n8728)
         );
  AOI21_X1 U9974 ( .B1(n9179), .B2(n8805), .A(n8728), .ZN(n8729) );
  OAI21_X1 U9975 ( .B1(n8730), .B2(n8808), .A(n8729), .ZN(P2_U3163) );
  XOR2_X1 U9976 ( .A(n8732), .B(n8731), .Z(n8738) );
  AOI22_X1 U9977 ( .A1(n9054), .A2(n8800), .B1(P2_REG3_REG_25__SCAN_IN), .B2(
        P2_U3151), .ZN(n8734) );
  NAND2_X1 U9978 ( .A1(n9027), .A2(n8819), .ZN(n8733) );
  OAI211_X1 U9979 ( .C1(n8735), .C2(n8803), .A(n8734), .B(n8733), .ZN(n8736)
         );
  AOI21_X1 U9980 ( .B1(n9162), .B2(n8805), .A(n8736), .ZN(n8737) );
  OAI21_X1 U9981 ( .B1(n8738), .B2(n8808), .A(n8737), .ZN(P2_U3165) );
  INV_X1 U9982 ( .A(n8739), .ZN(n9251) );
  OAI21_X1 U9983 ( .B1(n8740), .B2(n8743), .A(n8742), .ZN(n8744) );
  NAND2_X1 U9984 ( .A1(n8744), .A2(n8810), .ZN(n8749) );
  NAND2_X1 U9985 ( .A1(P2_REG3_REG_16__SCAN_IN), .A2(P2_U3151), .ZN(n10892) );
  OAI21_X1 U9986 ( .B1(n9118), .B2(n8803), .A(n10892), .ZN(n8747) );
  NOR2_X1 U9987 ( .A1(n8756), .A2(n8745), .ZN(n8746) );
  AOI211_X1 U9988 ( .C1(n8800), .C2(n8831), .A(n8747), .B(n8746), .ZN(n8748)
         );
  OAI211_X1 U9989 ( .C1(n9251), .C2(n8823), .A(n8749), .B(n8748), .ZN(P2_U3166) );
  XNOR2_X1 U9990 ( .A(n8751), .B(n8830), .ZN(n8752) );
  XNOR2_X1 U9991 ( .A(n8750), .B(n8752), .ZN(n8760) );
  NAND2_X1 U9992 ( .A1(P2_REG3_REG_17__SCAN_IN), .A2(P2_U3151), .ZN(n10912) );
  OAI21_X1 U9993 ( .B1(n8753), .B2(n8803), .A(n10912), .ZN(n8754) );
  AOI21_X1 U9994 ( .B1(n8800), .B2(n9135), .A(n8754), .ZN(n8755) );
  OAI21_X1 U9995 ( .B1(n9143), .B2(n8756), .A(n8755), .ZN(n8757) );
  AOI21_X1 U9996 ( .B1(n8758), .B2(n8805), .A(n8757), .ZN(n8759) );
  OAI21_X1 U9997 ( .B1(n8760), .B2(n8808), .A(n8759), .ZN(P2_U3168) );
  XOR2_X1 U9998 ( .A(n8762), .B(n8761), .Z(n8767) );
  AOI22_X1 U9999 ( .A1(n9065), .A2(n8800), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3151), .ZN(n8764) );
  NAND2_X1 U10000 ( .A1(n9047), .A2(n8819), .ZN(n8763) );
  OAI211_X1 U10001 ( .C1(n9044), .C2(n8803), .A(n8764), .B(n8763), .ZN(n8765)
         );
  AOI21_X1 U10002 ( .B1(n9039), .B2(n8805), .A(n8765), .ZN(n8766) );
  OAI21_X1 U10003 ( .B1(n8767), .B2(n8808), .A(n8766), .ZN(P2_U3169) );
  OAI21_X1 U10004 ( .B1(n8771), .B2(n8770), .A(n8769), .ZN(n8772) );
  NAND2_X1 U10005 ( .A1(n8772), .A2(n8810), .ZN(n8776) );
  AOI22_X1 U10006 ( .A1(n9064), .A2(n8814), .B1(P2_REG3_REG_20__SCAN_IN), .B2(
        P2_U3151), .ZN(n8773) );
  OAI21_X1 U10007 ( .B1(n9120), .B2(n8816), .A(n8773), .ZN(n8774) );
  AOI21_X1 U10008 ( .B1(n9092), .B2(n8819), .A(n8774), .ZN(n8775) );
  OAI211_X1 U10009 ( .C1(n9234), .C2(n8823), .A(n8776), .B(n8775), .ZN(
        P2_U3173) );
  AOI21_X1 U10010 ( .B1(n8777), .B2(n8778), .A(n8808), .ZN(n8780) );
  NAND2_X1 U10011 ( .A1(n8780), .A2(n8779), .ZN(n8784) );
  AOI22_X1 U10012 ( .A1(n9064), .A2(n8800), .B1(P2_REG3_REG_22__SCAN_IN), .B2(
        P2_U3151), .ZN(n8781) );
  OAI21_X1 U10013 ( .B1(n9045), .B2(n8803), .A(n8781), .ZN(n8782) );
  AOI21_X1 U10014 ( .B1(n9069), .B2(n8819), .A(n8782), .ZN(n8783) );
  OAI211_X1 U10015 ( .C1(n8785), .C2(n8823), .A(n8784), .B(n8783), .ZN(
        P2_U3175) );
  NAND2_X1 U10016 ( .A1(n8788), .A2(n8787), .ZN(n8790) );
  AOI21_X1 U10017 ( .B1(n8790), .B2(n8789), .A(n8808), .ZN(n8792) );
  NAND2_X1 U10018 ( .A1(n8792), .A2(n8791), .ZN(n8797) );
  INV_X1 U10019 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n8793) );
  NOR2_X1 U10020 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n8793), .ZN(n8915) );
  AOI21_X1 U10021 ( .B1(n8829), .B2(n8814), .A(n8915), .ZN(n8794) );
  OAI21_X1 U10022 ( .B1(n9118), .B2(n8816), .A(n8794), .ZN(n8795) );
  AOI21_X1 U10023 ( .B1(n9124), .B2(n8819), .A(n8795), .ZN(n8796) );
  OAI211_X1 U10024 ( .C1(n9242), .C2(n8823), .A(n8797), .B(n8796), .ZN(
        P2_U3178) );
  XOR2_X1 U10025 ( .A(n8799), .B(n8798), .Z(n8809) );
  AOI22_X1 U10026 ( .A1(n8828), .A2(n8800), .B1(P2_REG3_REG_26__SCAN_IN), .B2(
        P2_U3151), .ZN(n8802) );
  NAND2_X1 U10027 ( .A1(n9018), .A2(n8819), .ZN(n8801) );
  OAI211_X1 U10028 ( .C1(n9015), .C2(n8803), .A(n8802), .B(n8801), .ZN(n8804)
         );
  AOI21_X1 U10029 ( .B1(n8806), .B2(n8805), .A(n8804), .ZN(n8807) );
  OAI21_X1 U10030 ( .B1(n8809), .B2(n8808), .A(n8807), .ZN(P2_U3180) );
  OAI211_X1 U10031 ( .C1(n8813), .C2(n8812), .A(n8811), .B(n8810), .ZN(n8822)
         );
  NOR2_X1 U10032 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10000), .ZN(n10871) );
  AOI21_X1 U10033 ( .B1(n9135), .B2(n8814), .A(n10871), .ZN(n8815) );
  OAI21_X1 U10034 ( .B1(n8817), .B2(n8816), .A(n8815), .ZN(n8818) );
  AOI21_X1 U10035 ( .B1(n8820), .B2(n8819), .A(n8818), .ZN(n8821) );
  OAI211_X1 U10036 ( .C1(n8824), .C2(n8823), .A(n8822), .B(n8821), .ZN(
        P2_U3181) );
  MUX2_X1 U10037 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n8825), .S(P2_U3893), .Z(
        P2_U3521) );
  MUX2_X1 U10038 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n8826), .S(P2_U3893), .Z(
        P2_U3520) );
  MUX2_X1 U10039 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n9000), .S(P2_U3893), .Z(
        P2_U3519) );
  MUX2_X1 U10040 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n8827), .S(P2_U3893), .Z(
        P2_U3518) );
  MUX2_X1 U10041 ( .A(n9025), .B(P2_DATAO_REG_26__SCAN_IN), .S(n8913), .Z(
        P2_U3517) );
  MUX2_X1 U10042 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n8828), .S(P2_U3893), .Z(
        P2_U3516) );
  MUX2_X1 U10043 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n9054), .S(P2_U3893), .Z(
        P2_U3515) );
  MUX2_X1 U10044 ( .A(n9065), .B(P2_DATAO_REG_23__SCAN_IN), .S(n8913), .Z(
        P2_U3514) );
  MUX2_X1 U10045 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9075), .S(P2_U3893), .Z(
        P2_U3513) );
  MUX2_X1 U10046 ( .A(n9064), .B(P2_DATAO_REG_21__SCAN_IN), .S(n8913), .Z(
        P2_U3512) );
  MUX2_X1 U10047 ( .A(n9104), .B(P2_DATAO_REG_20__SCAN_IN), .S(n8913), .Z(
        P2_U3511) );
  MUX2_X1 U10048 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n8829), .S(P2_U3893), .Z(
        P2_U3510) );
  MUX2_X1 U10049 ( .A(n9134), .B(P2_DATAO_REG_18__SCAN_IN), .S(n8913), .Z(
        P2_U3509) );
  MUX2_X1 U10050 ( .A(n8830), .B(P2_DATAO_REG_17__SCAN_IN), .S(n8913), .Z(
        P2_U3508) );
  MUX2_X1 U10051 ( .A(n9135), .B(P2_DATAO_REG_16__SCAN_IN), .S(n8913), .Z(
        P2_U3507) );
  MUX2_X1 U10052 ( .A(n8831), .B(P2_DATAO_REG_15__SCAN_IN), .S(n8913), .Z(
        P2_U3506) );
  MUX2_X1 U10053 ( .A(n8832), .B(P2_DATAO_REG_14__SCAN_IN), .S(n8913), .Z(
        P2_U3505) );
  MUX2_X1 U10054 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n8833), .S(P2_U3893), .Z(
        P2_U3504) );
  MUX2_X1 U10055 ( .A(n8834), .B(P2_DATAO_REG_12__SCAN_IN), .S(n8913), .Z(
        P2_U3503) );
  MUX2_X1 U10056 ( .A(n8835), .B(P2_DATAO_REG_11__SCAN_IN), .S(n8913), .Z(
        P2_U3502) );
  MUX2_X1 U10057 ( .A(n8836), .B(P2_DATAO_REG_10__SCAN_IN), .S(n8913), .Z(
        P2_U3501) );
  MUX2_X1 U10058 ( .A(n8837), .B(P2_DATAO_REG_9__SCAN_IN), .S(n8913), .Z(
        P2_U3500) );
  MUX2_X1 U10059 ( .A(n8838), .B(P2_DATAO_REG_8__SCAN_IN), .S(n8913), .Z(
        P2_U3499) );
  MUX2_X1 U10060 ( .A(n8839), .B(P2_DATAO_REG_7__SCAN_IN), .S(n8913), .Z(
        P2_U3498) );
  MUX2_X1 U10061 ( .A(n8840), .B(P2_DATAO_REG_6__SCAN_IN), .S(n8913), .Z(
        P2_U3497) );
  MUX2_X1 U10062 ( .A(n8841), .B(P2_DATAO_REG_5__SCAN_IN), .S(n8913), .Z(
        P2_U3496) );
  MUX2_X1 U10063 ( .A(n8842), .B(P2_DATAO_REG_4__SCAN_IN), .S(n8913), .Z(
        P2_U3495) );
  MUX2_X1 U10064 ( .A(n8843), .B(P2_DATAO_REG_3__SCAN_IN), .S(n8913), .Z(
        P2_U3494) );
  MUX2_X1 U10065 ( .A(n8844), .B(P2_DATAO_REG_2__SCAN_IN), .S(n8913), .Z(
        P2_U3493) );
  MUX2_X1 U10066 ( .A(n6695), .B(P2_DATAO_REG_1__SCAN_IN), .S(n8913), .Z(
        P2_U3492) );
  OAI211_X1 U10067 ( .C1(n8847), .C2(n8846), .A(n8845), .B(n10904), .ZN(n8860)
         );
  AOI22_X1 U10068 ( .A1(n10896), .A2(n8848), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        P2_U3151), .ZN(n8859) );
  OAI21_X1 U10069 ( .B1(n8851), .B2(n8850), .A(n8849), .ZN(n8856) );
  OAI21_X1 U10070 ( .B1(n8854), .B2(n8853), .A(n8852), .ZN(n8855) );
  AOI22_X1 U10071 ( .A1(n10905), .A2(n8856), .B1(n10790), .B2(n8855), .ZN(
        n8858) );
  NAND2_X1 U10072 ( .A1(n10895), .A2(P2_ADDR_REG_2__SCAN_IN), .ZN(n8857) );
  NAND4_X1 U10073 ( .A1(n8860), .A2(n8859), .A3(n8858), .A4(n8857), .ZN(
        P2_U3184) );
  XNOR2_X1 U10074 ( .A(n8948), .B(P2_REG1_REG_18__SCAN_IN), .ZN(n8950) );
  AOI22_X1 U10075 ( .A1(n10879), .A2(n9207), .B1(P2_REG1_REG_16__SCAN_IN), 
        .B2(n8938), .ZN(n10882) );
  NAND2_X1 U10076 ( .A1(P2_REG1_REG_12__SCAN_IN), .A2(n8927), .ZN(n8867) );
  AOI22_X1 U10077 ( .A1(n10812), .A2(n8886), .B1(P2_REG1_REG_12__SCAN_IN), 
        .B2(n8927), .ZN(n10815) );
  INV_X1 U10078 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n8864) );
  MUX2_X1 U10079 ( .A(n8864), .B(P2_REG1_REG_10__SCAN_IN), .S(n10777), .Z(
        n10784) );
  OR2_X1 U10080 ( .A1(n8920), .A2(n8861), .ZN(n8863) );
  NAND2_X1 U10081 ( .A1(n10784), .A2(n10785), .ZN(n10783) );
  OAI21_X1 U10082 ( .B1(n10777), .B2(n8864), .A(n10783), .ZN(n8865) );
  NAND2_X1 U10083 ( .A1(n8898), .A2(n8865), .ZN(n8866) );
  XNOR2_X1 U10084 ( .A(n8865), .B(n10797), .ZN(n10802) );
  NAND2_X1 U10085 ( .A1(P2_REG1_REG_11__SCAN_IN), .A2(n10802), .ZN(n10801) );
  NAND2_X1 U10086 ( .A1(n5366), .A2(n8868), .ZN(n8869) );
  NAND2_X1 U10087 ( .A1(P2_REG1_REG_13__SCAN_IN), .A2(n10831), .ZN(n10830) );
  NAND2_X1 U10088 ( .A1(n8869), .A2(n10830), .ZN(n10847) );
  XNOR2_X1 U10089 ( .A(n10845), .B(P2_REG1_REG_14__SCAN_IN), .ZN(n10846) );
  AOI22_X1 U10090 ( .A1(n10847), .A2(n10846), .B1(P2_REG1_REG_14__SCAN_IN), 
        .B2(n8930), .ZN(n8870) );
  NAND2_X1 U10091 ( .A1(n8933), .A2(n8871), .ZN(n8872) );
  NAND2_X1 U10092 ( .A1(n10882), .A2(n10881), .ZN(n10880) );
  NAND2_X1 U10093 ( .A1(n8941), .A2(n8873), .ZN(n8874) );
  XOR2_X1 U10094 ( .A(n8950), .B(n8951), .Z(n8949) );
  OR2_X1 U10095 ( .A1(n6588), .A2(n9144), .ZN(n8876) );
  NAND2_X1 U10096 ( .A1(n6588), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n8875) );
  NAND2_X1 U10097 ( .A1(n8876), .A2(n8875), .ZN(n8877) );
  OR2_X1 U10098 ( .A1(n8877), .A2(n8941), .ZN(n8906) );
  XNOR2_X1 U10099 ( .A(n8877), .B(n10897), .ZN(n10902) );
  MUX2_X1 U10100 ( .A(n8936), .B(n9207), .S(n6588), .Z(n8878) );
  NAND2_X1 U10101 ( .A1(n10879), .A2(n8878), .ZN(n8905) );
  XNOR2_X1 U10102 ( .A(n8878), .B(n8938), .ZN(n10885) );
  MUX2_X1 U10103 ( .A(n8880), .B(n8879), .S(n6588), .Z(n8881) );
  NAND2_X1 U10104 ( .A1(n10863), .A2(n8881), .ZN(n8904) );
  XNOR2_X1 U10105 ( .A(n8881), .B(n8933), .ZN(n10868) );
  MUX2_X1 U10106 ( .A(P2_REG2_REG_14__SCAN_IN), .B(P2_REG1_REG_14__SCAN_IN), 
        .S(n6588), .Z(n8882) );
  OR2_X1 U10107 ( .A1(n8930), .A2(n8882), .ZN(n8903) );
  XNOR2_X1 U10108 ( .A(n8882), .B(n10845), .ZN(n10850) );
  MUX2_X1 U10109 ( .A(n8884), .B(n8883), .S(n6588), .Z(n8885) );
  NAND2_X1 U10110 ( .A1(n10829), .A2(n8885), .ZN(n8902) );
  XNOR2_X1 U10111 ( .A(n8885), .B(n5366), .ZN(n10834) );
  MUX2_X1 U10112 ( .A(n8887), .B(n8886), .S(n6588), .Z(n8888) );
  NAND2_X1 U10113 ( .A1(n10812), .A2(n8888), .ZN(n8901) );
  XNOR2_X1 U10114 ( .A(n8888), .B(n8927), .ZN(n10818) );
  MUX2_X1 U10115 ( .A(n8890), .B(n8889), .S(n6588), .Z(n8899) );
  NAND2_X1 U10116 ( .A1(n10797), .A2(n8899), .ZN(n8900) );
  AOI21_X1 U10117 ( .B1(n8893), .B2(n8892), .A(n8891), .ZN(n10782) );
  MUX2_X1 U10118 ( .A(n8894), .B(n8864), .S(n6588), .Z(n8895) );
  NAND2_X1 U10119 ( .A1(n8895), .A2(n10777), .ZN(n10779) );
  OR2_X1 U10120 ( .A1(n6588), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n8897) );
  NAND2_X1 U10121 ( .A1(n6588), .A2(n8864), .ZN(n8896) );
  AND3_X1 U10122 ( .A1(n8897), .A2(n8896), .A3(n8923), .ZN(n10778) );
  AOI21_X1 U10123 ( .B1(n10782), .B2(n10779), .A(n10778), .ZN(n10800) );
  XNOR2_X1 U10124 ( .A(n8899), .B(n8898), .ZN(n10799) );
  NAND2_X1 U10125 ( .A1(n10800), .A2(n10799), .ZN(n10798) );
  NAND2_X1 U10126 ( .A1(n8900), .A2(n10798), .ZN(n10817) );
  NAND2_X1 U10127 ( .A1(n10818), .A2(n10817), .ZN(n10816) );
  NAND2_X1 U10128 ( .A1(n8901), .A2(n10816), .ZN(n10833) );
  NAND2_X1 U10129 ( .A1(n10834), .A2(n10833), .ZN(n10832) );
  NAND2_X1 U10130 ( .A1(n8902), .A2(n10832), .ZN(n10849) );
  NAND2_X1 U10131 ( .A1(n10850), .A2(n10849), .ZN(n10848) );
  NAND2_X1 U10132 ( .A1(n8903), .A2(n10848), .ZN(n10867) );
  NAND2_X1 U10133 ( .A1(n10868), .A2(n10867), .ZN(n10866) );
  NAND2_X1 U10134 ( .A1(n8904), .A2(n10866), .ZN(n10884) );
  NAND2_X1 U10135 ( .A1(n10885), .A2(n10884), .ZN(n10883) );
  NAND2_X1 U10136 ( .A1(n8905), .A2(n10883), .ZN(n10901) );
  NAND2_X1 U10137 ( .A1(n10902), .A2(n10901), .ZN(n10900) );
  NAND2_X1 U10138 ( .A1(n8906), .A2(n10900), .ZN(n8910) );
  OR2_X1 U10139 ( .A1(n6588), .A2(n8916), .ZN(n8908) );
  NAND2_X1 U10140 ( .A1(n6588), .A2(P2_REG1_REG_18__SCAN_IN), .ZN(n8907) );
  AND2_X1 U10141 ( .A1(n8908), .A2(n8907), .ZN(n8909) );
  NAND2_X1 U10142 ( .A1(n8910), .A2(n8909), .ZN(n8964) );
  INV_X1 U10143 ( .A(n8964), .ZN(n8911) );
  NOR2_X1 U10144 ( .A1(n8910), .A2(n8909), .ZN(n8966) );
  OR2_X1 U10145 ( .A1(n8911), .A2(n8966), .ZN(n8914) );
  OAI21_X1 U10146 ( .B1(n8914), .B2(n8913), .A(n8912), .ZN(n8947) );
  NAND3_X1 U10147 ( .A1(n8914), .A2(n10904), .A3(n8965), .ZN(n8946) );
  INV_X1 U10148 ( .A(n8915), .ZN(n8945) );
  NAND2_X1 U10149 ( .A1(n10895), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n8944) );
  OR2_X1 U10150 ( .A1(n8948), .A2(n8916), .ZN(n8918) );
  NAND2_X1 U10151 ( .A1(n8948), .A2(n8916), .ZN(n8917) );
  AND2_X1 U10152 ( .A1(n8918), .A2(n8917), .ZN(n8959) );
  OAI22_X1 U10153 ( .A1(n8922), .A2(n8921), .B1(n8920), .B2(n8919), .ZN(n10789) );
  MUX2_X1 U10154 ( .A(n8894), .B(P2_REG2_REG_10__SCAN_IN), .S(n10777), .Z(
        n10788) );
  AOI21_X1 U10155 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n8923), .A(n10791), .ZN(
        n8924) );
  NOR2_X1 U10156 ( .A1(n10797), .A2(n8924), .ZN(n8925) );
  NAND2_X1 U10157 ( .A1(P2_REG2_REG_12__SCAN_IN), .A2(n8927), .ZN(n8926) );
  OAI21_X1 U10158 ( .B1(n8927), .B2(P2_REG2_REG_12__SCAN_IN), .A(n8926), .ZN(
        n10823) );
  MUX2_X1 U10159 ( .A(P2_REG2_REG_14__SCAN_IN), .B(n8929), .S(n10845), .Z(
        n10857) );
  NAND2_X1 U10160 ( .A1(n8930), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n8931) );
  NAND2_X1 U10161 ( .A1(n10854), .A2(n8931), .ZN(n8934) );
  INV_X1 U10162 ( .A(n8934), .ZN(n8932) );
  NOR2_X1 U10163 ( .A1(n10863), .A2(n8932), .ZN(n8935) );
  XNOR2_X1 U10164 ( .A(n8934), .B(n8933), .ZN(n10873) );
  NOR2_X1 U10165 ( .A1(n10873), .A2(n8880), .ZN(n10872) );
  NOR2_X1 U10166 ( .A1(n8938), .A2(n8936), .ZN(n8937) );
  AOI21_X1 U10167 ( .B1(n8936), .B2(n8938), .A(n8937), .ZN(n10888) );
  INV_X1 U10168 ( .A(n8953), .ZN(n8955) );
  INV_X1 U10169 ( .A(n8939), .ZN(n8940) );
  OAI21_X1 U10170 ( .B1(n8941), .B2(n8940), .A(n8953), .ZN(n10908) );
  NOR2_X1 U10171 ( .A1(n8955), .A2(n10907), .ZN(n8942) );
  XNOR2_X1 U10172 ( .A(n8959), .B(n8942), .ZN(n8943) );
  AOI22_X1 U10173 ( .A1(n8951), .A2(n8950), .B1(P2_REG1_REG_18__SCAN_IN), .B2(
        n8965), .ZN(n8952) );
  XNOR2_X1 U10174 ( .A(n8962), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n8967) );
  MUX2_X1 U10175 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n9109), .S(n8962), .Z(n8969) );
  NAND2_X1 U10176 ( .A1(n8953), .A2(n8916), .ZN(n8954) );
  AOI21_X1 U10177 ( .B1(n10896), .B2(n8962), .A(n8961), .ZN(n8963) );
  OAI21_X1 U10178 ( .B1(n8966), .B2(n8965), .A(n8964), .ZN(n8971) );
  INV_X1 U10179 ( .A(n8967), .ZN(n8968) );
  MUX2_X1 U10180 ( .A(n8969), .B(n8968), .S(n6588), .Z(n8970) );
  XNOR2_X1 U10181 ( .A(n8971), .B(n8970), .ZN(n8972) );
  NOR2_X1 U10182 ( .A1(n8972), .A2(n10772), .ZN(n8973) );
  INV_X1 U10183 ( .A(n8975), .ZN(n8976) );
  NOR2_X1 U10184 ( .A1(n8977), .A2(n8976), .ZN(n9212) );
  NOR2_X1 U10185 ( .A1(n8978), .A2(n9142), .ZN(n8985) );
  NOR3_X1 U10186 ( .A1(n9212), .A2(n9150), .A3(n8985), .ZN(n8981) );
  NOR2_X1 U10187 ( .A1(n9145), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8979) );
  OAI22_X1 U10188 ( .A1(n9214), .A2(n9141), .B1(n8981), .B2(n8979), .ZN(
        P2_U3202) );
  NOR2_X1 U10189 ( .A1(n9145), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8980) );
  OAI22_X1 U10190 ( .A1(n9217), .A2(n9141), .B1(n8981), .B2(n8980), .ZN(
        P2_U3203) );
  NAND2_X1 U10191 ( .A1(n8982), .A2(n9145), .ZN(n8987) );
  NOR2_X1 U10192 ( .A1(n8983), .A2(n9141), .ZN(n8984) );
  AOI211_X1 U10193 ( .C1(n9150), .C2(P2_REG2_REG_29__SCAN_IN), .A(n8985), .B(
        n8984), .ZN(n8986) );
  OAI211_X1 U10194 ( .C1(n8989), .C2(n8988), .A(n8987), .B(n8986), .ZN(
        P2_U3204) );
  INV_X1 U10195 ( .A(n8990), .ZN(n8997) );
  AOI22_X1 U10196 ( .A1(n8991), .A2(n9125), .B1(n9150), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n8992) );
  OAI21_X1 U10197 ( .B1(n8993), .B2(n9141), .A(n8992), .ZN(n8994) );
  AOI21_X1 U10198 ( .B1(n8995), .B2(n9148), .A(n8994), .ZN(n8996) );
  OAI21_X1 U10199 ( .B1(n8997), .B2(n9150), .A(n8996), .ZN(P2_U3205) );
  XNOR2_X1 U10200 ( .A(n8999), .B(n8998), .ZN(n9001) );
  INV_X1 U10201 ( .A(n9157), .ZN(n9002) );
  AOI21_X1 U10202 ( .B1(n9125), .B2(n9003), .A(n9002), .ZN(n9012) );
  NOR2_X1 U10203 ( .A1(n9005), .A2(n9004), .ZN(n9007) );
  OAI22_X1 U10204 ( .A1(n9009), .A2(n9141), .B1(n9008), .B2(n9145), .ZN(n9010)
         );
  AOI21_X1 U10205 ( .B1(n9156), .B2(n9148), .A(n9010), .ZN(n9011) );
  OAI21_X1 U10206 ( .B1(n9012), .B2(n9150), .A(n9011), .ZN(P2_U3206) );
  XNOR2_X1 U10207 ( .A(n9013), .B(n9016), .ZN(n9014) );
  OAI222_X1 U10208 ( .A1(n9121), .A2(n9015), .B1(n9119), .B2(n9044), .C1(n9116), .C2(n9014), .ZN(n9158) );
  INV_X1 U10209 ( .A(n9158), .ZN(n9022) );
  XNOR2_X1 U10210 ( .A(n9017), .B(n9016), .ZN(n9159) );
  AOI22_X1 U10211 ( .A1(n9018), .A2(n9125), .B1(n9150), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9019) );
  OAI21_X1 U10212 ( .B1(n9222), .B2(n9141), .A(n9019), .ZN(n9020) );
  AOI21_X1 U10213 ( .B1(n9159), .B2(n9148), .A(n9020), .ZN(n9021) );
  OAI21_X1 U10214 ( .B1(n9022), .B2(n9150), .A(n9021), .ZN(P2_U3207) );
  XNOR2_X1 U10215 ( .A(n9024), .B(n9023), .ZN(n9026) );
  AOI222_X1 U10216 ( .A1(n9130), .A2(n9026), .B1(n9054), .B2(n9136), .C1(n9025), .C2(n9133), .ZN(n9165) );
  INV_X1 U10217 ( .A(n9165), .ZN(n9031) );
  INV_X1 U10218 ( .A(n9027), .ZN(n9028) );
  OAI22_X1 U10219 ( .A1(n9029), .A2(n9040), .B1(n9028), .B2(n9142), .ZN(n9030)
         );
  OAI21_X1 U10220 ( .B1(n9031), .B2(n9030), .A(n9145), .ZN(n9037) );
  NAND2_X1 U10221 ( .A1(n9049), .A2(n9048), .ZN(n9033) );
  NAND2_X1 U10222 ( .A1(n9033), .A2(n9032), .ZN(n9035) );
  XNOR2_X1 U10223 ( .A(n9035), .B(n9034), .ZN(n9163) );
  NAND2_X1 U10224 ( .A1(n9163), .A2(n9148), .ZN(n9036) );
  OAI211_X1 U10225 ( .C1(n9145), .C2(n9038), .A(n9037), .B(n9036), .ZN(
        P2_U3208) );
  INV_X1 U10226 ( .A(n9039), .ZN(n9227) );
  NOR2_X1 U10227 ( .A1(n9227), .A2(n9040), .ZN(n9046) );
  XNOR2_X1 U10228 ( .A(n9042), .B(n9041), .ZN(n9043) );
  OAI222_X1 U10229 ( .A1(n9119), .A2(n9045), .B1(n9121), .B2(n9044), .C1(n9116), .C2(n9043), .ZN(n9166) );
  AOI211_X1 U10230 ( .C1(n9125), .C2(n9047), .A(n9046), .B(n9166), .ZN(n9051)
         );
  XNOR2_X1 U10231 ( .A(n9049), .B(n9048), .ZN(n9167) );
  AOI22_X1 U10232 ( .A1(n9167), .A2(n9148), .B1(P2_REG2_REG_24__SCAN_IN), .B2(
        n9150), .ZN(n9050) );
  OAI21_X1 U10233 ( .B1(n9051), .B2(n9150), .A(n9050), .ZN(P2_U3209) );
  XNOR2_X1 U10234 ( .A(n9053), .B(n9052), .ZN(n9055) );
  AOI222_X1 U10235 ( .A1(n9130), .A2(n9055), .B1(n9075), .B2(n9136), .C1(n9054), .C2(n9133), .ZN(n9172) );
  INV_X1 U10236 ( .A(n9056), .ZN(n9059) );
  OAI21_X1 U10237 ( .B1(n9059), .B2(n9058), .A(n9057), .ZN(n9170) );
  AOI22_X1 U10238 ( .A1(n9060), .A2(n9125), .B1(n9150), .B2(
        P2_REG2_REG_23__SCAN_IN), .ZN(n9061) );
  OAI21_X1 U10239 ( .B1(n9174), .B2(n9141), .A(n9061), .ZN(n9062) );
  AOI21_X1 U10240 ( .B1(n9170), .B2(n9148), .A(n9062), .ZN(n9063) );
  OAI21_X1 U10241 ( .B1(n9172), .B2(n9150), .A(n9063), .ZN(P2_U3210) );
  XNOR2_X1 U10242 ( .A(n5220), .B(n9067), .ZN(n9066) );
  AOI222_X1 U10243 ( .A1(n9130), .A2(n9066), .B1(n9065), .B2(n9133), .C1(n9064), .C2(n9136), .ZN(n9178) );
  XNOR2_X1 U10244 ( .A(n9068), .B(n9067), .ZN(n9176) );
  NAND2_X1 U10245 ( .A1(n9175), .A2(n9111), .ZN(n9071) );
  AOI22_X1 U10246 ( .A1(n9069), .A2(n9125), .B1(n9150), .B2(
        P2_REG2_REG_22__SCAN_IN), .ZN(n9070) );
  NAND2_X1 U10247 ( .A1(n9071), .A2(n9070), .ZN(n9072) );
  AOI21_X1 U10248 ( .B1(n9176), .B2(n9148), .A(n9072), .ZN(n9073) );
  OAI21_X1 U10249 ( .B1(n9178), .B2(n9150), .A(n9073), .ZN(P2_U3211) );
  XNOR2_X1 U10250 ( .A(n9074), .B(n9080), .ZN(n9079) );
  NAND2_X1 U10251 ( .A1(n9075), .A2(n9133), .ZN(n9076) );
  OAI21_X1 U10252 ( .B1(n9077), .B2(n9119), .A(n9076), .ZN(n9078) );
  AOI21_X1 U10253 ( .B1(n9079), .B2(n9130), .A(n9078), .ZN(n9183) );
  NAND2_X1 U10254 ( .A1(n9081), .A2(n9080), .ZN(n9082) );
  NAND2_X1 U10255 ( .A1(n9083), .A2(n9082), .ZN(n9181) );
  INV_X1 U10256 ( .A(n9179), .ZN(n9086) );
  AOI22_X1 U10257 ( .A1(n9125), .A2(n9084), .B1(n9150), .B2(
        P2_REG2_REG_21__SCAN_IN), .ZN(n9085) );
  OAI21_X1 U10258 ( .B1(n9086), .B2(n9141), .A(n9085), .ZN(n9087) );
  AOI21_X1 U10259 ( .B1(n9181), .B2(n9148), .A(n9087), .ZN(n9088) );
  OAI21_X1 U10260 ( .B1(n9183), .B2(n9150), .A(n9088), .ZN(P2_U3212) );
  AOI21_X1 U10261 ( .B1(n9093), .B2(n9089), .A(n5402), .ZN(n9090) );
  OAI222_X1 U10262 ( .A1(n9119), .A2(n9120), .B1(n9121), .B2(n9091), .C1(n9116), .C2(n9090), .ZN(n9184) );
  AOI21_X1 U10263 ( .B1(n9125), .B2(n9092), .A(n9184), .ZN(n9098) );
  XOR2_X1 U10264 ( .A(n9094), .B(n9093), .Z(n9185) );
  OAI22_X1 U10265 ( .A1(n9234), .A2(n9141), .B1(n9095), .B2(n9145), .ZN(n9096)
         );
  AOI21_X1 U10266 ( .B1(n9185), .B2(n9148), .A(n9096), .ZN(n9097) );
  OAI21_X1 U10267 ( .B1(n9098), .B2(n9150), .A(n9097), .ZN(P2_U3213) );
  OAI21_X1 U10268 ( .B1(n9100), .B2(n9102), .A(n9099), .ZN(n9189) );
  XNOR2_X1 U10269 ( .A(n9101), .B(n9102), .ZN(n9103) );
  NAND2_X1 U10270 ( .A1(n9103), .A2(n9130), .ZN(n9106) );
  AOI22_X1 U10271 ( .A1(n9104), .A2(n9133), .B1(n9136), .B2(n9134), .ZN(n9105)
         );
  NAND2_X1 U10272 ( .A1(n9106), .A2(n9105), .ZN(n9191) );
  NAND2_X1 U10273 ( .A1(n9191), .A2(n9145), .ZN(n9113) );
  INV_X1 U10274 ( .A(n9107), .ZN(n9108) );
  OAI22_X1 U10275 ( .A1(n9145), .A2(n9109), .B1(n9108), .B2(n9142), .ZN(n9110)
         );
  AOI21_X1 U10276 ( .B1(n9237), .B2(n9111), .A(n9110), .ZN(n9112) );
  OAI211_X1 U10277 ( .C1(n9189), .C2(n9114), .A(n9113), .B(n9112), .ZN(
        P2_U3214) );
  XNOR2_X1 U10278 ( .A(n9115), .B(n9123), .ZN(n9117) );
  OAI222_X1 U10279 ( .A1(n9121), .A2(n9120), .B1(n9119), .B2(n9118), .C1(n9117), .C2(n9116), .ZN(n9194) );
  INV_X1 U10280 ( .A(n9194), .ZN(n9129) );
  XNOR2_X1 U10281 ( .A(n9122), .B(n9123), .ZN(n9195) );
  AOI22_X1 U10282 ( .A1(n9150), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9125), .B2(
        n9124), .ZN(n9126) );
  OAI21_X1 U10283 ( .B1(n9242), .B2(n9141), .A(n9126), .ZN(n9127) );
  AOI21_X1 U10284 ( .B1(n9195), .B2(n9148), .A(n9127), .ZN(n9128) );
  OAI21_X1 U10285 ( .B1(n9129), .B2(n9150), .A(n9128), .ZN(P2_U3215) );
  OAI211_X1 U10286 ( .C1(n9132), .C2(n9140), .A(n9131), .B(n9130), .ZN(n9138)
         );
  AOI22_X1 U10287 ( .A1(n9136), .A2(n9135), .B1(n9134), .B2(n9133), .ZN(n9137)
         );
  NAND2_X1 U10288 ( .A1(n9138), .A2(n9137), .ZN(n9198) );
  INV_X1 U10289 ( .A(n9198), .ZN(n9151) );
  XNOR2_X1 U10290 ( .A(n9139), .B(n9140), .ZN(n9199) );
  NOR2_X1 U10291 ( .A1(n9246), .A2(n9141), .ZN(n9147) );
  OAI22_X1 U10292 ( .A1(n9145), .A2(n9144), .B1(n9143), .B2(n9142), .ZN(n9146)
         );
  AOI211_X1 U10293 ( .C1(n9199), .C2(n9148), .A(n9147), .B(n9146), .ZN(n9149)
         );
  OAI21_X1 U10294 ( .B1(n9151), .B2(n9150), .A(n9149), .ZN(P2_U3216) );
  NAND2_X1 U10295 ( .A1(n9212), .A2(n9206), .ZN(n9153) );
  NAND2_X1 U10296 ( .A1(n9210), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n9152) );
  OAI211_X1 U10297 ( .C1(n9214), .C2(n9209), .A(n9153), .B(n9152), .ZN(
        P2_U3490) );
  NAND2_X1 U10298 ( .A1(n9210), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n9154) );
  OAI211_X1 U10299 ( .C1(n9217), .C2(n9209), .A(n9154), .B(n9153), .ZN(
        P2_U3489) );
  AOI21_X1 U10300 ( .B1(n9159), .B2(n9204), .A(n9158), .ZN(n9219) );
  INV_X1 U10301 ( .A(P2_REG1_REG_26__SCAN_IN), .ZN(n9160) );
  MUX2_X1 U10302 ( .A(n9219), .B(n9160), .S(n9210), .Z(n9161) );
  OAI21_X1 U10303 ( .B1(n9222), .B2(n9209), .A(n9161), .ZN(P2_U3485) );
  AOI22_X1 U10304 ( .A1(n9163), .A2(n9204), .B1(n9180), .B2(n9162), .ZN(n9164)
         );
  NAND2_X1 U10305 ( .A1(n9165), .A2(n9164), .ZN(n9223) );
  MUX2_X1 U10306 ( .A(n9223), .B(P2_REG1_REG_25__SCAN_IN), .S(n9210), .Z(
        P2_U3484) );
  AOI21_X1 U10307 ( .B1(n9204), .B2(n9167), .A(n9166), .ZN(n9224) );
  INV_X1 U10308 ( .A(P2_REG1_REG_24__SCAN_IN), .ZN(n9168) );
  MUX2_X1 U10309 ( .A(n9224), .B(n9168), .S(n9210), .Z(n9169) );
  OAI21_X1 U10310 ( .B1(n9227), .B2(n9209), .A(n9169), .ZN(P2_U3483) );
  NAND2_X1 U10311 ( .A1(n9170), .A2(n9204), .ZN(n9171) );
  OAI211_X1 U10312 ( .C1(n9174), .C2(n9173), .A(n9172), .B(n9171), .ZN(n9228)
         );
  MUX2_X1 U10313 ( .A(n9228), .B(P2_REG1_REG_23__SCAN_IN), .S(n9210), .Z(
        P2_U3482) );
  AOI22_X1 U10314 ( .A1(n9176), .A2(n9204), .B1(n9180), .B2(n9175), .ZN(n9177)
         );
  NAND2_X1 U10315 ( .A1(n9178), .A2(n9177), .ZN(n9229) );
  MUX2_X1 U10316 ( .A(n9229), .B(P2_REG1_REG_22__SCAN_IN), .S(n9210), .Z(
        P2_U3481) );
  AOI22_X1 U10317 ( .A1(n9181), .A2(n9204), .B1(n9180), .B2(n9179), .ZN(n9182)
         );
  NAND2_X1 U10318 ( .A1(n9183), .A2(n9182), .ZN(n9230) );
  MUX2_X1 U10319 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9230), .S(n9206), .Z(
        P2_U3480) );
  INV_X1 U10320 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n9186) );
  AOI21_X1 U10321 ( .B1(n9185), .B2(n9204), .A(n9184), .ZN(n9231) );
  MUX2_X1 U10322 ( .A(n9186), .B(n9231), .S(n9206), .Z(n9187) );
  OAI21_X1 U10323 ( .B1(n9234), .B2(n9209), .A(n9187), .ZN(P2_U3479) );
  NOR2_X1 U10324 ( .A1(n9189), .A2(n9188), .ZN(n9190) );
  OR2_X1 U10325 ( .A1(n9191), .A2(n9190), .ZN(n9235) );
  MUX2_X1 U10326 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9235), .S(n9206), .Z(n9192) );
  AOI21_X1 U10327 ( .B1(n6400), .B2(n9237), .A(n9192), .ZN(n9193) );
  INV_X1 U10328 ( .A(n9193), .ZN(P2_U3478) );
  INV_X1 U10329 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9196) );
  AOI21_X1 U10330 ( .B1(n9204), .B2(n9195), .A(n9194), .ZN(n9239) );
  MUX2_X1 U10331 ( .A(n9196), .B(n9239), .S(n9206), .Z(n9197) );
  OAI21_X1 U10332 ( .B1(n9242), .B2(n9209), .A(n9197), .ZN(P2_U3477) );
  AOI21_X1 U10333 ( .B1(n9199), .B2(n9204), .A(n9198), .ZN(n9243) );
  MUX2_X1 U10334 ( .A(n9200), .B(n9243), .S(n9206), .Z(n9201) );
  OAI21_X1 U10335 ( .B1(n9246), .B2(n9209), .A(n9201), .ZN(P2_U3476) );
  INV_X1 U10336 ( .A(n9202), .ZN(n9205) );
  AOI21_X1 U10337 ( .B1(n9205), .B2(n9204), .A(n9203), .ZN(n9247) );
  MUX2_X1 U10338 ( .A(n9207), .B(n9247), .S(n9206), .Z(n9208) );
  OAI21_X1 U10339 ( .B1(n9251), .B2(n9209), .A(n9208), .ZN(P2_U3475) );
  MUX2_X1 U10340 ( .A(n9211), .B(P2_REG1_REG_0__SCAN_IN), .S(n9210), .Z(
        P2_U3459) );
  NAND2_X1 U10341 ( .A1(n6448), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n9213) );
  NAND2_X1 U10342 ( .A1(n9212), .A2(n11186), .ZN(n9215) );
  OAI211_X1 U10343 ( .C1(n9214), .C2(n9250), .A(n9213), .B(n9215), .ZN(
        P2_U3458) );
  NAND2_X1 U10344 ( .A1(n6448), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n9216) );
  OAI211_X1 U10345 ( .C1(n9217), .C2(n9250), .A(n9216), .B(n9215), .ZN(
        P2_U3457) );
  INV_X1 U10346 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n9220) );
  MUX2_X1 U10347 ( .A(n9220), .B(n9219), .S(n11186), .Z(n9221) );
  OAI21_X1 U10348 ( .B1(n9222), .B2(n9250), .A(n9221), .ZN(P2_U3453) );
  MUX2_X1 U10349 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9223), .S(n11186), .Z(
        P2_U3452) );
  INV_X1 U10350 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n9225) );
  MUX2_X1 U10351 ( .A(n9225), .B(n9224), .S(n11186), .Z(n9226) );
  OAI21_X1 U10352 ( .B1(n9227), .B2(n9250), .A(n9226), .ZN(P2_U3451) );
  MUX2_X1 U10353 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9228), .S(n11186), .Z(
        P2_U3450) );
  MUX2_X1 U10354 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9229), .S(n11186), .Z(
        P2_U3449) );
  MUX2_X1 U10355 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9230), .S(n11186), .Z(
        P2_U3448) );
  INV_X1 U10356 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n9232) );
  MUX2_X1 U10357 ( .A(n9232), .B(n9231), .S(n11186), .Z(n9233) );
  OAI21_X1 U10358 ( .B1(n9234), .B2(n9250), .A(n9233), .ZN(P2_U3447) );
  MUX2_X1 U10359 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9235), .S(n11186), .Z(
        n9236) );
  AOI21_X1 U10360 ( .B1(n6446), .B2(n9237), .A(n9236), .ZN(n9238) );
  INV_X1 U10361 ( .A(n9238), .ZN(P2_U3446) );
  MUX2_X1 U10362 ( .A(n9240), .B(n9239), .S(n11186), .Z(n9241) );
  OAI21_X1 U10363 ( .B1(n9242), .B2(n9250), .A(n9241), .ZN(P2_U3444) );
  INV_X1 U10364 ( .A(P2_REG0_REG_17__SCAN_IN), .ZN(n9244) );
  MUX2_X1 U10365 ( .A(n9244), .B(n9243), .S(n11186), .Z(n9245) );
  OAI21_X1 U10366 ( .B1(n9246), .B2(n9250), .A(n9245), .ZN(P2_U3441) );
  INV_X1 U10367 ( .A(P2_REG0_REG_16__SCAN_IN), .ZN(n9248) );
  MUX2_X1 U10368 ( .A(n9248), .B(n9247), .S(n11186), .Z(n9249) );
  OAI21_X1 U10369 ( .B1(n9251), .B2(n9250), .A(n9249), .ZN(P2_U3438) );
  INV_X1 U10370 ( .A(n9452), .ZN(n9258) );
  INV_X1 U10371 ( .A(n9252), .ZN(n9254) );
  NOR4_X1 U10372 ( .A1(n9254), .A2(P2_IR_REG_30__SCAN_IN), .A3(n9253), .A4(
        P2_U3151), .ZN(n9255) );
  AOI21_X1 U10373 ( .B1(n9256), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9255), .ZN(
        n9257) );
  OAI21_X1 U10374 ( .B1(n9258), .B2(n9262), .A(n9257), .ZN(P2_U3264) );
  OAI222_X1 U10375 ( .A1(n9262), .A2(n9261), .B1(P2_U3151), .B2(n9260), .C1(
        n9259), .C2(n9267), .ZN(P2_U3266) );
  NAND2_X1 U10376 ( .A1(n10519), .A2(n9263), .ZN(n9265) );
  OAI211_X1 U10377 ( .C1(n9267), .C2(n9266), .A(n9265), .B(n9264), .ZN(
        P2_U3267) );
  MUX2_X1 U10378 ( .A(n9268), .B(n10749), .S(P2_STATE_REG_SCAN_IN), .Z(
        P2_U3295) );
  AOI21_X1 U10379 ( .B1(n9375), .B2(n9270), .A(n9269), .ZN(n9271) );
  INV_X1 U10380 ( .A(n9272), .ZN(n10240) );
  INV_X1 U10381 ( .A(n10269), .ZN(n10432) );
  AOI22_X1 U10382 ( .A1(n9394), .A2(n10432), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9273) );
  OAI21_X1 U10383 ( .B1(n10401), .B2(n9391), .A(n9273), .ZN(n9274) );
  AOI21_X1 U10384 ( .B1(n10240), .B2(n9381), .A(n9274), .ZN(n9275) );
  OAI211_X1 U10385 ( .C1(n10419), .C2(n9385), .A(n9276), .B(n9275), .ZN(
        P1_U3214) );
  AOI21_X1 U10386 ( .B1(n9279), .B2(n9277), .A(n9278), .ZN(n9284) );
  AOI22_X1 U10387 ( .A1(n9367), .A2(n10445), .B1(P1_REG3_REG_23__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9281) );
  NAND2_X1 U10388 ( .A1(n9394), .A2(n10463), .ZN(n9280) );
  OAI211_X1 U10389 ( .C1(n9397), .C2(n10293), .A(n9281), .B(n9280), .ZN(n9282)
         );
  AOI21_X1 U10390 ( .B1(n10299), .B2(n9399), .A(n9282), .ZN(n9283) );
  OAI21_X1 U10391 ( .B1(n9284), .B2(n9402), .A(n9283), .ZN(P1_U3216) );
  XOR2_X1 U10392 ( .A(n9286), .B(n9285), .Z(n9291) );
  INV_X1 U10393 ( .A(n9432), .ZN(n10364) );
  NAND2_X1 U10394 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n10162)
         );
  OAI21_X1 U10395 ( .B1(n9391), .B2(n9435), .A(n10162), .ZN(n9287) );
  AOI21_X1 U10396 ( .B1(n9394), .B2(n10364), .A(n9287), .ZN(n9288) );
  OAI21_X1 U10397 ( .B1(n9397), .B2(n10356), .A(n9288), .ZN(n9289) );
  AOI21_X1 U10398 ( .B1(n10478), .B2(n9399), .A(n9289), .ZN(n9290) );
  OAI21_X1 U10399 ( .B1(n9291), .B2(n9402), .A(n9290), .ZN(P1_U3219) );
  AOI22_X1 U10400 ( .A1(n9394), .A2(n10462), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9293) );
  NAND2_X1 U10401 ( .A1(n9367), .A2(n10463), .ZN(n9292) );
  OAI211_X1 U10402 ( .C1(n9397), .C2(n10323), .A(n9293), .B(n9292), .ZN(n9299)
         );
  INV_X1 U10403 ( .A(n9294), .ZN(n9295) );
  AOI211_X1 U10404 ( .C1(n9297), .C2(n9296), .A(n9402), .B(n9295), .ZN(n9298)
         );
  AOI211_X1 U10405 ( .C1(n10331), .C2(n9399), .A(n9299), .B(n9298), .ZN(n9300)
         );
  INV_X1 U10406 ( .A(n9300), .ZN(P1_U3223) );
  OAI21_X1 U10407 ( .B1(n9303), .B2(n9302), .A(n9301), .ZN(n9304) );
  NAND2_X1 U10408 ( .A1(n9304), .A2(n9376), .ZN(n9309) );
  INV_X1 U10409 ( .A(n9305), .ZN(n10266) );
  AOI22_X1 U10410 ( .A1(n9367), .A2(n10432), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9306) );
  OAI21_X1 U10411 ( .B1(n10297), .B2(n9369), .A(n9306), .ZN(n9307) );
  AOI21_X1 U10412 ( .B1(n10266), .B2(n9381), .A(n9307), .ZN(n9308) );
  OAI211_X1 U10413 ( .C1(n10435), .C2(n9385), .A(n9309), .B(n9308), .ZN(
        P1_U3225) );
  NAND2_X1 U10414 ( .A1(n9311), .A2(n9310), .ZN(n9316) );
  INV_X1 U10415 ( .A(n9312), .ZN(n9387) );
  NOR2_X1 U10416 ( .A1(n9389), .A2(n9387), .ZN(n9314) );
  INV_X1 U10417 ( .A(n9389), .ZN(n9313) );
  OAI22_X1 U10418 ( .A1(n9314), .A2(n9386), .B1(n9313), .B2(n9312), .ZN(n9315)
         );
  XOR2_X1 U10419 ( .A(n9316), .B(n9315), .Z(n9324) );
  NOR2_X1 U10420 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9317), .ZN(n10118) );
  NOR2_X1 U10421 ( .A1(n9391), .A2(n10378), .ZN(n9318) );
  AOI211_X1 U10422 ( .C1(n9394), .C2(n9671), .A(n10118), .B(n9318), .ZN(n9319)
         );
  OAI21_X1 U10423 ( .B1(n9397), .B2(n9320), .A(n9319), .ZN(n9321) );
  AOI21_X1 U10424 ( .B1(n9322), .B2(n9399), .A(n9321), .ZN(n9323) );
  OAI21_X1 U10425 ( .B1(n9324), .B2(n9402), .A(n9323), .ZN(P1_U3226) );
  NAND2_X1 U10426 ( .A1(n9327), .A2(n9326), .ZN(n9328) );
  XNOR2_X1 U10427 ( .A(n9325), .B(n9328), .ZN(n9334) );
  NAND2_X1 U10428 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n10143)
         );
  OAI21_X1 U10429 ( .B1(n9369), .B2(n9390), .A(n10143), .ZN(n9329) );
  AOI21_X1 U10430 ( .B1(n9367), .B2(n10364), .A(n9329), .ZN(n9330) );
  OAI21_X1 U10431 ( .B1(n9331), .B2(n9397), .A(n9330), .ZN(n9332) );
  AOI21_X1 U10432 ( .B1(n10488), .B2(n9399), .A(n9332), .ZN(n9333) );
  OAI21_X1 U10433 ( .B1(n9334), .B2(n9402), .A(n9333), .ZN(P1_U3228) );
  INV_X1 U10434 ( .A(n9335), .ZN(n9336) );
  NOR2_X1 U10435 ( .A1(n9337), .A2(n9336), .ZN(n9338) );
  XNOR2_X1 U10436 ( .A(n5179), .B(n9338), .ZN(n9343) );
  AOI22_X1 U10437 ( .A1(n9367), .A2(n10424), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9340) );
  NAND2_X1 U10438 ( .A1(n9394), .A2(n10453), .ZN(n9339) );
  OAI211_X1 U10439 ( .C1(n9397), .C2(n10278), .A(n9340), .B(n9339), .ZN(n9341)
         );
  AOI21_X1 U10440 ( .B1(n10442), .B2(n9399), .A(n9341), .ZN(n9342) );
  OAI21_X1 U10441 ( .B1(n9343), .B2(n9402), .A(n9342), .ZN(P1_U3229) );
  XOR2_X1 U10442 ( .A(n9345), .B(n9344), .Z(n9350) );
  AOI22_X1 U10443 ( .A1(n9367), .A2(n10454), .B1(P1_REG3_REG_20__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9347) );
  INV_X1 U10444 ( .A(n10349), .ZN(n10375) );
  NAND2_X1 U10445 ( .A1(n9394), .A2(n10375), .ZN(n9346) );
  OAI211_X1 U10446 ( .C1(n9397), .C2(n10342), .A(n9347), .B(n9346), .ZN(n9348)
         );
  AOI21_X1 U10447 ( .B1(n10473), .B2(n9399), .A(n9348), .ZN(n9349) );
  OAI21_X1 U10448 ( .B1(n9350), .B2(n9402), .A(n9349), .ZN(P1_U3233) );
  INV_X1 U10449 ( .A(n9277), .ZN(n9357) );
  INV_X1 U10450 ( .A(n9351), .ZN(n9353) );
  NAND2_X1 U10451 ( .A1(n9353), .A2(n9352), .ZN(n9355) );
  AOI22_X1 U10452 ( .A1(n9357), .A2(n9356), .B1(n9355), .B2(n9354), .ZN(n9362)
         );
  AOI22_X1 U10453 ( .A1(n9394), .A2(n10454), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9359) );
  NAND2_X1 U10454 ( .A1(n9367), .A2(n10453), .ZN(n9358) );
  OAI211_X1 U10455 ( .C1(n9397), .C2(n10310), .A(n9359), .B(n9358), .ZN(n9360)
         );
  AOI21_X1 U10456 ( .B1(n10306), .B2(n9399), .A(n9360), .ZN(n9361) );
  OAI21_X1 U10457 ( .B1(n9362), .B2(n9402), .A(n9361), .ZN(P1_U3235) );
  NAND2_X1 U10458 ( .A1(n9364), .A2(n9363), .ZN(n9366) );
  XNOR2_X1 U10459 ( .A(n9366), .B(n9365), .ZN(n9373) );
  NOR2_X1 U10460 ( .A1(n9397), .A2(n10383), .ZN(n9371) );
  NAND2_X1 U10461 ( .A1(n9367), .A2(n10375), .ZN(n9368) );
  NAND2_X1 U10462 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n10731)
         );
  OAI211_X1 U10463 ( .C1(n9369), .C2(n10378), .A(n9368), .B(n10731), .ZN(n9370) );
  AOI211_X1 U10464 ( .C1(n10483), .C2(n9399), .A(n9371), .B(n9370), .ZN(n9372)
         );
  OAI21_X1 U10465 ( .B1(n9373), .B2(n9402), .A(n9372), .ZN(P1_U3238) );
  AND2_X1 U10466 ( .A1(n9301), .A2(n9374), .ZN(n9378) );
  OAI211_X1 U10467 ( .C1(n9378), .C2(n9377), .A(n9376), .B(n9375), .ZN(n9384)
         );
  INV_X1 U10468 ( .A(n10252), .ZN(n9382) );
  AOI22_X1 U10469 ( .A1(n9394), .A2(n10424), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n9379) );
  OAI21_X1 U10470 ( .B1(n10409), .B2(n9391), .A(n9379), .ZN(n9380) );
  AOI21_X1 U10471 ( .B1(n9382), .B2(n9381), .A(n9380), .ZN(n9383) );
  OAI211_X1 U10472 ( .C1(n5490), .C2(n9385), .A(n9384), .B(n9383), .ZN(
        P1_U3240) );
  XNOR2_X1 U10473 ( .A(n9387), .B(n9386), .ZN(n9388) );
  XNOR2_X1 U10474 ( .A(n9389), .B(n9388), .ZN(n9403) );
  NAND2_X1 U10475 ( .A1(P1_U3086), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10719)
         );
  INV_X1 U10476 ( .A(n10719), .ZN(n9393) );
  NOR2_X1 U10477 ( .A1(n9391), .A2(n9390), .ZN(n9392) );
  AOI211_X1 U10478 ( .C1(n9394), .C2(n11170), .A(n9393), .B(n9392), .ZN(n9395)
         );
  OAI21_X1 U10479 ( .B1(n9397), .B2(n9396), .A(n9395), .ZN(n9398) );
  AOI21_X1 U10480 ( .B1(n9400), .B2(n9399), .A(n9398), .ZN(n9401) );
  OAI21_X1 U10481 ( .B1(n9403), .B2(n9402), .A(n9401), .ZN(P1_U3241) );
  NOR3_X1 U10482 ( .A1(n10506), .A2(n10930), .A3(n9404), .ZN(n9668) );
  OAI21_X1 U10483 ( .B1(n9662), .B2(n6792), .A(P1_B_REG_SCAN_IN), .ZN(n9667)
         );
  NAND2_X1 U10484 ( .A1(n9405), .A2(n8029), .ZN(n9408) );
  OR2_X1 U10485 ( .A1(n5139), .A2(n9406), .ZN(n9407) );
  NOR2_X1 U10486 ( .A1(n10398), .A2(n10408), .ZN(n9472) );
  NOR2_X1 U10487 ( .A1(n10412), .A2(n10401), .ZN(n9475) );
  NOR2_X1 U10488 ( .A1(n9472), .A2(n9475), .ZN(n9461) );
  NAND2_X1 U10489 ( .A1(n10412), .A2(n10401), .ZN(n10188) );
  NAND2_X1 U10490 ( .A1(n10244), .A2(n10409), .ZN(n10187) );
  NAND2_X1 U10491 ( .A1(n10188), .A2(n10187), .ZN(n9462) );
  INV_X1 U10492 ( .A(n9462), .ZN(n9445) );
  NAND2_X1 U10493 ( .A1(n10442), .A2(n10297), .ZN(n9622) );
  INV_X1 U10494 ( .A(n10183), .ZN(n10182) );
  NAND2_X1 U10495 ( .A1(n10306), .A2(n10329), .ZN(n10180) );
  AND2_X1 U10496 ( .A1(n10182), .A2(n10180), .ZN(n9620) );
  NAND2_X1 U10497 ( .A1(n9622), .A2(n9620), .ZN(n9502) );
  INV_X1 U10498 ( .A(n9502), .ZN(n9441) );
  NAND2_X1 U10499 ( .A1(n10478), .A2(n10349), .ZN(n9608) );
  NAND2_X1 U10500 ( .A1(n9587), .A2(n9583), .ZN(n9579) );
  NAND2_X1 U10501 ( .A1(n9517), .A2(n9533), .ZN(n9529) );
  INV_X1 U10502 ( .A(n9529), .ZN(n9422) );
  INV_X1 U10503 ( .A(n9542), .ZN(n9411) );
  NAND2_X1 U10504 ( .A1(n7175), .A2(n10982), .ZN(n9478) );
  OAI211_X1 U10505 ( .C1(n10963), .C2(n9409), .A(n9655), .B(n9478), .ZN(n9410)
         );
  NAND3_X1 U10506 ( .A1(n9411), .A2(n9536), .A3(n9410), .ZN(n9413) );
  INV_X1 U10507 ( .A(n9543), .ZN(n9412) );
  AOI21_X1 U10508 ( .B1(n9413), .B2(n9540), .A(n9412), .ZN(n9414) );
  NAND2_X1 U10509 ( .A1(n9546), .A2(n9541), .ZN(n9537) );
  NOR2_X1 U10510 ( .A1(n9414), .A2(n9537), .ZN(n9416) );
  NAND2_X1 U10511 ( .A1(n9415), .A2(n9544), .ZN(n9550) );
  OAI21_X1 U10512 ( .B1(n9416), .B2(n9550), .A(n9552), .ZN(n9417) );
  AOI21_X1 U10513 ( .B1(n9559), .B2(n9417), .A(n9488), .ZN(n9420) );
  INV_X1 U10514 ( .A(n9418), .ZN(n9419) );
  OAI21_X1 U10515 ( .B1(n9420), .B2(n9419), .A(n9568), .ZN(n9421) );
  NAND2_X1 U10516 ( .A1(n9577), .A2(n9522), .ZN(n9520) );
  AOI21_X1 U10517 ( .B1(n9422), .B2(n9421), .A(n9520), .ZN(n9424) );
  AND2_X1 U10518 ( .A1(n9575), .A2(n9518), .ZN(n9581) );
  INV_X1 U10519 ( .A(n9581), .ZN(n9423) );
  NOR2_X1 U10520 ( .A1(n9424), .A2(n9423), .ZN(n9425) );
  NOR2_X1 U10521 ( .A1(n9579), .A2(n9425), .ZN(n9427) );
  AND2_X1 U10522 ( .A1(n9593), .A2(n9585), .ZN(n9578) );
  INV_X1 U10523 ( .A(n9578), .ZN(n9426) );
  OAI21_X1 U10524 ( .B1(n9427), .B2(n9426), .A(n9591), .ZN(n9430) );
  INV_X1 U10525 ( .A(n9595), .ZN(n9429) );
  INV_X1 U10526 ( .A(n9601), .ZN(n9428) );
  AOI211_X1 U10527 ( .C1(n9594), .C2(n9430), .A(n9429), .B(n9428), .ZN(n9433)
         );
  NAND2_X1 U10528 ( .A1(n10483), .A2(n9432), .ZN(n9604) );
  NAND2_X1 U10529 ( .A1(n9604), .A2(n9431), .ZN(n9597) );
  OAI21_X1 U10530 ( .B1(n9433), .B2(n9597), .A(n9602), .ZN(n9434) );
  OR2_X1 U10531 ( .A1(n10478), .A2(n10349), .ZN(n9455) );
  AND2_X1 U10532 ( .A1(n5159), .A2(n9455), .ZN(n9598) );
  AOI21_X1 U10533 ( .B1(n9608), .B2(n9434), .A(n5545), .ZN(n9437) );
  NAND2_X1 U10534 ( .A1(n10331), .A2(n10350), .ZN(n9516) );
  NAND2_X1 U10535 ( .A1(n10473), .A2(n9435), .ZN(n9609) );
  NAND2_X1 U10536 ( .A1(n9516), .A2(n9609), .ZN(n9436) );
  AND2_X1 U10537 ( .A1(n10466), .A2(n10454), .ZN(n9514) );
  OAI21_X1 U10538 ( .B1(n9437), .B2(n9436), .A(n5542), .ZN(n9440) );
  NAND2_X1 U10539 ( .A1(n10448), .A2(n10453), .ZN(n10181) );
  OR2_X1 U10540 ( .A1(n10306), .A2(n10329), .ZN(n9617) );
  AND2_X1 U10541 ( .A1(n10181), .A2(n9617), .ZN(n9513) );
  OAI21_X1 U10542 ( .B1(n9513), .B2(n10183), .A(n10184), .ZN(n9438) );
  AND2_X1 U10543 ( .A1(n10435), .A2(n10424), .ZN(n9476) );
  AOI21_X1 U10544 ( .B1(n9622), .B2(n9438), .A(n9476), .ZN(n9457) );
  INV_X1 U10545 ( .A(n9457), .ZN(n9439) );
  AOI21_X1 U10546 ( .B1(n9441), .B2(n9440), .A(n9439), .ZN(n9443) );
  NAND2_X1 U10547 ( .A1(n10257), .A2(n10269), .ZN(n10186) );
  AND2_X1 U10548 ( .A1(n10186), .A2(n10185), .ZN(n9459) );
  INV_X1 U10549 ( .A(n9459), .ZN(n9627) );
  NAND2_X1 U10550 ( .A1(n9633), .A2(n9628), .ZN(n9458) );
  INV_X1 U10551 ( .A(n9458), .ZN(n9442) );
  OAI21_X1 U10552 ( .B1(n9443), .B2(n9627), .A(n9442), .ZN(n9444) );
  NAND2_X1 U10553 ( .A1(n9445), .A2(n9444), .ZN(n9449) );
  OR2_X1 U10554 ( .A1(n5139), .A2(n10515), .ZN(n9447) );
  NOR2_X1 U10555 ( .A1(n10396), .A2(n10208), .ZN(n9474) );
  NOR2_X1 U10556 ( .A1(n9474), .A2(n9473), .ZN(n9465) );
  INV_X1 U10557 ( .A(n9465), .ZN(n9448) );
  AOI21_X1 U10558 ( .B1(n9461), .B2(n9449), .A(n9448), .ZN(n9453) );
  INV_X1 U10559 ( .A(n10208), .ZN(n9450) );
  OR2_X1 U10560 ( .A1(n10176), .A2(n9450), .ZN(n9467) );
  INV_X1 U10561 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n10510) );
  NOR2_X1 U10562 ( .A1(n5138), .A2(n10510), .ZN(n9451) );
  INV_X1 U10563 ( .A(n10393), .ZN(n10171) );
  INV_X1 U10564 ( .A(n10170), .ZN(n9466) );
  AND2_X1 U10565 ( .A1(n10393), .A2(n10170), .ZN(n9507) );
  INV_X1 U10566 ( .A(n9507), .ZN(n9649) );
  OAI21_X1 U10567 ( .B1(n9453), .B2(n9506), .A(n9649), .ZN(n9665) );
  NAND2_X1 U10568 ( .A1(n9454), .A2(n9601), .ZN(n10374) );
  OAI21_X1 U10569 ( .B1(n10179), .B2(n9502), .A(n9457), .ZN(n9460) );
  AOI21_X1 U10570 ( .B1(n9460), .B2(n9459), .A(n9458), .ZN(n9463) );
  OAI21_X1 U10571 ( .B1(n9463), .B2(n9462), .A(n9461), .ZN(n9464) );
  OAI211_X1 U10572 ( .C1(n10396), .C2(n10170), .A(n9465), .B(n9464), .ZN(n9468) );
  AOI21_X1 U10573 ( .B1(n9468), .B2(n9642), .A(n9507), .ZN(n9471) );
  INV_X1 U10574 ( .A(n9643), .ZN(n9470) );
  NOR3_X1 U10575 ( .A1(n9471), .A2(n9470), .A3(n9469), .ZN(n9508) );
  INV_X1 U10576 ( .A(n9472), .ZN(n9509) );
  NAND2_X1 U10577 ( .A1(n9509), .A2(n9510), .ZN(n10203) );
  INV_X1 U10578 ( .A(n9474), .ZN(n9504) );
  INV_X1 U10579 ( .A(n9475), .ZN(n9636) );
  NAND2_X1 U10580 ( .A1(n5159), .A2(n9609), .ZN(n10337) );
  INV_X1 U10581 ( .A(n10362), .ZN(n9499) );
  INV_X1 U10582 ( .A(n10985), .ZN(n9479) );
  INV_X1 U10583 ( .A(n9477), .ZN(n10986) );
  NAND2_X1 U10584 ( .A1(n10986), .A2(n9478), .ZN(n10976) );
  NOR4_X1 U10585 ( .A1(n9479), .A2(n7179), .A3(n10976), .A4(n9655), .ZN(n9485)
         );
  NOR4_X1 U10586 ( .A1(n9483), .A2(n9482), .A3(n9481), .A4(n9480), .ZN(n9484)
         );
  NAND4_X1 U10587 ( .A1(n9526), .A2(n9486), .A3(n9485), .A4(n9484), .ZN(n9487)
         );
  OR4_X1 U10588 ( .A1(n9490), .A2(n9489), .A3(n9488), .A4(n9487), .ZN(n9491)
         );
  NOR4_X1 U10589 ( .A1(n9494), .A2(n9493), .A3(n9492), .A4(n9491), .ZN(n9495)
         );
  NAND4_X1 U10590 ( .A1(n10191), .A2(n9497), .A3(n9496), .A4(n9495), .ZN(n9498) );
  NOR4_X1 U10591 ( .A1(n10337), .A2(n10370), .A3(n9499), .A4(n9498), .ZN(n9500) );
  NAND4_X1 U10592 ( .A1(n9513), .A2(n10184), .A3(n10319), .A4(n9500), .ZN(
        n9501) );
  NOR4_X1 U10593 ( .A1(n10249), .A2(n10262), .A3(n9502), .A4(n9501), .ZN(n9503) );
  NAND4_X1 U10594 ( .A1(n9504), .A2(n10236), .A3(n10220), .A4(n9503), .ZN(
        n9505) );
  OAI21_X1 U10595 ( .B1(n9508), .B2(n9654), .A(n10163), .ZN(n9661) );
  AND2_X1 U10596 ( .A1(n9647), .A2(n10158), .ZN(n9644) );
  INV_X1 U10597 ( .A(n9644), .ZN(n9640) );
  MUX2_X1 U10598 ( .A(n9510), .B(n9509), .S(n9640), .Z(n9638) );
  AND2_X1 U10599 ( .A1(n10185), .A2(n9622), .ZN(n9512) );
  NOR2_X1 U10600 ( .A1(n10262), .A2(n5539), .ZN(n9511) );
  MUX2_X1 U10601 ( .A(n9512), .B(n9511), .S(n9644), .Z(n9626) );
  INV_X1 U10602 ( .A(n9513), .ZN(n9616) );
  NOR2_X1 U10603 ( .A1(n9616), .A2(n9514), .ZN(n9515) );
  MUX2_X1 U10604 ( .A(n9516), .B(n9515), .S(n9644), .Z(n9615) );
  NAND2_X1 U10605 ( .A1(n9518), .A2(n9517), .ZN(n9519) );
  MUX2_X1 U10606 ( .A(n9520), .B(n9519), .S(n9644), .Z(n9521) );
  INV_X1 U10607 ( .A(n9521), .ZN(n9574) );
  INV_X1 U10608 ( .A(n9533), .ZN(n9524) );
  OAI211_X1 U10609 ( .C1(n9524), .C2(n9523), .A(n9522), .B(n9568), .ZN(n9525)
         );
  INV_X1 U10610 ( .A(n9525), .ZN(n9531) );
  INV_X1 U10611 ( .A(n9526), .ZN(n9527) );
  AND2_X1 U10612 ( .A1(n9568), .A2(n9527), .ZN(n9528) );
  NOR2_X1 U10613 ( .A1(n9529), .A2(n9528), .ZN(n9530) );
  MUX2_X1 U10614 ( .A(n9531), .B(n9530), .S(n9640), .Z(n9572) );
  AND2_X1 U10615 ( .A1(n9533), .A2(n9532), .ZN(n9534) );
  MUX2_X1 U10616 ( .A(n9535), .B(n9534), .S(n9644), .Z(n9570) );
  AND2_X1 U10617 ( .A1(n9543), .A2(n9536), .ZN(n9538) );
  AOI21_X1 U10618 ( .B1(n9539), .B2(n9538), .A(n9537), .ZN(n9549) );
  OAI211_X1 U10619 ( .C1(n9542), .C2(n7179), .A(n9541), .B(n9540), .ZN(n9545)
         );
  NAND3_X1 U10620 ( .A1(n9545), .A2(n9544), .A3(n9543), .ZN(n9547) );
  NAND2_X1 U10621 ( .A1(n9547), .A2(n9546), .ZN(n9548) );
  MUX2_X1 U10622 ( .A(n9549), .B(n9548), .S(n9644), .Z(n9558) );
  NAND2_X1 U10623 ( .A1(n9550), .A2(n9552), .ZN(n9551) );
  MUX2_X1 U10624 ( .A(n9552), .B(n9551), .S(n9640), .Z(n9555) );
  NAND3_X1 U10625 ( .A1(n9555), .A2(n9554), .A3(n9553), .ZN(n9556) );
  AOI21_X1 U10626 ( .B1(n9558), .B2(n9557), .A(n9556), .ZN(n9566) );
  OAI21_X1 U10627 ( .B1(n9562), .B2(n9559), .A(n11102), .ZN(n9564) );
  OAI21_X1 U10628 ( .B1(n9562), .B2(n9561), .A(n9560), .ZN(n9563) );
  MUX2_X1 U10629 ( .A(n9564), .B(n9563), .S(n9640), .Z(n9565) );
  OAI21_X1 U10630 ( .B1(n9566), .B2(n9565), .A(n11101), .ZN(n9567) );
  NAND4_X1 U10631 ( .A1(n9570), .A2(n9569), .A3(n9568), .A4(n9567), .ZN(n9571)
         );
  NAND2_X1 U10632 ( .A1(n9572), .A2(n9571), .ZN(n9573) );
  NAND2_X1 U10633 ( .A1(n9574), .A2(n9573), .ZN(n9582) );
  INV_X1 U10634 ( .A(n9575), .ZN(n9576) );
  AOI21_X1 U10635 ( .B1(n9582), .B2(n9577), .A(n9576), .ZN(n9580) );
  OAI211_X1 U10636 ( .C1(n9580), .C2(n9579), .A(n9578), .B(n9644), .ZN(n9590)
         );
  NAND2_X1 U10637 ( .A1(n9582), .A2(n9581), .ZN(n9584) );
  NAND2_X1 U10638 ( .A1(n9584), .A2(n9583), .ZN(n9586) );
  NAND2_X1 U10639 ( .A1(n9586), .A2(n9585), .ZN(n9588) );
  NAND4_X1 U10640 ( .A1(n9588), .A2(n9587), .A3(n9591), .A4(n9640), .ZN(n9589)
         );
  NAND2_X1 U10641 ( .A1(n9595), .A2(n9591), .ZN(n9592) );
  NAND2_X1 U10642 ( .A1(n9594), .A2(n9593), .ZN(n9596) );
  OAI211_X1 U10643 ( .C1(n9600), .C2(n9597), .A(n10362), .B(n9602), .ZN(n9599)
         );
  MUX2_X1 U10644 ( .A(n9599), .B(n9598), .S(n9644), .Z(n9607) );
  INV_X1 U10645 ( .A(n9600), .ZN(n9603) );
  NAND3_X1 U10646 ( .A1(n9603), .A2(n9602), .A3(n9601), .ZN(n9605) );
  NAND4_X1 U10647 ( .A1(n9605), .A2(n9644), .A3(n9604), .A4(n9608), .ZN(n9606)
         );
  AOI21_X1 U10648 ( .B1(n9607), .B2(n9606), .A(n9456), .ZN(n9613) );
  AOI21_X1 U10649 ( .B1(n9609), .B2(n9608), .A(n9644), .ZN(n9612) );
  NOR2_X1 U10650 ( .A1(n5159), .A2(n9644), .ZN(n9610) );
  NOR2_X1 U10651 ( .A1(n10321), .A2(n9610), .ZN(n9611) );
  OAI21_X1 U10652 ( .B1(n9613), .B2(n9612), .A(n9611), .ZN(n9614) );
  NAND2_X1 U10653 ( .A1(n9616), .A2(n9644), .ZN(n9618) );
  AOI21_X1 U10654 ( .B1(n9618), .B2(n10304), .A(n10183), .ZN(n9619) );
  INV_X1 U10655 ( .A(n9620), .ZN(n9621) );
  NOR2_X1 U10656 ( .A1(n9623), .A2(n9644), .ZN(n9624) );
  AOI21_X1 U10657 ( .B1(n9626), .B2(n9625), .A(n9624), .ZN(n9631) );
  NAND2_X1 U10658 ( .A1(n9627), .A2(n9644), .ZN(n9629) );
  MUX2_X1 U10659 ( .A(n9644), .B(n9629), .S(n9628), .Z(n9630) );
  OAI21_X1 U10660 ( .B1(n9631), .B2(n10249), .A(n9630), .ZN(n9632) );
  NAND2_X1 U10661 ( .A1(n9632), .A2(n10236), .ZN(n9635) );
  MUX2_X1 U10662 ( .A(n10187), .B(n9633), .S(n9640), .Z(n9634) );
  MUX2_X1 U10663 ( .A(n10188), .B(n9636), .S(n9644), .Z(n9637) );
  NAND2_X1 U10664 ( .A1(n10208), .A2(n10170), .ZN(n9639) );
  NAND3_X1 U10665 ( .A1(n10176), .A2(n9640), .A3(n9639), .ZN(n9641) );
  NAND2_X1 U10666 ( .A1(n9643), .A2(n9642), .ZN(n9645) );
  NAND2_X1 U10667 ( .A1(n9645), .A2(n9644), .ZN(n9646) );
  NAND2_X1 U10668 ( .A1(n9647), .A2(n9655), .ZN(n9657) );
  INV_X1 U10669 ( .A(n9657), .ZN(n9648) );
  INV_X1 U10670 ( .A(n9654), .ZN(n9660) );
  NAND2_X1 U10671 ( .A1(n9656), .A2(n9655), .ZN(n9659) );
  AOI21_X1 U10672 ( .B1(n9665), .B2(n9663), .A(n9662), .ZN(n9664) );
  MUX2_X1 U10673 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(n10416), .S(n10937), .Z(
        P1_U3582) );
  MUX2_X1 U10674 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n10425), .S(n10937), .Z(
        P1_U3581) );
  MUX2_X1 U10675 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n10432), .S(n10937), .Z(
        P1_U3580) );
  MUX2_X1 U10676 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n10424), .S(P1_U3973), .Z(
        P1_U3579) );
  MUX2_X1 U10677 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n10445), .S(n10937), .Z(
        P1_U3578) );
  MUX2_X1 U10678 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n10463), .S(P1_U3973), .Z(
        P1_U3576) );
  MUX2_X1 U10679 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n10454), .S(n10937), .Z(
        P1_U3575) );
  MUX2_X1 U10680 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n10462), .S(P1_U3973), .Z(
        P1_U3574) );
  MUX2_X1 U10681 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n10375), .S(P1_U3973), .Z(
        P1_U3573) );
  MUX2_X1 U10682 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n10364), .S(P1_U3973), .Z(
        P1_U3572) );
  MUX2_X1 U10683 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9670), .S(P1_U3973), .Z(
        P1_U3570) );
  MUX2_X1 U10684 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9671), .S(P1_U3973), .Z(
        P1_U3569) );
  MUX2_X1 U10685 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n11170), .S(P1_U3973), .Z(
        P1_U3568) );
  MUX2_X1 U10686 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9672), .S(P1_U3973), .Z(
        P1_U3567) );
  MUX2_X1 U10687 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n11171), .S(P1_U3973), .Z(
        P1_U3566) );
  MUX2_X1 U10688 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n11146), .S(P1_U3973), .Z(
        P1_U3565) );
  MUX2_X1 U10689 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n9673), .S(P1_U3973), .Z(
        P1_U3563) );
  MUX2_X1 U10690 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n11136), .S(P1_U3973), .Z(
        P1_U3562) );
  MUX2_X1 U10691 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n11065), .S(P1_U3973), .Z(
        P1_U3561) );
  MUX2_X1 U10692 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9674), .S(P1_U3973), .Z(
        P1_U3560) );
  MUX2_X1 U10693 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n11064), .S(P1_U3973), .Z(
        P1_U3559) );
  MUX2_X1 U10694 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n11019), .S(P1_U3973), .Z(
        P1_U3558) );
  MUX2_X1 U10695 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n5142), .S(P1_U3973), .Z(
        P1_U3557) );
  MUX2_X1 U10696 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n11020), .S(P1_U3973), .Z(
        P1_U3556) );
  MUX2_X1 U10697 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n11007), .S(n10937), .Z(
        P1_U3555) );
  MUX2_X1 U10698 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n7175), .S(n10937), .Z(
        P1_U3554) );
  XNOR2_X1 U10699 ( .A(n9676), .B(n9675), .ZN(n9686) );
  AOI22_X1 U10700 ( .A1(n10942), .A2(P1_ADDR_REG_10__SCAN_IN), .B1(
        P1_REG3_REG_10__SCAN_IN), .B2(P1_U3086), .ZN(n9682) );
  XOR2_X1 U10701 ( .A(n9679), .B(n9678), .Z(n9680) );
  NAND2_X1 U10702 ( .A1(n10954), .A2(n9680), .ZN(n9681) );
  OAI211_X1 U10703 ( .C1(n10949), .C2(n9683), .A(n9682), .B(n9681), .ZN(n9684)
         );
  AOI21_X1 U10704 ( .B1(n9686), .B2(n9685), .A(n9684), .ZN(n10110) );
  XNOR2_X1 U10705 ( .A(n9687), .B(keyinput_3), .ZN(n9700) );
  XNOR2_X1 U10706 ( .A(SI_31_), .B(keyinput_1), .ZN(n9690) );
  XNOR2_X1 U10707 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_0), .ZN(n9689) );
  XNOR2_X1 U10708 ( .A(SI_30_), .B(keyinput_2), .ZN(n9688) );
  OAI21_X1 U10709 ( .B1(n9690), .B2(n9689), .A(n9688), .ZN(n9699) );
  XNOR2_X1 U10710 ( .A(SI_25_), .B(keyinput_7), .ZN(n9692) );
  XNOR2_X1 U10711 ( .A(SI_28_), .B(keyinput_4), .ZN(n9691) );
  NOR2_X1 U10712 ( .A1(n9692), .A2(n9691), .ZN(n9697) );
  XNOR2_X1 U10713 ( .A(n9693), .B(keyinput_6), .ZN(n9696) );
  XNOR2_X1 U10714 ( .A(n9893), .B(keyinput_5), .ZN(n9695) );
  XNOR2_X1 U10715 ( .A(SI_24_), .B(keyinput_8), .ZN(n9694) );
  NAND4_X1 U10716 ( .A1(n9697), .A2(n9696), .A3(n9695), .A4(n9694), .ZN(n9698)
         );
  AOI21_X1 U10717 ( .B1(n9700), .B2(n9699), .A(n9698), .ZN(n9705) );
  XNOR2_X1 U10718 ( .A(n9701), .B(keyinput_9), .ZN(n9704) );
  XNOR2_X1 U10719 ( .A(n9702), .B(keyinput_10), .ZN(n9703) );
  OAI21_X1 U10720 ( .B1(n9705), .B2(n9704), .A(n9703), .ZN(n9710) );
  XNOR2_X1 U10721 ( .A(n9706), .B(keyinput_12), .ZN(n9709) );
  XNOR2_X1 U10722 ( .A(SI_21_), .B(keyinput_11), .ZN(n9708) );
  XNOR2_X1 U10723 ( .A(SI_19_), .B(keyinput_13), .ZN(n9707) );
  NAND4_X1 U10724 ( .A1(n9710), .A2(n9709), .A3(n9708), .A4(n9707), .ZN(n9713)
         );
  XNOR2_X1 U10725 ( .A(n9913), .B(keyinput_15), .ZN(n9712) );
  XNOR2_X1 U10726 ( .A(SI_18_), .B(keyinput_14), .ZN(n9711) );
  NAND3_X1 U10727 ( .A1(n9713), .A2(n9712), .A3(n9711), .ZN(n9720) );
  XNOR2_X1 U10728 ( .A(SI_16_), .B(keyinput_16), .ZN(n9719) );
  XNOR2_X1 U10729 ( .A(n9714), .B(keyinput_18), .ZN(n9717) );
  XNOR2_X1 U10730 ( .A(SI_13_), .B(keyinput_19), .ZN(n9716) );
  XNOR2_X1 U10731 ( .A(SI_15_), .B(keyinput_17), .ZN(n9715) );
  NAND3_X1 U10732 ( .A1(n9717), .A2(n9716), .A3(n9715), .ZN(n9718) );
  AOI21_X1 U10733 ( .B1(n9720), .B2(n9719), .A(n9718), .ZN(n9724) );
  XOR2_X1 U10734 ( .A(SI_12_), .B(keyinput_20), .Z(n9723) );
  XNOR2_X1 U10735 ( .A(n9923), .B(keyinput_22), .ZN(n9722) );
  XOR2_X1 U10736 ( .A(SI_11_), .B(keyinput_21), .Z(n9721) );
  OAI211_X1 U10737 ( .C1(n9724), .C2(n9723), .A(n9722), .B(n9721), .ZN(n9728)
         );
  XNOR2_X1 U10738 ( .A(n9725), .B(keyinput_24), .ZN(n9727) );
  XNOR2_X1 U10739 ( .A(SI_9_), .B(keyinput_23), .ZN(n9726) );
  NAND3_X1 U10740 ( .A1(n9728), .A2(n9727), .A3(n9726), .ZN(n9732) );
  XNOR2_X1 U10741 ( .A(n9932), .B(keyinput_25), .ZN(n9731) );
  XNOR2_X1 U10742 ( .A(n9729), .B(keyinput_26), .ZN(n9730) );
  AOI21_X1 U10743 ( .B1(n9732), .B2(n9731), .A(n9730), .ZN(n9741) );
  XNOR2_X1 U10744 ( .A(SI_5_), .B(keyinput_27), .ZN(n9740) );
  XOR2_X1 U10745 ( .A(SI_2_), .B(keyinput_30), .Z(n9735) );
  XNOR2_X1 U10746 ( .A(SI_0_), .B(keyinput_32), .ZN(n9734) );
  XNOR2_X1 U10747 ( .A(SI_4_), .B(keyinput_28), .ZN(n9733) );
  NAND3_X1 U10748 ( .A1(n9735), .A2(n9734), .A3(n9733), .ZN(n9738) );
  XNOR2_X1 U10749 ( .A(n9936), .B(keyinput_29), .ZN(n9737) );
  XNOR2_X1 U10750 ( .A(SI_1_), .B(keyinput_31), .ZN(n9736) );
  NOR3_X1 U10751 ( .A1(n9738), .A2(n9737), .A3(n9736), .ZN(n9739) );
  OAI21_X1 U10752 ( .B1(n9741), .B2(n9740), .A(n9739), .ZN(n9744) );
  XNOR2_X1 U10753 ( .A(P2_U3151), .B(keyinput_34), .ZN(n9743) );
  XNOR2_X1 U10754 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_33), .ZN(n9742) );
  NAND3_X1 U10755 ( .A1(n9744), .A2(n9743), .A3(n9742), .ZN(n9748) );
  XNOR2_X1 U10756 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_36), .ZN(n9747)
         );
  XNOR2_X1 U10757 ( .A(P2_REG3_REG_7__SCAN_IN), .B(keyinput_35), .ZN(n9746) );
  XNOR2_X1 U10758 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_37), .ZN(n9745)
         );
  NAND4_X1 U10759 ( .A1(n9748), .A2(n9747), .A3(n9746), .A4(n9745), .ZN(n9751)
         );
  XNOR2_X1 U10760 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_38), .ZN(n9750)
         );
  XNOR2_X1 U10761 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_39), .ZN(n9749)
         );
  AOI21_X1 U10762 ( .B1(n9751), .B2(n9750), .A(n9749), .ZN(n9755) );
  XNOR2_X1 U10763 ( .A(n9752), .B(keyinput_41), .ZN(n9754) );
  XNOR2_X1 U10764 ( .A(P2_REG3_REG_3__SCAN_IN), .B(keyinput_40), .ZN(n9753) );
  NOR3_X1 U10765 ( .A1(n9755), .A2(n9754), .A3(n9753), .ZN(n9758) );
  XNOR2_X1 U10766 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n9757)
         );
  XNOR2_X1 U10767 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_43), .ZN(n9756) );
  OAI21_X1 U10768 ( .B1(n9758), .B2(n9757), .A(n9756), .ZN(n9766) );
  XOR2_X1 U10769 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_44), .Z(n9765) );
  XOR2_X1 U10770 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_48), .Z(n9763) );
  XNOR2_X1 U10771 ( .A(n9759), .B(keyinput_47), .ZN(n9762) );
  XNOR2_X1 U10772 ( .A(n9966), .B(keyinput_45), .ZN(n9761) );
  XNOR2_X1 U10773 ( .A(P2_REG3_REG_12__SCAN_IN), .B(keyinput_46), .ZN(n9760)
         );
  NAND4_X1 U10774 ( .A1(n9763), .A2(n9762), .A3(n9761), .A4(n9760), .ZN(n9764)
         );
  AOI21_X1 U10775 ( .B1(n9766), .B2(n9765), .A(n9764), .ZN(n9770) );
  XNOR2_X1 U10776 ( .A(P2_REG3_REG_5__SCAN_IN), .B(keyinput_49), .ZN(n9769) );
  XNOR2_X1 U10777 ( .A(n9767), .B(keyinput_50), .ZN(n9768) );
  OAI21_X1 U10778 ( .B1(n9770), .B2(n9769), .A(n9768), .ZN(n9773) );
  XNOR2_X1 U10779 ( .A(n9979), .B(keyinput_51), .ZN(n9772) );
  XNOR2_X1 U10780 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_52), .ZN(n9771) );
  AOI21_X1 U10781 ( .B1(n9773), .B2(n9772), .A(n9771), .ZN(n9781) );
  XNOR2_X1 U10782 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput_53), .ZN(n9780) );
  INV_X1 U10783 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n9987) );
  AOI22_X1 U10784 ( .A1(n9987), .A2(keyinput_55), .B1(keyinput_58), .B2(n9984), 
        .ZN(n9774) );
  OAI221_X1 U10785 ( .B1(n9987), .B2(keyinput_55), .C1(n9984), .C2(keyinput_58), .A(n9774), .ZN(n9778) );
  INV_X1 U10786 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n9986) );
  AOI22_X1 U10787 ( .A1(n5738), .A2(keyinput_56), .B1(n9986), .B2(keyinput_57), 
        .ZN(n9775) );
  OAI221_X1 U10788 ( .B1(n5738), .B2(keyinput_56), .C1(n9986), .C2(keyinput_57), .A(n9775), .ZN(n9777) );
  XNOR2_X1 U10789 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_54), .ZN(n9776) );
  NOR3_X1 U10790 ( .A1(n9778), .A2(n9777), .A3(n9776), .ZN(n9779) );
  OAI21_X1 U10791 ( .B1(n9781), .B2(n9780), .A(n9779), .ZN(n9784) );
  XNOR2_X1 U10792 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_59), .ZN(n9783) );
  XOR2_X1 U10793 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_60), .Z(n9782) );
  AOI21_X1 U10794 ( .B1(n9784), .B2(n9783), .A(n9782), .ZN(n9793) );
  XOR2_X1 U10795 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_61), .Z(n9792) );
  INV_X1 U10796 ( .A(P2_B_REG_SCAN_IN), .ZN(n9786) );
  AOI22_X1 U10797 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(keyinput_63), .B1(n9786), 
        .B2(keyinput_64), .ZN(n9785) );
  OAI221_X1 U10798 ( .B1(P2_REG3_REG_15__SCAN_IN), .B2(keyinput_63), .C1(n9786), .C2(keyinput_64), .A(n9785), .ZN(n9790) );
  AOI22_X1 U10799 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(keyinput_65), .B1(
        n10515), .B2(keyinput_66), .ZN(n9787) );
  OAI221_X1 U10800 ( .B1(P2_DATAO_REG_31__SCAN_IN), .B2(keyinput_65), .C1(
        n10515), .C2(keyinput_66), .A(n9787), .ZN(n9789) );
  XNOR2_X1 U10801 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_62), .ZN(n9788)
         );
  NOR3_X1 U10802 ( .A1(n9790), .A2(n9789), .A3(n9788), .ZN(n9791) );
  OAI21_X1 U10803 ( .B1(n9793), .B2(n9792), .A(n9791), .ZN(n9796) );
  XNOR2_X1 U10804 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_67), .ZN(n9795)
         );
  XNOR2_X1 U10805 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_68), .ZN(n9794)
         );
  AOI21_X1 U10806 ( .B1(n9796), .B2(n9795), .A(n9794), .ZN(n9800) );
  XNOR2_X1 U10807 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_69), .ZN(n9799)
         );
  XNOR2_X1 U10808 ( .A(n9797), .B(keyinput_70), .ZN(n9798) );
  OAI21_X1 U10809 ( .B1(n9800), .B2(n9799), .A(n9798), .ZN(n9804) );
  XNOR2_X1 U10810 ( .A(n9801), .B(keyinput_72), .ZN(n9803) );
  XNOR2_X1 U10811 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(keyinput_71), .ZN(n9802)
         );
  NAND3_X1 U10812 ( .A1(n9804), .A2(n9803), .A3(n9802), .ZN(n9808) );
  XNOR2_X1 U10813 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(keyinput_73), .ZN(n9807)
         );
  XNOR2_X1 U10814 ( .A(n9805), .B(keyinput_74), .ZN(n9806) );
  AOI21_X1 U10815 ( .B1(n9808), .B2(n9807), .A(n9806), .ZN(n9811) );
  XOR2_X1 U10816 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_75), .Z(n9810) );
  XNOR2_X1 U10817 ( .A(n10021), .B(keyinput_76), .ZN(n9809) );
  NOR3_X1 U10818 ( .A1(n9811), .A2(n9810), .A3(n9809), .ZN(n9817) );
  XNOR2_X1 U10819 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_77), .ZN(n9816)
         );
  XOR2_X1 U10820 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_78), .Z(n9814) );
  XNOR2_X1 U10821 ( .A(n10025), .B(keyinput_80), .ZN(n9813) );
  XNOR2_X1 U10822 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_79), .ZN(n9812)
         );
  NOR3_X1 U10823 ( .A1(n9814), .A2(n9813), .A3(n9812), .ZN(n9815) );
  OAI21_X1 U10824 ( .B1(n9817), .B2(n9816), .A(n9815), .ZN(n9825) );
  XOR2_X1 U10825 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_81), .Z(n9821) );
  XNOR2_X1 U10826 ( .A(n10032), .B(keyinput_82), .ZN(n9820) );
  XNOR2_X1 U10827 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_84), .ZN(n9819)
         );
  XNOR2_X1 U10828 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_83), .ZN(n9818)
         );
  NOR4_X1 U10829 ( .A1(n9821), .A2(n9820), .A3(n9819), .A4(n9818), .ZN(n9824)
         );
  XOR2_X1 U10830 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_86), .Z(n9823) );
  XOR2_X1 U10831 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_85), .Z(n9822) );
  AOI211_X1 U10832 ( .C1(n9825), .C2(n9824), .A(n9823), .B(n9822), .ZN(n9828)
         );
  XOR2_X1 U10833 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_88), .Z(n9827) );
  XNOR2_X1 U10834 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_87), .ZN(n9826)
         );
  NOR3_X1 U10835 ( .A1(n9828), .A2(n9827), .A3(n9826), .ZN(n9831) );
  XNOR2_X1 U10836 ( .A(n5247), .B(keyinput_90), .ZN(n9830) );
  XNOR2_X1 U10837 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_89), .ZN(n9829)
         );
  NOR3_X1 U10838 ( .A1(n9831), .A2(n9830), .A3(n9829), .ZN(n9839) );
  XNOR2_X1 U10839 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_94), .ZN(n9838) );
  XNOR2_X1 U10840 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_95), .ZN(n9837) );
  XNOR2_X1 U10841 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_96), .ZN(n9835) );
  XNOR2_X1 U10842 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_93), .ZN(n9834) );
  XNOR2_X1 U10843 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_92), .ZN(n9833) );
  XNOR2_X1 U10844 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_91), .ZN(n9832) );
  NAND4_X1 U10845 ( .A1(n9835), .A2(n9834), .A3(n9833), .A4(n9832), .ZN(n9836)
         );
  NOR4_X1 U10846 ( .A1(n9839), .A2(n9838), .A3(n9837), .A4(n9836), .ZN(n9842)
         );
  XNOR2_X1 U10847 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_97), .ZN(n9841) );
  XNOR2_X1 U10848 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_98), .ZN(n9840) );
  NOR3_X1 U10849 ( .A1(n9842), .A2(n9841), .A3(n9840), .ZN(n9845) );
  XNOR2_X1 U10850 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_99), .ZN(n9844) );
  XNOR2_X1 U10851 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_100), .ZN(n9843) );
  NOR3_X1 U10852 ( .A1(n9845), .A2(n9844), .A3(n9843), .ZN(n9867) );
  XOR2_X1 U10853 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_103), .Z(n9850) );
  XNOR2_X1 U10854 ( .A(n10061), .B(keyinput_101), .ZN(n9849) );
  XNOR2_X1 U10855 ( .A(n9846), .B(keyinput_102), .ZN(n9848) );
  XNOR2_X1 U10856 ( .A(P1_IR_REG_14__SCAN_IN), .B(keyinput_104), .ZN(n9847) );
  NAND4_X1 U10857 ( .A1(n9850), .A2(n9849), .A3(n9848), .A4(n9847), .ZN(n9866)
         );
  OAI22_X1 U10858 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(keyinput_106), .B1(
        P1_IR_REG_20__SCAN_IN), .B2(keyinput_110), .ZN(n9851) );
  AOI221_X1 U10859 ( .B1(P1_IR_REG_16__SCAN_IN), .B2(keyinput_106), .C1(
        keyinput_110), .C2(P1_IR_REG_20__SCAN_IN), .A(n9851), .ZN(n9865) );
  OAI22_X1 U10860 ( .A1(n9853), .A2(keyinput_105), .B1(P1_IR_REG_21__SCAN_IN), 
        .B2(keyinput_111), .ZN(n9852) );
  AOI221_X1 U10861 ( .B1(n9853), .B2(keyinput_105), .C1(keyinput_111), .C2(
        P1_IR_REG_21__SCAN_IN), .A(n9852), .ZN(n9854) );
  INV_X1 U10862 ( .A(n9854), .ZN(n9863) );
  XNOR2_X1 U10863 ( .A(P1_IR_REG_23__SCAN_IN), .B(keyinput_113), .ZN(n9862) );
  XNOR2_X1 U10864 ( .A(P1_IR_REG_17__SCAN_IN), .B(keyinput_107), .ZN(n9861) );
  INV_X1 U10865 ( .A(keyinput_108), .ZN(n9855) );
  XNOR2_X1 U10866 ( .A(n9855), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9859) );
  INV_X1 U10867 ( .A(keyinput_112), .ZN(n9856) );
  XNOR2_X1 U10868 ( .A(n9856), .B(P1_IR_REG_22__SCAN_IN), .ZN(n9858) );
  XNOR2_X1 U10869 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_109), .ZN(n9857) );
  NAND3_X1 U10870 ( .A1(n9859), .A2(n9858), .A3(n9857), .ZN(n9860) );
  NOR4_X1 U10871 ( .A1(n9863), .A2(n9862), .A3(n9861), .A4(n9860), .ZN(n9864)
         );
  OAI211_X1 U10872 ( .C1(n9867), .C2(n9866), .A(n9865), .B(n9864), .ZN(n9871)
         );
  XNOR2_X1 U10873 ( .A(P1_IR_REG_24__SCAN_IN), .B(keyinput_114), .ZN(n9870) );
  XNOR2_X1 U10874 ( .A(n10083), .B(keyinput_115), .ZN(n9869) );
  XNOR2_X1 U10875 ( .A(P1_IR_REG_26__SCAN_IN), .B(keyinput_116), .ZN(n9868) );
  AOI211_X1 U10876 ( .C1(n9871), .C2(n9870), .A(n9869), .B(n9868), .ZN(n9874)
         );
  XNOR2_X1 U10877 ( .A(n10089), .B(keyinput_118), .ZN(n9873) );
  XNOR2_X1 U10878 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_117), .ZN(n9872) );
  NOR3_X1 U10879 ( .A1(n9874), .A2(n9873), .A3(n9872), .ZN(n9877) );
  XNOR2_X1 U10880 ( .A(n10093), .B(keyinput_119), .ZN(n9876) );
  INV_X1 U10881 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n10509) );
  XNOR2_X1 U10882 ( .A(n10509), .B(keyinput_120), .ZN(n9875) );
  NOR3_X1 U10883 ( .A1(n9877), .A2(n9876), .A3(n9875), .ZN(n9885) );
  INV_X1 U10884 ( .A(keyinput_121), .ZN(n9878) );
  XNOR2_X1 U10885 ( .A(n9878), .B(P1_IR_REG_31__SCAN_IN), .ZN(n9882) );
  XNOR2_X1 U10886 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_123), .ZN(n9881) );
  XNOR2_X1 U10887 ( .A(P1_D_REG_0__SCAN_IN), .B(keyinput_122), .ZN(n9880) );
  XNOR2_X1 U10888 ( .A(P1_D_REG_2__SCAN_IN), .B(keyinput_124), .ZN(n9879) );
  NAND4_X1 U10889 ( .A1(n9882), .A2(n9881), .A3(n9880), .A4(n9879), .ZN(n9884)
         );
  XNOR2_X1 U10890 ( .A(P1_D_REG_3__SCAN_IN), .B(keyinput_125), .ZN(n9883) );
  OAI21_X1 U10891 ( .B1(n9885), .B2(n9884), .A(n9883), .ZN(n9888) );
  XOR2_X1 U10892 ( .A(keyinput_127), .B(P1_D_REG_5__SCAN_IN), .Z(n9887) );
  XOR2_X1 U10893 ( .A(keyinput_126), .B(P1_D_REG_4__SCAN_IN), .Z(n9886) );
  NAND3_X1 U10894 ( .A1(n9888), .A2(n9887), .A3(n9886), .ZN(n10108) );
  XOR2_X1 U10895 ( .A(P1_D_REG_4__SCAN_IN), .B(keyinput_254), .Z(n10107) );
  XOR2_X1 U10896 ( .A(P1_D_REG_5__SCAN_IN), .B(keyinput_255), .Z(n10106) );
  XNOR2_X1 U10897 ( .A(P2_WR_REG_SCAN_IN), .B(keyinput_128), .ZN(n9892) );
  XNOR2_X1 U10898 ( .A(SI_31_), .B(keyinput_129), .ZN(n9891) );
  XNOR2_X1 U10899 ( .A(n9889), .B(keyinput_130), .ZN(n9890) );
  OAI21_X1 U10900 ( .B1(n9892), .B2(n9891), .A(n9890), .ZN(n9903) );
  XNOR2_X1 U10901 ( .A(SI_29_), .B(keyinput_131), .ZN(n9902) );
  XNOR2_X1 U10902 ( .A(n9893), .B(keyinput_133), .ZN(n9895) );
  XNOR2_X1 U10903 ( .A(SI_26_), .B(keyinput_134), .ZN(n9894) );
  NOR2_X1 U10904 ( .A1(n9895), .A2(n9894), .ZN(n9900) );
  XNOR2_X1 U10905 ( .A(n9896), .B(keyinput_135), .ZN(n9899) );
  XNOR2_X1 U10906 ( .A(SI_28_), .B(keyinput_132), .ZN(n9898) );
  XNOR2_X1 U10907 ( .A(SI_24_), .B(keyinput_136), .ZN(n9897) );
  NAND4_X1 U10908 ( .A1(n9900), .A2(n9899), .A3(n9898), .A4(n9897), .ZN(n9901)
         );
  AOI21_X1 U10909 ( .B1(n9903), .B2(n9902), .A(n9901), .ZN(n9906) );
  XNOR2_X1 U10910 ( .A(SI_23_), .B(keyinput_137), .ZN(n9905) );
  XNOR2_X1 U10911 ( .A(SI_22_), .B(keyinput_138), .ZN(n9904) );
  OAI21_X1 U10912 ( .B1(n9906), .B2(n9905), .A(n9904), .ZN(n9911) );
  XNOR2_X1 U10913 ( .A(n9907), .B(keyinput_141), .ZN(n9910) );
  XNOR2_X1 U10914 ( .A(SI_21_), .B(keyinput_139), .ZN(n9909) );
  XNOR2_X1 U10915 ( .A(SI_20_), .B(keyinput_140), .ZN(n9908) );
  NAND4_X1 U10916 ( .A1(n9911), .A2(n9910), .A3(n9909), .A4(n9908), .ZN(n9916)
         );
  XNOR2_X1 U10917 ( .A(n9912), .B(keyinput_142), .ZN(n9915) );
  XNOR2_X1 U10918 ( .A(n9913), .B(keyinput_143), .ZN(n9914) );
  NAND3_X1 U10919 ( .A1(n9916), .A2(n9915), .A3(n9914), .ZN(n9922) );
  XNOR2_X1 U10920 ( .A(SI_16_), .B(keyinput_144), .ZN(n9921) );
  XNOR2_X1 U10921 ( .A(SI_13_), .B(keyinput_147), .ZN(n9919) );
  XNOR2_X1 U10922 ( .A(SI_14_), .B(keyinput_146), .ZN(n9918) );
  XNOR2_X1 U10923 ( .A(SI_15_), .B(keyinput_145), .ZN(n9917) );
  NAND3_X1 U10924 ( .A1(n9919), .A2(n9918), .A3(n9917), .ZN(n9920) );
  AOI21_X1 U10925 ( .B1(n9922), .B2(n9921), .A(n9920), .ZN(n9927) );
  XOR2_X1 U10926 ( .A(SI_12_), .B(keyinput_148), .Z(n9926) );
  XNOR2_X1 U10927 ( .A(n9923), .B(keyinput_150), .ZN(n9925) );
  XNOR2_X1 U10928 ( .A(SI_11_), .B(keyinput_149), .ZN(n9924) );
  OAI211_X1 U10929 ( .C1(n9927), .C2(n9926), .A(n9925), .B(n9924), .ZN(n9931)
         );
  XNOR2_X1 U10930 ( .A(n9928), .B(keyinput_151), .ZN(n9930) );
  XNOR2_X1 U10931 ( .A(SI_8_), .B(keyinput_152), .ZN(n9929) );
  NAND3_X1 U10932 ( .A1(n9931), .A2(n9930), .A3(n9929), .ZN(n9935) );
  XNOR2_X1 U10933 ( .A(n9932), .B(keyinput_153), .ZN(n9934) );
  XNOR2_X1 U10934 ( .A(SI_6_), .B(keyinput_154), .ZN(n9933) );
  AOI21_X1 U10935 ( .B1(n9935), .B2(n9934), .A(n9933), .ZN(n9947) );
  XNOR2_X1 U10936 ( .A(SI_5_), .B(keyinput_155), .ZN(n9946) );
  XNOR2_X1 U10937 ( .A(n9936), .B(keyinput_157), .ZN(n9939) );
  XNOR2_X1 U10938 ( .A(SI_0_), .B(keyinput_160), .ZN(n9938) );
  XNOR2_X1 U10939 ( .A(SI_2_), .B(keyinput_158), .ZN(n9937) );
  NAND3_X1 U10940 ( .A1(n9939), .A2(n9938), .A3(n9937), .ZN(n9944) );
  XNOR2_X1 U10941 ( .A(n9940), .B(keyinput_159), .ZN(n9943) );
  XNOR2_X1 U10942 ( .A(n9941), .B(keyinput_156), .ZN(n9942) );
  NOR3_X1 U10943 ( .A1(n9944), .A2(n9943), .A3(n9942), .ZN(n9945) );
  OAI21_X1 U10944 ( .B1(n9947), .B2(n9946), .A(n9945), .ZN(n9950) );
  XNOR2_X1 U10945 ( .A(P2_U3151), .B(keyinput_162), .ZN(n9949) );
  XNOR2_X1 U10946 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_161), .ZN(n9948) );
  NAND3_X1 U10947 ( .A1(n9950), .A2(n9949), .A3(n9948), .ZN(n9955) );
  XNOR2_X1 U10948 ( .A(n9951), .B(keyinput_163), .ZN(n9954) );
  XNOR2_X1 U10949 ( .A(P2_REG3_REG_27__SCAN_IN), .B(keyinput_164), .ZN(n9953)
         );
  XNOR2_X1 U10950 ( .A(P2_REG3_REG_14__SCAN_IN), .B(keyinput_165), .ZN(n9952)
         );
  NAND4_X1 U10951 ( .A1(n9955), .A2(n9954), .A3(n9953), .A4(n9952), .ZN(n9958)
         );
  XOR2_X1 U10952 ( .A(P2_REG3_REG_23__SCAN_IN), .B(keyinput_166), .Z(n9957) );
  XNOR2_X1 U10953 ( .A(P2_REG3_REG_10__SCAN_IN), .B(keyinput_167), .ZN(n9956)
         );
  AOI21_X1 U10954 ( .B1(n9958), .B2(n9957), .A(n9956), .ZN(n9962) );
  XNOR2_X1 U10955 ( .A(n9959), .B(keyinput_168), .ZN(n9961) );
  XNOR2_X1 U10956 ( .A(P2_REG3_REG_19__SCAN_IN), .B(keyinput_169), .ZN(n9960)
         );
  NOR3_X1 U10957 ( .A1(n9962), .A2(n9961), .A3(n9960), .ZN(n9965) );
  XOR2_X1 U10958 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_170), .Z(n9964) );
  XNOR2_X1 U10959 ( .A(P2_REG3_REG_8__SCAN_IN), .B(keyinput_171), .ZN(n9963)
         );
  OAI21_X1 U10960 ( .B1(n9965), .B2(n9964), .A(n9963), .ZN(n9974) );
  XNOR2_X1 U10961 ( .A(P2_REG3_REG_1__SCAN_IN), .B(keyinput_172), .ZN(n9973)
         );
  XOR2_X1 U10962 ( .A(P2_REG3_REG_16__SCAN_IN), .B(keyinput_176), .Z(n9971) );
  XNOR2_X1 U10963 ( .A(n9966), .B(keyinput_173), .ZN(n9970) );
  XNOR2_X1 U10964 ( .A(n9967), .B(keyinput_174), .ZN(n9969) );
  XNOR2_X1 U10965 ( .A(P2_REG3_REG_25__SCAN_IN), .B(keyinput_175), .ZN(n9968)
         );
  NAND4_X1 U10966 ( .A1(n9971), .A2(n9970), .A3(n9969), .A4(n9968), .ZN(n9972)
         );
  AOI21_X1 U10967 ( .B1(n9974), .B2(n9973), .A(n9972), .ZN(n9978) );
  XNOR2_X1 U10968 ( .A(n9975), .B(keyinput_177), .ZN(n9977) );
  XNOR2_X1 U10969 ( .A(P2_REG3_REG_17__SCAN_IN), .B(keyinput_178), .ZN(n9976)
         );
  OAI21_X1 U10970 ( .B1(n9978), .B2(n9977), .A(n9976), .ZN(n9982) );
  XNOR2_X1 U10971 ( .A(n9979), .B(keyinput_179), .ZN(n9981) );
  XNOR2_X1 U10972 ( .A(P2_REG3_REG_4__SCAN_IN), .B(keyinput_180), .ZN(n9980)
         );
  AOI21_X1 U10973 ( .B1(n9982), .B2(n9981), .A(n9980), .ZN(n9993) );
  XNOR2_X1 U10974 ( .A(P2_REG3_REG_9__SCAN_IN), .B(keyinput_181), .ZN(n9992)
         );
  AOI22_X1 U10975 ( .A1(n5738), .A2(keyinput_184), .B1(keyinput_186), .B2(
        n9984), .ZN(n9983) );
  OAI221_X1 U10976 ( .B1(n5738), .B2(keyinput_184), .C1(n9984), .C2(
        keyinput_186), .A(n9983), .ZN(n9990) );
  AOI22_X1 U10977 ( .A1(n9987), .A2(keyinput_183), .B1(n9986), .B2(
        keyinput_185), .ZN(n9985) );
  OAI221_X1 U10978 ( .B1(n9987), .B2(keyinput_183), .C1(n9986), .C2(
        keyinput_185), .A(n9985), .ZN(n9989) );
  XNOR2_X1 U10979 ( .A(P2_REG3_REG_0__SCAN_IN), .B(keyinput_182), .ZN(n9988)
         );
  NOR3_X1 U10980 ( .A1(n9990), .A2(n9989), .A3(n9988), .ZN(n9991) );
  OAI21_X1 U10981 ( .B1(n9993), .B2(n9992), .A(n9991), .ZN(n9996) );
  XNOR2_X1 U10982 ( .A(P2_REG3_REG_2__SCAN_IN), .B(keyinput_187), .ZN(n9995)
         );
  XNOR2_X1 U10983 ( .A(P2_REG3_REG_18__SCAN_IN), .B(keyinput_188), .ZN(n9994)
         );
  AOI21_X1 U10984 ( .B1(n9996), .B2(n9995), .A(n9994), .ZN(n10006) );
  XNOR2_X1 U10985 ( .A(P2_REG3_REG_6__SCAN_IN), .B(keyinput_189), .ZN(n10005)
         );
  XOR2_X1 U10986 ( .A(P2_REG3_REG_26__SCAN_IN), .B(keyinput_190), .Z(n10003)
         );
  XNOR2_X1 U10987 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(keyinput_193), .ZN(n9999)
         );
  XNOR2_X1 U10988 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(keyinput_194), .ZN(n9998)
         );
  XNOR2_X1 U10989 ( .A(P2_B_REG_SCAN_IN), .B(keyinput_192), .ZN(n9997) );
  NAND3_X1 U10990 ( .A1(n9999), .A2(n9998), .A3(n9997), .ZN(n10002) );
  XNOR2_X1 U10991 ( .A(n10000), .B(keyinput_191), .ZN(n10001) );
  NOR3_X1 U10992 ( .A1(n10003), .A2(n10002), .A3(n10001), .ZN(n10004) );
  OAI21_X1 U10993 ( .B1(n10006), .B2(n10005), .A(n10004), .ZN(n10009) );
  XNOR2_X1 U10994 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(keyinput_195), .ZN(n10008) );
  XNOR2_X1 U10995 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(keyinput_196), .ZN(n10007) );
  AOI21_X1 U10996 ( .B1(n10009), .B2(n10008), .A(n10007), .ZN(n10012) );
  XNOR2_X1 U10997 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(keyinput_197), .ZN(n10011) );
  XNOR2_X1 U10998 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(keyinput_198), .ZN(n10010) );
  OAI21_X1 U10999 ( .B1(n10012), .B2(n10011), .A(n10010), .ZN(n10016) );
  XNOR2_X1 U11000 ( .A(n10013), .B(keyinput_199), .ZN(n10015) );
  XNOR2_X1 U11001 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(keyinput_200), .ZN(n10014) );
  NAND3_X1 U11002 ( .A1(n10016), .A2(n10015), .A3(n10014), .ZN(n10020) );
  XNOR2_X1 U11003 ( .A(n10017), .B(keyinput_201), .ZN(n10019) );
  XNOR2_X1 U11004 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(keyinput_202), .ZN(n10018) );
  AOI21_X1 U11005 ( .B1(n10020), .B2(n10019), .A(n10018), .ZN(n10024) );
  XOR2_X1 U11006 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(keyinput_203), .Z(n10023)
         );
  XNOR2_X1 U11007 ( .A(n10021), .B(keyinput_204), .ZN(n10022) );
  NOR3_X1 U11008 ( .A1(n10024), .A2(n10023), .A3(n10022), .ZN(n10031) );
  XNOR2_X1 U11009 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(keyinput_205), .ZN(n10030) );
  XNOR2_X1 U11010 ( .A(n10025), .B(keyinput_208), .ZN(n10028) );
  XNOR2_X1 U11011 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(keyinput_207), .ZN(n10027) );
  XNOR2_X1 U11012 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(keyinput_206), .ZN(n10026) );
  NOR3_X1 U11013 ( .A1(n10028), .A2(n10027), .A3(n10026), .ZN(n10029) );
  OAI21_X1 U11014 ( .B1(n10031), .B2(n10030), .A(n10029), .ZN(n10040) );
  XOR2_X1 U11015 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(keyinput_209), .Z(n10036)
         );
  XOR2_X1 U11016 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(keyinput_212), .Z(n10035)
         );
  XNOR2_X1 U11017 ( .A(n10032), .B(keyinput_210), .ZN(n10034) );
  XNOR2_X1 U11018 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(keyinput_211), .ZN(n10033) );
  NOR4_X1 U11019 ( .A1(n10036), .A2(n10035), .A3(n10034), .A4(n10033), .ZN(
        n10039) );
  XNOR2_X1 U11020 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(keyinput_214), .ZN(n10038) );
  XNOR2_X1 U11021 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(keyinput_213), .ZN(n10037) );
  AOI211_X1 U11022 ( .C1(n10040), .C2(n10039), .A(n10038), .B(n10037), .ZN(
        n10043) );
  XNOR2_X1 U11023 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(keyinput_215), .ZN(n10042)
         );
  XNOR2_X1 U11024 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(keyinput_216), .ZN(n10041)
         );
  NOR3_X1 U11025 ( .A1(n10043), .A2(n10042), .A3(n10041), .ZN(n10046) );
  XNOR2_X1 U11026 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(keyinput_217), .ZN(n10045)
         );
  XNOR2_X1 U11027 ( .A(P1_IR_REG_0__SCAN_IN), .B(keyinput_218), .ZN(n10044) );
  NOR3_X1 U11028 ( .A1(n10046), .A2(n10045), .A3(n10044), .ZN(n10054) );
  XNOR2_X1 U11029 ( .A(P1_IR_REG_2__SCAN_IN), .B(keyinput_220), .ZN(n10053) );
  XNOR2_X1 U11030 ( .A(P1_IR_REG_6__SCAN_IN), .B(keyinput_224), .ZN(n10052) );
  XOR2_X1 U11031 ( .A(P1_IR_REG_1__SCAN_IN), .B(keyinput_219), .Z(n10050) );
  XOR2_X1 U11032 ( .A(P1_IR_REG_3__SCAN_IN), .B(keyinput_221), .Z(n10049) );
  XNOR2_X1 U11033 ( .A(P1_IR_REG_4__SCAN_IN), .B(keyinput_222), .ZN(n10048) );
  XNOR2_X1 U11034 ( .A(P1_IR_REG_5__SCAN_IN), .B(keyinput_223), .ZN(n10047) );
  NAND4_X1 U11035 ( .A1(n10050), .A2(n10049), .A3(n10048), .A4(n10047), .ZN(
        n10051) );
  NOR4_X1 U11036 ( .A1(n10054), .A2(n10053), .A3(n10052), .A4(n10051), .ZN(
        n10057) );
  XNOR2_X1 U11037 ( .A(P1_IR_REG_7__SCAN_IN), .B(keyinput_225), .ZN(n10056) );
  XNOR2_X1 U11038 ( .A(P1_IR_REG_8__SCAN_IN), .B(keyinput_226), .ZN(n10055) );
  NOR3_X1 U11039 ( .A1(n10057), .A2(n10056), .A3(n10055), .ZN(n10060) );
  XOR2_X1 U11040 ( .A(P1_IR_REG_10__SCAN_IN), .B(keyinput_228), .Z(n10059) );
  XNOR2_X1 U11041 ( .A(P1_IR_REG_9__SCAN_IN), .B(keyinput_227), .ZN(n10058) );
  NOR3_X1 U11042 ( .A1(n10060), .A2(n10059), .A3(n10058), .ZN(n10081) );
  XNOR2_X1 U11043 ( .A(n10061), .B(keyinput_229), .ZN(n10066) );
  XNOR2_X1 U11044 ( .A(n10062), .B(keyinput_232), .ZN(n10065) );
  XNOR2_X1 U11045 ( .A(P1_IR_REG_13__SCAN_IN), .B(keyinput_231), .ZN(n10064)
         );
  XNOR2_X1 U11046 ( .A(P1_IR_REG_12__SCAN_IN), .B(keyinput_230), .ZN(n10063)
         );
  NAND4_X1 U11047 ( .A1(n10066), .A2(n10065), .A3(n10064), .A4(n10063), .ZN(
        n10080) );
  OAI22_X1 U11048 ( .A1(n10069), .A2(keyinput_240), .B1(keyinput_241), .B2(
        P1_IR_REG_23__SCAN_IN), .ZN(n10068) );
  AND2_X1 U11049 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(keyinput_241), .ZN(n10067)
         );
  AOI211_X1 U11050 ( .C1(keyinput_240), .C2(n10069), .A(n10068), .B(n10067), 
        .ZN(n10073) );
  XNOR2_X1 U11051 ( .A(P1_IR_REG_18__SCAN_IN), .B(keyinput_236), .ZN(n10072)
         );
  XNOR2_X1 U11052 ( .A(P1_IR_REG_20__SCAN_IN), .B(keyinput_238), .ZN(n10071)
         );
  XNOR2_X1 U11053 ( .A(P1_IR_REG_15__SCAN_IN), .B(keyinput_233), .ZN(n10070)
         );
  NAND4_X1 U11054 ( .A1(n10073), .A2(n10072), .A3(n10071), .A4(n10070), .ZN(
        n10078) );
  AOI22_X1 U11055 ( .A1(n7454), .A2(keyinput_235), .B1(keyinput_239), .B2(
        n6462), .ZN(n10074) );
  OAI221_X1 U11056 ( .B1(n7454), .B2(keyinput_235), .C1(n6462), .C2(
        keyinput_239), .A(n10074), .ZN(n10077) );
  XNOR2_X1 U11057 ( .A(P1_IR_REG_16__SCAN_IN), .B(keyinput_234), .ZN(n10076)
         );
  XNOR2_X1 U11058 ( .A(P1_IR_REG_19__SCAN_IN), .B(keyinput_237), .ZN(n10075)
         );
  NOR4_X1 U11059 ( .A1(n10078), .A2(n10077), .A3(n10076), .A4(n10075), .ZN(
        n10079) );
  OAI21_X1 U11060 ( .B1(n10081), .B2(n10080), .A(n10079), .ZN(n10088) );
  XNOR2_X1 U11061 ( .A(n10082), .B(keyinput_242), .ZN(n10087) );
  XNOR2_X1 U11062 ( .A(n10083), .B(keyinput_243), .ZN(n10086) );
  XNOR2_X1 U11063 ( .A(n10084), .B(keyinput_244), .ZN(n10085) );
  AOI211_X1 U11064 ( .C1(n10088), .C2(n10087), .A(n10086), .B(n10085), .ZN(
        n10092) );
  XNOR2_X1 U11065 ( .A(n10089), .B(keyinput_246), .ZN(n10091) );
  XNOR2_X1 U11066 ( .A(P1_IR_REG_27__SCAN_IN), .B(keyinput_245), .ZN(n10090)
         );
  NOR3_X1 U11067 ( .A1(n10092), .A2(n10091), .A3(n10090), .ZN(n10096) );
  XNOR2_X1 U11068 ( .A(n10093), .B(keyinput_247), .ZN(n10095) );
  XNOR2_X1 U11069 ( .A(P1_IR_REG_30__SCAN_IN), .B(keyinput_248), .ZN(n10094)
         );
  NOR3_X1 U11070 ( .A1(n10096), .A2(n10095), .A3(n10094), .ZN(n10104) );
  INV_X1 U11071 ( .A(P1_D_REG_2__SCAN_IN), .ZN(n10527) );
  XNOR2_X1 U11072 ( .A(n10527), .B(keyinput_252), .ZN(n10101) );
  XNOR2_X1 U11073 ( .A(n10097), .B(keyinput_250), .ZN(n10100) );
  XNOR2_X1 U11074 ( .A(P1_D_REG_1__SCAN_IN), .B(keyinput_251), .ZN(n10099) );
  XNOR2_X1 U11075 ( .A(P1_IR_REG_31__SCAN_IN), .B(keyinput_249), .ZN(n10098)
         );
  NAND4_X1 U11076 ( .A1(n10101), .A2(n10100), .A3(n10099), .A4(n10098), .ZN(
        n10103) );
  INV_X1 U11077 ( .A(P1_D_REG_3__SCAN_IN), .ZN(n10528) );
  XNOR2_X1 U11078 ( .A(n10528), .B(keyinput_253), .ZN(n10102) );
  OAI21_X1 U11079 ( .B1(n10104), .B2(n10103), .A(n10102), .ZN(n10105) );
  NAND4_X1 U11080 ( .A1(n10108), .A2(n10107), .A3(n10106), .A4(n10105), .ZN(
        n10109) );
  XOR2_X1 U11081 ( .A(n10110), .B(n10109), .Z(P1_U3253) );
  MUX2_X1 U11082 ( .A(n10111), .B(P1_REG1_REG_13__SCAN_IN), .S(n10743), .Z(
        n10736) );
  OAI21_X1 U11083 ( .B1(P1_REG1_REG_12__SCAN_IN), .B2(n10122), .A(n10112), 
        .ZN(n10737) );
  NOR2_X1 U11084 ( .A1(n10736), .A2(n10737), .ZN(n10735) );
  MUX2_X1 U11085 ( .A(n10113), .B(P1_REG1_REG_14__SCAN_IN), .S(n10699), .Z(
        n10703) );
  NOR2_X1 U11086 ( .A1(n10702), .A2(n10703), .ZN(n10701) );
  NOR2_X1 U11087 ( .A1(n10114), .A2(n5387), .ZN(n10115) );
  XNOR2_X1 U11088 ( .A(n5387), .B(n10114), .ZN(n10713) );
  NOR2_X1 U11089 ( .A1(n7993), .A2(n10713), .ZN(n10712) );
  NOR2_X1 U11090 ( .A1(n10115), .A2(n10712), .ZN(n10117) );
  AOI22_X1 U11091 ( .A1(n10140), .A2(P1_REG1_REG_16__SCAN_IN), .B1(n8019), 
        .B2(n10120), .ZN(n10116) );
  OAI21_X1 U11092 ( .B1(n10117), .B2(n10116), .A(n10139), .ZN(n10132) );
  AOI21_X1 U11093 ( .B1(n10942), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10118), 
        .ZN(n10119) );
  OAI21_X1 U11094 ( .B1(n10949), .B2(n10120), .A(n10119), .ZN(n10131) );
  OAI21_X1 U11095 ( .B1(n10122), .B2(P1_REG2_REG_12__SCAN_IN), .A(n10121), 
        .ZN(n10740) );
  NAND2_X1 U11096 ( .A1(n10743), .A2(P1_REG2_REG_13__SCAN_IN), .ZN(n10123) );
  OAI21_X1 U11097 ( .B1(n10743), .B2(P1_REG2_REG_13__SCAN_IN), .A(n10123), 
        .ZN(n10739) );
  NOR2_X1 U11098 ( .A1(n10740), .A2(n10739), .ZN(n10738) );
  NAND2_X1 U11099 ( .A1(n10699), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10124) );
  OAI21_X1 U11100 ( .B1(n10699), .B2(P1_REG2_REG_14__SCAN_IN), .A(n10124), 
        .ZN(n10695) );
  NOR2_X1 U11101 ( .A1(n10125), .A2(n5387), .ZN(n10126) );
  NOR2_X1 U11102 ( .A1(n8038), .A2(n10715), .ZN(n10714) );
  NOR2_X1 U11103 ( .A1(n10126), .A2(n10714), .ZN(n10129) );
  NAND2_X1 U11104 ( .A1(n10140), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n10127) );
  OAI21_X1 U11105 ( .B1(n10140), .B2(P1_REG2_REG_16__SCAN_IN), .A(n10127), 
        .ZN(n10128) );
  NOR2_X1 U11106 ( .A1(n10129), .A2(n10128), .ZN(n10135) );
  AOI211_X1 U11107 ( .C1(n10129), .C2(n10128), .A(n10135), .B(n10958), .ZN(
        n10130) );
  AOI211_X1 U11108 ( .C1(n10954), .C2(n10132), .A(n10131), .B(n10130), .ZN(
        n10133) );
  INV_X1 U11109 ( .A(n10133), .ZN(P1_U3259) );
  NOR2_X1 U11110 ( .A1(P1_REG2_REG_17__SCAN_IN), .A2(n10154), .ZN(n10134) );
  AOI21_X1 U11111 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n10154), .A(n10134), 
        .ZN(n10137) );
  AOI21_X1 U11112 ( .B1(P1_REG2_REG_16__SCAN_IN), .B2(n10140), .A(n10135), 
        .ZN(n10136) );
  NAND2_X1 U11113 ( .A1(n10137), .A2(n10136), .ZN(n10150) );
  OAI21_X1 U11114 ( .B1(n10137), .B2(n10136), .A(n10150), .ZN(n10138) );
  INV_X1 U11115 ( .A(n10138), .ZN(n10149) );
  AOI22_X1 U11116 ( .A1(n10145), .A2(n6519), .B1(P1_REG1_REG_17__SCAN_IN), 
        .B2(n10154), .ZN(n10142) );
  NAND2_X1 U11117 ( .A1(n10142), .A2(n10141), .ZN(n10153) );
  OAI21_X1 U11118 ( .B1(n10142), .B2(n10141), .A(n10153), .ZN(n10147) );
  NAND2_X1 U11119 ( .A1(n10942), .A2(P1_ADDR_REG_17__SCAN_IN), .ZN(n10144) );
  OAI211_X1 U11120 ( .C1(n10949), .C2(n10145), .A(n10144), .B(n10143), .ZN(
        n10146) );
  AOI21_X1 U11121 ( .B1(n10147), .B2(n10954), .A(n10146), .ZN(n10148) );
  OAI21_X1 U11122 ( .B1(n10149), .B2(n10958), .A(n10148), .ZN(P1_U3260) );
  OAI21_X1 U11123 ( .B1(P1_REG2_REG_17__SCAN_IN), .B2(n10154), .A(n10150), 
        .ZN(n10727) );
  XNOR2_X1 U11124 ( .A(n10730), .B(P1_REG2_REG_18__SCAN_IN), .ZN(n10726) );
  NOR2_X1 U11125 ( .A1(n10727), .A2(n10726), .ZN(n10725) );
  AOI21_X1 U11126 ( .B1(n10730), .B2(P1_REG2_REG_18__SCAN_IN), .A(n10725), 
        .ZN(n10152) );
  MUX2_X1 U11127 ( .A(n10357), .B(P1_REG2_REG_19__SCAN_IN), .S(n10158), .Z(
        n10151) );
  XNOR2_X1 U11128 ( .A(n10152), .B(n10151), .ZN(n10167) );
  OAI21_X1 U11129 ( .B1(P1_REG1_REG_17__SCAN_IN), .B2(n10154), .A(n10153), 
        .ZN(n10723) );
  NAND2_X1 U11130 ( .A1(n10730), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n10155) );
  OAI21_X1 U11131 ( .B1(n10730), .B2(P1_REG1_REG_18__SCAN_IN), .A(n10155), 
        .ZN(n10724) );
  INV_X1 U11132 ( .A(n10155), .ZN(n10156) );
  NOR2_X1 U11133 ( .A1(n10722), .A2(n10156), .ZN(n10160) );
  XNOR2_X1 U11134 ( .A(n10158), .B(n10157), .ZN(n10159) );
  XNOR2_X1 U11135 ( .A(n10160), .B(n10159), .ZN(n10165) );
  NAND2_X1 U11136 ( .A1(n10942), .A2(P1_ADDR_REG_19__SCAN_IN), .ZN(n10161) );
  OAI211_X1 U11137 ( .C1(n10949), .C2(n10163), .A(n10162), .B(n10161), .ZN(
        n10164) );
  AOI21_X1 U11138 ( .B1(n10165), .B2(n10954), .A(n10164), .ZN(n10166) );
  OAI21_X1 U11139 ( .B1(n10167), .B2(n10958), .A(n10166), .ZN(P1_U3262) );
  NAND2_X1 U11140 ( .A1(n10448), .A2(n10309), .ZN(n10292) );
  NAND2_X1 U11141 ( .A1(n10435), .A2(n10276), .ZN(n10265) );
  NAND2_X1 U11142 ( .A1(n10206), .A2(n10396), .ZN(n10174) );
  INV_X1 U11143 ( .A(P1_B_REG_SCAN_IN), .ZN(n10168) );
  NOR2_X1 U11144 ( .A1(n10522), .A2(n10168), .ZN(n10169) );
  NOR2_X1 U11145 ( .A1(n11107), .A2(n10169), .ZN(n10207) );
  NAND2_X1 U11146 ( .A1(n10170), .A2(n10207), .ZN(n10394) );
  NOR2_X1 U11147 ( .A1(n7171), .A2(n10394), .ZN(n10175) );
  AOI21_X1 U11148 ( .B1(n7171), .B2(P1_REG2_REG_31__SCAN_IN), .A(n10175), .ZN(
        n10173) );
  NAND2_X1 U11149 ( .A1(n10171), .A2(n11124), .ZN(n10172) );
  OAI211_X1 U11150 ( .C1(n10392), .C2(n10333), .A(n10173), .B(n10172), .ZN(
        P1_U3263) );
  OAI211_X1 U11151 ( .C1(n10206), .C2(n10396), .A(n5131), .B(n10174), .ZN(
        n10395) );
  AOI21_X1 U11152 ( .B1(n7171), .B2(P1_REG2_REG_30__SCAN_IN), .A(n10175), .ZN(
        n10178) );
  NAND2_X1 U11153 ( .A1(n10176), .A2(n11124), .ZN(n10177) );
  OAI211_X1 U11154 ( .C1(n10395), .C2(n10333), .A(n10178), .B(n10177), .ZN(
        P1_U3264) );
  INV_X1 U11155 ( .A(n10179), .ZN(n10305) );
  INV_X1 U11156 ( .A(n10188), .ZN(n10189) );
  INV_X1 U11157 ( .A(n10404), .ZN(n10217) );
  NAND2_X1 U11158 ( .A1(n10478), .A2(n10375), .ZN(n10193) );
  INV_X1 U11159 ( .A(n10478), .ZN(n10355) );
  INV_X1 U11160 ( .A(n10337), .ZN(n10346) );
  INV_X1 U11161 ( .A(n10304), .ZN(n10194) );
  NOR2_X1 U11162 ( .A1(n10299), .A2(n10453), .ZN(n10195) );
  INV_X1 U11163 ( .A(n10442), .ZN(n10277) );
  NOR2_X1 U11164 ( .A1(n10271), .A2(n10424), .ZN(n10197) );
  OAI22_X1 U11165 ( .A1(n10261), .A2(n10197), .B1(n10196), .B2(n10435), .ZN(
        n10248) );
  NOR2_X1 U11166 ( .A1(n5490), .A2(n10269), .ZN(n10198) );
  INV_X1 U11167 ( .A(n10236), .ZN(n10199) );
  NAND2_X1 U11168 ( .A1(n10419), .A2(n10409), .ZN(n10200) );
  NAND2_X1 U11169 ( .A1(n10412), .A2(n10416), .ZN(n10202) );
  INV_X1 U11170 ( .A(n10203), .ZN(n10204) );
  XNOR2_X1 U11171 ( .A(n10205), .B(n10204), .ZN(n10397) );
  NAND2_X1 U11172 ( .A1(n10397), .A2(n11129), .ZN(n10216) );
  AOI211_X1 U11173 ( .C1(n10398), .C2(n10224), .A(n11212), .B(n10206), .ZN(
        n10403) );
  NAND2_X1 U11174 ( .A1(n10398), .A2(n11124), .ZN(n10212) );
  NAND2_X1 U11175 ( .A1(n10208), .A2(n10207), .ZN(n10399) );
  OAI22_X1 U11176 ( .A1(n7171), .A2(n10399), .B1(n10209), .B2(n10968), .ZN(
        n10210) );
  AOI21_X1 U11177 ( .B1(P1_REG2_REG_29__SCAN_IN), .B2(n7171), .A(n10210), .ZN(
        n10211) );
  OAI211_X1 U11178 ( .C1(n10401), .C2(n10213), .A(n10212), .B(n10211), .ZN(
        n10214) );
  AOI21_X1 U11179 ( .B1(n10403), .B2(n11128), .A(n10214), .ZN(n10215) );
  OAI211_X1 U11180 ( .C1(n10233), .C2(n10217), .A(n10216), .B(n10215), .ZN(
        P1_U3356) );
  NAND2_X1 U11181 ( .A1(n10219), .A2(n10220), .ZN(n10221) );
  NAND2_X1 U11182 ( .A1(n10407), .A2(n11129), .ZN(n10232) );
  AOI21_X1 U11183 ( .B1(n10412), .B2(n10238), .A(n11212), .ZN(n10223) );
  NAND2_X1 U11184 ( .A1(n10412), .A2(n11124), .ZN(n10229) );
  OAI22_X1 U11185 ( .A1(n10367), .A2(n10226), .B1(n10225), .B2(n10968), .ZN(
        n10227) );
  AOI21_X1 U11186 ( .B1(n10326), .B2(n10425), .A(n10227), .ZN(n10228) );
  OAI211_X1 U11187 ( .C1(n10408), .C2(n10328), .A(n10229), .B(n10228), .ZN(
        n10230) );
  AOI21_X1 U11188 ( .B1(n10410), .B2(n11128), .A(n10230), .ZN(n10231) );
  OAI211_X1 U11189 ( .C1(n10414), .C2(n10233), .A(n10232), .B(n10231), .ZN(
        P1_U3265) );
  XNOR2_X1 U11190 ( .A(n10234), .B(n10236), .ZN(n10423) );
  OAI21_X1 U11191 ( .B1(n10237), .B2(n10236), .A(n10235), .ZN(n10421) );
  AOI21_X1 U11192 ( .B1(n10244), .B2(n5167), .A(n11212), .ZN(n10239) );
  NAND2_X1 U11193 ( .A1(n10239), .A2(n10238), .ZN(n10418) );
  AOI22_X1 U11194 ( .A1(n7171), .A2(P1_REG2_REG_27__SCAN_IN), .B1(n10240), 
        .B2(n11123), .ZN(n10242) );
  NAND2_X1 U11195 ( .A1(n10326), .A2(n10432), .ZN(n10241) );
  OAI211_X1 U11196 ( .C1(n10401), .C2(n10328), .A(n10242), .B(n10241), .ZN(
        n10243) );
  AOI21_X1 U11197 ( .B1(n10244), .B2(n11124), .A(n10243), .ZN(n10245) );
  OAI21_X1 U11198 ( .B1(n10418), .B2(n10333), .A(n10245), .ZN(n10246) );
  AOI21_X1 U11199 ( .B1(n10421), .B2(n10335), .A(n10246), .ZN(n10247) );
  OAI21_X1 U11200 ( .B1(n10423), .B2(n10391), .A(n10247), .ZN(P1_U3266) );
  XNOR2_X1 U11201 ( .A(n10248), .B(n10249), .ZN(n10431) );
  XNOR2_X1 U11202 ( .A(n10250), .B(n10249), .ZN(n10429) );
  AOI21_X1 U11203 ( .B1(n10265), .B2(n10257), .A(n11212), .ZN(n10251) );
  NAND2_X1 U11204 ( .A1(n10251), .A2(n5167), .ZN(n10427) );
  OAI22_X1 U11205 ( .A1(n10367), .A2(n10253), .B1(n10252), .B2(n10968), .ZN(
        n10254) );
  AOI21_X1 U11206 ( .B1(n10326), .B2(n10424), .A(n10254), .ZN(n10255) );
  OAI21_X1 U11207 ( .B1(n10409), .B2(n10328), .A(n10255), .ZN(n10256) );
  AOI21_X1 U11208 ( .B1(n10257), .B2(n11124), .A(n10256), .ZN(n10258) );
  OAI21_X1 U11209 ( .B1(n10427), .B2(n10333), .A(n10258), .ZN(n10259) );
  AOI21_X1 U11210 ( .B1(n10429), .B2(n10335), .A(n10259), .ZN(n10260) );
  OAI21_X1 U11211 ( .B1(n10431), .B2(n10391), .A(n10260), .ZN(P1_U3267) );
  XOR2_X1 U11212 ( .A(n10261), .B(n10262), .Z(n10439) );
  AOI21_X1 U11213 ( .B1(n10263), .B2(n10262), .A(n5197), .ZN(n10264) );
  INV_X1 U11214 ( .A(n10264), .ZN(n10437) );
  OAI211_X1 U11215 ( .C1(n10435), .C2(n10276), .A(n5131), .B(n10265), .ZN(
        n10434) );
  AOI22_X1 U11216 ( .A1(n7171), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n10266), 
        .B2(n11123), .ZN(n10268) );
  NAND2_X1 U11217 ( .A1(n10326), .A2(n10445), .ZN(n10267) );
  OAI211_X1 U11218 ( .C1(n10269), .C2(n10328), .A(n10268), .B(n10267), .ZN(
        n10270) );
  AOI21_X1 U11219 ( .B1(n10271), .B2(n11124), .A(n10270), .ZN(n10272) );
  OAI21_X1 U11220 ( .B1(n10434), .B2(n10333), .A(n10272), .ZN(n10273) );
  AOI21_X1 U11221 ( .B1(n10437), .B2(n10335), .A(n10273), .ZN(n10274) );
  OAI21_X1 U11222 ( .B1(n10439), .B2(n10391), .A(n10274), .ZN(P1_U3268) );
  XOR2_X1 U11223 ( .A(n10275), .B(n10283), .Z(n10444) );
  AOI211_X1 U11224 ( .C1(n10442), .C2(n10292), .A(n11212), .B(n10276), .ZN(
        n10441) );
  NOR2_X1 U11225 ( .A1(n10277), .A2(n10387), .ZN(n10281) );
  OAI22_X1 U11226 ( .A1(n10367), .A2(n10279), .B1(n10278), .B2(n10968), .ZN(
        n10280) );
  AOI211_X1 U11227 ( .C1(n10441), .C2(n11128), .A(n10281), .B(n10280), .ZN(
        n10288) );
  OAI211_X1 U11228 ( .C1(n10284), .C2(n10283), .A(n10282), .B(n11181), .ZN(
        n10286) );
  AOI22_X1 U11229 ( .A1(n11172), .A2(n10453), .B1(n10424), .B2(n11169), .ZN(
        n10285) );
  NAND2_X1 U11230 ( .A1(n10286), .A2(n10285), .ZN(n10440) );
  NAND2_X1 U11231 ( .A1(n10440), .A2(n10367), .ZN(n10287) );
  OAI211_X1 U11232 ( .C1(n10444), .C2(n10391), .A(n10288), .B(n10287), .ZN(
        P1_U3269) );
  XNOR2_X1 U11233 ( .A(n10289), .B(n10290), .ZN(n10452) );
  XNOR2_X1 U11234 ( .A(n10291), .B(n10290), .ZN(n10450) );
  OAI211_X1 U11235 ( .C1(n10448), .C2(n10309), .A(n5131), .B(n10292), .ZN(
        n10447) );
  OAI22_X1 U11236 ( .A1(n10358), .A2(n10294), .B1(n10293), .B2(n10968), .ZN(
        n10295) );
  AOI21_X1 U11237 ( .B1(n10326), .B2(n10463), .A(n10295), .ZN(n10296) );
  OAI21_X1 U11238 ( .B1(n10297), .B2(n10328), .A(n10296), .ZN(n10298) );
  AOI21_X1 U11239 ( .B1(n10299), .B2(n11124), .A(n10298), .ZN(n10300) );
  OAI21_X1 U11240 ( .B1(n10447), .B2(n10333), .A(n10300), .ZN(n10301) );
  AOI21_X1 U11241 ( .B1(n10450), .B2(n10335), .A(n10301), .ZN(n10302) );
  OAI21_X1 U11242 ( .B1(n10452), .B2(n10391), .A(n10302), .ZN(P1_U3270) );
  XNOR2_X1 U11243 ( .A(n10303), .B(n10304), .ZN(n10461) );
  XNOR2_X1 U11244 ( .A(n10305), .B(n10304), .ZN(n10459) );
  NAND2_X1 U11245 ( .A1(n10306), .A2(n5229), .ZN(n10307) );
  NAND2_X1 U11246 ( .A1(n10307), .A2(n5131), .ZN(n10308) );
  NOR2_X1 U11247 ( .A1(n10309), .A2(n10308), .ZN(n10458) );
  NAND2_X1 U11248 ( .A1(n10458), .A2(n11128), .ZN(n10316) );
  OAI22_X1 U11249 ( .A1(n10367), .A2(n10311), .B1(n10310), .B2(n10968), .ZN(
        n10314) );
  NOR2_X1 U11250 ( .A1(n10328), .A2(n10312), .ZN(n10313) );
  AOI211_X1 U11251 ( .C1(n10326), .C2(n10454), .A(n10314), .B(n10313), .ZN(
        n10315) );
  OAI211_X1 U11252 ( .C1(n10456), .C2(n10387), .A(n10316), .B(n10315), .ZN(
        n10317) );
  AOI21_X1 U11253 ( .B1(n10459), .B2(n10335), .A(n10317), .ZN(n10318) );
  OAI21_X1 U11254 ( .B1(n10461), .B2(n10391), .A(n10318), .ZN(P1_U3271) );
  XNOR2_X1 U11255 ( .A(n10320), .B(n10319), .ZN(n10470) );
  XNOR2_X1 U11256 ( .A(n10322), .B(n10321), .ZN(n10468) );
  OAI211_X1 U11257 ( .C1(n10466), .C2(n10339), .A(n5131), .B(n5229), .ZN(
        n10465) );
  OAI22_X1 U11258 ( .A1(n10358), .A2(n10324), .B1(n10323), .B2(n10968), .ZN(
        n10325) );
  AOI21_X1 U11259 ( .B1(n10326), .B2(n10462), .A(n10325), .ZN(n10327) );
  OAI21_X1 U11260 ( .B1(n10329), .B2(n10328), .A(n10327), .ZN(n10330) );
  AOI21_X1 U11261 ( .B1(n10331), .B2(n11124), .A(n10330), .ZN(n10332) );
  OAI21_X1 U11262 ( .B1(n10465), .B2(n10333), .A(n10332), .ZN(n10334) );
  AOI21_X1 U11263 ( .B1(n10468), .B2(n10335), .A(n10334), .ZN(n10336) );
  OAI21_X1 U11264 ( .B1(n10470), .B2(n10391), .A(n10336), .ZN(P1_U3272) );
  XNOR2_X1 U11265 ( .A(n10338), .B(n10337), .ZN(n10475) );
  INV_X1 U11266 ( .A(n10354), .ZN(n10340) );
  AOI211_X1 U11267 ( .C1(n10473), .C2(n10340), .A(n11212), .B(n10339), .ZN(
        n10472) );
  NOR2_X1 U11268 ( .A1(n10341), .A2(n10387), .ZN(n10345) );
  OAI22_X1 U11269 ( .A1(n10358), .A2(n10343), .B1(n10342), .B2(n10968), .ZN(
        n10344) );
  AOI211_X1 U11270 ( .C1(n10472), .C2(n11128), .A(n10345), .B(n10344), .ZN(
        n10352) );
  XNOR2_X1 U11271 ( .A(n10347), .B(n10346), .ZN(n10348) );
  OAI222_X1 U11272 ( .A1(n11107), .A2(n10350), .B1(n11109), .B2(n10349), .C1(
        n11104), .C2(n10348), .ZN(n10471) );
  NAND2_X1 U11273 ( .A1(n10471), .A2(n10367), .ZN(n10351) );
  OAI211_X1 U11274 ( .C1(n10475), .C2(n10391), .A(n10352), .B(n10351), .ZN(
        P1_U3273) );
  XNOR2_X1 U11275 ( .A(n10353), .B(n10362), .ZN(n10480) );
  AOI211_X1 U11276 ( .C1(n10478), .C2(n10379), .A(n11212), .B(n10354), .ZN(
        n10477) );
  NOR2_X1 U11277 ( .A1(n10355), .A2(n10387), .ZN(n10360) );
  OAI22_X1 U11278 ( .A1(n10358), .A2(n10357), .B1(n10356), .B2(n10968), .ZN(
        n10359) );
  AOI211_X1 U11279 ( .C1(n10477), .C2(n11128), .A(n10360), .B(n10359), .ZN(
        n10369) );
  OAI211_X1 U11280 ( .C1(n10363), .C2(n10362), .A(n10361), .B(n11181), .ZN(
        n10366) );
  AOI22_X1 U11281 ( .A1(n10364), .A2(n11172), .B1(n11169), .B2(n10462), .ZN(
        n10365) );
  NAND2_X1 U11282 ( .A1(n10366), .A2(n10365), .ZN(n10476) );
  NAND2_X1 U11283 ( .A1(n10476), .A2(n10367), .ZN(n10368) );
  OAI211_X1 U11284 ( .C1(n10480), .C2(n10391), .A(n10369), .B(n10368), .ZN(
        P1_U3274) );
  XNOR2_X1 U11285 ( .A(n10371), .B(n10370), .ZN(n10485) );
  OAI211_X1 U11286 ( .C1(n10374), .C2(n10373), .A(n10372), .B(n11181), .ZN(
        n10377) );
  NAND2_X1 U11287 ( .A1(n10375), .A2(n11169), .ZN(n10376) );
  OAI211_X1 U11288 ( .C1(n10378), .C2(n11109), .A(n10377), .B(n10376), .ZN(
        n10481) );
  INV_X1 U11289 ( .A(n10483), .ZN(n10388) );
  INV_X1 U11290 ( .A(n10379), .ZN(n10380) );
  AOI211_X1 U11291 ( .C1(n10483), .C2(n10382), .A(n11212), .B(n10380), .ZN(
        n10482) );
  NAND2_X1 U11292 ( .A1(n10482), .A2(n11128), .ZN(n10386) );
  INV_X1 U11293 ( .A(n10383), .ZN(n10384) );
  AOI22_X1 U11294 ( .A1(n7171), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n10384), 
        .B2(n11123), .ZN(n10385) );
  OAI211_X1 U11295 ( .C1(n10388), .C2(n10387), .A(n10386), .B(n10385), .ZN(
        n10389) );
  AOI21_X1 U11296 ( .B1(n10358), .B2(n10481), .A(n10389), .ZN(n10390) );
  OAI21_X1 U11297 ( .B1(n10485), .B2(n10391), .A(n10390), .ZN(P1_U3275) );
  MUX2_X1 U11298 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10491), .S(n11202), .Z(
        P1_U3553) );
  OAI211_X1 U11299 ( .C1(n10396), .C2(n11195), .A(n10395), .B(n10394), .ZN(
        n10492) );
  MUX2_X1 U11300 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10492), .S(n11202), .Z(
        P1_U3552) );
  NAND2_X1 U11301 ( .A1(n10397), .A2(n11199), .ZN(n10406) );
  NAND2_X1 U11302 ( .A1(n10398), .A2(n11147), .ZN(n10400) );
  OAI211_X1 U11303 ( .C1(n10401), .C2(n11109), .A(n10400), .B(n10399), .ZN(
        n10402) );
  NAND2_X1 U11304 ( .A1(n10406), .A2(n10405), .ZN(n10493) );
  MUX2_X1 U11305 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n10493), .S(n11202), .Z(
        P1_U3551) );
  OAI22_X1 U11306 ( .A1(n10409), .A2(n11109), .B1(n10408), .B2(n11107), .ZN(
        n10411) );
  AOI211_X1 U11307 ( .C1(n11147), .C2(n10412), .A(n10411), .B(n10410), .ZN(
        n10413) );
  MUX2_X1 U11308 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10494), .S(n11202), .Z(
        P1_U3550) );
  AOI22_X1 U11309 ( .A1(n11172), .A2(n10432), .B1(n10416), .B2(n11169), .ZN(
        n10417) );
  OAI211_X1 U11310 ( .C1(n10419), .C2(n11195), .A(n10418), .B(n10417), .ZN(
        n10420) );
  AOI21_X1 U11311 ( .B1(n10421), .B2(n11181), .A(n10420), .ZN(n10422) );
  OAI21_X1 U11312 ( .B1(n10423), .B2(n11176), .A(n10422), .ZN(n10495) );
  MUX2_X1 U11313 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10495), .S(n11202), .Z(
        P1_U3549) );
  AOI22_X1 U11314 ( .A1(n10425), .A2(n11169), .B1(n11172), .B2(n10424), .ZN(
        n10426) );
  OAI211_X1 U11315 ( .C1(n5490), .C2(n11195), .A(n10427), .B(n10426), .ZN(
        n10428) );
  AOI21_X1 U11316 ( .B1(n10429), .B2(n11181), .A(n10428), .ZN(n10430) );
  OAI21_X1 U11317 ( .B1(n10431), .B2(n11176), .A(n10430), .ZN(n10496) );
  MUX2_X1 U11318 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10496), .S(n11202), .Z(
        P1_U3548) );
  AOI22_X1 U11319 ( .A1(n11172), .A2(n10445), .B1(n10432), .B2(n11169), .ZN(
        n10433) );
  OAI211_X1 U11320 ( .C1(n10435), .C2(n11195), .A(n10434), .B(n10433), .ZN(
        n10436) );
  AOI21_X1 U11321 ( .B1(n10437), .B2(n11181), .A(n10436), .ZN(n10438) );
  OAI21_X1 U11322 ( .B1(n10439), .B2(n11176), .A(n10438), .ZN(n10497) );
  MUX2_X1 U11323 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10497), .S(n11202), .Z(
        P1_U3547) );
  AOI211_X1 U11324 ( .C1(n11147), .C2(n10442), .A(n10441), .B(n10440), .ZN(
        n10443) );
  OAI21_X1 U11325 ( .B1(n10444), .B2(n11176), .A(n10443), .ZN(n10498) );
  MUX2_X1 U11326 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10498), .S(n11202), .Z(
        P1_U3546) );
  AOI22_X1 U11327 ( .A1(n11172), .A2(n10463), .B1(n10445), .B2(n11169), .ZN(
        n10446) );
  OAI211_X1 U11328 ( .C1(n10448), .C2(n11195), .A(n10447), .B(n10446), .ZN(
        n10449) );
  AOI21_X1 U11329 ( .B1(n10450), .B2(n11181), .A(n10449), .ZN(n10451) );
  OAI21_X1 U11330 ( .B1(n10452), .B2(n11176), .A(n10451), .ZN(n10499) );
  MUX2_X1 U11331 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10499), .S(n11202), .Z(
        P1_U3545) );
  AOI22_X1 U11332 ( .A1(n11172), .A2(n10454), .B1(n10453), .B2(n11169), .ZN(
        n10455) );
  OAI21_X1 U11333 ( .B1(n10456), .B2(n11195), .A(n10455), .ZN(n10457) );
  AOI211_X1 U11334 ( .C1(n10459), .C2(n11181), .A(n10458), .B(n10457), .ZN(
        n10460) );
  OAI21_X1 U11335 ( .B1(n10461), .B2(n11176), .A(n10460), .ZN(n10500) );
  MUX2_X1 U11336 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10500), .S(n11202), .Z(
        P1_U3544) );
  AOI22_X1 U11337 ( .A1(n10463), .A2(n11169), .B1(n11172), .B2(n10462), .ZN(
        n10464) );
  OAI211_X1 U11338 ( .C1(n10466), .C2(n11195), .A(n10465), .B(n10464), .ZN(
        n10467) );
  AOI21_X1 U11339 ( .B1(n10468), .B2(n11181), .A(n10467), .ZN(n10469) );
  OAI21_X1 U11340 ( .B1(n10470), .B2(n11176), .A(n10469), .ZN(n10501) );
  MUX2_X1 U11341 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10501), .S(n11202), .Z(
        P1_U3543) );
  AOI211_X1 U11342 ( .C1(n11147), .C2(n10473), .A(n10472), .B(n10471), .ZN(
        n10474) );
  OAI21_X1 U11343 ( .B1(n10475), .B2(n11176), .A(n10474), .ZN(n10502) );
  MUX2_X1 U11344 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10502), .S(n11202), .Z(
        P1_U3542) );
  AOI211_X1 U11345 ( .C1(n11147), .C2(n10478), .A(n10477), .B(n10476), .ZN(
        n10479) );
  OAI21_X1 U11346 ( .B1(n10480), .B2(n11176), .A(n10479), .ZN(n10503) );
  MUX2_X1 U11347 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10503), .S(n11202), .Z(
        P1_U3541) );
  AOI211_X1 U11348 ( .C1(n11147), .C2(n10483), .A(n10482), .B(n10481), .ZN(
        n10484) );
  OAI21_X1 U11349 ( .B1(n10485), .B2(n11176), .A(n10484), .ZN(n10504) );
  MUX2_X1 U11350 ( .A(P1_REG1_REG_18__SCAN_IN), .B(n10504), .S(n11202), .Z(
        P1_U3540) );
  AOI211_X1 U11351 ( .C1(n11147), .C2(n10488), .A(n10487), .B(n10486), .ZN(
        n10489) );
  OAI21_X1 U11352 ( .B1(n10490), .B2(n11176), .A(n10489), .ZN(n10505) );
  MUX2_X1 U11353 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10505), .S(n11202), .Z(
        P1_U3539) );
  MUX2_X1 U11354 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10492), .S(n11206), .Z(
        P1_U3520) );
  MUX2_X1 U11355 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n10493), .S(n11206), .Z(
        P1_U3519) );
  MUX2_X1 U11356 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n10494), .S(n11206), .Z(
        P1_U3518) );
  MUX2_X1 U11357 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10495), .S(n11206), .Z(
        P1_U3517) );
  MUX2_X1 U11358 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10496), .S(n11206), .Z(
        P1_U3516) );
  MUX2_X1 U11359 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10497), .S(n11206), .Z(
        P1_U3515) );
  MUX2_X1 U11360 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10498), .S(n11206), .Z(
        P1_U3514) );
  MUX2_X1 U11361 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10499), .S(n11206), .Z(
        P1_U3513) );
  MUX2_X1 U11362 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10500), .S(n11206), .Z(
        P1_U3512) );
  MUX2_X1 U11363 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10501), .S(n11206), .Z(
        P1_U3511) );
  MUX2_X1 U11364 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10502), .S(n11206), .Z(
        P1_U3510) );
  MUX2_X1 U11365 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10503), .S(n11206), .Z(
        P1_U3509) );
  MUX2_X1 U11366 ( .A(P1_REG0_REG_18__SCAN_IN), .B(n10504), .S(n11206), .Z(
        P1_U3507) );
  MUX2_X1 U11367 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10505), .S(n11206), .Z(
        P1_U3504) );
  MUX2_X1 U11368 ( .A(n10507), .B(P1_D_REG_1__SCAN_IN), .S(n10506), .Z(
        P1_U3440) );
  NAND3_X1 U11369 ( .A1(n10509), .A2(P1_IR_REG_31__SCAN_IN), .A3(
        P1_STATE_REG_SCAN_IN), .ZN(n10511) );
  OAI22_X1 U11370 ( .A1(n10508), .A2(n10511), .B1(n10510), .B2(n5141), .ZN(
        n10512) );
  AOI21_X1 U11371 ( .B1(n9452), .B2(n10513), .A(n10512), .ZN(n10514) );
  INV_X1 U11372 ( .A(n10514), .ZN(P1_U3324) );
  OAI222_X1 U11373 ( .A1(P1_U3086), .A2(n10518), .B1(n10517), .B2(n10516), 
        .C1(n10515), .C2(n5141), .ZN(P1_U3325) );
  INV_X1 U11374 ( .A(n10519), .ZN(n10520) );
  OAI222_X1 U11375 ( .A1(n5141), .A2(n10521), .B1(n10517), .B2(n10520), .C1(
        n5145), .C2(P1_U3086), .ZN(P1_U3327) );
  OAI222_X1 U11376 ( .A1(n5141), .A2(n10524), .B1(n10517), .B2(n10523), .C1(
        P1_U3086), .C2(n10522), .ZN(P1_U3328) );
  INV_X1 U11377 ( .A(n10525), .ZN(n10526) );
  MUX2_X1 U11378 ( .A(n10526), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  NOR2_X1 U11379 ( .A1(n10529), .A2(n10527), .ZN(P1_U3323) );
  NOR2_X1 U11380 ( .A1(n10529), .A2(n10528), .ZN(P1_U3322) );
  AND2_X1 U11381 ( .A1(n10530), .A2(P1_D_REG_4__SCAN_IN), .ZN(P1_U3321) );
  AND2_X1 U11382 ( .A1(n10530), .A2(P1_D_REG_5__SCAN_IN), .ZN(P1_U3320) );
  AND2_X1 U11383 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10530), .ZN(P1_U3319) );
  AND2_X1 U11384 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10530), .ZN(P1_U3318) );
  AND2_X1 U11385 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10530), .ZN(P1_U3317) );
  AND2_X1 U11386 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10530), .ZN(P1_U3316) );
  AND2_X1 U11387 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10530), .ZN(P1_U3315) );
  AND2_X1 U11388 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10530), .ZN(P1_U3314) );
  AND2_X1 U11389 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10530), .ZN(P1_U3313) );
  AND2_X1 U11390 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10530), .ZN(P1_U3312) );
  AND2_X1 U11391 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10530), .ZN(P1_U3311) );
  AND2_X1 U11392 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10530), .ZN(P1_U3310) );
  AND2_X1 U11393 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10530), .ZN(P1_U3309) );
  AND2_X1 U11394 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10530), .ZN(P1_U3308) );
  AND2_X1 U11395 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10530), .ZN(P1_U3307) );
  AND2_X1 U11396 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10530), .ZN(P1_U3306) );
  AND2_X1 U11397 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10530), .ZN(P1_U3305) );
  AND2_X1 U11398 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10530), .ZN(P1_U3304) );
  AND2_X1 U11399 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10530), .ZN(P1_U3303) );
  AND2_X1 U11400 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10530), .ZN(P1_U3302) );
  AND2_X1 U11401 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10530), .ZN(P1_U3301) );
  AND2_X1 U11402 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10530), .ZN(P1_U3300) );
  AND2_X1 U11403 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10530), .ZN(P1_U3299) );
  AND2_X1 U11404 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10530), .ZN(P1_U3298) );
  AND2_X1 U11405 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10530), .ZN(P1_U3297) );
  AND2_X1 U11406 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10530), .ZN(P1_U3296) );
  AND2_X1 U11407 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10530), .ZN(P1_U3295) );
  AND2_X1 U11408 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10530), .ZN(P1_U3294) );
  XOR2_X1 U11409 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1068_U46) );
  OAI222_X1 U11410 ( .A1(n10535), .A2(n10534), .B1(n10535), .B2(n10533), .C1(
        n10532), .C2(n10531), .ZN(ADD_1068_U5) );
  AOI21_X1 U11411 ( .B1(n10538), .B2(n10537), .A(n10536), .ZN(ADD_1068_U54) );
  AOI21_X1 U11412 ( .B1(n10541), .B2(n10540), .A(n10539), .ZN(ADD_1068_U53) );
  OAI21_X1 U11413 ( .B1(n10544), .B2(n10543), .A(n10542), .ZN(ADD_1068_U52) );
  OAI21_X1 U11414 ( .B1(n10547), .B2(n10546), .A(n10545), .ZN(ADD_1068_U51) );
  OAI21_X1 U11415 ( .B1(n10550), .B2(n10549), .A(n10548), .ZN(ADD_1068_U50) );
  OAI21_X1 U11416 ( .B1(n10553), .B2(n10552), .A(n10551), .ZN(ADD_1068_U49) );
  OAI21_X1 U11417 ( .B1(n10556), .B2(n10555), .A(n10554), .ZN(ADD_1068_U48) );
  OAI21_X1 U11418 ( .B1(n10559), .B2(n10558), .A(n10557), .ZN(ADD_1068_U47) );
  OAI21_X1 U11419 ( .B1(n10562), .B2(n10561), .A(n10560), .ZN(ADD_1068_U63) );
  OAI21_X1 U11420 ( .B1(n10565), .B2(n10564), .A(n10563), .ZN(ADD_1068_U62) );
  OAI21_X1 U11421 ( .B1(n10568), .B2(n10567), .A(n10566), .ZN(ADD_1068_U61) );
  OAI21_X1 U11422 ( .B1(n10571), .B2(n10570), .A(n10569), .ZN(ADD_1068_U60) );
  OAI21_X1 U11423 ( .B1(n10574), .B2(n10573), .A(n10572), .ZN(ADD_1068_U59) );
  OAI21_X1 U11424 ( .B1(n10577), .B2(n10576), .A(n10575), .ZN(ADD_1068_U58) );
  OAI21_X1 U11425 ( .B1(n10580), .B2(n10579), .A(n10578), .ZN(ADD_1068_U57) );
  OAI21_X1 U11426 ( .B1(n10583), .B2(n10582), .A(n10581), .ZN(ADD_1068_U56) );
  OAI21_X1 U11427 ( .B1(n10586), .B2(n10585), .A(n10584), .ZN(ADD_1068_U55) );
  OR2_X1 U11428 ( .A1(n5145), .A2(n10587), .ZN(n10935) );
  OR2_X1 U11429 ( .A1(n10930), .A2(n10588), .ZN(n10589) );
  OAI21_X1 U11430 ( .B1(n10935), .B2(n10590), .A(n10589), .ZN(n10591) );
  INV_X1 U11431 ( .A(n10591), .ZN(n10592) );
  XOR2_X1 U11432 ( .A(n10592), .B(P1_IR_REG_0__SCAN_IN), .Z(n10595) );
  AOI22_X1 U11433 ( .A1(P1_ADDR_REG_0__SCAN_IN), .A2(n10942), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3086), .ZN(n10593) );
  OAI21_X1 U11434 ( .B1(n10595), .B2(n10594), .A(n10593), .ZN(P1_U3243) );
  AOI22_X1 U11435 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(n10942), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n10611) );
  NAND2_X1 U11436 ( .A1(n10596), .A2(n10933), .ZN(n10599) );
  INV_X1 U11437 ( .A(n10597), .ZN(n10598) );
  NAND2_X1 U11438 ( .A1(n10599), .A2(n10598), .ZN(n10608) );
  OR2_X1 U11439 ( .A1(n10949), .A2(n10600), .ZN(n10607) );
  INV_X1 U11440 ( .A(n10601), .ZN(n10605) );
  NAND2_X1 U11441 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n10602) );
  NAND2_X1 U11442 ( .A1(n10603), .A2(n10602), .ZN(n10604) );
  NAND3_X1 U11443 ( .A1(n10954), .A2(n10605), .A3(n10604), .ZN(n10606) );
  OAI211_X1 U11444 ( .C1(n10958), .C2(n10608), .A(n10607), .B(n10606), .ZN(
        n10609) );
  INV_X1 U11445 ( .A(n10609), .ZN(n10610) );
  NAND2_X1 U11446 ( .A1(n10611), .A2(n10610), .ZN(P1_U3244) );
  AOI211_X1 U11447 ( .C1(n10614), .C2(n10613), .A(n10612), .B(n10958), .ZN(
        n10619) );
  INV_X1 U11448 ( .A(n10954), .ZN(n10734) );
  AOI211_X1 U11449 ( .C1(n10617), .C2(n10616), .A(n10615), .B(n10734), .ZN(
        n10618) );
  AOI211_X1 U11450 ( .C1(n10744), .C2(n10620), .A(n10619), .B(n10618), .ZN(
        n10621) );
  INV_X1 U11451 ( .A(n10621), .ZN(n10623) );
  AOI211_X1 U11452 ( .C1(P1_ADDR_REG_3__SCAN_IN), .C2(n10942), .A(n10623), .B(
        n10622), .ZN(n10624) );
  INV_X1 U11453 ( .A(n10624), .ZN(P1_U3246) );
  INV_X1 U11454 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n10639) );
  NAND2_X1 U11455 ( .A1(n10626), .A2(n10625), .ZN(n10627) );
  NAND2_X1 U11456 ( .A1(n10627), .A2(n5378), .ZN(n10635) );
  OR2_X1 U11457 ( .A1(n10949), .A2(n10628), .ZN(n10634) );
  AOI21_X1 U11458 ( .B1(n10631), .B2(n10630), .A(n10629), .ZN(n10632) );
  NAND2_X1 U11459 ( .A1(n10954), .A2(n10632), .ZN(n10633) );
  OAI211_X1 U11460 ( .C1(n10958), .C2(n10635), .A(n10634), .B(n10633), .ZN(
        n10636) );
  INV_X1 U11461 ( .A(n10636), .ZN(n10638) );
  OAI211_X1 U11462 ( .C1(n10733), .C2(n10639), .A(n10638), .B(n10637), .ZN(
        P1_U3248) );
  AOI211_X1 U11463 ( .C1(n10642), .C2(n10641), .A(n10640), .B(n10958), .ZN(
        n10647) );
  AOI211_X1 U11464 ( .C1(n10645), .C2(n10644), .A(n10643), .B(n10734), .ZN(
        n10646) );
  AOI211_X1 U11465 ( .C1(n10744), .C2(n10648), .A(n10647), .B(n10646), .ZN(
        n10649) );
  INV_X1 U11466 ( .A(n10649), .ZN(n10651) );
  AOI211_X1 U11467 ( .C1(n10942), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n10651), .B(
        n10650), .ZN(n10652) );
  INV_X1 U11468 ( .A(n10652), .ZN(P1_U3249) );
  INV_X1 U11469 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n10668) );
  NAND2_X1 U11470 ( .A1(n10653), .A2(n5183), .ZN(n10656) );
  INV_X1 U11471 ( .A(n10654), .ZN(n10655) );
  NAND2_X1 U11472 ( .A1(n10656), .A2(n10655), .ZN(n10664) );
  OR2_X1 U11473 ( .A1(n10949), .A2(n10657), .ZN(n10663) );
  AOI21_X1 U11474 ( .B1(n10660), .B2(n10659), .A(n10658), .ZN(n10661) );
  NAND2_X1 U11475 ( .A1(n10954), .A2(n10661), .ZN(n10662) );
  OAI211_X1 U11476 ( .C1(n10958), .C2(n10664), .A(n10663), .B(n10662), .ZN(
        n10665) );
  INV_X1 U11477 ( .A(n10665), .ZN(n10667) );
  OAI211_X1 U11478 ( .C1(n10733), .C2(n10668), .A(n10667), .B(n10666), .ZN(
        P1_U3250) );
  AOI211_X1 U11479 ( .C1(n10671), .C2(n10670), .A(n10669), .B(n10958), .ZN(
        n10676) );
  AOI211_X1 U11480 ( .C1(n10674), .C2(n10673), .A(n10672), .B(n10734), .ZN(
        n10675) );
  AOI211_X1 U11481 ( .C1(n10744), .C2(n10677), .A(n10676), .B(n10675), .ZN(
        n10678) );
  INV_X1 U11482 ( .A(n10678), .ZN(n10680) );
  AOI211_X1 U11483 ( .C1(n10942), .C2(P1_ADDR_REG_8__SCAN_IN), .A(n10680), .B(
        n10679), .ZN(n10681) );
  INV_X1 U11484 ( .A(n10681), .ZN(P1_U3251) );
  INV_X1 U11485 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n10693) );
  AOI211_X1 U11486 ( .C1(n10684), .C2(n10683), .A(n10682), .B(n10734), .ZN(
        n10689) );
  AOI211_X1 U11487 ( .C1(n10687), .C2(n10686), .A(n10685), .B(n10958), .ZN(
        n10688) );
  AOI211_X1 U11488 ( .C1(n10744), .C2(n10690), .A(n10689), .B(n10688), .ZN(
        n10692) );
  OAI211_X1 U11489 ( .C1(n10733), .C2(n10693), .A(n10692), .B(n10691), .ZN(
        P1_U3254) );
  INV_X1 U11490 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n10711) );
  NAND2_X1 U11491 ( .A1(n10695), .A2(n10694), .ZN(n10698) );
  INV_X1 U11492 ( .A(n10696), .ZN(n10697) );
  NAND2_X1 U11493 ( .A1(n10698), .A2(n10697), .ZN(n10707) );
  INV_X1 U11494 ( .A(n10699), .ZN(n10700) );
  OR2_X1 U11495 ( .A1(n10949), .A2(n10700), .ZN(n10706) );
  AOI21_X1 U11496 ( .B1(n10703), .B2(n10702), .A(n10701), .ZN(n10704) );
  NAND2_X1 U11497 ( .A1(n10954), .A2(n10704), .ZN(n10705) );
  OAI211_X1 U11498 ( .C1(n10958), .C2(n10707), .A(n10706), .B(n10705), .ZN(
        n10708) );
  INV_X1 U11499 ( .A(n10708), .ZN(n10710) );
  OAI211_X1 U11500 ( .C1(n10733), .C2(n10711), .A(n10710), .B(n10709), .ZN(
        P1_U3257) );
  INV_X1 U11501 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n10721) );
  AOI211_X1 U11502 ( .C1(n10713), .C2(n7993), .A(n10712), .B(n10734), .ZN(
        n10717) );
  AOI211_X1 U11503 ( .C1(n10715), .C2(n8038), .A(n10714), .B(n10958), .ZN(
        n10716) );
  AOI211_X1 U11504 ( .C1(n10744), .C2(n10718), .A(n10717), .B(n10716), .ZN(
        n10720) );
  OAI211_X1 U11505 ( .C1(n10733), .C2(n10721), .A(n10720), .B(n10719), .ZN(
        P1_U3258) );
  INV_X1 U11506 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n10732) );
  AOI211_X1 U11507 ( .C1(n10724), .C2(n10723), .A(n10734), .B(n10722), .ZN(
        n10729) );
  AOI211_X1 U11508 ( .C1(n10727), .C2(n10726), .A(n10958), .B(n10725), .ZN(
        n10728) );
  AOI211_X1 U11509 ( .C1(n10737), .C2(n10736), .A(n10735), .B(n10734), .ZN(
        n10742) );
  AOI211_X1 U11510 ( .C1(n10740), .C2(n10739), .A(n10738), .B(n10958), .ZN(
        n10741) );
  AOI211_X1 U11511 ( .C1(n10744), .C2(n10743), .A(n10742), .B(n10741), .ZN(
        n10745) );
  INV_X1 U11512 ( .A(n10745), .ZN(n10747) );
  AOI211_X1 U11513 ( .C1(n10942), .C2(P1_ADDR_REG_13__SCAN_IN), .A(n10747), 
        .B(n10746), .ZN(n10748) );
  INV_X1 U11514 ( .A(n10748), .ZN(P1_U3256) );
  AOI22_X1 U11515 ( .A1(n10749), .A2(n10896), .B1(n10895), .B2(
        P2_ADDR_REG_0__SCAN_IN), .ZN(n10754) );
  XNOR2_X1 U11516 ( .A(n10750), .B(n10749), .ZN(n10751) );
  OAI21_X1 U11517 ( .B1(n10904), .B2(n10752), .A(n10751), .ZN(n10753) );
  OAI211_X1 U11518 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n10755), .A(n10754), .B(
        n10753), .ZN(P2_U3182) );
  AND3_X1 U11519 ( .A1(n10758), .A2(n10757), .A3(n10756), .ZN(n10759) );
  OAI21_X1 U11520 ( .B1(n10760), .B2(n10759), .A(n10790), .ZN(n10768) );
  OAI21_X1 U11521 ( .B1(n10763), .B2(n10762), .A(n10761), .ZN(n10764) );
  NAND2_X1 U11522 ( .A1(n10905), .A2(n10764), .ZN(n10767) );
  AOI21_X1 U11523 ( .B1(n10896), .B2(n5358), .A(n10765), .ZN(n10766) );
  AND3_X1 U11524 ( .A1(n10768), .A2(n10767), .A3(n10766), .ZN(n10776) );
  AOI21_X1 U11525 ( .B1(n10771), .B2(n10770), .A(n10769), .ZN(n10773) );
  NOR2_X1 U11526 ( .A1(n10773), .A2(n10772), .ZN(n10774) );
  AOI21_X1 U11527 ( .B1(n10895), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n10774), .ZN(
        n10775) );
  NAND2_X1 U11528 ( .A1(n10776), .A2(n10775), .ZN(P2_U3188) );
  AOI22_X1 U11529 ( .A1(n10895), .A2(P2_ADDR_REG_10__SCAN_IN), .B1(n10777), 
        .B2(n10896), .ZN(n10796) );
  INV_X1 U11530 ( .A(n10778), .ZN(n10780) );
  NAND2_X1 U11531 ( .A1(n10780), .A2(n10779), .ZN(n10781) );
  XNOR2_X1 U11532 ( .A(n10782), .B(n10781), .ZN(n10787) );
  OAI21_X1 U11533 ( .B1(n10785), .B2(n10784), .A(n10783), .ZN(n10786) );
  AOI22_X1 U11534 ( .A1(n10787), .A2(n10904), .B1(n10905), .B2(n10786), .ZN(
        n10795) );
  NAND2_X1 U11535 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(P2_U3151), .ZN(n10794)
         );
  NOR2_X1 U11536 ( .A1(n10789), .A2(n10788), .ZN(n10792) );
  OAI21_X1 U11537 ( .B1(n10792), .B2(n10791), .A(n10790), .ZN(n10793) );
  NAND4_X1 U11538 ( .A1(n10796), .A2(n10795), .A3(n10794), .A4(n10793), .ZN(
        P2_U3192) );
  AOI22_X1 U11539 ( .A1(n10797), .A2(n10896), .B1(n10895), .B2(
        P2_ADDR_REG_11__SCAN_IN), .ZN(n10811) );
  OAI21_X1 U11540 ( .B1(n10800), .B2(n10799), .A(n10798), .ZN(n10804) );
  OAI21_X1 U11541 ( .B1(P2_REG1_REG_11__SCAN_IN), .B2(n10802), .A(n10801), 
        .ZN(n10803) );
  AOI22_X1 U11542 ( .A1(n10804), .A2(n10904), .B1(n10905), .B2(n10803), .ZN(
        n10810) );
  NAND2_X1 U11543 ( .A1(P2_REG3_REG_11__SCAN_IN), .A2(P2_U3151), .ZN(n10809)
         );
  AOI21_X1 U11544 ( .B1(n10806), .B2(n8890), .A(n10805), .ZN(n10807) );
  OR2_X1 U11545 ( .A1(n10807), .A2(n10910), .ZN(n10808) );
  NAND4_X1 U11546 ( .A1(n10811), .A2(n10810), .A3(n10809), .A4(n10808), .ZN(
        P2_U3193) );
  AOI22_X1 U11547 ( .A1(n10812), .A2(n10896), .B1(n10895), .B2(
        P2_ADDR_REG_12__SCAN_IN), .ZN(n10828) );
  OAI21_X1 U11548 ( .B1(n10815), .B2(n10814), .A(n10813), .ZN(n10820) );
  OAI21_X1 U11549 ( .B1(n10818), .B2(n10817), .A(n10816), .ZN(n10819) );
  AOI22_X1 U11550 ( .A1(n10820), .A2(n10905), .B1(n10904), .B2(n10819), .ZN(
        n10827) );
  INV_X1 U11551 ( .A(n10821), .ZN(n10826) );
  AOI21_X1 U11552 ( .B1(n5231), .B2(n10823), .A(n10822), .ZN(n10824) );
  OR2_X1 U11553 ( .A1(n10824), .A2(n10910), .ZN(n10825) );
  NAND4_X1 U11554 ( .A1(n10828), .A2(n10827), .A3(n10826), .A4(n10825), .ZN(
        P2_U3194) );
  AOI22_X1 U11555 ( .A1(n10829), .A2(n10896), .B1(n10895), .B2(
        P2_ADDR_REG_13__SCAN_IN), .ZN(n10844) );
  OAI21_X1 U11556 ( .B1(P2_REG1_REG_13__SCAN_IN), .B2(n10831), .A(n10830), 
        .ZN(n10836) );
  OAI21_X1 U11557 ( .B1(n10834), .B2(n10833), .A(n10832), .ZN(n10835) );
  AOI22_X1 U11558 ( .A1(n10836), .A2(n10905), .B1(n10904), .B2(n10835), .ZN(
        n10843) );
  INV_X1 U11559 ( .A(n10837), .ZN(n10842) );
  AOI21_X1 U11560 ( .B1(n10839), .B2(n8884), .A(n10838), .ZN(n10840) );
  OR2_X1 U11561 ( .A1(n10910), .A2(n10840), .ZN(n10841) );
  NAND4_X1 U11562 ( .A1(n10844), .A2(n10843), .A3(n10842), .A4(n10841), .ZN(
        P2_U3195) );
  AOI22_X1 U11563 ( .A1(n10895), .A2(P2_ADDR_REG_14__SCAN_IN), .B1(n10845), 
        .B2(n10896), .ZN(n10862) );
  XNOR2_X1 U11564 ( .A(n10847), .B(n10846), .ZN(n10852) );
  OAI21_X1 U11565 ( .B1(n10850), .B2(n10849), .A(n10848), .ZN(n10851) );
  AOI22_X1 U11566 ( .A1(n10852), .A2(n10905), .B1(n10904), .B2(n10851), .ZN(
        n10861) );
  INV_X1 U11567 ( .A(n10853), .ZN(n10860) );
  INV_X1 U11568 ( .A(n10854), .ZN(n10855) );
  AOI21_X1 U11569 ( .B1(n10857), .B2(n10856), .A(n10855), .ZN(n10858) );
  OR2_X1 U11570 ( .A1(n10858), .A2(n10910), .ZN(n10859) );
  NAND4_X1 U11571 ( .A1(n10862), .A2(n10861), .A3(n10860), .A4(n10859), .ZN(
        P2_U3196) );
  AOI22_X1 U11572 ( .A1(n10863), .A2(n10896), .B1(n10895), .B2(
        P2_ADDR_REG_15__SCAN_IN), .ZN(n10878) );
  OAI21_X1 U11573 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n10865), .A(n10864), 
        .ZN(n10870) );
  OAI21_X1 U11574 ( .B1(n10868), .B2(n10867), .A(n10866), .ZN(n10869) );
  AOI22_X1 U11575 ( .A1(n10870), .A2(n10905), .B1(n10904), .B2(n10869), .ZN(
        n10877) );
  INV_X1 U11576 ( .A(n10871), .ZN(n10876) );
  AOI21_X1 U11577 ( .B1(n10873), .B2(n8880), .A(n10872), .ZN(n10874) );
  OR2_X1 U11578 ( .A1(n10874), .A2(n10910), .ZN(n10875) );
  NAND4_X1 U11579 ( .A1(n10878), .A2(n10877), .A3(n10876), .A4(n10875), .ZN(
        P2_U3197) );
  AOI22_X1 U11580 ( .A1(n10879), .A2(n10896), .B1(n10895), .B2(
        P2_ADDR_REG_16__SCAN_IN), .ZN(n10894) );
  OAI21_X1 U11581 ( .B1(n10882), .B2(n10881), .A(n10880), .ZN(n10887) );
  OAI21_X1 U11582 ( .B1(n10885), .B2(n10884), .A(n10883), .ZN(n10886) );
  AOI22_X1 U11583 ( .A1(n10887), .A2(n10905), .B1(n10904), .B2(n10886), .ZN(
        n10893) );
  AOI21_X1 U11584 ( .B1(n10889), .B2(n10888), .A(n5222), .ZN(n10890) );
  OR2_X1 U11585 ( .A1(n10890), .A2(n10910), .ZN(n10891) );
  NAND4_X1 U11586 ( .A1(n10894), .A2(n10893), .A3(n10892), .A4(n10891), .ZN(
        P2_U3198) );
  AOI22_X1 U11587 ( .A1(n10897), .A2(n10896), .B1(n10895), .B2(
        P2_ADDR_REG_17__SCAN_IN), .ZN(n10914) );
  OAI21_X1 U11588 ( .B1(P2_REG1_REG_17__SCAN_IN), .B2(n10899), .A(n10898), 
        .ZN(n10906) );
  OAI21_X1 U11589 ( .B1(n10902), .B2(n10901), .A(n10900), .ZN(n10903) );
  AOI22_X1 U11590 ( .A1(n10906), .A2(n10905), .B1(n10904), .B2(n10903), .ZN(
        n10913) );
  AOI21_X1 U11591 ( .B1(n10908), .B2(n9144), .A(n10907), .ZN(n10909) );
  OR2_X1 U11592 ( .A1(n10910), .A2(n10909), .ZN(n10911) );
  NAND4_X1 U11593 ( .A1(n10914), .A2(n10913), .A3(n10912), .A4(n10911), .ZN(
        P2_U3199) );
  XNOR2_X1 U11594 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  AOI22_X1 U11595 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(n10942), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n10940) );
  NAND2_X1 U11596 ( .A1(n10916), .A2(n10915), .ZN(n10919) );
  INV_X1 U11597 ( .A(n10917), .ZN(n10918) );
  NAND2_X1 U11598 ( .A1(n10919), .A2(n10918), .ZN(n10927) );
  OR2_X1 U11599 ( .A1(n10949), .A2(n10920), .ZN(n10926) );
  AOI21_X1 U11600 ( .B1(n10923), .B2(n10922), .A(n10921), .ZN(n10924) );
  NAND2_X1 U11601 ( .A1(n10954), .A2(n10924), .ZN(n10925) );
  OAI211_X1 U11602 ( .C1(n10958), .C2(n10927), .A(n10926), .B(n10925), .ZN(
        n10928) );
  INV_X1 U11603 ( .A(n10928), .ZN(n10939) );
  INV_X1 U11604 ( .A(n10929), .ZN(n10936) );
  INV_X1 U11605 ( .A(n10935), .ZN(n10931) );
  OAI22_X1 U11606 ( .A1(n10931), .A2(n5247), .B1(n10930), .B2(n10588), .ZN(
        n10932) );
  OAI21_X1 U11607 ( .B1(n10933), .B2(n5145), .A(n10932), .ZN(n10934) );
  OAI21_X1 U11608 ( .B1(n10936), .B2(n10935), .A(n10934), .ZN(n10938) );
  NAND2_X1 U11609 ( .A1(n10938), .A2(n10937), .ZN(n10960) );
  NAND3_X1 U11610 ( .A1(n10940), .A2(n10939), .A3(n10960), .ZN(P1_U3245) );
  AOI21_X1 U11611 ( .B1(P1_ADDR_REG_4__SCAN_IN), .B2(n10942), .A(n10941), .ZN(
        n10962) );
  NAND2_X1 U11612 ( .A1(n10944), .A2(n10943), .ZN(n10947) );
  INV_X1 U11613 ( .A(n10945), .ZN(n10946) );
  NAND2_X1 U11614 ( .A1(n10947), .A2(n10946), .ZN(n10957) );
  OR2_X1 U11615 ( .A1(n10949), .A2(n10948), .ZN(n10956) );
  AOI21_X1 U11616 ( .B1(n10952), .B2(n10951), .A(n10950), .ZN(n10953) );
  NAND2_X1 U11617 ( .A1(n10954), .A2(n10953), .ZN(n10955) );
  OAI211_X1 U11618 ( .C1(n10958), .C2(n10957), .A(n10956), .B(n10955), .ZN(
        n10959) );
  INV_X1 U11619 ( .A(n10959), .ZN(n10961) );
  NAND3_X1 U11620 ( .A1(n10962), .A2(n10961), .A3(n10960), .ZN(P1_U3247) );
  INV_X1 U11621 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n10969) );
  NOR2_X1 U11622 ( .A1(n10963), .A2(n11107), .ZN(n10973) );
  INV_X1 U11623 ( .A(n10973), .ZN(n10967) );
  NOR2_X1 U11624 ( .A1(n10982), .A2(n10964), .ZN(n10974) );
  NAND2_X1 U11625 ( .A1(n10974), .A2(n10965), .ZN(n10966) );
  OAI211_X1 U11626 ( .C1(n10969), .C2(n10968), .A(n10967), .B(n10966), .ZN(
        n10970) );
  AOI21_X1 U11627 ( .B1(n10971), .B2(n10976), .A(n10970), .ZN(n10972) );
  AOI22_X1 U11628 ( .A1(n7171), .A2(n10588), .B1(n10972), .B2(n10358), .ZN(
        P1_U3293) );
  NAND2_X1 U11629 ( .A1(n11176), .A2(n11104), .ZN(n10975) );
  AOI211_X1 U11630 ( .C1(n10976), .C2(n10975), .A(n10974), .B(n10973), .ZN(
        n10977) );
  AOI22_X1 U11631 ( .A1(n11202), .A2(n10977), .B1(n10590), .B2(n11201), .ZN(
        P1_U3522) );
  AOI22_X1 U11632 ( .A1(n11206), .A2(n10977), .B1(n6794), .B2(n11203), .ZN(
        P1_U3453) );
  INV_X1 U11633 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n10978) );
  AOI22_X1 U11634 ( .A1(n11186), .A2(n10979), .B1(n10978), .B2(n6448), .ZN(
        P2_U3393) );
  INV_X1 U11635 ( .A(n11091), .ZN(n11071) );
  XNOR2_X1 U11636 ( .A(n10985), .B(n10980), .ZN(n10994) );
  OAI211_X1 U11637 ( .C1(n10983), .C2(n10982), .A(n5131), .B(n10981), .ZN(
        n10997) );
  OAI21_X1 U11638 ( .B1(n10983), .B2(n11195), .A(n10997), .ZN(n10991) );
  INV_X1 U11639 ( .A(n10984), .ZN(n11095) );
  XNOR2_X1 U11640 ( .A(n10986), .B(n10985), .ZN(n10988) );
  AOI22_X1 U11641 ( .A1(n11172), .A2(n7175), .B1(n11020), .B2(n11169), .ZN(
        n10987) );
  OAI21_X1 U11642 ( .B1(n10988), .B2(n11104), .A(n10987), .ZN(n10989) );
  AOI21_X1 U11643 ( .B1(n11095), .B2(n10994), .A(n10989), .ZN(n11005) );
  INV_X1 U11644 ( .A(n11005), .ZN(n10990) );
  AOI211_X1 U11645 ( .C1(n11071), .C2(n10994), .A(n10991), .B(n10990), .ZN(
        n10993) );
  AOI22_X1 U11646 ( .A1(n11202), .A2(n10993), .B1(n10992), .B2(n11201), .ZN(
        P1_U3523) );
  AOI22_X1 U11647 ( .A1(n11206), .A2(n10993), .B1(n6761), .B2(n11203), .ZN(
        P1_U3456) );
  AOI22_X1 U11648 ( .A1(n11123), .A2(P1_REG3_REG_1__SCAN_IN), .B1(
        P1_REG2_REG_1__SCAN_IN), .B2(n7171), .ZN(n11004) );
  INV_X1 U11649 ( .A(n10994), .ZN(n11001) );
  INV_X1 U11650 ( .A(n10995), .ZN(n10996) );
  NAND2_X1 U11651 ( .A1(n10367), .A2(n10996), .ZN(n11076) );
  INV_X1 U11652 ( .A(n10997), .ZN(n10998) );
  NAND2_X1 U11653 ( .A1(n11128), .A2(n10998), .ZN(n11000) );
  NAND2_X1 U11654 ( .A1(n11124), .A2(n9409), .ZN(n10999) );
  OAI211_X1 U11655 ( .C1(n11001), .C2(n11076), .A(n11000), .B(n10999), .ZN(
        n11002) );
  INV_X1 U11656 ( .A(n11002), .ZN(n11003) );
  OAI211_X1 U11657 ( .C1(n7171), .C2(n11005), .A(n11004), .B(n11003), .ZN(
        P1_U3292) );
  AOI22_X1 U11658 ( .A1(n11172), .A2(n11007), .B1(n5142), .B2(n11169), .ZN(
        n11008) );
  OAI211_X1 U11659 ( .C1(n11010), .C2(n11195), .A(n11009), .B(n11008), .ZN(
        n11013) );
  NOR2_X1 U11660 ( .A1(n11011), .A2(n11104), .ZN(n11012) );
  AOI211_X1 U11661 ( .C1(n11199), .C2(n11014), .A(n11013), .B(n11012), .ZN(
        n11016) );
  AOI22_X1 U11662 ( .A1(n11202), .A2(n11016), .B1(n11015), .B2(n11201), .ZN(
        P1_U3524) );
  AOI22_X1 U11663 ( .A1(n11206), .A2(n11016), .B1(n6897), .B2(n11203), .ZN(
        P1_U3459) );
  INV_X1 U11664 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n11017) );
  AOI22_X1 U11665 ( .A1(n11186), .A2(n11018), .B1(n11017), .B2(n6448), .ZN(
        P2_U3396) );
  INV_X1 U11666 ( .A(n11027), .ZN(n11029) );
  AOI22_X1 U11667 ( .A1(n11172), .A2(n11020), .B1(n11019), .B2(n11169), .ZN(
        n11021) );
  OAI211_X1 U11668 ( .C1(n11023), .C2(n11195), .A(n11022), .B(n11021), .ZN(
        n11024) );
  INV_X1 U11669 ( .A(n11024), .ZN(n11026) );
  OAI211_X1 U11670 ( .C1(n11027), .C2(n11091), .A(n11026), .B(n11025), .ZN(
        n11028) );
  AOI21_X1 U11671 ( .B1(n11095), .B2(n11029), .A(n11028), .ZN(n11030) );
  AOI22_X1 U11672 ( .A1(n11202), .A2(n11030), .B1(n6967), .B2(n11201), .ZN(
        P1_U3525) );
  AOI22_X1 U11673 ( .A1(n11206), .A2(n11030), .B1(n6965), .B2(n11203), .ZN(
        P1_U3462) );
  INV_X1 U11674 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n11031) );
  AOI22_X1 U11675 ( .A1(n11186), .A2(n11032), .B1(n11031), .B2(n6448), .ZN(
        P2_U3399) );
  INV_X1 U11676 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n11033) );
  AOI22_X1 U11677 ( .A1(n11186), .A2(n11034), .B1(n11033), .B2(n6448), .ZN(
        P2_U3402) );
  OAI22_X1 U11678 ( .A1(n11036), .A2(n11109), .B1(n11035), .B2(n11107), .ZN(
        n11038) );
  AOI211_X1 U11679 ( .C1(n11147), .C2(n7004), .A(n11038), .B(n11037), .ZN(
        n11039) );
  OAI21_X1 U11680 ( .B1(n11040), .B2(n11176), .A(n11039), .ZN(n11041) );
  AOI21_X1 U11681 ( .B1(n11042), .B2(n11181), .A(n11041), .ZN(n11043) );
  AOI22_X1 U11682 ( .A1(n11202), .A2(n11043), .B1(n6865), .B2(n11201), .ZN(
        P1_U3526) );
  AOI22_X1 U11683 ( .A1(n11206), .A2(n11043), .B1(n6979), .B2(n11203), .ZN(
        P1_U3465) );
  INV_X1 U11684 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n11044) );
  AOI22_X1 U11685 ( .A1(n11186), .A2(n11045), .B1(n11044), .B2(n6448), .ZN(
        P2_U3405) );
  OAI22_X1 U11686 ( .A1(n11046), .A2(n11109), .B1(n11085), .B2(n11107), .ZN(
        n11047) );
  AOI21_X1 U11687 ( .B1(n11147), .B2(n11048), .A(n11047), .ZN(n11050) );
  OAI211_X1 U11688 ( .C1(n11051), .C2(n11176), .A(n11050), .B(n11049), .ZN(
        n11052) );
  AOI21_X1 U11689 ( .B1(n11053), .B2(n11181), .A(n11052), .ZN(n11054) );
  AOI22_X1 U11690 ( .A1(n11202), .A2(n11054), .B1(n7022), .B2(n11201), .ZN(
        P1_U3527) );
  AOI22_X1 U11691 ( .A1(n11206), .A2(n11054), .B1(n7023), .B2(n11203), .ZN(
        P1_U3468) );
  INV_X1 U11692 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n11055) );
  AOI22_X1 U11693 ( .A1(n11186), .A2(n11056), .B1(n11055), .B2(n6448), .ZN(
        P2_U3408) );
  XNOR2_X1 U11694 ( .A(n11057), .B(n11062), .ZN(n11080) );
  INV_X1 U11695 ( .A(n11058), .ZN(n11060) );
  OAI211_X1 U11696 ( .C1(n11060), .C2(n11061), .A(n5131), .B(n11059), .ZN(
        n11077) );
  OAI21_X1 U11697 ( .B1(n11061), .B2(n11195), .A(n11077), .ZN(n11070) );
  XNOR2_X1 U11698 ( .A(n11063), .B(n11062), .ZN(n11067) );
  AOI22_X1 U11699 ( .A1(n11065), .A2(n11169), .B1(n11172), .B2(n11064), .ZN(
        n11066) );
  OAI21_X1 U11700 ( .B1(n11067), .B2(n11104), .A(n11066), .ZN(n11068) );
  AOI21_X1 U11701 ( .B1(n11080), .B2(n11095), .A(n11068), .ZN(n11083) );
  INV_X1 U11702 ( .A(n11083), .ZN(n11069) );
  AOI211_X1 U11703 ( .C1(n11071), .C2(n11080), .A(n11070), .B(n11069), .ZN(
        n11072) );
  AOI22_X1 U11704 ( .A1(n11202), .A2(n11072), .B1(n6870), .B2(n11201), .ZN(
        P1_U3528) );
  AOI22_X1 U11705 ( .A1(n11206), .A2(n11072), .B1(n7299), .B2(n11203), .ZN(
        P1_U3471) );
  INV_X1 U11706 ( .A(n11073), .ZN(n11074) );
  AOI222_X1 U11707 ( .A1(n11075), .A2(n11124), .B1(P1_REG2_REG_6__SCAN_IN), 
        .B2(n7171), .C1(n11123), .C2(n11074), .ZN(n11082) );
  INV_X1 U11708 ( .A(n11076), .ZN(n11079) );
  INV_X1 U11709 ( .A(n11077), .ZN(n11078) );
  AOI22_X1 U11710 ( .A1(n11080), .A2(n11079), .B1(n11128), .B2(n11078), .ZN(
        n11081) );
  OAI211_X1 U11711 ( .C1(n7171), .C2(n11083), .A(n11082), .B(n11081), .ZN(
        P1_U3287) );
  INV_X1 U11712 ( .A(n11092), .ZN(n11094) );
  OAI22_X1 U11713 ( .A1(n11085), .A2(n11109), .B1(n11084), .B2(n11107), .ZN(
        n11087) );
  AOI211_X1 U11714 ( .C1(n11147), .C2(n11088), .A(n11087), .B(n11086), .ZN(
        n11090) );
  OAI211_X1 U11715 ( .C1(n11092), .C2(n11091), .A(n11090), .B(n11089), .ZN(
        n11093) );
  AOI21_X1 U11716 ( .B1(n11095), .B2(n11094), .A(n11093), .ZN(n11097) );
  INV_X1 U11717 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n11096) );
  AOI22_X1 U11718 ( .A1(n11202), .A2(n11097), .B1(n11096), .B2(n11201), .ZN(
        P1_U3529) );
  AOI22_X1 U11719 ( .A1(n11206), .A2(n11097), .B1(n7337), .B2(n11203), .ZN(
        P1_U3474) );
  XNOR2_X1 U11720 ( .A(n11099), .B(n11098), .ZN(n11130) );
  INV_X1 U11721 ( .A(n11100), .ZN(n11106) );
  AOI21_X1 U11722 ( .B1(n11103), .B2(n11102), .A(n11101), .ZN(n11105) );
  NOR3_X1 U11723 ( .A1(n11106), .A2(n11105), .A3(n11104), .ZN(n11112) );
  OAI22_X1 U11724 ( .A1(n11110), .A2(n11109), .B1(n11108), .B2(n11107), .ZN(
        n11111) );
  NOR2_X1 U11725 ( .A1(n11112), .A2(n11111), .ZN(n11133) );
  INV_X1 U11726 ( .A(n11113), .ZN(n11115) );
  OAI211_X1 U11727 ( .C1(n11117), .C2(n11116), .A(n11115), .B(n5131), .ZN(
        n11126) );
  OAI211_X1 U11728 ( .C1(n11117), .C2(n11195), .A(n11133), .B(n11126), .ZN(
        n11118) );
  AOI21_X1 U11729 ( .B1(n11199), .B2(n11130), .A(n11118), .ZN(n11120) );
  AOI22_X1 U11730 ( .A1(n11202), .A2(n11120), .B1(n7411), .B2(n11201), .ZN(
        P1_U3530) );
  INV_X1 U11731 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n11119) );
  AOI22_X1 U11732 ( .A1(n11206), .A2(n11120), .B1(n11119), .B2(n11203), .ZN(
        P1_U3477) );
  INV_X1 U11733 ( .A(n11121), .ZN(n11122) );
  AOI222_X1 U11734 ( .A1(n11125), .A2(n11124), .B1(P1_REG2_REG_8__SCAN_IN), 
        .B2(n7171), .C1(n11123), .C2(n11122), .ZN(n11132) );
  INV_X1 U11735 ( .A(n11126), .ZN(n11127) );
  AOI22_X1 U11736 ( .A1(n11130), .A2(n11129), .B1(n11128), .B2(n11127), .ZN(
        n11131) );
  OAI211_X1 U11737 ( .C1(n7171), .C2(n11133), .A(n11132), .B(n11131), .ZN(
        P1_U3285) );
  INV_X1 U11738 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n11134) );
  AOI22_X1 U11739 ( .A1(n11186), .A2(n11135), .B1(n11134), .B2(n6448), .ZN(
        P2_U3414) );
  AOI22_X1 U11740 ( .A1(n11137), .A2(n11147), .B1(n11172), .B2(n11136), .ZN(
        n11138) );
  OAI211_X1 U11741 ( .C1(n11140), .C2(n11176), .A(n11139), .B(n11138), .ZN(
        n11141) );
  AOI21_X1 U11742 ( .B1(n11181), .B2(n11142), .A(n11141), .ZN(n11145) );
  AOI22_X1 U11743 ( .A1(n11202), .A2(n11145), .B1(n11143), .B2(n11201), .ZN(
        P1_U3531) );
  INV_X1 U11744 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n11144) );
  AOI22_X1 U11745 ( .A1(n11206), .A2(n11145), .B1(n11144), .B2(n11203), .ZN(
        P1_U3480) );
  AOI22_X1 U11746 ( .A1(n11148), .A2(n11147), .B1(n11169), .B2(n11146), .ZN(
        n11150) );
  NAND3_X1 U11747 ( .A1(n11151), .A2(n11150), .A3(n11149), .ZN(n11152) );
  AOI21_X1 U11748 ( .B1(n11153), .B2(n11199), .A(n11152), .ZN(n11155) );
  AOI22_X1 U11749 ( .A1(n11202), .A2(n11155), .B1(n11154), .B2(n11201), .ZN(
        P1_U3532) );
  AOI22_X1 U11750 ( .A1(n11206), .A2(n11155), .B1(n6558), .B2(n11203), .ZN(
        P1_U3483) );
  AOI22_X1 U11751 ( .A1(n11186), .A2(n11156), .B1(n6042), .B2(n6448), .ZN(
        P2_U3420) );
  INV_X1 U11752 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n11157) );
  AOI22_X1 U11753 ( .A1(n11186), .A2(n11158), .B1(n11157), .B2(n6448), .ZN(
        P2_U3423) );
  INV_X1 U11754 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n11159) );
  AOI22_X1 U11755 ( .A1(n11186), .A2(n11160), .B1(n11159), .B2(n6448), .ZN(
        P2_U3426) );
  OAI211_X1 U11756 ( .C1(n11163), .C2(n11195), .A(n11162), .B(n11161), .ZN(
        n11164) );
  AOI21_X1 U11757 ( .B1(n11165), .B2(n11199), .A(n11164), .ZN(n11168) );
  AOI22_X1 U11758 ( .A1(n11202), .A2(n11168), .B1(n11166), .B2(n11201), .ZN(
        P1_U3534) );
  INV_X1 U11759 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n11167) );
  AOI22_X1 U11760 ( .A1(n11206), .A2(n11168), .B1(n11167), .B2(n11203), .ZN(
        P1_U3489) );
  AOI22_X1 U11761 ( .A1(n11172), .A2(n11171), .B1(n11170), .B2(n11169), .ZN(
        n11173) );
  OAI211_X1 U11762 ( .C1(n11175), .C2(n11195), .A(n11174), .B(n11173), .ZN(
        n11179) );
  NOR2_X1 U11763 ( .A1(n11177), .A2(n11176), .ZN(n11178) );
  AOI211_X1 U11764 ( .C1(n11181), .C2(n11180), .A(n11179), .B(n11178), .ZN(
        n11183) );
  AOI22_X1 U11765 ( .A1(n11202), .A2(n11183), .B1(n10111), .B2(n11201), .ZN(
        P1_U3535) );
  INV_X1 U11766 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n11182) );
  AOI22_X1 U11767 ( .A1(n11206), .A2(n11183), .B1(n11182), .B2(n11203), .ZN(
        P1_U3492) );
  INV_X1 U11768 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n11184) );
  AOI22_X1 U11769 ( .A1(n11186), .A2(n11185), .B1(n11184), .B2(n6448), .ZN(
        P2_U3429) );
  OAI21_X1 U11770 ( .B1(n11188), .B2(n11195), .A(n11187), .ZN(n11189) );
  AOI211_X1 U11771 ( .C1(n11191), .C2(n11199), .A(n11190), .B(n11189), .ZN(
        n11193) );
  AOI22_X1 U11772 ( .A1(n11202), .A2(n11193), .B1(n7993), .B2(n11201), .ZN(
        P1_U3537) );
  INV_X1 U11773 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n11192) );
  AOI22_X1 U11774 ( .A1(n11206), .A2(n11193), .B1(n11192), .B2(n11203), .ZN(
        P1_U3498) );
  OAI21_X1 U11775 ( .B1(n11196), .B2(n11195), .A(n11194), .ZN(n11197) );
  AOI211_X1 U11776 ( .C1(n11200), .C2(n11199), .A(n11198), .B(n11197), .ZN(
        n11205) );
  AOI22_X1 U11777 ( .A1(n11202), .A2(n11205), .B1(n8019), .B2(n11201), .ZN(
        P1_U3538) );
  INV_X1 U11778 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n11204) );
  AOI22_X1 U11779 ( .A1(n11206), .A2(n11205), .B1(n11204), .B2(n11203), .ZN(
        P1_U3501) );
  XNOR2_X1 U11780 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  OAI21_X1 U6659 ( .B1(n7399), .B2(n9557), .A(n5697), .ZN(n11057) );
  AOI21_X1 U6660 ( .B1(n11057), .B2(n11062), .A(n5696), .ZN(n7552) );
  CLKBUF_X1 U5202 ( .A(n5889), .Z(n5136) );
  CLKBUF_X1 U5211 ( .A(n5914), .Z(n6310) );
  INV_X1 U5212 ( .A(n6070), .ZN(n8468) );
  NAND2_X1 U5231 ( .A1(n6380), .A2(n5481), .ZN(n6348) );
  INV_X1 U5249 ( .A(n5143), .ZN(n6762) );
  CLKBUF_X1 U5269 ( .A(n5912), .Z(n6479) );
  CLKBUF_X1 U5324 ( .A(n6787), .Z(n5145) );
  OR2_X1 U5330 ( .A1(n10964), .A2(n9652), .ZN(n11212) );
endmodule

