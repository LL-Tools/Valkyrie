

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2134, n2135, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030;

  XNOR2_X1 U2376 ( .A(n2579), .B(n4978), .ZN(n4883) );
  CLKBUF_X2 U2377 ( .A(n2681), .Z(n3089) );
  OR2_X1 U2378 ( .A1(n3130), .A2(n3621), .ZN(n3135) );
  AOI21_X1 U2379 ( .B1(n3266), .B2(REG2_REG_6__SCAN_IN), .A(n2465), .ZN(n3291)
         );
  NAND4_X1 U2380 ( .A1(n2734), .A2(n2733), .A3(n2732), .A4(n2731), .ZN(n3511)
         );
  NAND4_X1 U2381 ( .A1(n2659), .A2(n2658), .A3(n2657), .A4(n2656), .ZN(n4936)
         );
  INV_X1 U2382 ( .A(n2767), .ZN(n2645) );
  AND2_X1 U2383 ( .A1(n3457), .A2(n2786), .ZN(n3849) );
  INV_X2 U2384 ( .A(n3006), .ZN(n3038) );
  OR2_X1 U2385 ( .A1(n4883), .A2(n2578), .ZN(n2586) );
  CLKBUF_X3 U2386 ( .A(n2680), .Z(n3040) );
  XNOR2_X1 U2388 ( .A(n2560), .B(n3227), .ZN(n4843) );
  OAI211_X1 U2389 ( .C1(n2210), .C2(n2208), .A(n3141), .B(n2207), .ZN(n3659)
         );
  CLKBUF_X3 U2390 ( .A(n2735), .Z(n2134) );
  AND4_X1 U2391 ( .A1(n2677), .A2(n2676), .A3(n2675), .A4(n2674), .ZN(n3121)
         );
  AOI21_X1 U2392 ( .B1(n4843), .B2(REG1_REG_4__SCAN_IN), .A(n2561), .ZN(n3279)
         );
  INV_X2 U2394 ( .A(n2532), .ZN(n2408) );
  NOR2_X2 U2395 ( .A1(n3537), .A2(n2416), .ZN(n2573) );
  XNOR2_X2 U2396 ( .A(n2476), .B(n4983), .ZN(n4859) );
  XNOR2_X2 U2397 ( .A(n2625), .B(IR_REG_30__SCAN_IN), .ZN(n2629) );
  XNOR2_X2 U2398 ( .A(n2514), .B(IR_REG_26__SCAN_IN), .ZN(n3244) );
  NOR2_X2 U2399 ( .A1(n3291), .A2(n3290), .ZN(n3289) );
  AND2_X1 U2400 ( .A1(n4292), .A2(n2623), .ZN(n3109) );
  CLKBUF_X2 U2401 ( .A(n2748), .Z(n3037) );
  XNOR2_X1 U2402 ( .A(n2520), .B(IR_REG_22__SCAN_IN), .ZN(n4828) );
  XNOR2_X1 U2403 ( .A(n2256), .B(n2626), .ZN(n2631) );
  INV_X1 U2404 ( .A(IR_REG_23__SCAN_IN), .ZN(n4003) );
  OR2_X1 U2405 ( .A1(n4634), .A2(n4411), .ZN(n3202) );
  OAI21_X1 U2406 ( .B1(n4863), .B2(n2362), .A(n2361), .ZN(n4871) );
  NAND3_X1 U2407 ( .A1(n2367), .A2(n2180), .A3(n2366), .ZN(n2484) );
  OR2_X1 U2408 ( .A1(n4853), .A2(n2571), .ZN(n2335) );
  AND2_X1 U2409 ( .A1(n3367), .A2(n3357), .ZN(n3457) );
  OR2_X1 U2410 ( .A1(n2568), .A2(n2566), .ZN(n2569) );
  NAND3_X1 U2411 ( .A1(n2346), .A2(n2345), .A3(n2347), .ZN(n2567) );
  NAND2_X1 U2412 ( .A1(n4932), .A2(n4933), .ZN(n4931) );
  NAND2_X2 U2413 ( .A1(n3419), .A2(n4691), .ZN(n4958) );
  XNOR2_X1 U2414 ( .A(n2464), .B(n4833), .ZN(n3266) );
  AND2_X1 U2415 ( .A1(n2344), .A2(n2171), .ZN(n2464) );
  NAND2_X1 U2416 ( .A1(n3164), .A2(n2302), .ZN(n4929) );
  INV_X1 U2417 ( .A(n2680), .ZN(n3009) );
  NAND2_X1 U2418 ( .A1(n4296), .A2(n4298), .ZN(n4703) );
  OAI211_X1 U2419 ( .C1(n2341), .C2(n2339), .A(n2342), .B(n2336), .ZN(n2344)
         );
  CLKBUF_X3 U2420 ( .A(n3168), .Z(n2135) );
  NAND4_X2 U2422 ( .A1(n2636), .A2(n2635), .A3(n2634), .A4(n2633), .ZN(n3119)
         );
  OR2_X1 U2423 ( .A1(n2137), .A2(n2627), .ZN(n2636) );
  INV_X1 U2424 ( .A(n2739), .ZN(n3033) );
  NAND2_X1 U2425 ( .A1(n3063), .A2(n4829), .ZN(n3422) );
  BUF_X4 U2426 ( .A(n2726), .Z(n2137) );
  NAND2_X1 U2427 ( .A1(n2203), .A2(n4827), .ZN(n2726) );
  XNOR2_X1 U2428 ( .A(n2557), .B(n3264), .ZN(n3258) );
  XNOR2_X1 U2429 ( .A(n2622), .B(n2621), .ZN(n3063) );
  NAND2_X2 U2430 ( .A1(n2629), .A2(n4827), .ZN(n2767) );
  INV_X1 U2431 ( .A(n2631), .ZN(n4827) );
  NAND2_X1 U2432 ( .A1(n2620), .A2(n2607), .ZN(n4433) );
  NAND2_X1 U2433 ( .A1(n2620), .A2(IR_REG_31__SCAN_IN), .ZN(n2622) );
  INV_X1 U2434 ( .A(n3276), .ZN(n2342) );
  NAND2_X1 U2435 ( .A1(n2258), .A2(n2257), .ZN(n2735) );
  BUF_X1 U2436 ( .A(n2631), .Z(n2632) );
  NAND2_X1 U2437 ( .A1(n2513), .A2(IR_REG_31__SCAN_IN), .ZN(n2514) );
  NAND2_X1 U2438 ( .A1(n2606), .A2(n2605), .ZN(n2620) );
  NAND2_X1 U2439 ( .A1(n2604), .A2(IR_REG_31__SCAN_IN), .ZN(n2606) );
  OR2_X1 U2440 ( .A1(n2521), .A2(IR_REG_21__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U2441 ( .A1(n3230), .A2(IR_REG_31__SCAN_IN), .ZN(n2625) );
  OAI21_X1 U2442 ( .B1(n2521), .B2(n2507), .A(IR_REG_31__SCAN_IN), .ZN(n2519)
         );
  AND2_X1 U2443 ( .A1(n2512), .A2(n2533), .ZN(n2526) );
  AND2_X1 U2444 ( .A1(n2530), .A2(n2528), .ZN(n2409) );
  AND4_X1 U2445 ( .A1(n2430), .A2(n2429), .A3(n2428), .A4(n2427), .ZN(n2530)
         );
  INV_X1 U2446 ( .A(IR_REG_29__SCAN_IN), .ZN(n2626) );
  INV_X1 U2447 ( .A(IR_REG_3__SCAN_IN), .ZN(n2453) );
  NOR2_X1 U2448 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2600)
         );
  INV_X1 U2449 ( .A(IR_REG_4__SCAN_IN), .ZN(n2456) );
  INV_X1 U2450 ( .A(IR_REG_2__SCAN_IN), .ZN(n2442) );
  NOR2_X1 U2451 ( .A1(IR_REG_24__SCAN_IN), .A2(IR_REG_22__SCAN_IN), .ZN(n2515)
         );
  NOR2_X1 U2452 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2430)
         );
  NOR2_X1 U2453 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2429)
         );
  NOR2_X1 U2454 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2428)
         );
  NOR2_X1 U2455 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2427)
         );
  INV_X1 U2456 ( .A(IR_REG_1__SCAN_IN), .ZN(n2377) );
  NOR2_X2 U2457 ( .A1(n3346), .A2(n2751), .ZN(n3356) );
  NOR2_X1 U2458 ( .A1(n4854), .A2(n4855), .ZN(n4853) );
  NAND2_X2 U2459 ( .A1(n2406), .A2(n2405), .ZN(n3886) );
  OR2_X2 U2460 ( .A1(n3909), .A2(n2418), .ZN(n2406) );
  XNOR2_X1 U2461 ( .A(n2562), .B(n4833), .ZN(n3265) );
  OAI21_X1 U2462 ( .B1(n2830), .B2(n3486), .A(n2724), .ZN(n2725) );
  OAI211_X1 U2463 ( .C1(n4273), .C2(n4271), .A(n4270), .B(n4272), .ZN(n3014)
         );
  OAI21_X2 U2464 ( .B1(n3550), .B2(n2394), .A(n2393), .ZN(n3862) );
  NAND2_X2 U2465 ( .A1(n2820), .A2(n3499), .ZN(n3550) );
  INV_X1 U2466 ( .A(n3119), .ZN(n4940) );
  INV_X2 U2467 ( .A(n2852), .ZN(n2830) );
  XNOR2_X2 U2468 ( .A(n2508), .B(IR_REG_24__SCAN_IN), .ZN(n3047) );
  XNOR2_X2 U2469 ( .A(n2517), .B(IR_REG_25__SCAN_IN), .ZN(n3045) );
  AOI21_X2 U2470 ( .B1(n3886), .B2(n2420), .A(n2985), .ZN(n4273) );
  AND2_X1 U2471 ( .A1(n2317), .A2(n3144), .ZN(n2316) );
  NAND2_X1 U2472 ( .A1(n3143), .A2(n3142), .ZN(n2317) );
  NAND2_X1 U2473 ( .A1(n4505), .A2(n3216), .ZN(n4502) );
  NAND2_X1 U2474 ( .A1(n2539), .A2(n2537), .ZN(n2257) );
  NAND2_X1 U2475 ( .A1(n2538), .A2(IR_REG_28__SCAN_IN), .ZN(n2258) );
  OR2_X1 U2476 ( .A1(n3026), .A2(n3990), .ZN(n4513) );
  INV_X1 U2477 ( .A(n2629), .ZN(n2203) );
  OR2_X1 U2478 ( .A1(n4872), .A2(n4864), .ZN(n2362) );
  INV_X1 U2479 ( .A(n4872), .ZN(n2360) );
  AND2_X1 U2480 ( .A1(n2221), .A2(n2177), .ZN(n2220) );
  NAND2_X1 U2481 ( .A1(n2218), .A2(n3160), .ZN(n2217) );
  INV_X1 U2482 ( .A(n2316), .ZN(n2314) );
  NAND2_X1 U2483 ( .A1(n3332), .A2(n2556), .ZN(n2557) );
  NOR2_X1 U2484 ( .A1(n2986), .A2(n4043), .ZN(n2995) );
  NAND2_X1 U2485 ( .A1(n4578), .A2(n4413), .ZN(n2243) );
  INV_X1 U2486 ( .A(n2943), .ZN(n2941) );
  AND2_X1 U2487 ( .A1(n2206), .A2(n2182), .ZN(n3760) );
  NAND2_X1 U2488 ( .A1(n3789), .A2(n3150), .ZN(n2206) );
  AND2_X1 U2489 ( .A1(n3140), .A2(n2170), .ZN(n2212) );
  INV_X1 U2490 ( .A(n2777), .ZN(n2283) );
  INV_X1 U2491 ( .A(n2224), .ZN(n2223) );
  OAI22_X1 U2492 ( .A1(n2225), .A2(n4703), .B1(n3559), .B2(n3121), .ZN(n2224)
         );
  NAND2_X1 U2493 ( .A1(n2160), .A2(n3120), .ZN(n2225) );
  XNOR2_X1 U2494 ( .A(n2652), .B(n3006), .ZN(n2669) );
  OR2_X1 U2495 ( .A1(n2876), .A2(n3734), .ZN(n2888) );
  INV_X1 U2496 ( .A(n2137), .ZN(n3028) );
  NOR2_X1 U2497 ( .A1(n3277), .A2(n2417), .ZN(n2562) );
  NAND2_X1 U2498 ( .A1(n4859), .A2(n2368), .ZN(n2367) );
  AND2_X1 U2499 ( .A1(n2369), .A2(REG2_REG_10__SCAN_IN), .ZN(n2368) );
  NAND2_X1 U2500 ( .A1(n2365), .A2(n2369), .ZN(n2366) );
  INV_X1 U2501 ( .A(n3542), .ZN(n2365) );
  AND2_X1 U2502 ( .A1(n2828), .A2(REG1_REG_13__SCAN_IN), .ZN(n2577) );
  OR2_X1 U2503 ( .A1(n2828), .A2(REG2_REG_13__SCAN_IN), .ZN(n2359) );
  NAND2_X1 U2504 ( .A1(n4499), .A2(n4506), .ZN(n2269) );
  NAND2_X1 U2505 ( .A1(n2152), .A2(n2323), .ZN(n2322) );
  NAND2_X1 U2506 ( .A1(n2324), .A2(n3162), .ZN(n2323) );
  INV_X1 U2507 ( .A(n4358), .ZN(n2324) );
  AND2_X1 U2508 ( .A1(n4657), .A2(n4643), .ZN(n3153) );
  AND4_X1 U2509 ( .A1(n2827), .A2(n2826), .A3(n2825), .A4(n2824), .ZN(n3689)
         );
  AND2_X1 U2510 ( .A1(n4510), .A2(n4509), .ZN(n4511) );
  NOR2_X1 U2511 ( .A1(n2320), .A2(n2319), .ZN(n4718) );
  NAND2_X1 U2512 ( .A1(n4353), .A2(n2322), .ZN(n2319) );
  NAND2_X1 U2513 ( .A1(n3215), .A2(n3216), .ZN(n4499) );
  NAND2_X1 U2514 ( .A1(n4699), .A2(n4998), .ZN(n5017) );
  AOI21_X1 U2515 ( .B1(n3086), .B2(n2645), .A(n3085), .ZN(n4355) );
  OAI21_X1 U2516 ( .B1(n2145), .B2(n3224), .A(n2268), .ZN(n2262) );
  NAND2_X1 U2517 ( .A1(n3224), .A2(REG1_REG_29__SCAN_IN), .ZN(n2268) );
  OR2_X1 U2518 ( .A1(n4936), .A2(n4947), .ZN(n4293) );
  AOI21_X1 U2519 ( .B1(n2316), .B2(n2313), .A(n2162), .ZN(n2312) );
  INV_X1 U2520 ( .A(n3142), .ZN(n2313) );
  AND2_X1 U2521 ( .A1(n2964), .A2(n2963), .ZN(n2981) );
  OR2_X1 U2522 ( .A1(n2134), .A2(n3024), .ZN(n4345) );
  NOR2_X1 U2523 ( .A1(n2300), .A2(n2942), .ZN(n2299) );
  AND2_X1 U2524 ( .A1(n2247), .A2(n2169), .ZN(n2246) );
  NOR2_X1 U2525 ( .A1(n4406), .A2(n2248), .ZN(n2247) );
  INV_X1 U2526 ( .A(n4404), .ZN(n2248) );
  NOR2_X1 U2527 ( .A1(n3177), .A2(n4312), .ZN(n2410) );
  NAND2_X1 U2528 ( .A1(n4301), .A2(n4302), .ZN(n2251) );
  OR2_X1 U2529 ( .A1(n3116), .A2(n3115), .ZN(n2302) );
  NAND2_X1 U2530 ( .A1(n3101), .A2(n3721), .ZN(n2282) );
  AND2_X1 U2531 ( .A1(n3767), .A2(n3764), .ZN(n3101) );
  OR2_X1 U2532 ( .A1(n2282), .A2(n3902), .ZN(n2281) );
  AND2_X1 U2533 ( .A1(n3579), .A2(n4683), .ZN(n2275) );
  OR2_X1 U2534 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_22__SCAN_IN), .ZN(n2507)
         );
  INV_X1 U2535 ( .A(IR_REG_6__SCAN_IN), .ZN(n2436) );
  AND2_X1 U2536 ( .A1(n3887), .A2(n3885), .ZN(n2407) );
  NAND2_X1 U2537 ( .A1(n2382), .A2(n2381), .ZN(n4234) );
  AOI21_X1 U2538 ( .B1(n2384), .B2(n2387), .A(n2181), .ZN(n2381) );
  NAND2_X1 U2539 ( .A1(n3396), .A2(n3397), .ZN(n2398) );
  NAND2_X1 U2540 ( .A1(n2401), .A2(n2400), .ZN(n2399) );
  INV_X1 U2541 ( .A(n3397), .ZN(n2400) );
  INV_X1 U2542 ( .A(n3396), .ZN(n2401) );
  AOI21_X1 U2543 ( .B1(n3009), .B2(n3119), .A(n2640), .ZN(n2644) );
  OR2_X1 U2544 ( .A1(n3062), .A2(n3416), .ZN(n3092) );
  INV_X1 U2545 ( .A(n4946), .ZN(n3073) );
  AND2_X1 U2546 ( .A1(n4828), .A2(n4829), .ZN(n3209) );
  OR2_X1 U2547 ( .A1(n3092), .A2(n3242), .ZN(n3082) );
  OAI21_X1 U2548 ( .B1(n4427), .B2(n2293), .A(n2292), .ZN(n2291) );
  AOI21_X1 U2549 ( .B1(n4487), .B2(n4430), .A(n4292), .ZN(n2292) );
  NAND2_X1 U2550 ( .A1(n2295), .A2(n2294), .ZN(n2293) );
  NAND2_X1 U2551 ( .A1(n4431), .A2(n4292), .ZN(n2290) );
  NAND2_X1 U2552 ( .A1(n4513), .A2(n3027), .ZN(n2301) );
  AND4_X1 U2553 ( .A1(n2813), .A2(n2812), .A3(n2811), .A4(n2810), .ZN(n3400)
         );
  NAND2_X1 U2554 ( .A1(n2559), .A2(n2558), .ZN(n2560) );
  OR2_X1 U2555 ( .A1(n2163), .A2(n4845), .ZN(n2341) );
  NAND2_X1 U2556 ( .A1(n2452), .A2(n2451), .ZN(n2458) );
  NAND2_X1 U2557 ( .A1(n4845), .A2(REG2_REG_4__SCAN_IN), .ZN(n2343) );
  INV_X1 U2558 ( .A(n2458), .ZN(n2339) );
  NOR2_X1 U2559 ( .A1(n2464), .A2(n3268), .ZN(n2465) );
  OR2_X1 U2560 ( .A1(n2565), .A2(n2411), .ZN(n2347) );
  NAND2_X1 U2561 ( .A1(n2563), .A2(n2348), .ZN(n2345) );
  INV_X1 U2562 ( .A(n3289), .ZN(n2194) );
  NOR2_X1 U2563 ( .A1(n2192), .A2(n3613), .ZN(n2191) );
  INV_X1 U2564 ( .A(n2195), .ZN(n2192) );
  OR2_X1 U2565 ( .A1(n3289), .A2(n2196), .ZN(n2193) );
  NAND2_X1 U2566 ( .A1(n2143), .A2(n2566), .ZN(n2196) );
  NAND2_X1 U2567 ( .A1(n3289), .A2(n4832), .ZN(n2190) );
  INV_X1 U2568 ( .A(n4983), .ZN(n2776) );
  NAND2_X1 U2569 ( .A1(n2363), .A2(REG1_REG_12__SCAN_IN), .ZN(n2364) );
  INV_X1 U2570 ( .A(n4863), .ZN(n2363) );
  NOR2_X1 U2571 ( .A1(n2579), .A2(n4978), .ZN(n4900) );
  OAI21_X1 U2572 ( .B1(n4474), .B2(REG2_REG_16__SCAN_IN), .A(n2496), .ZN(n4918) );
  NAND2_X1 U2573 ( .A1(n2202), .A2(n2200), .ZN(n4917) );
  AOI21_X1 U2574 ( .B1(n2496), .B2(REG2_REG_16__SCAN_IN), .A(n2201), .ZN(n2200) );
  NAND2_X1 U2575 ( .A1(n4474), .A2(n2496), .ZN(n2202) );
  NAND2_X1 U2576 ( .A1(n4918), .A2(n2354), .ZN(n2353) );
  NOR2_X1 U2577 ( .A1(n2201), .A2(n2183), .ZN(n2354) );
  OAI21_X1 U2578 ( .B1(n4578), .B2(n2234), .A(n2230), .ZN(n4503) );
  AOI21_X1 U2579 ( .B1(n2233), .B2(n2232), .A(n2231), .ZN(n2230) );
  INV_X1 U2580 ( .A(n4346), .ZN(n2231) );
  INV_X1 U2581 ( .A(n2239), .ZN(n2232) );
  INV_X1 U2582 ( .A(n4505), .ZN(n4538) );
  AND2_X1 U2583 ( .A1(n2243), .A2(n2241), .ZN(n4543) );
  AND2_X1 U2584 ( .A1(n2996), .A2(n2987), .ZN(n4571) );
  INV_X1 U2585 ( .A(n2222), .ZN(n2221) );
  OAI21_X1 U2586 ( .B1(n2139), .B2(n4620), .A(n2146), .ZN(n2222) );
  NAND2_X1 U2587 ( .A1(n2941), .A2(n2299), .ZN(n2968) );
  NAND2_X1 U2588 ( .A1(n3157), .A2(n2179), .ZN(n2305) );
  NAND2_X1 U2589 ( .A1(n2887), .A2(n2155), .ZN(n2943) );
  NAND2_X1 U2590 ( .A1(n4616), .A2(n4620), .ZN(n4615) );
  OAI21_X1 U2591 ( .B1(n3760), .B2(n3151), .A(n2205), .ZN(n2204) );
  INV_X1 U2592 ( .A(n3152), .ZN(n2205) );
  NAND2_X1 U2593 ( .A1(n2887), .A2(n2151), .ZN(n2928) );
  NAND2_X1 U2594 ( .A1(n3149), .A2(n3148), .ZN(n3789) );
  AND2_X1 U2595 ( .A1(n2424), .A2(n2309), .ZN(n2308) );
  NAND2_X1 U2596 ( .A1(n2283), .A2(n2156), .ZN(n2808) );
  OR2_X1 U2597 ( .A1(n2209), .A2(n2208), .ZN(n2207) );
  INV_X1 U2598 ( .A(n4379), .ZN(n2208) );
  NAND2_X1 U2599 ( .A1(n3406), .A2(n4372), .ZN(n3123) );
  NAND2_X1 U2600 ( .A1(n4947), .A2(n3379), .ZN(n4709) );
  NAND2_X1 U2601 ( .A1(n3116), .A2(n3115), .ZN(n3164) );
  CLKBUF_X1 U2602 ( .A(n3063), .Z(n3080) );
  NAND2_X1 U2603 ( .A1(n2269), .A2(n2138), .ZN(n2267) );
  NOR2_X1 U2604 ( .A1(n2142), .A2(n4535), .ZN(n3215) );
  NOR2_X1 U2605 ( .A1(n3049), .A2(n3048), .ZN(n3243) );
  INV_X1 U2606 ( .A(n3244), .ZN(n3048) );
  NAND2_X1 U2607 ( .A1(n2456), .A2(n2453), .ZN(n2229) );
  AND2_X1 U2608 ( .A1(n2501), .A2(n2600), .ZN(n2506) );
  NOR2_X1 U2609 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2501)
         );
  INV_X1 U2610 ( .A(n2531), .ZN(n2329) );
  INV_X1 U2611 ( .A(IR_REG_19__SCAN_IN), .ZN(n2605) );
  XNOR2_X1 U2612 ( .A(n2438), .B(IR_REG_13__SCAN_IN), .ZN(n2828) );
  INV_X1 U2613 ( .A(IR_REG_12__SCAN_IN), .ZN(n2481) );
  NOR2_X1 U2614 ( .A1(n2471), .A2(IR_REG_9__SCAN_IN), .ZN(n2473) );
  INV_X1 U2615 ( .A(IR_REG_10__SCAN_IN), .ZN(n2474) );
  OR3_X1 U2616 ( .A1(n2466), .A2(IR_REG_7__SCAN_IN), .A3(IR_REG_8__SCAN_IN), 
        .ZN(n2471) );
  NAND2_X1 U2617 ( .A1(n2377), .A2(n2374), .ZN(n2373) );
  NAND2_X1 U2618 ( .A1(n2174), .A2(n3551), .ZN(n2393) );
  NOR2_X1 U2619 ( .A1(n2174), .A2(n3551), .ZN(n2394) );
  NAND2_X1 U2620 ( .A1(n2383), .A2(n2388), .ZN(n3895) );
  NAND2_X1 U2621 ( .A1(n3731), .A2(n2390), .ZN(n2383) );
  INV_X1 U2622 ( .A(n4239), .ZN(n4657) );
  INV_X1 U2623 ( .A(n4552), .ZN(n4547) );
  INV_X1 U2624 ( .A(n4550), .ZN(n4442) );
  NAND2_X1 U2625 ( .A1(n3002), .A2(n3001), .ZN(n4566) );
  OR2_X1 U2626 ( .A1(n4553), .A2(n2767), .ZN(n3002) );
  OR2_X1 U2627 ( .A1(n4627), .A2(n2767), .ZN(n2949) );
  AND2_X1 U2628 ( .A1(n2546), .A2(n2544), .ZN(n3254) );
  NAND2_X1 U2629 ( .A1(n2352), .A2(n2351), .ZN(n2350) );
  NAND2_X1 U2630 ( .A1(n3265), .A2(REG1_REG_6__SCAN_IN), .ZN(n2352) );
  AND2_X1 U2631 ( .A1(n3254), .A2(n4838), .ZN(n4908) );
  NAND2_X1 U2632 ( .A1(n2371), .A2(n4473), .ZN(n2370) );
  OAI21_X1 U2633 ( .B1(n2159), .B2(n4646), .A(n4515), .ZN(n4516) );
  INV_X1 U2634 ( .A(n2269), .ZN(n2266) );
  INV_X1 U2635 ( .A(n2322), .ZN(n2318) );
  INV_X1 U2636 ( .A(n4719), .ZN(n4722) );
  NOR2_X1 U2637 ( .A1(n4499), .A2(n4506), .ZN(n4498) );
  INV_X1 U2638 ( .A(n2267), .ZN(n2265) );
  AOI21_X1 U2639 ( .B1(n4718), .B2(n2153), .A(n2176), .ZN(n2215) );
  AND2_X1 U2640 ( .A1(n2312), .A2(n2166), .ZN(n2310) );
  INV_X1 U2641 ( .A(n4305), .ZN(n2254) );
  INV_X1 U2642 ( .A(IR_REG_26__SCAN_IN), .ZN(n2527) );
  INV_X1 U2643 ( .A(IR_REG_27__SCAN_IN), .ZN(n2534) );
  INV_X1 U2644 ( .A(n2729), .ZN(n2284) );
  INV_X1 U2645 ( .A(n2909), .ZN(n2912) );
  INV_X1 U2646 ( .A(n2910), .ZN(n2911) );
  NAND2_X1 U2647 ( .A1(n4428), .A2(n4429), .ZN(n2295) );
  INV_X1 U2648 ( .A(n4426), .ZN(n2294) );
  INV_X1 U2649 ( .A(n2411), .ZN(n2348) );
  NAND2_X1 U2650 ( .A1(n4894), .A2(n2491), .ZN(n2495) );
  INV_X1 U2651 ( .A(n2238), .ZN(n2237) );
  OAI21_X1 U2652 ( .B1(n2241), .B2(n4421), .A(n4288), .ZN(n2238) );
  NOR2_X1 U2653 ( .A1(n2240), .A2(n4421), .ZN(n2239) );
  INV_X1 U2654 ( .A(n4413), .ZN(n2240) );
  NAND2_X1 U2655 ( .A1(n2221), .A2(n2219), .ZN(n2218) );
  AND2_X1 U2656 ( .A1(n2139), .A2(n2177), .ZN(n2219) );
  NOR2_X1 U2657 ( .A1(n4360), .A2(n2242), .ZN(n2241) );
  NAND2_X1 U2658 ( .A1(n2304), .A2(n3159), .ZN(n2303) );
  INV_X1 U2659 ( .A(n2305), .ZN(n2304) );
  NOR2_X1 U2660 ( .A1(n4092), .A2(n2297), .ZN(n2296) );
  INV_X1 U2661 ( .A(n2888), .ZN(n2887) );
  NAND2_X1 U2662 ( .A1(n2310), .A2(n2314), .ZN(n2309) );
  INV_X1 U2663 ( .A(n4929), .ZN(n4933) );
  INV_X1 U2664 ( .A(DATAI_21_), .ZN(n4036) );
  OR2_X1 U2665 ( .A1(n3659), .A2(n2314), .ZN(n2311) );
  INV_X1 U2666 ( .A(n3535), .ZN(n3176) );
  NAND2_X1 U2667 ( .A1(n2723), .A2(n3485), .ZN(n2272) );
  AND2_X1 U2668 ( .A1(n3568), .A2(n3413), .ZN(n3412) );
  INV_X1 U2669 ( .A(n3606), .ZN(n3167) );
  OAI211_X1 U2670 ( .C1(n3563), .C2(n2252), .A(n4317), .B(n2250), .ZN(n3510)
         );
  INV_X1 U2671 ( .A(n2253), .ZN(n2252) );
  NAND2_X1 U2672 ( .A1(n2251), .A2(n2253), .ZN(n2250) );
  NOR2_X1 U2673 ( .A1(n3599), .A2(n2254), .ZN(n2253) );
  AOI21_X1 U2674 ( .B1(n2526), .B2(n2527), .A(n2525), .ZN(n2538) );
  NAND2_X1 U2675 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2525) );
  INV_X1 U2676 ( .A(IR_REG_20__SCAN_IN), .ZN(n2621) );
  NAND3_X1 U2677 ( .A1(n2504), .A2(n2503), .A3(n2502), .ZN(n2601) );
  INV_X1 U2678 ( .A(IR_REG_17__SCAN_IN), .ZN(n2503) );
  INV_X1 U2679 ( .A(IR_REG_16__SCAN_IN), .ZN(n2502) );
  NAND2_X1 U2680 ( .A1(n2377), .A2(n2378), .ZN(n3927) );
  NAND2_X1 U2681 ( .A1(n2284), .A2(REG3_REG_7__SCAN_IN), .ZN(n2741) );
  AND2_X1 U2682 ( .A1(n3896), .A2(n2385), .ZN(n2384) );
  NAND2_X1 U2683 ( .A1(n2388), .A2(n2386), .ZN(n2385) );
  INV_X1 U2684 ( .A(n2390), .ZN(n2386) );
  INV_X1 U2685 ( .A(n2388), .ZN(n2387) );
  NOR2_X1 U2686 ( .A1(n4256), .A2(n2391), .ZN(n2390) );
  INV_X1 U2687 ( .A(n3732), .ZN(n2391) );
  AOI21_X1 U2688 ( .B1(n2389), .B2(n2392), .A(n2186), .ZN(n2388) );
  INV_X1 U2689 ( .A(n4256), .ZN(n2389) );
  INV_X1 U2690 ( .A(n2185), .ZN(n2392) );
  INV_X1 U2691 ( .A(n2697), .ZN(n2380) );
  AND2_X1 U2692 ( .A1(n3449), .A2(n3447), .ZN(n2693) );
  NAND2_X1 U2693 ( .A1(n2984), .A2(n2983), .ZN(n2985) );
  AND2_X1 U2694 ( .A1(n3209), .A2(n3076), .ZN(n3106) );
  INV_X1 U2695 ( .A(n4277), .ZN(n4260) );
  AND2_X1 U2696 ( .A1(n2882), .A2(n2881), .ZN(n3747) );
  OR2_X1 U2697 ( .A1(n2551), .A2(REG2_REG_1__SCAN_IN), .ZN(n2440) );
  NAND2_X1 U2698 ( .A1(n2555), .A2(n2554), .ZN(n3332) );
  OR2_X1 U2699 ( .A1(n2143), .A2(n2566), .ZN(n2195) );
  NAND2_X1 U2700 ( .A1(n4460), .A2(n2412), .ZN(n2476) );
  OAI211_X1 U2701 ( .C1(n2569), .C2(n2358), .A(n2356), .B(n2147), .ZN(n2570)
         );
  NOR2_X1 U2702 ( .A1(n2358), .A2(n2743), .ZN(n2357) );
  OR2_X1 U2703 ( .A1(n4898), .A2(n4897), .ZN(n4894) );
  NAND2_X1 U2704 ( .A1(n2581), .A2(n2580), .ZN(n2584) );
  NOR2_X1 U2705 ( .A1(n4513), .A2(n4691), .ZN(n4514) );
  INV_X1 U2706 ( .A(n2301), .ZN(n4521) );
  NOR2_X1 U2707 ( .A1(n3161), .A2(n2325), .ZN(n2320) );
  NAND2_X1 U2708 ( .A1(n2152), .A2(n4356), .ZN(n2325) );
  NAND2_X1 U2709 ( .A1(n2236), .A2(n2237), .ZN(n4533) );
  NAND2_X1 U2710 ( .A1(n4578), .A2(n2239), .ZN(n2236) );
  INV_X1 U2711 ( .A(n4345), .ZN(n4535) );
  AND2_X1 U2712 ( .A1(n3023), .A2(n3022), .ZN(n4550) );
  OR2_X1 U2713 ( .A1(n4530), .A2(n2767), .ZN(n3023) );
  AND2_X1 U2714 ( .A1(n2974), .A2(n2973), .ZN(n4564) );
  AND2_X1 U2715 ( .A1(n2243), .A2(n2244), .ZN(n4562) );
  AND2_X1 U2716 ( .A1(n2299), .A2(REG3_REG_24__SCAN_IN), .ZN(n2298) );
  AND2_X1 U2717 ( .A1(n2960), .A2(n2959), .ZN(n4581) );
  NAND2_X1 U2718 ( .A1(n2941), .A2(REG3_REG_22__SCAN_IN), .ZN(n2954) );
  NAND2_X1 U2719 ( .A1(n3195), .A2(n2247), .ZN(n4653) );
  AND2_X1 U2720 ( .A1(n2894), .A2(n2893), .ZN(n3900) );
  AND2_X1 U2721 ( .A1(n2906), .A2(n2905), .ZN(n4262) );
  AND2_X1 U2722 ( .A1(n2861), .A2(n2860), .ZN(n3817) );
  NAND2_X1 U2723 ( .A1(n2287), .A2(n2285), .ZN(n2876) );
  NOR2_X1 U2724 ( .A1(n2154), .A2(n2286), .ZN(n2285) );
  INV_X1 U2725 ( .A(n4215), .ZN(n3750) );
  NAND2_X1 U2726 ( .A1(n2287), .A2(n2141), .ZN(n2846) );
  NAND2_X1 U2727 ( .A1(n2287), .A2(REG3_REG_13__SCAN_IN), .ZN(n2834) );
  NOR2_X1 U2728 ( .A1(n2410), .A2(n3187), .ZN(n3188) );
  INV_X1 U2729 ( .A(n3190), .ZN(n4367) );
  INV_X1 U2730 ( .A(n2808), .ZN(n2807) );
  INV_X1 U2731 ( .A(n2158), .ZN(n2211) );
  OR2_X1 U2732 ( .A1(n2765), .A2(n2764), .ZN(n2777) );
  NAND2_X1 U2733 ( .A1(n2283), .A2(REG3_REG_10__SCAN_IN), .ZN(n2797) );
  INV_X1 U2734 ( .A(n3634), .ZN(n3626) );
  AND2_X1 U2735 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2699) );
  NAND2_X1 U2736 ( .A1(n2699), .A2(REG3_REG_5__SCAN_IN), .ZN(n2716) );
  NAND2_X1 U2737 ( .A1(n3563), .A2(n2255), .ZN(n2249) );
  INV_X1 U2738 ( .A(n2251), .ZN(n2255) );
  INV_X1 U2739 ( .A(n3516), .ZN(n3100) );
  NAND2_X1 U2740 ( .A1(n3563), .A2(n4301), .ZN(n3407) );
  INV_X1 U2741 ( .A(n4935), .ZN(n4618) );
  NOR2_X1 U2742 ( .A1(n3567), .A2(n4300), .ZN(n3568) );
  AND2_X1 U2743 ( .A1(n4927), .A2(n3118), .ZN(n4701) );
  OR2_X1 U2744 ( .A1(n3033), .A2(n2672), .ZN(n2676) );
  AND2_X1 U2745 ( .A1(n3208), .A2(n3207), .ZN(n4704) );
  INV_X1 U2746 ( .A(n4709), .ZN(n3099) );
  AND2_X1 U2747 ( .A1(n3209), .A2(n3340), .ZN(n4935) );
  NOR2_X1 U2748 ( .A1(n4998), .A2(n4829), .ZN(n3108) );
  AOI21_X1 U2749 ( .B1(n3243), .B2(n3247), .A(n3050), .ZN(n3417) );
  OR2_X1 U2750 ( .A1(n2137), .A2(n2646), .ZN(n2648) );
  NAND2_X1 U2751 ( .A1(n3209), .A2(n4838), .ZN(n4952) );
  INV_X1 U2752 ( .A(DATAI_0_), .ZN(n2259) );
  INV_X1 U2753 ( .A(n4354), .ZN(n4506) );
  INV_X1 U2754 ( .A(n4682), .ZN(n4937) );
  OR2_X1 U2755 ( .A1(n2134), .A2(n3036), .ZN(n3216) );
  OR2_X1 U2756 ( .A1(n2134), .A2(n3003), .ZN(n4552) );
  OR2_X1 U2757 ( .A1(n2134), .A2(n2993), .ZN(n4570) );
  OR2_X1 U2758 ( .A1(n2134), .A2(n4036), .ZN(n4643) );
  OR2_X1 U2759 ( .A1(n2281), .A2(n4667), .ZN(n2279) );
  NOR2_X1 U2760 ( .A1(n4771), .A2(n3821), .ZN(n3765) );
  NOR2_X1 U2761 ( .A1(n2144), .A2(n3688), .ZN(n2274) );
  NAND2_X1 U2762 ( .A1(n2273), .A2(n2275), .ZN(n3668) );
  NOR2_X1 U2763 ( .A1(n4690), .A2(n2144), .ZN(n3701) );
  INV_X1 U2764 ( .A(n2138), .ZN(n4779) );
  NOR2_X1 U2765 ( .A1(n3516), .A2(n2270), .ZN(n3632) );
  NAND2_X1 U2766 ( .A1(n2271), .A2(n3176), .ZN(n2270) );
  INV_X1 U2767 ( .A(n2272), .ZN(n2271) );
  NOR2_X1 U2768 ( .A1(n3516), .A2(n2272), .ZN(n3533) );
  NAND2_X1 U2769 ( .A1(n3100), .A2(n2723), .ZN(n3519) );
  OR2_X1 U2770 ( .A1(n4953), .A2(n4828), .ZN(n4998) );
  NAND2_X1 U2771 ( .A1(n2328), .A2(IR_REG_31__SCAN_IN), .ZN(n2256) );
  NOR2_X1 U2772 ( .A1(n2531), .A2(n2532), .ZN(n2333) );
  OR3_X1 U2773 ( .A1(n2488), .A2(IR_REG_16__SCAN_IN), .A3(IR_REG_15__SCAN_IN), 
        .ZN(n2497) );
  INV_X1 U2774 ( .A(IR_REG_11__SCAN_IN), .ZN(n2478) );
  INV_X1 U2775 ( .A(IR_REG_7__SCAN_IN), .ZN(n2467) );
  NAND2_X1 U2776 ( .A1(n2449), .A2(IR_REG_31__SCAN_IN), .ZN(n2454) );
  NAND2_X1 U2777 ( .A1(n2402), .A2(n2403), .ZN(n4221) );
  AND2_X1 U2778 ( .A1(n2407), .A2(n2404), .ZN(n2403) );
  NAND2_X1 U2779 ( .A1(n2405), .A2(n2418), .ZN(n2404) );
  INV_X1 U2780 ( .A(n3844), .ZN(n3902) );
  NAND2_X1 U2781 ( .A1(n3359), .A2(n2413), .ZN(n3357) );
  NAND2_X1 U2782 ( .A1(n4233), .A2(n4237), .ZN(n3909) );
  INV_X1 U2783 ( .A(n4283), .ZN(n3923) );
  INV_X1 U2784 ( .A(n2866), .ZN(n2875) );
  NAND2_X1 U2785 ( .A1(n3441), .A2(n2693), .ZN(n3448) );
  OR2_X1 U2786 ( .A1(n3092), .A2(n3090), .ZN(n4280) );
  INV_X1 U2787 ( .A(n4947), .ZN(n4942) );
  INV_X1 U2788 ( .A(n4280), .ZN(n4249) );
  NOR2_X1 U2789 ( .A1(n3500), .A2(n2396), .ZN(n2395) );
  INV_X1 U2790 ( .A(n2398), .ZN(n2396) );
  INV_X1 U2791 ( .A(n4285), .ZN(n4247) );
  INV_X1 U2792 ( .A(n3923), .ZN(n4252) );
  AND2_X1 U2793 ( .A1(n2992), .A2(n2991), .ZN(n4278) );
  INV_X1 U2794 ( .A(n3082), .ZN(n3065) );
  OAI21_X1 U2795 ( .B1(n3082), .B2(n4682), .A(n4691), .ZN(n4283) );
  INV_X1 U2796 ( .A(n2288), .ZN(n4434) );
  AOI21_X1 U2797 ( .B1(n4432), .B2(n3080), .A(n2289), .ZN(n2288) );
  AOI21_X1 U2798 ( .B1(n2291), .B2(n2290), .A(n3080), .ZN(n2289) );
  OAI21_X1 U2799 ( .B1(n2301), .B2(n2767), .A(n3035), .ZN(n4505) );
  INV_X1 U2800 ( .A(n4278), .ZN(n4583) );
  INV_X1 U2801 ( .A(n4564), .ZN(n4603) );
  INV_X1 U2802 ( .A(n4581), .ZN(n4624) );
  NAND2_X1 U2803 ( .A1(n2934), .A2(n2933), .ZN(n4239) );
  NAND2_X1 U2804 ( .A1(n2919), .A2(n2918), .ZN(n4636) );
  OR2_X1 U2805 ( .A1(n4668), .A2(n2767), .ZN(n2919) );
  INV_X1 U2806 ( .A(n4262), .ZN(n4655) );
  INV_X1 U2807 ( .A(n3900), .ZN(n3792) );
  INV_X1 U2808 ( .A(n3747), .ZN(n4259) );
  INV_X1 U2809 ( .A(n3817), .ZN(n3724) );
  INV_X1 U2810 ( .A(n3400), .ZN(n3695) );
  INV_X1 U2811 ( .A(n3121), .ZN(n4446) );
  OR2_X1 U2812 ( .A1(n2767), .A2(n2630), .ZN(n2634) );
  OR2_X1 U2813 ( .A1(n2137), .A2(n5021), .ZN(n2658) );
  OR2_X1 U2814 ( .A1(n2767), .A2(n2655), .ZN(n2659) );
  OAI21_X1 U2815 ( .B1(n2551), .B2(REG1_REG_1__SCAN_IN), .A(n2552), .ZN(n4452)
         );
  INV_X1 U2816 ( .A(n2343), .ZN(n2338) );
  XNOR2_X1 U2817 ( .A(n2567), .B(n2566), .ZN(n3301) );
  NAND2_X1 U2818 ( .A1(n3301), .A2(REG1_REG_8__SCAN_IN), .ZN(n3300) );
  NAND2_X1 U2819 ( .A1(n2198), .A2(n2197), .ZN(n4462) );
  NAND2_X1 U2820 ( .A1(n2194), .A2(n2143), .ZN(n2199) );
  NAND2_X1 U2821 ( .A1(n4462), .A2(n4461), .ZN(n4460) );
  XNOR2_X1 U2822 ( .A(n2570), .B(n2776), .ZN(n4854) );
  NAND2_X1 U2823 ( .A1(n4859), .A2(REG2_REG_10__SCAN_IN), .ZN(n4858) );
  AND2_X1 U2824 ( .A1(n2335), .A2(n2334), .ZN(n3537) );
  INV_X1 U2825 ( .A(n3538), .ZN(n2334) );
  INV_X1 U2826 ( .A(n2335), .ZN(n3539) );
  NAND2_X1 U2827 ( .A1(n2367), .A2(n2366), .ZN(n3540) );
  AND2_X1 U2828 ( .A1(n2364), .A2(n2575), .ZN(n4873) );
  NAND2_X1 U2829 ( .A1(n4867), .A2(n2485), .ZN(n4879) );
  XNOR2_X1 U2830 ( .A(n2486), .B(n4978), .ZN(n4886) );
  INV_X1 U2831 ( .A(n4908), .ZN(n4926) );
  NOR2_X1 U2832 ( .A1(n2611), .A2(n2355), .ZN(n2543) );
  NAND2_X1 U2833 ( .A1(n2353), .A2(n2187), .ZN(n2355) );
  AND2_X1 U2834 ( .A1(n2592), .A2(n2591), .ZN(n2599) );
  AND2_X1 U2835 ( .A1(n3254), .A2(n4435), .ZN(n4921) );
  NOR2_X1 U2836 ( .A1(n2321), .A2(n4358), .ZN(n4528) );
  OAI21_X1 U2837 ( .B1(n4616), .B2(n2139), .A(n2221), .ZN(n4559) );
  NAND2_X1 U2838 ( .A1(n2306), .A2(n2305), .ZN(n4576) );
  NAND2_X1 U2839 ( .A1(n4615), .A2(n2140), .ZN(n2306) );
  NAND2_X1 U2840 ( .A1(n4615), .A2(n3156), .ZN(n4594) );
  OR2_X1 U2841 ( .A1(n4625), .A2(n3155), .ZN(n4744) );
  OR2_X1 U2842 ( .A1(n3682), .A2(n3870), .ZN(n4771) );
  OR2_X1 U2843 ( .A1(n3659), .A2(n3143), .ZN(n2315) );
  NAND2_X1 U2844 ( .A1(n2214), .A2(n2158), .ZN(n2213) );
  INV_X1 U2845 ( .A(n4954), .ZN(n4691) );
  NAND2_X1 U2846 ( .A1(n3099), .A2(n3390), .ZN(n3567) );
  INV_X1 U2847 ( .A(n4646), .ZN(n4943) );
  AND2_X1 U2848 ( .A1(n4958), .A2(n3423), .ZN(n4955) );
  NAND2_X1 U2849 ( .A1(n4485), .A2(n4484), .ZN(n4793) );
  OR2_X1 U2850 ( .A1(n2267), .A2(n4498), .ZN(n2260) );
  OR2_X1 U2851 ( .A1(n3243), .A2(n3242), .ZN(n4974) );
  NOR2_X1 U2852 ( .A1(n2510), .A2(n2327), .ZN(n2330) );
  NOR2_X1 U2853 ( .A1(n2532), .A2(n2511), .ZN(n2326) );
  NAND2_X1 U2854 ( .A1(n2537), .A2(n2626), .ZN(n2327) );
  NAND2_X1 U2855 ( .A1(n2518), .A2(IR_REG_31__SCAN_IN), .ZN(n2508) );
  AND2_X1 U2856 ( .A1(n3078), .A2(STATE_REG_SCAN_IN), .ZN(n4975) );
  OR2_X1 U2857 ( .A1(n2606), .A2(n2605), .ZN(n2607) );
  INV_X1 U2858 ( .A(n2588), .ZN(n4976) );
  XNOR2_X1 U2859 ( .A(n2492), .B(IR_REG_15__SCAN_IN), .ZN(n4907) );
  INV_X1 U2860 ( .A(n2828), .ZN(n4980) );
  XNOR2_X1 U2861 ( .A(n2479), .B(n2478), .ZN(n3546) );
  XNOR2_X1 U2862 ( .A(n2475), .B(n2474), .ZN(n4983) );
  XNOR2_X1 U2863 ( .A(n2472), .B(IR_REG_9__SCAN_IN), .ZN(n4831) );
  AND2_X1 U2864 ( .A1(n2461), .A2(n2460), .ZN(n4834) );
  INV_X1 U2865 ( .A(n3286), .ZN(n2349) );
  NAND2_X1 U2866 ( .A1(n4516), .A2(n4958), .ZN(n4518) );
  NOR2_X1 U2867 ( .A1(n2414), .A2(n2415), .ZN(n3114) );
  INV_X1 U2868 ( .A(n2262), .ZN(n2261) );
  INV_X1 U2869 ( .A(n4498), .ZN(n2264) );
  OAI21_X1 U2870 ( .B1(n3225), .B2(n3224), .A(n2421), .ZN(U3546) );
  OR2_X1 U2871 ( .A1(n4523), .A2(n4761), .ZN(n3223) );
  NAND2_X1 U2872 ( .A1(n2227), .A2(n2226), .ZN(U3515) );
  NAND2_X1 U2873 ( .A1(n5019), .A2(REG0_REG_29__SCAN_IN), .ZN(n2226) );
  NAND2_X1 U2874 ( .A1(n2228), .A2(n5020), .ZN(n2227) );
  NAND2_X1 U2875 ( .A1(n2145), .A2(n2164), .ZN(n2228) );
  AND2_X1 U2876 ( .A1(n3219), .A2(n3218), .ZN(n3220) );
  NAND2_X1 U2877 ( .A1(n3159), .A2(n2140), .ZN(n2139) );
  AND2_X1 U2878 ( .A1(n3157), .A2(n3156), .ZN(n2140) );
  AND2_X1 U2879 ( .A1(REG3_REG_13__SCAN_IN), .A2(REG3_REG_14__SCAN_IN), .ZN(
        n2141) );
  OR3_X1 U2880 ( .A1(n4744), .A2(n2277), .A3(n4547), .ZN(n2142) );
  OR2_X1 U2881 ( .A1(n3285), .A2(n3492), .ZN(n2143) );
  XNOR2_X1 U2882 ( .A(n2457), .B(n2456), .ZN(n3227) );
  INV_X1 U2883 ( .A(n3227), .ZN(n4845) );
  NAND2_X1 U2884 ( .A1(n2275), .A2(n3182), .ZN(n2144) );
  AND2_X1 U2885 ( .A1(n2422), .A2(n2215), .ZN(n2145) );
  INV_X1 U2886 ( .A(n2276), .ZN(n4551) );
  NAND2_X1 U2887 ( .A1(n4624), .A2(n4606), .ZN(n3157) );
  NAND2_X1 U2888 ( .A1(n2807), .A2(REG3_REG_12__SCAN_IN), .ZN(n2822) );
  INV_X1 U2889 ( .A(n2822), .ZN(n2287) );
  AND2_X1 U2890 ( .A1(n2303), .A2(n2178), .ZN(n2146) );
  OR2_X1 U2891 ( .A1(n4464), .A2(n2768), .ZN(n2147) );
  AND2_X1 U2892 ( .A1(n2406), .A2(n2173), .ZN(n2148) );
  OR2_X1 U2893 ( .A1(n4690), .A2(n4689), .ZN(n2149) );
  INV_X1 U2894 ( .A(n4360), .ZN(n2244) );
  OR2_X1 U2895 ( .A1(n4771), .A2(n2281), .ZN(n2150) );
  AND2_X1 U2896 ( .A1(n2296), .A2(REG3_REG_20__SCAN_IN), .ZN(n2151) );
  NAND2_X1 U2897 ( .A1(n4442), .A2(n4535), .ZN(n2152) );
  AND2_X1 U2898 ( .A1(n4716), .A2(n5017), .ZN(n2153) );
  NAND2_X1 U2899 ( .A1(n2141), .A2(REG3_REG_15__SCAN_IN), .ZN(n2154) );
  INV_X1 U2900 ( .A(n2280), .ZN(n3766) );
  AND2_X1 U2901 ( .A1(n2151), .A2(REG3_REG_21__SCAN_IN), .ZN(n2155) );
  AND2_X1 U2902 ( .A1(REG3_REG_11__SCAN_IN), .A2(REG3_REG_10__SCAN_IN), .ZN(
        n2156) );
  INV_X1 U2903 ( .A(REG3_REG_14__SCAN_IN), .ZN(n2833) );
  OR2_X1 U2904 ( .A1(n2134), .A2(n2975), .ZN(n4589) );
  INV_X1 U2905 ( .A(n4958), .ZN(n4698) );
  NAND2_X2 U2906 ( .A1(n2637), .A2(n3226), .ZN(n2681) );
  INV_X1 U2907 ( .A(n3116), .ZN(n3117) );
  NAND2_X1 U2908 ( .A1(n3195), .A2(n4404), .ZN(n3756) );
  NAND2_X1 U2909 ( .A1(n2311), .A2(n2312), .ZN(n3678) );
  OR2_X1 U2910 ( .A1(n2822), .A2(n2154), .ZN(n2157) );
  NOR2_X1 U2911 ( .A1(n3479), .A2(n3139), .ZN(n2158) );
  OR2_X1 U2912 ( .A1(n3511), .A2(n3485), .ZN(n3170) );
  OR2_X1 U2913 ( .A1(n4498), .A2(n2266), .ZN(n2159) );
  OR2_X1 U2914 ( .A1(n4446), .A2(n4300), .ZN(n2160) );
  NAND2_X1 U2915 ( .A1(n2887), .A2(n2296), .ZN(n2161) );
  NAND2_X1 U2916 ( .A1(n2204), .A2(n4365), .ZN(n4632) );
  AOI21_X1 U2917 ( .B1(n3731), .B2(n3732), .A(n2392), .ZN(n4255) );
  NAND2_X1 U2918 ( .A1(n2315), .A2(n3142), .ZN(n3687) );
  AOI21_X1 U2919 ( .B1(n4616), .B2(n2220), .A(n2217), .ZN(n2216) );
  AND2_X1 U2920 ( .A1(n3688), .A2(n4444), .ZN(n2162) );
  AND2_X1 U2921 ( .A1(n3227), .A2(REG2_REG_4__SCAN_IN), .ZN(n2163) );
  NAND2_X1 U2922 ( .A1(n2373), .A2(n2375), .ZN(n2551) );
  AND2_X1 U2923 ( .A1(n4722), .A2(n2260), .ZN(n2164) );
  INV_X1 U2924 ( .A(n2234), .ZN(n2233) );
  NAND2_X1 U2925 ( .A1(n2237), .A2(n2235), .ZN(n2234) );
  MUX2_X1 U2926 ( .A(DATAI_3_), .B(n4835), .S(n2134), .Z(n4300) );
  NOR2_X1 U2927 ( .A1(n4689), .A2(n3577), .ZN(n2165) );
  INV_X1 U2928 ( .A(n4468), .ZN(n2358) );
  AND2_X1 U2929 ( .A1(n3742), .A2(n3190), .ZN(n2166) );
  AND2_X1 U2930 ( .A1(n4307), .A2(n3170), .ZN(n2167) );
  NAND2_X1 U2931 ( .A1(n2506), .A2(n2505), .ZN(n2511) );
  NOR2_X1 U2932 ( .A1(n2411), .A2(n2718), .ZN(n2168) );
  NAND2_X1 U2933 ( .A1(n4636), .A2(n3200), .ZN(n2169) );
  NAND2_X1 U2934 ( .A1(n4689), .A2(n3577), .ZN(n2170) );
  OR2_X1 U2935 ( .A1(n3281), .A2(n2462), .ZN(n2171) );
  INV_X1 U2936 ( .A(IR_REG_5__SCAN_IN), .ZN(n2528) );
  AND2_X1 U2937 ( .A1(REG3_REG_7__SCAN_IN), .A2(REG3_REG_8__SCAN_IN), .ZN(
        n2172) );
  INV_X1 U2938 ( .A(IR_REG_31__SCAN_IN), .ZN(n2535) );
  NAND2_X1 U2939 ( .A1(n3166), .A2(n4390), .ZN(n3563) );
  NOR2_X1 U2940 ( .A1(n4771), .A2(n2279), .ZN(n4642) );
  XNOR2_X1 U2941 ( .A(n4442), .B(n4345), .ZN(n4532) );
  INV_X1 U2942 ( .A(n4532), .ZN(n2235) );
  INV_X1 U2943 ( .A(IR_REG_14__SCAN_IN), .ZN(n2504) );
  NAND2_X1 U2944 ( .A1(n2940), .A2(n2939), .ZN(n2173) );
  NAND2_X1 U2945 ( .A1(n2249), .A2(n4305), .ZN(n3600) );
  NAND2_X1 U2946 ( .A1(n2397), .A2(n2398), .ZN(n3498) );
  NAND2_X1 U2947 ( .A1(n3169), .A2(n4307), .ZN(n3484) );
  NAND2_X1 U2948 ( .A1(n2213), .A2(n3140), .ZN(n4684) );
  XOR2_X1 U2949 ( .A(n2831), .B(n3006), .Z(n2174) );
  NAND2_X1 U2950 ( .A1(n4677), .A2(n4676), .ZN(n2175) );
  NOR3_X1 U2951 ( .A1(n4721), .A2(n4720), .A3(n5009), .ZN(n2176) );
  NAND2_X1 U2952 ( .A1(n4278), .A2(n4570), .ZN(n2177) );
  INV_X1 U2953 ( .A(n4359), .ZN(n2242) );
  NAND2_X1 U2954 ( .A1(n4868), .A2(REG2_REG_12__SCAN_IN), .ZN(n4867) );
  INV_X1 U2955 ( .A(n3688), .ZN(n3700) );
  OR2_X1 U2956 ( .A1(n4603), .A2(n3158), .ZN(n2178) );
  NOR2_X1 U2957 ( .A1(n4771), .A2(n2282), .ZN(n2280) );
  AND2_X1 U2958 ( .A1(n4581), .A2(n4600), .ZN(n2179) );
  OR2_X1 U2959 ( .A1(n3546), .A2(n4073), .ZN(n2180) );
  NOR2_X1 U2960 ( .A1(n4744), .A2(n2277), .ZN(n2276) );
  INV_X1 U2961 ( .A(n2278), .ZN(n4608) );
  NOR2_X1 U2962 ( .A1(n4744), .A2(n4606), .ZN(n2278) );
  NOR3_X1 U2963 ( .A1(n4744), .A2(n3158), .A3(n4606), .ZN(n4569) );
  AND2_X1 U2964 ( .A1(n4246), .A2(n2173), .ZN(n2405) );
  INV_X1 U2965 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2821) );
  AND2_X1 U2966 ( .A1(n2912), .A2(n2911), .ZN(n2181) );
  XNOR2_X1 U2967 ( .A(n2482), .B(n2481), .ZN(n4981) );
  NAND2_X1 U2968 ( .A1(n4603), .A2(n3158), .ZN(n3159) );
  INV_X1 U2969 ( .A(REG3_REG_11__SCAN_IN), .ZN(n4050) );
  OR2_X1 U2970 ( .A1(n2134), .A2(n2920), .ZN(n3200) );
  NAND2_X1 U2971 ( .A1(n4259), .A2(n3197), .ZN(n2182) );
  INV_X1 U2972 ( .A(IR_REG_0__SCAN_IN), .ZN(n2378) );
  INV_X1 U2973 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2286) );
  INV_X1 U2974 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2297) );
  XOR2_X1 U2975 ( .A(n3238), .B(REG2_REG_18__SCAN_IN), .Z(n2183) );
  INV_X1 U2976 ( .A(n4919), .ZN(n2201) );
  OR2_X1 U2977 ( .A1(n2134), .A2(n4046), .ZN(n4617) );
  NAND2_X1 U2978 ( .A1(n3442), .A2(n3443), .ZN(n3441) );
  AND2_X1 U2979 ( .A1(n4830), .A2(REG1_REG_16__SCAN_IN), .ZN(n2184) );
  NAND2_X1 U2980 ( .A1(n3448), .A2(n2697), .ZN(n3426) );
  NAND2_X1 U2981 ( .A1(n4700), .A2(n3120), .ZN(n3558) );
  OR2_X1 U2982 ( .A1(n2886), .A2(n2885), .ZN(n2185) );
  NOR2_X1 U2983 ( .A1(n2899), .A2(n2898), .ZN(n2186) );
  NAND2_X1 U2984 ( .A1(n4701), .A2(n4703), .ZN(n4700) );
  OR2_X1 U2985 ( .A1(n2183), .A2(n2500), .ZN(n2187) );
  INV_X1 U2986 ( .A(n4600), .ZN(n4606) );
  OR2_X1 U2987 ( .A1(n2134), .A2(n2961), .ZN(n4600) );
  AND2_X1 U2988 ( .A1(n2183), .A2(n2500), .ZN(n2188) );
  INV_X1 U2989 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4226) );
  AND2_X1 U2990 ( .A1(n2524), .A2(n2523), .ZN(n4829) );
  XNOR2_X1 U2991 ( .A(n2458), .B(n3227), .ZN(n4839) );
  AND2_X1 U2992 ( .A1(n2340), .A2(n2337), .ZN(n2189) );
  XNOR2_X1 U2993 ( .A(n2587), .B(n4830), .ZN(n2372) );
  XNOR2_X1 U2994 ( .A(n2495), .B(n4830), .ZN(n4474) );
  INV_X1 U2995 ( .A(n4830), .ZN(n2371) );
  OR2_X1 U2996 ( .A1(n2495), .A2(n4830), .ZN(n2496) );
  NAND3_X1 U2997 ( .A1(n2193), .A2(n2195), .A3(n2190), .ZN(n3297) );
  NAND3_X1 U2998 ( .A1(n2193), .A2(n2191), .A3(n2190), .ZN(n2198) );
  NAND2_X1 U2999 ( .A1(n2199), .A2(n4832), .ZN(n2197) );
  NOR2_X2 U3000 ( .A1(n4885), .A2(n2487), .ZN(n4898) );
  NOR2_X2 U3001 ( .A1(n4886), .A2(n4887), .ZN(n4885) );
  NOR2_X2 U3002 ( .A1(n2611), .A2(n2610), .ZN(n2613) );
  AND2_X2 U3003 ( .A1(n4917), .A2(n2188), .ZN(n2611) );
  NAND3_X1 U3004 ( .A1(n2442), .A2(n2378), .A3(n2377), .ZN(n2449) );
  OR2_X2 U3005 ( .A1(n2629), .A2(n4827), .ZN(n3308) );
  NAND2_X1 U3006 ( .A1(n2210), .A2(n2209), .ZN(n3587) );
  INV_X1 U3007 ( .A(n3509), .ZN(n2214) );
  AOI21_X2 U3008 ( .B1(n2212), .B2(n2211), .A(n2165), .ZN(n2209) );
  NAND2_X1 U3009 ( .A1(n2212), .A2(n3509), .ZN(n2210) );
  INV_X1 U3010 ( .A(n2216), .ZN(n3161) );
  OAI21_X1 U3011 ( .B1(n4701), .B2(n2225), .A(n2223), .ZN(n3406) );
  OR2_X2 U3012 ( .A1(n2449), .A2(n2229), .ZN(n2532) );
  NAND2_X1 U3013 ( .A1(n3169), .A2(n2167), .ZN(n3527) );
  NAND2_X1 U3014 ( .A1(n3527), .A2(n3174), .ZN(n3189) );
  NAND2_X1 U3015 ( .A1(n3195), .A2(n2246), .ZN(n2245) );
  NAND2_X1 U3016 ( .A1(n2245), .A2(n4409), .ZN(n4634) );
  MUX2_X1 U3017 ( .A(n3957), .B(n2551), .S(n2735), .Z(n3379) );
  MUX2_X1 U3018 ( .A(n2259), .B(n2378), .S(n2735), .Z(n4947) );
  OAI211_X1 U3019 ( .C1(n4722), .C2(n3224), .A(n2263), .B(n2261), .ZN(U3547)
         );
  NAND3_X1 U3020 ( .A1(n2265), .A2(n2264), .A3(n5030), .ZN(n2263) );
  INV_X1 U3021 ( .A(n4690), .ZN(n2273) );
  NAND2_X1 U3022 ( .A1(n2273), .A2(n2274), .ZN(n3682) );
  NAND3_X1 U3023 ( .A1(n4589), .A2(n4600), .A3(n4570), .ZN(n2277) );
  NAND2_X1 U3024 ( .A1(n2533), .A2(n2333), .ZN(n2624) );
  NAND2_X1 U3025 ( .A1(n2645), .A2(REG3_REG_1__SCAN_IN), .ZN(n2649) );
  NAND2_X1 U3026 ( .A1(n4403), .A2(n4367), .ZN(n3718) );
  NAND2_X1 U3027 ( .A1(n2284), .A2(n2172), .ZN(n2765) );
  NAND2_X1 U3028 ( .A1(n2887), .A2(REG3_REG_18__SCAN_IN), .ZN(n2900) );
  NAND2_X1 U3029 ( .A1(n2941), .A2(n2298), .ZN(n2986) );
  INV_X1 U3030 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2300) );
  NAND3_X1 U3031 ( .A1(n4295), .A2(n4294), .A3(n2302), .ZN(n4297) );
  NAND2_X1 U3032 ( .A1(n2307), .A2(n2308), .ZN(n3149) );
  NAND2_X1 U3033 ( .A1(n3659), .A2(n2310), .ZN(n2307) );
  OR2_X1 U3034 ( .A1(n2320), .A2(n2318), .ZN(n4494) );
  NOR2_X1 U3035 ( .A1(n3161), .A2(n4357), .ZN(n2321) );
  INV_X1 U3036 ( .A(n2511), .ZN(n2332) );
  NOR2_X1 U3037 ( .A1(n2510), .A2(IR_REG_28__SCAN_IN), .ZN(n2331) );
  NAND3_X1 U3038 ( .A1(n2329), .A2(n2330), .A3(n2326), .ZN(n3230) );
  NOR2_X1 U3039 ( .A1(n2511), .A2(n2510), .ZN(n2533) );
  NAND4_X1 U3040 ( .A1(n2329), .A2(n2408), .A3(n2332), .A4(n2331), .ZN(n2328)
         );
  NAND2_X1 U3041 ( .A1(n2339), .A2(n2343), .ZN(n2336) );
  NAND2_X1 U3042 ( .A1(n2339), .A2(n2338), .ZN(n2337) );
  NAND2_X1 U3043 ( .A1(n2341), .A2(n2458), .ZN(n2340) );
  INV_X1 U3044 ( .A(n2344), .ZN(n3275) );
  NAND2_X1 U3045 ( .A1(n3265), .A2(n2168), .ZN(n2346) );
  XNOR2_X1 U3046 ( .A(n2350), .B(n2349), .ZN(n3296) );
  INV_X1 U3047 ( .A(n2563), .ZN(n2351) );
  NAND2_X1 U3048 ( .A1(n3301), .A2(n2357), .ZN(n2356) );
  NAND2_X1 U3049 ( .A1(n4469), .A2(n4468), .ZN(n4467) );
  NAND2_X1 U3050 ( .A1(n3300), .A2(n2569), .ZN(n4469) );
  OAI21_X2 U3051 ( .B1(n4879), .B2(n4876), .A(n2359), .ZN(n2486) );
  NAND2_X1 U3052 ( .A1(n2576), .A2(n2360), .ZN(n2361) );
  INV_X1 U3053 ( .A(n2364), .ZN(n4862) );
  NAND2_X1 U3054 ( .A1(n2575), .A2(n2574), .ZN(n4863) );
  INV_X1 U3055 ( .A(n3541), .ZN(n2369) );
  AOI21_X2 U3056 ( .B1(n2587), .B2(n2370), .A(n2184), .ZN(n4915) );
  XNOR2_X1 U3057 ( .A(n2372), .B(n4473), .ZN(n4480) );
  NAND2_X1 U3058 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2374)
         );
  NAND3_X1 U3059 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .A3(
        IR_REG_1__SCAN_IN), .ZN(n2375) );
  NAND2_X1 U3060 ( .A1(n2376), .A2(n3376), .ZN(n3385) );
  NAND2_X1 U3061 ( .A1(n2667), .A2(n2666), .ZN(n2376) );
  XNOR2_X1 U3062 ( .A(n3376), .B(n2376), .ZN(n3383) );
  NAND2_X1 U3063 ( .A1(IR_REG_31__SCAN_IN), .A2(n3927), .ZN(n2443) );
  NAND3_X1 U3064 ( .A1(n3442), .A2(n2697), .A3(n3443), .ZN(n2379) );
  OAI211_X1 U3065 ( .C1(n2693), .C2(n2380), .A(n3427), .B(n2379), .ZN(n2713)
         );
  NAND2_X1 U3066 ( .A1(n3731), .A2(n2384), .ZN(n2382) );
  OAI21_X1 U3067 ( .B1(n3731), .B2(n2387), .A(n2384), .ZN(n3894) );
  INV_X1 U3068 ( .A(n3862), .ZN(n2844) );
  NAND2_X1 U3069 ( .A1(n2397), .A2(n2395), .ZN(n2820) );
  NAND2_X1 U3070 ( .A1(n3395), .A2(n2399), .ZN(n2397) );
  NAND2_X1 U3071 ( .A1(n3909), .A2(n2405), .ZN(n2402) );
  NOR2_X1 U3072 ( .A1(n2532), .A2(IR_REG_5__SCAN_IN), .ZN(n2435) );
  AND2_X2 U3073 ( .A1(n2408), .A2(n2409), .ZN(n2512) );
  NAND3_X1 U3074 ( .A1(n2409), .A2(n2408), .A3(n2332), .ZN(n2521) );
  NAND2_X1 U3075 ( .A1(n3632), .A2(n3626), .ZN(n4690) );
  NOR2_X1 U3076 ( .A1(n4719), .A2(n4514), .ZN(n4515) );
  INV_X1 U3077 ( .A(n2995), .ZN(n2996) );
  OAI21_X1 U3078 ( .B1(n2644), .B2(n2643), .A(n2671), .ZN(n3388) );
  INV_X1 U3079 ( .A(n2484), .ZN(n2483) );
  OAI21_X1 U3080 ( .B1(n2519), .B2(n4003), .A(n2518), .ZN(n3078) );
  NOR2_X1 U3081 ( .A1(n4871), .A2(n2577), .ZN(n2579) );
  XNOR2_X1 U3082 ( .A(n2484), .B(n4981), .ZN(n4868) );
  NAND2_X1 U3083 ( .A1(n3226), .A2(n4975), .ZN(n3242) );
  OR2_X1 U3084 ( .A1(n2638), .A2(REG2_REG_2__SCAN_IN), .ZN(n2444) );
  AND2_X1 U3085 ( .A1(n3285), .A2(n2564), .ZN(n2411) );
  INV_X2 U3086 ( .A(n4447), .ZN(U4043) );
  OR2_X1 U3087 ( .A1(n4464), .A2(n3636), .ZN(n2412) );
  NOR2_X1 U3088 ( .A1(n2763), .A2(n3361), .ZN(n2413) );
  AND2_X1 U3089 ( .A1(n5030), .A2(n4786), .ZN(n2414) );
  AND2_X1 U3090 ( .A1(n3224), .A2(REG1_REG_31__SCAN_IN), .ZN(n2415) );
  AND2_X1 U3091 ( .A1(n2572), .A2(REG1_REG_11__SCAN_IN), .ZN(n2416) );
  AND2_X1 U3092 ( .A1(n4834), .A2(REG1_REG_5__SCAN_IN), .ZN(n2417) );
  AND2_X1 U3093 ( .A1(n3907), .A2(n3906), .ZN(n2418) );
  XNOR2_X1 U3094 ( .A(REG1_REG_19__SCAN_IN), .B(n4433), .ZN(n2419) );
  INV_X1 U3095 ( .A(IR_REG_28__SCAN_IN), .ZN(n2537) );
  INV_X1 U3096 ( .A(n4430), .ZN(n3105) );
  AND2_X1 U3097 ( .A1(n2980), .A2(n2979), .ZN(n2420) );
  NAND2_X1 U3098 ( .A1(n2949), .A2(n2948), .ZN(n4639) );
  AND2_X1 U3099 ( .A1(n3223), .A2(n3222), .ZN(n2421) );
  NAND2_X1 U3100 ( .A1(n2519), .A2(n4003), .ZN(n2518) );
  INV_X1 U3101 ( .A(n5030), .ZN(n3224) );
  INV_X2 U3102 ( .A(n5019), .ZN(n5020) );
  OR2_X1 U3103 ( .A1(n4718), .A2(n4717), .ZN(n2422) );
  AND3_X1 U3104 ( .A1(n3066), .A2(n3069), .A3(n4247), .ZN(n2423) );
  AND2_X1 U3105 ( .A1(n3740), .A2(n4378), .ZN(n2424) );
  AND2_X1 U3106 ( .A1(n3096), .A2(n3095), .ZN(n2425) );
  NOR2_X1 U3107 ( .A1(n3242), .A2(n3106), .ZN(n2426) );
  INV_X1 U3108 ( .A(n4923), .ZN(n4902) );
  INV_X1 U3109 ( .A(n4224), .ZN(n2977) );
  AND3_X1 U3110 ( .A1(n2528), .A2(n2527), .A3(n2534), .ZN(n2529) );
  NAND2_X1 U3111 ( .A1(n2978), .A2(n2977), .ZN(n2979) );
  INV_X1 U3112 ( .A(n4589), .ZN(n3158) );
  INV_X1 U3113 ( .A(n3379), .ZN(n3115) );
  INV_X1 U3114 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4043) );
  INV_X1 U3115 ( .A(n3863), .ZN(n2843) );
  NAND2_X1 U3116 ( .A1(n2638), .A2(n2627), .ZN(n2553) );
  INV_X1 U3117 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2845) );
  OR2_X1 U3118 ( .A1(n3139), .A2(n3138), .ZN(n3140) );
  INV_X1 U3119 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4092) );
  NAND2_X1 U3120 ( .A1(n2762), .A2(n3467), .ZN(n3359) );
  AND2_X1 U3121 ( .A1(n2873), .A2(n4204), .ZN(n2874) );
  OAI21_X1 U3122 ( .B1(n2681), .B2(n3602), .A(n2688), .ZN(n2689) );
  INV_X1 U3123 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2927) );
  OAI22_X1 U3124 ( .A1(n4940), .A2(n2681), .B1(n3390), .B2(n2748), .ZN(n2642)
         );
  NAND2_X1 U3125 ( .A1(n2995), .A2(REG3_REG_26__SCAN_IN), .ZN(n3016) );
  OR2_X1 U3126 ( .A1(n4587), .A2(n2767), .ZN(n2974) );
  AND2_X1 U3127 ( .A1(n3238), .A2(REG2_REG_18__SCAN_IN), .ZN(n2610) );
  NAND2_X1 U3128 ( .A1(n4639), .A2(n3155), .ZN(n3156) );
  AND2_X1 U3129 ( .A1(n4657), .A2(n3910), .ZN(n4411) );
  INV_X1 U3130 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2764) );
  OR2_X1 U3131 ( .A1(n3092), .A2(n3091), .ZN(n4277) );
  NOR2_X1 U3132 ( .A1(n3089), .A2(n3088), .ZN(n4436) );
  OR2_X1 U3133 ( .A1(n4609), .A2(n2767), .ZN(n2960) );
  AND2_X1 U3134 ( .A1(n2560), .A2(n4845), .ZN(n2561) );
  INV_X1 U3135 ( .A(n4832), .ZN(n2566) );
  INV_X1 U3136 ( .A(REG3_REG_17__SCAN_IN), .ZN(n3734) );
  OR2_X1 U3137 ( .A1(n4639), .A2(n4617), .ZN(n4596) );
  NAND2_X1 U3138 ( .A1(n3073), .A2(n3072), .ZN(n4682) );
  INV_X1 U3139 ( .A(n3390), .ZN(n4710) );
  INV_X1 U3140 ( .A(n4952), .ZN(n4678) );
  AND2_X1 U3141 ( .A1(n3790), .A2(n3750), .ZN(n3764) );
  INV_X1 U3142 ( .A(n3485), .ZN(n3490) );
  INV_X1 U3143 ( .A(n3182), .ZN(n3667) );
  INV_X1 U3144 ( .A(n3579), .ZN(n3582) );
  INV_X1 U3145 ( .A(n4978), .ZN(n4890) );
  AND2_X1 U3146 ( .A1(n3254), .A2(n3339), .ZN(n4923) );
  AOI21_X1 U3147 ( .B1(n4632), .B2(n3154), .A(n3153), .ZN(n4616) );
  INV_X1 U31480 ( .A(n4704), .ZN(n4949) );
  AND2_X1 U31490 ( .A1(n3081), .A2(n3108), .ZN(n4954) );
  OAI22_X1 U3150 ( .A1(n3061), .A2(D_REG_0__SCAN_IN), .B1(n3047), .B2(n3244), 
        .ZN(n3416) );
  INV_X1 U3151 ( .A(n5017), .ZN(n5009) );
  OR3_X1 U3152 ( .A1(n3415), .A2(n3417), .A3(n3108), .ZN(n3214) );
  AND2_X1 U3153 ( .A1(n2546), .A2(n2545), .ZN(n4914) );
  NAND2_X1 U3154 ( .A1(n3065), .A2(n3064), .ZN(n4285) );
  INV_X1 U3155 ( .A(n3689), .ZN(n4444) );
  OR2_X1 U3156 ( .A1(n3226), .A2(n3245), .ZN(n4447) );
  INV_X1 U3157 ( .A(n4921), .ZN(n4896) );
  INV_X1 U3158 ( .A(n4914), .ZN(n4911) );
  OR2_X1 U3159 ( .A1(n3771), .A2(n4779), .ZN(n4646) );
  NAND2_X1 U3160 ( .A1(n4958), .A2(n3483), .ZN(n4649) );
  NAND2_X1 U3161 ( .A1(n5030), .A2(n2138), .ZN(n4761) );
  NAND2_X1 U3162 ( .A1(n5020), .A2(n2138), .ZN(n4820) );
  OR2_X1 U3163 ( .A1(n3214), .A2(n3213), .ZN(n5019) );
  INV_X1 U3164 ( .A(n4974), .ZN(n4973) );
  OR2_X1 U3165 ( .A1(n2434), .A2(n2433), .ZN(n4978) );
  OAI21_X1 U3166 ( .B1(n4788), .B2(n4761), .A(n3114), .ZN(U3549) );
  OAI21_X1 U3167 ( .B1(n3225), .B2(n5019), .A(n3220), .ZN(U3514) );
  INV_X2 U3168 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  NAND2_X1 U3169 ( .A1(n2512), .A2(n2504), .ZN(n2488) );
  OAI21_X1 U3170 ( .B1(n2497), .B2(IR_REG_17__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2431) );
  XNOR2_X1 U3171 ( .A(n2431), .B(IR_REG_18__SCAN_IN), .ZN(n3238) );
  NOR2_X1 U3172 ( .A1(n2512), .A2(n2535), .ZN(n2432) );
  MUX2_X1 U3173 ( .A(n2535), .B(n2432), .S(IR_REG_14__SCAN_IN), .Z(n2434) );
  INV_X1 U3174 ( .A(n2488), .ZN(n2433) );
  NAND2_X1 U3175 ( .A1(n2435), .A2(n2436), .ZN(n2466) );
  NAND2_X1 U3176 ( .A1(n2473), .A2(n2474), .ZN(n2477) );
  NAND2_X1 U3177 ( .A1(n2478), .A2(n2481), .ZN(n2437) );
  OAI21_X1 U3178 ( .B1(n2477), .B2(n2437), .A(IR_REG_31__SCAN_IN), .ZN(n2438)
         );
  INV_X1 U3179 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4877) );
  NOR2_X1 U3180 ( .A1(n4980), .A2(n4877), .ZN(n4876) );
  NAND2_X1 U3181 ( .A1(n2551), .A2(REG2_REG_1__SCAN_IN), .ZN(n2439) );
  NAND2_X1 U3182 ( .A1(n2440), .A2(n2439), .ZN(n4454) );
  AND2_X1 U3183 ( .A1(REG2_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2441)
         );
  NAND2_X1 U3184 ( .A1(n4454), .A2(n2441), .ZN(n3324) );
  INV_X1 U3185 ( .A(n2551), .ZN(n4837) );
  NAND2_X1 U3186 ( .A1(n4837), .A2(REG2_REG_1__SCAN_IN), .ZN(n3326) );
  NAND2_X1 U3187 ( .A1(n3324), .A2(n3326), .ZN(n2447) );
  XNOR2_X2 U3188 ( .A(n2443), .B(n2442), .ZN(n2638) );
  NAND2_X1 U3189 ( .A1(n2638), .A2(REG2_REG_2__SCAN_IN), .ZN(n2445) );
  INV_X1 U3190 ( .A(REG2_REG_2__SCAN_IN), .ZN(n4708) );
  NAND2_X1 U3191 ( .A1(n2445), .A2(n2444), .ZN(n2446) );
  NAND2_X1 U3192 ( .A1(n2447), .A2(n2446), .ZN(n3328) );
  INV_X1 U3193 ( .A(n2638), .ZN(n4836) );
  NAND2_X1 U3194 ( .A1(n4836), .A2(REG2_REG_2__SCAN_IN), .ZN(n2448) );
  NAND2_X1 U3195 ( .A1(n3328), .A2(n2448), .ZN(n2450) );
  XNOR2_X1 U3196 ( .A(n2454), .B(IR_REG_3__SCAN_IN), .ZN(n4835) );
  INV_X1 U3197 ( .A(n4835), .ZN(n3264) );
  XNOR2_X1 U3198 ( .A(n2450), .B(n3264), .ZN(n3259) );
  NAND2_X1 U3199 ( .A1(n3259), .A2(REG2_REG_3__SCAN_IN), .ZN(n2452) );
  NAND2_X1 U3200 ( .A1(n2450), .A2(n4835), .ZN(n2451) );
  NAND2_X1 U3201 ( .A1(n2454), .A2(n2453), .ZN(n2455) );
  NAND2_X1 U3202 ( .A1(n2455), .A2(IR_REG_31__SCAN_IN), .ZN(n2457) );
  INV_X1 U3203 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2462) );
  NAND2_X1 U3204 ( .A1(n2532), .A2(IR_REG_31__SCAN_IN), .ZN(n2459) );
  MUX2_X1 U3205 ( .A(n2459), .B(IR_REG_31__SCAN_IN), .S(n2528), .Z(n2461) );
  INV_X1 U3206 ( .A(n2435), .ZN(n2460) );
  MUX2_X1 U3207 ( .A(n2462), .B(REG2_REG_5__SCAN_IN), .S(n4834), .Z(n3276) );
  OR2_X1 U3208 ( .A1(n2435), .A2(n2535), .ZN(n2463) );
  XNOR2_X1 U3209 ( .A(n2463), .B(IR_REG_6__SCAN_IN), .ZN(n4833) );
  INV_X1 U32100 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3492) );
  NAND2_X1 U32110 ( .A1(n2466), .A2(IR_REG_31__SCAN_IN), .ZN(n2468) );
  XNOR2_X1 U32120 ( .A(n2468), .B(n2467), .ZN(n3285) );
  MUX2_X1 U32130 ( .A(REG2_REG_7__SCAN_IN), .B(n3492), .S(n3285), .Z(n3290) );
  INV_X1 U32140 ( .A(n3285), .ZN(n3294) );
  NAND2_X1 U32150 ( .A1(n2468), .A2(n2467), .ZN(n2469) );
  NAND2_X1 U32160 ( .A1(n2469), .A2(IR_REG_31__SCAN_IN), .ZN(n2470) );
  XNOR2_X1 U32170 ( .A(n2470), .B(IR_REG_8__SCAN_IN), .ZN(n4832) );
  INV_X1 U32180 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3613) );
  INV_X1 U32190 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3636) );
  NAND2_X1 U32200 ( .A1(n2471), .A2(IR_REG_31__SCAN_IN), .ZN(n2472) );
  MUX2_X1 U32210 ( .A(REG2_REG_9__SCAN_IN), .B(n3636), .S(n4831), .Z(n4461) );
  INV_X1 U32220 ( .A(n4831), .ZN(n4464) );
  OR2_X1 U32230 ( .A1(n2473), .A2(n2535), .ZN(n2475) );
  NAND2_X1 U32240 ( .A1(n2476), .A2(n2776), .ZN(n3542) );
  INV_X1 U32250 ( .A(REG2_REG_11__SCAN_IN), .ZN(n4073) );
  NAND2_X1 U32260 ( .A1(n2477), .A2(IR_REG_31__SCAN_IN), .ZN(n2479) );
  MUX2_X1 U32270 ( .A(REG2_REG_11__SCAN_IN), .B(n4073), .S(n3546), .Z(n3541)
         );
  INV_X1 U32280 ( .A(n3546), .ZN(n2572) );
  NAND2_X1 U32290 ( .A1(n2479), .A2(n2478), .ZN(n2480) );
  NAND2_X1 U32300 ( .A1(n2480), .A2(IR_REG_31__SCAN_IN), .ZN(n2482) );
  OR2_X1 U32310 ( .A1(n2483), .A2(n4981), .ZN(n2485) );
  NOR2_X1 U32320 ( .A1(n4978), .A2(n2486), .ZN(n2487) );
  INV_X1 U32330 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4887) );
  NAND2_X1 U32340 ( .A1(n2488), .A2(IR_REG_31__SCAN_IN), .ZN(n2492) );
  INV_X1 U32350 ( .A(REG2_REG_15__SCAN_IN), .ZN(n3802) );
  OR2_X1 U32360 ( .A1(n4907), .A2(n3802), .ZN(n2490) );
  NAND2_X1 U32370 ( .A1(n4907), .A2(n3802), .ZN(n2489) );
  AND2_X1 U32380 ( .A1(n2490), .A2(n2489), .ZN(n4897) );
  NAND2_X1 U32390 ( .A1(n4907), .A2(REG2_REG_15__SCAN_IN), .ZN(n2491) );
  INV_X1 U32400 ( .A(IR_REG_15__SCAN_IN), .ZN(n3956) );
  NAND2_X1 U32410 ( .A1(n2492), .A2(n3956), .ZN(n2493) );
  NAND2_X1 U32420 ( .A1(n2493), .A2(IR_REG_31__SCAN_IN), .ZN(n2494) );
  XNOR2_X1 U32430 ( .A(n2494), .B(IR_REG_16__SCAN_IN), .ZN(n4830) );
  NAND2_X1 U32440 ( .A1(n2497), .A2(IR_REG_31__SCAN_IN), .ZN(n2498) );
  XNOR2_X1 U32450 ( .A(n2498), .B(IR_REG_17__SCAN_IN), .ZN(n2588) );
  NOR2_X1 U32460 ( .A1(n2588), .A2(REG2_REG_17__SCAN_IN), .ZN(n2499) );
  AOI21_X1 U32470 ( .B1(REG2_REG_17__SCAN_IN), .B2(n2588), .A(n2499), .ZN(
        n4919) );
  OR2_X1 U32480 ( .A1(n2588), .A2(REG2_REG_17__SCAN_IN), .ZN(n2500) );
  INV_X1 U32490 ( .A(n2601), .ZN(n2505) );
  NOR2_X1 U32500 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2509) );
  NAND3_X1 U32510 ( .A1(n2515), .A2(n2509), .A3(n4003), .ZN(n2510) );
  INV_X1 U32520 ( .A(n2526), .ZN(n2513) );
  NAND2_X1 U32530 ( .A1(n2515), .A2(n4003), .ZN(n2516) );
  OAI21_X2 U32540 ( .B1(n2523), .B2(n2516), .A(IR_REG_31__SCAN_IN), .ZN(n2517)
         );
  NAND3_X2 U32550 ( .A1(n3047), .A2(n3244), .A3(n3045), .ZN(n3226) );
  OR2_X1 U32560 ( .A1(n3078), .A2(U3149), .ZN(n4439) );
  NAND2_X1 U32570 ( .A1(n3242), .A2(n4439), .ZN(n2546) );
  NAND2_X1 U32580 ( .A1(n2523), .A2(IR_REG_31__SCAN_IN), .ZN(n2520) );
  NAND2_X1 U32590 ( .A1(n2521), .A2(IR_REG_31__SCAN_IN), .ZN(n2522) );
  MUX2_X1 U32600 ( .A(IR_REG_31__SCAN_IN), .B(n2522), .S(IR_REG_21__SCAN_IN), 
        .Z(n2524) );
  NAND2_X1 U32610 ( .A1(n2530), .A2(n2529), .ZN(n2531) );
  NAND2_X1 U32620 ( .A1(n2535), .A2(n2534), .ZN(n2536) );
  NAND2_X1 U32630 ( .A1(n2624), .A2(n2536), .ZN(n2539) );
  AOI21_X1 U32640 ( .B1(n3209), .B2(n3078), .A(n2134), .ZN(n2544) );
  INV_X1 U32650 ( .A(n2538), .ZN(n2541) );
  INV_X1 U32660 ( .A(n2539), .ZN(n2540) );
  NAND2_X1 U32670 ( .A1(n2541), .A2(n2540), .ZN(n3339) );
  NAND2_X1 U32680 ( .A1(n2624), .A2(IR_REG_31__SCAN_IN), .ZN(n2542) );
  XNOR2_X1 U32690 ( .A(n2542), .B(n2537), .ZN(n4838) );
  NOR2_X1 U32700 ( .A1(n3339), .A2(n4838), .ZN(n4435) );
  NAND2_X1 U32710 ( .A1(n2543), .A2(n4921), .ZN(n2550) );
  INV_X1 U32720 ( .A(n3238), .ZN(n2895) );
  INV_X1 U32730 ( .A(n2544), .ZN(n2545) );
  NOR2_X1 U32740 ( .A1(n2297), .A2(STATE_REG_SCAN_IN), .ZN(n4258) );
  AOI21_X1 U32750 ( .B1(n4914), .B2(ADDR_REG_18__SCAN_IN), .A(n4258), .ZN(
        n2547) );
  OAI21_X1 U32760 ( .B1(n4926), .B2(n2895), .A(n2547), .ZN(n2548) );
  INV_X1 U32770 ( .A(n2548), .ZN(n2549) );
  NAND2_X1 U32780 ( .A1(n2550), .A2(n2549), .ZN(n2596) );
  NAND2_X1 U32790 ( .A1(n3238), .A2(REG1_REG_18__SCAN_IN), .ZN(n2597) );
  OAI21_X1 U32800 ( .B1(n3238), .B2(REG1_REG_18__SCAN_IN), .A(n2597), .ZN(
        n2594) );
  OR2_X1 U32810 ( .A1(n2588), .A2(REG1_REG_17__SCAN_IN), .ZN(n2589) );
  INV_X1 U32820 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4855) );
  INV_X1 U32830 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2646) );
  NAND2_X1 U32840 ( .A1(n2551), .A2(REG1_REG_1__SCAN_IN), .ZN(n2552) );
  AND2_X1 U32850 ( .A1(REG1_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n4453) );
  NAND2_X1 U32860 ( .A1(n4452), .A2(n4453), .ZN(n4451) );
  NAND2_X1 U32870 ( .A1(n4837), .A2(REG1_REG_1__SCAN_IN), .ZN(n3330) );
  NAND2_X1 U32880 ( .A1(n4451), .A2(n3330), .ZN(n2555) );
  INV_X1 U32890 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2627) );
  OAI21_X1 U32900 ( .B1(n2638), .B2(n2627), .A(n2553), .ZN(n3329) );
  INV_X1 U32910 ( .A(n3329), .ZN(n2554) );
  NAND2_X1 U32920 ( .A1(n4836), .A2(REG1_REG_2__SCAN_IN), .ZN(n2556) );
  NAND2_X1 U32930 ( .A1(n3258), .A2(REG1_REG_3__SCAN_IN), .ZN(n2559) );
  NAND2_X1 U32940 ( .A1(n2557), .A2(n4835), .ZN(n2558) );
  INV_X1 U32950 ( .A(REG1_REG_5__SCAN_IN), .ZN(n5027) );
  MUX2_X1 U32960 ( .A(n5027), .B(REG1_REG_5__SCAN_IN), .S(n4834), .Z(n3278) );
  NOR2_X1 U32970 ( .A1(n3279), .A2(n3278), .ZN(n3277) );
  NOR2_X1 U32980 ( .A1(n2562), .A2(n3268), .ZN(n2563) );
  NAND2_X1 U32990 ( .A1(n3294), .A2(REG1_REG_7__SCAN_IN), .ZN(n2565) );
  INV_X1 U33000 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2564) );
  INV_X1 U33010 ( .A(n2567), .ZN(n2568) );
  XOR2_X1 U33020 ( .A(REG1_REG_9__SCAN_IN), .B(n4831), .Z(n4468) );
  INV_X1 U33030 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2768) );
  AND2_X1 U33040 ( .A1(n2570), .A2(n2776), .ZN(n2571) );
  XOR2_X1 U33050 ( .A(REG1_REG_11__SCAN_IN), .B(n3546), .Z(n3538) );
  NOR2_X1 U33060 ( .A1(n2573), .A2(n4981), .ZN(n2576) );
  INV_X1 U33070 ( .A(n2576), .ZN(n2575) );
  NAND2_X1 U33080 ( .A1(n2573), .A2(n4981), .ZN(n2574) );
  INV_X1 U33090 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4864) );
  INV_X1 U33100 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3779) );
  AOI22_X1 U33110 ( .A1(n2828), .A2(n3779), .B1(REG1_REG_13__SCAN_IN), .B2(
        n4980), .ZN(n4872) );
  INV_X1 U33120 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4884) );
  NAND2_X1 U33130 ( .A1(n4907), .A2(REG1_REG_15__SCAN_IN), .ZN(n2580) );
  XNOR2_X1 U33140 ( .A(n4907), .B(REG1_REG_15__SCAN_IN), .ZN(n4903) );
  AND2_X1 U33150 ( .A1(n2580), .A2(n4903), .ZN(n2582) );
  OR2_X1 U33160 ( .A1(n4884), .A2(n2582), .ZN(n2578) );
  INV_X1 U33170 ( .A(n4900), .ZN(n2581) );
  INV_X1 U33180 ( .A(n2582), .ZN(n2583) );
  NAND2_X1 U33190 ( .A1(n2584), .A2(n2583), .ZN(n2585) );
  NAND2_X1 U33200 ( .A1(n2586), .A2(n2585), .ZN(n2587) );
  INV_X1 U33210 ( .A(REG1_REG_17__SCAN_IN), .ZN(n3798) );
  AOI22_X1 U33220 ( .A1(n2588), .A2(REG1_REG_17__SCAN_IN), .B1(n3798), .B2(
        n4976), .ZN(n4916) );
  NAND2_X1 U33230 ( .A1(n4915), .A2(n4916), .ZN(n2592) );
  NAND2_X1 U33240 ( .A1(n2589), .A2(n2592), .ZN(n2593) );
  INV_X1 U33250 ( .A(n2594), .ZN(n2590) );
  AND2_X1 U33260 ( .A1(n2590), .A2(n2589), .ZN(n2591) );
  AOI211_X1 U33270 ( .C1(n2594), .C2(n2593), .A(n2599), .B(n4902), .ZN(n2595)
         );
  OR2_X1 U33280 ( .A1(n2596), .A2(n2595), .ZN(U3258) );
  INV_X1 U33290 ( .A(n2597), .ZN(n2598) );
  NOR2_X2 U33300 ( .A1(n2599), .A2(n2598), .ZN(n2608) );
  INV_X1 U33310 ( .A(n2600), .ZN(n2602) );
  NOR2_X1 U33320 ( .A1(n2602), .A2(n2601), .ZN(n2603) );
  NAND2_X1 U33330 ( .A1(n2512), .A2(n2603), .ZN(n2604) );
  XNOR2_X1 U33340 ( .A(n2608), .B(n2419), .ZN(n2609) );
  NAND2_X1 U33350 ( .A1(n2609), .A2(n4923), .ZN(n2619) );
  INV_X1 U33360 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4188) );
  MUX2_X1 U33370 ( .A(n4188), .B(REG2_REG_19__SCAN_IN), .S(n4433), .Z(n2612)
         );
  XNOR2_X1 U33380 ( .A(n2613), .B(n2612), .ZN(n2614) );
  NAND2_X1 U33390 ( .A1(n2614), .A2(n4921), .ZN(n2618) );
  NAND2_X1 U33400 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3898) );
  NAND2_X1 U33410 ( .A1(n4914), .A2(ADDR_REG_19__SCAN_IN), .ZN(n2615) );
  OAI211_X1 U33420 ( .C1(n4926), .C2(n4433), .A(n3898), .B(n2615), .ZN(n2616)
         );
  INV_X1 U33430 ( .A(n2616), .ZN(n2617) );
  NAND3_X1 U33440 ( .A1(n2619), .A2(n2618), .A3(n2617), .ZN(U3259) );
  NAND2_X2 U33450 ( .A1(n3226), .A2(n3422), .ZN(n2748) );
  INV_X1 U33460 ( .A(n4829), .ZN(n4292) );
  INV_X1 U33470 ( .A(n3063), .ZN(n3072) );
  NOR2_X1 U33480 ( .A1(n4828), .A2(n3072), .ZN(n2623) );
  OR2_X2 U33490 ( .A1(n2748), .A2(n3109), .ZN(n2680) );
  INV_X1 U33500 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2628) );
  OR2_X1 U33510 ( .A1(n3308), .A2(n2628), .ZN(n2635) );
  INV_X1 U33520 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2630) );
  AND2_X4 U3353 ( .A1(n2629), .A2(n2632), .ZN(n2739) );
  NAND2_X1 U33540 ( .A1(n2739), .A2(REG2_REG_2__SCAN_IN), .ZN(n2633) );
  INV_X1 U3355 ( .A(n3422), .ZN(n2637) );
  INV_X1 U3356 ( .A(DATAI_2_), .ZN(n2639) );
  MUX2_X1 U3357 ( .A(n2639), .B(n2638), .S(n2735), .Z(n3390) );
  NOR2_X1 U3358 ( .A1(n2681), .A2(n3390), .ZN(n2640) );
  AND2_X1 U3359 ( .A1(n4828), .A2(n4433), .ZN(n3087) );
  INV_X1 U3360 ( .A(n3087), .ZN(n2641) );
  AND2_X2 U3361 ( .A1(n3422), .A2(n2641), .ZN(n3006) );
  XNOR2_X1 U3362 ( .A(n2642), .B(n3006), .ZN(n2643) );
  NAND2_X1 U3363 ( .A1(n2644), .A2(n2643), .ZN(n2671) );
  INV_X1 U3364 ( .A(REG0_REG_1__SCAN_IN), .ZN(n3955) );
  OR2_X1 U3365 ( .A1(n3308), .A2(n3955), .ZN(n2650) );
  NAND2_X1 U3366 ( .A1(n2739), .A2(REG2_REG_1__SCAN_IN), .ZN(n2647) );
  AND4_X2 U3367 ( .A1(n2650), .A2(n2649), .A3(n2648), .A4(n2647), .ZN(n3116)
         );
  INV_X1 U3368 ( .A(DATAI_1_), .ZN(n3957) );
  OR2_X1 U3369 ( .A1(n2748), .A2(n3379), .ZN(n2651) );
  OAI21_X1 U3370 ( .B1(n2681), .B2(n3116), .A(n2651), .ZN(n2652) );
  INV_X1 U3371 ( .A(n2669), .ZN(n2653) );
  OAI22_X1 U3372 ( .A1(n2680), .A2(n3116), .B1(n2681), .B2(n3379), .ZN(n2668)
         );
  NAND2_X1 U3373 ( .A1(n2653), .A2(n2668), .ZN(n3384) );
  INV_X1 U3374 ( .A(n3384), .ZN(n2654) );
  NOR2_X1 U3375 ( .A1(n3388), .A2(n2654), .ZN(n2670) );
  INV_X1 U3376 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2655) );
  INV_X1 U3377 ( .A(REG1_REG_0__SCAN_IN), .ZN(n5021) );
  NAND2_X1 U3378 ( .A1(n2739), .A2(REG2_REG_0__SCAN_IN), .ZN(n2657) );
  OR2_X1 U3379 ( .A1(n3308), .A2(n4987), .ZN(n2656) );
  INV_X1 U3380 ( .A(n4936), .ZN(n3378) );
  INV_X1 U3381 ( .A(n2681), .ZN(n2852) );
  INV_X1 U3382 ( .A(n3226), .ZN(n2660) );
  AOI22_X1 U3383 ( .A1(n2852), .A2(n4942), .B1(n2660), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2661) );
  OAI21_X1 U3384 ( .B1(n3040), .B2(n3378), .A(n2661), .ZN(n3338) );
  OR2_X1 U3385 ( .A1(n3378), .A2(n2681), .ZN(n2663) );
  OR2_X1 U3386 ( .A1(n2748), .A2(n4947), .ZN(n2662) );
  AND2_X1 U3387 ( .A1(n2663), .A2(n2662), .ZN(n2665) );
  OR2_X1 U3388 ( .A1(n3226), .A2(n5021), .ZN(n2664) );
  NAND2_X1 U3389 ( .A1(n2665), .A2(n2664), .ZN(n3337) );
  NAND2_X1 U3390 ( .A1(n3338), .A2(n3337), .ZN(n2667) );
  NAND2_X1 U3391 ( .A1(n2665), .A2(n3006), .ZN(n2666) );
  XNOR2_X1 U3392 ( .A(n2669), .B(n2668), .ZN(n3376) );
  NAND2_X1 U3393 ( .A1(n2670), .A2(n3385), .ZN(n3386) );
  NAND2_X1 U3394 ( .A1(n3386), .A2(n2671), .ZN(n3442) );
  INV_X1 U3395 ( .A(n4300), .ZN(n3559) );
  INV_X2 U3396 ( .A(n3308), .ZN(n3029) );
  NAND2_X1 U3397 ( .A1(n3029), .A2(REG0_REG_3__SCAN_IN), .ZN(n2677) );
  INV_X1 U3398 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2672) );
  OR2_X1 U3399 ( .A1(n2767), .A2(REG3_REG_3__SCAN_IN), .ZN(n2675) );
  INV_X1 U3400 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2673) );
  OR2_X1 U3401 ( .A1(n2137), .A2(n2673), .ZN(n2674) );
  OR2_X1 U3402 ( .A1(n2681), .A2(n3121), .ZN(n2678) );
  OAI21_X1 U3403 ( .B1(n2748), .B2(n3559), .A(n2678), .ZN(n2679) );
  XNOR2_X1 U3404 ( .A(n2679), .B(n3006), .ZN(n2691) );
  OAI22_X1 U3405 ( .A1(n3040), .A2(n3121), .B1(n2830), .B2(n3559), .ZN(n2690)
         );
  XNOR2_X1 U3406 ( .A(n2691), .B(n2690), .ZN(n3443) );
  INV_X1 U3407 ( .A(n2681), .ZN(n2838) );
  NAND2_X1 U3408 ( .A1(n2739), .A2(REG2_REG_4__SCAN_IN), .ZN(n2686) );
  INV_X1 U3409 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2682) );
  OR2_X1 U3410 ( .A1(n3308), .A2(n2682), .ZN(n2685) );
  XNOR2_X1 U3411 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(n3456) );
  OR2_X1 U3412 ( .A1(n2767), .A2(n3456), .ZN(n2684) );
  INV_X1 U3413 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4842) );
  OR2_X1 U3414 ( .A1(n2137), .A2(n4842), .ZN(n2683) );
  NAND4_X1 U3415 ( .A1(n2686), .A2(n2685), .A3(n2684), .A4(n2683), .ZN(n4445)
         );
  INV_X1 U3416 ( .A(n4445), .ZN(n3602) );
  INV_X1 U3417 ( .A(DATAI_4_), .ZN(n2687) );
  MUX2_X1 U3418 ( .A(n2687), .B(n3227), .S(n2134), .Z(n3413) );
  OR2_X1 U3419 ( .A1(n2748), .A2(n3413), .ZN(n2688) );
  XNOR2_X1 U3420 ( .A(n2689), .B(n3006), .ZN(n2694) );
  OAI22_X1 U3421 ( .A1(n3040), .A2(n3602), .B1(n2830), .B2(n3413), .ZN(n2695)
         );
  XNOR2_X1 U3422 ( .A(n2694), .B(n2695), .ZN(n3449) );
  INV_X1 U3423 ( .A(n2690), .ZN(n2692) );
  NAND2_X1 U3424 ( .A1(n2692), .A2(n2691), .ZN(n3447) );
  INV_X1 U3425 ( .A(n2694), .ZN(n2696) );
  NAND2_X1 U3426 ( .A1(n2696), .A2(n2695), .ZN(n2697) );
  NAND2_X1 U3427 ( .A1(n2739), .A2(REG2_REG_5__SCAN_IN), .ZN(n2706) );
  INV_X1 U3428 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2698) );
  OR2_X1 U3429 ( .A1(n3308), .A2(n2698), .ZN(n2705) );
  INV_X1 U3430 ( .A(n2699), .ZN(n2701) );
  INV_X1 U3431 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2700) );
  NAND2_X1 U3432 ( .A1(n2701), .A2(n2700), .ZN(n2702) );
  NAND2_X1 U3433 ( .A1(n2716), .A2(n2702), .ZN(n3607) );
  OR2_X1 U3434 ( .A1(n2767), .A2(n3607), .ZN(n2704) );
  OR2_X1 U3435 ( .A1(n2137), .A2(n5027), .ZN(n2703) );
  NAND4_X1 U3436 ( .A1(n2706), .A2(n2705), .A3(n2704), .A4(n2703), .ZN(n3349)
         );
  INV_X1 U3437 ( .A(n3349), .ZN(n3513) );
  MUX2_X1 U3438 ( .A(DATAI_5_), .B(n4834), .S(n2134), .Z(n3606) );
  OR2_X1 U3439 ( .A1(n3037), .A2(n3167), .ZN(n2707) );
  OAI21_X1 U3440 ( .B1(n2681), .B2(n3513), .A(n2707), .ZN(n2708) );
  XNOR2_X1 U3441 ( .A(n2708), .B(n3006), .ZN(n2709) );
  OAI22_X1 U3442 ( .A1(n3040), .A2(n3513), .B1(n2830), .B2(n3167), .ZN(n2710)
         );
  XNOR2_X1 U3443 ( .A(n2709), .B(n2710), .ZN(n3427) );
  INV_X1 U3444 ( .A(n2709), .ZN(n2711) );
  NAND2_X1 U3445 ( .A1(n2711), .A2(n2710), .ZN(n2712) );
  NAND2_X1 U3446 ( .A1(n2713), .A2(n2712), .ZN(n3346) );
  NAND2_X1 U3447 ( .A1(n3029), .A2(REG0_REG_6__SCAN_IN), .ZN(n2722) );
  INV_X1 U3448 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3591) );
  OR2_X1 U3449 ( .A1(n3033), .A2(n3591), .ZN(n2721) );
  INV_X1 U3450 ( .A(n2716), .ZN(n2714) );
  NAND2_X1 U3451 ( .A1(n2714), .A2(REG3_REG_6__SCAN_IN), .ZN(n2729) );
  INV_X1 U3452 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2715) );
  NAND2_X1 U3453 ( .A1(n2716), .A2(n2715), .ZN(n2717) );
  NAND2_X1 U3454 ( .A1(n2729), .A2(n2717), .ZN(n3590) );
  OR2_X1 U3455 ( .A1(n2767), .A2(n3590), .ZN(n2720) );
  INV_X1 U3456 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2718) );
  OR2_X1 U3457 ( .A1(n2137), .A2(n2718), .ZN(n2719) );
  NAND4_X1 U34580 ( .A1(n2722), .A2(n2721), .A3(n2720), .A4(n2719), .ZN(n3168)
         );
  INV_X1 U34590 ( .A(n2135), .ZN(n3486) );
  MUX2_X1 U3460 ( .A(DATAI_6_), .B(n4833), .S(n2134), .Z(n3517) );
  INV_X1 U3461 ( .A(n3517), .ZN(n2723) );
  OR2_X1 U3462 ( .A1(n2748), .A2(n2723), .ZN(n2724) );
  XNOR2_X1 U3463 ( .A(n2725), .B(n3038), .ZN(n2759) );
  OAI22_X1 U3464 ( .A1(n3040), .A2(n3486), .B1(n2681), .B2(n2723), .ZN(n2758)
         );
  AND2_X1 U3465 ( .A1(n2759), .A2(n2758), .ZN(n3466) );
  OR2_X1 U3466 ( .A1(n2137), .A2(n2564), .ZN(n2734) );
  INV_X1 U34670 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2727) );
  OR2_X1 U3468 ( .A1(n3308), .A2(n2727), .ZN(n2733) );
  NAND2_X1 U34690 ( .A1(n2739), .A2(REG2_REG_7__SCAN_IN), .ZN(n2732) );
  INV_X1 U3470 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2728) );
  NAND2_X1 U34710 ( .A1(n2729), .A2(n2728), .ZN(n2730) );
  NAND2_X1 U3472 ( .A1(n2741), .A2(n2730), .ZN(n3491) );
  OR2_X1 U34730 ( .A1(n2767), .A2(n3491), .ZN(n2731) );
  INV_X1 U3474 ( .A(n3511), .ZN(n3529) );
  INV_X1 U34750 ( .A(DATAI_7_), .ZN(n2736) );
  MUX2_X1 U3476 ( .A(n2736), .B(n3285), .S(n2735), .Z(n3485) );
  OR2_X1 U34770 ( .A1(n2748), .A2(n3485), .ZN(n2737) );
  OAI21_X1 U3478 ( .B1(n2681), .B2(n3529), .A(n2737), .ZN(n2738) );
  XNOR2_X1 U34790 ( .A(n2738), .B(n3038), .ZN(n2757) );
  OAI22_X1 U3480 ( .A1(n3040), .A2(n3529), .B1(n2830), .B2(n3485), .ZN(n2756)
         );
  AND2_X1 U34810 ( .A1(n2757), .A2(n2756), .ZN(n3361) );
  OR2_X1 U3482 ( .A1(n3466), .A2(n3361), .ZN(n3358) );
  NAND2_X1 U34830 ( .A1(n2739), .A2(REG2_REG_8__SCAN_IN), .ZN(n2747) );
  INV_X1 U3484 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2740) );
  OR2_X1 U34850 ( .A1(n3308), .A2(n2740), .ZN(n2746) );
  INV_X1 U3486 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3298) );
  NAND2_X1 U34870 ( .A1(n2741), .A2(n3298), .ZN(n2742) );
  NAND2_X1 U3488 ( .A1(n2765), .A2(n2742), .ZN(n3612) );
  OR2_X1 U34890 ( .A1(n2767), .A2(n3612), .ZN(n2745) );
  INV_X1 U3490 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2743) );
  OR2_X1 U34910 ( .A1(n2137), .A2(n2743), .ZN(n2744) );
  INV_X1 U3492 ( .A(n3629), .ZN(n3475) );
  MUX2_X1 U34930 ( .A(DATAI_8_), .B(n4832), .S(n2134), .Z(n3535) );
  OR2_X1 U3494 ( .A1(n2748), .A2(n3176), .ZN(n2749) );
  OAI21_X1 U34950 ( .B1(n2830), .B2(n3475), .A(n2749), .ZN(n2750) );
  XNOR2_X1 U3496 ( .A(n2750), .B(n3038), .ZN(n2753) );
  OAI22_X1 U34970 ( .A1(n3040), .A2(n3475), .B1(n2830), .B2(n3176), .ZN(n2752)
         );
  NAND2_X1 U3498 ( .A1(n2753), .A2(n2752), .ZN(n3365) );
  INV_X1 U34990 ( .A(n3365), .ZN(n2763) );
  OR2_X1 U3500 ( .A1(n3358), .A2(n2763), .ZN(n2751) );
  INV_X1 U35010 ( .A(n2752), .ZN(n2755) );
  INV_X1 U3502 ( .A(n2753), .ZN(n2754) );
  NAND2_X1 U35030 ( .A1(n2755), .A2(n2754), .ZN(n3367) );
  XNOR2_X1 U3504 ( .A(n2757), .B(n2756), .ZN(n3469) );
  INV_X1 U35050 ( .A(n3469), .ZN(n2762) );
  INV_X1 U35060 ( .A(n2758), .ZN(n2761) );
  INV_X1 U35070 ( .A(n2759), .ZN(n2760) );
  NAND2_X1 U35080 ( .A1(n2761), .A2(n2760), .ZN(n3467) );
  NAND2_X1 U35090 ( .A1(n2739), .A2(REG2_REG_9__SCAN_IN), .ZN(n2772) );
  INV_X1 U35100 ( .A(REG0_REG_9__SCAN_IN), .ZN(n4014) );
  OR2_X1 U35110 ( .A1(n3308), .A2(n4014), .ZN(n2771) );
  NAND2_X1 U35120 ( .A1(n2765), .A2(n2764), .ZN(n2766) );
  NAND2_X1 U35130 ( .A1(n2777), .A2(n2766), .ZN(n3635) );
  OR2_X1 U35140 ( .A1(n2767), .A2(n3635), .ZN(n2770) );
  OR2_X1 U35150 ( .A1(n2137), .A2(n2768), .ZN(n2769) );
  NAND4_X1 U35160 ( .A1(n2772), .A2(n2771), .A3(n2770), .A4(n2769), .ZN(n4680)
         );
  INV_X1 U35170 ( .A(n4680), .ZN(n3528) );
  MUX2_X1 U35180 ( .A(DATAI_9_), .B(n4831), .S(n2134), .Z(n3634) );
  OAI22_X1 U35190 ( .A1(n3040), .A2(n3528), .B1(n2830), .B2(n3626), .ZN(n2787)
         );
  INV_X1 U35200 ( .A(n2787), .ZN(n2775) );
  OR2_X1 U35210 ( .A1(n3037), .A2(n3626), .ZN(n2773) );
  OAI21_X1 U35220 ( .B1(n2681), .B2(n3528), .A(n2773), .ZN(n2774) );
  XNOR2_X1 U35230 ( .A(n2774), .B(n3006), .ZN(n2788) );
  NAND2_X1 U35240 ( .A1(n2775), .A2(n2788), .ZN(n2786) );
  MUX2_X1 U35250 ( .A(DATAI_10_), .B(n2776), .S(n2134), .Z(n4689) );
  INV_X1 U35260 ( .A(n4689), .ZN(n4683) );
  NAND2_X1 U35270 ( .A1(n3029), .A2(REG0_REG_10__SCAN_IN), .ZN(n2782) );
  INV_X1 U35280 ( .A(REG2_REG_10__SCAN_IN), .ZN(n4693) );
  OR2_X1 U35290 ( .A1(n3033), .A2(n4693), .ZN(n2781) );
  INV_X1 U35300 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4182) );
  NAND2_X1 U35310 ( .A1(n2777), .A2(n4182), .ZN(n2778) );
  NAND2_X1 U35320 ( .A1(n2797), .A2(n2778), .ZN(n4692) );
  OR2_X1 U35330 ( .A1(n2767), .A2(n4692), .ZN(n2780) );
  OR2_X1 U35340 ( .A1(n2137), .A2(n4855), .ZN(n2779) );
  NAND4_X1 U35350 ( .A1(n2782), .A2(n2781), .A3(n2780), .A4(n2779), .ZN(n3577)
         );
  INV_X1 U35360 ( .A(n3577), .ZN(n3627) );
  OR2_X1 U35370 ( .A1(n3627), .A2(n2681), .ZN(n2783) );
  OAI21_X1 U35380 ( .B1(n4683), .B2(n3037), .A(n2783), .ZN(n2784) );
  XNOR2_X1 U35390 ( .A(n2784), .B(n3038), .ZN(n2794) );
  OAI22_X1 U35400 ( .A1(n3040), .A2(n3627), .B1(n2681), .B2(n4683), .ZN(n2793)
         );
  XNOR2_X1 U35410 ( .A(n2794), .B(n2793), .ZN(n3853) );
  INV_X1 U35420 ( .A(n3853), .ZN(n2785) );
  NAND2_X1 U35430 ( .A1(n3849), .A2(n2785), .ZN(n2791) );
  INV_X1 U35440 ( .A(n2786), .ZN(n2789) );
  XNOR2_X1 U35450 ( .A(n2788), .B(n2787), .ZN(n3460) );
  OR2_X1 U35460 ( .A1(n2789), .A2(n3460), .ZN(n3851) );
  OR2_X1 U35470 ( .A1(n3853), .A2(n3851), .ZN(n2790) );
  OAI21_X1 U35480 ( .B1(n3356), .B2(n2791), .A(n2790), .ZN(n2792) );
  INV_X1 U35490 ( .A(n2792), .ZN(n3855) );
  NAND2_X1 U35500 ( .A1(n2794), .A2(n2793), .ZN(n2795) );
  NAND2_X1 U35510 ( .A1(n3855), .A2(n2795), .ZN(n3395) );
  NAND2_X1 U35520 ( .A1(n2739), .A2(REG2_REG_11__SCAN_IN), .ZN(n2803) );
  INV_X1 U35530 ( .A(REG0_REG_11__SCAN_IN), .ZN(n2796) );
  OR2_X1 U35540 ( .A1(n3308), .A2(n2796), .ZN(n2802) );
  NAND2_X1 U35550 ( .A1(n2797), .A2(n4050), .ZN(n2798) );
  NAND2_X1 U35560 ( .A1(n2808), .A2(n2798), .ZN(n3584) );
  OR2_X1 U35570 ( .A1(n2767), .A2(n3584), .ZN(n2801) );
  INV_X1 U35580 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2799) );
  OR2_X1 U35590 ( .A1(n2137), .A2(n2799), .ZN(n2800) );
  NAND4_X1 U35600 ( .A1(n2803), .A2(n2802), .A3(n2801), .A4(n2800), .ZN(n4679)
         );
  INV_X1 U35610 ( .A(n4679), .ZN(n3858) );
  INV_X1 U35620 ( .A(DATAI_11_), .ZN(n3240) );
  MUX2_X1 U35630 ( .A(n3240), .B(n3546), .S(n2134), .Z(n3579) );
  OR2_X1 U35640 ( .A1(n3037), .A2(n3579), .ZN(n2804) );
  OAI21_X1 U35650 ( .B1(n3089), .B2(n3858), .A(n2804), .ZN(n2805) );
  XNOR2_X1 U35660 ( .A(n2805), .B(n3038), .ZN(n3396) );
  OAI22_X1 U35670 ( .A1(n3040), .A2(n3858), .B1(n2830), .B2(n3579), .ZN(n3397)
         );
  INV_X1 U35680 ( .A(DATAI_12_), .ZN(n2806) );
  MUX2_X1 U35690 ( .A(n2806), .B(n4981), .S(n2134), .Z(n3182) );
  INV_X1 U35700 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4010) );
  OR2_X1 U35710 ( .A1(n3308), .A2(n4010), .ZN(n2813) );
  INV_X1 U35720 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3672) );
  OR2_X1 U35730 ( .A1(n3033), .A2(n3672), .ZN(n2812) );
  INV_X1 U35740 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4162) );
  NAND2_X1 U35750 ( .A1(n2808), .A2(n4162), .ZN(n2809) );
  NAND2_X1 U35760 ( .A1(n2822), .A2(n2809), .ZN(n3671) );
  OR2_X1 U35770 ( .A1(n2767), .A2(n3671), .ZN(n2811) );
  OR2_X1 U35780 ( .A1(n2137), .A2(n4864), .ZN(n2810) );
  OR2_X1 U35790 ( .A1(n3400), .A2(n2681), .ZN(n2814) );
  OAI21_X1 U35800 ( .B1(n3182), .B2(n3037), .A(n2814), .ZN(n2815) );
  XNOR2_X1 U35810 ( .A(n2815), .B(n3038), .ZN(n2816) );
  OAI22_X1 U3582 ( .A1(n3040), .A2(n3400), .B1(n3182), .B2(n2681), .ZN(n2817)
         );
  AND2_X1 U3583 ( .A1(n2816), .A2(n2817), .ZN(n3500) );
  INV_X1 U3584 ( .A(n2816), .ZN(n2819) );
  INV_X1 U3585 ( .A(n2817), .ZN(n2818) );
  NAND2_X1 U3586 ( .A1(n2819), .A2(n2818), .ZN(n3499) );
  NAND2_X1 U3587 ( .A1(n2822), .A2(n2821), .ZN(n2823) );
  NAND2_X1 U3588 ( .A1(n2834), .A2(n2823), .ZN(n3702) );
  OR2_X1 U3589 ( .A1(n3702), .A2(n2767), .ZN(n2827) );
  NAND2_X1 U3590 ( .A1(n3029), .A2(REG0_REG_13__SCAN_IN), .ZN(n2826) );
  NAND2_X1 U3591 ( .A1(n2739), .A2(REG2_REG_13__SCAN_IN), .ZN(n2825) );
  OR2_X1 U3592 ( .A1(n2137), .A2(n3779), .ZN(n2824) );
  INV_X1 U3593 ( .A(n3037), .ZN(n2839) );
  MUX2_X1 U3594 ( .A(DATAI_13_), .B(n2828), .S(n2134), .Z(n3688) );
  NAND2_X1 U3595 ( .A1(n2839), .A2(n3688), .ZN(n2829) );
  OAI21_X1 U3596 ( .B1(n3689), .B2(n2830), .A(n2829), .ZN(n2831) );
  NAND2_X1 U3597 ( .A1(n2838), .A2(n3688), .ZN(n2832) );
  OAI21_X1 U3598 ( .B1(n3040), .B2(n3689), .A(n2832), .ZN(n3551) );
  NAND2_X1 U3599 ( .A1(n2834), .A2(n2833), .ZN(n2835) );
  NAND2_X1 U3600 ( .A1(n2846), .A2(n2835), .ZN(n3867) );
  AOI22_X1 U3601 ( .A1(n3029), .A2(REG0_REG_14__SCAN_IN), .B1(n2739), .B2(
        REG2_REG_14__SCAN_IN), .ZN(n2837) );
  OR2_X1 U3602 ( .A1(n2137), .A2(n4884), .ZN(n2836) );
  OAI211_X1 U3603 ( .C1(n3867), .C2(n2767), .A(n2837), .B(n2836), .ZN(n3815)
         );
  NAND2_X1 U3604 ( .A1(n3815), .A2(n2838), .ZN(n2841) );
  MUX2_X1 U3605 ( .A(DATAI_14_), .B(n4890), .S(n2134), .Z(n3870) );
  NAND2_X1 U3606 ( .A1(n2839), .A2(n3870), .ZN(n2840) );
  NAND2_X1 U3607 ( .A1(n2841), .A2(n2840), .ZN(n2842) );
  XNOR2_X1 U3608 ( .A(n2842), .B(n3038), .ZN(n2865) );
  INV_X1 U3609 ( .A(n3815), .ZN(n3722) );
  INV_X1 U3610 ( .A(n3870), .ZN(n3145) );
  OAI22_X1 U3611 ( .A1(n3722), .A2(n3040), .B1(n3089), .B2(n3145), .ZN(n2864)
         );
  AND2_X1 U3612 ( .A1(n2865), .A2(n2864), .ZN(n3863) );
  NAND2_X1 U3613 ( .A1(n2844), .A2(n2843), .ZN(n3808) );
  INV_X1 U3614 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3979) );
  NAND2_X1 U3615 ( .A1(n2846), .A2(n2845), .ZN(n2847) );
  NAND2_X1 U3616 ( .A1(n2157), .A2(n2847), .ZN(n3818) );
  OR2_X1 U3617 ( .A1(n3818), .A2(n2767), .ZN(n2849) );
  AOI22_X1 U3618 ( .A1(n3029), .A2(REG0_REG_15__SCAN_IN), .B1(n2739), .B2(
        REG2_REG_15__SCAN_IN), .ZN(n2848) );
  OAI211_X1 U3619 ( .C1(n2137), .C2(n3979), .A(n2849), .B(n2848), .ZN(n4443)
         );
  NAND2_X1 U3620 ( .A1(n3009), .A2(n4443), .ZN(n2851) );
  MUX2_X1 U3621 ( .A(DATAI_15_), .B(n4907), .S(n2134), .Z(n3821) );
  INV_X1 U3622 ( .A(n3821), .ZN(n3721) );
  OR2_X1 U3623 ( .A1(n3089), .A2(n3721), .ZN(n2850) );
  NAND2_X1 U3624 ( .A1(n2851), .A2(n2850), .ZN(n2867) );
  NAND2_X1 U3625 ( .A1(n4443), .A2(n2852), .ZN(n2854) );
  OR2_X1 U3626 ( .A1(n3037), .A2(n3721), .ZN(n2853) );
  NAND2_X1 U3627 ( .A1(n2854), .A2(n2853), .ZN(n2855) );
  XNOR2_X1 U3628 ( .A(n2855), .B(n3038), .ZN(n3811) );
  NAND2_X1 U3629 ( .A1(n2157), .A2(n2286), .ZN(n2856) );
  NAND2_X1 U3630 ( .A1(n2876), .A2(n2856), .ZN(n4212) );
  OR2_X1 U3631 ( .A1(n4212), .A2(n2767), .ZN(n2861) );
  INV_X1 U3632 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4473) );
  NAND2_X1 U3633 ( .A1(n2739), .A2(REG2_REG_16__SCAN_IN), .ZN(n2858) );
  NAND2_X1 U3634 ( .A1(n3029), .A2(REG0_REG_16__SCAN_IN), .ZN(n2857) );
  OAI211_X1 U3635 ( .C1(n4473), .C2(n2137), .A(n2858), .B(n2857), .ZN(n2859)
         );
  INV_X1 U3636 ( .A(n2859), .ZN(n2860) );
  MUX2_X1 U3637 ( .A(DATAI_16_), .B(n4830), .S(n2134), .Z(n4215) );
  OAI22_X1 U3638 ( .A1(n3817), .A2(n2681), .B1(n3037), .B2(n3750), .ZN(n2862)
         );
  XNOR2_X1 U3639 ( .A(n2862), .B(n3006), .ZN(n2868) );
  NOR2_X1 U3640 ( .A1(n3089), .A2(n3750), .ZN(n2863) );
  AOI21_X1 U3641 ( .B1(n3724), .B2(n3009), .A(n2863), .ZN(n2869) );
  NAND2_X1 U3642 ( .A1(n2868), .A2(n2869), .ZN(n4204) );
  OR2_X1 U3643 ( .A1(n2865), .A2(n2864), .ZN(n3809) );
  OAI211_X1 U3644 ( .C1(n2867), .C2(n3811), .A(n4204), .B(n3809), .ZN(n2866)
         );
  INV_X1 U3645 ( .A(n2867), .ZN(n4207) );
  INV_X1 U3646 ( .A(n3811), .ZN(n2872) );
  INV_X1 U3647 ( .A(n2868), .ZN(n2871) );
  INV_X1 U3648 ( .A(n2869), .ZN(n2870) );
  NAND2_X1 U3649 ( .A1(n2871), .A2(n2870), .ZN(n4203) );
  OAI21_X1 U3650 ( .B1(n4207), .B2(n2872), .A(n4203), .ZN(n2873) );
  AOI21_X2 U3651 ( .B1(n3808), .B2(n2875), .A(n2874), .ZN(n3731) );
  NAND2_X1 U3652 ( .A1(n2876), .A2(n3734), .ZN(n2877) );
  AND2_X1 U3653 ( .A1(n2888), .A2(n2877), .ZN(n3826) );
  NAND2_X1 U3654 ( .A1(n3826), .A2(n2645), .ZN(n2882) );
  NAND2_X1 U3655 ( .A1(n3029), .A2(REG0_REG_17__SCAN_IN), .ZN(n2879) );
  INV_X1 U3656 ( .A(REG2_REG_17__SCAN_IN), .ZN(n3828) );
  OR2_X1 U3657 ( .A1(n3033), .A2(n3828), .ZN(n2878) );
  OAI211_X1 U3658 ( .C1(n3798), .C2(n2137), .A(n2879), .B(n2878), .ZN(n2880)
         );
  INV_X1 U3659 ( .A(n2880), .ZN(n2881) );
  INV_X1 U3660 ( .A(DATAI_17_), .ZN(n2883) );
  MUX2_X1 U3661 ( .A(n2883), .B(n4976), .S(n2134), .Z(n3790) );
  OAI22_X1 U3662 ( .A1(n3747), .A2(n3089), .B1(n3037), .B2(n3790), .ZN(n2884)
         );
  XNOR2_X1 U3663 ( .A(n2884), .B(n3038), .ZN(n2886) );
  OAI22_X1 U3664 ( .A1(n3747), .A2(n3040), .B1(n3089), .B2(n3790), .ZN(n2885)
         );
  NAND2_X1 U3665 ( .A1(n2886), .A2(n2885), .ZN(n3732) );
  NAND2_X1 U3666 ( .A1(n2888), .A2(n2297), .ZN(n2889) );
  NAND2_X1 U3667 ( .A1(n2900), .A2(n2889), .ZN(n4263) );
  OR2_X1 U3668 ( .A1(n4263), .A2(n2767), .ZN(n2894) );
  INV_X1 U3669 ( .A(REG0_REG_18__SCAN_IN), .ZN(n4053) );
  NAND2_X1 U3670 ( .A1(n3028), .A2(REG1_REG_18__SCAN_IN), .ZN(n2891) );
  NAND2_X1 U3671 ( .A1(n2739), .A2(REG2_REG_18__SCAN_IN), .ZN(n2890) );
  OAI211_X1 U3672 ( .C1(n3308), .C2(n4053), .A(n2891), .B(n2890), .ZN(n2892)
         );
  INV_X1 U3673 ( .A(n2892), .ZN(n2893) );
  INV_X1 U3674 ( .A(DATAI_18_), .ZN(n2896) );
  MUX2_X1 U3675 ( .A(n2896), .B(n2895), .S(n2134), .Z(n3767) );
  OAI22_X1 U3676 ( .A1(n3900), .A2(n3089), .B1(n3037), .B2(n3767), .ZN(n2897)
         );
  XNOR2_X1 U3677 ( .A(n2897), .B(n3038), .ZN(n2899) );
  OAI22_X1 U3678 ( .A1(n3900), .A2(n2680), .B1(n3089), .B2(n3767), .ZN(n2898)
         );
  AND2_X1 U3679 ( .A1(n2899), .A2(n2898), .ZN(n4256) );
  NAND2_X1 U3680 ( .A1(n2900), .A2(n4092), .ZN(n2901) );
  AND2_X1 U3681 ( .A1(n2161), .A2(n2901), .ZN(n3893) );
  NAND2_X1 U3682 ( .A1(n3893), .A2(n2645), .ZN(n2906) );
  INV_X1 U3683 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4818) );
  NAND2_X1 U3684 ( .A1(n2739), .A2(REG2_REG_19__SCAN_IN), .ZN(n2903) );
  NAND2_X1 U3685 ( .A1(n3028), .A2(REG1_REG_19__SCAN_IN), .ZN(n2902) );
  OAI211_X1 U3686 ( .C1(n3308), .C2(n4818), .A(n2903), .B(n2902), .ZN(n2904)
         );
  INV_X1 U3687 ( .A(n2904), .ZN(n2905) );
  INV_X1 U3688 ( .A(DATAI_19_), .ZN(n2907) );
  MUX2_X1 U3689 ( .A(n2907), .B(n4433), .S(n2134), .Z(n3844) );
  OAI22_X1 U3690 ( .A1(n4262), .A2(n3040), .B1(n3089), .B2(n3844), .ZN(n2910)
         );
  OAI22_X1 U3691 ( .A1(n4262), .A2(n3089), .B1(n3037), .B2(n3844), .ZN(n2908)
         );
  XNOR2_X1 U3692 ( .A(n2908), .B(n3038), .ZN(n2909) );
  XOR2_X1 U3693 ( .A(n2910), .B(n2909), .Z(n3896) );
  INV_X1 U3694 ( .A(REG3_REG_20__SCAN_IN), .ZN(n2913) );
  NAND2_X1 U3695 ( .A1(n2161), .A2(n2913), .ZN(n2914) );
  NAND2_X1 U3696 ( .A1(n2928), .A2(n2914), .ZN(n4668) );
  INV_X1 U3697 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4669) );
  NAND2_X1 U3698 ( .A1(n3028), .A2(REG1_REG_20__SCAN_IN), .ZN(n2916) );
  NAND2_X1 U3699 ( .A1(n3029), .A2(REG0_REG_20__SCAN_IN), .ZN(n2915) );
  OAI211_X1 U3700 ( .C1(n3033), .C2(n4669), .A(n2916), .B(n2915), .ZN(n2917)
         );
  INV_X1 U3701 ( .A(n2917), .ZN(n2918) );
  NAND2_X1 U3702 ( .A1(n4636), .A2(n2838), .ZN(n2922) );
  INV_X1 U3703 ( .A(DATAI_20_), .ZN(n2920) );
  OR2_X1 U3704 ( .A1(n3037), .A2(n3200), .ZN(n2921) );
  NAND2_X1 U3705 ( .A1(n2922), .A2(n2921), .ZN(n2923) );
  XNOR2_X1 U3706 ( .A(n2923), .B(n3006), .ZN(n2926) );
  NOR2_X1 U3707 ( .A1(n3089), .A2(n3200), .ZN(n2924) );
  AOI21_X1 U3708 ( .B1(n4636), .B2(n3009), .A(n2924), .ZN(n2925) );
  OR2_X1 U3709 ( .A1(n2926), .A2(n2925), .ZN(n4235) );
  NAND2_X1 U3710 ( .A1(n4234), .A2(n4235), .ZN(n4233) );
  NAND2_X1 U3711 ( .A1(n2926), .A2(n2925), .ZN(n4237) );
  NAND2_X1 U3712 ( .A1(n2928), .A2(n2927), .ZN(n2929) );
  AND2_X1 U3713 ( .A1(n2943), .A2(n2929), .ZN(n4644) );
  NAND2_X1 U3714 ( .A1(n4644), .A2(n2645), .ZN(n2934) );
  INV_X1 U3715 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4750) );
  NAND2_X1 U3716 ( .A1(n2739), .A2(REG2_REG_21__SCAN_IN), .ZN(n2931) );
  INV_X1 U3717 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4813) );
  OR2_X1 U3718 ( .A1(n3308), .A2(n4813), .ZN(n2930) );
  OAI211_X1 U3719 ( .C1(n4750), .C2(n2137), .A(n2931), .B(n2930), .ZN(n2932)
         );
  INV_X1 U3720 ( .A(n2932), .ZN(n2933) );
  NAND2_X1 U3721 ( .A1(n4239), .A2(n2838), .ZN(n2936) );
  OR2_X1 U3722 ( .A1(n3037), .A2(n4643), .ZN(n2935) );
  NAND2_X1 U3723 ( .A1(n2936), .A2(n2935), .ZN(n2937) );
  XNOR2_X1 U3724 ( .A(n2937), .B(n3006), .ZN(n3907) );
  NOR2_X1 U3725 ( .A1(n3089), .A2(n4643), .ZN(n2938) );
  AOI21_X1 U3726 ( .B1(n4239), .B2(n3009), .A(n2938), .ZN(n3906) );
  INV_X1 U3727 ( .A(n3907), .ZN(n2940) );
  INV_X1 U3728 ( .A(n3906), .ZN(n2939) );
  INV_X1 U3729 ( .A(REG3_REG_22__SCAN_IN), .ZN(n2942) );
  NAND2_X1 U3730 ( .A1(n2943), .A2(n2942), .ZN(n2944) );
  NAND2_X1 U3731 ( .A1(n2954), .A2(n2944), .ZN(n4627) );
  INV_X1 U3732 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4045) );
  NAND2_X1 U3733 ( .A1(n3028), .A2(REG1_REG_22__SCAN_IN), .ZN(n2946) );
  NAND2_X1 U3734 ( .A1(n2739), .A2(REG2_REG_22__SCAN_IN), .ZN(n2945) );
  OAI211_X1 U3735 ( .C1(n3308), .C2(n4045), .A(n2946), .B(n2945), .ZN(n2947)
         );
  INV_X1 U3736 ( .A(n2947), .ZN(n2948) );
  NAND2_X1 U3737 ( .A1(n4639), .A2(n2838), .ZN(n2951) );
  INV_X1 U3738 ( .A(DATAI_22_), .ZN(n4046) );
  OR2_X1 U3739 ( .A1(n3037), .A2(n4617), .ZN(n2950) );
  NAND2_X1 U3740 ( .A1(n2951), .A2(n2950), .ZN(n2952) );
  XNOR2_X1 U3741 ( .A(n2952), .B(n3038), .ZN(n2965) );
  NOR2_X1 U3742 ( .A1(n3089), .A2(n4617), .ZN(n2953) );
  AOI21_X1 U3743 ( .B1(n4639), .B2(n3009), .A(n2953), .ZN(n2966) );
  XNOR2_X1 U3744 ( .A(n2965), .B(n2966), .ZN(n4246) );
  NAND2_X1 U3745 ( .A1(n2954), .A2(n2300), .ZN(n2955) );
  NAND2_X1 U3746 ( .A1(n2968), .A2(n2955), .ZN(n4609) );
  INV_X1 U3747 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4741) );
  NAND2_X1 U3748 ( .A1(n3029), .A2(REG0_REG_23__SCAN_IN), .ZN(n2957) );
  NAND2_X1 U3749 ( .A1(n2739), .A2(REG2_REG_23__SCAN_IN), .ZN(n2956) );
  OAI211_X1 U3750 ( .C1(n2137), .C2(n4741), .A(n2957), .B(n2956), .ZN(n2958)
         );
  INV_X1 U3751 ( .A(n2958), .ZN(n2959) );
  INV_X1 U3752 ( .A(DATAI_23_), .ZN(n2961) );
  OAI22_X1 U3753 ( .A1(n4581), .A2(n3089), .B1(n3037), .B2(n4600), .ZN(n2962)
         );
  XNOR2_X1 U3754 ( .A(n2962), .B(n3006), .ZN(n3883) );
  OR2_X1 U3755 ( .A1(n4581), .A2(n2680), .ZN(n2964) );
  OR2_X1 U3756 ( .A1(n3089), .A2(n4600), .ZN(n2963) );
  INV_X1 U3757 ( .A(n2965), .ZN(n2967) );
  AND2_X1 U3758 ( .A1(n2967), .A2(n2966), .ZN(n3884) );
  AOI21_X1 U3759 ( .B1(n3883), .B2(n2981), .A(n3884), .ZN(n2980) );
  NAND2_X1 U3760 ( .A1(n2968), .A2(n4226), .ZN(n2969) );
  NAND2_X1 U3761 ( .A1(n2986), .A2(n2969), .ZN(n4587) );
  INV_X1 U3762 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4737) );
  NAND2_X1 U3763 ( .A1(n2739), .A2(REG2_REG_24__SCAN_IN), .ZN(n2971) );
  NAND2_X1 U3764 ( .A1(n3029), .A2(REG0_REG_24__SCAN_IN), .ZN(n2970) );
  OAI211_X1 U3765 ( .C1(n4737), .C2(n2137), .A(n2971), .B(n2970), .ZN(n2972)
         );
  INV_X1 U3766 ( .A(n2972), .ZN(n2973) );
  INV_X1 U3767 ( .A(DATAI_24_), .ZN(n2975) );
  OAI22_X1 U3768 ( .A1(n4564), .A2(n3089), .B1(n3037), .B2(n4589), .ZN(n2976)
         );
  XNOR2_X1 U3769 ( .A(n2976), .B(n3038), .ZN(n4222) );
  INV_X1 U3770 ( .A(n4222), .ZN(n2978) );
  OAI22_X1 U3771 ( .A1(n4564), .A2(n2680), .B1(n3089), .B2(n4589), .ZN(n4224)
         );
  NOR2_X1 U3772 ( .A1(n3883), .A2(n2981), .ZN(n4219) );
  OAI21_X1 U3773 ( .B1(n4219), .B2(n4224), .A(n4222), .ZN(n2984) );
  INV_X1 U3774 ( .A(n3883), .ZN(n2982) );
  INV_X1 U3775 ( .A(n2981), .ZN(n3882) );
  NAND3_X1 U3776 ( .A1(n2982), .A2(n4224), .A3(n3882), .ZN(n2983) );
  NAND2_X1 U3777 ( .A1(n2986), .A2(n4043), .ZN(n2987) );
  NAND2_X1 U3778 ( .A1(n4571), .A2(n2645), .ZN(n2992) );
  INV_X1 U3779 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4733) );
  NAND2_X1 U3780 ( .A1(n3029), .A2(REG0_REG_25__SCAN_IN), .ZN(n2989) );
  NAND2_X1 U3781 ( .A1(n2739), .A2(REG2_REG_25__SCAN_IN), .ZN(n2988) );
  OAI211_X1 U3782 ( .C1(n4733), .C2(n2137), .A(n2989), .B(n2988), .ZN(n2990)
         );
  INV_X1 U3783 ( .A(n2990), .ZN(n2991) );
  INV_X1 U3784 ( .A(DATAI_25_), .ZN(n2993) );
  OAI22_X1 U3785 ( .A1(n4278), .A2(n3089), .B1(n3037), .B2(n4570), .ZN(n2994)
         );
  XNOR2_X1 U3786 ( .A(n2994), .B(n3038), .ZN(n3011) );
  OAI22_X1 U3787 ( .A1(n4278), .A2(n2680), .B1(n3089), .B2(n4570), .ZN(n3010)
         );
  NOR2_X1 U3788 ( .A1(n3011), .A2(n3010), .ZN(n4271) );
  INV_X1 U3789 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4276) );
  NAND2_X1 U3790 ( .A1(n2996), .A2(n4276), .ZN(n2997) );
  NAND2_X1 U3791 ( .A1(n3016), .A2(n2997), .ZN(n4553) );
  INV_X1 U3792 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4729) );
  NAND2_X1 U3793 ( .A1(n3029), .A2(REG0_REG_26__SCAN_IN), .ZN(n2999) );
  NAND2_X1 U3794 ( .A1(n2739), .A2(REG2_REG_26__SCAN_IN), .ZN(n2998) );
  OAI211_X1 U3795 ( .C1(n4729), .C2(n2137), .A(n2999), .B(n2998), .ZN(n3000)
         );
  INV_X1 U3796 ( .A(n3000), .ZN(n3001) );
  NAND2_X1 U3797 ( .A1(n4566), .A2(n2838), .ZN(n3005) );
  INV_X1 U3798 ( .A(DATAI_26_), .ZN(n3003) );
  OR2_X1 U3799 ( .A1(n3037), .A2(n4552), .ZN(n3004) );
  NAND2_X1 U3800 ( .A1(n3005), .A2(n3004), .ZN(n3007) );
  XNOR2_X1 U3801 ( .A(n3007), .B(n3006), .ZN(n3013) );
  NOR2_X1 U3802 ( .A1(n3089), .A2(n4552), .ZN(n3008) );
  AOI21_X1 U3803 ( .B1(n4566), .B2(n3009), .A(n3008), .ZN(n3012) );
  OR2_X1 U3804 ( .A1(n3013), .A2(n3012), .ZN(n4270) );
  NAND2_X1 U3805 ( .A1(n3011), .A2(n3010), .ZN(n4272) );
  NAND2_X1 U3806 ( .A1(n3013), .A2(n3012), .ZN(n4269) );
  NAND2_X1 U3807 ( .A1(n3014), .A2(n4269), .ZN(n3874) );
  INV_X1 U3808 ( .A(n3016), .ZN(n3015) );
  NAND2_X1 U3809 ( .A1(n3015), .A2(REG3_REG_27__SCAN_IN), .ZN(n3026) );
  INV_X1 U3810 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3992) );
  NAND2_X1 U3811 ( .A1(n3016), .A2(n3992), .ZN(n3017) );
  NAND2_X1 U3812 ( .A1(n3026), .A2(n3017), .ZN(n4530) );
  INV_X1 U3813 ( .A(REG1_REG_27__SCAN_IN), .ZN(n3020) );
  NAND2_X1 U3814 ( .A1(n2739), .A2(REG2_REG_27__SCAN_IN), .ZN(n3019) );
  NAND2_X1 U3815 ( .A1(n3029), .A2(REG0_REG_27__SCAN_IN), .ZN(n3018) );
  OAI211_X1 U3816 ( .C1(n3020), .C2(n2137), .A(n3019), .B(n3018), .ZN(n3021)
         );
  INV_X1 U3817 ( .A(n3021), .ZN(n3022) );
  INV_X1 U3818 ( .A(DATAI_27_), .ZN(n3024) );
  OAI22_X1 U3819 ( .A1(n4550), .A2(n3089), .B1(n3037), .B2(n4345), .ZN(n3025)
         );
  XNOR2_X1 U3820 ( .A(n3025), .B(n3038), .ZN(n3044) );
  OAI22_X1 U3821 ( .A1(n4550), .A2(n3040), .B1(n3089), .B2(n4345), .ZN(n3043)
         );
  XNOR2_X1 U3822 ( .A(n3044), .B(n3043), .ZN(n3873) );
  NOR2_X2 U3823 ( .A1(n3874), .A2(n3873), .ZN(n3068) );
  INV_X1 U3824 ( .A(n3068), .ZN(n3067) );
  INV_X1 U3825 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3990) );
  NAND2_X1 U3826 ( .A1(n3026), .A2(n3990), .ZN(n3027) );
  INV_X1 U3827 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3032) );
  NAND2_X1 U3828 ( .A1(n3028), .A2(REG1_REG_28__SCAN_IN), .ZN(n3031) );
  NAND2_X1 U3829 ( .A1(n3029), .A2(REG0_REG_28__SCAN_IN), .ZN(n3030) );
  OAI211_X1 U3830 ( .C1(n3033), .C2(n3032), .A(n3031), .B(n3030), .ZN(n3034)
         );
  INV_X1 U3831 ( .A(n3034), .ZN(n3035) );
  INV_X1 U3832 ( .A(DATAI_28_), .ZN(n3036) );
  OAI22_X1 U3833 ( .A1(n4538), .A2(n3089), .B1(n3037), .B2(n3216), .ZN(n3039)
         );
  XNOR2_X1 U3834 ( .A(n3039), .B(n3038), .ZN(n3042) );
  OAI22_X1 U3835 ( .A1(n4538), .A2(n3040), .B1(n3089), .B2(n3216), .ZN(n3041)
         );
  XNOR2_X1 U3836 ( .A(n3042), .B(n3041), .ZN(n3071) );
  INV_X1 U3837 ( .A(n3071), .ZN(n3066) );
  NAND2_X1 U3838 ( .A1(n3044), .A2(n3043), .ZN(n3069) );
  INV_X1 U3839 ( .A(n3047), .ZN(n3248) );
  NOR2_X1 U3840 ( .A1(n3047), .A2(n3045), .ZN(n3046) );
  MUX2_X1 U3841 ( .A(n3047), .B(n3046), .S(B_REG_SCAN_IN), .Z(n3049) );
  INV_X1 U3842 ( .A(D_REG_1__SCAN_IN), .ZN(n3247) );
  NOR2_X1 U3843 ( .A1(n3045), .A2(n3244), .ZN(n3050) );
  INV_X1 U3844 ( .A(D_REG_27__SCAN_IN), .ZN(n4962) );
  INV_X1 U3845 ( .A(D_REG_21__SCAN_IN), .ZN(n4966) );
  INV_X1 U3846 ( .A(D_REG_23__SCAN_IN), .ZN(n4965) );
  INV_X1 U3847 ( .A(D_REG_25__SCAN_IN), .ZN(n4964) );
  NAND4_X1 U3848 ( .A1(n4962), .A2(n4966), .A3(n4965), .A4(n4964), .ZN(n3051)
         );
  NOR4_X1 U3849 ( .A1(D_REG_9__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(n3051), .ZN(n3933) );
  NOR4_X1 U3850 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_14__SCAN_IN), .ZN(n3052) );
  INV_X1 U3851 ( .A(D_REG_5__SCAN_IN), .ZN(n4971) );
  INV_X1 U3852 ( .A(D_REG_26__SCAN_IN), .ZN(n4963) );
  NAND3_X1 U3853 ( .A1(n3052), .A2(n4971), .A3(n4963), .ZN(n3058) );
  NOR4_X1 U3854 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_12__SCAN_IN), .ZN(n3056) );
  NOR4_X1 U3855 ( .A1(D_REG_13__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n3055) );
  NOR4_X1 U3856 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_22__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n3054) );
  NOR4_X1 U3857 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(D_REG_18__SCAN_IN), .ZN(n3053) );
  NAND4_X1 U3858 ( .A1(n3056), .A2(n3055), .A3(n3054), .A4(n3053), .ZN(n3057)
         );
  NOR3_X1 U3859 ( .A1(D_REG_29__SCAN_IN), .A2(n3058), .A3(n3057), .ZN(n3059)
         );
  NAND2_X1 U3860 ( .A1(n3933), .A2(n3059), .ZN(n3060) );
  NAND2_X1 U3861 ( .A1(n3243), .A2(n3060), .ZN(n3107) );
  NAND2_X1 U3862 ( .A1(n3417), .A2(n3107), .ZN(n3062) );
  INV_X1 U3863 ( .A(n3243), .ZN(n3061) );
  OR2_X1 U3864 ( .A1(n4829), .A2(n4828), .ZN(n4946) );
  NAND2_X1 U3865 ( .A1(n3080), .A2(n4433), .ZN(n3076) );
  AOI21_X1 U3866 ( .B1(n3073), .B2(n3076), .A(n3209), .ZN(n3064) );
  NAND2_X1 U3867 ( .A1(n3067), .A2(n2423), .ZN(n3098) );
  NAND3_X1 U3868 ( .A1(n3068), .A2(n4247), .A3(n3071), .ZN(n3097) );
  INV_X1 U3869 ( .A(n3069), .ZN(n3070) );
  NAND3_X1 U3870 ( .A1(n3071), .A2(n4247), .A3(n3070), .ZN(n3096) );
  NOR2_X1 U3871 ( .A1(n4946), .A2(n4433), .ZN(n3074) );
  NAND2_X1 U3872 ( .A1(n3074), .A2(n4682), .ZN(n3075) );
  NAND2_X1 U3873 ( .A1(n3092), .A2(n3075), .ZN(n3377) );
  INV_X1 U3874 ( .A(n3106), .ZN(n3077) );
  NAND4_X1 U3875 ( .A1(n3377), .A2(n3226), .A3(n3078), .A4(n3077), .ZN(n3079)
         );
  NAND2_X1 U3876 ( .A1(n3079), .A2(STATE_REG_SCAN_IN), .ZN(n4279) );
  INV_X1 U3877 ( .A(n4279), .ZN(n3920) );
  INV_X1 U3878 ( .A(n3242), .ZN(n3081) );
  INV_X1 U3879 ( .A(n4433), .ZN(n3414) );
  NAND2_X1 U3880 ( .A1(n3080), .A2(n3414), .ZN(n4953) );
  OAI22_X1 U3881 ( .A1(n3923), .A2(n3216), .B1(STATE_REG_SCAN_IN), .B2(n3990), 
        .ZN(n3094) );
  INV_X1 U3882 ( .A(n4513), .ZN(n3086) );
  INV_X1 U3883 ( .A(REG1_REG_29__SCAN_IN), .ZN(n4007) );
  NAND2_X1 U3884 ( .A1(n2739), .A2(REG2_REG_29__SCAN_IN), .ZN(n3084) );
  INV_X1 U3885 ( .A(REG0_REG_29__SCAN_IN), .ZN(n4039) );
  OR2_X1 U3886 ( .A1(n3308), .A2(n4039), .ZN(n3083) );
  OAI211_X1 U3887 ( .C1(n4007), .C2(n2137), .A(n3084), .B(n3083), .ZN(n3085)
         );
  NAND2_X1 U3888 ( .A1(n4975), .A2(n3087), .ZN(n3088) );
  NAND2_X1 U3889 ( .A1(n4436), .A2(n4838), .ZN(n3090) );
  INV_X1 U3890 ( .A(n4838), .ZN(n3340) );
  NAND2_X1 U3891 ( .A1(n4436), .A2(n3340), .ZN(n3091) );
  OAI22_X1 U3892 ( .A1(n4355), .A2(n4280), .B1(n4550), .B2(n4277), .ZN(n3093)
         );
  AOI211_X1 U3893 ( .C1(n4521), .C2(n3920), .A(n3094), .B(n3093), .ZN(n3095)
         );
  NAND3_X1 U3894 ( .A1(n3098), .A2(n3097), .A3(n2425), .ZN(U3217) );
  NAND2_X1 U3895 ( .A1(n3412), .A2(n3167), .ZN(n3516) );
  NAND2_X1 U3896 ( .A1(n4642), .A2(n4643), .ZN(n4625) );
  INV_X1 U3897 ( .A(DATAI_29_), .ZN(n3102) );
  OR2_X1 U3898 ( .A1(n2134), .A2(n3102), .ZN(n4354) );
  INV_X1 U3899 ( .A(DATAI_30_), .ZN(n3103) );
  OR2_X1 U3900 ( .A1(n2134), .A2(n3103), .ZN(n4483) );
  NAND2_X1 U3901 ( .A1(n4498), .A2(n4483), .ZN(n4485) );
  INV_X1 U3902 ( .A(DATAI_31_), .ZN(n3104) );
  OR2_X1 U3903 ( .A1(n2134), .A2(n3104), .ZN(n4430) );
  XNOR2_X1 U3904 ( .A(n4485), .B(n3105), .ZN(n4788) );
  NAND2_X1 U3905 ( .A1(n3107), .A2(n2426), .ZN(n3415) );
  NOR2_X4 U3906 ( .A1(n3214), .A2(n3416), .ZN(n5030) );
  INV_X1 U3907 ( .A(B_REG_SCAN_IN), .ZN(n4174) );
  NOR2_X1 U3908 ( .A1(n3339), .A2(n4174), .ZN(n3110) );
  NOR2_X1 U3909 ( .A1(n4952), .A2(n3110), .ZN(n4508) );
  INV_X1 U3910 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4148) );
  NAND2_X1 U3911 ( .A1(n2739), .A2(REG2_REG_31__SCAN_IN), .ZN(n3112) );
  INV_X1 U3912 ( .A(REG0_REG_31__SCAN_IN), .ZN(n4784) );
  OR2_X1 U3913 ( .A1(n3308), .A2(n4784), .ZN(n3111) );
  OAI211_X1 U3914 ( .C1(n2137), .C2(n4148), .A(n3112), .B(n3111), .ZN(n4441)
         );
  NAND2_X1 U3915 ( .A1(n4508), .A2(n4441), .ZN(n4489) );
  NAND2_X1 U3916 ( .A1(n4937), .A2(n3105), .ZN(n3113) );
  NAND2_X1 U3917 ( .A1(n4489), .A2(n3113), .ZN(n4786) );
  AND2_X1 U3918 ( .A1(n4936), .A2(n4942), .ZN(n4928) );
  NAND2_X1 U3919 ( .A1(n4929), .A2(n4928), .ZN(n4927) );
  NAND2_X1 U3920 ( .A1(n3117), .A2(n3115), .ZN(n3118) );
  OR2_X1 U3921 ( .A1(n3119), .A2(n3390), .ZN(n4296) );
  NAND2_X1 U3922 ( .A1(n3119), .A2(n3390), .ZN(n4298) );
  OR2_X1 U3923 ( .A1(n3119), .A2(n4710), .ZN(n3120) );
  OR2_X1 U3924 ( .A1(n4445), .A2(n3413), .ZN(n4302) );
  NAND2_X1 U3925 ( .A1(n4445), .A2(n3413), .ZN(n4305) );
  NAND2_X1 U3926 ( .A1(n4302), .A2(n4305), .ZN(n4372) );
  INV_X1 U3927 ( .A(n3413), .ZN(n3453) );
  NAND2_X1 U3928 ( .A1(n4445), .A2(n3453), .ZN(n3122) );
  NAND2_X1 U3929 ( .A1(n3123), .A2(n3122), .ZN(n3598) );
  AND2_X1 U3930 ( .A1(n3349), .A2(n3606), .ZN(n3124) );
  OAI22_X1 U3931 ( .A1(n3598), .A2(n3124), .B1(n3606), .B2(n3349), .ZN(n3509)
         );
  NOR2_X1 U3932 ( .A1(n2135), .A2(n3517), .ZN(n3479) );
  NAND2_X1 U3933 ( .A1(n4680), .A2(n3634), .ZN(n3136) );
  INV_X1 U3934 ( .A(n3136), .ZN(n3134) );
  NOR2_X1 U3935 ( .A1(n4680), .A2(n3634), .ZN(n3130) );
  OR2_X1 U3936 ( .A1(n3629), .A2(n3535), .ZN(n3129) );
  INV_X1 U3937 ( .A(n3129), .ZN(n3128) );
  AND2_X1 U3938 ( .A1(n3629), .A2(n3535), .ZN(n3126) );
  NAND2_X1 U3939 ( .A1(n3511), .A2(n3490), .ZN(n3524) );
  INV_X1 U3940 ( .A(n3524), .ZN(n3125) );
  NOR2_X1 U3941 ( .A1(n3126), .A2(n3125), .ZN(n3127) );
  OR2_X1 U3942 ( .A1(n3128), .A2(n3127), .ZN(n3621) );
  NAND2_X1 U3943 ( .A1(n3511), .A2(n3485), .ZN(n4311) );
  NAND2_X1 U3944 ( .A1(n3170), .A2(n4311), .ZN(n4373) );
  AND2_X1 U3945 ( .A1(n4373), .A2(n3129), .ZN(n3619) );
  INV_X1 U3946 ( .A(n3130), .ZN(n3131) );
  NAND2_X1 U3947 ( .A1(n3619), .A2(n3131), .ZN(n3132) );
  NAND2_X1 U3948 ( .A1(n3135), .A2(n3132), .ZN(n3133) );
  NOR2_X1 U3949 ( .A1(n3134), .A2(n3133), .ZN(n3139) );
  NAND2_X1 U3950 ( .A1(n2135), .A2(n3517), .ZN(n3480) );
  AND2_X1 U3951 ( .A1(n3480), .A2(n3135), .ZN(n3137) );
  AND2_X1 U3952 ( .A1(n3137), .A2(n3136), .ZN(n3138) );
  OR2_X1 U3953 ( .A1(n4679), .A2(n3579), .ZN(n3660) );
  NAND2_X1 U3954 ( .A1(n4679), .A2(n3579), .ZN(n3662) );
  NAND2_X1 U3955 ( .A1(n3660), .A2(n3662), .ZN(n4379) );
  NAND2_X1 U3956 ( .A1(n3858), .A2(n3579), .ZN(n3141) );
  AND2_X1 U3957 ( .A1(n3182), .A2(n3400), .ZN(n3143) );
  OR2_X1 U3958 ( .A1(n3182), .A2(n3400), .ZN(n3142) );
  NAND2_X1 U3959 ( .A1(n3700), .A2(n3689), .ZN(n3144) );
  NAND2_X1 U3960 ( .A1(n4443), .A2(n3821), .ZN(n3742) );
  OR2_X1 U3961 ( .A1(n3815), .A2(n3145), .ZN(n4329) );
  NAND2_X1 U3962 ( .A1(n3815), .A2(n3145), .ZN(n4315) );
  NAND2_X1 U3963 ( .A1(n4329), .A2(n4315), .ZN(n3190) );
  NOR2_X1 U3964 ( .A1(n3815), .A2(n3870), .ZN(n3716) );
  NAND2_X1 U3965 ( .A1(n3742), .A2(n3716), .ZN(n3147) );
  INV_X1 U3966 ( .A(n4443), .ZN(n4211) );
  NAND2_X1 U3967 ( .A1(n4211), .A2(n3721), .ZN(n3146) );
  AND2_X1 U3968 ( .A1(n3147), .A2(n3146), .ZN(n3740) );
  NAND2_X1 U3969 ( .A1(n3817), .A2(n4215), .ZN(n4407) );
  NAND2_X1 U3970 ( .A1(n3724), .A2(n3750), .ZN(n4404) );
  NAND2_X1 U3971 ( .A1(n4407), .A2(n4404), .ZN(n4378) );
  NAND2_X1 U3972 ( .A1(n3724), .A2(n4215), .ZN(n3148) );
  NAND2_X1 U3973 ( .A1(n3747), .A2(n3790), .ZN(n3150) );
  INV_X1 U3974 ( .A(n3790), .ZN(n3197) );
  NAND2_X1 U3975 ( .A1(n4262), .A2(n3844), .ZN(n4660) );
  NAND2_X1 U3976 ( .A1(n3900), .A2(n3767), .ZN(n3834) );
  NAND2_X1 U3977 ( .A1(n4660), .A2(n3834), .ZN(n3151) );
  INV_X1 U3978 ( .A(n3767), .ZN(n4266) );
  NAND2_X1 U3979 ( .A1(n3900), .A2(n4266), .ZN(n3836) );
  NAND2_X1 U3980 ( .A1(n3792), .A2(n3767), .ZN(n3837) );
  NAND2_X1 U3981 ( .A1(n3836), .A2(n3837), .ZN(n3761) );
  NAND2_X1 U3982 ( .A1(n4655), .A2(n3902), .ZN(n4658) );
  INV_X1 U3983 ( .A(n3200), .ZN(n4667) );
  NAND2_X1 U3984 ( .A1(n4636), .A2(n4667), .ZN(n4364) );
  OAI211_X1 U3985 ( .C1(n3151), .C2(n3761), .A(n4658), .B(n4364), .ZN(n3152)
         );
  INV_X1 U3986 ( .A(n4636), .ZN(n3913) );
  NAND2_X1 U3987 ( .A1(n3913), .A2(n3200), .ZN(n4365) );
  INV_X1 U3988 ( .A(n4643), .ZN(n3910) );
  NAND2_X1 U3989 ( .A1(n4239), .A2(n3910), .ZN(n3154) );
  NAND2_X1 U3990 ( .A1(n4639), .A2(n4617), .ZN(n3203) );
  NAND2_X1 U3991 ( .A1(n4596), .A2(n3203), .ZN(n4620) );
  INV_X1 U3992 ( .A(n4639), .ZN(n4601) );
  INV_X1 U3993 ( .A(n4617), .ZN(n3155) );
  INV_X1 U3994 ( .A(n4570), .ZN(n3205) );
  NAND2_X1 U3995 ( .A1(n4583), .A2(n3205), .ZN(n3160) );
  NAND2_X1 U3996 ( .A1(n4566), .A2(n4547), .ZN(n4356) );
  NOR2_X1 U3997 ( .A1(n4566), .A2(n4547), .ZN(n4358) );
  NAND2_X1 U3998 ( .A1(n4550), .A2(n4345), .ZN(n3162) );
  INV_X1 U3999 ( .A(n3216), .ZN(n4495) );
  NAND2_X1 U4000 ( .A1(n4538), .A2(n4495), .ZN(n4500) );
  NAND2_X1 U4001 ( .A1(n4500), .A2(n4502), .ZN(n4353) );
  XNOR2_X1 U4002 ( .A(n4494), .B(n4353), .ZN(n4520) );
  XNOR2_X1 U4003 ( .A(n3422), .B(n4828), .ZN(n3163) );
  NAND2_X1 U4004 ( .A1(n3163), .A2(n4433), .ZN(n4699) );
  INV_X1 U4005 ( .A(n4293), .ZN(n4932) );
  NAND2_X1 U4006 ( .A1(n4931), .A2(n3164), .ZN(n3165) );
  INV_X1 U4007 ( .A(n4703), .ZN(n4368) );
  NAND2_X1 U4008 ( .A1(n3165), .A2(n4368), .ZN(n3560) );
  NAND2_X1 U4009 ( .A1(n3560), .A2(n4296), .ZN(n3166) );
  XNOR2_X1 U4010 ( .A(n4446), .B(n4300), .ZN(n4390) );
  OR2_X1 U4011 ( .A1(n4446), .A2(n3559), .ZN(n4301) );
  AND2_X1 U4012 ( .A1(n3349), .A2(n3167), .ZN(n3599) );
  OR2_X1 U4013 ( .A1(n3349), .A2(n3167), .ZN(n4317) );
  NAND2_X1 U4014 ( .A1(n2135), .A2(n2723), .ZN(n4318) );
  NAND2_X1 U4015 ( .A1(n3510), .A2(n4318), .ZN(n3169) );
  OR2_X1 U4016 ( .A1(n2135), .A2(n2723), .ZN(n4307) );
  AND2_X1 U4017 ( .A1(n4680), .A2(n3626), .ZN(n4674) );
  NAND2_X1 U4018 ( .A1(n3577), .A2(n4683), .ZN(n4384) );
  INV_X1 U4019 ( .A(n4384), .ZN(n3179) );
  NOR2_X1 U4020 ( .A1(n4674), .A2(n3179), .ZN(n3171) );
  NAND2_X1 U4021 ( .A1(n3629), .A2(n3176), .ZN(n4310) );
  AND2_X1 U4022 ( .A1(n3171), .A2(n4310), .ZN(n3574) );
  NAND2_X1 U4023 ( .A1(n3700), .A2(n4444), .ZN(n3172) );
  NAND2_X1 U4024 ( .A1(n3182), .A2(n3695), .ZN(n3690) );
  NAND2_X1 U4025 ( .A1(n3172), .A2(n3690), .ZN(n3181) );
  INV_X1 U4026 ( .A(n3662), .ZN(n3173) );
  NOR2_X1 U4027 ( .A1(n3181), .A2(n3173), .ZN(n4327) );
  AND2_X1 U4028 ( .A1(n3574), .A2(n4327), .ZN(n3175) );
  AND2_X1 U4029 ( .A1(n4311), .A2(n3175), .ZN(n3174) );
  INV_X1 U4030 ( .A(n3175), .ZN(n3177) );
  OR2_X1 U4031 ( .A1(n3629), .A2(n3176), .ZN(n4312) );
  INV_X1 U4032 ( .A(n4327), .ZN(n3180) );
  OR2_X1 U4033 ( .A1(n4680), .A2(n3626), .ZN(n4676) );
  NAND2_X1 U4034 ( .A1(n3627), .A2(n4689), .ZN(n4385) );
  AND2_X1 U4035 ( .A1(n4676), .A2(n4385), .ZN(n3178) );
  OR2_X1 U4036 ( .A1(n3179), .A2(n3178), .ZN(n3575) );
  OR2_X1 U4037 ( .A1(n3180), .A2(n3575), .ZN(n3186) );
  INV_X1 U4038 ( .A(n3181), .ZN(n3185) );
  OR2_X1 U4039 ( .A1(n3182), .A2(n3695), .ZN(n3692) );
  NAND2_X1 U4040 ( .A1(n3692), .A2(n3660), .ZN(n3184) );
  AND2_X1 U4041 ( .A1(n3689), .A2(n3688), .ZN(n3183) );
  AOI21_X1 U4042 ( .B1(n3185), .B2(n3184), .A(n3183), .ZN(n4332) );
  NAND2_X1 U40430 ( .A1(n3186), .A2(n4332), .ZN(n3187) );
  NAND2_X1 U4044 ( .A1(n3189), .A2(n3188), .ZN(n4403) );
  NAND2_X1 U4045 ( .A1(n4211), .A2(n3821), .ZN(n4330) );
  NAND2_X1 U4046 ( .A1(n4443), .A2(n3721), .ZN(n4316) );
  NAND2_X1 U4047 ( .A1(n4330), .A2(n4316), .ZN(n3719) );
  INV_X1 U4048 ( .A(n4329), .ZN(n3191) );
  NOR2_X1 U4049 ( .A1(n3719), .A2(n3191), .ZN(n3192) );
  NAND2_X1 U4050 ( .A1(n3718), .A2(n3192), .ZN(n3193) );
  NAND2_X1 U4051 ( .A1(n3193), .A2(n4316), .ZN(n3745) );
  INV_X1 U4052 ( .A(n4378), .ZN(n3194) );
  NAND2_X1 U4053 ( .A1(n3745), .A2(n3194), .ZN(n3195) );
  NAND2_X1 U4054 ( .A1(n4655), .A2(n3844), .ZN(n3196) );
  NAND2_X1 U4055 ( .A1(n3196), .A2(n3837), .ZN(n3199) );
  AND2_X1 U4056 ( .A1(n4259), .A2(n3790), .ZN(n3786) );
  OR2_X1 U4057 ( .A1(n3199), .A2(n3786), .ZN(n4406) );
  NAND2_X1 U4058 ( .A1(n3747), .A2(n3197), .ZN(n3787) );
  AND2_X1 U4059 ( .A1(n3836), .A2(n3787), .ZN(n3198) );
  OAI22_X1 U4060 ( .A1(n3199), .A2(n3198), .B1(n4655), .B2(n3844), .ZN(n4651)
         );
  NOR2_X1 U4061 ( .A1(n4636), .A2(n3200), .ZN(n3201) );
  OR2_X1 U4062 ( .A1(n4651), .A2(n3201), .ZN(n4338) );
  NAND2_X1 U4063 ( .A1(n4338), .A2(n2169), .ZN(n4409) );
  NAND2_X1 U4064 ( .A1(n4239), .A2(n4643), .ZN(n4363) );
  NAND2_X1 U4065 ( .A1(n3202), .A2(n4363), .ZN(n4595) );
  NAND2_X1 U4066 ( .A1(n4595), .A2(n4596), .ZN(n3204) );
  NAND2_X1 U4067 ( .A1(n4624), .A2(n4600), .ZN(n4362) );
  AND2_X1 U4068 ( .A1(n4362), .A2(n3203), .ZN(n4290) );
  NAND2_X1 U4069 ( .A1(n3204), .A2(n4290), .ZN(n4578) );
  NAND2_X1 U4070 ( .A1(n4564), .A2(n3158), .ZN(n4361) );
  OR2_X1 U4071 ( .A1(n4624), .A2(n4600), .ZN(n4577) );
  AND2_X1 U4072 ( .A1(n4361), .A2(n4577), .ZN(n4413) );
  AND2_X1 U4073 ( .A1(n4603), .A2(n4589), .ZN(n4360) );
  NAND2_X1 U4074 ( .A1(n4583), .A2(n4570), .ZN(n4359) );
  INV_X1 U4075 ( .A(n4566), .ZN(n3875) );
  NAND2_X1 U4076 ( .A1(n3875), .A2(n4547), .ZN(n3206) );
  NAND2_X1 U4077 ( .A1(n4278), .A2(n3205), .ZN(n4541) );
  NAND2_X1 U4078 ( .A1(n3206), .A2(n4541), .ZN(n4421) );
  NAND2_X1 U4079 ( .A1(n4566), .A2(n4552), .ZN(n4288) );
  NAND2_X1 U4080 ( .A1(n4550), .A2(n4535), .ZN(n4346) );
  XNOR2_X1 U4081 ( .A(n4503), .B(n4353), .ZN(n3212) );
  NAND2_X1 U4082 ( .A1(n3072), .A2(n4829), .ZN(n3208) );
  NAND2_X1 U4083 ( .A1(n4828), .A2(n3414), .ZN(n3207) );
  OAI22_X1 U4084 ( .A1(n4355), .A2(n4952), .B1(n4682), .B2(n3216), .ZN(n3210)
         );
  AOI21_X1 U4085 ( .B1(n4935), .B2(n4442), .A(n3210), .ZN(n3211) );
  OAI21_X1 U4086 ( .B1(n3212), .B2(n4704), .A(n3211), .ZN(n4525) );
  AOI21_X1 U4087 ( .B1(n4520), .B2(n5017), .A(n4525), .ZN(n3225) );
  INV_X1 U4088 ( .A(n3416), .ZN(n3213) );
  OAI21_X1 U4089 ( .B1(n3215), .B2(n3216), .A(n4499), .ZN(n4523) );
  OR2_X1 U4090 ( .A1(n4523), .A2(n4820), .ZN(n3219) );
  INV_X1 U4091 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3217) );
  OR2_X1 U4092 ( .A1(n5020), .A2(n3217), .ZN(n3218) );
  INV_X1 U4093 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3221) );
  OR2_X1 U4094 ( .A1(n5030), .A2(n3221), .ZN(n3222) );
  INV_X1 U4095 ( .A(n4975), .ZN(n3245) );
  MUX2_X1 U4096 ( .A(n2687), .B(n3227), .S(STATE_REG_SCAN_IN), .Z(n3228) );
  INV_X1 U4097 ( .A(n3228), .ZN(U3348) );
  MUX2_X1 U4098 ( .A(n2736), .B(n3285), .S(STATE_REG_SCAN_IN), .Z(n3229) );
  INV_X1 U4099 ( .A(n3229), .ZN(U3345) );
  INV_X1 U4100 ( .A(IR_REG_30__SCAN_IN), .ZN(n4069) );
  NAND2_X1 U4101 ( .A1(IR_REG_31__SCAN_IN), .A2(n4069), .ZN(n3928) );
  OR3_X1 U4102 ( .A1(n3230), .A2(n3928), .A3(U3149), .ZN(n3231) );
  OAI21_X1 U4103 ( .B1(STATE_REG_SCAN_IN), .B2(n3104), .A(n3231), .ZN(U3321)
         );
  NAND2_X1 U4104 ( .A1(n3244), .A2(STATE_REG_SCAN_IN), .ZN(n3232) );
  OAI21_X1 U4105 ( .B1(STATE_REG_SCAN_IN), .B2(n3003), .A(n3232), .ZN(U3326)
         );
  NAND2_X1 U4106 ( .A1(n2629), .A2(STATE_REG_SCAN_IN), .ZN(n3233) );
  OAI21_X1 U4107 ( .B1(STATE_REG_SCAN_IN), .B2(n3103), .A(n3233), .ZN(U3322)
         );
  INV_X1 U4108 ( .A(n3339), .ZN(n3250) );
  NAND2_X1 U4109 ( .A1(n3250), .A2(STATE_REG_SCAN_IN), .ZN(n3234) );
  OAI21_X1 U4110 ( .B1(STATE_REG_SCAN_IN), .B2(n3024), .A(n3234), .ZN(U3325)
         );
  MUX2_X1 U4111 ( .A(n4433), .B(n2907), .S(U3149), .Z(n3235) );
  INV_X1 U4112 ( .A(n3235), .ZN(U3333) );
  NAND2_X1 U4113 ( .A1(n3072), .A2(STATE_REG_SCAN_IN), .ZN(n3236) );
  OAI21_X1 U4114 ( .B1(STATE_REG_SCAN_IN), .B2(n2920), .A(n3236), .ZN(U3332)
         );
  NAND2_X1 U4115 ( .A1(n3045), .A2(STATE_REG_SCAN_IN), .ZN(n3237) );
  OAI21_X1 U4116 ( .B1(STATE_REG_SCAN_IN), .B2(n2993), .A(n3237), .ZN(U3327)
         );
  NAND2_X1 U4117 ( .A1(n3238), .A2(STATE_REG_SCAN_IN), .ZN(n3239) );
  OAI21_X1 U4118 ( .B1(STATE_REG_SCAN_IN), .B2(n2896), .A(n3239), .ZN(U3334)
         );
  MUX2_X1 U4119 ( .A(n3240), .B(n3546), .S(STATE_REG_SCAN_IN), .Z(n3241) );
  INV_X1 U4120 ( .A(n3241), .ZN(U3341) );
  NOR2_X1 U4121 ( .A1(n3245), .A2(n3244), .ZN(n3249) );
  INV_X1 U4122 ( .A(n3045), .ZN(n3246) );
  AOI22_X1 U4123 ( .A1(n4974), .A2(n3247), .B1(n3249), .B2(n3246), .ZN(U3459)
         );
  INV_X1 U4124 ( .A(D_REG_0__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U4125 ( .A1(n4974), .A2(n4175), .B1(n3249), .B2(n3248), .ZN(U3458)
         );
  INV_X1 U4126 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n3257) );
  NAND3_X1 U4127 ( .A1(n4923), .A2(IR_REG_0__SCAN_IN), .A3(n5021), .ZN(n3256)
         );
  INV_X1 U4128 ( .A(REG2_REG_0__SCAN_IN), .ZN(n4957) );
  AOI21_X1 U4129 ( .B1(n3250), .B2(n4957), .A(n4838), .ZN(n3342) );
  OAI21_X1 U4130 ( .B1(n3250), .B2(REG1_REG_0__SCAN_IN), .A(n2378), .ZN(n3252)
         );
  NOR2_X1 U4131 ( .A1(n3342), .A2(IR_REG_0__SCAN_IN), .ZN(n3251) );
  AOI21_X1 U4132 ( .B1(n3342), .B2(n3252), .A(n3251), .ZN(n3253) );
  AOI22_X1 U4133 ( .A1(n3254), .A2(n3253), .B1(REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n3255) );
  OAI211_X1 U4134 ( .C1(n4911), .C2(n3257), .A(n3256), .B(n3255), .ZN(U3240)
         );
  XOR2_X1 U4135 ( .A(n3258), .B(REG1_REG_3__SCAN_IN), .Z(n3261) );
  XOR2_X1 U4136 ( .A(n3259), .B(REG2_REG_3__SCAN_IN), .Z(n3260) );
  AOI22_X1 U4137 ( .A1(n4923), .A2(n3261), .B1(n4921), .B2(n3260), .ZN(n3263)
         );
  INV_X1 U4138 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4186) );
  NOR2_X1 U4139 ( .A1(STATE_REG_SCAN_IN), .A2(n4186), .ZN(n3438) );
  AOI21_X1 U4140 ( .B1(n4914), .B2(ADDR_REG_3__SCAN_IN), .A(n3438), .ZN(n3262)
         );
  OAI211_X1 U4141 ( .C1(n3264), .C2(n4926), .A(n3263), .B(n3262), .ZN(U3243)
         );
  NOR2_X1 U4142 ( .A1(n4914), .A2(U4043), .ZN(U3148) );
  XNOR2_X1 U4143 ( .A(n3265), .B(REG1_REG_6__SCAN_IN), .ZN(n3272) );
  XNOR2_X1 U4144 ( .A(n3266), .B(n3591), .ZN(n3270) );
  INV_X1 U4145 ( .A(n4833), .ZN(n3268) );
  NAND2_X1 U4146 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3350) );
  NAND2_X1 U4147 ( .A1(n4914), .A2(ADDR_REG_6__SCAN_IN), .ZN(n3267) );
  OAI211_X1 U4148 ( .C1(n4926), .C2(n3268), .A(n3350), .B(n3267), .ZN(n3269)
         );
  AOI21_X1 U4149 ( .B1(n3270), .B2(n4921), .A(n3269), .ZN(n3271) );
  OAI21_X1 U4150 ( .B1(n3272), .B2(n4902), .A(n3271), .ZN(U3246) );
  INV_X1 U4151 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n4104) );
  NAND2_X1 U4152 ( .A1(U4043), .A2(n3629), .ZN(n3273) );
  OAI21_X1 U4153 ( .B1(U4043), .B2(n4104), .A(n3273), .ZN(U3558) );
  INV_X1 U4154 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n4106) );
  NAND2_X1 U4155 ( .A1(U4043), .A2(n4936), .ZN(n3274) );
  OAI21_X1 U4156 ( .B1(U4043), .B2(n4106), .A(n3274), .ZN(U3550) );
  AOI211_X1 U4157 ( .C1(n2189), .C2(n3276), .A(n3275), .B(n4896), .ZN(n3284)
         );
  AOI211_X1 U4158 ( .C1(n3279), .C2(n3278), .A(n3277), .B(n4902), .ZN(n3283)
         );
  INV_X1 U4159 ( .A(n4834), .ZN(n3281) );
  AND2_X1 U4160 ( .A1(U3149), .A2(REG3_REG_5__SCAN_IN), .ZN(n3428) );
  AOI21_X1 U4161 ( .B1(n4914), .B2(ADDR_REG_5__SCAN_IN), .A(n3428), .ZN(n3280)
         );
  OAI21_X1 U4162 ( .B1(n4926), .B2(n3281), .A(n3280), .ZN(n3282) );
  OR3_X1 U4163 ( .A1(n3284), .A2(n3283), .A3(n3282), .ZN(U3245) );
  MUX2_X1 U4164 ( .A(REG1_REG_7__SCAN_IN), .B(n2564), .S(n3285), .Z(n3286) );
  INV_X1 U4165 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n3288) );
  AND2_X1 U4166 ( .A1(U3149), .A2(REG3_REG_7__SCAN_IN), .ZN(n3473) );
  INV_X1 U4167 ( .A(n3473), .ZN(n3287) );
  OAI21_X1 U4168 ( .B1(n4911), .B2(n3288), .A(n3287), .ZN(n3293) );
  AOI211_X1 U4169 ( .C1(n3291), .C2(n3290), .A(n4896), .B(n3289), .ZN(n3292)
         );
  AOI211_X1 U4170 ( .C1(n4908), .C2(n3294), .A(n3293), .B(n3292), .ZN(n3295)
         );
  OAI21_X1 U4171 ( .B1(n4902), .B2(n3296), .A(n3295), .ZN(U3247) );
  XNOR2_X1 U4172 ( .A(n3297), .B(n3613), .ZN(n3304) );
  NOR2_X1 U4173 ( .A1(STATE_REG_SCAN_IN), .A2(n3298), .ZN(n3369) );
  NOR2_X1 U4174 ( .A1(n4926), .A2(n2566), .ZN(n3299) );
  AOI211_X1 U4175 ( .C1(n4914), .C2(ADDR_REG_8__SCAN_IN), .A(n3369), .B(n3299), 
        .ZN(n3303) );
  OAI211_X1 U4176 ( .C1(n3301), .C2(REG1_REG_8__SCAN_IN), .A(n3300), .B(n4923), 
        .ZN(n3302) );
  OAI211_X1 U4177 ( .C1(n3304), .C2(n4896), .A(n3303), .B(n3302), .ZN(U3248)
         );
  INV_X1 U4178 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n4118) );
  NAND2_X1 U4179 ( .A1(U4043), .A2(n3695), .ZN(n3305) );
  OAI21_X1 U4180 ( .B1(U4043), .B2(n4118), .A(n3305), .ZN(U3562) );
  INV_X1 U4181 ( .A(DATAO_REG_5__SCAN_IN), .ZN(n4129) );
  NAND2_X1 U4182 ( .A1(U4043), .A2(n3349), .ZN(n3306) );
  OAI21_X1 U4183 ( .B1(U4043), .B2(n4129), .A(n3306), .ZN(U3555) );
  INV_X1 U4184 ( .A(DATAO_REG_14__SCAN_IN), .ZN(n4133) );
  NAND2_X1 U4185 ( .A1(U4043), .A2(n3815), .ZN(n3307) );
  OAI21_X1 U4186 ( .B1(U4043), .B2(n4133), .A(n3307), .ZN(U3564) );
  INV_X1 U4187 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n4134) );
  INV_X1 U4188 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4038) );
  NAND2_X1 U4189 ( .A1(n2739), .A2(REG2_REG_30__SCAN_IN), .ZN(n3310) );
  INV_X1 U4190 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4789) );
  OR2_X1 U4191 ( .A1(n3308), .A2(n4789), .ZN(n3309) );
  OAI211_X1 U4192 ( .C1(n2137), .C2(n4038), .A(n3310), .B(n3309), .ZN(n4507)
         );
  NAND2_X1 U4193 ( .A1(U4043), .A2(n4507), .ZN(n3311) );
  OAI21_X1 U4194 ( .B1(U4043), .B2(n4134), .A(n3311), .ZN(U3580) );
  INV_X1 U4195 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n4137) );
  NAND2_X1 U4196 ( .A1(U4043), .A2(n3577), .ZN(n3312) );
  OAI21_X1 U4197 ( .B1(U4043), .B2(n4137), .A(n3312), .ZN(U3560) );
  INV_X1 U4198 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n4108) );
  NAND2_X1 U4199 ( .A1(U4043), .A2(n4680), .ZN(n3313) );
  OAI21_X1 U4200 ( .B1(U4043), .B2(n4108), .A(n3313), .ZN(U3559) );
  INV_X1 U4201 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n4136) );
  NAND2_X1 U4202 ( .A1(n4259), .A2(U4043), .ZN(n3314) );
  OAI21_X1 U4203 ( .B1(U4043), .B2(n4136), .A(n3314), .ZN(U3567) );
  INV_X1 U4204 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n4145) );
  NAND2_X1 U4205 ( .A1(n4239), .A2(U4043), .ZN(n3315) );
  OAI21_X1 U4206 ( .B1(U4043), .B2(n4145), .A(n3315), .ZN(U3571) );
  INV_X1 U4207 ( .A(DATAO_REG_16__SCAN_IN), .ZN(n4164) );
  NAND2_X1 U4208 ( .A1(n3724), .A2(U4043), .ZN(n3316) );
  OAI21_X1 U4209 ( .B1(U4043), .B2(n4164), .A(n3316), .ZN(U3566) );
  INV_X1 U4210 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n4165) );
  NAND2_X1 U4211 ( .A1(n3792), .A2(U4043), .ZN(n3317) );
  OAI21_X1 U4212 ( .B1(U4043), .B2(n4165), .A(n3317), .ZN(U3568) );
  INV_X1 U4213 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n4109) );
  NAND2_X1 U4214 ( .A1(n4655), .A2(U4043), .ZN(n3318) );
  OAI21_X1 U4215 ( .B1(U4043), .B2(n4109), .A(n3318), .ZN(U3569) );
  INV_X1 U4216 ( .A(DATAO_REG_7__SCAN_IN), .ZN(n4167) );
  NAND2_X1 U4217 ( .A1(U4043), .A2(n3511), .ZN(n3319) );
  OAI21_X1 U4218 ( .B1(U4043), .B2(n4167), .A(n3319), .ZN(U3557) );
  INV_X1 U4219 ( .A(DATAO_REG_6__SCAN_IN), .ZN(n4123) );
  NAND2_X1 U4220 ( .A1(U4043), .A2(n2135), .ZN(n3320) );
  OAI21_X1 U4221 ( .B1(U4043), .B2(n4123), .A(n3320), .ZN(U3556) );
  INV_X1 U4222 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n4103) );
  NAND2_X1 U4223 ( .A1(U4043), .A2(n3119), .ZN(n3321) );
  OAI21_X1 U4224 ( .B1(U4043), .B2(n4103), .A(n3321), .ZN(U3552) );
  INV_X1 U4225 ( .A(DATAO_REG_22__SCAN_IN), .ZN(n4116) );
  NAND2_X1 U4226 ( .A1(n4639), .A2(U4043), .ZN(n3323) );
  OAI21_X1 U4227 ( .B1(U4043), .B2(n4116), .A(n3323), .ZN(U3572) );
  AOI22_X1 U4228 ( .A1(n4914), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3336) );
  MUX2_X1 U4229 ( .A(REG2_REG_2__SCAN_IN), .B(n4708), .S(n2638), .Z(n3325) );
  NAND3_X1 U4230 ( .A1(n3324), .A2(n3326), .A3(n3325), .ZN(n3327) );
  NAND3_X1 U4231 ( .A1(n4921), .A2(n3328), .A3(n3327), .ZN(n3335) );
  NAND3_X1 U4232 ( .A1(n4451), .A2(n3330), .A3(n3329), .ZN(n3331) );
  NAND3_X1 U4233 ( .A1(n4923), .A2(n3332), .A3(n3331), .ZN(n3334) );
  NAND2_X1 U4234 ( .A1(n4908), .A2(n4836), .ZN(n3333) );
  AND4_X1 U4235 ( .A1(n3336), .A2(n3335), .A3(n3334), .A4(n3333), .ZN(n3345)
         );
  XNOR2_X1 U4236 ( .A(n3338), .B(n3337), .ZN(n3437) );
  NAND3_X1 U4237 ( .A1(n3437), .A2(n3340), .A3(n3339), .ZN(n3344) );
  NAND2_X1 U4238 ( .A1(n4435), .A2(REG2_REG_0__SCAN_IN), .ZN(n3341) );
  MUX2_X1 U4239 ( .A(n3342), .B(n3341), .S(IR_REG_0__SCAN_IN), .Z(n3343) );
  NAND3_X1 U4240 ( .A1(n3344), .A2(U4043), .A3(n3343), .ZN(n4851) );
  NAND2_X1 U4241 ( .A1(n3345), .A2(n4851), .ZN(U3242) );
  INV_X1 U4242 ( .A(n3467), .ZN(n3347) );
  NOR2_X1 U4243 ( .A1(n3347), .A2(n3466), .ZN(n3348) );
  XNOR2_X1 U4244 ( .A(n3346), .B(n3348), .ZN(n3355) );
  NAND2_X1 U4245 ( .A1(n4260), .A2(n3349), .ZN(n3351) );
  OAI211_X1 U4246 ( .C1(n3529), .C2(n4280), .A(n3351), .B(n3350), .ZN(n3353)
         );
  NOR2_X1 U4247 ( .A1(n4279), .A2(n3590), .ZN(n3352) );
  AOI211_X1 U4248 ( .C1(n3517), .C2(n4283), .A(n3353), .B(n3352), .ZN(n3354)
         );
  OAI21_X1 U4249 ( .B1(n3355), .B2(n4285), .A(n3354), .ZN(U3236) );
  INV_X1 U4250 ( .A(n3356), .ZN(n3850) );
  NAND2_X1 U4251 ( .A1(n3850), .A2(n3357), .ZN(n3368) );
  OR2_X1 U4252 ( .A1(n3346), .A2(n3358), .ZN(n3363) );
  INV_X1 U4253 ( .A(n3359), .ZN(n3360) );
  OR2_X1 U4254 ( .A1(n3361), .A2(n3360), .ZN(n3362) );
  NAND2_X1 U4255 ( .A1(n3363), .A2(n3362), .ZN(n3364) );
  AOI21_X1 U4256 ( .B1(n3367), .B2(n3365), .A(n3364), .ZN(n3366) );
  AOI21_X1 U4257 ( .B1(n3368), .B2(n3367), .A(n3366), .ZN(n3375) );
  NAND2_X1 U4258 ( .A1(n4260), .A2(n3511), .ZN(n3371) );
  INV_X1 U4259 ( .A(n3369), .ZN(n3370) );
  OAI211_X1 U4260 ( .C1(n3528), .C2(n4280), .A(n3371), .B(n3370), .ZN(n3373)
         );
  NOR2_X1 U4261 ( .A1(n4279), .A2(n3612), .ZN(n3372) );
  AOI211_X1 U4262 ( .C1(n3535), .C2(n4283), .A(n3373), .B(n3372), .ZN(n3374)
         );
  OAI21_X1 U4263 ( .B1(n3375), .B2(n4285), .A(n3374), .ZN(U3218) );
  NAND2_X1 U4264 ( .A1(n3377), .A2(n2426), .ZN(n3434) );
  OAI22_X1 U4265 ( .A1(n3378), .A2(n4277), .B1(n4280), .B2(n4940), .ZN(n3381)
         );
  NOR2_X1 U4266 ( .A1(n3923), .A2(n3379), .ZN(n3380) );
  AOI211_X1 U4267 ( .C1(REG3_REG_1__SCAN_IN), .C2(n3434), .A(n3381), .B(n3380), 
        .ZN(n3382) );
  OAI21_X1 U4268 ( .B1(n3383), .B2(n4285), .A(n3382), .ZN(U3219) );
  NAND2_X1 U4269 ( .A1(n3385), .A2(n3384), .ZN(n3389) );
  INV_X1 U4270 ( .A(n3386), .ZN(n3387) );
  AOI21_X1 U4271 ( .B1(n3389), .B2(n3388), .A(n3387), .ZN(n3394) );
  OAI22_X1 U4272 ( .A1(n3121), .A2(n4280), .B1(n4277), .B2(n3116), .ZN(n3392)
         );
  NOR2_X1 U4273 ( .A1(n3923), .A2(n3390), .ZN(n3391) );
  AOI211_X1 U4274 ( .C1(REG3_REG_2__SCAN_IN), .C2(n3434), .A(n3392), .B(n3391), 
        .ZN(n3393) );
  OAI21_X1 U4275 ( .B1(n3394), .B2(n4285), .A(n3393), .ZN(U3234) );
  XOR2_X1 U4276 ( .A(n3397), .B(n3396), .Z(n3398) );
  XNOR2_X1 U4277 ( .A(n3395), .B(n3398), .ZN(n3404) );
  NAND2_X1 U4278 ( .A1(n4260), .A2(n3577), .ZN(n3399) );
  NAND2_X1 U4279 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n3545) );
  OAI211_X1 U4280 ( .C1(n3400), .C2(n4280), .A(n3399), .B(n3545), .ZN(n3402)
         );
  NOR2_X1 U4281 ( .A1(n4279), .A2(n3584), .ZN(n3401) );
  AOI211_X1 U4282 ( .C1(n3582), .C2(n4283), .A(n3402), .B(n3401), .ZN(n3403)
         );
  OAI21_X1 U4283 ( .B1(n3404), .B2(n4285), .A(n3403), .ZN(U3233) );
  INV_X1 U4284 ( .A(DATAO_REG_24__SCAN_IN), .ZN(n4160) );
  NAND2_X1 U4285 ( .A1(n4603), .A2(U4043), .ZN(n3405) );
  OAI21_X1 U4286 ( .B1(U4043), .B2(n4160), .A(n3405), .ZN(U3574) );
  XNOR2_X1 U4287 ( .A(n3406), .B(n4372), .ZN(n3421) );
  XOR2_X1 U4288 ( .A(n4372), .B(n3407), .Z(n3410) );
  AOI22_X1 U4289 ( .A1(n4446), .A2(n4935), .B1(n3453), .B2(n4937), .ZN(n3408)
         );
  OAI21_X1 U4290 ( .B1(n3513), .B2(n4952), .A(n3408), .ZN(n3409) );
  AOI21_X1 U4291 ( .B1(n3410), .B2(n4949), .A(n3409), .ZN(n3411) );
  OAI21_X1 U4292 ( .B1(n4699), .B2(n3421), .A(n3411), .ZN(n5005) );
  INV_X1 U4293 ( .A(n3412), .ZN(n3605) );
  OAI211_X1 U4294 ( .C1(n3568), .C2(n3413), .A(n3605), .B(n2138), .ZN(n5004)
         );
  OAI22_X1 U4295 ( .A1(n5004), .A2(n3414), .B1(n4691), .B2(n3456), .ZN(n3420)
         );
  INV_X1 U4296 ( .A(n3415), .ZN(n3418) );
  NAND3_X1 U4297 ( .A1(n3418), .A2(n3417), .A3(n3416), .ZN(n3419) );
  OAI21_X1 U4298 ( .B1(n5005), .B2(n3420), .A(n4958), .ZN(n3425) );
  INV_X1 U4299 ( .A(n3421), .ZN(n5008) );
  OR2_X1 U4300 ( .A1(n3422), .A2(n4433), .ZN(n3482) );
  INV_X1 U4301 ( .A(n3482), .ZN(n3423) );
  AOI22_X1 U4302 ( .A1(n5008), .A2(n4955), .B1(REG2_REG_4__SCAN_IN), .B2(n4698), .ZN(n3424) );
  NAND2_X1 U4303 ( .A1(n3425), .A2(n3424), .ZN(U3286) );
  XNOR2_X1 U4304 ( .A(n3426), .B(n3427), .ZN(n3433) );
  AOI21_X1 U4305 ( .B1(n4260), .B2(n4445), .A(n3428), .ZN(n3429) );
  OAI21_X1 U4306 ( .B1(n3486), .B2(n4280), .A(n3429), .ZN(n3431) );
  NOR2_X1 U4307 ( .A1(n4279), .A2(n3607), .ZN(n3430) );
  AOI211_X1 U4308 ( .C1(n3606), .C2(n4252), .A(n3431), .B(n3430), .ZN(n3432)
         );
  OAI21_X1 U4309 ( .B1(n3433), .B2(n4285), .A(n3432), .ZN(U3224) );
  AOI22_X1 U4310 ( .A1(n4249), .A2(n3117), .B1(n3434), .B2(REG3_REG_0__SCAN_IN), .ZN(n3436) );
  NAND2_X1 U4311 ( .A1(n4252), .A2(n4942), .ZN(n3435) );
  OAI211_X1 U4312 ( .C1(n4285), .C2(n3437), .A(n3436), .B(n3435), .ZN(U3229)
         );
  AOI21_X1 U4313 ( .B1(n4260), .B2(n3119), .A(n3438), .ZN(n3439) );
  OAI21_X1 U4314 ( .B1(n3602), .B2(n4280), .A(n3439), .ZN(n3440) );
  AOI21_X1 U4315 ( .B1(n4300), .B2(n4252), .A(n3440), .ZN(n3446) );
  OAI21_X1 U4316 ( .B1(n3443), .B2(n3442), .A(n3441), .ZN(n3444) );
  NAND2_X1 U4317 ( .A1(n3444), .A2(n4247), .ZN(n3445) );
  OAI211_X1 U4318 ( .C1(REG3_REG_3__SCAN_IN), .C2(n4279), .A(n3446), .B(n3445), 
        .ZN(U3215) );
  AND2_X1 U4319 ( .A1(n3441), .A2(n3447), .ZN(n3450) );
  OAI211_X1 U4320 ( .C1(n3450), .C2(n3449), .A(n4247), .B(n3448), .ZN(n3455)
         );
  AND2_X1 U4321 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4846) );
  AOI21_X1 U4322 ( .B1(n4260), .B2(n4446), .A(n4846), .ZN(n3451) );
  OAI21_X1 U4323 ( .B1(n3513), .B2(n4280), .A(n3451), .ZN(n3452) );
  AOI21_X1 U4324 ( .B1(n3453), .B2(n4252), .A(n3452), .ZN(n3454) );
  OAI211_X1 U4325 ( .C1(n4279), .C2(n3456), .A(n3455), .B(n3454), .ZN(U3227)
         );
  NAND2_X1 U4326 ( .A1(n3850), .A2(n3457), .ZN(n3459) );
  NAND2_X1 U4327 ( .A1(n3459), .A2(n3460), .ZN(n3458) );
  OAI21_X1 U4328 ( .B1(n3460), .B2(n3459), .A(n3458), .ZN(n3461) );
  NAND2_X1 U4329 ( .A1(n3461), .A2(n4247), .ZN(n3465) );
  NAND2_X1 U4330 ( .A1(n4260), .A2(n3629), .ZN(n3462) );
  NAND2_X1 U4331 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4463) );
  OAI211_X1 U4332 ( .C1(n3627), .C2(n4280), .A(n3462), .B(n4463), .ZN(n3463)
         );
  AOI21_X1 U4333 ( .B1(n3634), .B2(n4252), .A(n3463), .ZN(n3464) );
  OAI211_X1 U4334 ( .C1(n4279), .C2(n3635), .A(n3465), .B(n3464), .ZN(U3228)
         );
  OR2_X1 U4335 ( .A1(n3346), .A2(n3466), .ZN(n3468) );
  NAND2_X1 U4336 ( .A1(n3468), .A2(n3467), .ZN(n3470) );
  AOI21_X1 U4337 ( .B1(n3470), .B2(n3469), .A(n4285), .ZN(n3472) );
  OR2_X1 U4338 ( .A1(n3470), .A2(n3469), .ZN(n3471) );
  NAND2_X1 U4339 ( .A1(n3472), .A2(n3471), .ZN(n3478) );
  AOI21_X1 U4340 ( .B1(n4260), .B2(n2135), .A(n3473), .ZN(n3474) );
  OAI21_X1 U4341 ( .B1(n3475), .B2(n4280), .A(n3474), .ZN(n3476) );
  AOI21_X1 U4342 ( .B1(n3490), .B2(n4252), .A(n3476), .ZN(n3477) );
  OAI211_X1 U4343 ( .C1(n4279), .C2(n3491), .A(n3478), .B(n3477), .ZN(U3210)
         );
  OR2_X1 U4344 ( .A1(n3509), .A2(n3479), .ZN(n3481) );
  NAND2_X1 U4345 ( .A1(n3481), .A2(n3480), .ZN(n3620) );
  INV_X1 U4346 ( .A(n4373), .ZN(n4308) );
  XNOR2_X1 U4347 ( .A(n3620), .B(n4308), .ZN(n5018) );
  INV_X1 U4348 ( .A(n5018), .ZN(n3497) );
  NAND2_X1 U4349 ( .A1(n4699), .A2(n3482), .ZN(n3483) );
  XNOR2_X1 U4350 ( .A(n3484), .B(n4373), .ZN(n3489) );
  OAI22_X1 U4351 ( .A1(n3486), .A2(n4618), .B1(n3485), .B2(n4682), .ZN(n3487)
         );
  AOI21_X1 U4352 ( .B1(n4678), .B2(n3629), .A(n3487), .ZN(n3488) );
  OAI21_X1 U4353 ( .B1(n3489), .B2(n4704), .A(n3488), .ZN(n5015) );
  NAND2_X1 U4354 ( .A1(n5015), .A2(n4958), .ZN(n3496) );
  AOI211_X1 U4355 ( .C1(n3490), .C2(n3519), .A(n4779), .B(n3533), .ZN(n5016)
         );
  NAND2_X1 U4356 ( .A1(n4958), .A2(n4433), .ZN(n3771) );
  INV_X1 U4357 ( .A(n3771), .ZN(n3494) );
  OAI22_X1 U4358 ( .A1(n4958), .A2(n3492), .B1(n3491), .B2(n4691), .ZN(n3493)
         );
  AOI21_X1 U4359 ( .B1(n5016), .B2(n3494), .A(n3493), .ZN(n3495) );
  OAI211_X1 U4360 ( .C1(n3497), .C2(n4649), .A(n3496), .B(n3495), .ZN(U3283)
         );
  INV_X1 U4361 ( .A(n3499), .ZN(n3501) );
  NOR2_X1 U4362 ( .A1(n3501), .A2(n3500), .ZN(n3502) );
  XNOR2_X1 U4363 ( .A(n3498), .B(n3502), .ZN(n3507) );
  AND2_X1 U4364 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n4866) );
  AOI21_X1 U4365 ( .B1(n4260), .B2(n4679), .A(n4866), .ZN(n3503) );
  OAI21_X1 U4366 ( .B1(n3689), .B2(n4280), .A(n3503), .ZN(n3505) );
  NOR2_X1 U4367 ( .A1(n4279), .A2(n3671), .ZN(n3504) );
  AOI211_X1 U4368 ( .C1(n3667), .C2(n4283), .A(n3505), .B(n3504), .ZN(n3506)
         );
  OAI21_X1 U4369 ( .B1(n3507), .B2(n4285), .A(n3506), .ZN(U3221) );
  INV_X1 U4370 ( .A(DATAO_REG_25__SCAN_IN), .ZN(n4130) );
  NAND2_X1 U4371 ( .A1(n4583), .A2(U4043), .ZN(n3508) );
  OAI21_X1 U4372 ( .B1(U4043), .B2(n4130), .A(n3508), .ZN(U3575) );
  AND2_X1 U4373 ( .A1(n4307), .A2(n4318), .ZN(n4370) );
  XNOR2_X1 U4374 ( .A(n3509), .B(n4370), .ZN(n3597) );
  XNOR2_X1 U4375 ( .A(n3510), .B(n4370), .ZN(n3515) );
  AOI22_X1 U4376 ( .A1(n4937), .A2(n3517), .B1(n3511), .B2(n4678), .ZN(n3512)
         );
  OAI21_X1 U4377 ( .B1(n3513), .B2(n4618), .A(n3512), .ZN(n3514) );
  AOI21_X1 U4378 ( .B1(n3515), .B2(n4949), .A(n3514), .ZN(n3592) );
  OAI21_X1 U4379 ( .B1(n3597), .B2(n5009), .A(n3592), .ZN(n3657) );
  NAND2_X1 U4380 ( .A1(n3516), .A2(n3517), .ZN(n3518) );
  NAND2_X1 U4381 ( .A1(n3519), .A2(n3518), .ZN(n3655) );
  INV_X1 U4382 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3520) );
  OAI22_X1 U4383 ( .A1(n4820), .A2(n3655), .B1(n5020), .B2(n3520), .ZN(n3521)
         );
  AOI21_X1 U4384 ( .B1(n3657), .B2(n5020), .A(n3521), .ZN(n3522) );
  INV_X1 U4385 ( .A(n3522), .ZN(U3479) );
  INV_X1 U4386 ( .A(DATAO_REG_26__SCAN_IN), .ZN(n4121) );
  NAND2_X1 U4387 ( .A1(n4566), .A2(U4043), .ZN(n3523) );
  OAI21_X1 U4388 ( .B1(U4043), .B2(n4121), .A(n3523), .ZN(U3576) );
  NAND2_X1 U4389 ( .A1(n4312), .A2(n4310), .ZN(n4383) );
  NAND2_X1 U4390 ( .A1(n3620), .A2(n4373), .ZN(n3525) );
  NAND2_X1 U4391 ( .A1(n3525), .A2(n3524), .ZN(n3526) );
  XOR2_X1 U4392 ( .A(n4383), .B(n3526), .Z(n3615) );
  NAND2_X1 U4393 ( .A1(n3527), .A2(n4311), .ZN(n3573) );
  XOR2_X1 U4394 ( .A(n4383), .B(n3573), .Z(n3532) );
  OAI22_X1 U4395 ( .A1(n3529), .A2(n4618), .B1(n3528), .B2(n4952), .ZN(n3530)
         );
  AOI21_X1 U4396 ( .B1(n3535), .B2(n4937), .A(n3530), .ZN(n3531) );
  OAI21_X1 U4397 ( .B1(n3532), .B2(n4704), .A(n3531), .ZN(n3611) );
  AOI21_X1 U4398 ( .B1(n3615), .B2(n5017), .A(n3611), .ZN(n3653) );
  INV_X1 U4399 ( .A(n3533), .ZN(n3534) );
  AOI21_X1 U4400 ( .B1(n3535), .B2(n3534), .A(n3632), .ZN(n3651) );
  INV_X1 U4401 ( .A(n4820), .ZN(n3643) );
  AOI22_X1 U4402 ( .A1(n3651), .A2(n3643), .B1(REG0_REG_8__SCAN_IN), .B2(n5019), .ZN(n3536) );
  OAI21_X1 U4403 ( .B1(n3653), .B2(n5019), .A(n3536), .ZN(U3483) );
  AOI211_X1 U4404 ( .C1(n3539), .C2(n3538), .A(n4902), .B(n3537), .ZN(n3549)
         );
  AND3_X1 U4405 ( .A1(n3542), .A2(n4858), .A3(n3541), .ZN(n3543) );
  NOR3_X1 U4406 ( .A1(n3540), .A2(n3543), .A3(n4896), .ZN(n3548) );
  NAND2_X1 U4407 ( .A1(n4914), .A2(ADDR_REG_11__SCAN_IN), .ZN(n3544) );
  OAI211_X1 U4408 ( .C1(n4926), .C2(n3546), .A(n3545), .B(n3544), .ZN(n3547)
         );
  OR3_X1 U4409 ( .A1(n3549), .A2(n3548), .A3(n3547), .ZN(U3251) );
  XNOR2_X1 U4410 ( .A(n2174), .B(n3551), .ZN(n3552) );
  XNOR2_X1 U4411 ( .A(n3550), .B(n3552), .ZN(n3557) );
  AND2_X1 U4412 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4875) );
  AOI21_X1 U4413 ( .B1(n4260), .B2(n3695), .A(n4875), .ZN(n3553) );
  OAI21_X1 U4414 ( .B1(n3722), .B2(n4280), .A(n3553), .ZN(n3555) );
  NOR2_X1 U4415 ( .A1(n4279), .A2(n3702), .ZN(n3554) );
  AOI211_X1 U4416 ( .C1(n3688), .C2(n4283), .A(n3555), .B(n3554), .ZN(n3556)
         );
  OAI21_X1 U4417 ( .B1(n3557), .B2(n4285), .A(n3556), .ZN(U3231) );
  XNOR2_X1 U4418 ( .A(n3558), .B(n4390), .ZN(n4999) );
  OAI22_X1 U4419 ( .A1(n4940), .A2(n4618), .B1(n3559), .B2(n4682), .ZN(n3565)
         );
  INV_X1 U4420 ( .A(n4390), .ZN(n3561) );
  NAND3_X1 U4421 ( .A1(n3560), .A2(n4296), .A3(n3561), .ZN(n3562) );
  AOI21_X1 U4422 ( .B1(n3563), .B2(n3562), .A(n4704), .ZN(n3564) );
  AOI211_X1 U4423 ( .C1(n4678), .C2(n4445), .A(n3565), .B(n3564), .ZN(n3566)
         );
  OAI21_X1 U4424 ( .B1(n4999), .B2(n4699), .A(n3566), .ZN(n5000) );
  INV_X1 U4425 ( .A(n5000), .ZN(n3572) );
  AOI21_X1 U4426 ( .B1(n4300), .B2(n3567), .A(n3568), .ZN(n5002) );
  INV_X1 U4427 ( .A(n4955), .ZN(n3707) );
  AOI22_X1 U4428 ( .A1(n4698), .A2(REG2_REG_3__SCAN_IN), .B1(n4954), .B2(n4186), .ZN(n3569) );
  OAI21_X1 U4429 ( .B1(n3707), .B2(n4999), .A(n3569), .ZN(n3570) );
  AOI21_X1 U4430 ( .B1(n4943), .B2(n5002), .A(n3570), .ZN(n3571) );
  OAI21_X1 U4431 ( .B1(n3572), .B2(n4698), .A(n3571), .ZN(U3287) );
  NAND2_X1 U4432 ( .A1(n3573), .A2(n4312), .ZN(n3625) );
  NAND2_X1 U4433 ( .A1(n3625), .A2(n3574), .ZN(n3576) );
  NAND2_X1 U4434 ( .A1(n3576), .A2(n3575), .ZN(n3663) );
  XOR2_X1 U4435 ( .A(n4379), .B(n3663), .Z(n3581) );
  AOI22_X1 U4436 ( .A1(n3695), .A2(n4678), .B1(n4935), .B2(n3577), .ZN(n3578)
         );
  OAI21_X1 U4437 ( .B1(n3579), .B2(n4682), .A(n3578), .ZN(n3580) );
  AOI21_X1 U4438 ( .B1(n3581), .B2(n4949), .A(n3580), .ZN(n4777) );
  NAND2_X1 U4439 ( .A1(n2149), .A2(n3582), .ZN(n3583) );
  NAND2_X1 U4440 ( .A1(n3668), .A2(n3583), .ZN(n4778) );
  INV_X1 U4441 ( .A(n4778), .ZN(n3586) );
  OAI22_X1 U4442 ( .A1(n4958), .A2(n4073), .B1(n3584), .B2(n4691), .ZN(n3585)
         );
  AOI21_X1 U4443 ( .B1(n3586), .B2(n4943), .A(n3585), .ZN(n3589) );
  XNOR2_X1 U4444 ( .A(n3587), .B(n4379), .ZN(n4775) );
  INV_X1 U4445 ( .A(n4649), .ZN(n3773) );
  NAND2_X1 U4446 ( .A1(n4775), .A2(n3773), .ZN(n3588) );
  OAI211_X1 U4447 ( .C1(n4777), .C2(n4698), .A(n3589), .B(n3588), .ZN(U3279)
         );
  INV_X1 U4448 ( .A(n3655), .ZN(n3595) );
  OAI22_X1 U4449 ( .A1(n4958), .A2(n3591), .B1(n3590), .B2(n4691), .ZN(n3594)
         );
  NOR2_X1 U4450 ( .A1(n3592), .A2(n4698), .ZN(n3593) );
  AOI211_X1 U4451 ( .C1(n3595), .C2(n4943), .A(n3594), .B(n3593), .ZN(n3596)
         );
  OAI21_X1 U4452 ( .B1(n4649), .B2(n3597), .A(n3596), .ZN(U3284) );
  INV_X1 U4453 ( .A(n3599), .ZN(n4304) );
  NAND2_X1 U4454 ( .A1(n4304), .A2(n4317), .ZN(n4386) );
  XNOR2_X1 U4455 ( .A(n3598), .B(n4386), .ZN(n5010) );
  XNOR2_X1 U4456 ( .A(n3600), .B(n4386), .ZN(n3604) );
  AOI22_X1 U4457 ( .A1(n4937), .A2(n3606), .B1(n2135), .B2(n4678), .ZN(n3601)
         );
  OAI21_X1 U4458 ( .B1(n3602), .B2(n4618), .A(n3601), .ZN(n3603) );
  AOI21_X1 U4459 ( .B1(n3604), .B2(n4949), .A(n3603), .ZN(n5011) );
  MUX2_X1 U4460 ( .A(n5011), .B(n2462), .S(n4698), .Z(n3610) );
  AOI21_X1 U4461 ( .B1(n3606), .B2(n3605), .A(n3100), .ZN(n5014) );
  INV_X1 U4462 ( .A(n3607), .ZN(n3608) );
  AOI22_X1 U4463 ( .A1(n4943), .A2(n5014), .B1(n3608), .B2(n4954), .ZN(n3609)
         );
  OAI211_X1 U4464 ( .C1(n4649), .C2(n5010), .A(n3610), .B(n3609), .ZN(U3285)
         );
  INV_X1 U4465 ( .A(n3611), .ZN(n3618) );
  OAI22_X1 U4466 ( .A1(n4958), .A2(n3613), .B1(n3612), .B2(n4691), .ZN(n3614)
         );
  AOI21_X1 U4467 ( .B1(n3651), .B2(n4943), .A(n3614), .ZN(n3617) );
  NAND2_X1 U4468 ( .A1(n3615), .A2(n3773), .ZN(n3616) );
  OAI211_X1 U4469 ( .C1(n3618), .C2(n4698), .A(n3617), .B(n3616), .ZN(U3282)
         );
  NAND2_X1 U4470 ( .A1(n3620), .A2(n3619), .ZN(n3622) );
  AND2_X1 U4471 ( .A1(n3622), .A2(n3621), .ZN(n3624) );
  INV_X1 U4472 ( .A(n4674), .ZN(n3623) );
  NAND2_X1 U4473 ( .A1(n3623), .A2(n4676), .ZN(n4387) );
  XNOR2_X1 U4474 ( .A(n3624), .B(n4387), .ZN(n3642) );
  INV_X1 U4475 ( .A(n3642), .ZN(n3640) );
  NAND2_X1 U4476 ( .A1(n3625), .A2(n4310), .ZN(n4675) );
  XOR2_X1 U4477 ( .A(n4387), .B(n4675), .Z(n3631) );
  OAI22_X1 U4478 ( .A1(n3627), .A2(n4952), .B1(n3626), .B2(n4682), .ZN(n3628)
         );
  AOI21_X1 U4479 ( .B1(n4935), .B2(n3629), .A(n3628), .ZN(n3630) );
  OAI21_X1 U4480 ( .B1(n3631), .B2(n4704), .A(n3630), .ZN(n3641) );
  NAND2_X1 U4481 ( .A1(n3641), .A2(n4958), .ZN(n3639) );
  INV_X1 U4482 ( .A(n3632), .ZN(n3633) );
  AOI21_X1 U4483 ( .B1(n3634), .B2(n3633), .A(n2273), .ZN(n3647) );
  OAI22_X1 U4484 ( .A1(n4958), .A2(n3636), .B1(n3635), .B2(n4691), .ZN(n3637)
         );
  AOI21_X1 U4485 ( .B1(n3647), .B2(n4943), .A(n3637), .ZN(n3638) );
  OAI211_X1 U4486 ( .C1(n3640), .C2(n4649), .A(n3639), .B(n3638), .ZN(U3281)
         );
  AOI21_X1 U4487 ( .B1(n5017), .B2(n3642), .A(n3641), .ZN(n3649) );
  AOI22_X1 U4488 ( .A1(n3647), .A2(n3643), .B1(REG0_REG_9__SCAN_IN), .B2(n5019), .ZN(n3644) );
  OAI21_X1 U4489 ( .B1(n3649), .B2(n5019), .A(n3644), .ZN(U3485) );
  INV_X1 U4490 ( .A(DATAO_REG_29__SCAN_IN), .ZN(n4101) );
  INV_X1 U4491 ( .A(n4355), .ZN(n3645) );
  NAND2_X1 U4492 ( .A1(n3645), .A2(U4043), .ZN(n3646) );
  OAI21_X1 U4493 ( .B1(U4043), .B2(n4101), .A(n3646), .ZN(U3579) );
  INV_X1 U4494 ( .A(n4761), .ZN(n3650) );
  AOI22_X1 U4495 ( .A1(n3647), .A2(n3650), .B1(REG1_REG_9__SCAN_IN), .B2(n3224), .ZN(n3648) );
  OAI21_X1 U4496 ( .B1(n3649), .B2(n3224), .A(n3648), .ZN(U3527) );
  AOI22_X1 U4497 ( .A1(n3651), .A2(n3650), .B1(REG1_REG_8__SCAN_IN), .B2(n3224), .ZN(n3652) );
  OAI21_X1 U4498 ( .B1(n3653), .B2(n3224), .A(n3652), .ZN(U3526) );
  INV_X1 U4499 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n4115) );
  NAND2_X1 U4500 ( .A1(n4505), .A2(U4043), .ZN(n3654) );
  OAI21_X1 U4501 ( .B1(n4115), .B2(U4043), .A(n3654), .ZN(U3578) );
  OAI22_X1 U4502 ( .A1(n4761), .A2(n3655), .B1(n5030), .B2(n2718), .ZN(n3656)
         );
  AOI21_X1 U4503 ( .B1(n3657), .B2(n5030), .A(n3656), .ZN(n3658) );
  INV_X1 U4504 ( .A(n3658), .ZN(U3524) );
  NAND2_X1 U4505 ( .A1(n3692), .A2(n3690), .ZN(n4392) );
  XNOR2_X1 U4506 ( .A(n3659), .B(n4392), .ZN(n3709) );
  INV_X1 U4507 ( .A(n3709), .ZN(n3676) );
  INV_X1 U4508 ( .A(n3660), .ZN(n3661) );
  AOI21_X1 U4509 ( .B1(n3663), .B2(n3662), .A(n3661), .ZN(n3693) );
  XOR2_X1 U4510 ( .A(n4392), .B(n3693), .Z(n3666) );
  OAI22_X1 U4511 ( .A1(n3689), .A2(n4952), .B1(n3858), .B2(n4618), .ZN(n3664)
         );
  AOI21_X1 U4512 ( .B1(n3667), .B2(n4937), .A(n3664), .ZN(n3665) );
  OAI21_X1 U4513 ( .B1(n3666), .B2(n4704), .A(n3665), .ZN(n3708) );
  INV_X1 U4514 ( .A(n3701), .ZN(n3670) );
  NAND2_X1 U4515 ( .A1(n3668), .A2(n3667), .ZN(n3669) );
  NAND2_X1 U4516 ( .A1(n3670), .A2(n3669), .ZN(n3713) );
  NOR2_X1 U4517 ( .A1(n3713), .A2(n4646), .ZN(n3674) );
  OAI22_X1 U4518 ( .A1(n4958), .A2(n3672), .B1(n3671), .B2(n4691), .ZN(n3673)
         );
  AOI211_X1 U4519 ( .C1(n3708), .C2(n4958), .A(n3674), .B(n3673), .ZN(n3675)
         );
  OAI21_X1 U4520 ( .B1(n3676), .B2(n4649), .A(n3675), .ZN(U3278) );
  OAI21_X1 U4521 ( .B1(n4367), .B2(n4403), .A(n3718), .ZN(n3681) );
  AOI22_X1 U4522 ( .A1(n4444), .A2(n4935), .B1(n3870), .B2(n4937), .ZN(n3677)
         );
  OAI21_X1 U4523 ( .B1(n4211), .B2(n4952), .A(n3677), .ZN(n3680) );
  NOR2_X1 U4524 ( .A1(n3678), .A2(n4367), .ZN(n3743) );
  AOI21_X1 U4525 ( .B1(n4367), .B2(n3678), .A(n3743), .ZN(n4774) );
  NOR2_X1 U4526 ( .A1(n4774), .A2(n4699), .ZN(n3679) );
  AOI211_X1 U4527 ( .C1(n4949), .C2(n3681), .A(n3680), .B(n3679), .ZN(n4773)
         );
  INV_X1 U4528 ( .A(n4774), .ZN(n3685) );
  NAND2_X1 U4529 ( .A1(n3682), .A2(n3870), .ZN(n4770) );
  AND3_X1 U4530 ( .A1(n4771), .A2(n4943), .A3(n4770), .ZN(n3684) );
  OAI22_X1 U4531 ( .A1(n4958), .A2(n4887), .B1(n3867), .B2(n4691), .ZN(n3683)
         );
  AOI211_X1 U4532 ( .C1(n3685), .C2(n4955), .A(n3684), .B(n3683), .ZN(n3686)
         );
  OAI21_X1 U4533 ( .B1(n4773), .B2(n4698), .A(n3686), .ZN(U3276) );
  XNOR2_X1 U4534 ( .A(n3689), .B(n3688), .ZN(n4393) );
  XNOR2_X1 U4535 ( .A(n3687), .B(n4393), .ZN(n3776) );
  INV_X1 U4536 ( .A(n3690), .ZN(n3691) );
  AOI21_X1 U4537 ( .B1(n3693), .B2(n3692), .A(n3691), .ZN(n3694) );
  XOR2_X1 U4538 ( .A(n4393), .B(n3694), .Z(n3698) );
  AOI22_X1 U4539 ( .A1(n3695), .A2(n4935), .B1(n3815), .B2(n4678), .ZN(n3696)
         );
  OAI21_X1 U4540 ( .B1(n3700), .B2(n4682), .A(n3696), .ZN(n3697) );
  AOI21_X1 U4541 ( .B1(n3698), .B2(n4949), .A(n3697), .ZN(n3699) );
  OAI21_X1 U4542 ( .B1(n3776), .B2(n4699), .A(n3699), .ZN(n3777) );
  NAND2_X1 U4543 ( .A1(n3777), .A2(n4958), .ZN(n3706) );
  OAI21_X1 U4544 ( .B1(n3701), .B2(n3700), .A(n3682), .ZN(n3784) );
  INV_X1 U4545 ( .A(n3784), .ZN(n3704) );
  OAI22_X1 U4546 ( .A1(n4958), .A2(n4877), .B1(n3702), .B2(n4691), .ZN(n3703)
         );
  AOI21_X1 U4547 ( .B1(n3704), .B2(n4943), .A(n3703), .ZN(n3705) );
  OAI211_X1 U4548 ( .C1(n3776), .C2(n3707), .A(n3706), .B(n3705), .ZN(U3277)
         );
  AOI21_X1 U4549 ( .B1(n5017), .B2(n3709), .A(n3708), .ZN(n3711) );
  MUX2_X1 U4550 ( .A(n4864), .B(n3711), .S(n5030), .Z(n3710) );
  OAI21_X1 U4551 ( .B1(n4761), .B2(n3713), .A(n3710), .ZN(U3530) );
  MUX2_X1 U4552 ( .A(n4010), .B(n3711), .S(n5020), .Z(n3712) );
  OAI21_X1 U4553 ( .B1(n3713), .B2(n4820), .A(n3712), .ZN(U3491) );
  INV_X1 U4554 ( .A(n4771), .ZN(n3715) );
  INV_X1 U4555 ( .A(n3765), .ZN(n3714) );
  OAI21_X1 U4556 ( .B1(n3715), .B2(n3721), .A(n3714), .ZN(n3801) );
  INV_X1 U4557 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3727) );
  NOR2_X1 U4558 ( .A1(n3743), .A2(n3716), .ZN(n3717) );
  INV_X1 U4559 ( .A(n3719), .ZN(n4369) );
  XNOR2_X1 U4560 ( .A(n3717), .B(n4369), .ZN(n3800) );
  NAND2_X1 U4561 ( .A1(n3718), .A2(n4329), .ZN(n3720) );
  XNOR2_X1 U4562 ( .A(n3720), .B(n3719), .ZN(n3726) );
  OAI22_X1 U4563 ( .A1(n3722), .A2(n4618), .B1(n3721), .B2(n4682), .ZN(n3723)
         );
  AOI21_X1 U4564 ( .B1(n3724), .B2(n4678), .A(n3723), .ZN(n3725) );
  OAI21_X1 U4565 ( .B1(n3726), .B2(n4704), .A(n3725), .ZN(n3805) );
  AOI21_X1 U4566 ( .B1(n3800), .B2(n5017), .A(n3805), .ZN(n3729) );
  MUX2_X1 U4567 ( .A(n3727), .B(n3729), .S(n5020), .Z(n3728) );
  OAI21_X1 U4568 ( .B1(n3801), .B2(n4820), .A(n3728), .ZN(U3497) );
  MUX2_X1 U4569 ( .A(n3979), .B(n3729), .S(n5030), .Z(n3730) );
  OAI21_X1 U4570 ( .B1(n4761), .B2(n3801), .A(n3730), .ZN(U3533) );
  NAND2_X1 U4571 ( .A1(n2185), .A2(n3732), .ZN(n3733) );
  XNOR2_X1 U4572 ( .A(n3731), .B(n3733), .ZN(n3739) );
  NOR2_X1 U4573 ( .A1(n3734), .A2(STATE_REG_SCAN_IN), .ZN(n4913) );
  NOR2_X1 U4574 ( .A1(n4277), .A2(n3817), .ZN(n3735) );
  AOI211_X1 U4575 ( .C1(n4249), .C2(n3792), .A(n4913), .B(n3735), .ZN(n3736)
         );
  OAI21_X1 U4576 ( .B1(n3923), .B2(n3790), .A(n3736), .ZN(n3737) );
  AOI21_X1 U4577 ( .B1(n3826), .B2(n3920), .A(n3737), .ZN(n3738) );
  OAI21_X1 U4578 ( .B1(n3739), .B2(n4285), .A(n3738), .ZN(U3225) );
  INV_X1 U4579 ( .A(n3740), .ZN(n3741) );
  AOI21_X1 U4580 ( .B1(n3743), .B2(n3742), .A(n3741), .ZN(n3744) );
  XNOR2_X1 U4581 ( .A(n3744), .B(n4378), .ZN(n4769) );
  XNOR2_X1 U4582 ( .A(n3745), .B(n4378), .ZN(n3749) );
  AOI22_X1 U4583 ( .A1(n4443), .A2(n4935), .B1(n4215), .B2(n4937), .ZN(n3746)
         );
  OAI21_X1 U4584 ( .B1(n3747), .B2(n4952), .A(n3746), .ZN(n3748) );
  AOI21_X1 U4585 ( .B1(n3749), .B2(n4949), .A(n3748), .ZN(n4768) );
  INV_X1 U4586 ( .A(n4768), .ZN(n3754) );
  NOR2_X1 U4587 ( .A1(n3765), .A2(n3750), .ZN(n4765) );
  AND2_X1 U4588 ( .A1(n3765), .A2(n3750), .ZN(n4766) );
  NOR3_X1 U4589 ( .A1(n4765), .A2(n4766), .A3(n4646), .ZN(n3753) );
  INV_X1 U4590 ( .A(REG2_REG_16__SCAN_IN), .ZN(n3751) );
  OAI22_X1 U4591 ( .A1(n4958), .A2(n3751), .B1(n4212), .B2(n4691), .ZN(n3752)
         );
  AOI211_X1 U4592 ( .C1(n3754), .C2(n4958), .A(n3753), .B(n3752), .ZN(n3755)
         );
  OAI21_X1 U4593 ( .B1(n4769), .B2(n4649), .A(n3755), .ZN(U3274) );
  OAI21_X1 U4594 ( .B1(n3756), .B2(n3786), .A(n3787), .ZN(n3839) );
  INV_X1 U4595 ( .A(n3761), .ZN(n4377) );
  XNOR2_X1 U4596 ( .A(n3839), .B(n4377), .ZN(n3759) );
  AOI22_X1 U4597 ( .A1(n4259), .A2(n4935), .B1(n4266), .B2(n4937), .ZN(n3757)
         );
  OAI21_X1 U4598 ( .B1(n4262), .B2(n4952), .A(n3757), .ZN(n3758) );
  AOI21_X1 U4599 ( .B1(n3759), .B2(n4949), .A(n3758), .ZN(n4763) );
  INV_X1 U4600 ( .A(n3760), .ZN(n3763) );
  NAND2_X1 U4601 ( .A1(n3760), .A2(n3761), .ZN(n3835) );
  INV_X1 U4602 ( .A(n3835), .ZN(n3762) );
  AOI21_X1 U4603 ( .B1(n4377), .B2(n3763), .A(n3762), .ZN(n4764) );
  INV_X1 U4604 ( .A(n4764), .ZN(n3774) );
  NAND2_X1 U4605 ( .A1(n3765), .A2(n3764), .ZN(n3785) );
  INV_X1 U4606 ( .A(n3785), .ZN(n3768) );
  OAI211_X1 U4607 ( .C1(n3768), .C2(n3767), .A(n2138), .B(n3766), .ZN(n4762)
         );
  INV_X1 U4608 ( .A(n4263), .ZN(n3769) );
  AOI22_X1 U4609 ( .A1(n4698), .A2(REG2_REG_18__SCAN_IN), .B1(n3769), .B2(
        n4954), .ZN(n3770) );
  OAI21_X1 U4610 ( .B1(n4762), .B2(n3771), .A(n3770), .ZN(n3772) );
  AOI21_X1 U4611 ( .B1(n3774), .B2(n3773), .A(n3772), .ZN(n3775) );
  OAI21_X1 U4612 ( .B1(n4698), .B2(n4763), .A(n3775), .ZN(U3272) );
  INV_X1 U4613 ( .A(n4998), .ZN(n5007) );
  INV_X1 U4614 ( .A(n3776), .ZN(n3778) );
  AOI21_X1 U4615 ( .B1(n5007), .B2(n3778), .A(n3777), .ZN(n3781) );
  MUX2_X1 U4616 ( .A(n3779), .B(n3781), .S(n5030), .Z(n3780) );
  OAI21_X1 U4617 ( .B1(n4761), .B2(n3784), .A(n3780), .ZN(U3531) );
  INV_X1 U4618 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3782) );
  MUX2_X1 U4619 ( .A(n3782), .B(n3781), .S(n5020), .Z(n3783) );
  OAI21_X1 U4620 ( .B1(n3784), .B2(n4820), .A(n3783), .ZN(U3493) );
  OAI21_X1 U4621 ( .B1(n4766), .B2(n3790), .A(n3785), .ZN(n3825) );
  INV_X1 U4622 ( .A(REG0_REG_17__SCAN_IN), .ZN(n3795) );
  INV_X1 U4623 ( .A(n3786), .ZN(n3788) );
  NAND2_X1 U4624 ( .A1(n3788), .A2(n3787), .ZN(n4380) );
  XOR2_X1 U4625 ( .A(n3789), .B(n4380), .Z(n3824) );
  XOR2_X1 U4626 ( .A(n3756), .B(n4380), .Z(n3794) );
  OAI22_X1 U4627 ( .A1(n3817), .A2(n4618), .B1(n3790), .B2(n4682), .ZN(n3791)
         );
  AOI21_X1 U4628 ( .B1(n3792), .B2(n4678), .A(n3791), .ZN(n3793) );
  OAI21_X1 U4629 ( .B1(n3794), .B2(n4704), .A(n3793), .ZN(n3831) );
  AOI21_X1 U4630 ( .B1(n3824), .B2(n5017), .A(n3831), .ZN(n3797) );
  MUX2_X1 U4631 ( .A(n3795), .B(n3797), .S(n5020), .Z(n3796) );
  OAI21_X1 U4632 ( .B1(n3825), .B2(n4820), .A(n3796), .ZN(U3501) );
  MUX2_X1 U4633 ( .A(n3798), .B(n3797), .S(n5030), .Z(n3799) );
  OAI21_X1 U4634 ( .B1(n4761), .B2(n3825), .A(n3799), .ZN(U3535) );
  INV_X1 U4635 ( .A(n3800), .ZN(n3807) );
  NOR2_X1 U4636 ( .A1(n3801), .A2(n4646), .ZN(n3804) );
  OAI22_X1 U4637 ( .A1(n4958), .A2(n3802), .B1(n3818), .B2(n4691), .ZN(n3803)
         );
  AOI211_X1 U4638 ( .C1(n3805), .C2(n4958), .A(n3804), .B(n3803), .ZN(n3806)
         );
  OAI21_X1 U4639 ( .B1(n3807), .B2(n4649), .A(n3806), .ZN(U3275) );
  INV_X1 U4640 ( .A(n3808), .ZN(n3810) );
  INV_X1 U4641 ( .A(n3809), .ZN(n3864) );
  NOR2_X1 U4642 ( .A1(n3810), .A2(n3864), .ZN(n3812) );
  NOR2_X1 U4643 ( .A1(n3812), .A2(n3811), .ZN(n4205) );
  INV_X1 U4644 ( .A(n4205), .ZN(n3813) );
  NAND2_X1 U4645 ( .A1(n3812), .A2(n3811), .ZN(n4206) );
  NAND2_X1 U4646 ( .A1(n3813), .A2(n4206), .ZN(n3814) );
  XNOR2_X1 U4647 ( .A(n3814), .B(n4207), .ZN(n3823) );
  NAND2_X1 U4648 ( .A1(n4260), .A2(n3815), .ZN(n3816) );
  NAND2_X1 U4649 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4909) );
  OAI211_X1 U4650 ( .C1(n3817), .C2(n4280), .A(n3816), .B(n4909), .ZN(n3820)
         );
  NOR2_X1 U4651 ( .A1(n4279), .A2(n3818), .ZN(n3819) );
  AOI211_X1 U4652 ( .C1(n3821), .C2(n4283), .A(n3820), .B(n3819), .ZN(n3822)
         );
  OAI21_X1 U4653 ( .B1(n3823), .B2(n4285), .A(n3822), .ZN(U3238) );
  INV_X1 U4654 ( .A(n3824), .ZN(n3833) );
  NOR2_X1 U4655 ( .A1(n3825), .A2(n4646), .ZN(n3830) );
  INV_X1 U4656 ( .A(n3826), .ZN(n3827) );
  OAI22_X1 U4657 ( .A1(n4958), .A2(n3828), .B1(n3827), .B2(n4691), .ZN(n3829)
         );
  AOI211_X1 U4658 ( .C1(n3831), .C2(n4958), .A(n3830), .B(n3829), .ZN(n3832)
         );
  OAI21_X1 U4659 ( .B1(n3833), .B2(n4649), .A(n3832), .ZN(U3273) );
  NAND2_X1 U4660 ( .A1(n4660), .A2(n4658), .ZN(n4375) );
  NAND2_X1 U4661 ( .A1(n3835), .A2(n3834), .ZN(n4659) );
  XOR2_X1 U4662 ( .A(n4375), .B(n4659), .Z(n4758) );
  INV_X1 U4663 ( .A(n4758), .ZN(n3848) );
  INV_X1 U4664 ( .A(n3836), .ZN(n3838) );
  OAI21_X1 U4665 ( .B1(n3839), .B2(n3838), .A(n3837), .ZN(n3840) );
  XNOR2_X1 U4666 ( .A(n3840), .B(n4375), .ZN(n3843) );
  OAI22_X1 U4667 ( .A1(n3900), .A2(n4618), .B1(n3844), .B2(n4682), .ZN(n3841)
         );
  AOI21_X1 U4668 ( .B1(n4636), .B2(n4678), .A(n3841), .ZN(n3842) );
  OAI21_X1 U4669 ( .B1(n3843), .B2(n4704), .A(n3842), .ZN(n4757) );
  OAI21_X1 U4670 ( .B1(n2280), .B2(n3844), .A(n2150), .ZN(n4821) );
  AOI22_X1 U4671 ( .A1(n4698), .A2(REG2_REG_19__SCAN_IN), .B1(n3893), .B2(
        n4954), .ZN(n3845) );
  OAI21_X1 U4672 ( .B1(n4821), .B2(n4646), .A(n3845), .ZN(n3846) );
  AOI21_X1 U4673 ( .B1(n4757), .B2(n4958), .A(n3846), .ZN(n3847) );
  OAI21_X1 U4674 ( .B1(n3848), .B2(n4649), .A(n3847), .ZN(U3271) );
  NAND2_X1 U4675 ( .A1(n3850), .A2(n3849), .ZN(n3852) );
  AND2_X1 U4676 ( .A1(n3852), .A2(n3851), .ZN(n3854) );
  AOI21_X1 U4677 ( .B1(n3854), .B2(n3853), .A(n4285), .ZN(n3856) );
  NAND2_X1 U4678 ( .A1(n3856), .A2(n3855), .ZN(n3861) );
  AND2_X1 U4679 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n4857) );
  AOI21_X1 U4680 ( .B1(n4260), .B2(n4680), .A(n4857), .ZN(n3857) );
  OAI21_X1 U4681 ( .B1(n3858), .B2(n4280), .A(n3857), .ZN(n3859) );
  AOI21_X1 U4682 ( .B1(n4689), .B2(n4252), .A(n3859), .ZN(n3860) );
  OAI211_X1 U4683 ( .C1(n4279), .C2(n4692), .A(n3861), .B(n3860), .ZN(U3214)
         );
  NOR2_X1 U4684 ( .A1(n3864), .A2(n3863), .ZN(n3865) );
  XNOR2_X1 U4685 ( .A(n3862), .B(n3865), .ZN(n3872) );
  NAND2_X1 U4686 ( .A1(n4260), .A2(n4444), .ZN(n3866) );
  NAND2_X1 U4687 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n4891) );
  OAI211_X1 U4688 ( .C1(n4211), .C2(n4280), .A(n3866), .B(n4891), .ZN(n3869)
         );
  NOR2_X1 U4689 ( .A1(n4279), .A2(n3867), .ZN(n3868) );
  AOI211_X1 U4690 ( .C1(n3870), .C2(n4283), .A(n3869), .B(n3868), .ZN(n3871)
         );
  OAI21_X1 U4691 ( .B1(n3872), .B2(n4285), .A(n3871), .ZN(U3212) );
  XNOR2_X1 U4692 ( .A(n3874), .B(n3873), .ZN(n3880) );
  OAI22_X1 U4693 ( .A1(n3875), .A2(n4277), .B1(STATE_REG_SCAN_IN), .B2(n3992), 
        .ZN(n3876) );
  AOI21_X1 U4694 ( .B1(n4535), .B2(n4252), .A(n3876), .ZN(n3877) );
  OAI21_X1 U4695 ( .B1(n4279), .B2(n4530), .A(n3877), .ZN(n3878) );
  AOI21_X1 U4696 ( .B1(n4249), .B2(n4505), .A(n3878), .ZN(n3879) );
  OAI21_X1 U4697 ( .B1(n3880), .B2(n4285), .A(n3879), .ZN(U3211) );
  INV_X1 U4698 ( .A(n3886), .ZN(n3881) );
  NOR2_X1 U4699 ( .A1(n3881), .A2(n3884), .ZN(n3888) );
  XNOR2_X1 U4700 ( .A(n3883), .B(n3882), .ZN(n3887) );
  INV_X1 U4701 ( .A(n3884), .ZN(n3885) );
  OAI211_X1 U4702 ( .C1(n3888), .C2(n3887), .A(n4247), .B(n4221), .ZN(n3892)
         );
  AOI22_X1 U4703 ( .A1(n4603), .A2(n4249), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3889) );
  OAI21_X1 U4704 ( .B1(n4601), .B2(n4277), .A(n3889), .ZN(n3890) );
  AOI21_X1 U4705 ( .B1(n4606), .B2(n4252), .A(n3890), .ZN(n3891) );
  OAI211_X1 U4706 ( .C1(n4279), .C2(n4609), .A(n3892), .B(n3891), .ZN(U3213)
         );
  INV_X1 U4707 ( .A(n3893), .ZN(n3905) );
  OAI21_X1 U4708 ( .B1(n3896), .B2(n3895), .A(n3894), .ZN(n3897) );
  NAND2_X1 U4709 ( .A1(n3897), .A2(n4247), .ZN(n3904) );
  NAND2_X1 U4710 ( .A1(n4249), .A2(n4636), .ZN(n3899) );
  OAI211_X1 U4711 ( .C1(n3900), .C2(n4277), .A(n3899), .B(n3898), .ZN(n3901)
         );
  AOI21_X1 U4712 ( .B1(n3902), .B2(n4252), .A(n3901), .ZN(n3903) );
  OAI211_X1 U4713 ( .C1(n4279), .C2(n3905), .A(n3904), .B(n3903), .ZN(U3216)
         );
  XNOR2_X1 U4714 ( .A(n3907), .B(n3906), .ZN(n3908) );
  XNOR2_X1 U4715 ( .A(n3909), .B(n3908), .ZN(n3916) );
  AOI22_X1 U4716 ( .A1(n4639), .A2(n4249), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3912) );
  NAND2_X1 U4717 ( .A1(n4252), .A2(n3910), .ZN(n3911) );
  OAI211_X1 U4718 ( .C1(n3913), .C2(n4277), .A(n3912), .B(n3911), .ZN(n3914)
         );
  AOI21_X1 U4719 ( .B1(n4644), .B2(n3920), .A(n3914), .ZN(n3915) );
  OAI21_X1 U4720 ( .B1(n3916), .B2(n4285), .A(n3915), .ZN(U3220) );
  INV_X1 U4721 ( .A(n4272), .ZN(n3917) );
  NOR2_X1 U4722 ( .A1(n4271), .A2(n3917), .ZN(n3918) );
  XNOR2_X1 U4723 ( .A(n4273), .B(n3918), .ZN(n3925) );
  OAI22_X1 U4724 ( .A1(n4564), .A2(n4277), .B1(STATE_REG_SCAN_IN), .B2(n4043), 
        .ZN(n3919) );
  AOI21_X1 U4725 ( .B1(n4566), .B2(n4249), .A(n3919), .ZN(n3922) );
  NAND2_X1 U4726 ( .A1(n4571), .A2(n3920), .ZN(n3921) );
  OAI211_X1 U4727 ( .C1(n3923), .C2(n4570), .A(n3922), .B(n3921), .ZN(n3924)
         );
  AOI21_X1 U4728 ( .B1(n3925), .B2(n4247), .A(n3924), .ZN(n4202) );
  NOR4_X1 U4729 ( .A1(REG3_REG_28__SCAN_IN), .A2(REG2_REG_20__SCAN_IN), .A3(
        REG2_REG_30__SCAN_IN), .A4(n4276), .ZN(n3949) );
  NOR4_X1 U4730 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        n2672), .A4(n2655), .ZN(n3948) );
  INV_X1 U4731 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n4063) );
  NOR4_X1 U4732 ( .A1(REG3_REG_1__SCAN_IN), .A2(ADDR_REG_7__SCAN_IN), .A3(
        n3591), .A4(n4063), .ZN(n3926) );
  NAND3_X1 U4733 ( .A1(DATAI_27_), .A2(REG2_REG_16__SCAN_IN), .A3(n3926), .ZN(
        n3935) );
  INV_X1 U4734 ( .A(n3927), .ZN(n3932) );
  INV_X1 U4735 ( .A(REG2_REG_25__SCAN_IN), .ZN(n3929) );
  NOR4_X1 U4736 ( .A1(n3929), .A2(n4188), .A3(n3928), .A4(REG2_REG_28__SCAN_IN), .ZN(n3931) );
  INV_X1 U4737 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n3930) );
  NAND4_X1 U4738 ( .A1(n3933), .A2(n3932), .A3(n3931), .A4(n3930), .ZN(n3934)
         );
  NOR4_X1 U4739 ( .A1(REG2_REG_10__SCAN_IN), .A2(REG2_REG_8__SCAN_IN), .A3(
        n3935), .A4(n3934), .ZN(n3947) );
  NAND4_X1 U4740 ( .A1(ADDR_REG_1__SCAN_IN), .A2(DATAO_REG_7__SCAN_IN), .A3(
        DATAO_REG_29__SCAN_IN), .A4(n4104), .ZN(n3945) );
  NAND4_X1 U4741 ( .A1(DATAO_REG_24__SCAN_IN), .A2(DATAO_REG_18__SCAN_IN), 
        .A3(n4162), .A4(n4164), .ZN(n3944) );
  INV_X1 U4742 ( .A(DATAI_16_), .ZN(n4143) );
  NAND4_X1 U4743 ( .A1(DATAO_REG_21__SCAN_IN), .A2(REG3_REG_18__SCAN_IN), .A3(
        ADDR_REG_0__SCAN_IN), .A4(n4148), .ZN(n3936) );
  NOR3_X1 U4744 ( .A1(DATAO_REG_17__SCAN_IN), .A2(n4143), .A3(n3936), .ZN(
        n3937) );
  NAND3_X1 U4745 ( .A1(DATAO_REG_10__SCAN_IN), .A2(n3937), .A3(n4133), .ZN(
        n3943) );
  NOR4_X1 U4746 ( .A1(DATAO_REG_22__SCAN_IN), .A2(ADDR_REG_2__SCAN_IN), .A3(
        n4108), .A4(n4115), .ZN(n3941) );
  NOR4_X1 U4747 ( .A1(DATAO_REG_2__SCAN_IN), .A2(DATAO_REG_0__SCAN_IN), .A3(
        ADDR_REG_14__SCAN_IN), .A4(n4109), .ZN(n3940) );
  NOR4_X1 U4748 ( .A1(ADDR_REG_15__SCAN_IN), .A2(DATAO_REG_5__SCAN_IN), .A3(
        n4130), .A4(n4134), .ZN(n3939) );
  NOR4_X1 U4749 ( .A1(DATAO_REG_26__SCAN_IN), .A2(DATAO_REG_12__SCAN_IN), .A3(
        DATAO_REG_6__SCAN_IN), .A4(n2286), .ZN(n3938) );
  NAND4_X1 U4750 ( .A1(n3941), .A2(n3940), .A3(n3939), .A4(n3938), .ZN(n3942)
         );
  NOR4_X1 U4751 ( .A1(n3945), .A2(n3944), .A3(n3943), .A4(n3942), .ZN(n3946)
         );
  NAND4_X1 U4752 ( .A1(n3949), .A2(n3948), .A3(n3947), .A4(n3946), .ZN(n3977)
         );
  NAND4_X1 U4753 ( .A1(D_REG_14__SCAN_IN), .A2(REG1_REG_21__SCAN_IN), .A3(
        n4733), .A4(n4036), .ZN(n3950) );
  NOR3_X1 U4754 ( .A1(REG0_REG_21__SCAN_IN), .A2(REG0_REG_15__SCAN_IN), .A3(
        n3950), .ZN(n3961) );
  NOR4_X1 U4755 ( .A1(IR_REG_3__SCAN_IN), .A2(REG0_REG_7__SCAN_IN), .A3(
        REG0_REG_4__SCAN_IN), .A4(n4014), .ZN(n3954) );
  INV_X1 U4756 ( .A(DATAI_10_), .ZN(n4982) );
  NAND4_X1 U4757 ( .A1(REG0_REG_12__SCAN_IN), .A2(REG1_REG_10__SCAN_IN), .A3(
        n4864), .A4(n4982), .ZN(n3952) );
  INV_X1 U4758 ( .A(DATAI_8_), .ZN(n4086) );
  NAND4_X1 U4759 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_10__SCAN_IN), .A3(
        DATAI_6_), .A4(n4086), .ZN(n3951) );
  NOR2_X1 U4760 ( .A1(n3952), .A2(n3951), .ZN(n3953) );
  NAND4_X1 U4761 ( .A1(n3955), .A2(n4039), .A3(n3954), .A4(n3953), .ZN(n3959)
         );
  NAND4_X1 U4762 ( .A1(n3956), .A2(IR_REG_6__SCAN_IN), .A3(IR_REG_11__SCAN_IN), 
        .A4(DATAI_2_), .ZN(n3958) );
  NOR4_X1 U4763 ( .A1(n3959), .A2(n3958), .A3(REG1_REG_29__SCAN_IN), .A4(n3957), .ZN(n3960) );
  NAND2_X1 U4764 ( .A1(n3961), .A2(n3960), .ZN(n3964) );
  NOR4_X1 U4765 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG2_REG_15__SCAN_IN), .A3(
        REG1_REG_30__SCAN_IN), .A4(n3636), .ZN(n3962) );
  NAND3_X1 U4766 ( .A1(REG2_REG_29__SCAN_IN), .A2(REG2_REG_11__SCAN_IN), .A3(
        n3962), .ZN(n3963) );
  NOR2_X1 U4767 ( .A1(n3964), .A2(n3963), .ZN(n3975) );
  NAND4_X1 U4768 ( .A1(IR_REG_13__SCAN_IN), .A2(REG0_REG_18__SCAN_IN), .A3(
        n2504), .A4(n2896), .ZN(n3968) );
  INV_X1 U4769 ( .A(DATAI_13_), .ZN(n4979) );
  NAND4_X1 U4770 ( .A1(REG3_REG_11__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .A3(
        DATAI_9_), .A4(n4979), .ZN(n3967) );
  NAND4_X1 U4771 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .A3(
        DATAI_30_), .A4(n4003), .ZN(n3966) );
  NAND4_X1 U4772 ( .A1(DATAI_22_), .A2(REG0_REG_22__SCAN_IN), .A3(
        REG0_REG_19__SCAN_IN), .A4(n4092), .ZN(n3965) );
  NOR4_X1 U4773 ( .A1(n3968), .A2(n3967), .A3(n3966), .A4(n3965), .ZN(n3974)
         );
  NAND4_X1 U4774 ( .A1(REG1_REG_1__SCAN_IN), .A2(n5027), .A3(n5021), .A4(n3979), .ZN(n3972) );
  INV_X1 U4775 ( .A(ADDR_REG_13__SCAN_IN), .ZN(n3981) );
  NAND4_X1 U4776 ( .A1(ADDR_REG_10__SCAN_IN), .A2(ADDR_REG_12__SCAN_IN), .A3(
        n3672), .A4(n3981), .ZN(n3971) );
  NAND4_X1 U4777 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_31__SCAN_IN), .A3(
        D_REG_3__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n3970) );
  NAND4_X1 U4778 ( .A1(D_REG_0__SCAN_IN), .A2(D_REG_5__SCAN_IN), .A3(
        REG1_REG_26__SCAN_IN), .A4(n4174), .ZN(n3969) );
  NOR4_X1 U4779 ( .A1(n3972), .A2(n3971), .A3(n3970), .A4(n3969), .ZN(n3973)
         );
  NAND3_X1 U4780 ( .A1(n3975), .A2(n3974), .A3(n3973), .ZN(n3976) );
  OAI21_X1 U4781 ( .B1(n3977), .B2(n3976), .A(n4182), .ZN(n4200) );
  INV_X1 U4782 ( .A(keyinput8), .ZN(n4199) );
  AOI22_X1 U4783 ( .A1(n3979), .A2(keyinput127), .B1(n5021), .B2(keyinput16), 
        .ZN(n3978) );
  OAI221_X1 U4784 ( .B1(n3979), .B2(keyinput127), .C1(n5021), .C2(keyinput16), 
        .A(n3978), .ZN(n3988) );
  INV_X1 U4785 ( .A(ADDR_REG_12__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4786 ( .A1(n3982), .A2(keyinput87), .B1(keyinput12), .B2(n3981), 
        .ZN(n3980) );
  OAI221_X1 U4787 ( .B1(n3982), .B2(keyinput87), .C1(n3981), .C2(keyinput12), 
        .A(n3980), .ZN(n3987) );
  AOI22_X1 U4788 ( .A1(n3802), .A2(keyinput3), .B1(n3636), .B2(keyinput83), 
        .ZN(n3983) );
  OAI221_X1 U4789 ( .B1(n3802), .B2(keyinput3), .C1(n3636), .C2(keyinput83), 
        .A(n3983), .ZN(n3986) );
  AOI22_X1 U4790 ( .A1(n2646), .A2(keyinput62), .B1(n5027), .B2(keyinput119), 
        .ZN(n3984) );
  OAI221_X1 U4791 ( .B1(n2646), .B2(keyinput62), .C1(n5027), .C2(keyinput119), 
        .A(n3984), .ZN(n3985) );
  NOR4_X1 U4792 ( .A1(n3988), .A2(n3987), .A3(n3986), .A4(n3985), .ZN(n4000)
         );
  INV_X1 U4793 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4492) );
  AOI22_X1 U4794 ( .A1(n3990), .A2(keyinput113), .B1(keyinput60), .B2(n4492), 
        .ZN(n3989) );
  OAI221_X1 U4795 ( .B1(n3990), .B2(keyinput113), .C1(n4492), .C2(keyinput60), 
        .A(n3989), .ZN(n3998) );
  AOI22_X1 U4796 ( .A1(n3992), .A2(keyinput4), .B1(keyinput54), .B2(n4276), 
        .ZN(n3991) );
  OAI221_X1 U4797 ( .B1(n3992), .B2(keyinput4), .C1(n4276), .C2(keyinput54), 
        .A(n3991), .ZN(n3997) );
  INV_X1 U4798 ( .A(REG3_REG_1__SCAN_IN), .ZN(n4448) );
  AOI22_X1 U4799 ( .A1(n3024), .A2(keyinput44), .B1(keyinput110), .B2(n4448), 
        .ZN(n3993) );
  OAI221_X1 U4800 ( .B1(n3024), .B2(keyinput44), .C1(n4448), .C2(keyinput110), 
        .A(n3993), .ZN(n3996) );
  AOI22_X1 U4801 ( .A1(n4669), .A2(keyinput18), .B1(keyinput9), .B2(n3751), 
        .ZN(n3994) );
  OAI221_X1 U4802 ( .B1(n4669), .B2(keyinput18), .C1(n3751), .C2(keyinput9), 
        .A(n3994), .ZN(n3995) );
  NOR4_X1 U4803 ( .A1(n3998), .A2(n3997), .A3(n3996), .A4(n3995), .ZN(n3999)
         );
  NAND2_X1 U4804 ( .A1(n4000), .A2(n3999), .ZN(n4198) );
  AOI22_X1 U4805 ( .A1(n2478), .A2(keyinput85), .B1(keyinput89), .B2(n4864), 
        .ZN(n4001) );
  OAI221_X1 U4806 ( .B1(n2478), .B2(keyinput85), .C1(n4864), .C2(keyinput89), 
        .A(n4001), .ZN(n4005) );
  AOI22_X1 U4807 ( .A1(n2621), .A2(keyinput82), .B1(n4003), .B2(keyinput47), 
        .ZN(n4002) );
  OAI221_X1 U4808 ( .B1(n2621), .B2(keyinput82), .C1(n4003), .C2(keyinput47), 
        .A(n4002), .ZN(n4004) );
  NOR2_X1 U4809 ( .A1(n4005), .A2(n4004), .ZN(n4034) );
  INV_X1 U4810 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4811 ( .A1(n4008), .A2(keyinput13), .B1(n4007), .B2(keyinput36), 
        .ZN(n4006) );
  OAI221_X1 U4812 ( .B1(n4008), .B2(keyinput13), .C1(n4007), .C2(keyinput36), 
        .A(n4006), .ZN(n4012) );
  AOI22_X1 U4813 ( .A1(n4010), .A2(keyinput92), .B1(keyinput91), .B2(n4855), 
        .ZN(n4009) );
  OAI221_X1 U4814 ( .B1(n4010), .B2(keyinput92), .C1(n4855), .C2(keyinput91), 
        .A(n4009), .ZN(n4011) );
  NOR2_X1 U4815 ( .A1(n4012), .A2(n4011), .ZN(n4033) );
  AOI22_X1 U4816 ( .A1(n2727), .A2(keyinput63), .B1(n4014), .B2(keyinput97), 
        .ZN(n4013) );
  OAI221_X1 U4817 ( .B1(n2727), .B2(keyinput63), .C1(n4014), .C2(keyinput97), 
        .A(n4013), .ZN(n4020) );
  XNOR2_X1 U4818 ( .A(IR_REG_0__SCAN_IN), .B(keyinput59), .ZN(n4018) );
  XNOR2_X1 U4819 ( .A(IR_REG_3__SCAN_IN), .B(keyinput115), .ZN(n4017) );
  XNOR2_X1 U4820 ( .A(IR_REG_1__SCAN_IN), .B(keyinput56), .ZN(n4016) );
  XNOR2_X1 U4821 ( .A(IR_REG_13__SCAN_IN), .B(keyinput53), .ZN(n4015) );
  NAND4_X1 U4822 ( .A1(n4018), .A2(n4017), .A3(n4016), .A4(n4015), .ZN(n4019)
         );
  NOR2_X1 U4823 ( .A1(n4020), .A2(n4019), .ZN(n4032) );
  XNOR2_X1 U4824 ( .A(IR_REG_9__SCAN_IN), .B(keyinput46), .ZN(n4024) );
  XNOR2_X1 U4825 ( .A(IR_REG_22__SCAN_IN), .B(keyinput88), .ZN(n4023) );
  XNOR2_X1 U4826 ( .A(REG0_REG_15__SCAN_IN), .B(keyinput98), .ZN(n4022) );
  XNOR2_X1 U4827 ( .A(IR_REG_31__SCAN_IN), .B(keyinput64), .ZN(n4021) );
  NAND4_X1 U4828 ( .A1(n4024), .A2(n4023), .A3(n4022), .A4(n4021), .ZN(n4030)
         );
  XNOR2_X1 U4829 ( .A(DATAI_1_), .B(keyinput112), .ZN(n4028) );
  XNOR2_X1 U4830 ( .A(IR_REG_15__SCAN_IN), .B(keyinput77), .ZN(n4027) );
  XNOR2_X1 U4831 ( .A(DATAI_2_), .B(keyinput105), .ZN(n4026) );
  XNOR2_X1 U4832 ( .A(IR_REG_6__SCAN_IN), .B(keyinput1), .ZN(n4025) );
  NAND4_X1 U4833 ( .A1(n4028), .A2(n4027), .A3(n4026), .A4(n4025), .ZN(n4029)
         );
  NOR2_X1 U4834 ( .A1(n4030), .A2(n4029), .ZN(n4031) );
  NAND4_X1 U4835 ( .A1(n4034), .A2(n4033), .A3(n4032), .A4(n4031), .ZN(n4060)
         );
  AOI22_X1 U4836 ( .A1(n4733), .A2(keyinput25), .B1(keyinput111), .B2(n4036), 
        .ZN(n4035) );
  OAI221_X1 U4837 ( .B1(n4733), .B2(keyinput25), .C1(n4036), .C2(keyinput111), 
        .A(n4035), .ZN(n4041) );
  AOI22_X1 U4838 ( .A1(n4039), .A2(keyinput117), .B1(keyinput86), .B2(n4038), 
        .ZN(n4037) );
  OAI221_X1 U4839 ( .B1(n4039), .B2(keyinput117), .C1(n4038), .C2(keyinput86), 
        .A(n4037), .ZN(n4040) );
  NOR2_X1 U4840 ( .A1(n4041), .A2(n4040), .ZN(n4058) );
  AOI22_X1 U4841 ( .A1(n4043), .A2(keyinput68), .B1(keyinput58), .B2(n4729), 
        .ZN(n4042) );
  OAI221_X1 U4842 ( .B1(n4043), .B2(keyinput68), .C1(n4729), .C2(keyinput58), 
        .A(n4042), .ZN(n4048) );
  AOI22_X1 U4843 ( .A1(n4046), .A2(keyinput11), .B1(keyinput72), .B2(n4045), 
        .ZN(n4044) );
  OAI221_X1 U4844 ( .B1(n4046), .B2(keyinput11), .C1(n4045), .C2(keyinput72), 
        .A(n4044), .ZN(n4047) );
  NOR2_X1 U4845 ( .A1(n4048), .A2(n4047), .ZN(n4057) );
  AOI22_X1 U4846 ( .A1(n4050), .A2(keyinput5), .B1(keyinput120), .B2(n4979), 
        .ZN(n4049) );
  OAI221_X1 U4847 ( .B1(n4050), .B2(keyinput5), .C1(n4979), .C2(keyinput120), 
        .A(n4049), .ZN(n4051) );
  INV_X1 U4848 ( .A(n4051), .ZN(n4056) );
  AOI22_X1 U4849 ( .A1(n4053), .A2(keyinput7), .B1(n2896), .B2(keyinput70), 
        .ZN(n4052) );
  OAI221_X1 U4850 ( .B1(n4053), .B2(keyinput7), .C1(n2896), .C2(keyinput70), 
        .A(n4052), .ZN(n4054) );
  INV_X1 U4851 ( .A(n4054), .ZN(n4055) );
  NAND4_X1 U4852 ( .A1(n4058), .A2(n4057), .A3(n4056), .A4(n4055), .ZN(n4059)
         );
  NOR2_X1 U4853 ( .A1(n4060), .A2(n4059), .ZN(n4099) );
  AOI22_X1 U4854 ( .A1(n3613), .A2(keyinput114), .B1(n4693), .B2(keyinput15), 
        .ZN(n4061) );
  OAI221_X1 U4855 ( .B1(n3613), .B2(keyinput114), .C1(n4693), .C2(keyinput15), 
        .A(n4061), .ZN(n4082) );
  AOI22_X1 U4856 ( .A1(n4982), .A2(keyinput76), .B1(n2474), .B2(keyinput42), 
        .ZN(n4062) );
  OAI221_X1 U4857 ( .B1(n4982), .B2(keyinput76), .C1(n2474), .C2(keyinput42), 
        .A(n4062), .ZN(n4081) );
  XNOR2_X1 U4858 ( .A(keyinput123), .B(n4063), .ZN(n4065) );
  XNOR2_X1 U4859 ( .A(keyinput108), .B(n3955), .ZN(n4064) );
  NOR2_X1 U4860 ( .A1(n4065), .A2(n4064), .ZN(n4079) );
  INV_X1 U4861 ( .A(DATAI_6_), .ZN(n4066) );
  XNOR2_X1 U4862 ( .A(keyinput99), .B(n4066), .ZN(n4068) );
  XNOR2_X1 U4863 ( .A(keyinput101), .B(n2504), .ZN(n4067) );
  NOR2_X1 U4864 ( .A1(n4068), .A2(n4067), .ZN(n4078) );
  XNOR2_X1 U4865 ( .A(keyinput69), .B(n4069), .ZN(n4071) );
  XNOR2_X1 U4866 ( .A(keyinput57), .B(n2682), .ZN(n4070) );
  NOR2_X1 U4867 ( .A1(n4071), .A2(n4070), .ZN(n4077) );
  INV_X1 U4868 ( .A(DATAI_9_), .ZN(n4072) );
  XNOR2_X1 U4869 ( .A(keyinput65), .B(n4072), .ZN(n4075) );
  XNOR2_X1 U4870 ( .A(keyinput35), .B(n4073), .ZN(n4074) );
  NOR2_X1 U4871 ( .A1(n4075), .A2(n4074), .ZN(n4076) );
  NAND4_X1 U4872 ( .A1(n4079), .A2(n4078), .A3(n4077), .A4(n4076), .ZN(n4080)
         );
  NOR3_X1 U4873 ( .A1(n4082), .A2(n4081), .A3(n4080), .ZN(n4098) );
  INV_X1 U4874 ( .A(ADDR_REG_10__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U4875 ( .A1(n4084), .A2(keyinput39), .B1(n3672), .B2(keyinput19), 
        .ZN(n4083) );
  OAI221_X1 U4876 ( .B1(n4084), .B2(keyinput39), .C1(n3672), .C2(keyinput19), 
        .A(n4083), .ZN(n4088) );
  AOI22_X1 U4877 ( .A1(n4086), .A2(keyinput22), .B1(n2467), .B2(keyinput0), 
        .ZN(n4085) );
  OAI221_X1 U4878 ( .B1(n4086), .B2(keyinput22), .C1(n2467), .C2(keyinput0), 
        .A(n4085), .ZN(n4087) );
  NOR2_X1 U4879 ( .A1(n4088), .A2(n4087), .ZN(n4097) );
  AOI22_X1 U4880 ( .A1(n3591), .A2(keyinput21), .B1(keyinput52), .B2(n3288), 
        .ZN(n4089) );
  OAI221_X1 U4881 ( .B1(n3591), .B2(keyinput21), .C1(n3288), .C2(keyinput52), 
        .A(n4089), .ZN(n4095) );
  AOI22_X1 U4882 ( .A1(n4750), .A2(keyinput126), .B1(n4813), .B2(keyinput2), 
        .ZN(n4090) );
  OAI221_X1 U4883 ( .B1(n4750), .B2(keyinput126), .C1(n4813), .C2(keyinput2), 
        .A(n4090), .ZN(n4094) );
  AOI22_X1 U4884 ( .A1(n4818), .A2(keyinput96), .B1(n4092), .B2(keyinput125), 
        .ZN(n4091) );
  OAI221_X1 U4885 ( .B1(n4818), .B2(keyinput96), .C1(n4092), .C2(keyinput125), 
        .A(n4091), .ZN(n4093) );
  NOR3_X1 U4886 ( .A1(n4095), .A2(n4094), .A3(n4093), .ZN(n4096) );
  NAND4_X1 U4887 ( .A1(n4099), .A2(n4098), .A3(n4097), .A4(n4096), .ZN(n4158)
         );
  INV_X1 U4888 ( .A(D_REG_10__SCAN_IN), .ZN(n4968) );
  AOI22_X1 U4889 ( .A1(n4968), .A2(keyinput26), .B1(keyinput29), .B2(n4101), 
        .ZN(n4100) );
  OAI221_X1 U4890 ( .B1(n4968), .B2(keyinput26), .C1(n4101), .C2(keyinput29), 
        .A(n4100), .ZN(n4113) );
  AOI22_X1 U4891 ( .A1(n4104), .A2(keyinput28), .B1(keyinput41), .B2(n4103), 
        .ZN(n4102) );
  OAI221_X1 U4892 ( .B1(n4104), .B2(keyinput28), .C1(n4103), .C2(keyinput41), 
        .A(n4102), .ZN(n4112) );
  INV_X1 U4893 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n4893) );
  AOI22_X1 U4894 ( .A1(n4106), .A2(keyinput40), .B1(keyinput33), .B2(n4893), 
        .ZN(n4105) );
  OAI221_X1 U4895 ( .B1(n4106), .B2(keyinput40), .C1(n4893), .C2(keyinput33), 
        .A(n4105), .ZN(n4111) );
  AOI22_X1 U4896 ( .A1(n4109), .A2(keyinput32), .B1(keyinput34), .B2(n4108), 
        .ZN(n4107) );
  OAI221_X1 U4897 ( .B1(n4109), .B2(keyinput32), .C1(n4108), .C2(keyinput34), 
        .A(n4107), .ZN(n4110) );
  NOR4_X1 U4898 ( .A1(n4113), .A2(n4112), .A3(n4111), .A4(n4110), .ZN(n4156)
         );
  AOI22_X1 U4899 ( .A1(n4116), .A2(keyinput37), .B1(keyinput6), .B2(n4115), 
        .ZN(n4114) );
  OAI221_X1 U4900 ( .B1(n4116), .B2(keyinput37), .C1(n4115), .C2(keyinput6), 
        .A(n4114), .ZN(n4127) );
  INV_X1 U4901 ( .A(ADDR_REG_2__SCAN_IN), .ZN(n4119) );
  AOI22_X1 U4902 ( .A1(n4119), .A2(keyinput17), .B1(keyinput14), .B2(n4118), 
        .ZN(n4117) );
  OAI221_X1 U4903 ( .B1(n4119), .B2(keyinput17), .C1(n4118), .C2(keyinput14), 
        .A(n4117), .ZN(n4126) );
  AOI22_X1 U4904 ( .A1(n4121), .A2(keyinput124), .B1(n2286), .B2(keyinput116), 
        .ZN(n4120) );
  OAI221_X1 U4905 ( .B1(n4121), .B2(keyinput124), .C1(n2286), .C2(keyinput116), 
        .A(n4120), .ZN(n4125) );
  AOI22_X1 U4906 ( .A1(n4123), .A2(keyinput118), .B1(n4962), .B2(keyinput106), 
        .ZN(n4122) );
  OAI221_X1 U4907 ( .B1(n4123), .B2(keyinput118), .C1(n4962), .C2(keyinput106), 
        .A(n4122), .ZN(n4124) );
  NOR4_X1 U4908 ( .A1(n4127), .A2(n4126), .A3(n4125), .A4(n4124), .ZN(n4155)
         );
  AOI22_X1 U4909 ( .A1(n4130), .A2(keyinput109), .B1(keyinput100), .B2(n4129), 
        .ZN(n4128) );
  OAI221_X1 U4910 ( .B1(n4130), .B2(keyinput109), .C1(n4129), .C2(keyinput100), 
        .A(n4128), .ZN(n4141) );
  INV_X1 U4911 ( .A(ADDR_REG_15__SCAN_IN), .ZN(n4912) );
  AOI22_X1 U4912 ( .A1(n4966), .A2(keyinput102), .B1(keyinput90), .B2(n4912), 
        .ZN(n4131) );
  OAI221_X1 U4913 ( .B1(n4966), .B2(keyinput102), .C1(n4912), .C2(keyinput90), 
        .A(n4131), .ZN(n4140) );
  AOI22_X1 U4914 ( .A1(n4134), .A2(keyinput93), .B1(keyinput84), .B2(n4133), 
        .ZN(n4132) );
  OAI221_X1 U4915 ( .B1(n4134), .B2(keyinput93), .C1(n4133), .C2(keyinput84), 
        .A(n4132), .ZN(n4139) );
  AOI22_X1 U4916 ( .A1(n4137), .A2(keyinput81), .B1(keyinput80), .B2(n4136), 
        .ZN(n4135) );
  OAI221_X1 U4917 ( .B1(n4137), .B2(keyinput81), .C1(n4136), .C2(keyinput80), 
        .A(n4135), .ZN(n4138) );
  NOR4_X1 U4918 ( .A1(n4141), .A2(n4140), .A3(n4139), .A4(n4138), .ZN(n4154)
         );
  AOI22_X1 U4919 ( .A1(n4143), .A2(keyinput78), .B1(n4965), .B2(keyinput74), 
        .ZN(n4142) );
  OAI221_X1 U4920 ( .B1(n4143), .B2(keyinput78), .C1(n4965), .C2(keyinput74), 
        .A(n4142), .ZN(n4152) );
  AOI22_X1 U4921 ( .A1(n4145), .A2(keyinput73), .B1(n2297), .B2(keyinput66), 
        .ZN(n4144) );
  OAI221_X1 U4922 ( .B1(n4145), .B2(keyinput73), .C1(n2297), .C2(keyinput66), 
        .A(n4144), .ZN(n4151) );
  AOI22_X1 U4923 ( .A1(n4964), .A2(keyinput61), .B1(keyinput50), .B2(n3257), 
        .ZN(n4146) );
  OAI221_X1 U4924 ( .B1(n4964), .B2(keyinput61), .C1(n3257), .C2(keyinput50), 
        .A(n4146), .ZN(n4150) );
  INV_X1 U4925 ( .A(D_REG_9__SCAN_IN), .ZN(n4969) );
  AOI22_X1 U4926 ( .A1(n4969), .A2(keyinput48), .B1(keyinput45), .B2(n4148), 
        .ZN(n4147) );
  OAI221_X1 U4927 ( .B1(n4969), .B2(keyinput48), .C1(n4148), .C2(keyinput45), 
        .A(n4147), .ZN(n4149) );
  NOR4_X1 U4928 ( .A1(n4152), .A2(n4151), .A3(n4150), .A4(n4149), .ZN(n4153)
         );
  NAND4_X1 U4929 ( .A1(n4156), .A2(n4155), .A3(n4154), .A4(n4153), .ZN(n4157)
         );
  NOR2_X1 U4930 ( .A1(n4158), .A2(n4157), .ZN(n4196) );
  AOI22_X1 U4931 ( .A1(n3103), .A2(keyinput55), .B1(keyinput43), .B2(n4160), 
        .ZN(n4159) );
  OAI221_X1 U4932 ( .B1(n3103), .B2(keyinput55), .C1(n4160), .C2(keyinput43), 
        .A(n4159), .ZN(n4171) );
  INV_X1 U4933 ( .A(D_REG_30__SCAN_IN), .ZN(n4961) );
  AOI22_X1 U4934 ( .A1(n4961), .A2(keyinput23), .B1(keyinput103), .B2(n4162), 
        .ZN(n4161) );
  OAI221_X1 U4935 ( .B1(n4961), .B2(keyinput23), .C1(n4162), .C2(keyinput103), 
        .A(n4161), .ZN(n4170) );
  AOI22_X1 U4936 ( .A1(n4165), .A2(keyinput79), .B1(keyinput95), .B2(n4164), 
        .ZN(n4163) );
  OAI221_X1 U4937 ( .B1(n4165), .B2(keyinput79), .C1(n4164), .C2(keyinput95), 
        .A(n4163), .ZN(n4169) );
  INV_X1 U4938 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n4449) );
  AOI22_X1 U4939 ( .A1(n4167), .A2(keyinput51), .B1(keyinput71), .B2(n4449), 
        .ZN(n4166) );
  OAI221_X1 U4940 ( .B1(n4167), .B2(keyinput51), .C1(n4449), .C2(keyinput71), 
        .A(n4166), .ZN(n4168) );
  NOR4_X1 U4941 ( .A1(n4171), .A2(n4170), .A3(n4169), .A4(n4168), .ZN(n4195)
         );
  AOI22_X1 U4942 ( .A1(n4971), .A2(keyinput24), .B1(keyinput104), .B2(n4963), 
        .ZN(n4172) );
  OAI221_X1 U4943 ( .B1(n4971), .B2(keyinput24), .C1(n4963), .C2(keyinput104), 
        .A(n4172), .ZN(n4181) );
  AOI22_X1 U4944 ( .A1(n4175), .A2(keyinput49), .B1(keyinput31), .B2(n4174), 
        .ZN(n4173) );
  OAI221_X1 U4945 ( .B1(n4175), .B2(keyinput49), .C1(n4174), .C2(keyinput31), 
        .A(n4173), .ZN(n4180) );
  INV_X1 U4946 ( .A(D_REG_8__SCAN_IN), .ZN(n4970) );
  INV_X1 U4947 ( .A(D_REG_14__SCAN_IN), .ZN(n4967) );
  AOI22_X1 U4948 ( .A1(n4970), .A2(keyinput107), .B1(keyinput121), .B2(n4967), 
        .ZN(n4176) );
  OAI221_X1 U4949 ( .B1(n4970), .B2(keyinput107), .C1(n4967), .C2(keyinput121), 
        .A(n4176), .ZN(n4179) );
  INV_X1 U4950 ( .A(D_REG_31__SCAN_IN), .ZN(n4960) );
  INV_X1 U4951 ( .A(D_REG_3__SCAN_IN), .ZN(n4972) );
  AOI22_X1 U4952 ( .A1(n4960), .A2(keyinput38), .B1(keyinput20), .B2(n4972), 
        .ZN(n4177) );
  OAI221_X1 U4953 ( .B1(n4960), .B2(keyinput38), .C1(n4972), .C2(keyinput20), 
        .A(n4177), .ZN(n4178) );
  NOR4_X1 U4954 ( .A1(n4181), .A2(n4180), .A3(n4179), .A4(n4178), .ZN(n4194)
         );
  AOI22_X1 U4955 ( .A1(keyinput94), .A2(n3930), .B1(keyinput8), .B2(n4182), 
        .ZN(n4183) );
  OAI21_X1 U4956 ( .B1(n3930), .B2(keyinput94), .A(n4183), .ZN(n4192) );
  AOI22_X1 U4957 ( .A1(n3032), .A2(keyinput30), .B1(keyinput122), .B2(n3929), 
        .ZN(n4184) );
  OAI221_X1 U4958 ( .B1(n3032), .B2(keyinput30), .C1(n3929), .C2(keyinput122), 
        .A(n4184), .ZN(n4191) );
  AOI22_X1 U4959 ( .A1(n4186), .A2(keyinput75), .B1(keyinput10), .B2(n2655), 
        .ZN(n4185) );
  OAI221_X1 U4960 ( .B1(n4186), .B2(keyinput75), .C1(n2655), .C2(keyinput10), 
        .A(n4185), .ZN(n4190) );
  AOI22_X1 U4961 ( .A1(n4188), .A2(keyinput67), .B1(keyinput27), .B2(n2672), 
        .ZN(n4187) );
  OAI221_X1 U4962 ( .B1(n4188), .B2(keyinput67), .C1(n2672), .C2(keyinput27), 
        .A(n4187), .ZN(n4189) );
  NOR4_X1 U4963 ( .A1(n4192), .A2(n4191), .A3(n4190), .A4(n4189), .ZN(n4193)
         );
  NAND4_X1 U4964 ( .A1(n4196), .A2(n4195), .A3(n4194), .A4(n4193), .ZN(n4197)
         );
  AOI211_X1 U4965 ( .C1(n4200), .C2(n4199), .A(n4198), .B(n4197), .ZN(n4201)
         );
  XNOR2_X1 U4966 ( .A(n4202), .B(n4201), .ZN(U3222) );
  NAND2_X1 U4967 ( .A1(n4204), .A2(n4203), .ZN(n4209) );
  AOI21_X1 U4968 ( .B1(n4207), .B2(n4206), .A(n4205), .ZN(n4208) );
  XOR2_X1 U4969 ( .A(n4209), .B(n4208), .Z(n4217) );
  NOR2_X1 U4970 ( .A1(n2286), .A2(STATE_REG_SCAN_IN), .ZN(n4475) );
  AOI21_X1 U4971 ( .B1(n4249), .B2(n4259), .A(n4475), .ZN(n4210) );
  OAI21_X1 U4972 ( .B1(n4211), .B2(n4277), .A(n4210), .ZN(n4214) );
  NOR2_X1 U4973 ( .A1(n4279), .A2(n4212), .ZN(n4213) );
  AOI211_X1 U4974 ( .C1(n4215), .C2(n4283), .A(n4214), .B(n4213), .ZN(n4216)
         );
  OAI21_X1 U4975 ( .B1(n4217), .B2(n4285), .A(n4216), .ZN(U3223) );
  INV_X1 U4976 ( .A(n4219), .ZN(n4218) );
  NAND2_X1 U4977 ( .A1(n4221), .A2(n4218), .ZN(n4223) );
  NOR2_X1 U4978 ( .A1(n4219), .A2(n4222), .ZN(n4220) );
  AOI22_X1 U4979 ( .A1(n4223), .A2(n4222), .B1(n4221), .B2(n4220), .ZN(n4225)
         );
  XNOR2_X1 U4980 ( .A(n4225), .B(n2977), .ZN(n4231) );
  OAI22_X1 U4981 ( .A1(n4581), .A2(n4277), .B1(STATE_REG_SCAN_IN), .B2(n4226), 
        .ZN(n4227) );
  AOI21_X1 U4982 ( .B1(n4583), .B2(n4249), .A(n4227), .ZN(n4229) );
  NAND2_X1 U4983 ( .A1(n4252), .A2(n3158), .ZN(n4228) );
  OAI211_X1 U4984 ( .C1(n4279), .C2(n4587), .A(n4229), .B(n4228), .ZN(n4230)
         );
  AOI21_X1 U4985 ( .B1(n4231), .B2(n4247), .A(n4230), .ZN(n4232) );
  INV_X1 U4986 ( .A(n4232), .ZN(U3226) );
  INV_X1 U4987 ( .A(n4233), .ZN(n4238) );
  AOI21_X1 U4988 ( .B1(n4237), .B2(n4235), .A(n4234), .ZN(n4236) );
  AOI21_X1 U4989 ( .B1(n4238), .B2(n4237), .A(n4236), .ZN(n4245) );
  NAND2_X1 U4990 ( .A1(n4239), .A2(n4249), .ZN(n4241) );
  NAND2_X1 U4991 ( .A1(U3149), .A2(REG3_REG_20__SCAN_IN), .ZN(n4240) );
  OAI211_X1 U4992 ( .C1(n4262), .C2(n4277), .A(n4241), .B(n4240), .ZN(n4243)
         );
  NOR2_X1 U4993 ( .A1(n4279), .A2(n4668), .ZN(n4242) );
  AOI211_X1 U4994 ( .C1(n4667), .C2(n4252), .A(n4243), .B(n4242), .ZN(n4244)
         );
  OAI21_X1 U4995 ( .B1(n4245), .B2(n4285), .A(n4244), .ZN(U3230) );
  OAI21_X1 U4996 ( .B1(n4246), .B2(n2148), .A(n3886), .ZN(n4248) );
  NAND2_X1 U4997 ( .A1(n4248), .A2(n4247), .ZN(n4254) );
  AOI22_X1 U4998 ( .A1(n4624), .A2(n4249), .B1(REG3_REG_22__SCAN_IN), .B2(
        U3149), .ZN(n4250) );
  OAI21_X1 U4999 ( .B1(n4657), .B2(n4277), .A(n4250), .ZN(n4251) );
  AOI21_X1 U5000 ( .B1(n3155), .B2(n4252), .A(n4251), .ZN(n4253) );
  OAI211_X1 U5001 ( .C1(n4279), .C2(n4627), .A(n4254), .B(n4253), .ZN(U3232)
         );
  NOR2_X1 U5002 ( .A1(n2186), .A2(n4256), .ZN(n4257) );
  XNOR2_X1 U5003 ( .A(n4255), .B(n4257), .ZN(n4268) );
  AOI21_X1 U5004 ( .B1(n4260), .B2(n4259), .A(n4258), .ZN(n4261) );
  OAI21_X1 U5005 ( .B1(n4262), .B2(n4280), .A(n4261), .ZN(n4265) );
  NOR2_X1 U5006 ( .A1(n4279), .A2(n4263), .ZN(n4264) );
  AOI211_X1 U5007 ( .C1(n4266), .C2(n4283), .A(n4265), .B(n4264), .ZN(n4267)
         );
  OAI21_X1 U5008 ( .B1(n4268), .B2(n4285), .A(n4267), .ZN(U3235) );
  NAND2_X1 U5009 ( .A1(n4270), .A2(n4269), .ZN(n4275) );
  AOI21_X1 U5010 ( .B1(n4273), .B2(n4272), .A(n4271), .ZN(n4274) );
  XOR2_X1 U5011 ( .A(n4275), .B(n4274), .Z(n4286) );
  OAI22_X1 U5012 ( .A1(n4278), .A2(n4277), .B1(STATE_REG_SCAN_IN), .B2(n4276), 
        .ZN(n4282) );
  OAI22_X1 U5013 ( .A1(n4550), .A2(n4280), .B1(n4279), .B2(n4553), .ZN(n4281)
         );
  AOI211_X1 U5014 ( .C1(n4547), .C2(n4283), .A(n4282), .B(n4281), .ZN(n4284)
         );
  OAI21_X1 U5015 ( .B1(n4286), .B2(n4285), .A(n4284), .ZN(U3237) );
  OR2_X1 U5016 ( .A1(n4355), .A2(n4506), .ZN(n4287) );
  NAND2_X1 U5017 ( .A1(n4502), .A2(n4287), .ZN(n4348) );
  INV_X1 U5018 ( .A(n4288), .ZN(n4289) );
  NOR2_X1 U5019 ( .A1(n4348), .A2(n4289), .ZN(n4424) );
  INV_X1 U5020 ( .A(n4424), .ZN(n4344) );
  INV_X1 U5021 ( .A(n4290), .ZN(n4291) );
  AOI211_X1 U5022 ( .C1(n4413), .C2(n4291), .A(n4360), .B(n2242), .ZN(n4416)
         );
  INV_X1 U5023 ( .A(n4411), .ZN(n4341) );
  NAND2_X1 U5024 ( .A1(n4293), .A2(n4292), .ZN(n4295) );
  AND2_X1 U5025 ( .A1(n4947), .A2(n4936), .ZN(n4366) );
  INV_X1 U5026 ( .A(n4366), .ZN(n4294) );
  NAND3_X1 U5027 ( .A1(n4297), .A2(n4296), .A3(n3164), .ZN(n4299) );
  OAI211_X1 U5028 ( .C1(n4300), .C2(n3121), .A(n4299), .B(n4298), .ZN(n4303)
         );
  NAND3_X1 U5029 ( .A1(n4303), .A2(n4302), .A3(n4301), .ZN(n4306) );
  NAND4_X1 U5030 ( .A1(n4306), .A2(n4305), .A3(n4304), .A4(n4318), .ZN(n4309)
         );
  NAND3_X1 U5031 ( .A1(n4309), .A2(n4308), .A3(n4307), .ZN(n4314) );
  AND2_X1 U5032 ( .A1(n4311), .A2(n4310), .ZN(n4320) );
  NAND2_X1 U5033 ( .A1(n4676), .A2(n4312), .ZN(n4313) );
  AOI21_X1 U5034 ( .B1(n4314), .B2(n4320), .A(n4313), .ZN(n4325) );
  NAND2_X1 U5035 ( .A1(n4316), .A2(n4315), .ZN(n4324) );
  NAND2_X1 U5036 ( .A1(n4324), .A2(n4330), .ZN(n4401) );
  INV_X1 U5037 ( .A(n4401), .ZN(n4323) );
  INV_X1 U5038 ( .A(n4317), .ZN(n4319) );
  NAND3_X1 U5039 ( .A1(n4320), .A2(n4319), .A3(n4318), .ZN(n4321) );
  AND2_X1 U5040 ( .A1(n4321), .A2(n4385), .ZN(n4322) );
  OAI22_X1 U5041 ( .A1(n4325), .A2(n4324), .B1(n4323), .B2(n4322), .ZN(n4328)
         );
  NAND2_X1 U5042 ( .A1(n4385), .A2(n4674), .ZN(n4326) );
  NAND4_X1 U5043 ( .A1(n4328), .A2(n4327), .A3(n4384), .A4(n4326), .ZN(n4335)
         );
  NAND2_X1 U5044 ( .A1(n4330), .A2(n4329), .ZN(n4402) );
  INV_X1 U5045 ( .A(n4402), .ZN(n4331) );
  NAND2_X1 U5046 ( .A1(n4332), .A2(n4331), .ZN(n4333) );
  NAND2_X1 U5047 ( .A1(n4333), .A2(n4401), .ZN(n4334) );
  NAND2_X1 U5048 ( .A1(n4335), .A2(n4334), .ZN(n4336) );
  NAND2_X1 U5049 ( .A1(n4336), .A2(n4404), .ZN(n4337) );
  AOI21_X1 U5050 ( .B1(n4337), .B2(n4407), .A(n4406), .ZN(n4339) );
  OAI211_X1 U5051 ( .C1(n4339), .C2(n4338), .A(n4363), .B(n2169), .ZN(n4340)
         );
  NAND4_X1 U5052 ( .A1(n4413), .A2(n4596), .A3(n4341), .A4(n4340), .ZN(n4342)
         );
  AOI21_X1 U5053 ( .B1(n4416), .B2(n4342), .A(n4421), .ZN(n4343) );
  AOI211_X1 U5054 ( .C1(n4442), .C2(n4345), .A(n4344), .B(n4343), .ZN(n4352)
         );
  AND2_X1 U5055 ( .A1(n4500), .A2(n4346), .ZN(n4418) );
  NAND2_X1 U5056 ( .A1(n4441), .A2(n4430), .ZN(n4349) );
  OR2_X1 U5057 ( .A1(n4507), .A2(n4483), .ZN(n4347) );
  NAND2_X1 U5058 ( .A1(n4349), .A2(n4347), .ZN(n4381) );
  AOI21_X1 U5059 ( .B1(n4355), .B2(n4506), .A(n4381), .ZN(n4419) );
  OAI21_X1 U5060 ( .B1(n4418), .B2(n4348), .A(n4419), .ZN(n4423) );
  INV_X1 U5061 ( .A(n4349), .ZN(n4351) );
  NAND2_X1 U5062 ( .A1(n4507), .A2(n4483), .ZN(n4425) );
  OAI21_X1 U5063 ( .B1(n4441), .B2(n4430), .A(n4425), .ZN(n4382) );
  INV_X1 U5064 ( .A(n4382), .ZN(n4350) );
  OAI22_X1 U5065 ( .A1(n4352), .A2(n4423), .B1(n4351), .B2(n4350), .ZN(n4432)
         );
  INV_X1 U5066 ( .A(n4353), .ZN(n4493) );
  XNOR2_X1 U5067 ( .A(n4355), .B(n4354), .ZN(n4716) );
  INV_X1 U5068 ( .A(n4356), .ZN(n4357) );
  NOR2_X1 U5069 ( .A1(n4358), .A2(n4357), .ZN(n4544) );
  NAND2_X1 U5070 ( .A1(n4541), .A2(n4359), .ZN(n4560) );
  NAND2_X1 U5071 ( .A1(n2244), .A2(n4361), .ZN(n4579) );
  NAND2_X1 U5072 ( .A1(n4577), .A2(n4362), .ZN(n4599) );
  INV_X1 U5073 ( .A(n4599), .ZN(n4398) );
  INV_X1 U5074 ( .A(n4620), .ZN(n4397) );
  INV_X1 U5075 ( .A(n4363), .ZN(n4414) );
  NOR2_X1 U5076 ( .A1(n4411), .A2(n4414), .ZN(n4633) );
  NAND2_X1 U5077 ( .A1(n4365), .A2(n4364), .ZN(n4662) );
  NOR2_X1 U5078 ( .A1(n4366), .A2(n4932), .ZN(n4948) );
  NAND4_X1 U5079 ( .A1(n4369), .A2(n4368), .A3(n4367), .A4(n4948), .ZN(n4374)
         );
  NAND2_X1 U5080 ( .A1(n4933), .A2(n4370), .ZN(n4371) );
  NOR4_X1 U5081 ( .A1(n4374), .A2(n4373), .A3(n4372), .A4(n4371), .ZN(n4376)
         );
  NAND4_X1 U5082 ( .A1(n4662), .A2(n4377), .A3(n4376), .A4(n4375), .ZN(n4395)
         );
  NOR3_X1 U5083 ( .A1(n4380), .A2(n4379), .A3(n4378), .ZN(n4391) );
  NOR3_X1 U5084 ( .A1(n4383), .A2(n4382), .A3(n4381), .ZN(n4389) );
  NAND2_X1 U5085 ( .A1(n4385), .A2(n4384), .ZN(n4685) );
  NOR3_X1 U5086 ( .A1(n4387), .A2(n4386), .A3(n4685), .ZN(n4388) );
  NAND4_X1 U5087 ( .A1(n4391), .A2(n4390), .A3(n4389), .A4(n4388), .ZN(n4394)
         );
  NOR4_X1 U5088 ( .A1(n4395), .A2(n4394), .A3(n4393), .A4(n4392), .ZN(n4396)
         );
  NAND4_X1 U5089 ( .A1(n4398), .A2(n4397), .A3(n4633), .A4(n4396), .ZN(n4399)
         );
  NOR4_X1 U5090 ( .A1(n4544), .A2(n4560), .A3(n4579), .A4(n4399), .ZN(n4400)
         );
  NAND4_X1 U5091 ( .A1(n4493), .A2(n2235), .A3(n4716), .A4(n4400), .ZN(n4431)
         );
  INV_X1 U5092 ( .A(n4483), .ZN(n4487) );
  OAI21_X1 U5093 ( .B1(n4403), .B2(n4402), .A(n4401), .ZN(n4408) );
  NAND2_X1 U5094 ( .A1(n2169), .A2(n4404), .ZN(n4405) );
  AOI211_X1 U5095 ( .C1(n4408), .C2(n4407), .A(n4406), .B(n4405), .ZN(n4412)
         );
  INV_X1 U5096 ( .A(n4409), .ZN(n4410) );
  NOR3_X1 U5097 ( .A1(n4412), .A2(n4411), .A3(n4410), .ZN(n4415) );
  OAI211_X1 U5098 ( .C1(n4415), .C2(n4414), .A(n4413), .B(n4596), .ZN(n4417)
         );
  NAND2_X1 U5099 ( .A1(n4417), .A2(n4416), .ZN(n4429) );
  INV_X1 U5100 ( .A(n4418), .ZN(n4422) );
  INV_X1 U5101 ( .A(n4419), .ZN(n4420) );
  NOR3_X1 U5102 ( .A1(n4422), .A2(n4421), .A3(n4420), .ZN(n4428) );
  AOI21_X1 U5103 ( .B1(n2235), .B2(n4424), .A(n4423), .ZN(n4427) );
  AOI21_X1 U5104 ( .B1(n4425), .B2(n4441), .A(n4430), .ZN(n4426) );
  XNOR2_X1 U5105 ( .A(n4434), .B(n4433), .ZN(n4440) );
  NAND2_X1 U5106 ( .A1(n4436), .A2(n4435), .ZN(n4437) );
  OAI211_X1 U5107 ( .C1(n4828), .C2(n4439), .A(n4437), .B(B_REG_SCAN_IN), .ZN(
        n4438) );
  OAI21_X1 U5108 ( .B1(n4440), .B2(n4439), .A(n4438), .ZN(U3239) );
  MUX2_X1 U5109 ( .A(n4441), .B(DATAO_REG_31__SCAN_IN), .S(n4447), .Z(U3581)
         );
  MUX2_X1 U5110 ( .A(n4442), .B(DATAO_REG_27__SCAN_IN), .S(n4447), .Z(U3577)
         );
  MUX2_X1 U5111 ( .A(n4624), .B(DATAO_REG_23__SCAN_IN), .S(n4447), .Z(U3573)
         );
  MUX2_X1 U5112 ( .A(n4636), .B(DATAO_REG_20__SCAN_IN), .S(n4447), .Z(U3570)
         );
  MUX2_X1 U5113 ( .A(n4443), .B(DATAO_REG_15__SCAN_IN), .S(n4447), .Z(U3565)
         );
  MUX2_X1 U5114 ( .A(n4444), .B(DATAO_REG_13__SCAN_IN), .S(n4447), .Z(U3563)
         );
  MUX2_X1 U5115 ( .A(n4679), .B(DATAO_REG_11__SCAN_IN), .S(n4447), .Z(U3561)
         );
  MUX2_X1 U5116 ( .A(n4445), .B(DATAO_REG_4__SCAN_IN), .S(n4447), .Z(U3554) );
  MUX2_X1 U5117 ( .A(n4446), .B(DATAO_REG_3__SCAN_IN), .S(n4447), .Z(U3553) );
  MUX2_X1 U5118 ( .A(n3117), .B(DATAO_REG_1__SCAN_IN), .S(n4447), .Z(U3551) );
  OAI22_X1 U5119 ( .A1(n4911), .A2(n4449), .B1(STATE_REG_SCAN_IN), .B2(n4448), 
        .ZN(n4450) );
  AOI21_X1 U5120 ( .B1(n4837), .B2(n4908), .A(n4450), .ZN(n4459) );
  OAI211_X1 U5121 ( .C1(n4453), .C2(n4452), .A(n4923), .B(n4451), .ZN(n4458)
         );
  INV_X1 U5122 ( .A(n4454), .ZN(n4455) );
  OAI21_X1 U5123 ( .B1(n4957), .B2(n2378), .A(n4455), .ZN(n4456) );
  NAND3_X1 U5124 ( .A1(n4921), .A2(n3324), .A3(n4456), .ZN(n4457) );
  NAND3_X1 U5125 ( .A1(n4459), .A2(n4458), .A3(n4457), .ZN(U3241) );
  OAI211_X1 U5126 ( .C1(n4462), .C2(n4461), .A(n4460), .B(n4921), .ZN(n4472)
         );
  INV_X1 U5127 ( .A(n4463), .ZN(n4466) );
  NOR2_X1 U5128 ( .A1(n4926), .A2(n4464), .ZN(n4465) );
  AOI211_X1 U5129 ( .C1(n4914), .C2(ADDR_REG_9__SCAN_IN), .A(n4466), .B(n4465), 
        .ZN(n4471) );
  OAI211_X1 U5130 ( .C1(n4469), .C2(n4468), .A(n4467), .B(n4923), .ZN(n4470)
         );
  NAND3_X1 U5131 ( .A1(n4472), .A2(n4471), .A3(n4470), .ZN(U3249) );
  XOR2_X1 U5132 ( .A(n3751), .B(n4474), .Z(n4478) );
  AOI21_X1 U5133 ( .B1(n4914), .B2(ADDR_REG_16__SCAN_IN), .A(n4475), .ZN(n4476) );
  OAI21_X1 U5134 ( .B1(n4926), .B2(n2371), .A(n4476), .ZN(n4477) );
  AOI21_X1 U5135 ( .B1(n4478), .B2(n4921), .A(n4477), .ZN(n4479) );
  OAI21_X1 U5136 ( .B1(n4480), .B2(n4902), .A(n4479), .ZN(U3256) );
  NAND2_X1 U5137 ( .A1(n4958), .A2(n4786), .ZN(n4482) );
  NAND2_X1 U5138 ( .A1(n4698), .A2(REG2_REG_31__SCAN_IN), .ZN(n4481) );
  OAI211_X1 U5139 ( .C1(n4788), .C2(n4646), .A(n4482), .B(n4481), .ZN(U3260)
         );
  OR2_X1 U5140 ( .A1(n4498), .A2(n4483), .ZN(n4484) );
  INV_X1 U5141 ( .A(n4793), .ZN(n4486) );
  NAND2_X1 U5142 ( .A1(n4486), .A2(n4943), .ZN(n4491) );
  NAND2_X1 U5143 ( .A1(n4937), .A2(n4487), .ZN(n4488) );
  NAND2_X1 U5144 ( .A1(n4489), .A2(n4488), .ZN(n4791) );
  NAND2_X1 U5145 ( .A1(n4958), .A2(n4791), .ZN(n4490) );
  OAI211_X1 U5146 ( .C1(n4958), .C2(n4492), .A(n4491), .B(n4490), .ZN(U3261)
         );
  NAND2_X1 U5147 ( .A1(n4505), .A2(n4495), .ZN(n4720) );
  INV_X1 U5148 ( .A(n4720), .ZN(n4496) );
  NOR2_X1 U5149 ( .A1(n4718), .A2(n4496), .ZN(n4497) );
  XNOR2_X1 U5150 ( .A(n4497), .B(n4716), .ZN(n4519) );
  INV_X1 U5151 ( .A(n4500), .ZN(n4501) );
  AOI21_X1 U5152 ( .B1(n4503), .B2(n4502), .A(n4501), .ZN(n4504) );
  XNOR2_X1 U5153 ( .A(n4504), .B(n4716), .ZN(n4512) );
  NAND2_X1 U5154 ( .A1(n4505), .A2(n4935), .ZN(n4510) );
  AOI22_X1 U5155 ( .A1(n4508), .A2(n4507), .B1(n4937), .B2(n4506), .ZN(n4509)
         );
  OAI21_X1 U5156 ( .B1(n4512), .B2(n4704), .A(n4511), .ZN(n4719) );
  NAND2_X1 U5157 ( .A1(n4698), .A2(REG2_REG_29__SCAN_IN), .ZN(n4517) );
  OAI211_X1 U5158 ( .C1(n4519), .C2(n4649), .A(n4518), .B(n4517), .ZN(U3354)
         );
  INV_X1 U5159 ( .A(n4520), .ZN(n4527) );
  AOI22_X1 U5160 ( .A1(n4521), .A2(n4954), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4698), .ZN(n4522) );
  OAI21_X1 U5161 ( .B1(n4523), .B2(n4646), .A(n4522), .ZN(n4524) );
  AOI21_X1 U5162 ( .B1(n4525), .B2(n4958), .A(n4524), .ZN(n4526) );
  OAI21_X1 U5163 ( .B1(n4527), .B2(n4649), .A(n4526), .ZN(U3262) );
  XNOR2_X1 U5164 ( .A(n4528), .B(n4532), .ZN(n4726) );
  AOI21_X1 U5165 ( .B1(n4535), .B2(n2142), .A(n3215), .ZN(n4724) );
  INV_X1 U5166 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4529) );
  OAI22_X1 U5167 ( .A1(n4530), .A2(n4691), .B1(n4529), .B2(n4958), .ZN(n4531)
         );
  AOI21_X1 U5168 ( .B1(n4724), .B2(n4943), .A(n4531), .ZN(n4540) );
  XNOR2_X1 U5169 ( .A(n4533), .B(n4532), .ZN(n4534) );
  NAND2_X1 U5170 ( .A1(n4534), .A2(n4949), .ZN(n4537) );
  AOI22_X1 U5171 ( .A1(n4566), .A2(n4935), .B1(n4937), .B2(n4535), .ZN(n4536)
         );
  OAI211_X1 U5172 ( .C1(n4538), .C2(n4952), .A(n4537), .B(n4536), .ZN(n4723)
         );
  NAND2_X1 U5173 ( .A1(n4723), .A2(n4958), .ZN(n4539) );
  OAI211_X1 U5174 ( .C1(n4726), .C2(n4649), .A(n4540), .B(n4539), .ZN(U3263)
         );
  XNOR2_X1 U5175 ( .A(n2216), .B(n4544), .ZN(n4728) );
  INV_X1 U5176 ( .A(n4728), .ZN(n4558) );
  INV_X1 U5177 ( .A(n4541), .ZN(n4542) );
  NOR2_X1 U5178 ( .A1(n4543), .A2(n4542), .ZN(n4545) );
  XNOR2_X1 U5179 ( .A(n4545), .B(n4544), .ZN(n4546) );
  NAND2_X1 U5180 ( .A1(n4546), .A2(n4949), .ZN(n4549) );
  AOI22_X1 U5181 ( .A1(n4583), .A2(n4935), .B1(n4547), .B2(n4937), .ZN(n4548)
         );
  OAI211_X1 U5182 ( .C1(n4550), .C2(n4952), .A(n4549), .B(n4548), .ZN(n4727)
         );
  OAI21_X1 U5183 ( .B1(n2276), .B2(n4552), .A(n2142), .ZN(n4798) );
  INV_X1 U5184 ( .A(n4553), .ZN(n4554) );
  AOI22_X1 U5185 ( .A1(n4554), .A2(n4954), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4698), .ZN(n4555) );
  OAI21_X1 U5186 ( .B1(n4798), .B2(n4646), .A(n4555), .ZN(n4556) );
  AOI21_X1 U5187 ( .B1(n4727), .B2(n4958), .A(n4556), .ZN(n4557) );
  OAI21_X1 U5188 ( .B1(n4558), .B2(n4649), .A(n4557), .ZN(U3264) );
  XNOR2_X1 U5189 ( .A(n4559), .B(n4560), .ZN(n4732) );
  INV_X1 U5190 ( .A(n4732), .ZN(n4575) );
  INV_X1 U5191 ( .A(n4560), .ZN(n4561) );
  XNOR2_X1 U5192 ( .A(n4562), .B(n4561), .ZN(n4563) );
  NAND2_X1 U5193 ( .A1(n4563), .A2(n4949), .ZN(n4568) );
  OAI22_X1 U5194 ( .A1(n4564), .A2(n4618), .B1(n4682), .B2(n4570), .ZN(n4565)
         );
  AOI21_X1 U5195 ( .B1(n4566), .B2(n4678), .A(n4565), .ZN(n4567) );
  NAND2_X1 U5196 ( .A1(n4568), .A2(n4567), .ZN(n4731) );
  OAI21_X1 U5197 ( .B1(n4569), .B2(n4570), .A(n4551), .ZN(n4802) );
  AOI22_X1 U5198 ( .A1(n4571), .A2(n4954), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4698), .ZN(n4572) );
  OAI21_X1 U5199 ( .B1(n4802), .B2(n4646), .A(n4572), .ZN(n4573) );
  AOI21_X1 U5200 ( .B1(n4731), .B2(n4958), .A(n4573), .ZN(n4574) );
  OAI21_X1 U5201 ( .B1(n4575), .B2(n4649), .A(n4574), .ZN(U3265) );
  XNOR2_X1 U5202 ( .A(n4576), .B(n4579), .ZN(n4736) );
  INV_X1 U5203 ( .A(n4736), .ZN(n4593) );
  NAND2_X1 U5204 ( .A1(n4578), .A2(n4577), .ZN(n4580) );
  XNOR2_X1 U5205 ( .A(n4580), .B(n4579), .ZN(n4585) );
  OAI22_X1 U5206 ( .A1(n4581), .A2(n4618), .B1(n4589), .B2(n4682), .ZN(n4582)
         );
  AOI21_X1 U5207 ( .B1(n4583), .B2(n4678), .A(n4582), .ZN(n4584) );
  OAI21_X1 U5208 ( .B1(n4585), .B2(n4704), .A(n4584), .ZN(n4735) );
  INV_X1 U5209 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4586) );
  OAI22_X1 U5210 ( .A1(n4587), .A2(n4691), .B1(n4586), .B2(n4958), .ZN(n4591)
         );
  INV_X1 U5211 ( .A(n4569), .ZN(n4588) );
  OAI21_X1 U5212 ( .B1(n2278), .B2(n4589), .A(n4588), .ZN(n4806) );
  NOR2_X1 U5213 ( .A1(n4806), .A2(n4646), .ZN(n4590) );
  AOI211_X1 U5214 ( .C1(n4958), .C2(n4735), .A(n4591), .B(n4590), .ZN(n4592)
         );
  OAI21_X1 U5215 ( .B1(n4593), .B2(n4649), .A(n4592), .ZN(U3266) );
  XOR2_X1 U5216 ( .A(n4594), .B(n4599), .Z(n4740) );
  INV_X1 U5217 ( .A(n4740), .ZN(n4614) );
  NOR2_X1 U5218 ( .A1(n4595), .A2(n4620), .ZN(n4619) );
  INV_X1 U5219 ( .A(n4596), .ZN(n4597) );
  NOR2_X1 U5220 ( .A1(n4619), .A2(n4597), .ZN(n4598) );
  XOR2_X1 U5221 ( .A(n4599), .B(n4598), .Z(n4605) );
  OAI22_X1 U5222 ( .A1(n4601), .A2(n4618), .B1(n4682), .B2(n4600), .ZN(n4602)
         );
  AOI21_X1 U5223 ( .B1(n4603), .B2(n4678), .A(n4602), .ZN(n4604) );
  OAI21_X1 U5224 ( .B1(n4605), .B2(n4704), .A(n4604), .ZN(n4739) );
  NAND2_X1 U5225 ( .A1(n4744), .A2(n4606), .ZN(n4607) );
  NAND2_X1 U5226 ( .A1(n4608), .A2(n4607), .ZN(n4810) );
  INV_X1 U5227 ( .A(n4609), .ZN(n4610) );
  AOI22_X1 U5228 ( .A1(n4610), .A2(n4954), .B1(REG2_REG_23__SCAN_IN), .B2(
        n4698), .ZN(n4611) );
  OAI21_X1 U5229 ( .B1(n4810), .B2(n4646), .A(n4611), .ZN(n4612) );
  AOI21_X1 U5230 ( .B1(n4739), .B2(n4958), .A(n4612), .ZN(n4613) );
  OAI21_X1 U5231 ( .B1(n4614), .B2(n4649), .A(n4613), .ZN(U3267) );
  OAI21_X1 U5232 ( .B1(n4616), .B2(n4620), .A(n4615), .ZN(n4747) );
  OAI22_X1 U5233 ( .A1(n4657), .A2(n4618), .B1(n4617), .B2(n4682), .ZN(n4623)
         );
  AOI21_X1 U5234 ( .B1(n4620), .B2(n4595), .A(n4619), .ZN(n4621) );
  NOR2_X1 U5235 ( .A1(n4621), .A2(n4704), .ZN(n4622) );
  AOI211_X1 U5236 ( .C1(n4678), .C2(n4624), .A(n4623), .B(n4622), .ZN(n4746)
         );
  INV_X1 U5237 ( .A(n4746), .ZN(n4630) );
  NAND2_X1 U5238 ( .A1(n4625), .A2(n3155), .ZN(n4743) );
  AND3_X1 U5239 ( .A1(n4744), .A2(n4943), .A3(n4743), .ZN(n4629) );
  INV_X1 U5240 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4626) );
  OAI22_X1 U5241 ( .A1(n4627), .A2(n4691), .B1(n4626), .B2(n4958), .ZN(n4628)
         );
  AOI211_X1 U5242 ( .C1(n4630), .C2(n4958), .A(n4629), .B(n4628), .ZN(n4631)
         );
  OAI21_X1 U5243 ( .B1(n4649), .B2(n4747), .A(n4631), .ZN(U3268) );
  XOR2_X1 U5244 ( .A(n4633), .B(n4632), .Z(n4749) );
  INV_X1 U5245 ( .A(n4749), .ZN(n4650) );
  XNOR2_X1 U5246 ( .A(n4634), .B(n4633), .ZN(n4635) );
  NAND2_X1 U5247 ( .A1(n4635), .A2(n4949), .ZN(n4641) );
  NAND2_X1 U5248 ( .A1(n4636), .A2(n4935), .ZN(n4637) );
  OAI21_X1 U5249 ( .B1(n4682), .B2(n4643), .A(n4637), .ZN(n4638) );
  AOI21_X1 U5250 ( .B1(n4639), .B2(n4678), .A(n4638), .ZN(n4640) );
  NAND2_X1 U5251 ( .A1(n4641), .A2(n4640), .ZN(n4748) );
  OAI21_X1 U5252 ( .B1(n4642), .B2(n4643), .A(n4625), .ZN(n4815) );
  AOI22_X1 U5253 ( .A1(n4698), .A2(REG2_REG_21__SCAN_IN), .B1(n4644), .B2(
        n4954), .ZN(n4645) );
  OAI21_X1 U5254 ( .B1(n4815), .B2(n4646), .A(n4645), .ZN(n4647) );
  AOI21_X1 U5255 ( .B1(n4748), .B2(n4958), .A(n4647), .ZN(n4648) );
  OAI21_X1 U5256 ( .B1(n4650), .B2(n4649), .A(n4648), .ZN(U3269) );
  INV_X1 U5257 ( .A(n4651), .ZN(n4652) );
  NAND2_X1 U5258 ( .A1(n4653), .A2(n4652), .ZN(n4654) );
  XNOR2_X1 U5259 ( .A(n4654), .B(n4662), .ZN(n4666) );
  AOI22_X1 U5260 ( .A1(n4655), .A2(n4935), .B1(n4667), .B2(n4937), .ZN(n4656)
         );
  OAI21_X1 U5261 ( .B1(n4657), .B2(n4952), .A(n4656), .ZN(n4665) );
  NAND2_X1 U5262 ( .A1(n4659), .A2(n4658), .ZN(n4661) );
  NAND2_X1 U5263 ( .A1(n4661), .A2(n4660), .ZN(n4663) );
  XNOR2_X1 U5264 ( .A(n4663), .B(n4662), .ZN(n4756) );
  NOR2_X1 U5265 ( .A1(n4756), .A2(n4699), .ZN(n4664) );
  AOI211_X1 U5266 ( .C1(n4949), .C2(n4666), .A(n4665), .B(n4664), .ZN(n4755)
         );
  INV_X1 U5267 ( .A(n4756), .ZN(n4672) );
  INV_X1 U5268 ( .A(n4642), .ZN(n4753) );
  NAND2_X1 U5269 ( .A1(n2150), .A2(n4667), .ZN(n4752) );
  AND3_X1 U5270 ( .A1(n4753), .A2(n4943), .A3(n4752), .ZN(n4671) );
  OAI22_X1 U5271 ( .A1(n4958), .A2(n4669), .B1(n4668), .B2(n4691), .ZN(n4670)
         );
  AOI211_X1 U5272 ( .C1(n4672), .C2(n4955), .A(n4671), .B(n4670), .ZN(n4673)
         );
  OAI21_X1 U5273 ( .B1(n4755), .B2(n4698), .A(n4673), .ZN(U3270) );
  OR2_X1 U5274 ( .A1(n4675), .A2(n4674), .ZN(n4677) );
  XOR2_X1 U5275 ( .A(n2175), .B(n4685), .Z(n4688) );
  AOI22_X1 U5276 ( .A1(n4935), .A2(n4680), .B1(n4679), .B2(n4678), .ZN(n4681)
         );
  OAI21_X1 U5277 ( .B1(n4683), .B2(n4682), .A(n4681), .ZN(n4687) );
  XNOR2_X1 U5278 ( .A(n4684), .B(n4685), .ZN(n4783) );
  NOR2_X1 U5279 ( .A1(n4783), .A2(n4699), .ZN(n4686) );
  AOI211_X1 U5280 ( .C1(n4688), .C2(n4949), .A(n4687), .B(n4686), .ZN(n4782)
         );
  INV_X1 U5281 ( .A(n4783), .ZN(n4696) );
  NAND2_X1 U5282 ( .A1(n4690), .A2(n4689), .ZN(n4780) );
  AND3_X1 U5283 ( .A1(n2149), .A2(n4943), .A3(n4780), .ZN(n4695) );
  OAI22_X1 U5284 ( .A1(n4958), .A2(n4693), .B1(n4692), .B2(n4691), .ZN(n4694)
         );
  AOI211_X1 U5285 ( .C1(n4696), .C2(n4955), .A(n4695), .B(n4694), .ZN(n4697)
         );
  OAI21_X1 U5286 ( .B1(n4782), .B2(n4698), .A(n4697), .ZN(U3280) );
  INV_X1 U5287 ( .A(n4699), .ZN(n4950) );
  OAI21_X1 U5288 ( .B1(n4701), .B2(n4703), .A(n4700), .ZN(n4992) );
  AOI22_X1 U5289 ( .A1(n4710), .A2(n4937), .B1(n3117), .B2(n4935), .ZN(n4702)
         );
  OAI21_X1 U5290 ( .B1(n3121), .B2(n4952), .A(n4702), .ZN(n4707) );
  NAND3_X1 U5291 ( .A1(n4931), .A2(n4703), .A3(n3164), .ZN(n4705) );
  AOI21_X1 U5292 ( .B1(n3560), .B2(n4705), .A(n4704), .ZN(n4706) );
  AOI211_X1 U5293 ( .C1(n4950), .C2(n4992), .A(n4707), .B(n4706), .ZN(n4995)
         );
  MUX2_X1 U5294 ( .A(n4708), .B(n4995), .S(n4958), .Z(n4713) );
  AOI22_X1 U5295 ( .A1(n4955), .A2(n4992), .B1(REG3_REG_2__SCAN_IN), .B2(n4954), .ZN(n4712) );
  NAND2_X1 U5296 ( .A1(n4709), .A2(n4710), .ZN(n4993) );
  NAND3_X1 U5297 ( .A1(n4943), .A2(n3567), .A3(n4993), .ZN(n4711) );
  NAND3_X1 U5298 ( .A1(n4713), .A2(n4712), .A3(n4711), .ZN(U3288) );
  NAND2_X1 U5299 ( .A1(n5030), .A2(n4791), .ZN(n4715) );
  NAND2_X1 U5300 ( .A1(n3224), .A2(REG1_REG_30__SCAN_IN), .ZN(n4714) );
  OAI211_X1 U5301 ( .C1(n4793), .C2(n4761), .A(n4715), .B(n4714), .ZN(U3548)
         );
  INV_X1 U5302 ( .A(n4716), .ZN(n4721) );
  NAND3_X1 U5303 ( .A1(n4720), .A2(n5017), .A3(n4721), .ZN(n4717) );
  AOI21_X1 U5304 ( .B1(n2138), .B2(n4724), .A(n4723), .ZN(n4725) );
  OAI21_X1 U5305 ( .B1(n4726), .B2(n5009), .A(n4725), .ZN(n4794) );
  MUX2_X1 U5306 ( .A(REG1_REG_27__SCAN_IN), .B(n4794), .S(n5030), .Z(U3545) );
  AOI21_X1 U5307 ( .B1(n4728), .B2(n5017), .A(n4727), .ZN(n4795) );
  MUX2_X1 U5308 ( .A(n4729), .B(n4795), .S(n5030), .Z(n4730) );
  OAI21_X1 U5309 ( .B1(n4761), .B2(n4798), .A(n4730), .ZN(U3544) );
  AOI21_X1 U5310 ( .B1(n4732), .B2(n5017), .A(n4731), .ZN(n4799) );
  MUX2_X1 U5311 ( .A(n4733), .B(n4799), .S(n5030), .Z(n4734) );
  OAI21_X1 U5312 ( .B1(n4761), .B2(n4802), .A(n4734), .ZN(U3543) );
  AOI21_X1 U5313 ( .B1(n4736), .B2(n5017), .A(n4735), .ZN(n4803) );
  MUX2_X1 U5314 ( .A(n4737), .B(n4803), .S(n5030), .Z(n4738) );
  OAI21_X1 U5315 ( .B1(n4761), .B2(n4806), .A(n4738), .ZN(U3542) );
  AOI21_X1 U5316 ( .B1(n4740), .B2(n5017), .A(n4739), .ZN(n4807) );
  MUX2_X1 U5317 ( .A(n4741), .B(n4807), .S(n5030), .Z(n4742) );
  OAI21_X1 U5318 ( .B1(n4761), .B2(n4810), .A(n4742), .ZN(U3541) );
  NAND3_X1 U5319 ( .A1(n4744), .A2(n2138), .A3(n4743), .ZN(n4745) );
  OAI211_X1 U5320 ( .C1(n5009), .C2(n4747), .A(n4746), .B(n4745), .ZN(n4811)
         );
  MUX2_X1 U5321 ( .A(REG1_REG_22__SCAN_IN), .B(n4811), .S(n5030), .Z(U3540) );
  AOI21_X1 U5322 ( .B1(n4749), .B2(n5017), .A(n4748), .ZN(n4812) );
  MUX2_X1 U5323 ( .A(n4750), .B(n4812), .S(n5030), .Z(n4751) );
  OAI21_X1 U5324 ( .B1(n4761), .B2(n4815), .A(n4751), .ZN(U3539) );
  NAND3_X1 U5325 ( .A1(n4753), .A2(n2138), .A3(n4752), .ZN(n4754) );
  OAI211_X1 U5326 ( .C1(n4756), .C2(n4998), .A(n4755), .B(n4754), .ZN(n4816)
         );
  MUX2_X1 U5327 ( .A(REG1_REG_20__SCAN_IN), .B(n4816), .S(n5030), .Z(U3538) );
  INV_X1 U5328 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4759) );
  AOI21_X1 U5329 ( .B1(n4758), .B2(n5017), .A(n4757), .ZN(n4817) );
  MUX2_X1 U5330 ( .A(n4759), .B(n4817), .S(n5030), .Z(n4760) );
  OAI21_X1 U5331 ( .B1(n4761), .B2(n4821), .A(n4760), .ZN(U3537) );
  OAI211_X1 U5332 ( .C1(n4764), .C2(n5009), .A(n4763), .B(n4762), .ZN(n4822)
         );
  MUX2_X1 U5333 ( .A(REG1_REG_18__SCAN_IN), .B(n4822), .S(n5030), .Z(U3536) );
  OR3_X1 U5334 ( .A1(n4766), .A2(n4765), .A3(n4779), .ZN(n4767) );
  OAI211_X1 U5335 ( .C1(n4769), .C2(n5009), .A(n4768), .B(n4767), .ZN(n4823)
         );
  MUX2_X1 U5336 ( .A(REG1_REG_16__SCAN_IN), .B(n4823), .S(n5030), .Z(U3534) );
  NAND3_X1 U5337 ( .A1(n4771), .A2(n2138), .A3(n4770), .ZN(n4772) );
  OAI211_X1 U5338 ( .C1(n4774), .C2(n4998), .A(n4773), .B(n4772), .ZN(n4824)
         );
  MUX2_X1 U5339 ( .A(REG1_REG_14__SCAN_IN), .B(n4824), .S(n5030), .Z(U3532) );
  NAND2_X1 U5340 ( .A1(n4775), .A2(n5017), .ZN(n4776) );
  OAI211_X1 U5341 ( .C1(n4779), .C2(n4778), .A(n4777), .B(n4776), .ZN(n4825)
         );
  MUX2_X1 U5342 ( .A(REG1_REG_11__SCAN_IN), .B(n4825), .S(n5030), .Z(U3529) );
  NAND3_X1 U5343 ( .A1(n2149), .A2(n2138), .A3(n4780), .ZN(n4781) );
  OAI211_X1 U5344 ( .C1(n4783), .C2(n4998), .A(n4782), .B(n4781), .ZN(n4826)
         );
  MUX2_X1 U5345 ( .A(REG1_REG_10__SCAN_IN), .B(n4826), .S(n5030), .Z(U3528) );
  NOR2_X1 U5346 ( .A1(n5020), .A2(n4784), .ZN(n4785) );
  AOI21_X1 U5347 ( .B1(n5020), .B2(n4786), .A(n4785), .ZN(n4787) );
  OAI21_X1 U5348 ( .B1(n4788), .B2(n4820), .A(n4787), .ZN(U3517) );
  NOR2_X1 U5349 ( .A1(n5020), .A2(n4789), .ZN(n4790) );
  AOI21_X1 U5350 ( .B1(n5020), .B2(n4791), .A(n4790), .ZN(n4792) );
  OAI21_X1 U5351 ( .B1(n4793), .B2(n4820), .A(n4792), .ZN(U3516) );
  MUX2_X1 U5352 ( .A(REG0_REG_27__SCAN_IN), .B(n4794), .S(n5020), .Z(U3513) );
  INV_X1 U5353 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4796) );
  MUX2_X1 U5354 ( .A(n4796), .B(n4795), .S(n5020), .Z(n4797) );
  OAI21_X1 U5355 ( .B1(n4798), .B2(n4820), .A(n4797), .ZN(U3512) );
  INV_X1 U5356 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4800) );
  MUX2_X1 U5357 ( .A(n4800), .B(n4799), .S(n5020), .Z(n4801) );
  OAI21_X1 U5358 ( .B1(n4802), .B2(n4820), .A(n4801), .ZN(U3511) );
  INV_X1 U5359 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4804) );
  MUX2_X1 U5360 ( .A(n4804), .B(n4803), .S(n5020), .Z(n4805) );
  OAI21_X1 U5361 ( .B1(n4806), .B2(n4820), .A(n4805), .ZN(U3510) );
  INV_X1 U5362 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4808) );
  MUX2_X1 U5363 ( .A(n4808), .B(n4807), .S(n5020), .Z(n4809) );
  OAI21_X1 U5364 ( .B1(n4810), .B2(n4820), .A(n4809), .ZN(U3509) );
  MUX2_X1 U5365 ( .A(REG0_REG_22__SCAN_IN), .B(n4811), .S(n5020), .Z(U3508) );
  MUX2_X1 U5366 ( .A(n4813), .B(n4812), .S(n5020), .Z(n4814) );
  OAI21_X1 U5367 ( .B1(n4815), .B2(n4820), .A(n4814), .ZN(U3507) );
  MUX2_X1 U5368 ( .A(REG0_REG_20__SCAN_IN), .B(n4816), .S(n5020), .Z(U3506) );
  MUX2_X1 U5369 ( .A(n4818), .B(n4817), .S(n5020), .Z(n4819) );
  OAI21_X1 U5370 ( .B1(n4821), .B2(n4820), .A(n4819), .ZN(U3505) );
  MUX2_X1 U5371 ( .A(REG0_REG_18__SCAN_IN), .B(n4822), .S(n5020), .Z(U3503) );
  MUX2_X1 U5372 ( .A(REG0_REG_16__SCAN_IN), .B(n4823), .S(n5020), .Z(U3499) );
  MUX2_X1 U5373 ( .A(REG0_REG_14__SCAN_IN), .B(n4824), .S(n5020), .Z(U3495) );
  MUX2_X1 U5374 ( .A(REG0_REG_11__SCAN_IN), .B(n4825), .S(n5020), .Z(U3489) );
  MUX2_X1 U5375 ( .A(REG0_REG_10__SCAN_IN), .B(n4826), .S(n5020), .Z(U3487) );
  MUX2_X1 U5376 ( .A(DATAI_29_), .B(n4827), .S(STATE_REG_SCAN_IN), .Z(U3323)
         );
  MUX2_X1 U5377 ( .A(n3047), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5378 ( .A(n4828), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5379 ( .A(n4829), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5380 ( .A(DATAI_16_), .B(n4830), .S(STATE_REG_SCAN_IN), .Z(U3336)
         );
  MUX2_X1 U5381 ( .A(DATAI_15_), .B(n4907), .S(STATE_REG_SCAN_IN), .Z(U3337)
         );
  MUX2_X1 U5382 ( .A(n4831), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5383 ( .A(DATAI_8_), .B(n4832), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5384 ( .A(n4833), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5385 ( .A(n4834), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5386 ( .A(DATAI_3_), .B(n4835), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5387 ( .A(n4836), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5388 ( .A(n4837), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5389 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  AOI22_X1 U5390 ( .A1(STATE_REG_SCAN_IN), .A2(n4838), .B1(n3036), .B2(U3149), 
        .ZN(U3324) );
  INV_X1 U5391 ( .A(REG2_REG_4__SCAN_IN), .ZN(n4840) );
  XNOR2_X1 U5392 ( .A(n4839), .B(n4840), .ZN(n4841) );
  NAND2_X1 U5393 ( .A1(n4921), .A2(n4841), .ZN(n4850) );
  XNOR2_X1 U5394 ( .A(n4843), .B(n4842), .ZN(n4844) );
  NAND2_X1 U5395 ( .A1(n4923), .A2(n4844), .ZN(n4849) );
  NAND2_X1 U5396 ( .A1(n4908), .A2(n4845), .ZN(n4848) );
  AOI21_X1 U5397 ( .B1(n4914), .B2(ADDR_REG_4__SCAN_IN), .A(n4846), .ZN(n4847)
         );
  AND4_X1 U5398 ( .A1(n4850), .A2(n4849), .A3(n4848), .A4(n4847), .ZN(n4852)
         );
  NAND2_X1 U5399 ( .A1(n4852), .A2(n4851), .ZN(U3244) );
  AOI211_X1 U5400 ( .C1(n4855), .C2(n4854), .A(n4853), .B(n4902), .ZN(n4856)
         );
  AOI211_X1 U5401 ( .C1(n4914), .C2(ADDR_REG_10__SCAN_IN), .A(n4857), .B(n4856), .ZN(n4861) );
  OAI211_X1 U5402 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4859), .A(n4921), .B(n4858), .ZN(n4860) );
  OAI211_X1 U5403 ( .C1(n4926), .C2(n4983), .A(n4861), .B(n4860), .ZN(U3250)
         );
  AOI211_X1 U5404 ( .C1(n4864), .C2(n4863), .A(n4862), .B(n4902), .ZN(n4865)
         );
  AOI211_X1 U5405 ( .C1(n4914), .C2(ADDR_REG_12__SCAN_IN), .A(n4866), .B(n4865), .ZN(n4870) );
  OAI211_X1 U5406 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4868), .A(n4921), .B(n4867), .ZN(n4869) );
  OAI211_X1 U5407 ( .C1(n4926), .C2(n4981), .A(n4870), .B(n4869), .ZN(U3252)
         );
  AOI211_X1 U5408 ( .C1(n4873), .C2(n4872), .A(n4871), .B(n4902), .ZN(n4874)
         );
  AOI211_X1 U5409 ( .C1(ADDR_REG_13__SCAN_IN), .C2(n4914), .A(n4875), .B(n4874), .ZN(n4882) );
  AOI21_X1 U5410 ( .B1(n4980), .B2(n4877), .A(n4876), .ZN(n4880) );
  AOI21_X1 U5411 ( .B1(n4880), .B2(n4879), .A(n4896), .ZN(n4878) );
  OAI21_X1 U5412 ( .B1(n4880), .B2(n4879), .A(n4878), .ZN(n4881) );
  OAI211_X1 U5413 ( .C1(n4926), .C2(n4980), .A(n4882), .B(n4881), .ZN(U3253)
         );
  NOR2_X1 U5414 ( .A1(n4884), .A2(n4883), .ZN(n4899) );
  AOI211_X1 U5415 ( .C1(n4884), .C2(n4883), .A(n4899), .B(n4902), .ZN(n4889)
         );
  AOI211_X1 U5416 ( .C1(n4887), .C2(n4886), .A(n4885), .B(n4896), .ZN(n4888)
         );
  AOI211_X1 U5417 ( .C1(n4908), .C2(n4890), .A(n4889), .B(n4888), .ZN(n4892)
         );
  OAI211_X1 U5418 ( .C1(n4893), .C2(n4911), .A(n4892), .B(n4891), .ZN(U3254)
         );
  INV_X1 U5419 ( .A(n4894), .ZN(n4895) );
  AOI211_X1 U5420 ( .C1(n4898), .C2(n4897), .A(n4896), .B(n4895), .ZN(n4906)
         );
  NOR2_X1 U5421 ( .A1(n4900), .A2(n4899), .ZN(n4904) );
  NOR2_X1 U5422 ( .A1(n4904), .A2(n4903), .ZN(n4901) );
  AOI211_X1 U5423 ( .C1(n4904), .C2(n4903), .A(n4902), .B(n4901), .ZN(n4905)
         );
  AOI211_X1 U5424 ( .C1(n4908), .C2(n4907), .A(n4906), .B(n4905), .ZN(n4910)
         );
  OAI211_X1 U5425 ( .C1(n4912), .C2(n4911), .A(n4910), .B(n4909), .ZN(U3255)
         );
  AOI21_X1 U5426 ( .B1(n4914), .B2(ADDR_REG_17__SCAN_IN), .A(n4913), .ZN(n4925) );
  OAI21_X1 U5427 ( .B1(n4916), .B2(n4915), .A(n2592), .ZN(n4922) );
  OAI21_X1 U5428 ( .B1(n4919), .B2(n4918), .A(n4917), .ZN(n4920) );
  AOI22_X1 U5429 ( .A1(n4923), .A2(n4922), .B1(n4921), .B2(n4920), .ZN(n4924)
         );
  OAI211_X1 U5430 ( .C1(n4976), .C2(n4926), .A(n4925), .B(n4924), .ZN(U3257)
         );
  OAI21_X1 U5431 ( .B1(n4929), .B2(n4928), .A(n4927), .ZN(n4930) );
  INV_X1 U5432 ( .A(n4930), .ZN(n4989) );
  OAI21_X1 U5433 ( .B1(n4933), .B2(n4932), .A(n4931), .ZN(n4934) );
  NAND2_X1 U5434 ( .A1(n4934), .A2(n4949), .ZN(n4939) );
  AOI22_X1 U5435 ( .A1(n3115), .A2(n4937), .B1(n4936), .B2(n4935), .ZN(n4938)
         );
  OAI211_X1 U5436 ( .C1(n4940), .C2(n4952), .A(n4939), .B(n4938), .ZN(n4941)
         );
  AOI21_X1 U5437 ( .B1(n4950), .B2(n4989), .A(n4941), .ZN(n4991) );
  AOI22_X1 U5438 ( .A1(REG2_REG_1__SCAN_IN), .A2(n4698), .B1(
        REG3_REG_1__SCAN_IN), .B2(n4954), .ZN(n4945) );
  AOI21_X1 U5439 ( .B1(n3115), .B2(n4942), .A(n3099), .ZN(n4988) );
  AOI22_X1 U5440 ( .A1(n4943), .A2(n4988), .B1(n4955), .B2(n4989), .ZN(n4944)
         );
  OAI211_X1 U5441 ( .C1(n4698), .C2(n4991), .A(n4945), .B(n4944), .ZN(U3289)
         );
  NOR2_X1 U5442 ( .A1(n4947), .A2(n4946), .ZN(n4985) );
  INV_X1 U5443 ( .A(n4948), .ZN(n4986) );
  OAI21_X1 U5444 ( .B1(n4950), .B2(n4949), .A(n4986), .ZN(n4951) );
  OAI21_X1 U5445 ( .B1(n3116), .B2(n4952), .A(n4951), .ZN(n4984) );
  AOI21_X1 U5446 ( .B1(n4985), .B2(n4953), .A(n4984), .ZN(n4959) );
  AOI22_X1 U5447 ( .A1(n4955), .A2(n4986), .B1(REG3_REG_0__SCAN_IN), .B2(n4954), .ZN(n4956) );
  OAI221_X1 U5448 ( .B1(n4698), .B2(n4959), .C1(n4958), .C2(n4957), .A(n4956), 
        .ZN(U3290) );
  NOR2_X1 U5449 ( .A1(n4973), .A2(n4960), .ZN(U3291) );
  NOR2_X1 U5450 ( .A1(n4973), .A2(n4961), .ZN(U3292) );
  AND2_X1 U5451 ( .A1(D_REG_29__SCAN_IN), .A2(n4974), .ZN(U3293) );
  AND2_X1 U5452 ( .A1(D_REG_28__SCAN_IN), .A2(n4974), .ZN(U3294) );
  NOR2_X1 U5453 ( .A1(n4973), .A2(n4962), .ZN(U3295) );
  NOR2_X1 U5454 ( .A1(n4973), .A2(n4963), .ZN(U3296) );
  NOR2_X1 U5455 ( .A1(n4973), .A2(n4964), .ZN(U3297) );
  AND2_X1 U5456 ( .A1(D_REG_24__SCAN_IN), .A2(n4974), .ZN(U3298) );
  NOR2_X1 U5457 ( .A1(n4973), .A2(n4965), .ZN(U3299) );
  AND2_X1 U5458 ( .A1(D_REG_22__SCAN_IN), .A2(n4974), .ZN(U3300) );
  NOR2_X1 U5459 ( .A1(n4973), .A2(n4966), .ZN(U3301) );
  AND2_X1 U5460 ( .A1(D_REG_20__SCAN_IN), .A2(n4974), .ZN(U3302) );
  AND2_X1 U5461 ( .A1(D_REG_19__SCAN_IN), .A2(n4974), .ZN(U3303) );
  AND2_X1 U5462 ( .A1(D_REG_18__SCAN_IN), .A2(n4974), .ZN(U3304) );
  AND2_X1 U5463 ( .A1(D_REG_17__SCAN_IN), .A2(n4974), .ZN(U3305) );
  AND2_X1 U5464 ( .A1(D_REG_16__SCAN_IN), .A2(n4974), .ZN(U3306) );
  AND2_X1 U5465 ( .A1(D_REG_15__SCAN_IN), .A2(n4974), .ZN(U3307) );
  NOR2_X1 U5466 ( .A1(n4973), .A2(n4967), .ZN(U3308) );
  AND2_X1 U5467 ( .A1(D_REG_13__SCAN_IN), .A2(n4974), .ZN(U3309) );
  AND2_X1 U5468 ( .A1(D_REG_12__SCAN_IN), .A2(n4974), .ZN(U3310) );
  AND2_X1 U5469 ( .A1(D_REG_11__SCAN_IN), .A2(n4974), .ZN(U3311) );
  NOR2_X1 U5470 ( .A1(n4973), .A2(n4968), .ZN(U3312) );
  NOR2_X1 U5471 ( .A1(n4973), .A2(n4969), .ZN(U3313) );
  NOR2_X1 U5472 ( .A1(n4973), .A2(n4970), .ZN(U3314) );
  AND2_X1 U5473 ( .A1(D_REG_7__SCAN_IN), .A2(n4974), .ZN(U3315) );
  AND2_X1 U5474 ( .A1(D_REG_6__SCAN_IN), .A2(n4974), .ZN(U3316) );
  NOR2_X1 U5475 ( .A1(n4973), .A2(n4971), .ZN(U3317) );
  AND2_X1 U5476 ( .A1(D_REG_4__SCAN_IN), .A2(n4974), .ZN(U3318) );
  NOR2_X1 U5477 ( .A1(n4973), .A2(n4972), .ZN(U3319) );
  AND2_X1 U5478 ( .A1(D_REG_2__SCAN_IN), .A2(n4974), .ZN(U3320) );
  AOI21_X1 U5479 ( .B1(U3149), .B2(n2961), .A(n4975), .ZN(U3329) );
  AOI22_X1 U5480 ( .A1(STATE_REG_SCAN_IN), .A2(n4976), .B1(n2883), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5481 ( .A(DATAI_14_), .ZN(n4977) );
  AOI22_X1 U5482 ( .A1(STATE_REG_SCAN_IN), .A2(n4978), .B1(n4977), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5483 ( .A1(STATE_REG_SCAN_IN), .A2(n4980), .B1(n4979), .B2(U3149), 
        .ZN(U3339) );
  AOI22_X1 U5484 ( .A1(STATE_REG_SCAN_IN), .A2(n4981), .B1(n2806), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5485 ( .A1(STATE_REG_SCAN_IN), .A2(n4983), .B1(n4982), .B2(U3149), 
        .ZN(U3342) );
  AOI211_X1 U5486 ( .C1(n5007), .C2(n4986), .A(n4985), .B(n4984), .ZN(n5022)
         );
  INV_X1 U5487 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4987) );
  AOI22_X1 U5488 ( .A1(n5020), .A2(n5022), .B1(n4987), .B2(n5019), .ZN(U3467)
         );
  AOI22_X1 U5489 ( .A1(n4989), .A2(n5007), .B1(n4988), .B2(n2138), .ZN(n4990)
         );
  AND2_X1 U5490 ( .A1(n4991), .A2(n4990), .ZN(n5023) );
  AOI22_X1 U5491 ( .A1(n5020), .A2(n5023), .B1(n3955), .B2(n5019), .ZN(U3469)
         );
  INV_X1 U5492 ( .A(n4992), .ZN(n4996) );
  NAND3_X1 U5493 ( .A1(n3567), .A2(n2138), .A3(n4993), .ZN(n4994) );
  OAI211_X1 U5494 ( .C1(n4996), .C2(n4998), .A(n4995), .B(n4994), .ZN(n4997)
         );
  INV_X1 U5495 ( .A(n4997), .ZN(n5024) );
  AOI22_X1 U5496 ( .A1(n5020), .A2(n5024), .B1(n2628), .B2(n5019), .ZN(U3471)
         );
  NOR2_X1 U5497 ( .A1(n4999), .A2(n4998), .ZN(n5001) );
  AOI211_X1 U5498 ( .C1(n2138), .C2(n5002), .A(n5001), .B(n5000), .ZN(n5025)
         );
  INV_X1 U5499 ( .A(REG0_REG_3__SCAN_IN), .ZN(n5003) );
  AOI22_X1 U5500 ( .A1(n5020), .A2(n5025), .B1(n5003), .B2(n5019), .ZN(U3473)
         );
  INV_X1 U5501 ( .A(n5004), .ZN(n5006) );
  AOI211_X1 U5502 ( .C1(n5008), .C2(n5007), .A(n5006), .B(n5005), .ZN(n5026)
         );
  AOI22_X1 U5503 ( .A1(n5020), .A2(n5026), .B1(n2682), .B2(n5019), .ZN(U3475)
         );
  NOR2_X1 U5504 ( .A1(n5010), .A2(n5009), .ZN(n5013) );
  INV_X1 U5505 ( .A(n5011), .ZN(n5012) );
  AOI211_X1 U5506 ( .C1(n2138), .C2(n5014), .A(n5013), .B(n5012), .ZN(n5028)
         );
  AOI22_X1 U5507 ( .A1(n5020), .A2(n5028), .B1(n2698), .B2(n5019), .ZN(U3477)
         );
  AOI211_X1 U5508 ( .C1(n5018), .C2(n5017), .A(n5016), .B(n5015), .ZN(n5029)
         );
  AOI22_X1 U5509 ( .A1(n5020), .A2(n5029), .B1(n2727), .B2(n5019), .ZN(U3481)
         );
  AOI22_X1 U5510 ( .A1(n5030), .A2(n5022), .B1(n5021), .B2(n3224), .ZN(U3518)
         );
  AOI22_X1 U5511 ( .A1(n5030), .A2(n5023), .B1(n2646), .B2(n3224), .ZN(U3519)
         );
  AOI22_X1 U5512 ( .A1(n5030), .A2(n5024), .B1(n2627), .B2(n3224), .ZN(U3520)
         );
  AOI22_X1 U5513 ( .A1(n5030), .A2(n5025), .B1(n2673), .B2(n3224), .ZN(U3521)
         );
  AOI22_X1 U5514 ( .A1(n5030), .A2(n5026), .B1(n4842), .B2(n3224), .ZN(U3522)
         );
  AOI22_X1 U5515 ( .A1(n5030), .A2(n5028), .B1(n5027), .B2(n3224), .ZN(U3523)
         );
  AOI22_X1 U5516 ( .A1(n5030), .A2(n5029), .B1(n2564), .B2(n3224), .ZN(U3525)
         );
  NAND4_X1 U2387 ( .A1(n2747), .A2(n2746), .A3(n2745), .A4(n2744), .ZN(n3629)
         );
  CLKBUF_X1 U2393 ( .A(n3109), .Z(n2138) );
endmodule

